/* Verilog module written by vlog2Verilog (qflow) */

module array16(
    input [15:0] a,
    input [15:0] b,
    output [31:0] c
);

wire vdd = 1'b1;
wire gnd = 1'b0;

wire \z4.z1.z2.z1.a  ;
wire [15:0] a ;
wire [15:0] b ;
wire [31:0] c ;
wire _1677_ ;
wire _1257_ ;
wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire \z1.z4.z1.z2.c  ;
wire _397_ ;
wire \z1.z1.z1.z1.c  ;
wire _2903_ ;
wire _1295_ ;
wire _3021_ ;
wire _2712_ ;
wire \z1.z4.z2.z1.s  ;
wire \z3.z1.z4.z1.b  ;
wire _2941_ ;
wire _2521_ ;
wire _2101_ ;
wire \z1.z2.z4.z2.s  ;
wire \z4.z4.z3.z1.s  ;
wire _703_ ;
wire \z2.z4.z1.z1.a  ;
wire _1389_ ;
wire _2750_ ;
wire _2330_ ;
wire _19_ ;
wire _1601_ ;
wire \z2.z2.z3.z2.a  ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire \z3.z2.z1.z1.c  ;
wire _1198_ ;
wire _1830_ ;
wire _1410_ ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _57_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _2844_ ;
wire _2424_ ;
wire _2004_ ;
wire \z1.z4.z3.z1.b  ;
wire _606_ ;
wire _2653_ ;
wire _2233_ ;
wire _3018_ ;
wire _1924_ ;
wire _1504_ ;
wire _835_ ;
wire _415_ ;
wire [3:0] \z1.z2.q1  ;
wire _2709_ ;
wire _95_ ;
wire \z4.z3.z3.z2.a  ;
wire _2882_ ;
wire _2462_ ;
wire _2042_ ;
wire \z3.z1.z1.z2.s  ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2938_ ;
wire _2518_ ;
wire _2691_ ;
wire _2271_ ;
wire _1962_ ;
wire _1542_ ;
wire _1122_ ;
wire \z1.z3.z2.z2.c  ;
wire _873_ ;
wire _453_ ;
wire _2747_ ;
wire _2327_ ;
wire _2080_ ;
wire _929_ ;
wire _509_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _2976_ ;
wire _2556_ ;
wire _2136_ ;
wire _1827_ ;
wire _1407_ ;
wire _738_ ;
wire _318_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _2785_ ;
wire _2365_ ;
wire \z1.z3.z3.z1.s  ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _2594_ ;
wire _2174_ ;
wire \z4.z3.z4.z1.s  ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire \z2.z3.z2.z1.a  ;
wire _776_ ;
wire _356_ ;
wire \z3.z4.z2.z2.c  ;
wire \z2.z1.z4.z2.a  ;
wire \z3.z1.z2.z1.c  ;
wire _1674_ ;
wire _1254_ ;
wire _585_ ;
wire _165_ ;
wire _2879_ ;
wire _2459_ ;
wire _2039_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _2900_ ;
wire _1292_ ;
wire _2497_ ;
wire _2077_ ;
wire \z1.z3.z4.z1.b  ;
wire _1768_ ;
wire _1348_ ;
wire _679_ ;
wire _259_ ;
wire \z4.z4.z2.z1.a  ;
wire \z4.z2.z4.z2.a  ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _700_ ;
wire _1386_ ;
wire \z1.z4.z1.z1.c  ;
wire _297_ ;
wire _16_ ;
wire \z1.z2.z3.z2.c  ;
wire _2803_ ;
wire _1195_ ;
wire \z3.z4.z4.z1.b  ;
wire _2612_ ;
wire _54_ ;
wire _2841_ ;
wire _2421_ ;
wire _2001_ ;
wire \z1.z2.z4.z1.s  ;
wire [3:0] \z3.z1.q2  ;
wire _603_ ;
wire _1289_ ;
wire _2650_ ;
wire _2230_ ;
wire _3015_ ;
wire \z1.z3.z1.z2.s  ;
wire _1921_ ;
wire _1501_ ;
wire \z2.z2.z3.z1.a  ;
wire [3:0] \z2.z4.q1  ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _92_ ;
wire \z3.z3.z3.z2.c  ;
wire _1098_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _2935_ ;
wire _2515_ ;
wire [31:0] _3053_ ;
wire _870_ ;
wire _450_ ;
wire _2744_ ;
wire _2324_ ;
wire _926_ ;
wire _506_ ;
wire _2973_ ;
wire _2553_ ;
wire _2133_ ;
wire _1824_ ;
wire _1404_ ;
wire _735_ ;
wire _315_ ;
wire \z3.z4.z1.z2.s  ;
wire _2609_ ;
wire \z4.z3.z3.z1.a  ;
wire _2782_ ;
wire _2362_ ;
wire \z3.z1.z1.z1.s  ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2838_ ;
wire _2418_ ;
wire _2591_ ;
wire _2171_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire \z1.z3.z2.z1.c  ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _1918_ ;
wire \z1.z1.z4.z2.c  ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _2876_ ;
wire _2456_ ;
wire _2036_ ;
wire _1727_ ;
wire _1307_ ;
wire _638_ ;
wire _218_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _2685_ ;
wire _2265_ ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _2494_ ;
wire _2074_ ;
wire _1765_ ;
wire _1345_ ;
wire \z2.z4.z4.z2.a  ;
wire _676_ ;
wire _256_ ;
wire \z3.z4.z2.z1.c  ;
wire \z1.z2.z2.z2.s  ;
wire \z2.z1.z4.z1.a  ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire \z3.z2.z4.z2.c  ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _1383_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire _13_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _1192_ ;
wire \z2.z2.z1.z1.b  ;
wire _2397_ ;
wire _1668_ ;
wire _1248_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire \z3.z3.z2.z2.s  ;
wire _51_ ;
wire \z4.z2.z4.z1.a  ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire [3:0] \z4.z3.q2  ;
wire _600_ ;
wire _1286_ ;
wire _197_ ;
wire _3012_ ;
wire \z4.z3.z1.z2.a  ;
wire \z1.z2.z3.z1.c  ;
wire _2703_ ;
wire _1095_ ;
wire _2932_ ;
wire _2512_ ;
wire _3050_ ;
wire _2741_ ;
wire _2321_ ;
wire _7_ ;
wire _923_ ;
wire _503_ ;
wire _1189_ ;
wire _2970_ ;
wire _2550_ ;
wire _2130_ ;
wire \z1.z3.z1.z1.s  ;
wire _1821_ ;
wire _1401_ ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire \z3.z3.z3.z1.c  ;
wire \z1.z1.z3.z2.s  ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2835_ ;
wire _2415_ ;
wire _770_ ;
wire _350_ ;
wire _2644_ ;
wire _2224_ ;
wire _3009_ ;
wire _1915_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire \z2.z1.z2.z1.b  ;
wire _2873_ ;
wire _2453_ ;
wire _2033_ ;
wire _1724_ ;
wire _1304_ ;
wire _635_ ;
wire _215_ ;
wire \z3.z4.z1.z1.s  ;
wire _2929_ ;
wire _2509_ ;
wire _2682_ ;
wire _2262_ ;
wire _3047_ ;
wire \z3.z2.z3.z2.s  ;
wire _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire \z1.z2.z1.z2.a  ;
wire _2491_ ;
wire _2071_ ;
wire _1762_ ;
wire _1342_ ;
wire \z1.z4.z4.z2.c  ;
wire _673_ ;
wire _253_ ;
wire _2967_ ;
wire _2547_ ;
wire _2127_ ;
wire \z4.z2.z2.z2.a  ;
wire [3:0] \z3.z4.q3  ;
wire _1818_ ;
wire \z1.z1.z4.z1.c  ;
wire _729_ ;
wire _309_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _2776_ ;
wire _2356_ ;
wire _1627_ ;
wire _1207_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _1380_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _10_ ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _2394_ ;
wire [3:0] \z2.z2.q2  ;
wire _1665_ ;
wire _1245_ ;
wire \z2.z4.z4.z1.a  ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire \z1.z2.z2.z1.s  ;
wire _1894_ ;
wire _1474_ ;
wire _1054_ ;
wire \z3.z2.z4.z1.c  ;
wire _385_ ;
wire _2679_ ;
wire _2259_ ;
wire _1283_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire \z3.z3.z1.z2.c  ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _1092_ ;
wire _2297_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire \z3.z3.z2.z1.s  ;
wire _1797_ ;
wire _1377_ ;
wire _288_ ;
wire _4_ ;
wire [7:0] \z3.q1  ;
wire \z3.z1.z4.z2.s  ;
wire _920_ ;
wire _500_ ;
wire \z1.z1.z2.z2.a  ;
wire _1186_ ;
wire \z4.z3.z1.z1.a  ;
wire _2603_ ;
wire \z4.z1.z3.z2.a  ;
wire _45_ ;
wire _2832_ ;
wire _2412_ ;
wire _2641_ ;
wire _2221_ ;
wire _3006_ ;
wire _1912_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _1089_ ;
wire _2870_ ;
wire _2450_ ;
wire _2030_ ;
wire [15:0] q0 ;
wire [15:0] q1 ;
wire [15:0] q2 ;
wire [15:0] q3 ;
wire \z1.z4.z3.z2.s  ;
wire _1721_ ;
wire _1301_ ;
wire _632_ ;
wire _212_ ;
wire _2926_ ;
wire _2506_ ;
wire [3:0] \z1.z3.q3  ;
wire \z1.z1.z3.z1.s  ;
wire _3044_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _2964_ ;
wire _2544_ ;
wire _2124_ ;
wire \z3.z2.z2.z2.c  ;
wire \z2.z4.z2.z1.b  ;
wire _1815_ ;
wire _726_ ;
wire _306_ ;
wire _2773_ ;
wire _2353_ ;
wire _1624_ ;
wire _1204_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2829_ ;
wire _2409_ ;
wire [3:0] \z4.z1.q3  ;
wire _2582_ ;
wire _2162_ ;
wire \z3.z2.z3.z1.s  ;
wire _1853_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire \z1.z2.z1.z1.a  ;
wire _2391_ ;
wire _1909_ ;
wire _1662_ ;
wire _1242_ ;
wire \z1.z4.z4.z1.c  ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2867_ ;
wire _2447_ ;
wire _2027_ ;
wire \z4.z2.z2.z1.a  ;
wire _1718_ ;
wire _629_ ;
wire _209_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _858_ ;
wire _438_ ;
wire _1280_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _2294_ ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire \z1.z3.z4.z2.s  ;
wire _1794_ ;
wire _1374_ ;
wire _285_ ;
wire _2999_ ;
wire _2579_ ;
wire _2159_ ;
wire _1_ ;
wire _1183_ ;
wire _2388_ ;
wire \z3.z3.z1.z1.c  ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire \z3.z1.z3.z2.c  ;
wire \z2.z3.z3.z1.b  ;
wire _2197_ ;
wire _42_ ;
wire _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire \z3.z4.z4.z2.s  ;
wire _1697_ ;
wire _1277_ ;
wire _188_ ;
wire _3003_ ;
wire \z1.z4.z2.z2.a  ;
wire \z3.z1.z4.z1.s  ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire \z1.z1.z2.z1.a  ;
wire _1086_ ;
wire \z4.z4.z3.z2.a  ;
wire _2923_ ;
wire _2503_ ;
wire \z4.z1.z3.z1.a  ;
wire _3041_ ;
wire _2732_ ;
wire _2312_ ;
wire _914_ ;
wire _2961_ ;
wire _2541_ ;
wire _2121_ ;
wire _1812_ ;
wire _723_ ;
wire _303_ ;
wire _2770_ ;
wire _2350_ ;
wire \z1.z4.z3.z1.s  ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2826_ ;
wire _2406_ ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire _1906_ ;
wire _817_ ;
wire _77_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _2864_ ;
wire _2444_ ;
wire _2024_ ;
wire \z3.z2.z2.z1.c  ;
wire _1715_ ;
wire _626_ ;
wire _206_ ;
wire \z2.z2.z4.z1.b  ;
wire _2673_ ;
wire _2253_ ;
wire _3038_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire [7:0] \z1.q2  ;
wire _2729_ ;
wire _2309_ ;
wire _2482_ ;
wire _2062_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _2958_ ;
wire _2538_ ;
wire _2118_ ;
wire \z1.z3.z3.z2.a  ;
wire _2291_ ;
wire _1809_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire \z4.z3.z4.z2.a  ;
wire _1618_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _1791_ ;
wire _1371_ ;
wire _282_ ;
wire _2996_ ;
wire _2576_ ;
wire _2156_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _758_ ;
wire _338_ ;
wire _1180_ ;
wire _2385_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _2194_ ;
wire \z4.z1.z1.z1.b  ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire \z2.z2.z1.z2.s  ;
wire _376_ ;
wire \z1.z3.z4.z1.s  ;
wire _1694_ ;
wire _1274_ ;
wire _185_ ;
wire _2899_ ;
wire _2479_ ;
wire _2059_ ;
wire _3000_ ;
wire [3:0] \z3.z2.q1  ;
wire _1083_ ;
wire _2288_ ;
wire \z3.z4.z3.z2.c  ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2920_ ;
wire _2500_ ;
wire \z3.z1.z3.z1.c  ;
wire _2097_ ;
wire _1788_ ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire \z3.z4.z4.z1.s  ;
wire _1597_ ;
wire _1177_ ;
wire \z1.z4.z2.z1.a  ;
wire _720_ ;
wire _300_ ;
wire \z1.z2.z4.z2.a  ;
wire \z4.z4.z3.z1.a  ;
wire _36_ ;
wire _2823_ ;
wire _2403_ ;
wire _2632_ ;
wire _2212_ ;
wire _1903_ ;
wire _814_ ;
wire _74_ ;
wire _2861_ ;
wire _2441_ ;
wire _2021_ ;
wire _1712_ ;
wire _623_ ;
wire _203_ ;
wire _2917_ ;
wire _2670_ ;
wire _2250_ ;
wire _3035_ ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire \z2.z1.z2.z2.s  ;
wire _2726_ ;
wire _2306_ ;
wire _908_ ;
wire _1750_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire _2955_ ;
wire _2535_ ;
wire _2115_ ;
wire \z3.z1.z1.z2.a  ;
wire _1806_ ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _2764_ ;
wire _2344_ ;
wire \z3.z3.z4.z2.c  ;
wire _1615_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _2993_ ;
wire _2573_ ;
wire _2153_ ;
wire _1844_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _2629_ ;
wire _2209_ ;
wire _2382_ ;
wire \z2.z3.z1.z1.b  ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2858_ ;
wire _2438_ ;
wire _2018_ ;
wire \z1.z3.z3.z1.a  ;
wire _2191_ ;
wire [3:0] \z1.z1.q1  ;
wire _1709_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire \z4.z3.z4.z1.a  ;
wire _1938_ ;
wire _1518_ ;
wire _849_ ;
wire _429_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _2896_ ;
wire _2476_ ;
wire _2056_ ;
wire [3:0] \z4.z4.q1  ;
wire _1747_ ;
wire _1327_ ;
wire _658_ ;
wire _238_ ;
wire _1080_ ;
wire _2285_ ;
wire \z4.z4.z1.z1.b  ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _2094_ ;
wire _1785_ ;
wire _1365_ ;
wire _696_ ;
wire \z2.z2.z1.z1.s  ;
wire _276_ ;
wire _1594_ ;
wire _1174_ ;
wire _2799_ ;
wire _2379_ ;
wire [15:0] \z4.q3  ;
wire _2188_ ;
wire \z3.z4.z3.z1.c  ;
wire _33_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2820_ ;
wire _2400_ ;
wire _1688_ ;
wire _1268_ ;
wire _599_ ;
wire _179_ ;
wire _1900_ ;
wire _811_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire \z2.z2.z2.z1.b  ;
wire _620_ ;
wire _200_ ;
wire _2914_ ;
wire \z1.z2.z4.z1.a  ;
wire _3032_ ;
wire _2723_ ;
wire _2303_ ;
wire \z1.z3.z1.z2.a  ;
wire _905_ ;
wire _2952_ ;
wire _2532_ ;
wire _2112_ ;
wire _1803_ ;
wire \z2.z1.z1.z2.c  ;
wire _714_ ;
wire _2761_ ;
wire _2341_ ;
wire _1612_ ;
wire \z4.z3.z2.z1.b  ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _2817_ ;
wire _2990_ ;
wire _2570_ ;
wire _2150_ ;
wire \z2.z4.z2.z2.s  ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire \z2.z1.z2.z1.s  ;
wire _2626_ ;
wire _2206_ ;
wire _808_ ;
wire _68_ ;
wire _1650_ ;
wire _1230_ ;
wire \z3.z4.z1.z2.a  ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2855_ ;
wire _2435_ ;
wire _2015_ ;
wire [3:0] \z2.z3.q1  ;
wire \z3.z1.z1.z1.a  ;
wire _1706_ ;
wire _617_ ;
wire \z4.z2.z1.z2.c  ;
wire _790_ ;
wire _370_ ;
wire _2664_ ;
wire _2244_ ;
wire _3029_ ;
wire \z3.z3.z4.z1.c  ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _2893_ ;
wire _2473_ ;
wire _2053_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _2949_ ;
wire _2529_ ;
wire _2109_ ;
wire _2282_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire \z2.z1.z3.z1.b  ;
wire _2091_ ;
wire _1609_ ;
wire _1782_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _2987_ ;
wire _2567_ ;
wire _2147_ ;
wire _1838_ ;
wire _1418_ ;
wire _749_ ;
wire _329_ ;
wire _1591_ ;
wire _1171_ ;
wire _2796_ ;
wire _2376_ ;
wire \z1.z2.z2.z2.a  ;
wire [7:0] \z4.q0  ;
wire _1647_ ;
wire _1227_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _2185_ ;
wire _30_ ;
wire _1876_ ;
wire _1456_ ;
wire _1036_ ;
wire _787_ ;
wire _367_ ;
wire \z4.z2.z3.z1.b  ;
wire _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire \z2.z3.z3.z2.s  ;
wire _1494_ ;
wire _1074_ ;
wire _2699_ ;
wire _2279_ ;
wire \z3.z3.z2.z2.a  ;
wire _2911_ ;
wire _2088_ ;
wire \z4.z1.z2.z2.c  ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire [3:0] \z1.z4.q2  ;
wire _902_ ;
wire _1588_ ;
wire _1168_ ;
wire _499_ ;
wire _1800_ ;
wire _711_ ;
wire _1397_ ;
wire _27_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _2623_ ;
wire _2203_ ;
wire [3:0] \z4.z2.q2  ;
wire \z1.z3.z1.z1.a  ;
wire _805_ ;
wire _65_ ;
wire \z2.z4.z1.z2.c  ;
wire _2852_ ;
wire _2432_ ;
wire _2012_ ;
wire \z1.z1.z3.z2.a  ;
wire _1703_ ;
wire \z2.z1.z1.z1.c  ;
wire _614_ ;
wire _2908_ ;
wire _2661_ ;
wire _2241_ ;
wire _3026_ ;
wire _1932_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _2890_ ;
wire _2470_ ;
wire _2050_ ;
wire \z2.z4.z2.z1.s  ;
wire \z4.z1.z4.z1.b  ;
wire _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _2946_ ;
wire _2526_ ;
wire \z2.z2.z4.z2.s  ;
wire _2106_ ;
wire _708_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire \z3.z4.z1.z1.a  ;
wire _881_ ;
wire _461_ ;
wire _2755_ ;
wire _2335_ ;
wire \z3.z2.z3.z2.a  ;
wire _1606_ ;
wire _937_ ;
wire _517_ ;
wire \z4.z2.z1.z1.c  ;
wire _690_ ;
wire _270_ ;
wire _2984_ ;
wire _2564_ ;
wire _2144_ ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _2793_ ;
wire _2373_ ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2849_ ;
wire _2429_ ;
wire _2009_ ;
wire _2182_ ;
wire \z2.z4.z3.z1.b  ;
wire _1873_ ;
wire _1453_ ;
wire _1033_ ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _1929_ ;
wire _1509_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _2887_ ;
wire _2467_ ;
wire _2047_ ;
wire \z4.z1.z1.z2.s  ;
wire _1738_ ;
wire _1318_ ;
wire _649_ ;
wire _229_ ;
wire _1491_ ;
wire _1071_ ;
wire _2696_ ;
wire _2276_ ;
wire \z1.z2.z2.z1.a  ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire \z2.z3.z2.z2.c  ;
wire _878_ ;
wire _458_ ;
wire [3:0] \z3.z3.q3  ;
wire _2085_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire \z2.z3.z3.z1.s  ;
wire _1394_ ;
wire [3:0] \z2.z1.q2  ;
wire _2599_ ;
wire _2179_ ;
wire _24_ ;
wire \z3.z3.z2.z1.a  ;
wire _2811_ ;
wire \z4.z4.z2.z2.c  ;
wire \z3.z1.z4.z2.a  ;
wire \z4.z1.z2.z1.c  ;
wire _1679_ ;
wire _1259_ ;
wire _2620_ ;
wire _2200_ ;
wire _802_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _399_ ;
wire _1700_ ;
wire _611_ ;
wire _2905_ ;
wire _1297_ ;
wire _3023_ ;
wire \z2.z3.z4.z1.b  ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _2943_ ;
wire _2523_ ;
wire _2103_ ;
wire [7:0] \z2.q1  ;
wire \z1.z4.z3.z2.a  ;
wire _705_ ;
wire \z2.z4.z1.z1.c  ;
wire _2752_ ;
wire _2332_ ;
wire \z1.z1.z3.z1.a  ;
wire _1603_ ;
wire \z2.z2.z3.z2.c  ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire _2981_ ;
wire _2561_ ;
wire _2141_ ;
wire _1832_ ;
wire _1412_ ;
wire \z4.z4.z4.z1.b  ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _2790_ ;
wire _2370_ ;
wire _59_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2846_ ;
wire _2426_ ;
wire \z2.z2.z4.z1.s  ;
wire _2006_ ;
wire _608_ ;
wire _1870_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire \z2.z3.z1.z2.s  ;
wire \z3.z2.z3.z1.a  ;
wire _1926_ ;
wire _1506_ ;
wire _837_ ;
wire _417_ ;
wire [3:0] \z1.z2.q3  ;
wire _97_ ;
wire \z4.z3.z3.z2.c  ;
wire _590_ ;
wire _170_ ;
wire _2884_ ;
wire _2464_ ;
wire _2044_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire _2693_ ;
wire _2273_ ;
wire _1964_ ;
wire _1544_ ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _2082_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _2978_ ;
wire _2558_ ;
wire _2138_ ;
wire _1829_ ;
wire _1409_ ;
wire \z4.z4.z1.z2.s  ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _2787_ ;
wire _2367_ ;
wire \z4.z1.z1.z1.s  ;
wire _1638_ ;
wire _1218_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _1391_ ;
wire _2596_ ;
wire _2176_ ;
wire \z1.z3.z4.z2.a  ;
wire _21_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire \z2.z3.z2.z1.c  ;
wire _778_ ;
wire _358_ ;
wire \z2.z1.z4.z2.c  ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _1485_ ;
wire _1065_ ;
wire _396_ ;
wire \z1.z1.z1.z1.b  ;
wire _2902_ ;
wire _1294_ ;
wire _2499_ ;
wire _2079_ ;
wire _3020_ ;
wire \z3.z4.z4.z2.a  ;
wire _2711_ ;
wire \z4.z4.z2.z1.c  ;
wire \z2.z2.z2.z2.s  ;
wire \z3.z1.z4.z1.a  ;
wire \z4.z2.z4.z2.c  ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _2940_ ;
wire _2520_ ;
wire _2100_ ;
wire _702_ ;
wire _1388_ ;
wire _299_ ;
wire _18_ ;
wire _1600_ ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire \z3.z2.z1.z1.b  ;
wire _1197_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire \z4.z3.z2.z2.s  ;
wire _56_ ;
wire _2843_ ;
wire _2423_ ;
wire _2003_ ;
wire \z1.z4.z3.z1.a  ;
wire _605_ ;
wire _2652_ ;
wire _2232_ ;
wire _3017_ ;
wire _1923_ ;
wire _1503_ ;
wire \z2.z2.z3.z1.c  ;
wire [3:0] \z2.z4.q3  ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _2881_ ;
wire _2461_ ;
wire _2041_ ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _2937_ ;
wire _2517_ ;
wire _2690_ ;
wire _2270_ ;
wire _1961_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire _928_ ;
wire _508_ ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _2975_ ;
wire _2555_ ;
wire _2135_ ;
wire \z2.z3.z1.z1.s  ;
wire _1826_ ;
wire _1406_ ;
wire _737_ ;
wire _317_ ;
wire \z4.z3.z3.z1.c  ;
wire _490_ ;
wire _2784_ ;
wire _2364_ ;
wire \z2.z1.z3.z2.s  ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _2593_ ;
wire _2173_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _2649_ ;
wire _2229_ ;
wire \z3.z1.z2.z1.b  ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _2878_ ;
wire _2458_ ;
wire _2038_ ;
wire _1729_ ;
wire _1309_ ;
wire \z4.z4.z1.z1.s  ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _2687_ ;
wire _2267_ ;
wire \z4.z2.z3.z2.s  ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _869_ ;
wire _449_ ;
wire _1291_ ;
wire \z2.z2.z1.z2.a  ;
wire _2496_ ;
wire _2076_ ;
wire \z1.z3.z4.z1.a  ;
wire _1767_ ;
wire _1347_ ;
wire \z2.z4.z4.z2.c  ;
wire _678_ ;
wire _258_ ;
wire \z2.z1.z4.z1.c  ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _1385_ ;
wire \z1.z4.z1.z1.b  ;
wire _296_ ;
wire _15_ ;
wire _2802_ ;
wire _1194_ ;
wire _2399_ ;
wire \z3.z4.z4.z1.a  ;
wire _2611_ ;
wire \z2.z2.z2.z1.s  ;
wire _53_ ;
wire \z4.z2.z4.z1.c  ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _2840_ ;
wire _2420_ ;
wire _2000_ ;
wire [3:0] \z3.z1.q1  ;
wire _602_ ;
wire _1288_ ;
wire _199_ ;
wire _3014_ ;
wire \z4.z3.z1.z2.c  ;
wire _1920_ ;
wire _1500_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _91_ ;
wire _1097_ ;
wire _640_ ;
wire _220_ ;
wire _2934_ ;
wire _2514_ ;
wire _3052_ ;
wire \z4.z3.z2.z1.s  ;
wire _2743_ ;
wire _2323_ ;
wire _9_ ;
wire \z4.z1.z4.z2.s  ;
wire _925_ ;
wire _505_ ;
wire \z2.z1.z2.z2.a  ;
wire _2972_ ;
wire _2552_ ;
wire _2132_ ;
wire _1823_ ;
wire _1403_ ;
wire _734_ ;
wire _314_ ;
wire _2608_ ;
wire _2781_ ;
wire _2361_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2837_ ;
wire _2417_ ;
wire _2590_ ;
wire _2170_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire \z1.z3.z2.z1.b  ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire _1917_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _2875_ ;
wire _2455_ ;
wire _2035_ ;
wire \z2.z4.z3.z2.s  ;
wire _1726_ ;
wire _1306_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _2684_ ;
wire _2264_ ;
wire \z2.z1.z3.z1.s  ;
wire _3049_ ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire \z1.z2.z1.z2.c  ;
wire _2493_ ;
wire _2073_ ;
wire _1764_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _2969_ ;
wire _2549_ ;
wire _2129_ ;
wire \z4.z2.z2.z2.c  ;
wire \z3.z4.z2.z1.b  ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _1629_ ;
wire _1209_ ;
wire _1382_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire \z4.z2.z3.z1.s  ;
wire _12_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _769_ ;
wire _349_ ;
wire _1191_ ;
wire \z2.z2.z1.z1.a  ;
wire _2396_ ;
wire _1667_ ;
wire _1247_ ;
wire \z2.z4.z4.z1.c  ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire [3:0] \z4.z3.q1  ;
wire _1285_ ;
wire _196_ ;
wire _3011_ ;
wire \z1.z2.z3.z1.b  ;
wire _2702_ ;
wire _1094_ ;
wire _2299_ ;
wire _2931_ ;
wire _2511_ ;
wire \z2.z3.z4.z2.s  ;
wire _1799_ ;
wire _1379_ ;
wire _2740_ ;
wire _2320_ ;
wire _6_ ;
wire [15:0] \z3.q3  ;
wire _922_ ;
wire _502_ ;
wire \z1.z1.z2.z2.c  ;
wire _1188_ ;
wire \z4.z3.z1.z1.c  ;
wire _1820_ ;
wire _1400_ ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire \z4.z1.z3.z2.c  ;
wire \z3.z3.z3.z1.b  ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2834_ ;
wire _2414_ ;
wire \z4.z4.z4.z2.s  ;
wire _2643_ ;
wire _2223_ ;
wire _3008_ ;
wire \z2.z4.z2.z2.a  ;
wire \z4.z1.z4.z1.s  ;
wire _1914_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire \z2.z1.z2.z1.a  ;
wire _2872_ ;
wire _2452_ ;
wire _2032_ ;
wire _1723_ ;
wire _1303_ ;
wire _634_ ;
wire _214_ ;
wire _2928_ ;
wire _2508_ ;
wire _2681_ ;
wire _2261_ ;
wire _3046_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _2490_ ;
wire _2070_ ;
wire _919_ ;
wire _1761_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _2966_ ;
wire _2546_ ;
wire _2126_ ;
wire [3:0] \z3.z4.q2  ;
wire _1817_ ;
wire \z1.z1.z4.z1.b  ;
wire _728_ ;
wire _308_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _2775_ ;
wire _2355_ ;
wire \z2.z4.z3.z1.s  ;
wire _1626_ ;
wire _1206_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _2584_ ;
wire _2164_ ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire \z1.z2.z1.z1.c  ;
wire _2393_ ;
wire [3:0] \z2.z2.q1  ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2869_ ;
wire _2449_ ;
wire _2029_ ;
wire \z4.z2.z2.z1.c  ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire \z3.z2.z4.z1.b  ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _1282_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _1758_ ;
wire _1338_ ;
wire _669_ ;
wire _249_ ;
wire _1091_ ;
wire \z2.z3.z3.z2.a  ;
wire _2296_ ;
wire \z1.z1.z1.z2.s  ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _1796_ ;
wire _1376_ ;
wire _287_ ;
wire _3_ ;
wire [7:0] \z3.q0  ;
wire _1185_ ;
wire _2602_ ;
wire _2199_ ;
wire _44_ ;
wire _2831_ ;
wire _2411_ ;
wire \z3.z2.z1.z2.s  ;
wire \z2.z3.z4.z1.s  ;
wire _1699_ ;
wire _1279_ ;
wire _2640_ ;
wire _2220_ ;
wire _3005_ ;
wire \z1.z4.z2.z2.c  ;
wire _1911_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire \z1.z1.z2.z1.c  ;
wire _1088_ ;
wire \z4.z4.z3.z2.c  ;
wire _1720_ ;
wire _1300_ ;
wire _631_ ;
wire _211_ ;
wire _2925_ ;
wire _2505_ ;
wire [3:0] \z1.z3.q2  ;
wire \z4.z1.z3.z1.c  ;
wire _3043_ ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _916_ ;
wire \z4.z4.z4.z1.s  ;
wire _2963_ ;
wire _2543_ ;
wire _2123_ ;
wire \z2.z4.z2.z1.a  ;
wire _1814_ ;
wire _725_ ;
wire _305_ ;
wire \z2.z2.z4.z2.a  ;
wire _2772_ ;
wire _2352_ ;
wire _1623_ ;
wire _1203_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2828_ ;
wire _2408_ ;
wire [3:0] \z4.z1.q2  ;
wire _2581_ ;
wire _2161_ ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _2390_ ;
wire _1908_ ;
wire _819_ ;
wire _79_ ;
wire _1661_ ;
wire _1241_ ;
wire \z1.z4.z4.z1.b  ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2866_ ;
wire _2446_ ;
wire _2026_ ;
wire _1717_ ;
wire _628_ ;
wire _208_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire \z3.z1.z2.z2.s  ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _2484_ ;
wire _2064_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire \z1.z3.z3.z2.c  ;
wire _2293_ ;
wire \z4.z1.z1.z2.a  ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire \z4.z3.z4.z2.c  ;
wire _1793_ ;
wire _1373_ ;
wire _284_ ;
wire _2998_ ;
wire _2578_ ;
wire _2158_ ;
wire _0_ ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _1182_ ;
wire _2387_ ;
wire \z3.z3.z1.z1.b  ;
wire _1658_ ;
wire _1238_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire \z1.z4.z1.z2.s  ;
wire \z2.z3.z3.z1.a  ;
wire _2196_ ;
wire \z1.z1.z1.z1.s  ;
wire _41_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _1696_ ;
wire _1276_ ;
wire _187_ ;
wire _3002_ ;
wire [3:0] \z3.z2.q3  ;
wire _1085_ ;
wire _2922_ ;
wire _2502_ ;
wire _2099_ ;
wire _3040_ ;
wire _2731_ ;
wire _2311_ ;
wire \z3.z2.z1.z1.s  ;
wire _913_ ;
wire _1599_ ;
wire _1179_ ;
wire _2960_ ;
wire _2540_ ;
wire _2120_ ;
wire \z1.z4.z2.z1.c  ;
wire _1811_ ;
wire _722_ ;
wire _302_ ;
wire \z1.z2.z4.z2.c  ;
wire \z4.z4.z3.z1.c  ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2825_ ;
wire _2405_ ;
wire _760_ ;
wire _340_ ;
wire _2634_ ;
wire _2214_ ;
wire _1905_ ;
wire _816_ ;
wire _76_ ;
wire _2863_ ;
wire _2443_ ;
wire _2023_ ;
wire \z3.z2.z2.z1.b  ;
wire _1714_ ;
wire _625_ ;
wire _205_ ;
wire _2919_ ;
wire \z1.z3.z2.z2.s  ;
wire \z2.z2.z4.z1.a  ;
wire _2672_ ;
wire _2252_ ;
wire _3037_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire [7:0] \z1.q1  ;
wire _2728_ ;
wire _2308_ ;
wire _2481_ ;
wire _2061_ ;
wire \z2.z3.z1.z2.a  ;
wire _1752_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _2957_ ;
wire _2537_ ;
wire _2117_ ;
wire _2290_ ;
wire \z3.z1.z1.z2.c  ;
wire _1808_ ;
wire _719_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _1617_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _1790_ ;
wire _1370_ ;
wire _281_ ;
wire _2995_ ;
wire _2575_ ;
wire _2155_ ;
wire \z3.z4.z2.z2.s  ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire \z3.z1.z2.z1.s  ;
wire _757_ ;
wire _337_ ;
wire _2384_ ;
wire \z4.z4.z1.z2.a  ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire \z1.z3.z3.z1.c  ;
wire _2193_ ;
wire \z4.z1.z1.z1.a  ;
wire [3:0] \z1.z1.q3  ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire \z4.z3.z4.z1.c  ;
wire _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _2898_ ;
wire _2478_ ;
wire _2058_ ;
wire [3:0] \z4.z4.q3  ;
wire _1749_ ;
wire _1329_ ;
wire _1082_ ;
wire _2287_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _889_ ;
wire _469_ ;
wire \z1.z4.z1.z1.s  ;
wire \z3.z1.z3.z1.b  ;
wire _2096_ ;
wire \z1.z2.z3.z2.s  ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _1596_ ;
wire _1176_ ;
wire \z2.z2.z2.z2.a  ;
wire _35_ ;
wire _2822_ ;
wire _2402_ ;
wire _2631_ ;
wire _2211_ ;
wire \z3.z3.z3.z2.s  ;
wire _1902_ ;
wire _813_ ;
wire _73_ ;
wire _1499_ ;
wire _1079_ ;
wire _2860_ ;
wire _2440_ ;
wire _2020_ ;
wire _1711_ ;
wire \z4.z3.z2.z2.a  ;
wire _622_ ;
wire _202_ ;
wire _2916_ ;
wire \z1.z2.z4.z1.c  ;
wire _3034_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _2725_ ;
wire _2305_ ;
wire \z1.z3.z1.z2.c  ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _2954_ ;
wire _2534_ ;
wire _2114_ ;
wire _1805_ ;
wire _716_ ;
wire _2763_ ;
wire _2343_ ;
wire _1614_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2819_ ;
wire \z1.z3.z2.z1.s  ;
wire _2992_ ;
wire _2572_ ;
wire _2152_ ;
wire \z1.z1.z4.z2.s  ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _2628_ ;
wire _2208_ ;
wire _2381_ ;
wire \z2.z3.z1.z1.a  ;
wire _1652_ ;
wire _1232_ ;
wire \z3.z4.z1.z2.c  ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2857_ ;
wire _2437_ ;
wire _2017_ ;
wire \z2.z1.z3.z2.a  ;
wire _2190_ ;
wire [3:0] \z2.z3.q3  ;
wire \z3.z1.z1.z1.c  ;
wire _1708_ ;
wire _619_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire _1937_ ;
wire _1517_ ;
wire _848_ ;
wire _428_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _2895_ ;
wire _2475_ ;
wire _2055_ ;
wire \z3.z4.z2.z1.s  ;
wire _1746_ ;
wire _1326_ ;
wire \z3.z2.z4.z2.s  ;
wire _657_ ;
wire _237_ ;
wire _2284_ ;
wire \z4.z4.z1.z1.a  ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _2093_ ;
wire \z4.z2.z3.z2.a  ;
wire _1784_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _2989_ ;
wire _2569_ ;
wire _2149_ ;
wire _1593_ ;
wire _1173_ ;
wire _2798_ ;
wire _2378_ ;
wire \z1.z2.z2.z2.c  ;
wire [7:0] \z4.q2  ;
wire _1649_ ;
wire _1229_ ;
wire _2187_ ;
wire \z3.z4.z3.z1.b  ;
wire _32_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _789_ ;
wire _369_ ;
wire \z1.z2.z3.z1.s  ;
wire _1687_ ;
wire _1267_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire \z2.z2.z2.z1.a  ;
wire \z3.z3.z2.z2.c  ;
wire _2913_ ;
wire _3031_ ;
wire _2722_ ;
wire _2302_ ;
wire _904_ ;
wire _2951_ ;
wire _2531_ ;
wire _2111_ ;
wire \z3.z3.z3.z1.s  ;
wire _1802_ ;
wire _713_ ;
wire _1399_ ;
wire _2760_ ;
wire _2340_ ;
wire _29_ ;
wire _1611_ ;
wire \z4.z3.z2.z1.a  ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _2816_ ;
wire \z4.z1.z4.z2.a  ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire \z1.z3.z1.z1.c  ;
wire _807_ ;
wire _67_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _2854_ ;
wire _2434_ ;
wire _2014_ ;
wire \z1.z1.z3.z2.c  ;
wire _1705_ ;
wire _616_ ;
wire _2663_ ;
wire _2243_ ;
wire _3028_ ;
wire \z3.z3.z4.z1.b  ;
wire _1934_ ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire \z1.z4.z4.z2.s  ;
wire _2892_ ;
wire _2472_ ;
wire _2052_ ;
wire \z1.z1.z4.z1.s  ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire _2948_ ;
wire _2528_ ;
wire _2108_ ;
wire _2281_ ;
wire \z2.z4.z3.z2.a  ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire \z3.z4.z1.z1.c  ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire \z2.z1.z3.z1.a  ;
wire _2090_ ;
wire \z3.z2.z3.z2.c  ;
wire _1608_ ;
wire _939_ ;
wire _519_ ;
wire _1781_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _2986_ ;
wire _2566_ ;
wire _2146_ ;
wire _1837_ ;
wire _1417_ ;
wire _748_ ;
wire _328_ ;
wire _1590_ ;
wire _1170_ ;
wire _2795_ ;
wire _2375_ ;
wire _1646_ ;
wire _1226_ ;
wire \z3.z2.z4.z1.s  ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _2184_ ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire \z3.z3.z1.z2.s  ;
wire \z4.z2.z3.z1.a  ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _2889_ ;
wire _2469_ ;
wire _2049_ ;
wire _1493_ ;
wire _1073_ ;
wire _2698_ ;
wire _2278_ ;
wire \z1.z2.z2.z1.c  ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2910_ ;
wire _2087_ ;
wire _1778_ ;
wire _1358_ ;
wire _689_ ;
wire _269_ ;
wire [3:0] \z1.z4.q1  ;
wire _901_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _710_ ;
wire _1396_ ;
wire \z2.z3.z4.z2.a  ;
wire _26_ ;
wire \z3.z3.z2.z1.c  ;
wire _2813_ ;
wire \z3.z1.z4.z2.c  ;
wire _2622_ ;
wire _2202_ ;
wire [3:0] \z4.z2.q1  ;
wire _804_ ;
wire _64_ ;
wire _2851_ ;
wire _2431_ ;
wire _2011_ ;
wire _1702_ ;
wire \z2.z1.z1.z1.b  ;
wire _613_ ;
wire _2907_ ;
wire _1299_ ;
wire _2660_ ;
wire _2240_ ;
wire _3025_ ;
wire _1931_ ;
wire _1511_ ;
wire \z4.z4.z4.z2.a  ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire \z3.z2.z2.z2.s  ;
wire \z4.z1.z4.z1.a  ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _2945_ ;
wire _2525_ ;
wire _2105_ ;
wire [15:0] \z2.q3  ;
wire \z1.z4.z3.z2.c  ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _2754_ ;
wire _2334_ ;
wire \z1.z1.z3.z1.c  ;
wire _1605_ ;
wire _936_ ;
wire _516_ ;
wire \z4.z2.z1.z1.b  ;
wire _2983_ ;
wire _2563_ ;
wire _2143_ ;
wire _1834_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire \z1.z4.z4.z1.s  ;
wire _2792_ ;
wire _2372_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2848_ ;
wire _2428_ ;
wire _2008_ ;
wire _2181_ ;
wire \z2.z4.z3.z1.a  ;
wire _1872_ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _2657_ ;
wire _2237_ ;
wire \z3.z2.z3.z1.c  ;
wire _1928_ ;
wire _1508_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _2886_ ;
wire _2466_ ;
wire _2046_ ;
wire _1737_ ;
wire _1317_ ;
wire _648_ ;
wire _228_ ;
wire _1490_ ;
wire _1070_ ;
wire _2695_ ;
wire _2275_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire [3:0] \z3.z3.q2  ;
wire _2084_ ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire \z3.z3.z1.z1.s  ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire \z3.z1.z3.z2.s  ;
wire _2789_ ;
wire _2369_ ;
wire \z1.z1.z1.z2.a  ;
wire _1393_ ;
wire [3:0] \z2.z1.q1  ;
wire _2598_ ;
wire _2178_ ;
wire \z1.z3.z4.z2.c  ;
wire _23_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire \z4.z1.z2.z1.b  ;
wire _1678_ ;
wire _1258_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _610_ ;
wire _2904_ ;
wire \z3.z2.z1.z2.a  ;
wire _1296_ ;
wire _3022_ ;
wire \z2.z3.z4.z1.a  ;
wire \z3.z4.z4.z2.c  ;
wire _2713_ ;
wire \z3.z1.z4.z1.c  ;
wire _2942_ ;
wire _2522_ ;
wire _2102_ ;
wire [7:0] \z2.q0  ;
wire _704_ ;
wire \z2.z4.z1.z1.b  ;
wire _2751_ ;
wire _2331_ ;
wire _1602_ ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _1199_ ;
wire _2980_ ;
wire _2560_ ;
wire _2140_ ;
wire _1831_ ;
wire _1411_ ;
wire \z4.z4.z4.z1.a  ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire \z3.z2.z2.z1.s  ;
wire _58_ ;
wire _1640_ ;
wire _1220_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2845_ ;
wire _2425_ ;
wire _2005_ ;
wire \z1.z4.z3.z1.c  ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _2654_ ;
wire _2234_ ;
wire _3019_ ;
wire _1925_ ;
wire _1505_ ;
wire _836_ ;
wire _416_ ;
wire [3:0] \z1.z2.q2  ;
wire _96_ ;
wire _2883_ ;
wire _2463_ ;
wire _2043_ ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _2939_ ;
wire _2519_ ;
wire _2692_ ;
wire _2272_ ;
wire _1963_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _2081_ ;
wire \z3.z1.z2.z2.a  ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _2977_ ;
wire _2557_ ;
wire _2137_ ;
wire _1828_ ;
wire _1408_ ;
wire _739_ ;
wire _319_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _2786_ ;
wire _2366_ ;
wire _1637_ ;
wire _1217_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _1390_ ;
wire _2595_ ;
wire _2175_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire \z2.z3.z2.z1.b  ;
wire _777_ ;
wire _357_ ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire \z3.z4.z3.z2.s  ;
wire _1484_ ;
wire _1064_ ;
wire \z1.z4.z1.z2.a  ;
wire _395_ ;
wire \z3.z1.z3.z1.s  ;
wire _2689_ ;
wire _2269_ ;
wire \z1.z1.z1.z1.a  ;
wire _2901_ ;
wire _1293_ ;
wire \z2.z2.z1.z2.c  ;
wire _2498_ ;
wire _2078_ ;
wire \z1.z3.z4.z1.c  ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire \z4.z4.z2.z1.b  ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _701_ ;
wire _1387_ ;
wire _298_ ;
wire _17_ ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire \z3.z2.z1.z1.a  ;
wire _1196_ ;
wire \z3.z4.z4.z1.c  ;
wire _2613_ ;
wire _55_ ;
wire _2842_ ;
wire _2422_ ;
wire _2002_ ;
wire [3:0] \z3.z1.q3  ;
wire _604_ ;
wire _2651_ ;
wire _2231_ ;
wire _3016_ ;
wire _1922_ ;
wire _1502_ ;
wire \z2.z2.z3.z1.b  ;
wire [3:0] \z2.z4.q2  ;
wire _833_ ;
wire _413_ ;
wire _2707_ ;
wire _93_ ;
wire _1099_ ;
wire _2880_ ;
wire _2460_ ;
wire _2040_ ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _2936_ ;
wire _2516_ ;
wire \z3.z3.z4.z2.s  ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire \z1.z3.z2.z2.a  ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire _927_ ;
wire _507_ ;
wire \z2.z1.z2.z2.c  ;
wire _680_ ;
wire _260_ ;
wire _2974_ ;
wire _2554_ ;
wire _2134_ ;
wire _1825_ ;
wire _1405_ ;
wire _736_ ;
wire _316_ ;
wire \z4.z3.z3.z1.b  ;
wire _2783_ ;
wire _2363_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2839_ ;
wire _2419_ ;
wire _2592_ ;
wire _2172_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire \z3.z4.z2.z2.a  ;
wire _1919_ ;
wire \z3.z1.z2.z1.a  ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _2877_ ;
wire _2457_ ;
wire _2037_ ;
wire _1728_ ;
wire _1308_ ;
wire _639_ ;
wire _219_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire _2686_ ;
wire _2266_ ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _868_ ;
wire _448_ ;
wire _1290_ ;
wire _2495_ ;
wire _2075_ ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire \z2.z1.z4.z1.b  ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire \z3.z4.z3.z1.s  ;
wire _1384_ ;
wire \z1.z4.z1.z1.a  ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire _14_ ;
wire \z1.z2.z3.z2.a  ;
wire _2801_ ;
wire _1193_ ;
wire \z2.z2.z1.z1.c  ;
wire _2398_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _52_ ;
wire \z4.z2.z4.z1.b  ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire _389_ ;
wire [3:0] \z4.z3.q3  ;
wire _601_ ;
wire _1287_ ;
wire _198_ ;
wire _3013_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _90_ ;
wire \z3.z3.z3.z2.a  ;
wire _1096_ ;
wire \z2.z1.z1.z2.s  ;
wire _2933_ ;
wire _2513_ ;
wire _3051_ ;
wire _2742_ ;
wire _2322_ ;
wire _8_ ;
wire _924_ ;
wire _504_ ;
wire _2971_ ;
wire _2551_ ;
wire _2131_ ;
wire _1822_ ;
wire _1402_ ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _2780_ ;
wire _2360_ ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire \z4.z2.z1.z2.s  ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2836_ ;
wire _2416_ ;
wire \z3.z3.z4.z1.s  ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire \z1.z3.z2.z1.a  ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire \z2.z4.z2.z2.c  ;
wire _1916_ ;
wire \z1.z1.z4.z2.a  ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire \z2.z1.z2.z1.c  ;
wire _580_ ;
wire _160_ ;
wire _2874_ ;
wire _2454_ ;
wire _2034_ ;
wire _1725_ ;
wire _1305_ ;
wire _636_ ;
wire _216_ ;
wire _2683_ ;
wire _2263_ ;
wire _3048_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _2492_ ;
wire _2072_ ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _2968_ ;
wire _2548_ ;
wire _2128_ ;
wire \z3.z4.z2.z1.a  ;
wire _1819_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire \z3.z2.z4.z2.a  ;
wire _483_ ;
wire _2777_ ;
wire _2357_ ;
wire _1628_ ;
wire _1208_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _1381_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _11_ ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _768_ ;
wire _348_ ;
wire _1190_ ;
wire _2395_ ;
wire [3:0] \z2.z2.q3  ;
wire _1666_ ;
wire _1246_ ;
wire \z2.z4.z4.z1.b  ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire \z4.z1.z2.z2.s  ;
wire _1284_ ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _3010_ ;
wire \z1.z2.z3.z1.a  ;
wire _2701_ ;
wire _1093_ ;
wire \z2.z3.z3.z2.c  ;
wire _2298_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2930_ ;
wire _2510_ ;
wire _1798_ ;
wire _1378_ ;
wire _289_ ;
wire _5_ ;
wire [7:0] \z3.q2  ;
wire _921_ ;
wire _501_ ;
wire _1187_ ;
wire \z4.z3.z1.z1.b  ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire \z2.z4.z1.z2.s  ;
wire \z3.z3.z3.z1.a  ;
wire \z2.z1.z1.z1.s  ;
wire _46_ ;
wire _2833_ ;
wire _2413_ ;
wire _2642_ ;
wire _2222_ ;
wire _3007_ ;
wire _1913_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _2871_ ;
wire _2451_ ;
wire _2031_ ;
wire _1722_ ;
wire _1302_ ;
wire _633_ ;
wire _213_ ;
wire _2927_ ;
wire _2507_ ;
wire _2680_ ;
wire _2260_ ;
wire _3045_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire \z4.z2.z1.z1.s  ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire _918_ ;
wire _1760_ ;
wire _1340_ ;
wire \z1.z4.z4.z2.a  ;
wire _671_ ;
wire _251_ ;
wire _2965_ ;
wire _2545_ ;
wire _2125_ ;
wire [3:0] \z3.z4.q1  ;
wire \z2.z4.z2.z1.c  ;
wire _1816_ ;
wire \z1.z1.z4.z1.a  ;
wire _727_ ;
wire _307_ ;
wire \z2.z2.z4.z2.c  ;
wire _480_ ;
wire _2774_ ;
wire _2354_ ;
wire _1625_ ;
wire _1205_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _2583_ ;
wire _2163_ ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire \z1.z2.z1.z1.b  ;
wire _2392_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2868_ ;
wire _2448_ ;
wire _2028_ ;
wire \z4.z2.z2.z1.b  ;
wire _1719_ ;
wire \z2.z3.z2.z2.s  ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire \z3.z2.z4.z1.a  ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire _1948_ ;
wire _1528_ ;
wire _1108_ ;
wire _859_ ;
wire _439_ ;
wire _1281_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire \z3.z3.z1.z2.a  ;
wire _1757_ ;
wire _1337_ ;
wire _668_ ;
wire _248_ ;
wire _1090_ ;
wire _2295_ ;
wire \z4.z1.z1.z2.c  ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _1795_ ;
wire _1375_ ;
wire \z4.z4.z2.z2.s  ;
wire _286_ ;
wire _2_ ;
wire \z4.z1.z2.z1.s  ;
wire _1184_ ;
wire _2389_ ;
wire _2601_ ;
wire \z2.z3.z3.z1.c  ;
wire _2198_ ;
wire _43_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2830_ ;
wire _2410_ ;
wire _1698_ ;
wire _1278_ ;
wire _189_ ;
wire _3004_ ;
wire _1910_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire \z1.z1.z2.z1.b  ;
wire _1087_ ;
wire _630_ ;
wire _210_ ;
wire _2924_ ;
wire _2504_ ;
wire \z2.z4.z1.z1.s  ;
wire [3:0] \z1.z3.q1  ;
wire \z4.z1.z3.z1.b  ;
wire _3042_ ;
wire \z2.z2.z3.z2.s  ;
wire _2733_ ;
wire _2313_ ;
wire _915_ ;
wire _2962_ ;
wire _2542_ ;
wire _2122_ ;
wire \z3.z2.z2.z2.a  ;
wire _1813_ ;
wire _724_ ;
wire _304_ ;
wire _2771_ ;
wire _2351_ ;
wire _1622_ ;
wire _1202_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _2827_ ;
wire _2407_ ;
wire [3:0] \z4.z1.q1  ;
wire _2580_ ;
wire _2160_ ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire \z4.z3.z3.z2.s  ;
wire _2636_ ;
wire _2216_ ;
wire _1907_ ;
wire _818_ ;
wire _78_ ;
wire _1660_ ;
wire _1240_ ;
wire \z1.z4.z4.z1.a  ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2865_ ;
wire _2445_ ;
wire _2025_ ;
wire _1716_ ;
wire _627_ ;
wire _207_ ;
wire \z2.z2.z4.z1.c  ;
wire _380_ ;
wire _2674_ ;
wire _2254_ ;
wire _3039_ ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire [15:0] \z1.q3  ;
wire _2483_ ;
wire _2063_ ;
wire \z2.z3.z1.z2.c  ;
wire _1754_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _2959_ ;
wire _2539_ ;
wire _2119_ ;
wire _2292_ ;
wire _1983_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire _1619_ ;
wire \z2.z3.z2.z1.s  ;
wire _1792_ ;
wire _1372_ ;
wire _283_ ;
wire _2997_ ;
wire _2577_ ;
wire _2157_ ;
wire \z2.z1.z4.z2.s  ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _759_ ;
wire _339_ ;
wire _1181_ ;
wire _2386_ ;
wire \z3.z3.z1.z1.a  ;
wire \z4.z4.z1.z2.c  ;
wire _1657_ ;
wire _1237_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire \z3.z1.z3.z2.a  ;
wire _2195_ ;
wire \z4.z1.z1.z1.c  ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire _1695_ ;
wire _1275_ ;
wire \z4.z4.z2.z1.s  ;
wire _186_ ;
wire _3001_ ;
wire [3:0] \z3.z2.q2  ;
wire \z4.z2.z4.z2.s  ;
wire _1084_ ;
wire _2289_ ;
wire _2921_ ;
wire _2501_ ;
wire _2098_ ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire _912_ ;
wire _1598_ ;
wire _1178_ ;
wire \z2.z2.z2.z2.c  ;
wire \z1.z4.z2.z1.b  ;
wire _1810_ ;
wire _721_ ;
wire _301_ ;
wire \z4.z4.z3.z1.b  ;
wire _37_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2824_ ;
wire _2404_ ;
wire \z2.z2.z3.z1.s  ;
wire _2633_ ;
wire _2213_ ;
wire _1904_ ;
wire _815_ ;
wire _75_ ;
wire _2862_ ;
wire _2442_ ;
wire _2022_ ;
wire \z3.z2.z2.z1.a  ;
wire _1713_ ;
wire \z4.z3.z2.z2.c  ;
wire _624_ ;
wire _204_ ;
wire _2918_ ;
wire _2671_ ;
wire _2251_ ;
wire _3036_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire [7:0] \z1.q0  ;
wire _2727_ ;
wire _2307_ ;
wire _2480_ ;
wire _2060_ ;
wire _909_ ;
wire _1751_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire \z4.z3.z3.z1.s  ;
wire _2956_ ;
wire _2536_ ;
wire _2116_ ;
wire _1807_ ;
wire _718_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _1616_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _2994_ ;
wire _2574_ ;
wire _2154_ ;
wire _1845_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _2383_ ;
wire \z2.z3.z1.z1.c  ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2859_ ;
wire _2439_ ;
wire _2019_ ;
wire \z2.z1.z3.z2.c  ;
wire \z1.z3.z3.z1.b  ;
wire _2192_ ;
wire [3:0] \z1.z1.q2  ;
wire _1883_ ;
wire _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire \z4.z3.z4.z1.b  ;
wire _1939_ ;
wire _1519_ ;
wire \z2.z4.z4.z2.s  ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _2897_ ;
wire _2477_ ;
wire _2057_ ;
wire \z2.z1.z4.z1.s  ;
wire [3:0] \z4.z4.q2  ;
wire _1748_ ;
wire _1328_ ;
wire _659_ ;
wire _239_ ;
wire _1081_ ;
wire _2286_ ;
wire \z3.z4.z3.z2.a  ;
wire \z4.z4.z1.z1.c  ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _888_ ;
wire _468_ ;
wire \z3.z1.z3.z1.a  ;
wire _2095_ ;
wire \z4.z2.z3.z2.c  ;
wire _1786_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _1595_ ;
wire _1175_ ;
wire \z4.z2.z4.z1.s  ;
wire _2189_ ;
wire _34_ ;
wire _2821_ ;
wire _2401_ ;
wire \z4.z3.z1.z2.s  ;
wire _1689_ ;
wire _1269_ ;
wire _2630_ ;
wire _2210_ ;
wire _1901_ ;
wire _812_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire \z2.z2.z2.z1.c  ;
wire _1710_ ;
wire _621_ ;
wire _201_ ;
wire _2915_ ;
wire \z1.z2.z4.z1.b  ;
wire _3033_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _906_ ;
wire _2953_ ;
wire _2533_ ;
wire _2113_ ;
wire _1804_ ;
wire _715_ ;
wire _2762_ ;
wire _2342_ ;
wire \z3.z3.z4.z2.a  ;
wire _1613_ ;
wire \z4.z3.z2.z1.c  ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2818_ ;
wire _2991_ ;
wire _2571_ ;
wire _2151_ ;
wire \z4.z1.z4.z2.c  ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire _2627_ ;
wire _2207_ ;
wire _2380_ ;
wire _809_ ;
wire _69_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2856_ ;
wire _2436_ ;
wire _2016_ ;
wire [3:0] \z2.z3.q2  ;
wire \z3.z1.z1.z1.b  ;
wire _1707_ ;
wire _618_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire \z1.z2.z1.z2.s  ;
wire _1936_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _2894_ ;
wire _2474_ ;
wire _2054_ ;
wire \z4.z2.z2.z2.s  ;
wire _1745_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _2283_ ;
wire \z2.z4.z3.z2.c  ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _2759_ ;
wire _2339_ ;
wire \z2.z1.z3.z1.c  ;
wire _2092_ ;
wire _1783_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _2988_ ;
wire _2568_ ;
wire _2148_ ;
wire _1839_ ;
wire _1419_ ;
wire \z2.z4.z4.z1.s  ;
wire _1592_ ;
wire _1172_ ;
wire _2797_ ;
wire _2377_ ;
wire [7:0] \z4.q1  ;
wire _1648_ ;
wire _1228_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _2186_ ;
wire \z3.z4.z3.z1.a  ;
wire _31_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _788_ ;
wire _368_ ;
wire \z4.z2.z3.z1.c  ;
wire _1686_ ;
wire _1266_ ;
wire _597_ ;
wire _177_ ;
wire _1495_ ;
wire _1075_ ;
wire _2912_ ;
wire _2089_ ;
wire _3030_ ;
wire _2721_ ;
wire _2301_ ;
wire \z1.z1.z2.z2.s  ;
wire [3:0] \z1.z4.q3  ;
wire \z4.z3.z1.z1.s  ;
wire _903_ ;
wire _1589_ ;
wire _1169_ ;
wire _2950_ ;
wire _2530_ ;
wire _2110_ ;
wire \z4.z1.z3.z2.s  ;
wire _1801_ ;
wire \z2.z1.z1.z2.a  ;
wire _712_ ;
wire _1398_ ;
wire \z2.z3.z4.z2.c  ;
wire _28_ ;
wire _1610_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire _750_ ;
wire _330_ ;
wire _2624_ ;
wire _2204_ ;
wire [3:0] \z4.z2.q3  ;
wire \z1.z3.z1.z1.b  ;
wire _806_ ;
wire _66_ ;
wire _2853_ ;
wire _2433_ ;
wire _2013_ ;
wire _1704_ ;
wire _615_ ;
wire _2909_ ;
wire \z4.z2.z1.z2.a  ;
wire _2662_ ;
wire _2242_ ;
wire _3027_ ;
wire \z3.z3.z4.z1.a  ;
wire _1933_ ;
wire _1513_ ;
wire \z4.z4.z4.z2.c  ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire _2891_ ;
wire _2471_ ;
wire _2051_ ;
wire \z4.z1.z4.z1.c  ;
wire _1742_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire _2947_ ;
wire _2527_ ;
wire _2107_ ;
wire _2280_ ;
wire _709_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire \z3.z4.z1.z1.b  ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire _1607_ ;
wire _938_ ;
wire _518_ ;
wire _1780_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _2985_ ;
wire _2565_ ;
wire _2145_ ;
wire \z1.z2.z1.z1.s  ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _2794_ ;
wire _2374_ ;
wire \z4.z2.z2.z1.s  ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _2183_ ;
wire \z2.z4.z3.z1.c  ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _2888_ ;
wire _2468_ ;
wire _2048_ ;
wire _1739_ ;
wire _1319_ ;
wire _1492_ ;
wire _1072_ ;
wire _2697_ ;
wire _2277_ ;
wire \z1.z2.z2.z1.b  ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _879_ ;
wire _459_ ;
wire _2086_ ;
wire \z4.z1.z2.z2.a  ;
wire _1777_ ;
wire _1357_ ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire \z1.z1.z1.z2.c  ;
wire _1395_ ;
wire [3:0] \z2.z1.q3  ;
wire _25_ ;
wire \z3.z3.z2.z1.b  ;
wire _2812_ ;
wire \z1.z4.z2.z2.s  ;
wire _2621_ ;
wire _2201_ ;
wire \z1.z1.z2.z1.s  ;
wire \z4.z4.z3.z2.s  ;
wire _803_ ;
wire _63_ ;
wire \z2.z4.z1.z2.a  ;
wire _1489_ ;
wire _1069_ ;
wire _2850_ ;
wire _2430_ ;
wire _2010_ ;
wire \z4.z1.z3.z1.s  ;
wire _1701_ ;
wire \z2.z1.z1.z1.a  ;
wire _612_ ;
wire _2906_ ;
wire \z3.z2.z1.z2.c  ;
wire _1298_ ;
wire _3024_ ;
wire \z2.z3.z4.z1.c  ;
wire _1930_ ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _650_ ;
wire _230_ ;
wire _2944_ ;
wire _2524_ ;
wire _2104_ ;
wire [7:0] \z2.q2  ;
wire _706_ ;
wire _2753_ ;
wire _2333_ ;
wire \z1.z1.z3.z1.b  ;
wire _1604_ ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire \z4.z2.z1.z1.a  ;
wire _2982_ ;
wire _2562_ ;
wire _2142_ ;
wire _1833_ ;
wire _1413_ ;
wire \z4.z4.z4.z1.c  ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _2791_ ;
wire _2371_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _2847_ ;
wire _2427_ ;
wire _2007_ ;
wire _2180_ ;
wire _609_ ;
wire _1871_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire \z3.z2.z3.z1.b  ;
wire _1927_ ;
wire _1507_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _2885_ ;
wire _2465_ ;
wire _2045_ ;
wire \z1.z3.z3.z2.s  ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _2694_ ;
wire _2274_ ;
wire \z4.z3.z4.z2.s  ;
wire _1965_ ;
wire _1545_ ;
wire _1125_ ;
wire \z2.z3.z2.z2.a  ;
wire _876_ ;
wire _456_ ;
wire [3:0] \z3.z3.q1  ;
wire _2083_ ;
wire \z3.z1.z2.z2.c  ;
wire _1774_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _2979_ ;
wire _2559_ ;
wire _2139_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire _1639_ ;
wire _1219_ ;
wire _1392_ ;
wire _2597_ ;
wire _2177_ ;
wire _22_ ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _779_ ;
wire _359_ ;
wire \z4.z4.z2.z2.a  ;

NOR2X1 _3054_ (
    .A(q1[0]),
    .B(q0[8]),
    .Y(_415_)
);

NAND2X1 _3055_ (
    .A(q1[0]),
    .B(q0[8]),
    .Y(_416_)
);

INVX1 _3056_ (
    .A(_416_),
    .Y(_417_)
);

OR2X2 _3057_ (
    .A(_417_),
    .B(_415_),
    .Y(_418_)
);

INVX1 _3058_ (
    .A(_418_),
    .Y(_419_)
);

AND2X2 _3059_ (
    .A(_419_),
    .B(q2[0]),
    .Y(_420_)
);

NOR2X1 _3060_ (
    .A(q2[0]),
    .B(_419_),
    .Y(_421_)
);

NOR2X1 _3061_ (
    .A(_421_),
    .B(_420_),
    .Y(_3053_[8])
);

NAND2X1 _3062_ (
    .A(\z2.z1.z1.z1.s ),
    .B(q0[9]),
    .Y(_422_)
);

OR2X2 _3063_ (
    .A(\z2.z1.z1.z1.s ),
    .B(q0[9]),
    .Y(_423_)
);

NAND2X1 _3064_ (
    .A(_422_),
    .B(_423_),
    .Y(_424_)
);

NOR2X1 _3065_ (
    .A(_416_),
    .B(_424_),
    .Y(_425_)
);

AOI21X1 _3066_ (
    .A(_422_),
    .B(_423_),
    .C(_417_),
    .Y(_426_)
);

NOR2X1 _3067_ (
    .A(_426_),
    .B(_425_),
    .Y(_427_)
);

NAND2X1 _3068_ (
    .A(\z3.z1.z1.z1.s ),
    .B(_427_),
    .Y(_428_)
);

OR2X2 _3069_ (
    .A(_427_),
    .B(\z3.z1.z1.z1.s ),
    .Y(_429_)
);

NAND3X1 _3070_ (
    .A(_420_),
    .B(_428_),
    .C(_429_),
    .Y(_430_)
);

INVX1 _3071_ (
    .A(_430_),
    .Y(_431_)
);

INVX1 _3072_ (
    .A(_428_),
    .Y(_432_)
);

NOR2X1 _3073_ (
    .A(\z2.z1.z1.z1.s ),
    .B(q0[9]),
    .Y(_0_)
);

OAI21X1 _3074_ (
    .A(_416_),
    .B(_0_),
    .C(_422_),
    .Y(_1_)
);

NOR2X1 _3075_ (
    .A(q1[2]),
    .B(q0[10]),
    .Y(_2_)
);

AND2X2 _3076_ (
    .A(q1[2]),
    .B(q0[10]),
    .Y(_3_)
);

NOR2X1 _3077_ (
    .A(_2_),
    .B(_3_),
    .Y(_4_)
);

NAND2X1 _3078_ (
    .A(_1_),
    .B(_4_),
    .Y(_5_)
);

OR2X2 _3079_ (
    .A(_4_),
    .B(_1_),
    .Y(_6_)
);

NAND3X1 _3080_ (
    .A(q2[2]),
    .B(_5_),
    .C(_6_),
    .Y(_7_)
);

INVX1 _3081_ (
    .A(q2[2]),
    .Y(_8_)
);

NAND2X1 _3082_ (
    .A(_5_),
    .B(_6_),
    .Y(_9_)
);

NAND2X1 _3083_ (
    .A(_8_),
    .B(_9_),
    .Y(_10_)
);

AOI21X1 _3084_ (
    .A(_7_),
    .B(_10_),
    .C(_432_),
    .Y(_11_)
);

NAND3X1 _3085_ (
    .A(_7_),
    .B(_10_),
    .C(_432_),
    .Y(_12_)
);

INVX1 _3086_ (
    .A(_12_),
    .Y(_13_)
);

NOR2X1 _3087_ (
    .A(_11_),
    .B(_13_),
    .Y(_14_)
);

NAND2X1 _3088_ (
    .A(_431_),
    .B(_14_),
    .Y(_15_)
);

INVX1 _3089_ (
    .A(_15_),
    .Y(_16_)
);

NOR2X1 _3090_ (
    .A(_431_),
    .B(_14_),
    .Y(_17_)
);

NOR2X1 _3091_ (
    .A(_17_),
    .B(_16_),
    .Y(_3053_[10])
);

NAND2X1 _3092_ (
    .A(q1[2]),
    .B(q0[10]),
    .Y(_18_)
);

INVX1 _3093_ (
    .A(q1[3]),
    .Y(_19_)
);

NAND2X1 _3094_ (
    .A(q0[11]),
    .B(_19_),
    .Y(_20_)
);

INVX1 _3095_ (
    .A(q0[11]),
    .Y(_21_)
);

NAND2X1 _3096_ (
    .A(q1[3]),
    .B(_21_),
    .Y(_22_)
);

NAND2X1 _3097_ (
    .A(_20_),
    .B(_22_),
    .Y(_23_)
);

NAND3X1 _3098_ (
    .A(_18_),
    .B(_23_),
    .C(_5_),
    .Y(_24_)
);

NAND2X1 _3099_ (
    .A(_18_),
    .B(_5_),
    .Y(_25_)
);

NAND3X1 _3100_ (
    .A(_20_),
    .B(_22_),
    .C(_25_),
    .Y(_26_)
);

NAND2X1 _3101_ (
    .A(_24_),
    .B(_26_),
    .Y(_27_)
);

NAND2X1 _3102_ (
    .A(q2[3]),
    .B(_27_),
    .Y(_28_)
);

INVX1 _3103_ (
    .A(q2[3]),
    .Y(_29_)
);

NAND3X1 _3104_ (
    .A(_29_),
    .B(_24_),
    .C(_26_),
    .Y(_30_)
);

NAND2X1 _3105_ (
    .A(_30_),
    .B(_28_),
    .Y(_31_)
);

OAI21X1 _3106_ (
    .A(_8_),
    .B(_9_),
    .C(_31_),
    .Y(_32_)
);

INVX1 _3107_ (
    .A(_7_),
    .Y(_33_)
);

NAND3X1 _3108_ (
    .A(_33_),
    .B(_30_),
    .C(_28_),
    .Y(_34_)
);

NAND2X1 _3109_ (
    .A(_34_),
    .B(_32_),
    .Y(_35_)
);

OAI21X1 _3110_ (
    .A(_13_),
    .B(_16_),
    .C(_35_),
    .Y(_36_)
);

OAI21X1 _3111_ (
    .A(_430_),
    .B(_11_),
    .C(_12_),
    .Y(_37_)
);

OR2X2 _3112_ (
    .A(_35_),
    .B(_37_),
    .Y(_38_)
);

NAND2X1 _3113_ (
    .A(_38_),
    .B(_36_),
    .Y(_3053_[11])
);

INVX1 _3114_ (
    .A(_34_),
    .Y(_39_)
);

AOI21X1 _3115_ (
    .A(_37_),
    .B(_32_),
    .C(_39_),
    .Y(_40_)
);

INVX1 _3116_ (
    .A(_28_),
    .Y(_41_)
);

INVX1 _3117_ (
    .A(q2[4]),
    .Y(_42_)
);

NAND3X1 _3118_ (
    .A(_1_),
    .B(_23_),
    .C(_4_),
    .Y(_43_)
);

AOI21X1 _3119_ (
    .A(_19_),
    .B(_21_),
    .C(_18_),
    .Y(_44_)
);

AOI21X1 _3120_ (
    .A(q1[3]),
    .B(q0[11]),
    .C(_44_),
    .Y(_45_)
);

INVX1 _3121_ (
    .A(q1[4]),
    .Y(_46_)
);

INVX1 _3122_ (
    .A(q0[12]),
    .Y(_47_)
);

NAND2X1 _3123_ (
    .A(_46_),
    .B(_47_),
    .Y(_48_)
);

NAND2X1 _3124_ (
    .A(q1[4]),
    .B(q0[12]),
    .Y(_49_)
);

NAND2X1 _3125_ (
    .A(_49_),
    .B(_48_),
    .Y(_50_)
);

AOI21X1 _3126_ (
    .A(_43_),
    .B(_45_),
    .C(_50_),
    .Y(_51_)
);

INVX1 _3127_ (
    .A(_51_),
    .Y(_52_)
);

AND2X2 _3128_ (
    .A(_43_),
    .B(_45_),
    .Y(_53_)
);

NOR2X1 _3129_ (
    .A(q1[4]),
    .B(q0[12]),
    .Y(_54_)
);

AND2X2 _3130_ (
    .A(q1[4]),
    .B(q0[12]),
    .Y(_55_)
);

OAI21X1 _3131_ (
    .A(_54_),
    .B(_55_),
    .C(_53_),
    .Y(_56_)
);

NAND2X1 _3132_ (
    .A(_52_),
    .B(_56_),
    .Y(_57_)
);

OR2X2 _3133_ (
    .A(_57_),
    .B(_42_),
    .Y(_58_)
);

AOI21X1 _3134_ (
    .A(_56_),
    .B(_52_),
    .C(q2[4]),
    .Y(_59_)
);

INVX1 _3135_ (
    .A(_59_),
    .Y(_60_)
);

NAND3X1 _3136_ (
    .A(_41_),
    .B(_60_),
    .C(_58_),
    .Y(_61_)
);

NOR2X1 _3137_ (
    .A(_42_),
    .B(_57_),
    .Y(_62_)
);

OAI21X1 _3138_ (
    .A(_59_),
    .B(_62_),
    .C(_28_),
    .Y(_63_)
);

NAND2X1 _3139_ (
    .A(_63_),
    .B(_61_),
    .Y(_64_)
);

NOR2X1 _3140_ (
    .A(_64_),
    .B(_40_),
    .Y(_65_)
);

AND2X2 _3141_ (
    .A(_40_),
    .B(_64_),
    .Y(_66_)
);

NOR2X1 _3142_ (
    .A(_65_),
    .B(_66_),
    .Y(_3053_[12])
);

OAI21X1 _3143_ (
    .A(_64_),
    .B(_40_),
    .C(_61_),
    .Y(_67_)
);

INVX1 _3144_ (
    .A(q2[5]),
    .Y(_68_)
);

NAND2X1 _3145_ (
    .A(q1[5]),
    .B(q0[13]),
    .Y(_69_)
);

INVX1 _3146_ (
    .A(q1[5]),
    .Y(_70_)
);

INVX1 _3147_ (
    .A(q0[13]),
    .Y(_71_)
);

NAND2X1 _3148_ (
    .A(_70_),
    .B(_71_),
    .Y(_72_)
);

NAND2X1 _3149_ (
    .A(_69_),
    .B(_72_),
    .Y(_73_)
);

OAI21X1 _3150_ (
    .A(_46_),
    .B(_47_),
    .C(_73_),
    .Y(_74_)
);

NAND2X1 _3151_ (
    .A(q0[13]),
    .B(_70_),
    .Y(_75_)
);

NAND2X1 _3152_ (
    .A(q1[5]),
    .B(_71_),
    .Y(_76_)
);

NAND2X1 _3153_ (
    .A(_75_),
    .B(_76_),
    .Y(_77_)
);

OAI21X1 _3154_ (
    .A(_55_),
    .B(_51_),
    .C(_77_),
    .Y(_78_)
);

OAI21X1 _3155_ (
    .A(_51_),
    .B(_74_),
    .C(_78_),
    .Y(_79_)
);

NOR2X1 _3156_ (
    .A(_68_),
    .B(_79_),
    .Y(_80_)
);

AND2X2 _3157_ (
    .A(_79_),
    .B(_68_),
    .Y(_81_)
);

OAI21X1 _3158_ (
    .A(_80_),
    .B(_81_),
    .C(_58_),
    .Y(_82_)
);

OR2X2 _3159_ (
    .A(_79_),
    .B(_68_),
    .Y(_83_)
);

NAND2X1 _3160_ (
    .A(_68_),
    .B(_79_),
    .Y(_84_)
);

NAND3X1 _3161_ (
    .A(_62_),
    .B(_84_),
    .C(_83_),
    .Y(_85_)
);

NAND2X1 _3162_ (
    .A(_82_),
    .B(_85_),
    .Y(_86_)
);

NAND2X1 _3163_ (
    .A(_86_),
    .B(_67_),
    .Y(_87_)
);

OR2X2 _3164_ (
    .A(_67_),
    .B(_86_),
    .Y(_88_)
);

NAND2X1 _3165_ (
    .A(_87_),
    .B(_88_),
    .Y(_3053_[13])
);

NOR3X1 _3166_ (
    .A(_64_),
    .B(_40_),
    .C(_86_),
    .Y(_89_)
);

OAI21X1 _3167_ (
    .A(_61_),
    .B(_86_),
    .C(_85_),
    .Y(_90_)
);

NOR2X1 _3168_ (
    .A(_54_),
    .B(_55_),
    .Y(_91_)
);

NAND2X1 _3169_ (
    .A(_77_),
    .B(_91_),
    .Y(_92_)
);

AOI21X1 _3170_ (
    .A(_43_),
    .B(_45_),
    .C(_92_),
    .Y(_93_)
);

NOR2X1 _3171_ (
    .A(q1[5]),
    .B(q0[13]),
    .Y(_94_)
);

OAI21X1 _3172_ (
    .A(_49_),
    .B(_94_),
    .C(_69_),
    .Y(_95_)
);

NOR2X1 _3173_ (
    .A(q1[6]),
    .B(q0[14]),
    .Y(_96_)
);

AND2X2 _3174_ (
    .A(q1[6]),
    .B(q0[14]),
    .Y(_97_)
);

NOR2X1 _3175_ (
    .A(_96_),
    .B(_97_),
    .Y(_98_)
);

OAI21X1 _3176_ (
    .A(_95_),
    .B(_93_),
    .C(_98_),
    .Y(_99_)
);

INVX1 _3177_ (
    .A(q1[6]),
    .Y(_100_)
);

INVX1 _3178_ (
    .A(q0[14]),
    .Y(_101_)
);

NAND2X1 _3179_ (
    .A(_100_),
    .B(_101_),
    .Y(_102_)
);

NAND2X1 _3180_ (
    .A(q1[6]),
    .B(q0[14]),
    .Y(_103_)
);

NAND2X1 _3181_ (
    .A(_103_),
    .B(_102_),
    .Y(_104_)
);

NAND3X1 _3182_ (
    .A(_69_),
    .B(_104_),
    .C(_78_),
    .Y(_105_)
);

NAND3X1 _3183_ (
    .A(q2[6]),
    .B(_99_),
    .C(_105_),
    .Y(_106_)
);

INVX1 _3184_ (
    .A(q2[6]),
    .Y(_107_)
);

NAND2X1 _3185_ (
    .A(_99_),
    .B(_105_),
    .Y(_108_)
);

NAND2X1 _3186_ (
    .A(_107_),
    .B(_108_),
    .Y(_109_)
);

NAND2X1 _3187_ (
    .A(_106_),
    .B(_109_),
    .Y(_110_)
);

OR2X2 _3188_ (
    .A(_110_),
    .B(_83_),
    .Y(_111_)
);

OAI21X1 _3189_ (
    .A(_68_),
    .B(_79_),
    .C(_110_),
    .Y(_112_)
);

AND2X2 _3190_ (
    .A(_111_),
    .B(_112_),
    .Y(_113_)
);

OAI21X1 _3191_ (
    .A(_90_),
    .B(_89_),
    .C(_113_),
    .Y(_114_)
);

INVX1 _3192_ (
    .A(_85_),
    .Y(_115_)
);

AOI21X1 _3193_ (
    .A(_67_),
    .B(_82_),
    .C(_115_),
    .Y(_116_)
);

NAND2X1 _3194_ (
    .A(_112_),
    .B(_111_),
    .Y(_117_)
);

NAND2X1 _3195_ (
    .A(_117_),
    .B(_116_),
    .Y(_118_)
);

AND2X2 _3196_ (
    .A(_118_),
    .B(_114_),
    .Y(_3053_[14])
);

OAI21X1 _3197_ (
    .A(_117_),
    .B(_116_),
    .C(_111_),
    .Y(_119_)
);

OAI21X1 _3198_ (
    .A(_100_),
    .B(_101_),
    .C(_99_),
    .Y(_120_)
);

INVX1 _3199_ (
    .A(q1[7]),
    .Y(_121_)
);

NAND2X1 _3200_ (
    .A(q0[15]),
    .B(_121_),
    .Y(_122_)
);

INVX1 _3201_ (
    .A(q0[15]),
    .Y(_123_)
);

NAND2X1 _3202_ (
    .A(q1[7]),
    .B(_123_),
    .Y(_124_)
);

NAND2X1 _3203_ (
    .A(_122_),
    .B(_124_),
    .Y(_125_)
);

NAND2X1 _3204_ (
    .A(_125_),
    .B(_120_),
    .Y(_126_)
);

OR2X2 _3205_ (
    .A(_120_),
    .B(_125_),
    .Y(_127_)
);

NAND3X1 _3206_ (
    .A(q2[7]),
    .B(_126_),
    .C(_127_),
    .Y(_128_)
);

INVX1 _3207_ (
    .A(q2[7]),
    .Y(_129_)
);

NAND2X1 _3208_ (
    .A(q1[7]),
    .B(q0[15]),
    .Y(_130_)
);

NAND2X1 _3209_ (
    .A(_121_),
    .B(_123_),
    .Y(_131_)
);

NAND2X1 _3210_ (
    .A(_130_),
    .B(_131_),
    .Y(_132_)
);

NAND2X1 _3211_ (
    .A(_132_),
    .B(_120_),
    .Y(_133_)
);

OR2X2 _3212_ (
    .A(_120_),
    .B(_132_),
    .Y(_134_)
);

NAND3X1 _3213_ (
    .A(_129_),
    .B(_133_),
    .C(_134_),
    .Y(_135_)
);

NAND2X1 _3214_ (
    .A(_128_),
    .B(_135_),
    .Y(_136_)
);

OAI21X1 _3215_ (
    .A(_107_),
    .B(_108_),
    .C(_136_),
    .Y(_137_)
);

INVX1 _3216_ (
    .A(_106_),
    .Y(_138_)
);

NAND3X1 _3217_ (
    .A(_138_),
    .B(_128_),
    .C(_135_),
    .Y(_139_)
);

NAND2X1 _3218_ (
    .A(_139_),
    .B(_137_),
    .Y(_140_)
);

OR2X2 _3219_ (
    .A(_119_),
    .B(_140_),
    .Y(_141_)
);

NAND2X1 _3220_ (
    .A(_140_),
    .B(_119_),
    .Y(_142_)
);

NAND2X1 _3221_ (
    .A(_142_),
    .B(_141_),
    .Y(_3053_[15])
);

AOI21X1 _3222_ (
    .A(_134_),
    .B(_133_),
    .C(_129_),
    .Y(_143_)
);

NOR2X1 _3223_ (
    .A(_50_),
    .B(_73_),
    .Y(_144_)
);

NOR2X1 _3224_ (
    .A(_104_),
    .B(_132_),
    .Y(_145_)
);

NAND2X1 _3225_ (
    .A(_144_),
    .B(_145_),
    .Y(_146_)
);

OAI21X1 _3226_ (
    .A(q1[7]),
    .B(q0[15]),
    .C(_97_),
    .Y(_147_)
);

OAI21X1 _3227_ (
    .A(_121_),
    .B(_123_),
    .C(_147_),
    .Y(_148_)
);

AOI21X1 _3228_ (
    .A(_145_),
    .B(_95_),
    .C(_148_),
    .Y(_149_)
);

OAI21X1 _3229_ (
    .A(_146_),
    .B(_53_),
    .C(_149_),
    .Y(_150_)
);

NAND2X1 _3230_ (
    .A(q1[8]),
    .B(_150_),
    .Y(_151_)
);

INVX1 _3231_ (
    .A(q1[8]),
    .Y(_152_)
);

NAND2X1 _3232_ (
    .A(_45_),
    .B(_43_),
    .Y(_153_)
);

NAND2X1 _3233_ (
    .A(_125_),
    .B(_98_),
    .Y(_154_)
);

NOR2X1 _3234_ (
    .A(_92_),
    .B(_154_),
    .Y(_155_)
);

NAND3X1 _3235_ (
    .A(_95_),
    .B(_125_),
    .C(_98_),
    .Y(_156_)
);

NAND3X1 _3236_ (
    .A(_130_),
    .B(_147_),
    .C(_156_),
    .Y(_157_)
);

AOI21X1 _3237_ (
    .A(_155_),
    .B(_153_),
    .C(_157_),
    .Y(_158_)
);

NAND2X1 _3238_ (
    .A(_152_),
    .B(_158_),
    .Y(_159_)
);

NAND2X1 _3239_ (
    .A(q3[0]),
    .B(q2[8]),
    .Y(_160_)
);

INVX1 _3240_ (
    .A(q3[0]),
    .Y(_161_)
);

INVX1 _3241_ (
    .A(q2[8]),
    .Y(_162_)
);

NAND2X1 _3242_ (
    .A(_161_),
    .B(_162_),
    .Y(_163_)
);

NAND2X1 _3243_ (
    .A(_160_),
    .B(_163_),
    .Y(_164_)
);

INVX1 _3244_ (
    .A(_164_),
    .Y(_165_)
);

NAND3X1 _3245_ (
    .A(_165_),
    .B(_159_),
    .C(_151_),
    .Y(_166_)
);

NAND3X1 _3246_ (
    .A(_144_),
    .B(_145_),
    .C(_153_),
    .Y(_167_)
);

AOI21X1 _3247_ (
    .A(_167_),
    .B(_149_),
    .C(_152_),
    .Y(_168_)
);

INVX1 _3248_ (
    .A(_159_),
    .Y(_169_)
);

OAI21X1 _3249_ (
    .A(_168_),
    .B(_169_),
    .C(_164_),
    .Y(_170_)
);

NAND3X1 _3250_ (
    .A(_166_),
    .B(_170_),
    .C(_143_),
    .Y(_171_)
);

NAND2X1 _3251_ (
    .A(_166_),
    .B(_170_),
    .Y(_172_)
);

NAND2X1 _3252_ (
    .A(_128_),
    .B(_172_),
    .Y(_173_)
);

AND2X2 _3253_ (
    .A(_171_),
    .B(_173_),
    .Y(_174_)
);

AND2X2 _3254_ (
    .A(_111_),
    .B(_139_),
    .Y(_175_)
);

OAI21X1 _3255_ (
    .A(_117_),
    .B(_116_),
    .C(_175_),
    .Y(_176_)
);

NAND2X1 _3256_ (
    .A(_137_),
    .B(_176_),
    .Y(_177_)
);

NAND2X1 _3257_ (
    .A(_174_),
    .B(_177_),
    .Y(_178_)
);

INVX1 _3258_ (
    .A(_174_),
    .Y(_179_)
);

AOI22X1 _3259_ (
    .A(_106_),
    .B(_136_),
    .C(_114_),
    .D(_175_),
    .Y(_180_)
);

NAND2X1 _3260_ (
    .A(_179_),
    .B(_180_),
    .Y(_181_)
);

NAND2X1 _3261_ (
    .A(_181_),
    .B(_178_),
    .Y(_3053_[16])
);

OAI21X1 _3262_ (
    .A(_179_),
    .B(_177_),
    .C(_171_),
    .Y(_182_)
);

OAI21X1 _3263_ (
    .A(_161_),
    .B(_162_),
    .C(_166_),
    .Y(_183_)
);

NAND3X1 _3264_ (
    .A(q1[8]),
    .B(q1[9]),
    .C(_150_),
    .Y(_184_)
);

INVX1 _3265_ (
    .A(q1[9]),
    .Y(_185_)
);

OAI21X1 _3266_ (
    .A(_152_),
    .B(_158_),
    .C(_185_),
    .Y(_186_)
);

INVX1 _3267_ (
    .A(\z4.z1.z1.z1.s ),
    .Y(_187_)
);

INVX1 _3268_ (
    .A(q2[9]),
    .Y(_188_)
);

NAND2X1 _3269_ (
    .A(_187_),
    .B(_188_),
    .Y(_189_)
);

NAND2X1 _3270_ (
    .A(\z4.z1.z1.z1.s ),
    .B(q2[9]),
    .Y(_190_)
);

NAND2X1 _3271_ (
    .A(_190_),
    .B(_189_),
    .Y(_191_)
);

INVX1 _3272_ (
    .A(_191_),
    .Y(_192_)
);

NAND3X1 _3273_ (
    .A(_192_),
    .B(_184_),
    .C(_186_),
    .Y(_193_)
);

NAND2X1 _3274_ (
    .A(_184_),
    .B(_186_),
    .Y(_194_)
);

NAND2X1 _3275_ (
    .A(_191_),
    .B(_194_),
    .Y(_195_)
);

NAND3X1 _3276_ (
    .A(_193_),
    .B(_183_),
    .C(_195_),
    .Y(_196_)
);

INVX1 _3277_ (
    .A(_196_),
    .Y(_197_)
);

AOI21X1 _3278_ (
    .A(_195_),
    .B(_193_),
    .C(_183_),
    .Y(_198_)
);

NOR2X1 _3279_ (
    .A(_198_),
    .B(_197_),
    .Y(_199_)
);

OR2X2 _3280_ (
    .A(_182_),
    .B(_199_),
    .Y(_200_)
);

NAND2X1 _3281_ (
    .A(_199_),
    .B(_182_),
    .Y(_201_)
);

AND2X2 _3282_ (
    .A(_200_),
    .B(_201_),
    .Y(_3053_[17])
);

AOI21X1 _3283_ (
    .A(_171_),
    .B(_196_),
    .C(_198_),
    .Y(_202_)
);

INVX1 _3284_ (
    .A(_202_),
    .Y(_203_)
);

NAND2X1 _3285_ (
    .A(_199_),
    .B(_174_),
    .Y(_204_)
);

OAI21X1 _3286_ (
    .A(_204_),
    .B(_177_),
    .C(_203_),
    .Y(_205_)
);

OAI21X1 _3287_ (
    .A(_187_),
    .B(_188_),
    .C(_193_),
    .Y(_206_)
);

NAND3X1 _3288_ (
    .A(q1[9]),
    .B(q1[10]),
    .C(_168_),
    .Y(_207_)
);

INVX1 _3289_ (
    .A(q1[10]),
    .Y(_208_)
);

NAND2X1 _3290_ (
    .A(_208_),
    .B(_184_),
    .Y(_209_)
);

INVX1 _3291_ (
    .A(q3[2]),
    .Y(_210_)
);

INVX1 _3292_ (
    .A(q2[10]),
    .Y(_211_)
);

NAND2X1 _3293_ (
    .A(_210_),
    .B(_211_),
    .Y(_212_)
);

NAND2X1 _3294_ (
    .A(q3[2]),
    .B(q2[10]),
    .Y(_213_)
);

NAND2X1 _3295_ (
    .A(_213_),
    .B(_212_),
    .Y(_214_)
);

INVX1 _3296_ (
    .A(_214_),
    .Y(_215_)
);

NAND3X1 _3297_ (
    .A(_207_),
    .B(_215_),
    .C(_209_),
    .Y(_216_)
);

AOI21X1 _3298_ (
    .A(_209_),
    .B(_207_),
    .C(_215_),
    .Y(_217_)
);

INVX1 _3299_ (
    .A(_217_),
    .Y(_218_)
);

NAND3X1 _3300_ (
    .A(_206_),
    .B(_216_),
    .C(_218_),
    .Y(_219_)
);

INVX1 _3301_ (
    .A(_206_),
    .Y(_220_)
);

INVX1 _3302_ (
    .A(_216_),
    .Y(_221_)
);

OAI21X1 _3303_ (
    .A(_217_),
    .B(_221_),
    .C(_220_),
    .Y(_222_)
);

AND2X2 _3304_ (
    .A(_219_),
    .B(_222_),
    .Y(_223_)
);

NAND2X1 _3305_ (
    .A(_223_),
    .B(_205_),
    .Y(_224_)
);

OR2X2 _3306_ (
    .A(_205_),
    .B(_223_),
    .Y(_225_)
);

AND2X2 _3307_ (
    .A(_225_),
    .B(_224_),
    .Y(_3053_[18])
);

NAND2X1 _3308_ (
    .A(_219_),
    .B(_224_),
    .Y(_226_)
);

OAI21X1 _3309_ (
    .A(_210_),
    .B(_211_),
    .C(_216_),
    .Y(_227_)
);

NOR3X1 _3310_ (
    .A(_152_),
    .B(_185_),
    .C(_158_),
    .Y(_228_)
);

NAND3X1 _3311_ (
    .A(q1[10]),
    .B(q1[11]),
    .C(_228_),
    .Y(_229_)
);

INVX1 _3312_ (
    .A(q1[11]),
    .Y(_230_)
);

OAI21X1 _3313_ (
    .A(_208_),
    .B(_184_),
    .C(_230_),
    .Y(_231_)
);

NOR2X1 _3314_ (
    .A(q3[3]),
    .B(q2[11]),
    .Y(_232_)
);

INVX1 _3315_ (
    .A(q3[3]),
    .Y(_233_)
);

INVX1 _3316_ (
    .A(q2[11]),
    .Y(_234_)
);

NOR2X1 _3317_ (
    .A(_233_),
    .B(_234_),
    .Y(_235_)
);

NOR2X1 _3318_ (
    .A(_232_),
    .B(_235_),
    .Y(_236_)
);

NAND3X1 _3319_ (
    .A(_231_),
    .B(_236_),
    .C(_229_),
    .Y(_237_)
);

NAND2X1 _3320_ (
    .A(_231_),
    .B(_229_),
    .Y(_238_)
);

OAI21X1 _3321_ (
    .A(_232_),
    .B(_235_),
    .C(_238_),
    .Y(_239_)
);

NAND3X1 _3322_ (
    .A(_227_),
    .B(_237_),
    .C(_239_),
    .Y(_240_)
);

AND2X2 _3323_ (
    .A(_216_),
    .B(_213_),
    .Y(_241_)
);

INVX1 _3324_ (
    .A(_236_),
    .Y(_242_)
);

NAND3X1 _3325_ (
    .A(_231_),
    .B(_242_),
    .C(_229_),
    .Y(_243_)
);

NAND2X1 _3326_ (
    .A(_236_),
    .B(_238_),
    .Y(_244_)
);

NAND3X1 _3327_ (
    .A(_243_),
    .B(_241_),
    .C(_244_),
    .Y(_245_)
);

NAND2X1 _3328_ (
    .A(_245_),
    .B(_240_),
    .Y(_246_)
);

OR2X2 _3329_ (
    .A(_226_),
    .B(_246_),
    .Y(_247_)
);

NAND2X1 _3330_ (
    .A(_246_),
    .B(_226_),
    .Y(_248_)
);

NAND2X1 _3331_ (
    .A(_248_),
    .B(_247_),
    .Y(_3053_[19])
);

NAND2X1 _3332_ (
    .A(_222_),
    .B(_219_),
    .Y(_249_)
);

NOR3X1 _3333_ (
    .A(_249_),
    .B(_246_),
    .C(_204_),
    .Y(_250_)
);

AND2X2 _3334_ (
    .A(_240_),
    .B(_245_),
    .Y(_251_)
);

NAND3X1 _3335_ (
    .A(_202_),
    .B(_223_),
    .C(_251_),
    .Y(_252_)
);

INVX1 _3336_ (
    .A(_219_),
    .Y(_253_)
);

NAND2X1 _3337_ (
    .A(_253_),
    .B(_251_),
    .Y(_254_)
);

NAND3X1 _3338_ (
    .A(_240_),
    .B(_254_),
    .C(_252_),
    .Y(_255_)
);

AOI21X1 _3339_ (
    .A(_180_),
    .B(_250_),
    .C(_255_),
    .Y(_256_)
);

OAI21X1 _3340_ (
    .A(_233_),
    .B(_234_),
    .C(_237_),
    .Y(_257_)
);

NOR2X1 _3341_ (
    .A(_208_),
    .B(_184_),
    .Y(_258_)
);

NAND3X1 _3342_ (
    .A(q1[11]),
    .B(q1[12]),
    .C(_258_),
    .Y(_259_)
);

INVX1 _3343_ (
    .A(q1[12]),
    .Y(_260_)
);

OAI21X1 _3344_ (
    .A(_230_),
    .B(_207_),
    .C(_260_),
    .Y(_261_)
);

INVX1 _3345_ (
    .A(q3[4]),
    .Y(_262_)
);

INVX1 _3346_ (
    .A(q2[12]),
    .Y(_263_)
);

NAND2X1 _3347_ (
    .A(_262_),
    .B(_263_),
    .Y(_264_)
);

NAND2X1 _3348_ (
    .A(q3[4]),
    .B(q2[12]),
    .Y(_265_)
);

NAND2X1 _3349_ (
    .A(_265_),
    .B(_264_),
    .Y(_266_)
);

INVX1 _3350_ (
    .A(_266_),
    .Y(_267_)
);

NAND3X1 _3351_ (
    .A(_261_),
    .B(_267_),
    .C(_259_),
    .Y(_268_)
);

AOI21X1 _3352_ (
    .A(_259_),
    .B(_261_),
    .C(_267_),
    .Y(_269_)
);

INVX1 _3353_ (
    .A(_269_),
    .Y(_270_)
);

NAND3X1 _3354_ (
    .A(_257_),
    .B(_268_),
    .C(_270_),
    .Y(_271_)
);

INVX1 _3355_ (
    .A(_257_),
    .Y(_272_)
);

INVX1 _3356_ (
    .A(_268_),
    .Y(_273_)
);

OAI21X1 _3357_ (
    .A(_269_),
    .B(_273_),
    .C(_272_),
    .Y(_274_)
);

NAND2X1 _3358_ (
    .A(_274_),
    .B(_271_),
    .Y(_275_)
);

NOR2X1 _3359_ (
    .A(_275_),
    .B(_256_),
    .Y(_276_)
);

AND2X2 _3360_ (
    .A(_256_),
    .B(_275_),
    .Y(_277_)
);

NOR2X1 _3361_ (
    .A(_276_),
    .B(_277_),
    .Y(_3053_[20])
);

OAI21X1 _3362_ (
    .A(_275_),
    .B(_256_),
    .C(_271_),
    .Y(_278_)
);

OAI21X1 _3363_ (
    .A(_262_),
    .B(_263_),
    .C(_268_),
    .Y(_279_)
);

NOR2X1 _3364_ (
    .A(_230_),
    .B(_207_),
    .Y(_280_)
);

NAND3X1 _3365_ (
    .A(q1[12]),
    .B(q1[13]),
    .C(_280_),
    .Y(_281_)
);

INVX1 _3366_ (
    .A(q1[13]),
    .Y(_282_)
);

OAI21X1 _3367_ (
    .A(_260_),
    .B(_229_),
    .C(_282_),
    .Y(_283_)
);

NOR2X1 _3368_ (
    .A(q3[5]),
    .B(q2[13]),
    .Y(_284_)
);

INVX1 _3369_ (
    .A(q3[5]),
    .Y(_285_)
);

INVX1 _3370_ (
    .A(q2[13]),
    .Y(_286_)
);

NOR2X1 _3371_ (
    .A(_285_),
    .B(_286_),
    .Y(_287_)
);

NOR2X1 _3372_ (
    .A(_284_),
    .B(_287_),
    .Y(_288_)
);

NAND3X1 _3373_ (
    .A(_288_),
    .B(_283_),
    .C(_281_),
    .Y(_289_)
);

NOR3X1 _3374_ (
    .A(_260_),
    .B(_282_),
    .C(_229_),
    .Y(_290_)
);

AOI21X1 _3375_ (
    .A(_280_),
    .B(q1[12]),
    .C(q1[13]),
    .Y(_291_)
);

INVX1 _3376_ (
    .A(_288_),
    .Y(_292_)
);

OAI21X1 _3377_ (
    .A(_291_),
    .B(_290_),
    .C(_292_),
    .Y(_293_)
);

NAND3X1 _3378_ (
    .A(_279_),
    .B(_289_),
    .C(_293_),
    .Y(_294_)
);

AND2X2 _3379_ (
    .A(_268_),
    .B(_265_),
    .Y(_295_)
);

NAND3X1 _3380_ (
    .A(_292_),
    .B(_283_),
    .C(_281_),
    .Y(_296_)
);

OAI21X1 _3381_ (
    .A(_291_),
    .B(_290_),
    .C(_288_),
    .Y(_297_)
);

NAND3X1 _3382_ (
    .A(_296_),
    .B(_297_),
    .C(_295_),
    .Y(_298_)
);

NAND2X1 _3383_ (
    .A(_294_),
    .B(_298_),
    .Y(_299_)
);

OR2X2 _3384_ (
    .A(_278_),
    .B(_299_),
    .Y(_300_)
);

NAND2X1 _3385_ (
    .A(_299_),
    .B(_278_),
    .Y(_301_)
);

NAND2X1 _3386_ (
    .A(_301_),
    .B(_300_),
    .Y(_3053_[21])
);

NOR2X1 _3387_ (
    .A(_249_),
    .B(_246_),
    .Y(_302_)
);

NAND3X1 _3388_ (
    .A(_174_),
    .B(_199_),
    .C(_302_),
    .Y(_303_)
);

OAI21X1 _3389_ (
    .A(_219_),
    .B(_246_),
    .C(_240_),
    .Y(_304_)
);

AOI21X1 _3390_ (
    .A(_302_),
    .B(_202_),
    .C(_304_),
    .Y(_305_)
);

OAI21X1 _3391_ (
    .A(_303_),
    .B(_177_),
    .C(_305_),
    .Y(_306_)
);

OAI21X1 _3392_ (
    .A(_271_),
    .B(_299_),
    .C(_294_),
    .Y(_307_)
);

NOR2X1 _3393_ (
    .A(_275_),
    .B(_299_),
    .Y(_308_)
);

AOI21X1 _3394_ (
    .A(_306_),
    .B(_308_),
    .C(_307_),
    .Y(_309_)
);

OAI21X1 _3395_ (
    .A(_285_),
    .B(_286_),
    .C(_289_),
    .Y(_310_)
);

NOR3X1 _3396_ (
    .A(_230_),
    .B(_260_),
    .C(_207_),
    .Y(_311_)
);

NAND3X1 _3397_ (
    .A(q1[13]),
    .B(q1[14]),
    .C(_311_),
    .Y(_312_)
);

INVX1 _3398_ (
    .A(q1[14]),
    .Y(_313_)
);

OAI21X1 _3399_ (
    .A(_282_),
    .B(_259_),
    .C(_313_),
    .Y(_314_)
);

INVX1 _3400_ (
    .A(q3[6]),
    .Y(_315_)
);

INVX1 _3401_ (
    .A(q2[14]),
    .Y(_316_)
);

NAND2X1 _3402_ (
    .A(_315_),
    .B(_316_),
    .Y(_317_)
);

NAND2X1 _3403_ (
    .A(q3[6]),
    .B(q2[14]),
    .Y(_318_)
);

NAND2X1 _3404_ (
    .A(_318_),
    .B(_317_),
    .Y(_319_)
);

INVX1 _3405_ (
    .A(_319_),
    .Y(_320_)
);

NAND3X1 _3406_ (
    .A(_312_),
    .B(_320_),
    .C(_314_),
    .Y(_321_)
);

AOI21X1 _3407_ (
    .A(_314_),
    .B(_312_),
    .C(_320_),
    .Y(_322_)
);

INVX1 _3408_ (
    .A(_322_),
    .Y(_323_)
);

NAND3X1 _3409_ (
    .A(_310_),
    .B(_321_),
    .C(_323_),
    .Y(_324_)
);

INVX1 _3410_ (
    .A(_310_),
    .Y(_325_)
);

INVX1 _3411_ (
    .A(_321_),
    .Y(_326_)
);

OAI21X1 _3412_ (
    .A(_322_),
    .B(_326_),
    .C(_325_),
    .Y(_327_)
);

NAND2X1 _3413_ (
    .A(_324_),
    .B(_327_),
    .Y(_328_)
);

NOR2X1 _3414_ (
    .A(_328_),
    .B(_309_),
    .Y(_329_)
);

AND2X2 _3415_ (
    .A(_309_),
    .B(_328_),
    .Y(_330_)
);

NOR2X1 _3416_ (
    .A(_329_),
    .B(_330_),
    .Y(_3053_[22])
);

INVX1 _3417_ (
    .A(_324_),
    .Y(_331_)
);

NOR2X1 _3418_ (
    .A(_331_),
    .B(_329_),
    .Y(_332_)
);

OAI21X1 _3419_ (
    .A(_315_),
    .B(_316_),
    .C(_321_),
    .Y(_333_)
);

INVX1 _3420_ (
    .A(q3[7]),
    .Y(_334_)
);

INVX1 _3421_ (
    .A(q2[15]),
    .Y(_335_)
);

NAND2X1 _3422_ (
    .A(_334_),
    .B(_335_),
    .Y(_336_)
);

NAND2X1 _3423_ (
    .A(q3[7]),
    .B(q2[15]),
    .Y(_337_)
);

NAND2X1 _3424_ (
    .A(_337_),
    .B(_336_),
    .Y(_338_)
);

INVX1 _3425_ (
    .A(_338_),
    .Y(_339_)
);

INVX1 _3426_ (
    .A(q1[15]),
    .Y(_340_)
);

OAI21X1 _3427_ (
    .A(_313_),
    .B(_281_),
    .C(_340_),
    .Y(_341_)
);

NAND3X1 _3428_ (
    .A(q1[14]),
    .B(q1[15]),
    .C(_290_),
    .Y(_342_)
);

NAND3X1 _3429_ (
    .A(_339_),
    .B(_341_),
    .C(_342_),
    .Y(_343_)
);

OAI21X1 _3430_ (
    .A(_313_),
    .B(_281_),
    .C(q1[15]),
    .Y(_344_)
);

NAND3X1 _3431_ (
    .A(q1[14]),
    .B(_340_),
    .C(_290_),
    .Y(_345_)
);

NAND3X1 _3432_ (
    .A(_338_),
    .B(_344_),
    .C(_345_),
    .Y(_346_)
);

NAND3X1 _3433_ (
    .A(_343_),
    .B(_346_),
    .C(_333_),
    .Y(_347_)
);

AND2X2 _3434_ (
    .A(_321_),
    .B(_318_),
    .Y(_348_)
);

AOI21X1 _3435_ (
    .A(_345_),
    .B(_344_),
    .C(_338_),
    .Y(_349_)
);

AOI21X1 _3436_ (
    .A(_342_),
    .B(_341_),
    .C(_339_),
    .Y(_350_)
);

OAI21X1 _3437_ (
    .A(_349_),
    .B(_350_),
    .C(_348_),
    .Y(_351_)
);

AND2X2 _3438_ (
    .A(_351_),
    .B(_347_),
    .Y(_352_)
);

NAND2X1 _3439_ (
    .A(_352_),
    .B(_332_),
    .Y(_353_)
);

NAND2X1 _3440_ (
    .A(_347_),
    .B(_351_),
    .Y(_354_)
);

OAI21X1 _3441_ (
    .A(_331_),
    .B(_329_),
    .C(_354_),
    .Y(_355_)
);

NAND2X1 _3442_ (
    .A(_355_),
    .B(_353_),
    .Y(_3053_[23])
);

AND2X2 _3443_ (
    .A(_327_),
    .B(_324_),
    .Y(_356_)
);

NAND3X1 _3444_ (
    .A(_307_),
    .B(_356_),
    .C(_352_),
    .Y(_357_)
);

NAND2X1 _3445_ (
    .A(_331_),
    .B(_352_),
    .Y(_358_)
);

NAND3X1 _3446_ (
    .A(_347_),
    .B(_358_),
    .C(_357_),
    .Y(_359_)
);

NAND3X1 _3447_ (
    .A(_308_),
    .B(_356_),
    .C(_352_),
    .Y(_360_)
);

NOR2X1 _3448_ (
    .A(_256_),
    .B(_360_),
    .Y(_361_)
);

OAI21X1 _3449_ (
    .A(_334_),
    .B(_335_),
    .C(_343_),
    .Y(_362_)
);

NAND2X1 _3450_ (
    .A(q3[8]),
    .B(_362_),
    .Y(_363_)
);

OR2X2 _3451_ (
    .A(_362_),
    .B(q3[8]),
    .Y(_364_)
);

AND2X2 _3452_ (
    .A(_364_),
    .B(_363_),
    .Y(_365_)
);

OAI21X1 _3453_ (
    .A(_359_),
    .B(_361_),
    .C(_365_),
    .Y(_366_)
);

NOR2X1 _3454_ (
    .A(_328_),
    .B(_354_),
    .Y(_367_)
);

OAI21X1 _3455_ (
    .A(_324_),
    .B(_354_),
    .C(_347_),
    .Y(_368_)
);

AOI21X1 _3456_ (
    .A(_367_),
    .B(_307_),
    .C(_368_),
    .Y(_369_)
);

OAI21X1 _3457_ (
    .A(_256_),
    .B(_360_),
    .C(_369_),
    .Y(_370_)
);

OR2X2 _3458_ (
    .A(_370_),
    .B(_365_),
    .Y(_371_)
);

AND2X2 _3459_ (
    .A(_371_),
    .B(_366_),
    .Y(_3053_[24])
);

INVX1 _3460_ (
    .A(q3[9]),
    .Y(_372_)
);

NAND2X1 _3461_ (
    .A(_363_),
    .B(_366_),
    .Y(_373_)
);

NAND2X1 _3462_ (
    .A(_372_),
    .B(_373_),
    .Y(_374_)
);

NAND3X1 _3463_ (
    .A(q3[9]),
    .B(_363_),
    .C(_366_),
    .Y(_375_)
);

NAND2X1 _3464_ (
    .A(_375_),
    .B(_374_),
    .Y(_3053_[25])
);

INVX1 _3465_ (
    .A(q3[10]),
    .Y(_376_)
);

NOR2X1 _3466_ (
    .A(_372_),
    .B(_376_),
    .Y(_377_)
);

NAND2X1 _3467_ (
    .A(_377_),
    .B(_373_),
    .Y(_378_)
);

NOR2X1 _3468_ (
    .A(_372_),
    .B(_363_),
    .Y(_379_)
);

NAND3X1 _3469_ (
    .A(q3[9]),
    .B(_363_),
    .C(_364_),
    .Y(_380_)
);

INVX1 _3470_ (
    .A(_380_),
    .Y(_381_)
);

AOI21X1 _3471_ (
    .A(_370_),
    .B(_381_),
    .C(_379_),
    .Y(_382_)
);

NAND2X1 _3472_ (
    .A(_376_),
    .B(_382_),
    .Y(_383_)
);

AND2X2 _3473_ (
    .A(_378_),
    .B(_383_),
    .Y(_3053_[26])
);

OAI21X1 _3474_ (
    .A(_376_),
    .B(_382_),
    .C(q3[11]),
    .Y(_384_)
);

INVX1 _3475_ (
    .A(q3[11]),
    .Y(_385_)
);

NAND3X1 _3476_ (
    .A(_385_),
    .B(_377_),
    .C(_373_),
    .Y(_386_)
);

NAND2X1 _3477_ (
    .A(_386_),
    .B(_384_),
    .Y(_3053_[27])
);

INVX1 _3478_ (
    .A(q3[12]),
    .Y(_387_)
);

NOR2X1 _3479_ (
    .A(_376_),
    .B(_385_),
    .Y(_388_)
);

NAND2X1 _3480_ (
    .A(_388_),
    .B(_379_),
    .Y(_389_)
);

INVX1 _3481_ (
    .A(_389_),
    .Y(_390_)
);

NAND3X1 _3482_ (
    .A(_308_),
    .B(_367_),
    .C(_306_),
    .Y(_391_)
);

NAND3X1 _3483_ (
    .A(q3[9]),
    .B(_388_),
    .C(_365_),
    .Y(_392_)
);

AOI21X1 _3484_ (
    .A(_369_),
    .B(_391_),
    .C(_392_),
    .Y(_393_)
);

OAI21X1 _3485_ (
    .A(_390_),
    .B(_393_),
    .C(_387_),
    .Y(_394_)
);

INVX1 _3486_ (
    .A(_388_),
    .Y(_395_)
);

NOR2X1 _3487_ (
    .A(_395_),
    .B(_380_),
    .Y(_396_)
);

AOI21X1 _3488_ (
    .A(_370_),
    .B(_396_),
    .C(_390_),
    .Y(_397_)
);

NAND2X1 _3489_ (
    .A(q3[12]),
    .B(_397_),
    .Y(_398_)
);

NAND2X1 _3490_ (
    .A(_394_),
    .B(_398_),
    .Y(_3053_[28])
);

OAI21X1 _3491_ (
    .A(_387_),
    .B(_397_),
    .C(q3[13]),
    .Y(_399_)
);

INVX1 _3492_ (
    .A(q3[13]),
    .Y(_400_)
);

OAI21X1 _3493_ (
    .A(_359_),
    .B(_361_),
    .C(_396_),
    .Y(_401_)
);

NAND2X1 _3494_ (
    .A(_389_),
    .B(_401_),
    .Y(_402_)
);

NAND3X1 _3495_ (
    .A(q3[12]),
    .B(_400_),
    .C(_402_),
    .Y(_403_)
);

NAND2X1 _3496_ (
    .A(_403_),
    .B(_399_),
    .Y(_3053_[29])
);

INVX1 _3497_ (
    .A(q3[14]),
    .Y(_404_)
);

NOR2X1 _3498_ (
    .A(_387_),
    .B(_400_),
    .Y(_405_)
);

INVX1 _3499_ (
    .A(_405_),
    .Y(_406_)
);

AOI21X1 _3500_ (
    .A(_401_),
    .B(_389_),
    .C(_406_),
    .Y(_407_)
);

NAND2X1 _3501_ (
    .A(_404_),
    .B(_407_),
    .Y(_408_)
);

OAI21X1 _3502_ (
    .A(_406_),
    .B(_397_),
    .C(q3[14]),
    .Y(_409_)
);

NAND2X1 _3503_ (
    .A(_409_),
    .B(_408_),
    .Y(_3053_[30])
);

OAI21X1 _3504_ (
    .A(_390_),
    .B(_393_),
    .C(_405_),
    .Y(_410_)
);

OAI21X1 _3505_ (
    .A(_404_),
    .B(_410_),
    .C(q3[15]),
    .Y(_411_)
);

INVX1 _3506_ (
    .A(q3[15]),
    .Y(_412_)
);

NAND3X1 _3507_ (
    .A(q3[14]),
    .B(_412_),
    .C(_407_),
    .Y(_413_)
);

NAND2X1 _3508_ (
    .A(_413_),
    .B(_411_),
    .Y(_3053_[31])
);

AOI21X1 _3509_ (
    .A(_429_),
    .B(_428_),
    .C(_420_),
    .Y(_414_)
);

NOR2X1 _3510_ (
    .A(_414_),
    .B(_431_),
    .Y(_3053_[9])
);

OR2X2 _3511_ (
    .A(\z1.q1 [0]),
    .B(\z1.q0 [4]),
    .Y(_575_)
);

NAND2X1 _3512_ (
    .A(\z1.q1 [0]),
    .B(\z1.q0 [4]),
    .Y(_576_)
);

NAND2X1 _3513_ (
    .A(_576_),
    .B(_575_),
    .Y(_577_)
);

INVX1 _3514_ (
    .A(_577_),
    .Y(_578_)
);

AND2X2 _3515_ (
    .A(_578_),
    .B(\z1.q2 [0]),
    .Y(_579_)
);

NOR2X1 _3516_ (
    .A(\z1.q2 [0]),
    .B(_578_),
    .Y(_580_)
);

NOR2X1 _3517_ (
    .A(_580_),
    .B(_579_),
    .Y(q0[4])
);

INVX1 _3518_ (
    .A(\z1.z3.z1.z1.s ),
    .Y(_581_)
);

INVX1 _3519_ (
    .A(_576_),
    .Y(_582_)
);

NAND2X1 _3520_ (
    .A(\z1.z2.z1.z1.s ),
    .B(\z1.q0 [5]),
    .Y(_583_)
);

OR2X2 _3521_ (
    .A(\z1.z2.z1.z1.s ),
    .B(\z1.q0 [5]),
    .Y(_584_)
);

NAND3X1 _3522_ (
    .A(_583_),
    .B(_584_),
    .C(_582_),
    .Y(_585_)
);

AND2X2 _3523_ (
    .A(\z1.z2.z1.z1.s ),
    .B(\z1.q0 [5]),
    .Y(_586_)
);

NOR2X1 _3524_ (
    .A(\z1.z2.z1.z1.s ),
    .B(\z1.q0 [5]),
    .Y(_587_)
);

OAI21X1 _3525_ (
    .A(_587_),
    .B(_586_),
    .C(_576_),
    .Y(_588_)
);

NAND2X1 _3526_ (
    .A(_588_),
    .B(_585_),
    .Y(_589_)
);

OR2X2 _3527_ (
    .A(_589_),
    .B(_581_),
    .Y(_590_)
);

NAND2X1 _3528_ (
    .A(_581_),
    .B(_589_),
    .Y(_591_)
);

AND2X2 _3529_ (
    .A(_590_),
    .B(_591_),
    .Y(_592_)
);

NAND2X1 _3530_ (
    .A(_579_),
    .B(_592_),
    .Y(_593_)
);

INVX1 _3531_ (
    .A(_590_),
    .Y(_594_)
);

OAI21X1 _3532_ (
    .A(_576_),
    .B(_587_),
    .C(_583_),
    .Y(_595_)
);

INVX1 _3533_ (
    .A(\z1.q0 [6]),
    .Y(_596_)
);

NOR2X1 _3534_ (
    .A(\z1.q1 [2]),
    .B(_596_),
    .Y(_597_)
);

INVX1 _3535_ (
    .A(\z1.q1 [2]),
    .Y(_598_)
);

NOR2X1 _3536_ (
    .A(\z1.q0 [6]),
    .B(_598_),
    .Y(_599_)
);

OAI21X1 _3537_ (
    .A(_597_),
    .B(_599_),
    .C(_595_),
    .Y(_600_)
);

NAND2X1 _3538_ (
    .A(\z1.q0 [6]),
    .B(_598_),
    .Y(_601_)
);

NAND2X1 _3539_ (
    .A(\z1.q1 [2]),
    .B(_596_),
    .Y(_602_)
);

NAND2X1 _3540_ (
    .A(_601_),
    .B(_602_),
    .Y(_603_)
);

OR2X2 _3541_ (
    .A(_603_),
    .B(_595_),
    .Y(_604_)
);

NAND3X1 _3542_ (
    .A(\z1.q2 [2]),
    .B(_600_),
    .C(_604_),
    .Y(_605_)
);

INVX1 _3543_ (
    .A(\z1.q2 [2]),
    .Y(_606_)
);

NAND2X1 _3544_ (
    .A(_600_),
    .B(_604_),
    .Y(_607_)
);

NAND2X1 _3545_ (
    .A(_606_),
    .B(_607_),
    .Y(_608_)
);

AOI21X1 _3546_ (
    .A(_608_),
    .B(_605_),
    .C(_594_),
    .Y(_609_)
);

INVX1 _3547_ (
    .A(_609_),
    .Y(_610_)
);

NAND3X1 _3548_ (
    .A(_605_),
    .B(_608_),
    .C(_594_),
    .Y(_611_)
);

NAND3X1 _3549_ (
    .A(_593_),
    .B(_611_),
    .C(_610_),
    .Y(_612_)
);

INVX1 _3550_ (
    .A(_593_),
    .Y(_613_)
);

INVX1 _3551_ (
    .A(_611_),
    .Y(_614_)
);

OAI21X1 _3552_ (
    .A(_609_),
    .B(_614_),
    .C(_613_),
    .Y(_615_)
);

NAND2X1 _3553_ (
    .A(_612_),
    .B(_615_),
    .Y(q0[6])
);

OAI21X1 _3554_ (
    .A(_609_),
    .B(_593_),
    .C(_611_),
    .Y(_616_)
);

INVX1 _3555_ (
    .A(_605_),
    .Y(_617_)
);

INVX1 _3556_ (
    .A(\z1.q2 [3]),
    .Y(_618_)
);

INVX1 _3557_ (
    .A(\z1.q0 [7]),
    .Y(_619_)
);

NOR2X1 _3558_ (
    .A(\z1.q1 [3]),
    .B(_619_),
    .Y(_620_)
);

INVX1 _3559_ (
    .A(\z1.q1 [3]),
    .Y(_621_)
);

NOR2X1 _3560_ (
    .A(\z1.q0 [7]),
    .B(_621_),
    .Y(_622_)
);

NAND2X1 _3561_ (
    .A(\z1.q1 [2]),
    .B(\z1.q0 [6]),
    .Y(_623_)
);

INVX1 _3562_ (
    .A(_623_),
    .Y(_624_)
);

AOI21X1 _3563_ (
    .A(_603_),
    .B(_595_),
    .C(_624_),
    .Y(_625_)
);

OAI21X1 _3564_ (
    .A(_620_),
    .B(_622_),
    .C(_625_),
    .Y(_626_)
);

NAND2X1 _3565_ (
    .A(\z1.q1 [3]),
    .B(\z1.q0 [7]),
    .Y(_627_)
);

INVX1 _3566_ (
    .A(_627_),
    .Y(_628_)
);

NOR2X1 _3567_ (
    .A(\z1.q1 [3]),
    .B(\z1.q0 [7]),
    .Y(_629_)
);

INVX1 _3568_ (
    .A(_625_),
    .Y(_630_)
);

OAI21X1 _3569_ (
    .A(_628_),
    .B(_629_),
    .C(_630_),
    .Y(_631_)
);

AOI21X1 _3570_ (
    .A(_631_),
    .B(_626_),
    .C(_618_),
    .Y(_433_)
);

INVX1 _3571_ (
    .A(_433_),
    .Y(_434_)
);

NAND3X1 _3572_ (
    .A(_618_),
    .B(_626_),
    .C(_631_),
    .Y(_435_)
);

AOI21X1 _3573_ (
    .A(_434_),
    .B(_435_),
    .C(_617_),
    .Y(_436_)
);

NAND3X1 _3574_ (
    .A(_617_),
    .B(_435_),
    .C(_434_),
    .Y(_437_)
);

INVX1 _3575_ (
    .A(_437_),
    .Y(_438_)
);

OAI21X1 _3576_ (
    .A(_436_),
    .B(_438_),
    .C(_616_),
    .Y(_439_)
);

INVX1 _3577_ (
    .A(_616_),
    .Y(_440_)
);

NAND2X1 _3578_ (
    .A(_435_),
    .B(_434_),
    .Y(_441_)
);

OAI21X1 _3579_ (
    .A(_606_),
    .B(_607_),
    .C(_441_),
    .Y(_442_)
);

NAND3X1 _3580_ (
    .A(_437_),
    .B(_440_),
    .C(_442_),
    .Y(_443_)
);

NAND2X1 _3581_ (
    .A(_443_),
    .B(_439_),
    .Y(q0[7])
);

AOI21X1 _3582_ (
    .A(_442_),
    .B(_616_),
    .C(_438_),
    .Y(_444_)
);

AOI21X1 _3583_ (
    .A(_582_),
    .B(_584_),
    .C(_586_),
    .Y(_445_)
);

OAI22X1 _3584_ (
    .A(_597_),
    .B(_599_),
    .C(_620_),
    .D(_622_),
    .Y(_446_)
);

OAI21X1 _3585_ (
    .A(_623_),
    .B(_629_),
    .C(_627_),
    .Y(_447_)
);

INVX1 _3586_ (
    .A(_447_),
    .Y(_448_)
);

OAI21X1 _3587_ (
    .A(_445_),
    .B(_446_),
    .C(_448_),
    .Y(_449_)
);

NAND2X1 _3588_ (
    .A(\z1.q1 [4]),
    .B(_449_),
    .Y(_450_)
);

INVX1 _3589_ (
    .A(\z1.q1 [4]),
    .Y(_451_)
);

NAND2X1 _3590_ (
    .A(\z1.q0 [7]),
    .B(_621_),
    .Y(_452_)
);

NAND2X1 _3591_ (
    .A(\z1.q1 [3]),
    .B(_619_),
    .Y(_453_)
);

NAND2X1 _3592_ (
    .A(_452_),
    .B(_453_),
    .Y(_454_)
);

NAND3X1 _3593_ (
    .A(_595_),
    .B(_603_),
    .C(_454_),
    .Y(_455_)
);

NAND3X1 _3594_ (
    .A(_451_),
    .B(_448_),
    .C(_455_),
    .Y(_456_)
);

NAND2X1 _3595_ (
    .A(\z1.q3 [0]),
    .B(\z1.q2 [4]),
    .Y(_457_)
);

INVX1 _3596_ (
    .A(\z1.q3 [0]),
    .Y(_458_)
);

INVX1 _3597_ (
    .A(\z1.q2 [4]),
    .Y(_459_)
);

NAND2X1 _3598_ (
    .A(_458_),
    .B(_459_),
    .Y(_460_)
);

NAND2X1 _3599_ (
    .A(_457_),
    .B(_460_),
    .Y(_461_)
);

INVX1 _3600_ (
    .A(_461_),
    .Y(_462_)
);

NAND3X1 _3601_ (
    .A(_456_),
    .B(_462_),
    .C(_450_),
    .Y(_463_)
);

AOI21X1 _3602_ (
    .A(_455_),
    .B(_448_),
    .C(_451_),
    .Y(_464_)
);

INVX1 _3603_ (
    .A(_456_),
    .Y(_465_)
);

OAI21X1 _3604_ (
    .A(_464_),
    .B(_465_),
    .C(_461_),
    .Y(_466_)
);

NAND3X1 _3605_ (
    .A(_463_),
    .B(_466_),
    .C(_433_),
    .Y(_467_)
);

NAND2X1 _3606_ (
    .A(_463_),
    .B(_466_),
    .Y(_468_)
);

NAND2X1 _3607_ (
    .A(_468_),
    .B(_434_),
    .Y(_469_)
);

AND2X2 _3608_ (
    .A(_469_),
    .B(_467_),
    .Y(_470_)
);

NAND2X1 _3609_ (
    .A(_470_),
    .B(_444_),
    .Y(_471_)
);

OAI21X1 _3610_ (
    .A(_436_),
    .B(_440_),
    .C(_437_),
    .Y(_472_)
);

NAND2X1 _3611_ (
    .A(_467_),
    .B(_469_),
    .Y(_473_)
);

NAND2X1 _3612_ (
    .A(_473_),
    .B(_472_),
    .Y(_474_)
);

NAND2X1 _3613_ (
    .A(_471_),
    .B(_474_),
    .Y(q0[8])
);

OAI21X1 _3614_ (
    .A(_473_),
    .B(_444_),
    .C(_467_),
    .Y(_475_)
);

OAI21X1 _3615_ (
    .A(_458_),
    .B(_459_),
    .C(_463_),
    .Y(_476_)
);

NAND3X1 _3616_ (
    .A(\z1.q1 [4]),
    .B(\z1.q1 [5]),
    .C(_449_),
    .Y(_477_)
);

INVX1 _3617_ (
    .A(\z1.q1 [5]),
    .Y(_478_)
);

AOI22X1 _3618_ (
    .A(_601_),
    .B(_602_),
    .C(_452_),
    .D(_453_),
    .Y(_479_)
);

AOI21X1 _3619_ (
    .A(_479_),
    .B(_595_),
    .C(_447_),
    .Y(_480_)
);

OAI21X1 _3620_ (
    .A(_451_),
    .B(_480_),
    .C(_478_),
    .Y(_481_)
);

INVX1 _3621_ (
    .A(\z1.z4.z1.z1.s ),
    .Y(_482_)
);

INVX1 _3622_ (
    .A(\z1.q2 [5]),
    .Y(_483_)
);

NAND2X1 _3623_ (
    .A(_482_),
    .B(_483_),
    .Y(_484_)
);

NAND2X1 _3624_ (
    .A(\z1.z4.z1.z1.s ),
    .B(\z1.q2 [5]),
    .Y(_485_)
);

AND2X2 _3625_ (
    .A(_484_),
    .B(_485_),
    .Y(_486_)
);

NAND3X1 _3626_ (
    .A(_486_),
    .B(_481_),
    .C(_477_),
    .Y(_487_)
);

AOI21X1 _3627_ (
    .A(_477_),
    .B(_481_),
    .C(_486_),
    .Y(_488_)
);

INVX1 _3628_ (
    .A(_488_),
    .Y(_489_)
);

NAND3X1 _3629_ (
    .A(_487_),
    .B(_476_),
    .C(_489_),
    .Y(_490_)
);

AND2X2 _3630_ (
    .A(_463_),
    .B(_457_),
    .Y(_491_)
);

INVX1 _3631_ (
    .A(_487_),
    .Y(_492_)
);

OAI21X1 _3632_ (
    .A(_492_),
    .B(_488_),
    .C(_491_),
    .Y(_493_)
);

NAND2X1 _3633_ (
    .A(_490_),
    .B(_493_),
    .Y(_494_)
);

OR2X2 _3634_ (
    .A(_475_),
    .B(_494_),
    .Y(_495_)
);

NAND2X1 _3635_ (
    .A(_494_),
    .B(_475_),
    .Y(_496_)
);

NAND2X1 _3636_ (
    .A(_496_),
    .B(_495_),
    .Y(q0[9])
);

NAND3X1 _3637_ (
    .A(_490_),
    .B(_493_),
    .C(_470_),
    .Y(_497_)
);

OAI21X1 _3638_ (
    .A(_434_),
    .B(_468_),
    .C(_490_),
    .Y(_498_)
);

NAND2X1 _3639_ (
    .A(_493_),
    .B(_498_),
    .Y(_499_)
);

OAI21X1 _3640_ (
    .A(_444_),
    .B(_497_),
    .C(_499_),
    .Y(_500_)
);

OAI21X1 _3641_ (
    .A(_482_),
    .B(_483_),
    .C(_487_),
    .Y(_501_)
);

NAND3X1 _3642_ (
    .A(\z1.q1 [5]),
    .B(\z1.q1 [6]),
    .C(_464_),
    .Y(_502_)
);

INVX1 _3643_ (
    .A(\z1.q1 [6]),
    .Y(_503_)
);

NAND2X1 _3644_ (
    .A(_503_),
    .B(_477_),
    .Y(_504_)
);

INVX1 _3645_ (
    .A(\z1.q3 [2]),
    .Y(_505_)
);

INVX1 _3646_ (
    .A(\z1.q2 [6]),
    .Y(_506_)
);

NAND2X1 _3647_ (
    .A(_505_),
    .B(_506_),
    .Y(_507_)
);

NAND2X1 _3648_ (
    .A(\z1.q3 [2]),
    .B(\z1.q2 [6]),
    .Y(_508_)
);

NAND2X1 _3649_ (
    .A(_508_),
    .B(_507_),
    .Y(_509_)
);

INVX1 _3650_ (
    .A(_509_),
    .Y(_510_)
);

NAND3X1 _3651_ (
    .A(_502_),
    .B(_510_),
    .C(_504_),
    .Y(_511_)
);

AOI21X1 _3652_ (
    .A(_504_),
    .B(_502_),
    .C(_510_),
    .Y(_512_)
);

INVX1 _3653_ (
    .A(_512_),
    .Y(_513_)
);

NAND3X1 _3654_ (
    .A(_501_),
    .B(_511_),
    .C(_513_),
    .Y(_514_)
);

INVX1 _3655_ (
    .A(_501_),
    .Y(_515_)
);

INVX1 _3656_ (
    .A(_511_),
    .Y(_516_)
);

OAI21X1 _3657_ (
    .A(_512_),
    .B(_516_),
    .C(_515_),
    .Y(_517_)
);

NAND2X1 _3658_ (
    .A(_517_),
    .B(_514_),
    .Y(_518_)
);

NAND2X1 _3659_ (
    .A(_518_),
    .B(_500_),
    .Y(_519_)
);

NOR2X1 _3660_ (
    .A(_473_),
    .B(_494_),
    .Y(_520_)
);

AOI22X1 _3661_ (
    .A(_493_),
    .B(_498_),
    .C(_520_),
    .D(_472_),
    .Y(_521_)
);

AND2X2 _3662_ (
    .A(_514_),
    .B(_517_),
    .Y(_522_)
);

NAND2X1 _3663_ (
    .A(_522_),
    .B(_521_),
    .Y(_523_)
);

NAND2X1 _3664_ (
    .A(_519_),
    .B(_523_),
    .Y(q0[10])
);

OAI21X1 _3665_ (
    .A(_518_),
    .B(_521_),
    .C(_514_),
    .Y(_524_)
);

OAI21X1 _3666_ (
    .A(_505_),
    .B(_506_),
    .C(_511_),
    .Y(_525_)
);

NOR2X1 _3667_ (
    .A(\z1.q3 [3]),
    .B(\z1.q2 [7]),
    .Y(_526_)
);

INVX1 _3668_ (
    .A(\z1.q3 [3]),
    .Y(_527_)
);

INVX1 _3669_ (
    .A(\z1.q2 [7]),
    .Y(_528_)
);

NOR2X1 _3670_ (
    .A(_527_),
    .B(_528_),
    .Y(_529_)
);

NOR2X1 _3671_ (
    .A(_526_),
    .B(_529_),
    .Y(_530_)
);

INVX1 _3672_ (
    .A(\z1.q1 [7]),
    .Y(_531_)
);

OAI21X1 _3673_ (
    .A(_503_),
    .B(_477_),
    .C(_531_),
    .Y(_532_)
);

AND2X2 _3674_ (
    .A(_464_),
    .B(\z1.q1 [5]),
    .Y(_533_)
);

NAND3X1 _3675_ (
    .A(\z1.q1 [6]),
    .B(\z1.q1 [7]),
    .C(_533_),
    .Y(_534_)
);

NAND3X1 _3676_ (
    .A(_530_),
    .B(_532_),
    .C(_534_),
    .Y(_535_)
);

INVX1 _3677_ (
    .A(_530_),
    .Y(_536_)
);

OAI21X1 _3678_ (
    .A(_503_),
    .B(_477_),
    .C(\z1.q1 [7]),
    .Y(_537_)
);

NAND3X1 _3679_ (
    .A(\z1.q1 [6]),
    .B(_531_),
    .C(_533_),
    .Y(_538_)
);

NAND3X1 _3680_ (
    .A(_536_),
    .B(_537_),
    .C(_538_),
    .Y(_539_)
);

NAND3X1 _3681_ (
    .A(_535_),
    .B(_539_),
    .C(_525_),
    .Y(_540_)
);

AND2X2 _3682_ (
    .A(_511_),
    .B(_508_),
    .Y(_541_)
);

NAND2X1 _3683_ (
    .A(_535_),
    .B(_539_),
    .Y(_542_)
);

NAND2X1 _3684_ (
    .A(_541_),
    .B(_542_),
    .Y(_543_)
);

NAND2X1 _3685_ (
    .A(_540_),
    .B(_543_),
    .Y(_544_)
);

OR2X2 _3686_ (
    .A(_524_),
    .B(_544_),
    .Y(_545_)
);

NAND2X1 _3687_ (
    .A(_544_),
    .B(_524_),
    .Y(_546_)
);

NAND2X1 _3688_ (
    .A(_546_),
    .B(_545_),
    .Y(q0[11])
);

OAI21X1 _3689_ (
    .A(_541_),
    .B(_542_),
    .C(_514_),
    .Y(_547_)
);

NAND2X1 _3690_ (
    .A(_543_),
    .B(_547_),
    .Y(_548_)
);

NAND3X1 _3691_ (
    .A(_540_),
    .B(_543_),
    .C(_522_),
    .Y(_549_)
);

OAI21X1 _3692_ (
    .A(_549_),
    .B(_521_),
    .C(_548_),
    .Y(_550_)
);

OAI21X1 _3693_ (
    .A(_527_),
    .B(_528_),
    .C(_535_),
    .Y(_551_)
);

NAND2X1 _3694_ (
    .A(\z1.q3 [4]),
    .B(_551_),
    .Y(_552_)
);

OR2X2 _3695_ (
    .A(_551_),
    .B(\z1.q3 [4]),
    .Y(_553_)
);

NAND3X1 _3696_ (
    .A(_552_),
    .B(_553_),
    .C(_550_),
    .Y(_554_)
);

NOR2X1 _3697_ (
    .A(_518_),
    .B(_544_),
    .Y(_555_)
);

AOI22X1 _3698_ (
    .A(_543_),
    .B(_547_),
    .C(_555_),
    .D(_500_),
    .Y(_556_)
);

NAND2X1 _3699_ (
    .A(_552_),
    .B(_553_),
    .Y(_557_)
);

NAND2X1 _3700_ (
    .A(_557_),
    .B(_556_),
    .Y(_558_)
);

AND2X2 _3701_ (
    .A(_554_),
    .B(_558_),
    .Y(q0[12])
);

INVX1 _3702_ (
    .A(\z1.q3 [5]),
    .Y(_559_)
);

OAI21X1 _3703_ (
    .A(_557_),
    .B(_556_),
    .C(_552_),
    .Y(_560_)
);

NAND2X1 _3704_ (
    .A(_559_),
    .B(_560_),
    .Y(_561_)
);

NAND3X1 _3705_ (
    .A(\z1.q3 [5]),
    .B(_552_),
    .C(_554_),
    .Y(_562_)
);

NAND2X1 _3706_ (
    .A(_562_),
    .B(_561_),
    .Y(q0[13])
);

INVX1 _3707_ (
    .A(\z1.q3 [6]),
    .Y(_563_)
);

NAND3X1 _3708_ (
    .A(\z1.q3 [5]),
    .B(_552_),
    .C(_553_),
    .Y(_564_)
);

OAI22X1 _3709_ (
    .A(_559_),
    .B(_552_),
    .C(_564_),
    .D(_556_),
    .Y(_565_)
);

NAND2X1 _3710_ (
    .A(_563_),
    .B(_565_),
    .Y(_566_)
);

INVX1 _3711_ (
    .A(_552_),
    .Y(_567_)
);

INVX1 _3712_ (
    .A(_564_),
    .Y(_568_)
);

AOI22X1 _3713_ (
    .A(\z1.q3 [5]),
    .B(_567_),
    .C(_550_),
    .D(_568_),
    .Y(_569_)
);

NAND2X1 _3714_ (
    .A(\z1.q3 [6]),
    .B(_569_),
    .Y(_570_)
);

NAND2X1 _3715_ (
    .A(_570_),
    .B(_566_),
    .Y(q0[14])
);

OAI21X1 _3716_ (
    .A(_563_),
    .B(_569_),
    .C(\z1.q3 [7]),
    .Y(_571_)
);

INVX1 _3717_ (
    .A(\z1.q3 [7]),
    .Y(_572_)
);

NAND3X1 _3718_ (
    .A(\z1.q3 [6]),
    .B(_572_),
    .C(_565_),
    .Y(_573_)
);

NAND2X1 _3719_ (
    .A(_573_),
    .B(_571_),
    .Y(q0[15])
);

NOR2X1 _3720_ (
    .A(_579_),
    .B(_592_),
    .Y(_574_)
);

NOR2X1 _3721_ (
    .A(_574_),
    .B(_613_),
    .Y(q0[5])
);

NOR2X1 _3722_ (
    .A(\z1.z1.q1 [0]),
    .B(\z1.z1.z1.z2.s ),
    .Y(_639_)
);

AND2X2 _3723_ (
    .A(\z1.z1.q1 [0]),
    .B(\z1.z1.z1.z2.s ),
    .Y(_640_)
);

NOR2X1 _3724_ (
    .A(_639_),
    .B(_640_),
    .Y(_641_)
);

NAND2X1 _3725_ (
    .A(\z1.z1.q2 [0]),
    .B(_641_),
    .Y(_642_)
);

INVX1 _3726_ (
    .A(_642_),
    .Y(_643_)
);

NOR2X1 _3727_ (
    .A(\z1.z1.q2 [0]),
    .B(_641_),
    .Y(_644_)
);

NOR2X1 _3728_ (
    .A(_644_),
    .B(_643_),
    .Y(q0[2])
);

NAND2X1 _3729_ (
    .A(\z1.z1.q1 [0]),
    .B(\z1.z1.z1.z2.s ),
    .Y(_645_)
);

NOR2X1 _3730_ (
    .A(\z1.z1.z2.z1.s ),
    .B(\z1.z1.z1.z2.c ),
    .Y(_646_)
);

NAND2X1 _3731_ (
    .A(\z1.z1.z2.z1.s ),
    .B(\z1.z1.z1.z2.c ),
    .Y(_647_)
);

INVX1 _3732_ (
    .A(_647_),
    .Y(_648_)
);

OAI21X1 _3733_ (
    .A(_646_),
    .B(_648_),
    .C(_645_),
    .Y(_649_)
);

INVX1 _3734_ (
    .A(\z1.z1.z2.z1.s ),
    .Y(_650_)
);

INVX1 _3735_ (
    .A(\z1.z1.z1.z2.c ),
    .Y(_651_)
);

NAND2X1 _3736_ (
    .A(_650_),
    .B(_651_),
    .Y(_652_)
);

NAND3X1 _3737_ (
    .A(_640_),
    .B(_647_),
    .C(_652_),
    .Y(_653_)
);

NAND3X1 _3738_ (
    .A(\z1.z1.z3.z1.s ),
    .B(_653_),
    .C(_649_),
    .Y(_654_)
);

INVX1 _3739_ (
    .A(\z1.z1.z3.z1.s ),
    .Y(_655_)
);

NAND2X1 _3740_ (
    .A(_653_),
    .B(_649_),
    .Y(_656_)
);

NAND2X1 _3741_ (
    .A(_655_),
    .B(_656_),
    .Y(_657_)
);

NAND3X1 _3742_ (
    .A(_643_),
    .B(_654_),
    .C(_657_),
    .Y(_658_)
);

INVX1 _3743_ (
    .A(_658_),
    .Y(_659_)
);

INVX1 _3744_ (
    .A(_654_),
    .Y(_660_)
);

OAI21X1 _3745_ (
    .A(_645_),
    .B(_646_),
    .C(_647_),
    .Y(_661_)
);

NAND2X1 _3746_ (
    .A(\z1.z1.z2.z2.s ),
    .B(_661_),
    .Y(_662_)
);

INVX1 _3747_ (
    .A(\z1.z1.z2.z2.s ),
    .Y(_663_)
);

NAND3X1 _3748_ (
    .A(_663_),
    .B(_647_),
    .C(_653_),
    .Y(_664_)
);

NAND2X1 _3749_ (
    .A(\z1.z1.q3 [0]),
    .B(\z1.z1.z3.z2.s ),
    .Y(_665_)
);

INVX1 _3750_ (
    .A(\z1.z1.q3 [0]),
    .Y(_666_)
);

INVX1 _3751_ (
    .A(\z1.z1.z3.z2.s ),
    .Y(_667_)
);

NAND2X1 _3752_ (
    .A(_666_),
    .B(_667_),
    .Y(_668_)
);

NAND2X1 _3753_ (
    .A(_665_),
    .B(_668_),
    .Y(_669_)
);

INVX1 _3754_ (
    .A(_669_),
    .Y(_670_)
);

NAND3X1 _3755_ (
    .A(_662_),
    .B(_670_),
    .C(_664_),
    .Y(_671_)
);

AND2X2 _3756_ (
    .A(_661_),
    .B(\z1.z1.z2.z2.s ),
    .Y(_672_)
);

NOR2X1 _3757_ (
    .A(\z1.z1.z2.z2.s ),
    .B(_661_),
    .Y(_673_)
);

OAI21X1 _3758_ (
    .A(_673_),
    .B(_672_),
    .C(_669_),
    .Y(_674_)
);

NAND3X1 _3759_ (
    .A(_660_),
    .B(_671_),
    .C(_674_),
    .Y(_675_)
);

INVX1 _3760_ (
    .A(_671_),
    .Y(_676_)
);

AOI21X1 _3761_ (
    .A(_664_),
    .B(_662_),
    .C(_670_),
    .Y(_677_)
);

OAI21X1 _3762_ (
    .A(_677_),
    .B(_676_),
    .C(_654_),
    .Y(_678_)
);

NAND3X1 _3763_ (
    .A(_659_),
    .B(_675_),
    .C(_678_),
    .Y(_679_)
);

INVX1 _3764_ (
    .A(_675_),
    .Y(_680_)
);

INVX1 _3765_ (
    .A(_656_),
    .Y(_681_)
);

AOI22X1 _3766_ (
    .A(\z1.z1.z3.z1.s ),
    .B(_681_),
    .C(_674_),
    .D(_671_),
    .Y(_682_)
);

OAI21X1 _3767_ (
    .A(_682_),
    .B(_680_),
    .C(_658_),
    .Y(_683_)
);

AND2X2 _3768_ (
    .A(_683_),
    .B(_679_),
    .Y(\z1.q0 [4])
);

OAI21X1 _3769_ (
    .A(_658_),
    .B(_682_),
    .C(_675_),
    .Y(_684_)
);

OAI21X1 _3770_ (
    .A(_666_),
    .B(_667_),
    .C(_671_),
    .Y(_685_)
);

NAND2X1 _3771_ (
    .A(\z1.z1.z4.z1.s ),
    .B(\z1.z1.z3.z2.c ),
    .Y(_686_)
);

OR2X2 _3772_ (
    .A(\z1.z1.z4.z1.s ),
    .B(\z1.z1.z3.z2.c ),
    .Y(_687_)
);

NAND2X1 _3773_ (
    .A(_686_),
    .B(_687_),
    .Y(_688_)
);

INVX1 _3774_ (
    .A(_688_),
    .Y(_689_)
);

NAND2X1 _3775_ (
    .A(\z1.z1.z2.z2.c ),
    .B(_672_),
    .Y(_690_)
);

INVX1 _3776_ (
    .A(\z1.z1.z2.z2.c ),
    .Y(_691_)
);

NAND2X1 _3777_ (
    .A(_691_),
    .B(_662_),
    .Y(_692_)
);

NAND3X1 _3778_ (
    .A(_689_),
    .B(_692_),
    .C(_690_),
    .Y(_693_)
);

NAND2X1 _3779_ (
    .A(\z1.z1.z2.z2.c ),
    .B(_662_),
    .Y(_694_)
);

NAND2X1 _3780_ (
    .A(_691_),
    .B(_672_),
    .Y(_695_)
);

NAND3X1 _3781_ (
    .A(_688_),
    .B(_694_),
    .C(_695_),
    .Y(_696_)
);

NAND3X1 _3782_ (
    .A(_685_),
    .B(_693_),
    .C(_696_),
    .Y(_697_)
);

INVX1 _3783_ (
    .A(_685_),
    .Y(_698_)
);

AOI21X1 _3784_ (
    .A(_695_),
    .B(_694_),
    .C(_688_),
    .Y(_699_)
);

AOI21X1 _3785_ (
    .A(_690_),
    .B(_692_),
    .C(_689_),
    .Y(_700_)
);

OAI21X1 _3786_ (
    .A(_699_),
    .B(_700_),
    .C(_698_),
    .Y(_701_)
);

NAND2X1 _3787_ (
    .A(_697_),
    .B(_701_),
    .Y(_702_)
);

NAND2X1 _3788_ (
    .A(_684_),
    .B(_702_),
    .Y(_703_)
);

OR2X2 _3789_ (
    .A(_702_),
    .B(_684_),
    .Y(_704_)
);

NAND2X1 _3790_ (
    .A(_703_),
    .B(_704_),
    .Y(\z1.q0 [5])
);

INVX1 _3791_ (
    .A(\z1.z1.z4.z2.s ),
    .Y(_705_)
);

INVX1 _3792_ (
    .A(_686_),
    .Y(_706_)
);

OAI21X1 _3793_ (
    .A(_706_),
    .B(_699_),
    .C(_705_),
    .Y(_707_)
);

NAND3X1 _3794_ (
    .A(\z1.z1.z4.z2.s ),
    .B(_686_),
    .C(_693_),
    .Y(_708_)
);

NAND2X1 _3795_ (
    .A(_701_),
    .B(_684_),
    .Y(_709_)
);

AOI22X1 _3796_ (
    .A(_707_),
    .B(_708_),
    .C(_709_),
    .D(_697_),
    .Y(_710_)
);

NAND2X1 _3797_ (
    .A(_708_),
    .B(_707_),
    .Y(_711_)
);

NAND3X1 _3798_ (
    .A(_675_),
    .B(_697_),
    .C(_679_),
    .Y(_712_)
);

AOI21X1 _3799_ (
    .A(_712_),
    .B(_701_),
    .C(_711_),
    .Y(_713_)
);

NOR2X1 _3800_ (
    .A(_710_),
    .B(_713_),
    .Y(\z1.q0 [6])
);

OAI21X1 _3801_ (
    .A(_706_),
    .B(_699_),
    .C(\z1.z1.z4.z2.s ),
    .Y(_632_)
);

NAND3X1 _3802_ (
    .A(_701_),
    .B(_711_),
    .C(_712_),
    .Y(_633_)
);

NAND3X1 _3803_ (
    .A(\z1.z1.z4.z2.c ),
    .B(_632_),
    .C(_633_),
    .Y(_634_)
);

INVX1 _3804_ (
    .A(\z1.z1.z4.z2.c ),
    .Y(_635_)
);

INVX1 _3805_ (
    .A(_632_),
    .Y(_636_)
);

OAI21X1 _3806_ (
    .A(_636_),
    .B(_710_),
    .C(_635_),
    .Y(_637_)
);

NAND2X1 _3807_ (
    .A(_634_),
    .B(_637_),
    .Y(\z1.q0 [7])
);

AOI21X1 _3808_ (
    .A(_657_),
    .B(_654_),
    .C(_643_),
    .Y(_638_)
);

NOR2X1 _3809_ (
    .A(_638_),
    .B(_659_),
    .Y(q0[3])
);

AND2X2 _3810_ (
    .A(b[0]),
    .B(a[0]),
    .Y(q0[0])
);

AND2X2 _3811_ (
    .A(b[0]),
    .B(a[1]),
    .Y(\z1.z1.z1.z1.a )
);

AND2X2 _3812_ (
    .A(a[0]),
    .B(b[1]),
    .Y(\z1.z1.z1.z1.b )
);

AND2X2 _3813_ (
    .A(a[1]),
    .B(b[1]),
    .Y(\z1.z1.z1.z2.a )
);

INVX1 _3814_ (
    .A(\z1.z1.z1.z1.b ),
    .Y(_714_)
);

NAND2X1 _3815_ (
    .A(\z1.z1.z1.z1.a ),
    .B(_714_),
    .Y(_715_)
);

INVX1 _3816_ (
    .A(\z1.z1.z1.z1.a ),
    .Y(_716_)
);

NAND2X1 _3817_ (
    .A(\z1.z1.z1.z1.b ),
    .B(_716_),
    .Y(_717_)
);

NAND2X1 _3818_ (
    .A(_715_),
    .B(_717_),
    .Y(\z1.z1.z1.z1.s )
);

NOR2X1 _3819_ (
    .A(_714_),
    .B(_716_),
    .Y(\z1.z1.z1.z1.c )
);

INVX1 _3820_ (
    .A(\z1.z1.z1.z1.c ),
    .Y(_718_)
);

NAND2X1 _3821_ (
    .A(\z1.z1.z1.z2.a ),
    .B(_718_),
    .Y(_719_)
);

INVX1 _3822_ (
    .A(\z1.z1.z1.z2.a ),
    .Y(_720_)
);

NAND2X1 _3823_ (
    .A(\z1.z1.z1.z1.c ),
    .B(_720_),
    .Y(_721_)
);

NAND2X1 _3824_ (
    .A(_719_),
    .B(_721_),
    .Y(\z1.z1.z1.z2.s )
);

NOR2X1 _3825_ (
    .A(_718_),
    .B(_720_),
    .Y(\z1.z1.z1.z2.c )
);

AND2X2 _3826_ (
    .A(b[0]),
    .B(a[2]),
    .Y(\z1.z1.q1 [0])
);

AND2X2 _3827_ (
    .A(b[0]),
    .B(a[3]),
    .Y(\z1.z1.z2.z1.a )
);

AND2X2 _3828_ (
    .A(a[2]),
    .B(b[1]),
    .Y(\z1.z1.z2.z1.b )
);

AND2X2 _3829_ (
    .A(a[3]),
    .B(b[1]),
    .Y(\z1.z1.z2.z2.a )
);

INVX1 _3830_ (
    .A(\z1.z1.z2.z1.b ),
    .Y(_722_)
);

NAND2X1 _3831_ (
    .A(\z1.z1.z2.z1.a ),
    .B(_722_),
    .Y(_723_)
);

INVX1 _3832_ (
    .A(\z1.z1.z2.z1.a ),
    .Y(_724_)
);

NAND2X1 _3833_ (
    .A(\z1.z1.z2.z1.b ),
    .B(_724_),
    .Y(_725_)
);

NAND2X1 _3834_ (
    .A(_723_),
    .B(_725_),
    .Y(\z1.z1.z2.z1.s )
);

NOR2X1 _3835_ (
    .A(_722_),
    .B(_724_),
    .Y(\z1.z1.z2.z1.c )
);

INVX1 _3836_ (
    .A(\z1.z1.z2.z1.c ),
    .Y(_726_)
);

NAND2X1 _3837_ (
    .A(\z1.z1.z2.z2.a ),
    .B(_726_),
    .Y(_727_)
);

INVX1 _3838_ (
    .A(\z1.z1.z2.z2.a ),
    .Y(_728_)
);

NAND2X1 _3839_ (
    .A(\z1.z1.z2.z1.c ),
    .B(_728_),
    .Y(_729_)
);

NAND2X1 _3840_ (
    .A(_727_),
    .B(_729_),
    .Y(\z1.z1.z2.z2.s )
);

NOR2X1 _3841_ (
    .A(_726_),
    .B(_728_),
    .Y(\z1.z1.z2.z2.c )
);

AND2X2 _3842_ (
    .A(b[2]),
    .B(a[0]),
    .Y(\z1.z1.q2 [0])
);

AND2X2 _3843_ (
    .A(b[2]),
    .B(a[1]),
    .Y(\z1.z1.z3.z1.a )
);

AND2X2 _3844_ (
    .A(a[0]),
    .B(b[3]),
    .Y(\z1.z1.z3.z1.b )
);

AND2X2 _3845_ (
    .A(a[1]),
    .B(b[3]),
    .Y(\z1.z1.z3.z2.a )
);

INVX1 _3846_ (
    .A(\z1.z1.z3.z1.b ),
    .Y(_730_)
);

NAND2X1 _3847_ (
    .A(\z1.z1.z3.z1.a ),
    .B(_730_),
    .Y(_731_)
);

INVX1 _3848_ (
    .A(\z1.z1.z3.z1.a ),
    .Y(_732_)
);

NAND2X1 _3849_ (
    .A(\z1.z1.z3.z1.b ),
    .B(_732_),
    .Y(_733_)
);

NAND2X1 _3850_ (
    .A(_731_),
    .B(_733_),
    .Y(\z1.z1.z3.z1.s )
);

NOR2X1 _3851_ (
    .A(_730_),
    .B(_732_),
    .Y(\z1.z1.z3.z1.c )
);

INVX1 _3852_ (
    .A(\z1.z1.z3.z1.c ),
    .Y(_734_)
);

NAND2X1 _3853_ (
    .A(\z1.z1.z3.z2.a ),
    .B(_734_),
    .Y(_735_)
);

INVX1 _3854_ (
    .A(\z1.z1.z3.z2.a ),
    .Y(_736_)
);

NAND2X1 _3855_ (
    .A(\z1.z1.z3.z1.c ),
    .B(_736_),
    .Y(_737_)
);

NAND2X1 _3856_ (
    .A(_735_),
    .B(_737_),
    .Y(\z1.z1.z3.z2.s )
);

NOR2X1 _3857_ (
    .A(_734_),
    .B(_736_),
    .Y(\z1.z1.z3.z2.c )
);

AND2X2 _3858_ (
    .A(b[2]),
    .B(a[2]),
    .Y(\z1.z1.q3 [0])
);

AND2X2 _3859_ (
    .A(b[2]),
    .B(a[3]),
    .Y(\z1.z1.z4.z1.a )
);

AND2X2 _3860_ (
    .A(a[2]),
    .B(b[3]),
    .Y(\z1.z1.z4.z1.b )
);

AND2X2 _3861_ (
    .A(a[3]),
    .B(b[3]),
    .Y(\z1.z1.z4.z2.a )
);

INVX1 _3862_ (
    .A(\z1.z1.z4.z1.b ),
    .Y(_738_)
);

NAND2X1 _3863_ (
    .A(\z1.z1.z4.z1.a ),
    .B(_738_),
    .Y(_739_)
);

INVX1 _3864_ (
    .A(\z1.z1.z4.z1.a ),
    .Y(_740_)
);

NAND2X1 _3865_ (
    .A(\z1.z1.z4.z1.b ),
    .B(_740_),
    .Y(_741_)
);

NAND2X1 _3866_ (
    .A(_739_),
    .B(_741_),
    .Y(\z1.z1.z4.z1.s )
);

NOR2X1 _3867_ (
    .A(_738_),
    .B(_740_),
    .Y(\z1.z1.z4.z1.c )
);

INVX1 _3868_ (
    .A(\z1.z1.z4.z1.c ),
    .Y(_742_)
);

NAND2X1 _3869_ (
    .A(\z1.z1.z4.z2.a ),
    .B(_742_),
    .Y(_743_)
);

INVX1 _3870_ (
    .A(\z1.z1.z4.z2.a ),
    .Y(_744_)
);

NAND2X1 _3871_ (
    .A(\z1.z1.z4.z1.c ),
    .B(_744_),
    .Y(_745_)
);

NAND2X1 _3872_ (
    .A(_743_),
    .B(_745_),
    .Y(\z1.z1.z4.z2.s )
);

NOR2X1 _3873_ (
    .A(_742_),
    .B(_744_),
    .Y(\z1.z1.z4.z2.c )
);

NOR2X1 _3874_ (
    .A(\z1.z2.q1 [0]),
    .B(\z1.z2.z1.z2.s ),
    .Y(_753_)
);

AND2X2 _3875_ (
    .A(\z1.z2.q1 [0]),
    .B(\z1.z2.z1.z2.s ),
    .Y(_754_)
);

NOR2X1 _3876_ (
    .A(_753_),
    .B(_754_),
    .Y(_755_)
);

NAND2X1 _3877_ (
    .A(\z1.z2.q2 [0]),
    .B(_755_),
    .Y(_756_)
);

INVX1 _3878_ (
    .A(_756_),
    .Y(_757_)
);

NOR2X1 _3879_ (
    .A(\z1.z2.q2 [0]),
    .B(_755_),
    .Y(_758_)
);

NOR2X1 _3880_ (
    .A(_758_),
    .B(_757_),
    .Y(\z1.q1 [2])
);

NAND2X1 _3881_ (
    .A(\z1.z2.q1 [0]),
    .B(\z1.z2.z1.z2.s ),
    .Y(_759_)
);

NOR2X1 _3882_ (
    .A(\z1.z2.z2.z1.s ),
    .B(\z1.z2.z1.z2.c ),
    .Y(_760_)
);

NAND2X1 _3883_ (
    .A(\z1.z2.z2.z1.s ),
    .B(\z1.z2.z1.z2.c ),
    .Y(_761_)
);

INVX1 _3884_ (
    .A(_761_),
    .Y(_762_)
);

OAI21X1 _3885_ (
    .A(_760_),
    .B(_762_),
    .C(_759_),
    .Y(_763_)
);

INVX1 _3886_ (
    .A(\z1.z2.z2.z1.s ),
    .Y(_764_)
);

INVX1 _3887_ (
    .A(\z1.z2.z1.z2.c ),
    .Y(_765_)
);

NAND2X1 _3888_ (
    .A(_764_),
    .B(_765_),
    .Y(_766_)
);

NAND3X1 _3889_ (
    .A(_754_),
    .B(_761_),
    .C(_766_),
    .Y(_767_)
);

NAND3X1 _3890_ (
    .A(\z1.z2.z3.z1.s ),
    .B(_767_),
    .C(_763_),
    .Y(_768_)
);

INVX1 _3891_ (
    .A(\z1.z2.z3.z1.s ),
    .Y(_769_)
);

NAND2X1 _3892_ (
    .A(_767_),
    .B(_763_),
    .Y(_770_)
);

NAND2X1 _3893_ (
    .A(_769_),
    .B(_770_),
    .Y(_771_)
);

NAND3X1 _3894_ (
    .A(_757_),
    .B(_768_),
    .C(_771_),
    .Y(_772_)
);

INVX1 _3895_ (
    .A(_772_),
    .Y(_773_)
);

INVX1 _3896_ (
    .A(_768_),
    .Y(_774_)
);

OAI21X1 _3897_ (
    .A(_759_),
    .B(_760_),
    .C(_761_),
    .Y(_775_)
);

NAND2X1 _3898_ (
    .A(\z1.z2.z2.z2.s ),
    .B(_775_),
    .Y(_776_)
);

INVX1 _3899_ (
    .A(\z1.z2.z2.z2.s ),
    .Y(_777_)
);

NAND3X1 _3900_ (
    .A(_777_),
    .B(_761_),
    .C(_767_),
    .Y(_778_)
);

NAND2X1 _3901_ (
    .A(\z1.z2.q3 [0]),
    .B(\z1.z2.z3.z2.s ),
    .Y(_779_)
);

INVX1 _3902_ (
    .A(\z1.z2.q3 [0]),
    .Y(_780_)
);

INVX1 _3903_ (
    .A(\z1.z2.z3.z2.s ),
    .Y(_781_)
);

NAND2X1 _3904_ (
    .A(_780_),
    .B(_781_),
    .Y(_782_)
);

NAND2X1 _3905_ (
    .A(_779_),
    .B(_782_),
    .Y(_783_)
);

INVX1 _3906_ (
    .A(_783_),
    .Y(_784_)
);

NAND3X1 _3907_ (
    .A(_776_),
    .B(_784_),
    .C(_778_),
    .Y(_785_)
);

AND2X2 _3908_ (
    .A(_775_),
    .B(\z1.z2.z2.z2.s ),
    .Y(_786_)
);

NOR2X1 _3909_ (
    .A(\z1.z2.z2.z2.s ),
    .B(_775_),
    .Y(_787_)
);

OAI21X1 _3910_ (
    .A(_787_),
    .B(_786_),
    .C(_783_),
    .Y(_788_)
);

NAND3X1 _3911_ (
    .A(_774_),
    .B(_785_),
    .C(_788_),
    .Y(_789_)
);

INVX1 _3912_ (
    .A(_785_),
    .Y(_790_)
);

AOI21X1 _3913_ (
    .A(_778_),
    .B(_776_),
    .C(_784_),
    .Y(_791_)
);

OAI21X1 _3914_ (
    .A(_791_),
    .B(_790_),
    .C(_768_),
    .Y(_792_)
);

NAND3X1 _3915_ (
    .A(_773_),
    .B(_789_),
    .C(_792_),
    .Y(_793_)
);

INVX1 _3916_ (
    .A(_789_),
    .Y(_794_)
);

INVX1 _3917_ (
    .A(_770_),
    .Y(_795_)
);

AOI22X1 _3918_ (
    .A(\z1.z2.z3.z1.s ),
    .B(_795_),
    .C(_788_),
    .D(_785_),
    .Y(_796_)
);

OAI21X1 _3919_ (
    .A(_796_),
    .B(_794_),
    .C(_772_),
    .Y(_797_)
);

AND2X2 _3920_ (
    .A(_797_),
    .B(_793_),
    .Y(\z1.q1 [4])
);

OAI21X1 _3921_ (
    .A(_772_),
    .B(_796_),
    .C(_789_),
    .Y(_798_)
);

OAI21X1 _3922_ (
    .A(_780_),
    .B(_781_),
    .C(_785_),
    .Y(_799_)
);

NAND2X1 _3923_ (
    .A(\z1.z2.z4.z1.s ),
    .B(\z1.z2.z3.z2.c ),
    .Y(_800_)
);

OR2X2 _3924_ (
    .A(\z1.z2.z4.z1.s ),
    .B(\z1.z2.z3.z2.c ),
    .Y(_801_)
);

NAND2X1 _3925_ (
    .A(_800_),
    .B(_801_),
    .Y(_802_)
);

INVX1 _3926_ (
    .A(_802_),
    .Y(_803_)
);

NAND2X1 _3927_ (
    .A(\z1.z2.z2.z2.c ),
    .B(_786_),
    .Y(_804_)
);

INVX1 _3928_ (
    .A(\z1.z2.z2.z2.c ),
    .Y(_805_)
);

NAND2X1 _3929_ (
    .A(_805_),
    .B(_776_),
    .Y(_806_)
);

NAND3X1 _3930_ (
    .A(_803_),
    .B(_806_),
    .C(_804_),
    .Y(_807_)
);

NAND2X1 _3931_ (
    .A(\z1.z2.z2.z2.c ),
    .B(_776_),
    .Y(_808_)
);

NAND2X1 _3932_ (
    .A(_805_),
    .B(_786_),
    .Y(_809_)
);

NAND3X1 _3933_ (
    .A(_802_),
    .B(_808_),
    .C(_809_),
    .Y(_810_)
);

NAND3X1 _3934_ (
    .A(_799_),
    .B(_807_),
    .C(_810_),
    .Y(_811_)
);

INVX1 _3935_ (
    .A(_799_),
    .Y(_812_)
);

AOI21X1 _3936_ (
    .A(_809_),
    .B(_808_),
    .C(_802_),
    .Y(_813_)
);

AOI21X1 _3937_ (
    .A(_804_),
    .B(_806_),
    .C(_803_),
    .Y(_814_)
);

OAI21X1 _3938_ (
    .A(_813_),
    .B(_814_),
    .C(_812_),
    .Y(_815_)
);

NAND2X1 _3939_ (
    .A(_811_),
    .B(_815_),
    .Y(_816_)
);

NAND2X1 _3940_ (
    .A(_798_),
    .B(_816_),
    .Y(_817_)
);

OR2X2 _3941_ (
    .A(_816_),
    .B(_798_),
    .Y(_818_)
);

NAND2X1 _3942_ (
    .A(_817_),
    .B(_818_),
    .Y(\z1.q1 [5])
);

INVX1 _3943_ (
    .A(\z1.z2.z4.z2.s ),
    .Y(_819_)
);

INVX1 _3944_ (
    .A(_800_),
    .Y(_820_)
);

OAI21X1 _3945_ (
    .A(_820_),
    .B(_813_),
    .C(_819_),
    .Y(_821_)
);

NAND3X1 _3946_ (
    .A(\z1.z2.z4.z2.s ),
    .B(_800_),
    .C(_807_),
    .Y(_822_)
);

NAND2X1 _3947_ (
    .A(_815_),
    .B(_798_),
    .Y(_823_)
);

AOI22X1 _3948_ (
    .A(_821_),
    .B(_822_),
    .C(_823_),
    .D(_811_),
    .Y(_824_)
);

NAND2X1 _3949_ (
    .A(_822_),
    .B(_821_),
    .Y(_825_)
);

NAND3X1 _3950_ (
    .A(_789_),
    .B(_811_),
    .C(_793_),
    .Y(_826_)
);

AOI21X1 _3951_ (
    .A(_826_),
    .B(_815_),
    .C(_825_),
    .Y(_827_)
);

NOR2X1 _3952_ (
    .A(_824_),
    .B(_827_),
    .Y(\z1.q1 [6])
);

OAI21X1 _3953_ (
    .A(_820_),
    .B(_813_),
    .C(\z1.z2.z4.z2.s ),
    .Y(_746_)
);

NAND3X1 _3954_ (
    .A(_815_),
    .B(_825_),
    .C(_826_),
    .Y(_747_)
);

NAND3X1 _3955_ (
    .A(\z1.z2.z4.z2.c ),
    .B(_746_),
    .C(_747_),
    .Y(_748_)
);

INVX1 _3956_ (
    .A(\z1.z2.z4.z2.c ),
    .Y(_749_)
);

INVX1 _3957_ (
    .A(_746_),
    .Y(_750_)
);

OAI21X1 _3958_ (
    .A(_750_),
    .B(_824_),
    .C(_749_),
    .Y(_751_)
);

NAND2X1 _3959_ (
    .A(_748_),
    .B(_751_),
    .Y(\z1.q1 [7])
);

AOI21X1 _3960_ (
    .A(_771_),
    .B(_768_),
    .C(_757_),
    .Y(_752_)
);

NOR2X1 _3961_ (
    .A(_752_),
    .B(_773_),
    .Y(\z1.q1 [3])
);

AND2X2 _3962_ (
    .A(b[0]),
    .B(a[4]),
    .Y(\z1.q1 [0])
);

AND2X2 _3963_ (
    .A(b[0]),
    .B(a[5]),
    .Y(\z1.z2.z1.z1.a )
);

AND2X2 _3964_ (
    .A(a[4]),
    .B(b[1]),
    .Y(\z1.z2.z1.z1.b )
);

AND2X2 _3965_ (
    .A(a[5]),
    .B(b[1]),
    .Y(\z1.z2.z1.z2.a )
);

INVX1 _3966_ (
    .A(\z1.z2.z1.z1.b ),
    .Y(_828_)
);

NAND2X1 _3967_ (
    .A(\z1.z2.z1.z1.a ),
    .B(_828_),
    .Y(_829_)
);

INVX1 _3968_ (
    .A(\z1.z2.z1.z1.a ),
    .Y(_830_)
);

NAND2X1 _3969_ (
    .A(\z1.z2.z1.z1.b ),
    .B(_830_),
    .Y(_831_)
);

NAND2X1 _3970_ (
    .A(_829_),
    .B(_831_),
    .Y(\z1.z2.z1.z1.s )
);

NOR2X1 _3971_ (
    .A(_828_),
    .B(_830_),
    .Y(\z1.z2.z1.z1.c )
);

INVX1 _3972_ (
    .A(\z1.z2.z1.z1.c ),
    .Y(_832_)
);

NAND2X1 _3973_ (
    .A(\z1.z2.z1.z2.a ),
    .B(_832_),
    .Y(_833_)
);

INVX1 _3974_ (
    .A(\z1.z2.z1.z2.a ),
    .Y(_834_)
);

NAND2X1 _3975_ (
    .A(\z1.z2.z1.z1.c ),
    .B(_834_),
    .Y(_835_)
);

NAND2X1 _3976_ (
    .A(_833_),
    .B(_835_),
    .Y(\z1.z2.z1.z2.s )
);

NOR2X1 _3977_ (
    .A(_832_),
    .B(_834_),
    .Y(\z1.z2.z1.z2.c )
);

AND2X2 _3978_ (
    .A(b[0]),
    .B(a[6]),
    .Y(\z1.z2.q1 [0])
);

AND2X2 _3979_ (
    .A(b[0]),
    .B(a[7]),
    .Y(\z1.z2.z2.z1.a )
);

AND2X2 _3980_ (
    .A(a[6]),
    .B(b[1]),
    .Y(\z1.z2.z2.z1.b )
);

AND2X2 _3981_ (
    .A(a[7]),
    .B(b[1]),
    .Y(\z1.z2.z2.z2.a )
);

INVX1 _3982_ (
    .A(\z1.z2.z2.z1.b ),
    .Y(_836_)
);

NAND2X1 _3983_ (
    .A(\z1.z2.z2.z1.a ),
    .B(_836_),
    .Y(_837_)
);

INVX1 _3984_ (
    .A(\z1.z2.z2.z1.a ),
    .Y(_838_)
);

NAND2X1 _3985_ (
    .A(\z1.z2.z2.z1.b ),
    .B(_838_),
    .Y(_839_)
);

NAND2X1 _3986_ (
    .A(_837_),
    .B(_839_),
    .Y(\z1.z2.z2.z1.s )
);

NOR2X1 _3987_ (
    .A(_836_),
    .B(_838_),
    .Y(\z1.z2.z2.z1.c )
);

INVX1 _3988_ (
    .A(\z1.z2.z2.z1.c ),
    .Y(_840_)
);

NAND2X1 _3989_ (
    .A(\z1.z2.z2.z2.a ),
    .B(_840_),
    .Y(_841_)
);

INVX1 _3990_ (
    .A(\z1.z2.z2.z2.a ),
    .Y(_842_)
);

NAND2X1 _3991_ (
    .A(\z1.z2.z2.z1.c ),
    .B(_842_),
    .Y(_843_)
);

NAND2X1 _3992_ (
    .A(_841_),
    .B(_843_),
    .Y(\z1.z2.z2.z2.s )
);

NOR2X1 _3993_ (
    .A(_840_),
    .B(_842_),
    .Y(\z1.z2.z2.z2.c )
);

AND2X2 _3994_ (
    .A(b[2]),
    .B(a[4]),
    .Y(\z1.z2.q2 [0])
);

AND2X2 _3995_ (
    .A(b[2]),
    .B(a[5]),
    .Y(\z1.z2.z3.z1.a )
);

AND2X2 _3996_ (
    .A(a[4]),
    .B(b[3]),
    .Y(\z1.z2.z3.z1.b )
);

AND2X2 _3997_ (
    .A(a[5]),
    .B(b[3]),
    .Y(\z1.z2.z3.z2.a )
);

INVX1 _3998_ (
    .A(\z1.z2.z3.z1.b ),
    .Y(_844_)
);

NAND2X1 _3999_ (
    .A(\z1.z2.z3.z1.a ),
    .B(_844_),
    .Y(_845_)
);

INVX1 _4000_ (
    .A(\z1.z2.z3.z1.a ),
    .Y(_846_)
);

NAND2X1 _4001_ (
    .A(\z1.z2.z3.z1.b ),
    .B(_846_),
    .Y(_847_)
);

NAND2X1 _4002_ (
    .A(_845_),
    .B(_847_),
    .Y(\z1.z2.z3.z1.s )
);

NOR2X1 _4003_ (
    .A(_844_),
    .B(_846_),
    .Y(\z1.z2.z3.z1.c )
);

INVX1 _4004_ (
    .A(\z1.z2.z3.z1.c ),
    .Y(_848_)
);

NAND2X1 _4005_ (
    .A(\z1.z2.z3.z2.a ),
    .B(_848_),
    .Y(_849_)
);

INVX1 _4006_ (
    .A(\z1.z2.z3.z2.a ),
    .Y(_850_)
);

NAND2X1 _4007_ (
    .A(\z1.z2.z3.z1.c ),
    .B(_850_),
    .Y(_851_)
);

NAND2X1 _4008_ (
    .A(_849_),
    .B(_851_),
    .Y(\z1.z2.z3.z2.s )
);

NOR2X1 _4009_ (
    .A(_848_),
    .B(_850_),
    .Y(\z1.z2.z3.z2.c )
);

AND2X2 _4010_ (
    .A(b[2]),
    .B(a[6]),
    .Y(\z1.z2.q3 [0])
);

AND2X2 _4011_ (
    .A(b[2]),
    .B(a[7]),
    .Y(\z1.z2.z4.z1.a )
);

AND2X2 _4012_ (
    .A(a[6]),
    .B(b[3]),
    .Y(\z1.z2.z4.z1.b )
);

AND2X2 _4013_ (
    .A(a[7]),
    .B(b[3]),
    .Y(\z1.z2.z4.z2.a )
);

INVX1 _4014_ (
    .A(\z1.z2.z4.z1.b ),
    .Y(_852_)
);

NAND2X1 _4015_ (
    .A(\z1.z2.z4.z1.a ),
    .B(_852_),
    .Y(_853_)
);

INVX1 _4016_ (
    .A(\z1.z2.z4.z1.a ),
    .Y(_854_)
);

NAND2X1 _4017_ (
    .A(\z1.z2.z4.z1.b ),
    .B(_854_),
    .Y(_855_)
);

NAND2X1 _4018_ (
    .A(_853_),
    .B(_855_),
    .Y(\z1.z2.z4.z1.s )
);

NOR2X1 _4019_ (
    .A(_852_),
    .B(_854_),
    .Y(\z1.z2.z4.z1.c )
);

INVX1 _4020_ (
    .A(\z1.z2.z4.z1.c ),
    .Y(_856_)
);

NAND2X1 _4021_ (
    .A(\z1.z2.z4.z2.a ),
    .B(_856_),
    .Y(_857_)
);

INVX1 _4022_ (
    .A(\z1.z2.z4.z2.a ),
    .Y(_858_)
);

NAND2X1 _4023_ (
    .A(\z1.z2.z4.z1.c ),
    .B(_858_),
    .Y(_859_)
);

NAND2X1 _4024_ (
    .A(_857_),
    .B(_859_),
    .Y(\z1.z2.z4.z2.s )
);

NOR2X1 _4025_ (
    .A(_856_),
    .B(_858_),
    .Y(\z1.z2.z4.z2.c )
);

NOR2X1 _4026_ (
    .A(\z1.z3.q1 [0]),
    .B(\z1.z3.z1.z2.s ),
    .Y(_867_)
);

AND2X2 _4027_ (
    .A(\z1.z3.q1 [0]),
    .B(\z1.z3.z1.z2.s ),
    .Y(_868_)
);

NOR2X1 _4028_ (
    .A(_867_),
    .B(_868_),
    .Y(_869_)
);

NAND2X1 _4029_ (
    .A(\z1.z3.q2 [0]),
    .B(_869_),
    .Y(_870_)
);

INVX1 _4030_ (
    .A(_870_),
    .Y(_871_)
);

NOR2X1 _4031_ (
    .A(\z1.z3.q2 [0]),
    .B(_869_),
    .Y(_872_)
);

NOR2X1 _4032_ (
    .A(_872_),
    .B(_871_),
    .Y(\z1.q2 [2])
);

NAND2X1 _4033_ (
    .A(\z1.z3.q1 [0]),
    .B(\z1.z3.z1.z2.s ),
    .Y(_873_)
);

NOR2X1 _4034_ (
    .A(\z1.z3.z2.z1.s ),
    .B(\z1.z3.z1.z2.c ),
    .Y(_874_)
);

NAND2X1 _4035_ (
    .A(\z1.z3.z2.z1.s ),
    .B(\z1.z3.z1.z2.c ),
    .Y(_875_)
);

INVX1 _4036_ (
    .A(_875_),
    .Y(_876_)
);

OAI21X1 _4037_ (
    .A(_874_),
    .B(_876_),
    .C(_873_),
    .Y(_877_)
);

INVX1 _4038_ (
    .A(\z1.z3.z2.z1.s ),
    .Y(_878_)
);

INVX1 _4039_ (
    .A(\z1.z3.z1.z2.c ),
    .Y(_879_)
);

NAND2X1 _4040_ (
    .A(_878_),
    .B(_879_),
    .Y(_880_)
);

NAND3X1 _4041_ (
    .A(_868_),
    .B(_875_),
    .C(_880_),
    .Y(_881_)
);

NAND3X1 _4042_ (
    .A(\z1.z3.z3.z1.s ),
    .B(_881_),
    .C(_877_),
    .Y(_882_)
);

INVX1 _4043_ (
    .A(\z1.z3.z3.z1.s ),
    .Y(_883_)
);

NAND2X1 _4044_ (
    .A(_881_),
    .B(_877_),
    .Y(_884_)
);

NAND2X1 _4045_ (
    .A(_883_),
    .B(_884_),
    .Y(_885_)
);

NAND3X1 _4046_ (
    .A(_871_),
    .B(_882_),
    .C(_885_),
    .Y(_886_)
);

INVX1 _4047_ (
    .A(_886_),
    .Y(_887_)
);

INVX1 _4048_ (
    .A(_882_),
    .Y(_888_)
);

OAI21X1 _4049_ (
    .A(_873_),
    .B(_874_),
    .C(_875_),
    .Y(_889_)
);

NAND2X1 _4050_ (
    .A(\z1.z3.z2.z2.s ),
    .B(_889_),
    .Y(_890_)
);

INVX1 _4051_ (
    .A(\z1.z3.z2.z2.s ),
    .Y(_891_)
);

NAND3X1 _4052_ (
    .A(_891_),
    .B(_875_),
    .C(_881_),
    .Y(_892_)
);

NAND2X1 _4053_ (
    .A(\z1.z3.q3 [0]),
    .B(\z1.z3.z3.z2.s ),
    .Y(_893_)
);

INVX1 _4054_ (
    .A(\z1.z3.q3 [0]),
    .Y(_894_)
);

INVX1 _4055_ (
    .A(\z1.z3.z3.z2.s ),
    .Y(_895_)
);

NAND2X1 _4056_ (
    .A(_894_),
    .B(_895_),
    .Y(_896_)
);

NAND2X1 _4057_ (
    .A(_893_),
    .B(_896_),
    .Y(_897_)
);

INVX1 _4058_ (
    .A(_897_),
    .Y(_898_)
);

NAND3X1 _4059_ (
    .A(_890_),
    .B(_898_),
    .C(_892_),
    .Y(_899_)
);

AND2X2 _4060_ (
    .A(_889_),
    .B(\z1.z3.z2.z2.s ),
    .Y(_900_)
);

NOR2X1 _4061_ (
    .A(\z1.z3.z2.z2.s ),
    .B(_889_),
    .Y(_901_)
);

OAI21X1 _4062_ (
    .A(_901_),
    .B(_900_),
    .C(_897_),
    .Y(_902_)
);

NAND3X1 _4063_ (
    .A(_888_),
    .B(_899_),
    .C(_902_),
    .Y(_903_)
);

INVX1 _4064_ (
    .A(_899_),
    .Y(_904_)
);

AOI21X1 _4065_ (
    .A(_892_),
    .B(_890_),
    .C(_898_),
    .Y(_905_)
);

OAI21X1 _4066_ (
    .A(_905_),
    .B(_904_),
    .C(_882_),
    .Y(_906_)
);

NAND3X1 _4067_ (
    .A(_887_),
    .B(_903_),
    .C(_906_),
    .Y(_907_)
);

INVX1 _4068_ (
    .A(_903_),
    .Y(_908_)
);

INVX1 _4069_ (
    .A(_884_),
    .Y(_909_)
);

AOI22X1 _4070_ (
    .A(\z1.z3.z3.z1.s ),
    .B(_909_),
    .C(_902_),
    .D(_899_),
    .Y(_910_)
);

OAI21X1 _4071_ (
    .A(_910_),
    .B(_908_),
    .C(_886_),
    .Y(_911_)
);

AND2X2 _4072_ (
    .A(_911_),
    .B(_907_),
    .Y(\z1.q2 [4])
);

OAI21X1 _4073_ (
    .A(_886_),
    .B(_910_),
    .C(_903_),
    .Y(_912_)
);

OAI21X1 _4074_ (
    .A(_894_),
    .B(_895_),
    .C(_899_),
    .Y(_913_)
);

NAND2X1 _4075_ (
    .A(\z1.z3.z4.z1.s ),
    .B(\z1.z3.z3.z2.c ),
    .Y(_914_)
);

OR2X2 _4076_ (
    .A(\z1.z3.z4.z1.s ),
    .B(\z1.z3.z3.z2.c ),
    .Y(_915_)
);

NAND2X1 _4077_ (
    .A(_914_),
    .B(_915_),
    .Y(_916_)
);

INVX1 _4078_ (
    .A(_916_),
    .Y(_917_)
);

NAND2X1 _4079_ (
    .A(\z1.z3.z2.z2.c ),
    .B(_900_),
    .Y(_918_)
);

INVX1 _4080_ (
    .A(\z1.z3.z2.z2.c ),
    .Y(_919_)
);

NAND2X1 _4081_ (
    .A(_919_),
    .B(_890_),
    .Y(_920_)
);

NAND3X1 _4082_ (
    .A(_917_),
    .B(_920_),
    .C(_918_),
    .Y(_921_)
);

NAND2X1 _4083_ (
    .A(\z1.z3.z2.z2.c ),
    .B(_890_),
    .Y(_922_)
);

NAND2X1 _4084_ (
    .A(_919_),
    .B(_900_),
    .Y(_923_)
);

NAND3X1 _4085_ (
    .A(_916_),
    .B(_922_),
    .C(_923_),
    .Y(_924_)
);

NAND3X1 _4086_ (
    .A(_913_),
    .B(_921_),
    .C(_924_),
    .Y(_925_)
);

INVX1 _4087_ (
    .A(_913_),
    .Y(_926_)
);

AOI21X1 _4088_ (
    .A(_923_),
    .B(_922_),
    .C(_916_),
    .Y(_927_)
);

AOI21X1 _4089_ (
    .A(_918_),
    .B(_920_),
    .C(_917_),
    .Y(_928_)
);

OAI21X1 _4090_ (
    .A(_927_),
    .B(_928_),
    .C(_926_),
    .Y(_929_)
);

NAND2X1 _4091_ (
    .A(_925_),
    .B(_929_),
    .Y(_930_)
);

NAND2X1 _4092_ (
    .A(_912_),
    .B(_930_),
    .Y(_931_)
);

OR2X2 _4093_ (
    .A(_930_),
    .B(_912_),
    .Y(_932_)
);

NAND2X1 _4094_ (
    .A(_931_),
    .B(_932_),
    .Y(\z1.q2 [5])
);

INVX1 _4095_ (
    .A(\z1.z3.z4.z2.s ),
    .Y(_933_)
);

INVX1 _4096_ (
    .A(_914_),
    .Y(_934_)
);

OAI21X1 _4097_ (
    .A(_934_),
    .B(_927_),
    .C(_933_),
    .Y(_935_)
);

NAND3X1 _4098_ (
    .A(\z1.z3.z4.z2.s ),
    .B(_914_),
    .C(_921_),
    .Y(_936_)
);

NAND2X1 _4099_ (
    .A(_929_),
    .B(_912_),
    .Y(_937_)
);

AOI22X1 _4100_ (
    .A(_935_),
    .B(_936_),
    .C(_937_),
    .D(_925_),
    .Y(_938_)
);

NAND2X1 _4101_ (
    .A(_936_),
    .B(_935_),
    .Y(_939_)
);

NAND3X1 _4102_ (
    .A(_903_),
    .B(_925_),
    .C(_907_),
    .Y(_940_)
);

AOI21X1 _4103_ (
    .A(_940_),
    .B(_929_),
    .C(_939_),
    .Y(_941_)
);

NOR2X1 _4104_ (
    .A(_938_),
    .B(_941_),
    .Y(\z1.q2 [6])
);

OAI21X1 _4105_ (
    .A(_934_),
    .B(_927_),
    .C(\z1.z3.z4.z2.s ),
    .Y(_860_)
);

NAND3X1 _4106_ (
    .A(_929_),
    .B(_939_),
    .C(_940_),
    .Y(_861_)
);

NAND3X1 _4107_ (
    .A(\z1.z3.z4.z2.c ),
    .B(_860_),
    .C(_861_),
    .Y(_862_)
);

INVX1 _4108_ (
    .A(\z1.z3.z4.z2.c ),
    .Y(_863_)
);

INVX1 _4109_ (
    .A(_860_),
    .Y(_864_)
);

OAI21X1 _4110_ (
    .A(_864_),
    .B(_938_),
    .C(_863_),
    .Y(_865_)
);

NAND2X1 _4111_ (
    .A(_862_),
    .B(_865_),
    .Y(\z1.q2 [7])
);

AOI21X1 _4112_ (
    .A(_885_),
    .B(_882_),
    .C(_871_),
    .Y(_866_)
);

NOR2X1 _4113_ (
    .A(_866_),
    .B(_887_),
    .Y(\z1.q2 [3])
);

AND2X2 _4114_ (
    .A(b[4]),
    .B(a[0]),
    .Y(\z1.q2 [0])
);

AND2X2 _4115_ (
    .A(b[4]),
    .B(a[1]),
    .Y(\z1.z3.z1.z1.a )
);

AND2X2 _4116_ (
    .A(a[0]),
    .B(b[5]),
    .Y(\z1.z3.z1.z1.b )
);

AND2X2 _4117_ (
    .A(a[1]),
    .B(b[5]),
    .Y(\z1.z3.z1.z2.a )
);

INVX1 _4118_ (
    .A(\z1.z3.z1.z1.b ),
    .Y(_942_)
);

NAND2X1 _4119_ (
    .A(\z1.z3.z1.z1.a ),
    .B(_942_),
    .Y(_943_)
);

INVX1 _4120_ (
    .A(\z1.z3.z1.z1.a ),
    .Y(_944_)
);

NAND2X1 _4121_ (
    .A(\z1.z3.z1.z1.b ),
    .B(_944_),
    .Y(_945_)
);

NAND2X1 _4122_ (
    .A(_943_),
    .B(_945_),
    .Y(\z1.z3.z1.z1.s )
);

NOR2X1 _4123_ (
    .A(_942_),
    .B(_944_),
    .Y(\z1.z3.z1.z1.c )
);

INVX1 _4124_ (
    .A(\z1.z3.z1.z1.c ),
    .Y(_946_)
);

NAND2X1 _4125_ (
    .A(\z1.z3.z1.z2.a ),
    .B(_946_),
    .Y(_947_)
);

INVX1 _4126_ (
    .A(\z1.z3.z1.z2.a ),
    .Y(_948_)
);

NAND2X1 _4127_ (
    .A(\z1.z3.z1.z1.c ),
    .B(_948_),
    .Y(_949_)
);

NAND2X1 _4128_ (
    .A(_947_),
    .B(_949_),
    .Y(\z1.z3.z1.z2.s )
);

NOR2X1 _4129_ (
    .A(_946_),
    .B(_948_),
    .Y(\z1.z3.z1.z2.c )
);

AND2X2 _4130_ (
    .A(b[4]),
    .B(a[2]),
    .Y(\z1.z3.q1 [0])
);

AND2X2 _4131_ (
    .A(b[4]),
    .B(a[3]),
    .Y(\z1.z3.z2.z1.a )
);

AND2X2 _4132_ (
    .A(a[2]),
    .B(b[5]),
    .Y(\z1.z3.z2.z1.b )
);

AND2X2 _4133_ (
    .A(a[3]),
    .B(b[5]),
    .Y(\z1.z3.z2.z2.a )
);

INVX1 _4134_ (
    .A(\z1.z3.z2.z1.b ),
    .Y(_950_)
);

NAND2X1 _4135_ (
    .A(\z1.z3.z2.z1.a ),
    .B(_950_),
    .Y(_951_)
);

INVX1 _4136_ (
    .A(\z1.z3.z2.z1.a ),
    .Y(_952_)
);

NAND2X1 _4137_ (
    .A(\z1.z3.z2.z1.b ),
    .B(_952_),
    .Y(_953_)
);

NAND2X1 _4138_ (
    .A(_951_),
    .B(_953_),
    .Y(\z1.z3.z2.z1.s )
);

NOR2X1 _4139_ (
    .A(_950_),
    .B(_952_),
    .Y(\z1.z3.z2.z1.c )
);

INVX1 _4140_ (
    .A(\z1.z3.z2.z1.c ),
    .Y(_954_)
);

NAND2X1 _4141_ (
    .A(\z1.z3.z2.z2.a ),
    .B(_954_),
    .Y(_955_)
);

INVX1 _4142_ (
    .A(\z1.z3.z2.z2.a ),
    .Y(_956_)
);

NAND2X1 _4143_ (
    .A(\z1.z3.z2.z1.c ),
    .B(_956_),
    .Y(_957_)
);

NAND2X1 _4144_ (
    .A(_955_),
    .B(_957_),
    .Y(\z1.z3.z2.z2.s )
);

NOR2X1 _4145_ (
    .A(_954_),
    .B(_956_),
    .Y(\z1.z3.z2.z2.c )
);

AND2X2 _4146_ (
    .A(b[6]),
    .B(a[0]),
    .Y(\z1.z3.q2 [0])
);

AND2X2 _4147_ (
    .A(b[6]),
    .B(a[1]),
    .Y(\z1.z3.z3.z1.a )
);

AND2X2 _4148_ (
    .A(a[0]),
    .B(b[7]),
    .Y(\z1.z3.z3.z1.b )
);

AND2X2 _4149_ (
    .A(a[1]),
    .B(b[7]),
    .Y(\z1.z3.z3.z2.a )
);

INVX1 _4150_ (
    .A(\z1.z3.z3.z1.b ),
    .Y(_958_)
);

NAND2X1 _4151_ (
    .A(\z1.z3.z3.z1.a ),
    .B(_958_),
    .Y(_959_)
);

INVX1 _4152_ (
    .A(\z1.z3.z3.z1.a ),
    .Y(_960_)
);

NAND2X1 _4153_ (
    .A(\z1.z3.z3.z1.b ),
    .B(_960_),
    .Y(_961_)
);

NAND2X1 _4154_ (
    .A(_959_),
    .B(_961_),
    .Y(\z1.z3.z3.z1.s )
);

NOR2X1 _4155_ (
    .A(_958_),
    .B(_960_),
    .Y(\z1.z3.z3.z1.c )
);

INVX1 _4156_ (
    .A(\z1.z3.z3.z1.c ),
    .Y(_962_)
);

NAND2X1 _4157_ (
    .A(\z1.z3.z3.z2.a ),
    .B(_962_),
    .Y(_963_)
);

INVX1 _4158_ (
    .A(\z1.z3.z3.z2.a ),
    .Y(_964_)
);

NAND2X1 _4159_ (
    .A(\z1.z3.z3.z1.c ),
    .B(_964_),
    .Y(_965_)
);

NAND2X1 _4160_ (
    .A(_963_),
    .B(_965_),
    .Y(\z1.z3.z3.z2.s )
);

NOR2X1 _4161_ (
    .A(_962_),
    .B(_964_),
    .Y(\z1.z3.z3.z2.c )
);

AND2X2 _4162_ (
    .A(b[6]),
    .B(a[2]),
    .Y(\z1.z3.q3 [0])
);

AND2X2 _4163_ (
    .A(b[6]),
    .B(a[3]),
    .Y(\z1.z3.z4.z1.a )
);

AND2X2 _4164_ (
    .A(a[2]),
    .B(b[7]),
    .Y(\z1.z3.z4.z1.b )
);

AND2X2 _4165_ (
    .A(a[3]),
    .B(b[7]),
    .Y(\z1.z3.z4.z2.a )
);

INVX1 _4166_ (
    .A(\z1.z3.z4.z1.b ),
    .Y(_966_)
);

NAND2X1 _4167_ (
    .A(\z1.z3.z4.z1.a ),
    .B(_966_),
    .Y(_967_)
);

INVX1 _4168_ (
    .A(\z1.z3.z4.z1.a ),
    .Y(_968_)
);

NAND2X1 _4169_ (
    .A(\z1.z3.z4.z1.b ),
    .B(_968_),
    .Y(_969_)
);

NAND2X1 _4170_ (
    .A(_967_),
    .B(_969_),
    .Y(\z1.z3.z4.z1.s )
);

NOR2X1 _4171_ (
    .A(_966_),
    .B(_968_),
    .Y(\z1.z3.z4.z1.c )
);

INVX1 _4172_ (
    .A(\z1.z3.z4.z1.c ),
    .Y(_970_)
);

NAND2X1 _4173_ (
    .A(\z1.z3.z4.z2.a ),
    .B(_970_),
    .Y(_971_)
);

INVX1 _4174_ (
    .A(\z1.z3.z4.z2.a ),
    .Y(_972_)
);

NAND2X1 _4175_ (
    .A(\z1.z3.z4.z1.c ),
    .B(_972_),
    .Y(_973_)
);

NAND2X1 _4176_ (
    .A(_971_),
    .B(_973_),
    .Y(\z1.z3.z4.z2.s )
);

NOR2X1 _4177_ (
    .A(_970_),
    .B(_972_),
    .Y(\z1.z3.z4.z2.c )
);

NOR2X1 _4178_ (
    .A(\z1.z4.q1 [0]),
    .B(\z1.z4.z1.z2.s ),
    .Y(_981_)
);

AND2X2 _4179_ (
    .A(\z1.z4.q1 [0]),
    .B(\z1.z4.z1.z2.s ),
    .Y(_982_)
);

NOR2X1 _4180_ (
    .A(_981_),
    .B(_982_),
    .Y(_983_)
);

NAND2X1 _4181_ (
    .A(\z1.z4.q2 [0]),
    .B(_983_),
    .Y(_984_)
);

INVX1 _4182_ (
    .A(_984_),
    .Y(_985_)
);

NOR2X1 _4183_ (
    .A(\z1.z4.q2 [0]),
    .B(_983_),
    .Y(_986_)
);

NOR2X1 _4184_ (
    .A(_986_),
    .B(_985_),
    .Y(\z1.q3 [2])
);

NAND2X1 _4185_ (
    .A(\z1.z4.q1 [0]),
    .B(\z1.z4.z1.z2.s ),
    .Y(_987_)
);

NOR2X1 _4186_ (
    .A(\z1.z4.z2.z1.s ),
    .B(\z1.z4.z1.z2.c ),
    .Y(_988_)
);

NAND2X1 _4187_ (
    .A(\z1.z4.z2.z1.s ),
    .B(\z1.z4.z1.z2.c ),
    .Y(_989_)
);

INVX1 _4188_ (
    .A(_989_),
    .Y(_990_)
);

OAI21X1 _4189_ (
    .A(_988_),
    .B(_990_),
    .C(_987_),
    .Y(_991_)
);

INVX1 _4190_ (
    .A(\z1.z4.z2.z1.s ),
    .Y(_992_)
);

INVX1 _4191_ (
    .A(\z1.z4.z1.z2.c ),
    .Y(_993_)
);

NAND2X1 _4192_ (
    .A(_992_),
    .B(_993_),
    .Y(_994_)
);

NAND3X1 _4193_ (
    .A(_982_),
    .B(_989_),
    .C(_994_),
    .Y(_995_)
);

NAND3X1 _4194_ (
    .A(\z1.z4.z3.z1.s ),
    .B(_995_),
    .C(_991_),
    .Y(_996_)
);

INVX1 _4195_ (
    .A(\z1.z4.z3.z1.s ),
    .Y(_997_)
);

NAND2X1 _4196_ (
    .A(_995_),
    .B(_991_),
    .Y(_998_)
);

NAND2X1 _4197_ (
    .A(_997_),
    .B(_998_),
    .Y(_999_)
);

NAND3X1 _4198_ (
    .A(_985_),
    .B(_996_),
    .C(_999_),
    .Y(_1000_)
);

INVX1 _4199_ (
    .A(_1000_),
    .Y(_1001_)
);

INVX1 _4200_ (
    .A(_996_),
    .Y(_1002_)
);

OAI21X1 _4201_ (
    .A(_987_),
    .B(_988_),
    .C(_989_),
    .Y(_1003_)
);

NAND2X1 _4202_ (
    .A(\z1.z4.z2.z2.s ),
    .B(_1003_),
    .Y(_1004_)
);

INVX1 _4203_ (
    .A(\z1.z4.z2.z2.s ),
    .Y(_1005_)
);

NAND3X1 _4204_ (
    .A(_1005_),
    .B(_989_),
    .C(_995_),
    .Y(_1006_)
);

NAND2X1 _4205_ (
    .A(\z1.z4.q3 [0]),
    .B(\z1.z4.z3.z2.s ),
    .Y(_1007_)
);

INVX1 _4206_ (
    .A(\z1.z4.q3 [0]),
    .Y(_1008_)
);

INVX1 _4207_ (
    .A(\z1.z4.z3.z2.s ),
    .Y(_1009_)
);

NAND2X1 _4208_ (
    .A(_1008_),
    .B(_1009_),
    .Y(_1010_)
);

NAND2X1 _4209_ (
    .A(_1007_),
    .B(_1010_),
    .Y(_1011_)
);

INVX1 _4210_ (
    .A(_1011_),
    .Y(_1012_)
);

NAND3X1 _4211_ (
    .A(_1004_),
    .B(_1012_),
    .C(_1006_),
    .Y(_1013_)
);

AND2X2 _4212_ (
    .A(_1003_),
    .B(\z1.z4.z2.z2.s ),
    .Y(_1014_)
);

NOR2X1 _4213_ (
    .A(\z1.z4.z2.z2.s ),
    .B(_1003_),
    .Y(_1015_)
);

OAI21X1 _4214_ (
    .A(_1015_),
    .B(_1014_),
    .C(_1011_),
    .Y(_1016_)
);

NAND3X1 _4215_ (
    .A(_1002_),
    .B(_1013_),
    .C(_1016_),
    .Y(_1017_)
);

INVX1 _4216_ (
    .A(_1013_),
    .Y(_1018_)
);

AOI21X1 _4217_ (
    .A(_1006_),
    .B(_1004_),
    .C(_1012_),
    .Y(_1019_)
);

OAI21X1 _4218_ (
    .A(_1019_),
    .B(_1018_),
    .C(_996_),
    .Y(_1020_)
);

NAND3X1 _4219_ (
    .A(_1001_),
    .B(_1017_),
    .C(_1020_),
    .Y(_1021_)
);

INVX1 _4220_ (
    .A(_1017_),
    .Y(_1022_)
);

INVX1 _4221_ (
    .A(_998_),
    .Y(_1023_)
);

AOI22X1 _4222_ (
    .A(\z1.z4.z3.z1.s ),
    .B(_1023_),
    .C(_1016_),
    .D(_1013_),
    .Y(_1024_)
);

OAI21X1 _4223_ (
    .A(_1024_),
    .B(_1022_),
    .C(_1000_),
    .Y(_1025_)
);

AND2X2 _4224_ (
    .A(_1025_),
    .B(_1021_),
    .Y(\z1.q3 [4])
);

OAI21X1 _4225_ (
    .A(_1000_),
    .B(_1024_),
    .C(_1017_),
    .Y(_1026_)
);

OAI21X1 _4226_ (
    .A(_1008_),
    .B(_1009_),
    .C(_1013_),
    .Y(_1027_)
);

NAND2X1 _4227_ (
    .A(\z1.z4.z4.z1.s ),
    .B(\z1.z4.z3.z2.c ),
    .Y(_1028_)
);

OR2X2 _4228_ (
    .A(\z1.z4.z4.z1.s ),
    .B(\z1.z4.z3.z2.c ),
    .Y(_1029_)
);

NAND2X1 _4229_ (
    .A(_1028_),
    .B(_1029_),
    .Y(_1030_)
);

INVX1 _4230_ (
    .A(_1030_),
    .Y(_1031_)
);

NAND2X1 _4231_ (
    .A(\z1.z4.z2.z2.c ),
    .B(_1014_),
    .Y(_1032_)
);

INVX1 _4232_ (
    .A(\z1.z4.z2.z2.c ),
    .Y(_1033_)
);

NAND2X1 _4233_ (
    .A(_1033_),
    .B(_1004_),
    .Y(_1034_)
);

NAND3X1 _4234_ (
    .A(_1031_),
    .B(_1034_),
    .C(_1032_),
    .Y(_1035_)
);

NAND2X1 _4235_ (
    .A(\z1.z4.z2.z2.c ),
    .B(_1004_),
    .Y(_1036_)
);

NAND2X1 _4236_ (
    .A(_1033_),
    .B(_1014_),
    .Y(_1037_)
);

NAND3X1 _4237_ (
    .A(_1030_),
    .B(_1036_),
    .C(_1037_),
    .Y(_1038_)
);

NAND3X1 _4238_ (
    .A(_1027_),
    .B(_1035_),
    .C(_1038_),
    .Y(_1039_)
);

INVX1 _4239_ (
    .A(_1027_),
    .Y(_1040_)
);

AOI21X1 _4240_ (
    .A(_1037_),
    .B(_1036_),
    .C(_1030_),
    .Y(_1041_)
);

AOI21X1 _4241_ (
    .A(_1032_),
    .B(_1034_),
    .C(_1031_),
    .Y(_1042_)
);

OAI21X1 _4242_ (
    .A(_1041_),
    .B(_1042_),
    .C(_1040_),
    .Y(_1043_)
);

NAND2X1 _4243_ (
    .A(_1039_),
    .B(_1043_),
    .Y(_1044_)
);

NAND2X1 _4244_ (
    .A(_1026_),
    .B(_1044_),
    .Y(_1045_)
);

OR2X2 _4245_ (
    .A(_1044_),
    .B(_1026_),
    .Y(_1046_)
);

NAND2X1 _4246_ (
    .A(_1045_),
    .B(_1046_),
    .Y(\z1.q3 [5])
);

INVX1 _4247_ (
    .A(\z1.z4.z4.z2.s ),
    .Y(_1047_)
);

INVX1 _4248_ (
    .A(_1028_),
    .Y(_1048_)
);

OAI21X1 _4249_ (
    .A(_1048_),
    .B(_1041_),
    .C(_1047_),
    .Y(_1049_)
);

NAND3X1 _4250_ (
    .A(\z1.z4.z4.z2.s ),
    .B(_1028_),
    .C(_1035_),
    .Y(_1050_)
);

NAND2X1 _4251_ (
    .A(_1043_),
    .B(_1026_),
    .Y(_1051_)
);

AOI22X1 _4252_ (
    .A(_1049_),
    .B(_1050_),
    .C(_1051_),
    .D(_1039_),
    .Y(_1052_)
);

NAND2X1 _4253_ (
    .A(_1050_),
    .B(_1049_),
    .Y(_1053_)
);

NAND3X1 _4254_ (
    .A(_1017_),
    .B(_1039_),
    .C(_1021_),
    .Y(_1054_)
);

AOI21X1 _4255_ (
    .A(_1054_),
    .B(_1043_),
    .C(_1053_),
    .Y(_1055_)
);

NOR2X1 _4256_ (
    .A(_1052_),
    .B(_1055_),
    .Y(\z1.q3 [6])
);

OAI21X1 _4257_ (
    .A(_1048_),
    .B(_1041_),
    .C(\z1.z4.z4.z2.s ),
    .Y(_974_)
);

NAND3X1 _4258_ (
    .A(_1043_),
    .B(_1053_),
    .C(_1054_),
    .Y(_975_)
);

NAND3X1 _4259_ (
    .A(\z1.z4.z4.z2.c ),
    .B(_974_),
    .C(_975_),
    .Y(_976_)
);

INVX1 _4260_ (
    .A(\z1.z4.z4.z2.c ),
    .Y(_977_)
);

INVX1 _4261_ (
    .A(_974_),
    .Y(_978_)
);

OAI21X1 _4262_ (
    .A(_978_),
    .B(_1052_),
    .C(_977_),
    .Y(_979_)
);

NAND2X1 _4263_ (
    .A(_976_),
    .B(_979_),
    .Y(\z1.q3 [7])
);

AOI21X1 _4264_ (
    .A(_999_),
    .B(_996_),
    .C(_985_),
    .Y(_980_)
);

NOR2X1 _4265_ (
    .A(_980_),
    .B(_1001_),
    .Y(\z1.q3 [3])
);

AND2X2 _4266_ (
    .A(b[4]),
    .B(a[4]),
    .Y(\z1.q3 [0])
);

AND2X2 _4267_ (
    .A(b[4]),
    .B(a[5]),
    .Y(\z1.z4.z1.z1.a )
);

AND2X2 _4268_ (
    .A(a[4]),
    .B(b[5]),
    .Y(\z1.z4.z1.z1.b )
);

AND2X2 _4269_ (
    .A(a[5]),
    .B(b[5]),
    .Y(\z1.z4.z1.z2.a )
);

INVX1 _4270_ (
    .A(\z1.z4.z1.z1.b ),
    .Y(_1056_)
);

NAND2X1 _4271_ (
    .A(\z1.z4.z1.z1.a ),
    .B(_1056_),
    .Y(_1057_)
);

INVX1 _4272_ (
    .A(\z1.z4.z1.z1.a ),
    .Y(_1058_)
);

NAND2X1 _4273_ (
    .A(\z1.z4.z1.z1.b ),
    .B(_1058_),
    .Y(_1059_)
);

NAND2X1 _4274_ (
    .A(_1057_),
    .B(_1059_),
    .Y(\z1.z4.z1.z1.s )
);

NOR2X1 _4275_ (
    .A(_1056_),
    .B(_1058_),
    .Y(\z1.z4.z1.z1.c )
);

INVX1 _4276_ (
    .A(\z1.z4.z1.z1.c ),
    .Y(_1060_)
);

NAND2X1 _4277_ (
    .A(\z1.z4.z1.z2.a ),
    .B(_1060_),
    .Y(_1061_)
);

INVX1 _4278_ (
    .A(\z1.z4.z1.z2.a ),
    .Y(_1062_)
);

NAND2X1 _4279_ (
    .A(\z1.z4.z1.z1.c ),
    .B(_1062_),
    .Y(_1063_)
);

NAND2X1 _4280_ (
    .A(_1061_),
    .B(_1063_),
    .Y(\z1.z4.z1.z2.s )
);

NOR2X1 _4281_ (
    .A(_1060_),
    .B(_1062_),
    .Y(\z1.z4.z1.z2.c )
);

AND2X2 _4282_ (
    .A(b[4]),
    .B(a[6]),
    .Y(\z1.z4.q1 [0])
);

AND2X2 _4283_ (
    .A(b[4]),
    .B(a[7]),
    .Y(\z1.z4.z2.z1.a )
);

AND2X2 _4284_ (
    .A(a[6]),
    .B(b[5]),
    .Y(\z1.z4.z2.z1.b )
);

AND2X2 _4285_ (
    .A(a[7]),
    .B(b[5]),
    .Y(\z1.z4.z2.z2.a )
);

INVX1 _4286_ (
    .A(\z1.z4.z2.z1.b ),
    .Y(_1064_)
);

NAND2X1 _4287_ (
    .A(\z1.z4.z2.z1.a ),
    .B(_1064_),
    .Y(_1065_)
);

INVX1 _4288_ (
    .A(\z1.z4.z2.z1.a ),
    .Y(_1066_)
);

NAND2X1 _4289_ (
    .A(\z1.z4.z2.z1.b ),
    .B(_1066_),
    .Y(_1067_)
);

NAND2X1 _4290_ (
    .A(_1065_),
    .B(_1067_),
    .Y(\z1.z4.z2.z1.s )
);

NOR2X1 _4291_ (
    .A(_1064_),
    .B(_1066_),
    .Y(\z1.z4.z2.z1.c )
);

INVX1 _4292_ (
    .A(\z1.z4.z2.z1.c ),
    .Y(_1068_)
);

NAND2X1 _4293_ (
    .A(\z1.z4.z2.z2.a ),
    .B(_1068_),
    .Y(_1069_)
);

INVX1 _4294_ (
    .A(\z1.z4.z2.z2.a ),
    .Y(_1070_)
);

NAND2X1 _4295_ (
    .A(\z1.z4.z2.z1.c ),
    .B(_1070_),
    .Y(_1071_)
);

NAND2X1 _4296_ (
    .A(_1069_),
    .B(_1071_),
    .Y(\z1.z4.z2.z2.s )
);

NOR2X1 _4297_ (
    .A(_1068_),
    .B(_1070_),
    .Y(\z1.z4.z2.z2.c )
);

AND2X2 _4298_ (
    .A(b[6]),
    .B(a[4]),
    .Y(\z1.z4.q2 [0])
);

AND2X2 _4299_ (
    .A(b[6]),
    .B(a[5]),
    .Y(\z1.z4.z3.z1.a )
);

AND2X2 _4300_ (
    .A(a[4]),
    .B(b[7]),
    .Y(\z1.z4.z3.z1.b )
);

AND2X2 _4301_ (
    .A(a[5]),
    .B(b[7]),
    .Y(\z1.z4.z3.z2.a )
);

INVX1 _4302_ (
    .A(\z1.z4.z3.z1.b ),
    .Y(_1072_)
);

NAND2X1 _4303_ (
    .A(\z1.z4.z3.z1.a ),
    .B(_1072_),
    .Y(_1073_)
);

INVX1 _4304_ (
    .A(\z1.z4.z3.z1.a ),
    .Y(_1074_)
);

NAND2X1 _4305_ (
    .A(\z1.z4.z3.z1.b ),
    .B(_1074_),
    .Y(_1075_)
);

NAND2X1 _4306_ (
    .A(_1073_),
    .B(_1075_),
    .Y(\z1.z4.z3.z1.s )
);

NOR2X1 _4307_ (
    .A(_1072_),
    .B(_1074_),
    .Y(\z1.z4.z3.z1.c )
);

INVX1 _4308_ (
    .A(\z1.z4.z3.z1.c ),
    .Y(_1076_)
);

NAND2X1 _4309_ (
    .A(\z1.z4.z3.z2.a ),
    .B(_1076_),
    .Y(_1077_)
);

INVX1 _4310_ (
    .A(\z1.z4.z3.z2.a ),
    .Y(_1078_)
);

NAND2X1 _4311_ (
    .A(\z1.z4.z3.z1.c ),
    .B(_1078_),
    .Y(_1079_)
);

NAND2X1 _4312_ (
    .A(_1077_),
    .B(_1079_),
    .Y(\z1.z4.z3.z2.s )
);

NOR2X1 _4313_ (
    .A(_1076_),
    .B(_1078_),
    .Y(\z1.z4.z3.z2.c )
);

AND2X2 _4314_ (
    .A(b[6]),
    .B(a[6]),
    .Y(\z1.z4.q3 [0])
);

AND2X2 _4315_ (
    .A(b[6]),
    .B(a[7]),
    .Y(\z1.z4.z4.z1.a )
);

AND2X2 _4316_ (
    .A(a[6]),
    .B(b[7]),
    .Y(\z1.z4.z4.z1.b )
);

AND2X2 _4317_ (
    .A(a[7]),
    .B(b[7]),
    .Y(\z1.z4.z4.z2.a )
);

INVX1 _4318_ (
    .A(\z1.z4.z4.z1.b ),
    .Y(_1080_)
);

NAND2X1 _4319_ (
    .A(\z1.z4.z4.z1.a ),
    .B(_1080_),
    .Y(_1081_)
);

INVX1 _4320_ (
    .A(\z1.z4.z4.z1.a ),
    .Y(_1082_)
);

NAND2X1 _4321_ (
    .A(\z1.z4.z4.z1.b ),
    .B(_1082_),
    .Y(_1083_)
);

NAND2X1 _4322_ (
    .A(_1081_),
    .B(_1083_),
    .Y(\z1.z4.z4.z1.s )
);

NOR2X1 _4323_ (
    .A(_1080_),
    .B(_1082_),
    .Y(\z1.z4.z4.z1.c )
);

INVX1 _4324_ (
    .A(\z1.z4.z4.z1.c ),
    .Y(_1084_)
);

NAND2X1 _4325_ (
    .A(\z1.z4.z4.z2.a ),
    .B(_1084_),
    .Y(_1085_)
);

INVX1 _4326_ (
    .A(\z1.z4.z4.z2.a ),
    .Y(_1086_)
);

NAND2X1 _4327_ (
    .A(\z1.z4.z4.z1.c ),
    .B(_1086_),
    .Y(_1087_)
);

NAND2X1 _4328_ (
    .A(_1085_),
    .B(_1087_),
    .Y(\z1.z4.z4.z2.s )
);

NOR2X1 _4329_ (
    .A(_1084_),
    .B(_1086_),
    .Y(\z1.z4.z4.z2.c )
);

OR2X2 _4330_ (
    .A(\z2.q1 [0]),
    .B(\z2.q0 [4]),
    .Y(_1230_)
);

NAND2X1 _4331_ (
    .A(\z2.q1 [0]),
    .B(\z2.q0 [4]),
    .Y(_1231_)
);

NAND2X1 _4332_ (
    .A(_1231_),
    .B(_1230_),
    .Y(_1232_)
);

INVX1 _4333_ (
    .A(_1232_),
    .Y(_1233_)
);

AND2X2 _4334_ (
    .A(_1233_),
    .B(\z2.q2 [0]),
    .Y(_1234_)
);

NOR2X1 _4335_ (
    .A(\z2.q2 [0]),
    .B(_1233_),
    .Y(_1235_)
);

NOR2X1 _4336_ (
    .A(_1235_),
    .B(_1234_),
    .Y(q1[4])
);

INVX1 _4337_ (
    .A(\z2.z3.z1.z1.s ),
    .Y(_1236_)
);

INVX1 _4338_ (
    .A(_1231_),
    .Y(_1237_)
);

NAND2X1 _4339_ (
    .A(\z2.z2.z1.z1.s ),
    .B(\z2.q0 [5]),
    .Y(_1238_)
);

OR2X2 _4340_ (
    .A(\z2.z2.z1.z1.s ),
    .B(\z2.q0 [5]),
    .Y(_1239_)
);

NAND3X1 _4341_ (
    .A(_1238_),
    .B(_1239_),
    .C(_1237_),
    .Y(_1240_)
);

AND2X2 _4342_ (
    .A(\z2.z2.z1.z1.s ),
    .B(\z2.q0 [5]),
    .Y(_1241_)
);

NOR2X1 _4343_ (
    .A(\z2.z2.z1.z1.s ),
    .B(\z2.q0 [5]),
    .Y(_1242_)
);

OAI21X1 _4344_ (
    .A(_1242_),
    .B(_1241_),
    .C(_1231_),
    .Y(_1243_)
);

NAND2X1 _4345_ (
    .A(_1243_),
    .B(_1240_),
    .Y(_1244_)
);

OR2X2 _4346_ (
    .A(_1244_),
    .B(_1236_),
    .Y(_1245_)
);

NAND2X1 _4347_ (
    .A(_1236_),
    .B(_1244_),
    .Y(_1246_)
);

AND2X2 _4348_ (
    .A(_1245_),
    .B(_1246_),
    .Y(_1247_)
);

NAND2X1 _4349_ (
    .A(_1234_),
    .B(_1247_),
    .Y(_1248_)
);

INVX1 _4350_ (
    .A(_1245_),
    .Y(_1249_)
);

OAI21X1 _4351_ (
    .A(_1231_),
    .B(_1242_),
    .C(_1238_),
    .Y(_1250_)
);

INVX1 _4352_ (
    .A(\z2.q0 [6]),
    .Y(_1251_)
);

NOR2X1 _4353_ (
    .A(\z2.q1 [2]),
    .B(_1251_),
    .Y(_1252_)
);

INVX1 _4354_ (
    .A(\z2.q1 [2]),
    .Y(_1253_)
);

NOR2X1 _4355_ (
    .A(\z2.q0 [6]),
    .B(_1253_),
    .Y(_1254_)
);

OAI21X1 _4356_ (
    .A(_1252_),
    .B(_1254_),
    .C(_1250_),
    .Y(_1255_)
);

NAND2X1 _4357_ (
    .A(\z2.q0 [6]),
    .B(_1253_),
    .Y(_1256_)
);

NAND2X1 _4358_ (
    .A(\z2.q1 [2]),
    .B(_1251_),
    .Y(_1257_)
);

NAND2X1 _4359_ (
    .A(_1256_),
    .B(_1257_),
    .Y(_1258_)
);

OR2X2 _4360_ (
    .A(_1258_),
    .B(_1250_),
    .Y(_1259_)
);

NAND3X1 _4361_ (
    .A(\z2.q2 [2]),
    .B(_1255_),
    .C(_1259_),
    .Y(_1260_)
);

INVX1 _4362_ (
    .A(\z2.q2 [2]),
    .Y(_1261_)
);

NAND2X1 _4363_ (
    .A(_1255_),
    .B(_1259_),
    .Y(_1262_)
);

NAND2X1 _4364_ (
    .A(_1261_),
    .B(_1262_),
    .Y(_1263_)
);

AOI21X1 _4365_ (
    .A(_1263_),
    .B(_1260_),
    .C(_1249_),
    .Y(_1264_)
);

INVX1 _4366_ (
    .A(_1264_),
    .Y(_1265_)
);

NAND3X1 _4367_ (
    .A(_1260_),
    .B(_1263_),
    .C(_1249_),
    .Y(_1266_)
);

NAND3X1 _4368_ (
    .A(_1248_),
    .B(_1266_),
    .C(_1265_),
    .Y(_1267_)
);

INVX1 _4369_ (
    .A(_1248_),
    .Y(_1268_)
);

INVX1 _4370_ (
    .A(_1266_),
    .Y(_1269_)
);

OAI21X1 _4371_ (
    .A(_1264_),
    .B(_1269_),
    .C(_1268_),
    .Y(_1270_)
);

NAND2X1 _4372_ (
    .A(_1267_),
    .B(_1270_),
    .Y(q1[6])
);

OAI21X1 _4373_ (
    .A(_1264_),
    .B(_1248_),
    .C(_1266_),
    .Y(_1271_)
);

INVX1 _4374_ (
    .A(_1260_),
    .Y(_1272_)
);

INVX1 _4375_ (
    .A(\z2.q2 [3]),
    .Y(_1273_)
);

INVX1 _4376_ (
    .A(\z2.q0 [7]),
    .Y(_1274_)
);

NOR2X1 _4377_ (
    .A(\z2.q1 [3]),
    .B(_1274_),
    .Y(_1275_)
);

INVX1 _4378_ (
    .A(\z2.q1 [3]),
    .Y(_1276_)
);

NOR2X1 _4379_ (
    .A(\z2.q0 [7]),
    .B(_1276_),
    .Y(_1277_)
);

NAND2X1 _4380_ (
    .A(\z2.q1 [2]),
    .B(\z2.q0 [6]),
    .Y(_1278_)
);

INVX1 _4381_ (
    .A(_1278_),
    .Y(_1279_)
);

AOI21X1 _4382_ (
    .A(_1258_),
    .B(_1250_),
    .C(_1279_),
    .Y(_1280_)
);

OAI21X1 _4383_ (
    .A(_1275_),
    .B(_1277_),
    .C(_1280_),
    .Y(_1281_)
);

NAND2X1 _4384_ (
    .A(\z2.q1 [3]),
    .B(\z2.q0 [7]),
    .Y(_1282_)
);

INVX1 _4385_ (
    .A(_1282_),
    .Y(_1283_)
);

NOR2X1 _4386_ (
    .A(\z2.q1 [3]),
    .B(\z2.q0 [7]),
    .Y(_1284_)
);

INVX1 _4387_ (
    .A(_1280_),
    .Y(_1285_)
);

OAI21X1 _4388_ (
    .A(_1283_),
    .B(_1284_),
    .C(_1285_),
    .Y(_1286_)
);

AOI21X1 _4389_ (
    .A(_1286_),
    .B(_1281_),
    .C(_1273_),
    .Y(_1088_)
);

INVX1 _4390_ (
    .A(_1088_),
    .Y(_1089_)
);

NAND3X1 _4391_ (
    .A(_1273_),
    .B(_1281_),
    .C(_1286_),
    .Y(_1090_)
);

AOI21X1 _4392_ (
    .A(_1089_),
    .B(_1090_),
    .C(_1272_),
    .Y(_1091_)
);

NAND3X1 _4393_ (
    .A(_1272_),
    .B(_1090_),
    .C(_1089_),
    .Y(_1092_)
);

INVX1 _4394_ (
    .A(_1092_),
    .Y(_1093_)
);

OAI21X1 _4395_ (
    .A(_1091_),
    .B(_1093_),
    .C(_1271_),
    .Y(_1094_)
);

INVX1 _4396_ (
    .A(_1271_),
    .Y(_1095_)
);

NAND2X1 _4397_ (
    .A(_1090_),
    .B(_1089_),
    .Y(_1096_)
);

OAI21X1 _4398_ (
    .A(_1261_),
    .B(_1262_),
    .C(_1096_),
    .Y(_1097_)
);

NAND3X1 _4399_ (
    .A(_1092_),
    .B(_1095_),
    .C(_1097_),
    .Y(_1098_)
);

NAND2X1 _4400_ (
    .A(_1098_),
    .B(_1094_),
    .Y(q1[7])
);

AOI21X1 _4401_ (
    .A(_1097_),
    .B(_1271_),
    .C(_1093_),
    .Y(_1099_)
);

AOI21X1 _4402_ (
    .A(_1237_),
    .B(_1239_),
    .C(_1241_),
    .Y(_1100_)
);

OAI22X1 _4403_ (
    .A(_1252_),
    .B(_1254_),
    .C(_1275_),
    .D(_1277_),
    .Y(_1101_)
);

OAI21X1 _4404_ (
    .A(_1278_),
    .B(_1284_),
    .C(_1282_),
    .Y(_1102_)
);

INVX1 _4405_ (
    .A(_1102_),
    .Y(_1103_)
);

OAI21X1 _4406_ (
    .A(_1100_),
    .B(_1101_),
    .C(_1103_),
    .Y(_1104_)
);

NAND2X1 _4407_ (
    .A(\z2.q1 [4]),
    .B(_1104_),
    .Y(_1105_)
);

INVX1 _4408_ (
    .A(\z2.q1 [4]),
    .Y(_1106_)
);

NAND2X1 _4409_ (
    .A(\z2.q0 [7]),
    .B(_1276_),
    .Y(_1107_)
);

NAND2X1 _4410_ (
    .A(\z2.q1 [3]),
    .B(_1274_),
    .Y(_1108_)
);

NAND2X1 _4411_ (
    .A(_1107_),
    .B(_1108_),
    .Y(_1109_)
);

NAND3X1 _4412_ (
    .A(_1250_),
    .B(_1258_),
    .C(_1109_),
    .Y(_1110_)
);

NAND3X1 _4413_ (
    .A(_1106_),
    .B(_1103_),
    .C(_1110_),
    .Y(_1111_)
);

NAND2X1 _4414_ (
    .A(\z2.q3 [0]),
    .B(\z2.q2 [4]),
    .Y(_1112_)
);

INVX1 _4415_ (
    .A(\z2.q3 [0]),
    .Y(_1113_)
);

INVX1 _4416_ (
    .A(\z2.q2 [4]),
    .Y(_1114_)
);

NAND2X1 _4417_ (
    .A(_1113_),
    .B(_1114_),
    .Y(_1115_)
);

NAND2X1 _4418_ (
    .A(_1112_),
    .B(_1115_),
    .Y(_1116_)
);

INVX1 _4419_ (
    .A(_1116_),
    .Y(_1117_)
);

NAND3X1 _4420_ (
    .A(_1111_),
    .B(_1117_),
    .C(_1105_),
    .Y(_1118_)
);

AOI21X1 _4421_ (
    .A(_1110_),
    .B(_1103_),
    .C(_1106_),
    .Y(_1119_)
);

INVX1 _4422_ (
    .A(_1111_),
    .Y(_1120_)
);

OAI21X1 _4423_ (
    .A(_1119_),
    .B(_1120_),
    .C(_1116_),
    .Y(_1121_)
);

NAND3X1 _4424_ (
    .A(_1118_),
    .B(_1121_),
    .C(_1088_),
    .Y(_1122_)
);

NAND2X1 _4425_ (
    .A(_1118_),
    .B(_1121_),
    .Y(_1123_)
);

NAND2X1 _4426_ (
    .A(_1123_),
    .B(_1089_),
    .Y(_1124_)
);

AND2X2 _4427_ (
    .A(_1124_),
    .B(_1122_),
    .Y(_1125_)
);

NAND2X1 _4428_ (
    .A(_1125_),
    .B(_1099_),
    .Y(_1126_)
);

OAI21X1 _4429_ (
    .A(_1091_),
    .B(_1095_),
    .C(_1092_),
    .Y(_1127_)
);

NAND2X1 _4430_ (
    .A(_1122_),
    .B(_1124_),
    .Y(_1128_)
);

NAND2X1 _4431_ (
    .A(_1128_),
    .B(_1127_),
    .Y(_1129_)
);

NAND2X1 _4432_ (
    .A(_1126_),
    .B(_1129_),
    .Y(q1[8])
);

OAI21X1 _4433_ (
    .A(_1128_),
    .B(_1099_),
    .C(_1122_),
    .Y(_1130_)
);

OAI21X1 _4434_ (
    .A(_1113_),
    .B(_1114_),
    .C(_1118_),
    .Y(_1131_)
);

NAND3X1 _4435_ (
    .A(\z2.q1 [4]),
    .B(\z2.q1 [5]),
    .C(_1104_),
    .Y(_1132_)
);

INVX1 _4436_ (
    .A(\z2.q1 [5]),
    .Y(_1133_)
);

AOI22X1 _4437_ (
    .A(_1256_),
    .B(_1257_),
    .C(_1107_),
    .D(_1108_),
    .Y(_1134_)
);

AOI21X1 _4438_ (
    .A(_1134_),
    .B(_1250_),
    .C(_1102_),
    .Y(_1135_)
);

OAI21X1 _4439_ (
    .A(_1106_),
    .B(_1135_),
    .C(_1133_),
    .Y(_1136_)
);

INVX1 _4440_ (
    .A(\z2.z4.z1.z1.s ),
    .Y(_1137_)
);

INVX1 _4441_ (
    .A(\z2.q2 [5]),
    .Y(_1138_)
);

NAND2X1 _4442_ (
    .A(_1137_),
    .B(_1138_),
    .Y(_1139_)
);

NAND2X1 _4443_ (
    .A(\z2.z4.z1.z1.s ),
    .B(\z2.q2 [5]),
    .Y(_1140_)
);

AND2X2 _4444_ (
    .A(_1139_),
    .B(_1140_),
    .Y(_1141_)
);

NAND3X1 _4445_ (
    .A(_1141_),
    .B(_1136_),
    .C(_1132_),
    .Y(_1142_)
);

AOI21X1 _4446_ (
    .A(_1132_),
    .B(_1136_),
    .C(_1141_),
    .Y(_1143_)
);

INVX1 _4447_ (
    .A(_1143_),
    .Y(_1144_)
);

NAND3X1 _4448_ (
    .A(_1142_),
    .B(_1131_),
    .C(_1144_),
    .Y(_1145_)
);

AND2X2 _4449_ (
    .A(_1118_),
    .B(_1112_),
    .Y(_1146_)
);

INVX1 _4450_ (
    .A(_1142_),
    .Y(_1147_)
);

OAI21X1 _4451_ (
    .A(_1147_),
    .B(_1143_),
    .C(_1146_),
    .Y(_1148_)
);

NAND2X1 _4452_ (
    .A(_1145_),
    .B(_1148_),
    .Y(_1149_)
);

OR2X2 _4453_ (
    .A(_1130_),
    .B(_1149_),
    .Y(_1150_)
);

NAND2X1 _4454_ (
    .A(_1149_),
    .B(_1130_),
    .Y(_1151_)
);

NAND2X1 _4455_ (
    .A(_1151_),
    .B(_1150_),
    .Y(q1[9])
);

NAND3X1 _4456_ (
    .A(_1145_),
    .B(_1148_),
    .C(_1125_),
    .Y(_1152_)
);

OAI21X1 _4457_ (
    .A(_1089_),
    .B(_1123_),
    .C(_1145_),
    .Y(_1153_)
);

NAND2X1 _4458_ (
    .A(_1148_),
    .B(_1153_),
    .Y(_1154_)
);

OAI21X1 _4459_ (
    .A(_1099_),
    .B(_1152_),
    .C(_1154_),
    .Y(_1155_)
);

OAI21X1 _4460_ (
    .A(_1137_),
    .B(_1138_),
    .C(_1142_),
    .Y(_1156_)
);

NAND3X1 _4461_ (
    .A(\z2.q1 [5]),
    .B(\z2.q1 [6]),
    .C(_1119_),
    .Y(_1157_)
);

INVX1 _4462_ (
    .A(\z2.q1 [6]),
    .Y(_1158_)
);

NAND2X1 _4463_ (
    .A(_1158_),
    .B(_1132_),
    .Y(_1159_)
);

INVX1 _4464_ (
    .A(\z2.q3 [2]),
    .Y(_1160_)
);

INVX1 _4465_ (
    .A(\z2.q2 [6]),
    .Y(_1161_)
);

NAND2X1 _4466_ (
    .A(_1160_),
    .B(_1161_),
    .Y(_1162_)
);

NAND2X1 _4467_ (
    .A(\z2.q3 [2]),
    .B(\z2.q2 [6]),
    .Y(_1163_)
);

NAND2X1 _4468_ (
    .A(_1163_),
    .B(_1162_),
    .Y(_1164_)
);

INVX1 _4469_ (
    .A(_1164_),
    .Y(_1165_)
);

NAND3X1 _4470_ (
    .A(_1157_),
    .B(_1165_),
    .C(_1159_),
    .Y(_1166_)
);

AOI21X1 _4471_ (
    .A(_1159_),
    .B(_1157_),
    .C(_1165_),
    .Y(_1167_)
);

INVX1 _4472_ (
    .A(_1167_),
    .Y(_1168_)
);

NAND3X1 _4473_ (
    .A(_1156_),
    .B(_1166_),
    .C(_1168_),
    .Y(_1169_)
);

INVX1 _4474_ (
    .A(_1156_),
    .Y(_1170_)
);

INVX1 _4475_ (
    .A(_1166_),
    .Y(_1171_)
);

OAI21X1 _4476_ (
    .A(_1167_),
    .B(_1171_),
    .C(_1170_),
    .Y(_1172_)
);

NAND2X1 _4477_ (
    .A(_1172_),
    .B(_1169_),
    .Y(_1173_)
);

NAND2X1 _4478_ (
    .A(_1173_),
    .B(_1155_),
    .Y(_1174_)
);

NOR2X1 _4479_ (
    .A(_1128_),
    .B(_1149_),
    .Y(_1175_)
);

AOI22X1 _4480_ (
    .A(_1148_),
    .B(_1153_),
    .C(_1175_),
    .D(_1127_),
    .Y(_1176_)
);

AND2X2 _4481_ (
    .A(_1169_),
    .B(_1172_),
    .Y(_1177_)
);

NAND2X1 _4482_ (
    .A(_1177_),
    .B(_1176_),
    .Y(_1178_)
);

NAND2X1 _4483_ (
    .A(_1174_),
    .B(_1178_),
    .Y(q1[10])
);

OAI21X1 _4484_ (
    .A(_1173_),
    .B(_1176_),
    .C(_1169_),
    .Y(_1179_)
);

OAI21X1 _4485_ (
    .A(_1160_),
    .B(_1161_),
    .C(_1166_),
    .Y(_1180_)
);

NOR2X1 _4486_ (
    .A(\z2.q3 [3]),
    .B(\z2.q2 [7]),
    .Y(_1181_)
);

INVX1 _4487_ (
    .A(\z2.q3 [3]),
    .Y(_1182_)
);

INVX1 _4488_ (
    .A(\z2.q2 [7]),
    .Y(_1183_)
);

NOR2X1 _4489_ (
    .A(_1182_),
    .B(_1183_),
    .Y(_1184_)
);

NOR2X1 _4490_ (
    .A(_1181_),
    .B(_1184_),
    .Y(_1185_)
);

INVX1 _4491_ (
    .A(\z2.q1 [7]),
    .Y(_1186_)
);

OAI21X1 _4492_ (
    .A(_1158_),
    .B(_1132_),
    .C(_1186_),
    .Y(_1187_)
);

AND2X2 _4493_ (
    .A(_1119_),
    .B(\z2.q1 [5]),
    .Y(_1188_)
);

NAND3X1 _4494_ (
    .A(\z2.q1 [6]),
    .B(\z2.q1 [7]),
    .C(_1188_),
    .Y(_1189_)
);

NAND3X1 _4495_ (
    .A(_1185_),
    .B(_1187_),
    .C(_1189_),
    .Y(_1190_)
);

INVX1 _4496_ (
    .A(_1185_),
    .Y(_1191_)
);

OAI21X1 _4497_ (
    .A(_1158_),
    .B(_1132_),
    .C(\z2.q1 [7]),
    .Y(_1192_)
);

NAND3X1 _4498_ (
    .A(\z2.q1 [6]),
    .B(_1186_),
    .C(_1188_),
    .Y(_1193_)
);

NAND3X1 _4499_ (
    .A(_1191_),
    .B(_1192_),
    .C(_1193_),
    .Y(_1194_)
);

NAND3X1 _4500_ (
    .A(_1190_),
    .B(_1194_),
    .C(_1180_),
    .Y(_1195_)
);

AND2X2 _4501_ (
    .A(_1166_),
    .B(_1163_),
    .Y(_1196_)
);

NAND2X1 _4502_ (
    .A(_1190_),
    .B(_1194_),
    .Y(_1197_)
);

NAND2X1 _4503_ (
    .A(_1196_),
    .B(_1197_),
    .Y(_1198_)
);

NAND2X1 _4504_ (
    .A(_1195_),
    .B(_1198_),
    .Y(_1199_)
);

OR2X2 _4505_ (
    .A(_1179_),
    .B(_1199_),
    .Y(_1200_)
);

NAND2X1 _4506_ (
    .A(_1199_),
    .B(_1179_),
    .Y(_1201_)
);

NAND2X1 _4507_ (
    .A(_1201_),
    .B(_1200_),
    .Y(q1[11])
);

OAI21X1 _4508_ (
    .A(_1196_),
    .B(_1197_),
    .C(_1169_),
    .Y(_1202_)
);

NAND2X1 _4509_ (
    .A(_1198_),
    .B(_1202_),
    .Y(_1203_)
);

NAND3X1 _4510_ (
    .A(_1195_),
    .B(_1198_),
    .C(_1177_),
    .Y(_1204_)
);

OAI21X1 _4511_ (
    .A(_1204_),
    .B(_1176_),
    .C(_1203_),
    .Y(_1205_)
);

OAI21X1 _4512_ (
    .A(_1182_),
    .B(_1183_),
    .C(_1190_),
    .Y(_1206_)
);

NAND2X1 _4513_ (
    .A(\z2.q3 [4]),
    .B(_1206_),
    .Y(_1207_)
);

OR2X2 _4514_ (
    .A(_1206_),
    .B(\z2.q3 [4]),
    .Y(_1208_)
);

NAND3X1 _4515_ (
    .A(_1207_),
    .B(_1208_),
    .C(_1205_),
    .Y(_1209_)
);

NOR2X1 _4516_ (
    .A(_1173_),
    .B(_1199_),
    .Y(_1210_)
);

AOI22X1 _4517_ (
    .A(_1198_),
    .B(_1202_),
    .C(_1210_),
    .D(_1155_),
    .Y(_1211_)
);

NAND2X1 _4518_ (
    .A(_1207_),
    .B(_1208_),
    .Y(_1212_)
);

NAND2X1 _4519_ (
    .A(_1212_),
    .B(_1211_),
    .Y(_1213_)
);

AND2X2 _4520_ (
    .A(_1209_),
    .B(_1213_),
    .Y(q1[12])
);

INVX1 _4521_ (
    .A(\z2.q3 [5]),
    .Y(_1214_)
);

OAI21X1 _4522_ (
    .A(_1212_),
    .B(_1211_),
    .C(_1207_),
    .Y(_1215_)
);

NAND2X1 _4523_ (
    .A(_1214_),
    .B(_1215_),
    .Y(_1216_)
);

NAND3X1 _4524_ (
    .A(\z2.q3 [5]),
    .B(_1207_),
    .C(_1209_),
    .Y(_1217_)
);

NAND2X1 _4525_ (
    .A(_1217_),
    .B(_1216_),
    .Y(q1[13])
);

INVX1 _4526_ (
    .A(\z2.q3 [6]),
    .Y(_1218_)
);

NAND3X1 _4527_ (
    .A(\z2.q3 [5]),
    .B(_1207_),
    .C(_1208_),
    .Y(_1219_)
);

OAI22X1 _4528_ (
    .A(_1214_),
    .B(_1207_),
    .C(_1219_),
    .D(_1211_),
    .Y(_1220_)
);

NAND2X1 _4529_ (
    .A(_1218_),
    .B(_1220_),
    .Y(_1221_)
);

INVX1 _4530_ (
    .A(_1207_),
    .Y(_1222_)
);

INVX1 _4531_ (
    .A(_1219_),
    .Y(_1223_)
);

AOI22X1 _4532_ (
    .A(\z2.q3 [5]),
    .B(_1222_),
    .C(_1205_),
    .D(_1223_),
    .Y(_1224_)
);

NAND2X1 _4533_ (
    .A(\z2.q3 [6]),
    .B(_1224_),
    .Y(_1225_)
);

NAND2X1 _4534_ (
    .A(_1225_),
    .B(_1221_),
    .Y(q1[14])
);

OAI21X1 _4535_ (
    .A(_1218_),
    .B(_1224_),
    .C(\z2.q3 [7]),
    .Y(_1226_)
);

INVX1 _4536_ (
    .A(\z2.q3 [7]),
    .Y(_1227_)
);

NAND3X1 _4537_ (
    .A(\z2.q3 [6]),
    .B(_1227_),
    .C(_1220_),
    .Y(_1228_)
);

NAND2X1 _4538_ (
    .A(_1228_),
    .B(_1226_),
    .Y(q1[15])
);

NOR2X1 _4539_ (
    .A(_1234_),
    .B(_1247_),
    .Y(_1229_)
);

NOR2X1 _4540_ (
    .A(_1229_),
    .B(_1268_),
    .Y(q1[5])
);

NOR2X1 _4541_ (
    .A(\z2.z1.q1 [0]),
    .B(\z2.z1.z1.z2.s ),
    .Y(_1294_)
);

AND2X2 _4542_ (
    .A(\z2.z1.q1 [0]),
    .B(\z2.z1.z1.z2.s ),
    .Y(_1295_)
);

NOR2X1 _4543_ (
    .A(_1294_),
    .B(_1295_),
    .Y(_1296_)
);

NAND2X1 _4544_ (
    .A(\z2.z1.q2 [0]),
    .B(_1296_),
    .Y(_1297_)
);

INVX1 _4545_ (
    .A(_1297_),
    .Y(_1298_)
);

NOR2X1 _4546_ (
    .A(\z2.z1.q2 [0]),
    .B(_1296_),
    .Y(_1299_)
);

NOR2X1 _4547_ (
    .A(_1299_),
    .B(_1298_),
    .Y(q1[2])
);

NAND2X1 _4548_ (
    .A(\z2.z1.q1 [0]),
    .B(\z2.z1.z1.z2.s ),
    .Y(_1300_)
);

NOR2X1 _4549_ (
    .A(\z2.z1.z2.z1.s ),
    .B(\z2.z1.z1.z2.c ),
    .Y(_1301_)
);

NAND2X1 _4550_ (
    .A(\z2.z1.z2.z1.s ),
    .B(\z2.z1.z1.z2.c ),
    .Y(_1302_)
);

INVX1 _4551_ (
    .A(_1302_),
    .Y(_1303_)
);

OAI21X1 _4552_ (
    .A(_1301_),
    .B(_1303_),
    .C(_1300_),
    .Y(_1304_)
);

INVX1 _4553_ (
    .A(\z2.z1.z2.z1.s ),
    .Y(_1305_)
);

INVX1 _4554_ (
    .A(\z2.z1.z1.z2.c ),
    .Y(_1306_)
);

NAND2X1 _4555_ (
    .A(_1305_),
    .B(_1306_),
    .Y(_1307_)
);

NAND3X1 _4556_ (
    .A(_1295_),
    .B(_1302_),
    .C(_1307_),
    .Y(_1308_)
);

NAND3X1 _4557_ (
    .A(\z2.z1.z3.z1.s ),
    .B(_1308_),
    .C(_1304_),
    .Y(_1309_)
);

INVX1 _4558_ (
    .A(\z2.z1.z3.z1.s ),
    .Y(_1310_)
);

NAND2X1 _4559_ (
    .A(_1308_),
    .B(_1304_),
    .Y(_1311_)
);

NAND2X1 _4560_ (
    .A(_1310_),
    .B(_1311_),
    .Y(_1312_)
);

NAND3X1 _4561_ (
    .A(_1298_),
    .B(_1309_),
    .C(_1312_),
    .Y(_1313_)
);

INVX1 _4562_ (
    .A(_1313_),
    .Y(_1314_)
);

INVX1 _4563_ (
    .A(_1309_),
    .Y(_1315_)
);

OAI21X1 _4564_ (
    .A(_1300_),
    .B(_1301_),
    .C(_1302_),
    .Y(_1316_)
);

NAND2X1 _4565_ (
    .A(\z2.z1.z2.z2.s ),
    .B(_1316_),
    .Y(_1317_)
);

INVX1 _4566_ (
    .A(\z2.z1.z2.z2.s ),
    .Y(_1318_)
);

NAND3X1 _4567_ (
    .A(_1318_),
    .B(_1302_),
    .C(_1308_),
    .Y(_1319_)
);

NAND2X1 _4568_ (
    .A(\z2.z1.q3 [0]),
    .B(\z2.z1.z3.z2.s ),
    .Y(_1320_)
);

INVX1 _4569_ (
    .A(\z2.z1.q3 [0]),
    .Y(_1321_)
);

INVX1 _4570_ (
    .A(\z2.z1.z3.z2.s ),
    .Y(_1322_)
);

NAND2X1 _4571_ (
    .A(_1321_),
    .B(_1322_),
    .Y(_1323_)
);

NAND2X1 _4572_ (
    .A(_1320_),
    .B(_1323_),
    .Y(_1324_)
);

INVX1 _4573_ (
    .A(_1324_),
    .Y(_1325_)
);

NAND3X1 _4574_ (
    .A(_1317_),
    .B(_1325_),
    .C(_1319_),
    .Y(_1326_)
);

AND2X2 _4575_ (
    .A(_1316_),
    .B(\z2.z1.z2.z2.s ),
    .Y(_1327_)
);

NOR2X1 _4576_ (
    .A(\z2.z1.z2.z2.s ),
    .B(_1316_),
    .Y(_1328_)
);

OAI21X1 _4577_ (
    .A(_1328_),
    .B(_1327_),
    .C(_1324_),
    .Y(_1329_)
);

NAND3X1 _4578_ (
    .A(_1315_),
    .B(_1326_),
    .C(_1329_),
    .Y(_1330_)
);

INVX1 _4579_ (
    .A(_1326_),
    .Y(_1331_)
);

AOI21X1 _4580_ (
    .A(_1319_),
    .B(_1317_),
    .C(_1325_),
    .Y(_1332_)
);

OAI21X1 _4581_ (
    .A(_1332_),
    .B(_1331_),
    .C(_1309_),
    .Y(_1333_)
);

NAND3X1 _4582_ (
    .A(_1314_),
    .B(_1330_),
    .C(_1333_),
    .Y(_1334_)
);

INVX1 _4583_ (
    .A(_1330_),
    .Y(_1335_)
);

INVX1 _4584_ (
    .A(_1311_),
    .Y(_1336_)
);

AOI22X1 _4585_ (
    .A(\z2.z1.z3.z1.s ),
    .B(_1336_),
    .C(_1329_),
    .D(_1326_),
    .Y(_1337_)
);

OAI21X1 _4586_ (
    .A(_1337_),
    .B(_1335_),
    .C(_1313_),
    .Y(_1338_)
);

AND2X2 _4587_ (
    .A(_1338_),
    .B(_1334_),
    .Y(\z2.q0 [4])
);

OAI21X1 _4588_ (
    .A(_1313_),
    .B(_1337_),
    .C(_1330_),
    .Y(_1339_)
);

OAI21X1 _4589_ (
    .A(_1321_),
    .B(_1322_),
    .C(_1326_),
    .Y(_1340_)
);

NAND2X1 _4590_ (
    .A(\z2.z1.z4.z1.s ),
    .B(\z2.z1.z3.z2.c ),
    .Y(_1341_)
);

OR2X2 _4591_ (
    .A(\z2.z1.z4.z1.s ),
    .B(\z2.z1.z3.z2.c ),
    .Y(_1342_)
);

NAND2X1 _4592_ (
    .A(_1341_),
    .B(_1342_),
    .Y(_1343_)
);

INVX1 _4593_ (
    .A(_1343_),
    .Y(_1344_)
);

NAND2X1 _4594_ (
    .A(\z2.z1.z2.z2.c ),
    .B(_1327_),
    .Y(_1345_)
);

INVX1 _4595_ (
    .A(\z2.z1.z2.z2.c ),
    .Y(_1346_)
);

NAND2X1 _4596_ (
    .A(_1346_),
    .B(_1317_),
    .Y(_1347_)
);

NAND3X1 _4597_ (
    .A(_1344_),
    .B(_1347_),
    .C(_1345_),
    .Y(_1348_)
);

NAND2X1 _4598_ (
    .A(\z2.z1.z2.z2.c ),
    .B(_1317_),
    .Y(_1349_)
);

NAND2X1 _4599_ (
    .A(_1346_),
    .B(_1327_),
    .Y(_1350_)
);

NAND3X1 _4600_ (
    .A(_1343_),
    .B(_1349_),
    .C(_1350_),
    .Y(_1351_)
);

NAND3X1 _4601_ (
    .A(_1340_),
    .B(_1348_),
    .C(_1351_),
    .Y(_1352_)
);

INVX1 _4602_ (
    .A(_1340_),
    .Y(_1353_)
);

AOI21X1 _4603_ (
    .A(_1350_),
    .B(_1349_),
    .C(_1343_),
    .Y(_1354_)
);

AOI21X1 _4604_ (
    .A(_1345_),
    .B(_1347_),
    .C(_1344_),
    .Y(_1355_)
);

OAI21X1 _4605_ (
    .A(_1354_),
    .B(_1355_),
    .C(_1353_),
    .Y(_1356_)
);

NAND2X1 _4606_ (
    .A(_1352_),
    .B(_1356_),
    .Y(_1357_)
);

NAND2X1 _4607_ (
    .A(_1339_),
    .B(_1357_),
    .Y(_1358_)
);

OR2X2 _4608_ (
    .A(_1357_),
    .B(_1339_),
    .Y(_1359_)
);

NAND2X1 _4609_ (
    .A(_1358_),
    .B(_1359_),
    .Y(\z2.q0 [5])
);

INVX1 _4610_ (
    .A(\z2.z1.z4.z2.s ),
    .Y(_1360_)
);

INVX1 _4611_ (
    .A(_1341_),
    .Y(_1361_)
);

OAI21X1 _4612_ (
    .A(_1361_),
    .B(_1354_),
    .C(_1360_),
    .Y(_1362_)
);

NAND3X1 _4613_ (
    .A(\z2.z1.z4.z2.s ),
    .B(_1341_),
    .C(_1348_),
    .Y(_1363_)
);

NAND2X1 _4614_ (
    .A(_1356_),
    .B(_1339_),
    .Y(_1364_)
);

AOI22X1 _4615_ (
    .A(_1362_),
    .B(_1363_),
    .C(_1364_),
    .D(_1352_),
    .Y(_1365_)
);

NAND2X1 _4616_ (
    .A(_1363_),
    .B(_1362_),
    .Y(_1366_)
);

NAND3X1 _4617_ (
    .A(_1330_),
    .B(_1352_),
    .C(_1334_),
    .Y(_1367_)
);

AOI21X1 _4618_ (
    .A(_1367_),
    .B(_1356_),
    .C(_1366_),
    .Y(_1368_)
);

NOR2X1 _4619_ (
    .A(_1365_),
    .B(_1368_),
    .Y(\z2.q0 [6])
);

OAI21X1 _4620_ (
    .A(_1361_),
    .B(_1354_),
    .C(\z2.z1.z4.z2.s ),
    .Y(_1287_)
);

NAND3X1 _4621_ (
    .A(_1356_),
    .B(_1366_),
    .C(_1367_),
    .Y(_1288_)
);

NAND3X1 _4622_ (
    .A(\z2.z1.z4.z2.c ),
    .B(_1287_),
    .C(_1288_),
    .Y(_1289_)
);

INVX1 _4623_ (
    .A(\z2.z1.z4.z2.c ),
    .Y(_1290_)
);

INVX1 _4624_ (
    .A(_1287_),
    .Y(_1291_)
);

OAI21X1 _4625_ (
    .A(_1291_),
    .B(_1365_),
    .C(_1290_),
    .Y(_1292_)
);

NAND2X1 _4626_ (
    .A(_1289_),
    .B(_1292_),
    .Y(\z2.q0 [7])
);

AOI21X1 _4627_ (
    .A(_1312_),
    .B(_1309_),
    .C(_1298_),
    .Y(_1293_)
);

NOR2X1 _4628_ (
    .A(_1293_),
    .B(_1314_),
    .Y(q1[3])
);

AND2X2 _4629_ (
    .A(b[0]),
    .B(a[8]),
    .Y(q1[0])
);

AND2X2 _4630_ (
    .A(b[0]),
    .B(a[9]),
    .Y(\z2.z1.z1.z1.a )
);

AND2X2 _4631_ (
    .A(a[8]),
    .B(b[1]),
    .Y(\z2.z1.z1.z1.b )
);

AND2X2 _4632_ (
    .A(a[9]),
    .B(b[1]),
    .Y(\z2.z1.z1.z2.a )
);

INVX1 _4633_ (
    .A(\z2.z1.z1.z1.b ),
    .Y(_1369_)
);

NAND2X1 _4634_ (
    .A(\z2.z1.z1.z1.a ),
    .B(_1369_),
    .Y(_1370_)
);

INVX1 _4635_ (
    .A(\z2.z1.z1.z1.a ),
    .Y(_1371_)
);

NAND2X1 _4636_ (
    .A(\z2.z1.z1.z1.b ),
    .B(_1371_),
    .Y(_1372_)
);

NAND2X1 _4637_ (
    .A(_1370_),
    .B(_1372_),
    .Y(\z2.z1.z1.z1.s )
);

NOR2X1 _4638_ (
    .A(_1369_),
    .B(_1371_),
    .Y(\z2.z1.z1.z1.c )
);

INVX1 _4639_ (
    .A(\z2.z1.z1.z1.c ),
    .Y(_1373_)
);

NAND2X1 _4640_ (
    .A(\z2.z1.z1.z2.a ),
    .B(_1373_),
    .Y(_1374_)
);

INVX1 _4641_ (
    .A(\z2.z1.z1.z2.a ),
    .Y(_1375_)
);

NAND2X1 _4642_ (
    .A(\z2.z1.z1.z1.c ),
    .B(_1375_),
    .Y(_1376_)
);

NAND2X1 _4643_ (
    .A(_1374_),
    .B(_1376_),
    .Y(\z2.z1.z1.z2.s )
);

NOR2X1 _4644_ (
    .A(_1373_),
    .B(_1375_),
    .Y(\z2.z1.z1.z2.c )
);

AND2X2 _4645_ (
    .A(b[0]),
    .B(a[10]),
    .Y(\z2.z1.q1 [0])
);

AND2X2 _4646_ (
    .A(b[0]),
    .B(a[11]),
    .Y(\z2.z1.z2.z1.a )
);

AND2X2 _4647_ (
    .A(a[10]),
    .B(b[1]),
    .Y(\z2.z1.z2.z1.b )
);

AND2X2 _4648_ (
    .A(a[11]),
    .B(b[1]),
    .Y(\z2.z1.z2.z2.a )
);

INVX1 _4649_ (
    .A(\z2.z1.z2.z1.b ),
    .Y(_1377_)
);

NAND2X1 _4650_ (
    .A(\z2.z1.z2.z1.a ),
    .B(_1377_),
    .Y(_1378_)
);

INVX1 _4651_ (
    .A(\z2.z1.z2.z1.a ),
    .Y(_1379_)
);

NAND2X1 _4652_ (
    .A(\z2.z1.z2.z1.b ),
    .B(_1379_),
    .Y(_1380_)
);

NAND2X1 _4653_ (
    .A(_1378_),
    .B(_1380_),
    .Y(\z2.z1.z2.z1.s )
);

NOR2X1 _4654_ (
    .A(_1377_),
    .B(_1379_),
    .Y(\z2.z1.z2.z1.c )
);

INVX1 _4655_ (
    .A(\z2.z1.z2.z1.c ),
    .Y(_1381_)
);

NAND2X1 _4656_ (
    .A(\z2.z1.z2.z2.a ),
    .B(_1381_),
    .Y(_1382_)
);

INVX1 _4657_ (
    .A(\z2.z1.z2.z2.a ),
    .Y(_1383_)
);

NAND2X1 _4658_ (
    .A(\z2.z1.z2.z1.c ),
    .B(_1383_),
    .Y(_1384_)
);

NAND2X1 _4659_ (
    .A(_1382_),
    .B(_1384_),
    .Y(\z2.z1.z2.z2.s )
);

NOR2X1 _4660_ (
    .A(_1381_),
    .B(_1383_),
    .Y(\z2.z1.z2.z2.c )
);

AND2X2 _4661_ (
    .A(b[2]),
    .B(a[8]),
    .Y(\z2.z1.q2 [0])
);

AND2X2 _4662_ (
    .A(b[2]),
    .B(a[9]),
    .Y(\z2.z1.z3.z1.a )
);

AND2X2 _4663_ (
    .A(a[8]),
    .B(b[3]),
    .Y(\z2.z1.z3.z1.b )
);

AND2X2 _4664_ (
    .A(a[9]),
    .B(b[3]),
    .Y(\z2.z1.z3.z2.a )
);

INVX1 _4665_ (
    .A(\z2.z1.z3.z1.b ),
    .Y(_1385_)
);

NAND2X1 _4666_ (
    .A(\z2.z1.z3.z1.a ),
    .B(_1385_),
    .Y(_1386_)
);

INVX1 _4667_ (
    .A(\z2.z1.z3.z1.a ),
    .Y(_1387_)
);

NAND2X1 _4668_ (
    .A(\z2.z1.z3.z1.b ),
    .B(_1387_),
    .Y(_1388_)
);

NAND2X1 _4669_ (
    .A(_1386_),
    .B(_1388_),
    .Y(\z2.z1.z3.z1.s )
);

NOR2X1 _4670_ (
    .A(_1385_),
    .B(_1387_),
    .Y(\z2.z1.z3.z1.c )
);

INVX1 _4671_ (
    .A(\z2.z1.z3.z1.c ),
    .Y(_1389_)
);

NAND2X1 _4672_ (
    .A(\z2.z1.z3.z2.a ),
    .B(_1389_),
    .Y(_1390_)
);

INVX1 _4673_ (
    .A(\z2.z1.z3.z2.a ),
    .Y(_1391_)
);

NAND2X1 _4674_ (
    .A(\z2.z1.z3.z1.c ),
    .B(_1391_),
    .Y(_1392_)
);

NAND2X1 _4675_ (
    .A(_1390_),
    .B(_1392_),
    .Y(\z2.z1.z3.z2.s )
);

NOR2X1 _4676_ (
    .A(_1389_),
    .B(_1391_),
    .Y(\z2.z1.z3.z2.c )
);

AND2X2 _4677_ (
    .A(b[2]),
    .B(a[10]),
    .Y(\z2.z1.q3 [0])
);

AND2X2 _4678_ (
    .A(b[2]),
    .B(a[11]),
    .Y(\z2.z1.z4.z1.a )
);

AND2X2 _4679_ (
    .A(a[10]),
    .B(b[3]),
    .Y(\z2.z1.z4.z1.b )
);

AND2X2 _4680_ (
    .A(a[11]),
    .B(b[3]),
    .Y(\z2.z1.z4.z2.a )
);

INVX1 _4681_ (
    .A(\z2.z1.z4.z1.b ),
    .Y(_1393_)
);

NAND2X1 _4682_ (
    .A(\z2.z1.z4.z1.a ),
    .B(_1393_),
    .Y(_1394_)
);

INVX1 _4683_ (
    .A(\z2.z1.z4.z1.a ),
    .Y(_1395_)
);

NAND2X1 _4684_ (
    .A(\z2.z1.z4.z1.b ),
    .B(_1395_),
    .Y(_1396_)
);

NAND2X1 _4685_ (
    .A(_1394_),
    .B(_1396_),
    .Y(\z2.z1.z4.z1.s )
);

NOR2X1 _4686_ (
    .A(_1393_),
    .B(_1395_),
    .Y(\z2.z1.z4.z1.c )
);

INVX1 _4687_ (
    .A(\z2.z1.z4.z1.c ),
    .Y(_1397_)
);

NAND2X1 _4688_ (
    .A(\z2.z1.z4.z2.a ),
    .B(_1397_),
    .Y(_1398_)
);

INVX1 _4689_ (
    .A(\z2.z1.z4.z2.a ),
    .Y(_1399_)
);

NAND2X1 _4690_ (
    .A(\z2.z1.z4.z1.c ),
    .B(_1399_),
    .Y(_1400_)
);

NAND2X1 _4691_ (
    .A(_1398_),
    .B(_1400_),
    .Y(\z2.z1.z4.z2.s )
);

NOR2X1 _4692_ (
    .A(_1397_),
    .B(_1399_),
    .Y(\z2.z1.z4.z2.c )
);

NOR2X1 _4693_ (
    .A(\z2.z2.q1 [0]),
    .B(\z2.z2.z1.z2.s ),
    .Y(_1408_)
);

AND2X2 _4694_ (
    .A(\z2.z2.q1 [0]),
    .B(\z2.z2.z1.z2.s ),
    .Y(_1409_)
);

NOR2X1 _4695_ (
    .A(_1408_),
    .B(_1409_),
    .Y(_1410_)
);

NAND2X1 _4696_ (
    .A(\z2.z2.q2 [0]),
    .B(_1410_),
    .Y(_1411_)
);

INVX1 _4697_ (
    .A(_1411_),
    .Y(_1412_)
);

NOR2X1 _4698_ (
    .A(\z2.z2.q2 [0]),
    .B(_1410_),
    .Y(_1413_)
);

NOR2X1 _4699_ (
    .A(_1413_),
    .B(_1412_),
    .Y(\z2.q1 [2])
);

NAND2X1 _4700_ (
    .A(\z2.z2.q1 [0]),
    .B(\z2.z2.z1.z2.s ),
    .Y(_1414_)
);

NOR2X1 _4701_ (
    .A(\z2.z2.z2.z1.s ),
    .B(\z2.z2.z1.z2.c ),
    .Y(_1415_)
);

NAND2X1 _4702_ (
    .A(\z2.z2.z2.z1.s ),
    .B(\z2.z2.z1.z2.c ),
    .Y(_1416_)
);

INVX1 _4703_ (
    .A(_1416_),
    .Y(_1417_)
);

OAI21X1 _4704_ (
    .A(_1415_),
    .B(_1417_),
    .C(_1414_),
    .Y(_1418_)
);

INVX1 _4705_ (
    .A(\z2.z2.z2.z1.s ),
    .Y(_1419_)
);

INVX1 _4706_ (
    .A(\z2.z2.z1.z2.c ),
    .Y(_1420_)
);

NAND2X1 _4707_ (
    .A(_1419_),
    .B(_1420_),
    .Y(_1421_)
);

NAND3X1 _4708_ (
    .A(_1409_),
    .B(_1416_),
    .C(_1421_),
    .Y(_1422_)
);

NAND3X1 _4709_ (
    .A(\z2.z2.z3.z1.s ),
    .B(_1422_),
    .C(_1418_),
    .Y(_1423_)
);

INVX1 _4710_ (
    .A(\z2.z2.z3.z1.s ),
    .Y(_1424_)
);

NAND2X1 _4711_ (
    .A(_1422_),
    .B(_1418_),
    .Y(_1425_)
);

NAND2X1 _4712_ (
    .A(_1424_),
    .B(_1425_),
    .Y(_1426_)
);

NAND3X1 _4713_ (
    .A(_1412_),
    .B(_1423_),
    .C(_1426_),
    .Y(_1427_)
);

INVX1 _4714_ (
    .A(_1427_),
    .Y(_1428_)
);

INVX1 _4715_ (
    .A(_1423_),
    .Y(_1429_)
);

OAI21X1 _4716_ (
    .A(_1414_),
    .B(_1415_),
    .C(_1416_),
    .Y(_1430_)
);

NAND2X1 _4717_ (
    .A(\z2.z2.z2.z2.s ),
    .B(_1430_),
    .Y(_1431_)
);

INVX1 _4718_ (
    .A(\z2.z2.z2.z2.s ),
    .Y(_1432_)
);

NAND3X1 _4719_ (
    .A(_1432_),
    .B(_1416_),
    .C(_1422_),
    .Y(_1433_)
);

NAND2X1 _4720_ (
    .A(\z2.z2.q3 [0]),
    .B(\z2.z2.z3.z2.s ),
    .Y(_1434_)
);

INVX1 _4721_ (
    .A(\z2.z2.q3 [0]),
    .Y(_1435_)
);

INVX1 _4722_ (
    .A(\z2.z2.z3.z2.s ),
    .Y(_1436_)
);

NAND2X1 _4723_ (
    .A(_1435_),
    .B(_1436_),
    .Y(_1437_)
);

NAND2X1 _4724_ (
    .A(_1434_),
    .B(_1437_),
    .Y(_1438_)
);

INVX1 _4725_ (
    .A(_1438_),
    .Y(_1439_)
);

NAND3X1 _4726_ (
    .A(_1431_),
    .B(_1439_),
    .C(_1433_),
    .Y(_1440_)
);

AND2X2 _4727_ (
    .A(_1430_),
    .B(\z2.z2.z2.z2.s ),
    .Y(_1441_)
);

NOR2X1 _4728_ (
    .A(\z2.z2.z2.z2.s ),
    .B(_1430_),
    .Y(_1442_)
);

OAI21X1 _4729_ (
    .A(_1442_),
    .B(_1441_),
    .C(_1438_),
    .Y(_1443_)
);

NAND3X1 _4730_ (
    .A(_1429_),
    .B(_1440_),
    .C(_1443_),
    .Y(_1444_)
);

INVX1 _4731_ (
    .A(_1440_),
    .Y(_1445_)
);

AOI21X1 _4732_ (
    .A(_1433_),
    .B(_1431_),
    .C(_1439_),
    .Y(_1446_)
);

OAI21X1 _4733_ (
    .A(_1446_),
    .B(_1445_),
    .C(_1423_),
    .Y(_1447_)
);

NAND3X1 _4734_ (
    .A(_1428_),
    .B(_1444_),
    .C(_1447_),
    .Y(_1448_)
);

INVX1 _4735_ (
    .A(_1444_),
    .Y(_1449_)
);

INVX1 _4736_ (
    .A(_1425_),
    .Y(_1450_)
);

AOI22X1 _4737_ (
    .A(\z2.z2.z3.z1.s ),
    .B(_1450_),
    .C(_1443_),
    .D(_1440_),
    .Y(_1451_)
);

OAI21X1 _4738_ (
    .A(_1451_),
    .B(_1449_),
    .C(_1427_),
    .Y(_1452_)
);

AND2X2 _4739_ (
    .A(_1452_),
    .B(_1448_),
    .Y(\z2.q1 [4])
);

OAI21X1 _4740_ (
    .A(_1427_),
    .B(_1451_),
    .C(_1444_),
    .Y(_1453_)
);

OAI21X1 _4741_ (
    .A(_1435_),
    .B(_1436_),
    .C(_1440_),
    .Y(_1454_)
);

NAND2X1 _4742_ (
    .A(\z2.z2.z4.z1.s ),
    .B(\z2.z2.z3.z2.c ),
    .Y(_1455_)
);

OR2X2 _4743_ (
    .A(\z2.z2.z4.z1.s ),
    .B(\z2.z2.z3.z2.c ),
    .Y(_1456_)
);

NAND2X1 _4744_ (
    .A(_1455_),
    .B(_1456_),
    .Y(_1457_)
);

INVX1 _4745_ (
    .A(_1457_),
    .Y(_1458_)
);

NAND2X1 _4746_ (
    .A(\z2.z2.z2.z2.c ),
    .B(_1441_),
    .Y(_1459_)
);

INVX1 _4747_ (
    .A(\z2.z2.z2.z2.c ),
    .Y(_1460_)
);

NAND2X1 _4748_ (
    .A(_1460_),
    .B(_1431_),
    .Y(_1461_)
);

NAND3X1 _4749_ (
    .A(_1458_),
    .B(_1461_),
    .C(_1459_),
    .Y(_1462_)
);

NAND2X1 _4750_ (
    .A(\z2.z2.z2.z2.c ),
    .B(_1431_),
    .Y(_1463_)
);

NAND2X1 _4751_ (
    .A(_1460_),
    .B(_1441_),
    .Y(_1464_)
);

NAND3X1 _4752_ (
    .A(_1457_),
    .B(_1463_),
    .C(_1464_),
    .Y(_1465_)
);

NAND3X1 _4753_ (
    .A(_1454_),
    .B(_1462_),
    .C(_1465_),
    .Y(_1466_)
);

INVX1 _4754_ (
    .A(_1454_),
    .Y(_1467_)
);

AOI21X1 _4755_ (
    .A(_1464_),
    .B(_1463_),
    .C(_1457_),
    .Y(_1468_)
);

AOI21X1 _4756_ (
    .A(_1459_),
    .B(_1461_),
    .C(_1458_),
    .Y(_1469_)
);

OAI21X1 _4757_ (
    .A(_1468_),
    .B(_1469_),
    .C(_1467_),
    .Y(_1470_)
);

NAND2X1 _4758_ (
    .A(_1466_),
    .B(_1470_),
    .Y(_1471_)
);

NAND2X1 _4759_ (
    .A(_1453_),
    .B(_1471_),
    .Y(_1472_)
);

OR2X2 _4760_ (
    .A(_1471_),
    .B(_1453_),
    .Y(_1473_)
);

NAND2X1 _4761_ (
    .A(_1472_),
    .B(_1473_),
    .Y(\z2.q1 [5])
);

INVX1 _4762_ (
    .A(\z2.z2.z4.z2.s ),
    .Y(_1474_)
);

INVX1 _4763_ (
    .A(_1455_),
    .Y(_1475_)
);

OAI21X1 _4764_ (
    .A(_1475_),
    .B(_1468_),
    .C(_1474_),
    .Y(_1476_)
);

NAND3X1 _4765_ (
    .A(\z2.z2.z4.z2.s ),
    .B(_1455_),
    .C(_1462_),
    .Y(_1477_)
);

NAND2X1 _4766_ (
    .A(_1470_),
    .B(_1453_),
    .Y(_1478_)
);

AOI22X1 _4767_ (
    .A(_1476_),
    .B(_1477_),
    .C(_1478_),
    .D(_1466_),
    .Y(_1479_)
);

NAND2X1 _4768_ (
    .A(_1477_),
    .B(_1476_),
    .Y(_1480_)
);

NAND3X1 _4769_ (
    .A(_1444_),
    .B(_1466_),
    .C(_1448_),
    .Y(_1481_)
);

AOI21X1 _4770_ (
    .A(_1481_),
    .B(_1470_),
    .C(_1480_),
    .Y(_1482_)
);

NOR2X1 _4771_ (
    .A(_1479_),
    .B(_1482_),
    .Y(\z2.q1 [6])
);

OAI21X1 _4772_ (
    .A(_1475_),
    .B(_1468_),
    .C(\z2.z2.z4.z2.s ),
    .Y(_1401_)
);

NAND3X1 _4773_ (
    .A(_1470_),
    .B(_1480_),
    .C(_1481_),
    .Y(_1402_)
);

NAND3X1 _4774_ (
    .A(\z2.z2.z4.z2.c ),
    .B(_1401_),
    .C(_1402_),
    .Y(_1403_)
);

INVX1 _4775_ (
    .A(\z2.z2.z4.z2.c ),
    .Y(_1404_)
);

INVX1 _4776_ (
    .A(_1401_),
    .Y(_1405_)
);

OAI21X1 _4777_ (
    .A(_1405_),
    .B(_1479_),
    .C(_1404_),
    .Y(_1406_)
);

NAND2X1 _4778_ (
    .A(_1403_),
    .B(_1406_),
    .Y(\z2.q1 [7])
);

AOI21X1 _4779_ (
    .A(_1426_),
    .B(_1423_),
    .C(_1412_),
    .Y(_1407_)
);

NOR2X1 _4780_ (
    .A(_1407_),
    .B(_1428_),
    .Y(\z2.q1 [3])
);

AND2X2 _4781_ (
    .A(b[0]),
    .B(a[12]),
    .Y(\z2.q1 [0])
);

AND2X2 _4782_ (
    .A(b[0]),
    .B(a[13]),
    .Y(\z2.z2.z1.z1.a )
);

AND2X2 _4783_ (
    .A(a[12]),
    .B(b[1]),
    .Y(\z2.z2.z1.z1.b )
);

AND2X2 _4784_ (
    .A(a[13]),
    .B(b[1]),
    .Y(\z2.z2.z1.z2.a )
);

INVX1 _4785_ (
    .A(\z2.z2.z1.z1.b ),
    .Y(_1483_)
);

NAND2X1 _4786_ (
    .A(\z2.z2.z1.z1.a ),
    .B(_1483_),
    .Y(_1484_)
);

INVX1 _4787_ (
    .A(\z2.z2.z1.z1.a ),
    .Y(_1485_)
);

NAND2X1 _4788_ (
    .A(\z2.z2.z1.z1.b ),
    .B(_1485_),
    .Y(_1486_)
);

NAND2X1 _4789_ (
    .A(_1484_),
    .B(_1486_),
    .Y(\z2.z2.z1.z1.s )
);

NOR2X1 _4790_ (
    .A(_1483_),
    .B(_1485_),
    .Y(\z2.z2.z1.z1.c )
);

INVX1 _4791_ (
    .A(\z2.z2.z1.z1.c ),
    .Y(_1487_)
);

NAND2X1 _4792_ (
    .A(\z2.z2.z1.z2.a ),
    .B(_1487_),
    .Y(_1488_)
);

INVX1 _4793_ (
    .A(\z2.z2.z1.z2.a ),
    .Y(_1489_)
);

NAND2X1 _4794_ (
    .A(\z2.z2.z1.z1.c ),
    .B(_1489_),
    .Y(_1490_)
);

NAND2X1 _4795_ (
    .A(_1488_),
    .B(_1490_),
    .Y(\z2.z2.z1.z2.s )
);

NOR2X1 _4796_ (
    .A(_1487_),
    .B(_1489_),
    .Y(\z2.z2.z1.z2.c )
);

AND2X2 _4797_ (
    .A(b[0]),
    .B(a[14]),
    .Y(\z2.z2.q1 [0])
);

AND2X2 _4798_ (
    .A(b[0]),
    .B(a[15]),
    .Y(\z2.z2.z2.z1.a )
);

AND2X2 _4799_ (
    .A(a[14]),
    .B(b[1]),
    .Y(\z2.z2.z2.z1.b )
);

AND2X2 _4800_ (
    .A(a[15]),
    .B(b[1]),
    .Y(\z2.z2.z2.z2.a )
);

INVX1 _4801_ (
    .A(\z2.z2.z2.z1.b ),
    .Y(_1491_)
);

NAND2X1 _4802_ (
    .A(\z2.z2.z2.z1.a ),
    .B(_1491_),
    .Y(_1492_)
);

INVX1 _4803_ (
    .A(\z2.z2.z2.z1.a ),
    .Y(_1493_)
);

NAND2X1 _4804_ (
    .A(\z2.z2.z2.z1.b ),
    .B(_1493_),
    .Y(_1494_)
);

NAND2X1 _4805_ (
    .A(_1492_),
    .B(_1494_),
    .Y(\z2.z2.z2.z1.s )
);

NOR2X1 _4806_ (
    .A(_1491_),
    .B(_1493_),
    .Y(\z2.z2.z2.z1.c )
);

INVX1 _4807_ (
    .A(\z2.z2.z2.z1.c ),
    .Y(_1495_)
);

NAND2X1 _4808_ (
    .A(\z2.z2.z2.z2.a ),
    .B(_1495_),
    .Y(_1496_)
);

INVX1 _4809_ (
    .A(\z2.z2.z2.z2.a ),
    .Y(_1497_)
);

NAND2X1 _4810_ (
    .A(\z2.z2.z2.z1.c ),
    .B(_1497_),
    .Y(_1498_)
);

NAND2X1 _4811_ (
    .A(_1496_),
    .B(_1498_),
    .Y(\z2.z2.z2.z2.s )
);

NOR2X1 _4812_ (
    .A(_1495_),
    .B(_1497_),
    .Y(\z2.z2.z2.z2.c )
);

AND2X2 _4813_ (
    .A(b[2]),
    .B(a[12]),
    .Y(\z2.z2.q2 [0])
);

AND2X2 _4814_ (
    .A(b[2]),
    .B(a[13]),
    .Y(\z2.z2.z3.z1.a )
);

AND2X2 _4815_ (
    .A(a[12]),
    .B(b[3]),
    .Y(\z2.z2.z3.z1.b )
);

AND2X2 _4816_ (
    .A(a[13]),
    .B(b[3]),
    .Y(\z2.z2.z3.z2.a )
);

INVX1 _4817_ (
    .A(\z2.z2.z3.z1.b ),
    .Y(_1499_)
);

NAND2X1 _4818_ (
    .A(\z2.z2.z3.z1.a ),
    .B(_1499_),
    .Y(_1500_)
);

INVX1 _4819_ (
    .A(\z2.z2.z3.z1.a ),
    .Y(_1501_)
);

NAND2X1 _4820_ (
    .A(\z2.z2.z3.z1.b ),
    .B(_1501_),
    .Y(_1502_)
);

NAND2X1 _4821_ (
    .A(_1500_),
    .B(_1502_),
    .Y(\z2.z2.z3.z1.s )
);

NOR2X1 _4822_ (
    .A(_1499_),
    .B(_1501_),
    .Y(\z2.z2.z3.z1.c )
);

INVX1 _4823_ (
    .A(\z2.z2.z3.z1.c ),
    .Y(_1503_)
);

NAND2X1 _4824_ (
    .A(\z2.z2.z3.z2.a ),
    .B(_1503_),
    .Y(_1504_)
);

INVX1 _4825_ (
    .A(\z2.z2.z3.z2.a ),
    .Y(_1505_)
);

NAND2X1 _4826_ (
    .A(\z2.z2.z3.z1.c ),
    .B(_1505_),
    .Y(_1506_)
);

NAND2X1 _4827_ (
    .A(_1504_),
    .B(_1506_),
    .Y(\z2.z2.z3.z2.s )
);

NOR2X1 _4828_ (
    .A(_1503_),
    .B(_1505_),
    .Y(\z2.z2.z3.z2.c )
);

AND2X2 _4829_ (
    .A(b[2]),
    .B(a[14]),
    .Y(\z2.z2.q3 [0])
);

AND2X2 _4830_ (
    .A(b[2]),
    .B(a[15]),
    .Y(\z2.z2.z4.z1.a )
);

AND2X2 _4831_ (
    .A(a[14]),
    .B(b[3]),
    .Y(\z2.z2.z4.z1.b )
);

AND2X2 _4832_ (
    .A(a[15]),
    .B(b[3]),
    .Y(\z2.z2.z4.z2.a )
);

INVX1 _4833_ (
    .A(\z2.z2.z4.z1.b ),
    .Y(_1507_)
);

NAND2X1 _4834_ (
    .A(\z2.z2.z4.z1.a ),
    .B(_1507_),
    .Y(_1508_)
);

INVX1 _4835_ (
    .A(\z2.z2.z4.z1.a ),
    .Y(_1509_)
);

NAND2X1 _4836_ (
    .A(\z2.z2.z4.z1.b ),
    .B(_1509_),
    .Y(_1510_)
);

NAND2X1 _4837_ (
    .A(_1508_),
    .B(_1510_),
    .Y(\z2.z2.z4.z1.s )
);

NOR2X1 _4838_ (
    .A(_1507_),
    .B(_1509_),
    .Y(\z2.z2.z4.z1.c )
);

INVX1 _4839_ (
    .A(\z2.z2.z4.z1.c ),
    .Y(_1511_)
);

NAND2X1 _4840_ (
    .A(\z2.z2.z4.z2.a ),
    .B(_1511_),
    .Y(_1512_)
);

INVX1 _4841_ (
    .A(\z2.z2.z4.z2.a ),
    .Y(_1513_)
);

NAND2X1 _4842_ (
    .A(\z2.z2.z4.z1.c ),
    .B(_1513_),
    .Y(_1514_)
);

NAND2X1 _4843_ (
    .A(_1512_),
    .B(_1514_),
    .Y(\z2.z2.z4.z2.s )
);

NOR2X1 _4844_ (
    .A(_1511_),
    .B(_1513_),
    .Y(\z2.z2.z4.z2.c )
);

NOR2X1 _4845_ (
    .A(\z2.z3.q1 [0]),
    .B(\z2.z3.z1.z2.s ),
    .Y(_1522_)
);

AND2X2 _4846_ (
    .A(\z2.z3.q1 [0]),
    .B(\z2.z3.z1.z2.s ),
    .Y(_1523_)
);

NOR2X1 _4847_ (
    .A(_1522_),
    .B(_1523_),
    .Y(_1524_)
);

NAND2X1 _4848_ (
    .A(\z2.z3.q2 [0]),
    .B(_1524_),
    .Y(_1525_)
);

INVX1 _4849_ (
    .A(_1525_),
    .Y(_1526_)
);

NOR2X1 _4850_ (
    .A(\z2.z3.q2 [0]),
    .B(_1524_),
    .Y(_1527_)
);

NOR2X1 _4851_ (
    .A(_1527_),
    .B(_1526_),
    .Y(\z2.q2 [2])
);

NAND2X1 _4852_ (
    .A(\z2.z3.q1 [0]),
    .B(\z2.z3.z1.z2.s ),
    .Y(_1528_)
);

NOR2X1 _4853_ (
    .A(\z2.z3.z2.z1.s ),
    .B(\z2.z3.z1.z2.c ),
    .Y(_1529_)
);

NAND2X1 _4854_ (
    .A(\z2.z3.z2.z1.s ),
    .B(\z2.z3.z1.z2.c ),
    .Y(_1530_)
);

INVX1 _4855_ (
    .A(_1530_),
    .Y(_1531_)
);

OAI21X1 _4856_ (
    .A(_1529_),
    .B(_1531_),
    .C(_1528_),
    .Y(_1532_)
);

INVX1 _4857_ (
    .A(\z2.z3.z2.z1.s ),
    .Y(_1533_)
);

INVX1 _4858_ (
    .A(\z2.z3.z1.z2.c ),
    .Y(_1534_)
);

NAND2X1 _4859_ (
    .A(_1533_),
    .B(_1534_),
    .Y(_1535_)
);

NAND3X1 _4860_ (
    .A(_1523_),
    .B(_1530_),
    .C(_1535_),
    .Y(_1536_)
);

NAND3X1 _4861_ (
    .A(\z2.z3.z3.z1.s ),
    .B(_1536_),
    .C(_1532_),
    .Y(_1537_)
);

INVX1 _4862_ (
    .A(\z2.z3.z3.z1.s ),
    .Y(_1538_)
);

NAND2X1 _4863_ (
    .A(_1536_),
    .B(_1532_),
    .Y(_1539_)
);

NAND2X1 _4864_ (
    .A(_1538_),
    .B(_1539_),
    .Y(_1540_)
);

NAND3X1 _4865_ (
    .A(_1526_),
    .B(_1537_),
    .C(_1540_),
    .Y(_1541_)
);

INVX1 _4866_ (
    .A(_1541_),
    .Y(_1542_)
);

INVX1 _4867_ (
    .A(_1537_),
    .Y(_1543_)
);

OAI21X1 _4868_ (
    .A(_1528_),
    .B(_1529_),
    .C(_1530_),
    .Y(_1544_)
);

NAND2X1 _4869_ (
    .A(\z2.z3.z2.z2.s ),
    .B(_1544_),
    .Y(_1545_)
);

INVX1 _4870_ (
    .A(\z2.z3.z2.z2.s ),
    .Y(_1546_)
);

NAND3X1 _4871_ (
    .A(_1546_),
    .B(_1530_),
    .C(_1536_),
    .Y(_1547_)
);

NAND2X1 _4872_ (
    .A(\z2.z3.q3 [0]),
    .B(\z2.z3.z3.z2.s ),
    .Y(_1548_)
);

INVX1 _4873_ (
    .A(\z2.z3.q3 [0]),
    .Y(_1549_)
);

INVX1 _4874_ (
    .A(\z2.z3.z3.z2.s ),
    .Y(_1550_)
);

NAND2X1 _4875_ (
    .A(_1549_),
    .B(_1550_),
    .Y(_1551_)
);

NAND2X1 _4876_ (
    .A(_1548_),
    .B(_1551_),
    .Y(_1552_)
);

INVX1 _4877_ (
    .A(_1552_),
    .Y(_1553_)
);

NAND3X1 _4878_ (
    .A(_1545_),
    .B(_1553_),
    .C(_1547_),
    .Y(_1554_)
);

AND2X2 _4879_ (
    .A(_1544_),
    .B(\z2.z3.z2.z2.s ),
    .Y(_1555_)
);

NOR2X1 _4880_ (
    .A(\z2.z3.z2.z2.s ),
    .B(_1544_),
    .Y(_1556_)
);

OAI21X1 _4881_ (
    .A(_1556_),
    .B(_1555_),
    .C(_1552_),
    .Y(_1557_)
);

NAND3X1 _4882_ (
    .A(_1543_),
    .B(_1554_),
    .C(_1557_),
    .Y(_1558_)
);

INVX1 _4883_ (
    .A(_1554_),
    .Y(_1559_)
);

AOI21X1 _4884_ (
    .A(_1547_),
    .B(_1545_),
    .C(_1553_),
    .Y(_1560_)
);

OAI21X1 _4885_ (
    .A(_1560_),
    .B(_1559_),
    .C(_1537_),
    .Y(_1561_)
);

NAND3X1 _4886_ (
    .A(_1542_),
    .B(_1558_),
    .C(_1561_),
    .Y(_1562_)
);

INVX1 _4887_ (
    .A(_1558_),
    .Y(_1563_)
);

INVX1 _4888_ (
    .A(_1539_),
    .Y(_1564_)
);

AOI22X1 _4889_ (
    .A(\z2.z3.z3.z1.s ),
    .B(_1564_),
    .C(_1557_),
    .D(_1554_),
    .Y(_1565_)
);

OAI21X1 _4890_ (
    .A(_1565_),
    .B(_1563_),
    .C(_1541_),
    .Y(_1566_)
);

AND2X2 _4891_ (
    .A(_1566_),
    .B(_1562_),
    .Y(\z2.q2 [4])
);

OAI21X1 _4892_ (
    .A(_1541_),
    .B(_1565_),
    .C(_1558_),
    .Y(_1567_)
);

OAI21X1 _4893_ (
    .A(_1549_),
    .B(_1550_),
    .C(_1554_),
    .Y(_1568_)
);

NAND2X1 _4894_ (
    .A(\z2.z3.z4.z1.s ),
    .B(\z2.z3.z3.z2.c ),
    .Y(_1569_)
);

OR2X2 _4895_ (
    .A(\z2.z3.z4.z1.s ),
    .B(\z2.z3.z3.z2.c ),
    .Y(_1570_)
);

NAND2X1 _4896_ (
    .A(_1569_),
    .B(_1570_),
    .Y(_1571_)
);

INVX1 _4897_ (
    .A(_1571_),
    .Y(_1572_)
);

NAND2X1 _4898_ (
    .A(\z2.z3.z2.z2.c ),
    .B(_1555_),
    .Y(_1573_)
);

INVX1 _4899_ (
    .A(\z2.z3.z2.z2.c ),
    .Y(_1574_)
);

NAND2X1 _4900_ (
    .A(_1574_),
    .B(_1545_),
    .Y(_1575_)
);

NAND3X1 _4901_ (
    .A(_1572_),
    .B(_1575_),
    .C(_1573_),
    .Y(_1576_)
);

NAND2X1 _4902_ (
    .A(\z2.z3.z2.z2.c ),
    .B(_1545_),
    .Y(_1577_)
);

NAND2X1 _4903_ (
    .A(_1574_),
    .B(_1555_),
    .Y(_1578_)
);

NAND3X1 _4904_ (
    .A(_1571_),
    .B(_1577_),
    .C(_1578_),
    .Y(_1579_)
);

NAND3X1 _4905_ (
    .A(_1568_),
    .B(_1576_),
    .C(_1579_),
    .Y(_1580_)
);

INVX1 _4906_ (
    .A(_1568_),
    .Y(_1581_)
);

AOI21X1 _4907_ (
    .A(_1578_),
    .B(_1577_),
    .C(_1571_),
    .Y(_1582_)
);

AOI21X1 _4908_ (
    .A(_1573_),
    .B(_1575_),
    .C(_1572_),
    .Y(_1583_)
);

OAI21X1 _4909_ (
    .A(_1582_),
    .B(_1583_),
    .C(_1581_),
    .Y(_1584_)
);

NAND2X1 _4910_ (
    .A(_1580_),
    .B(_1584_),
    .Y(_1585_)
);

NAND2X1 _4911_ (
    .A(_1567_),
    .B(_1585_),
    .Y(_1586_)
);

OR2X2 _4912_ (
    .A(_1585_),
    .B(_1567_),
    .Y(_1587_)
);

NAND2X1 _4913_ (
    .A(_1586_),
    .B(_1587_),
    .Y(\z2.q2 [5])
);

INVX1 _4914_ (
    .A(\z2.z3.z4.z2.s ),
    .Y(_1588_)
);

INVX1 _4915_ (
    .A(_1569_),
    .Y(_1589_)
);

OAI21X1 _4916_ (
    .A(_1589_),
    .B(_1582_),
    .C(_1588_),
    .Y(_1590_)
);

NAND3X1 _4917_ (
    .A(\z2.z3.z4.z2.s ),
    .B(_1569_),
    .C(_1576_),
    .Y(_1591_)
);

NAND2X1 _4918_ (
    .A(_1584_),
    .B(_1567_),
    .Y(_1592_)
);

AOI22X1 _4919_ (
    .A(_1590_),
    .B(_1591_),
    .C(_1592_),
    .D(_1580_),
    .Y(_1593_)
);

NAND2X1 _4920_ (
    .A(_1591_),
    .B(_1590_),
    .Y(_1594_)
);

NAND3X1 _4921_ (
    .A(_1558_),
    .B(_1580_),
    .C(_1562_),
    .Y(_1595_)
);

AOI21X1 _4922_ (
    .A(_1595_),
    .B(_1584_),
    .C(_1594_),
    .Y(_1596_)
);

NOR2X1 _4923_ (
    .A(_1593_),
    .B(_1596_),
    .Y(\z2.q2 [6])
);

OAI21X1 _4924_ (
    .A(_1589_),
    .B(_1582_),
    .C(\z2.z3.z4.z2.s ),
    .Y(_1515_)
);

NAND3X1 _4925_ (
    .A(_1584_),
    .B(_1594_),
    .C(_1595_),
    .Y(_1516_)
);

NAND3X1 _4926_ (
    .A(\z2.z3.z4.z2.c ),
    .B(_1515_),
    .C(_1516_),
    .Y(_1517_)
);

INVX1 _4927_ (
    .A(\z2.z3.z4.z2.c ),
    .Y(_1518_)
);

INVX1 _4928_ (
    .A(_1515_),
    .Y(_1519_)
);

OAI21X1 _4929_ (
    .A(_1519_),
    .B(_1593_),
    .C(_1518_),
    .Y(_1520_)
);

NAND2X1 _4930_ (
    .A(_1517_),
    .B(_1520_),
    .Y(\z2.q2 [7])
);

AOI21X1 _4931_ (
    .A(_1540_),
    .B(_1537_),
    .C(_1526_),
    .Y(_1521_)
);

NOR2X1 _4932_ (
    .A(_1521_),
    .B(_1542_),
    .Y(\z2.q2 [3])
);

AND2X2 _4933_ (
    .A(b[4]),
    .B(a[8]),
    .Y(\z2.q2 [0])
);

AND2X2 _4934_ (
    .A(b[4]),
    .B(a[9]),
    .Y(\z2.z3.z1.z1.a )
);

AND2X2 _4935_ (
    .A(a[8]),
    .B(b[5]),
    .Y(\z2.z3.z1.z1.b )
);

AND2X2 _4936_ (
    .A(a[9]),
    .B(b[5]),
    .Y(\z2.z3.z1.z2.a )
);

INVX1 _4937_ (
    .A(\z2.z3.z1.z1.b ),
    .Y(_1597_)
);

NAND2X1 _4938_ (
    .A(\z2.z3.z1.z1.a ),
    .B(_1597_),
    .Y(_1598_)
);

INVX1 _4939_ (
    .A(\z2.z3.z1.z1.a ),
    .Y(_1599_)
);

NAND2X1 _4940_ (
    .A(\z2.z3.z1.z1.b ),
    .B(_1599_),
    .Y(_1600_)
);

NAND2X1 _4941_ (
    .A(_1598_),
    .B(_1600_),
    .Y(\z2.z3.z1.z1.s )
);

NOR2X1 _4942_ (
    .A(_1597_),
    .B(_1599_),
    .Y(\z2.z3.z1.z1.c )
);

INVX1 _4943_ (
    .A(\z2.z3.z1.z1.c ),
    .Y(_1601_)
);

NAND2X1 _4944_ (
    .A(\z2.z3.z1.z2.a ),
    .B(_1601_),
    .Y(_1602_)
);

INVX1 _4945_ (
    .A(\z2.z3.z1.z2.a ),
    .Y(_1603_)
);

NAND2X1 _4946_ (
    .A(\z2.z3.z1.z1.c ),
    .B(_1603_),
    .Y(_1604_)
);

NAND2X1 _4947_ (
    .A(_1602_),
    .B(_1604_),
    .Y(\z2.z3.z1.z2.s )
);

NOR2X1 _4948_ (
    .A(_1601_),
    .B(_1603_),
    .Y(\z2.z3.z1.z2.c )
);

AND2X2 _4949_ (
    .A(b[4]),
    .B(a[10]),
    .Y(\z2.z3.q1 [0])
);

AND2X2 _4950_ (
    .A(b[4]),
    .B(a[11]),
    .Y(\z2.z3.z2.z1.a )
);

AND2X2 _4951_ (
    .A(a[10]),
    .B(b[5]),
    .Y(\z2.z3.z2.z1.b )
);

AND2X2 _4952_ (
    .A(a[11]),
    .B(b[5]),
    .Y(\z2.z3.z2.z2.a )
);

INVX1 _4953_ (
    .A(\z2.z3.z2.z1.b ),
    .Y(_1605_)
);

NAND2X1 _4954_ (
    .A(\z2.z3.z2.z1.a ),
    .B(_1605_),
    .Y(_1606_)
);

INVX1 _4955_ (
    .A(\z2.z3.z2.z1.a ),
    .Y(_1607_)
);

NAND2X1 _4956_ (
    .A(\z2.z3.z2.z1.b ),
    .B(_1607_),
    .Y(_1608_)
);

NAND2X1 _4957_ (
    .A(_1606_),
    .B(_1608_),
    .Y(\z2.z3.z2.z1.s )
);

NOR2X1 _4958_ (
    .A(_1605_),
    .B(_1607_),
    .Y(\z2.z3.z2.z1.c )
);

INVX1 _4959_ (
    .A(\z2.z3.z2.z1.c ),
    .Y(_1609_)
);

NAND2X1 _4960_ (
    .A(\z2.z3.z2.z2.a ),
    .B(_1609_),
    .Y(_1610_)
);

INVX1 _4961_ (
    .A(\z2.z3.z2.z2.a ),
    .Y(_1611_)
);

NAND2X1 _4962_ (
    .A(\z2.z3.z2.z1.c ),
    .B(_1611_),
    .Y(_1612_)
);

NAND2X1 _4963_ (
    .A(_1610_),
    .B(_1612_),
    .Y(\z2.z3.z2.z2.s )
);

NOR2X1 _4964_ (
    .A(_1609_),
    .B(_1611_),
    .Y(\z2.z3.z2.z2.c )
);

AND2X2 _4965_ (
    .A(b[6]),
    .B(a[8]),
    .Y(\z2.z3.q2 [0])
);

AND2X2 _4966_ (
    .A(b[6]),
    .B(a[9]),
    .Y(\z2.z3.z3.z1.a )
);

AND2X2 _4967_ (
    .A(a[8]),
    .B(b[7]),
    .Y(\z2.z3.z3.z1.b )
);

AND2X2 _4968_ (
    .A(a[9]),
    .B(b[7]),
    .Y(\z2.z3.z3.z2.a )
);

INVX1 _4969_ (
    .A(\z2.z3.z3.z1.b ),
    .Y(_1613_)
);

NAND2X1 _4970_ (
    .A(\z2.z3.z3.z1.a ),
    .B(_1613_),
    .Y(_1614_)
);

INVX1 _4971_ (
    .A(\z2.z3.z3.z1.a ),
    .Y(_1615_)
);

NAND2X1 _4972_ (
    .A(\z2.z3.z3.z1.b ),
    .B(_1615_),
    .Y(_1616_)
);

NAND2X1 _4973_ (
    .A(_1614_),
    .B(_1616_),
    .Y(\z2.z3.z3.z1.s )
);

NOR2X1 _4974_ (
    .A(_1613_),
    .B(_1615_),
    .Y(\z2.z3.z3.z1.c )
);

INVX1 _4975_ (
    .A(\z2.z3.z3.z1.c ),
    .Y(_1617_)
);

NAND2X1 _4976_ (
    .A(\z2.z3.z3.z2.a ),
    .B(_1617_),
    .Y(_1618_)
);

INVX1 _4977_ (
    .A(\z2.z3.z3.z2.a ),
    .Y(_1619_)
);

NAND2X1 _4978_ (
    .A(\z2.z3.z3.z1.c ),
    .B(_1619_),
    .Y(_1620_)
);

NAND2X1 _4979_ (
    .A(_1618_),
    .B(_1620_),
    .Y(\z2.z3.z3.z2.s )
);

NOR2X1 _4980_ (
    .A(_1617_),
    .B(_1619_),
    .Y(\z2.z3.z3.z2.c )
);

AND2X2 _4981_ (
    .A(b[6]),
    .B(a[10]),
    .Y(\z2.z3.q3 [0])
);

AND2X2 _4982_ (
    .A(b[6]),
    .B(a[11]),
    .Y(\z2.z3.z4.z1.a )
);

AND2X2 _4983_ (
    .A(a[10]),
    .B(b[7]),
    .Y(\z2.z3.z4.z1.b )
);

AND2X2 _4984_ (
    .A(a[11]),
    .B(b[7]),
    .Y(\z2.z3.z4.z2.a )
);

INVX1 _4985_ (
    .A(\z2.z3.z4.z1.b ),
    .Y(_1621_)
);

NAND2X1 _4986_ (
    .A(\z2.z3.z4.z1.a ),
    .B(_1621_),
    .Y(_1622_)
);

INVX1 _4987_ (
    .A(\z2.z3.z4.z1.a ),
    .Y(_1623_)
);

NAND2X1 _4988_ (
    .A(\z2.z3.z4.z1.b ),
    .B(_1623_),
    .Y(_1624_)
);

NAND2X1 _4989_ (
    .A(_1622_),
    .B(_1624_),
    .Y(\z2.z3.z4.z1.s )
);

NOR2X1 _4990_ (
    .A(_1621_),
    .B(_1623_),
    .Y(\z2.z3.z4.z1.c )
);

INVX1 _4991_ (
    .A(\z2.z3.z4.z1.c ),
    .Y(_1625_)
);

NAND2X1 _4992_ (
    .A(\z2.z3.z4.z2.a ),
    .B(_1625_),
    .Y(_1626_)
);

INVX1 _4993_ (
    .A(\z2.z3.z4.z2.a ),
    .Y(_1627_)
);

NAND2X1 _4994_ (
    .A(\z2.z3.z4.z1.c ),
    .B(_1627_),
    .Y(_1628_)
);

NAND2X1 _4995_ (
    .A(_1626_),
    .B(_1628_),
    .Y(\z2.z3.z4.z2.s )
);

NOR2X1 _4996_ (
    .A(_1625_),
    .B(_1627_),
    .Y(\z2.z3.z4.z2.c )
);

NOR2X1 _4997_ (
    .A(\z2.z4.q1 [0]),
    .B(\z2.z4.z1.z2.s ),
    .Y(_1636_)
);

AND2X2 _4998_ (
    .A(\z2.z4.q1 [0]),
    .B(\z2.z4.z1.z2.s ),
    .Y(_1637_)
);

NOR2X1 _4999_ (
    .A(_1636_),
    .B(_1637_),
    .Y(_1638_)
);

NAND2X1 _5000_ (
    .A(\z2.z4.q2 [0]),
    .B(_1638_),
    .Y(_1639_)
);

INVX1 _5001_ (
    .A(_1639_),
    .Y(_1640_)
);

NOR2X1 _5002_ (
    .A(\z2.z4.q2 [0]),
    .B(_1638_),
    .Y(_1641_)
);

NOR2X1 _5003_ (
    .A(_1641_),
    .B(_1640_),
    .Y(\z2.q3 [2])
);

NAND2X1 _5004_ (
    .A(\z2.z4.q1 [0]),
    .B(\z2.z4.z1.z2.s ),
    .Y(_1642_)
);

NOR2X1 _5005_ (
    .A(\z2.z4.z2.z1.s ),
    .B(\z2.z4.z1.z2.c ),
    .Y(_1643_)
);

NAND2X1 _5006_ (
    .A(\z2.z4.z2.z1.s ),
    .B(\z2.z4.z1.z2.c ),
    .Y(_1644_)
);

INVX1 _5007_ (
    .A(_1644_),
    .Y(_1645_)
);

OAI21X1 _5008_ (
    .A(_1643_),
    .B(_1645_),
    .C(_1642_),
    .Y(_1646_)
);

INVX1 _5009_ (
    .A(\z2.z4.z2.z1.s ),
    .Y(_1647_)
);

INVX1 _5010_ (
    .A(\z2.z4.z1.z2.c ),
    .Y(_1648_)
);

NAND2X1 _5011_ (
    .A(_1647_),
    .B(_1648_),
    .Y(_1649_)
);

NAND3X1 _5012_ (
    .A(_1637_),
    .B(_1644_),
    .C(_1649_),
    .Y(_1650_)
);

NAND3X1 _5013_ (
    .A(\z2.z4.z3.z1.s ),
    .B(_1650_),
    .C(_1646_),
    .Y(_1651_)
);

INVX1 _5014_ (
    .A(\z2.z4.z3.z1.s ),
    .Y(_1652_)
);

NAND2X1 _5015_ (
    .A(_1650_),
    .B(_1646_),
    .Y(_1653_)
);

NAND2X1 _5016_ (
    .A(_1652_),
    .B(_1653_),
    .Y(_1654_)
);

NAND3X1 _5017_ (
    .A(_1640_),
    .B(_1651_),
    .C(_1654_),
    .Y(_1655_)
);

INVX1 _5018_ (
    .A(_1655_),
    .Y(_1656_)
);

INVX1 _5019_ (
    .A(_1651_),
    .Y(_1657_)
);

OAI21X1 _5020_ (
    .A(_1642_),
    .B(_1643_),
    .C(_1644_),
    .Y(_1658_)
);

NAND2X1 _5021_ (
    .A(\z2.z4.z2.z2.s ),
    .B(_1658_),
    .Y(_1659_)
);

INVX1 _5022_ (
    .A(\z2.z4.z2.z2.s ),
    .Y(_1660_)
);

NAND3X1 _5023_ (
    .A(_1660_),
    .B(_1644_),
    .C(_1650_),
    .Y(_1661_)
);

NAND2X1 _5024_ (
    .A(\z2.z4.q3 [0]),
    .B(\z2.z4.z3.z2.s ),
    .Y(_1662_)
);

INVX1 _5025_ (
    .A(\z2.z4.q3 [0]),
    .Y(_1663_)
);

INVX1 _5026_ (
    .A(\z2.z4.z3.z2.s ),
    .Y(_1664_)
);

NAND2X1 _5027_ (
    .A(_1663_),
    .B(_1664_),
    .Y(_1665_)
);

NAND2X1 _5028_ (
    .A(_1662_),
    .B(_1665_),
    .Y(_1666_)
);

INVX1 _5029_ (
    .A(_1666_),
    .Y(_1667_)
);

NAND3X1 _5030_ (
    .A(_1659_),
    .B(_1667_),
    .C(_1661_),
    .Y(_1668_)
);

AND2X2 _5031_ (
    .A(_1658_),
    .B(\z2.z4.z2.z2.s ),
    .Y(_1669_)
);

NOR2X1 _5032_ (
    .A(\z2.z4.z2.z2.s ),
    .B(_1658_),
    .Y(_1670_)
);

OAI21X1 _5033_ (
    .A(_1670_),
    .B(_1669_),
    .C(_1666_),
    .Y(_1671_)
);

NAND3X1 _5034_ (
    .A(_1657_),
    .B(_1668_),
    .C(_1671_),
    .Y(_1672_)
);

INVX1 _5035_ (
    .A(_1668_),
    .Y(_1673_)
);

AOI21X1 _5036_ (
    .A(_1661_),
    .B(_1659_),
    .C(_1667_),
    .Y(_1674_)
);

OAI21X1 _5037_ (
    .A(_1674_),
    .B(_1673_),
    .C(_1651_),
    .Y(_1675_)
);

NAND3X1 _5038_ (
    .A(_1656_),
    .B(_1672_),
    .C(_1675_),
    .Y(_1676_)
);

INVX1 _5039_ (
    .A(_1672_),
    .Y(_1677_)
);

INVX1 _5040_ (
    .A(_1653_),
    .Y(_1678_)
);

AOI22X1 _5041_ (
    .A(\z2.z4.z3.z1.s ),
    .B(_1678_),
    .C(_1671_),
    .D(_1668_),
    .Y(_1679_)
);

OAI21X1 _5042_ (
    .A(_1679_),
    .B(_1677_),
    .C(_1655_),
    .Y(_1680_)
);

AND2X2 _5043_ (
    .A(_1680_),
    .B(_1676_),
    .Y(\z2.q3 [4])
);

OAI21X1 _5044_ (
    .A(_1655_),
    .B(_1679_),
    .C(_1672_),
    .Y(_1681_)
);

OAI21X1 _5045_ (
    .A(_1663_),
    .B(_1664_),
    .C(_1668_),
    .Y(_1682_)
);

NAND2X1 _5046_ (
    .A(\z2.z4.z4.z1.s ),
    .B(\z2.z4.z3.z2.c ),
    .Y(_1683_)
);

OR2X2 _5047_ (
    .A(\z2.z4.z4.z1.s ),
    .B(\z2.z4.z3.z2.c ),
    .Y(_1684_)
);

NAND2X1 _5048_ (
    .A(_1683_),
    .B(_1684_),
    .Y(_1685_)
);

INVX1 _5049_ (
    .A(_1685_),
    .Y(_1686_)
);

NAND2X1 _5050_ (
    .A(\z2.z4.z2.z2.c ),
    .B(_1669_),
    .Y(_1687_)
);

INVX1 _5051_ (
    .A(\z2.z4.z2.z2.c ),
    .Y(_1688_)
);

NAND2X1 _5052_ (
    .A(_1688_),
    .B(_1659_),
    .Y(_1689_)
);

NAND3X1 _5053_ (
    .A(_1686_),
    .B(_1689_),
    .C(_1687_),
    .Y(_1690_)
);

NAND2X1 _5054_ (
    .A(\z2.z4.z2.z2.c ),
    .B(_1659_),
    .Y(_1691_)
);

NAND2X1 _5055_ (
    .A(_1688_),
    .B(_1669_),
    .Y(_1692_)
);

NAND3X1 _5056_ (
    .A(_1685_),
    .B(_1691_),
    .C(_1692_),
    .Y(_1693_)
);

NAND3X1 _5057_ (
    .A(_1682_),
    .B(_1690_),
    .C(_1693_),
    .Y(_1694_)
);

INVX1 _5058_ (
    .A(_1682_),
    .Y(_1695_)
);

AOI21X1 _5059_ (
    .A(_1692_),
    .B(_1691_),
    .C(_1685_),
    .Y(_1696_)
);

AOI21X1 _5060_ (
    .A(_1687_),
    .B(_1689_),
    .C(_1686_),
    .Y(_1697_)
);

OAI21X1 _5061_ (
    .A(_1696_),
    .B(_1697_),
    .C(_1695_),
    .Y(_1698_)
);

NAND2X1 _5062_ (
    .A(_1694_),
    .B(_1698_),
    .Y(_1699_)
);

NAND2X1 _5063_ (
    .A(_1681_),
    .B(_1699_),
    .Y(_1700_)
);

OR2X2 _5064_ (
    .A(_1699_),
    .B(_1681_),
    .Y(_1701_)
);

NAND2X1 _5065_ (
    .A(_1700_),
    .B(_1701_),
    .Y(\z2.q3 [5])
);

INVX1 _5066_ (
    .A(\z2.z4.z4.z2.s ),
    .Y(_1702_)
);

INVX1 _5067_ (
    .A(_1683_),
    .Y(_1703_)
);

OAI21X1 _5068_ (
    .A(_1703_),
    .B(_1696_),
    .C(_1702_),
    .Y(_1704_)
);

NAND3X1 _5069_ (
    .A(\z2.z4.z4.z2.s ),
    .B(_1683_),
    .C(_1690_),
    .Y(_1705_)
);

NAND2X1 _5070_ (
    .A(_1698_),
    .B(_1681_),
    .Y(_1706_)
);

AOI22X1 _5071_ (
    .A(_1704_),
    .B(_1705_),
    .C(_1706_),
    .D(_1694_),
    .Y(_1707_)
);

NAND2X1 _5072_ (
    .A(_1705_),
    .B(_1704_),
    .Y(_1708_)
);

NAND3X1 _5073_ (
    .A(_1672_),
    .B(_1694_),
    .C(_1676_),
    .Y(_1709_)
);

AOI21X1 _5074_ (
    .A(_1709_),
    .B(_1698_),
    .C(_1708_),
    .Y(_1710_)
);

NOR2X1 _5075_ (
    .A(_1707_),
    .B(_1710_),
    .Y(\z2.q3 [6])
);

OAI21X1 _5076_ (
    .A(_1703_),
    .B(_1696_),
    .C(\z2.z4.z4.z2.s ),
    .Y(_1629_)
);

NAND3X1 _5077_ (
    .A(_1698_),
    .B(_1708_),
    .C(_1709_),
    .Y(_1630_)
);

NAND3X1 _5078_ (
    .A(\z2.z4.z4.z2.c ),
    .B(_1629_),
    .C(_1630_),
    .Y(_1631_)
);

INVX1 _5079_ (
    .A(\z2.z4.z4.z2.c ),
    .Y(_1632_)
);

INVX1 _5080_ (
    .A(_1629_),
    .Y(_1633_)
);

OAI21X1 _5081_ (
    .A(_1633_),
    .B(_1707_),
    .C(_1632_),
    .Y(_1634_)
);

NAND2X1 _5082_ (
    .A(_1631_),
    .B(_1634_),
    .Y(\z2.q3 [7])
);

AOI21X1 _5083_ (
    .A(_1654_),
    .B(_1651_),
    .C(_1640_),
    .Y(_1635_)
);

NOR2X1 _5084_ (
    .A(_1635_),
    .B(_1656_),
    .Y(\z2.q3 [3])
);

AND2X2 _5085_ (
    .A(b[4]),
    .B(a[12]),
    .Y(\z2.q3 [0])
);

AND2X2 _5086_ (
    .A(b[4]),
    .B(a[13]),
    .Y(\z2.z4.z1.z1.a )
);

AND2X2 _5087_ (
    .A(a[12]),
    .B(b[5]),
    .Y(\z2.z4.z1.z1.b )
);

AND2X2 _5088_ (
    .A(a[13]),
    .B(b[5]),
    .Y(\z2.z4.z1.z2.a )
);

INVX1 _5089_ (
    .A(\z2.z4.z1.z1.b ),
    .Y(_1711_)
);

NAND2X1 _5090_ (
    .A(\z2.z4.z1.z1.a ),
    .B(_1711_),
    .Y(_1712_)
);

INVX1 _5091_ (
    .A(\z2.z4.z1.z1.a ),
    .Y(_1713_)
);

NAND2X1 _5092_ (
    .A(\z2.z4.z1.z1.b ),
    .B(_1713_),
    .Y(_1714_)
);

NAND2X1 _5093_ (
    .A(_1712_),
    .B(_1714_),
    .Y(\z2.z4.z1.z1.s )
);

NOR2X1 _5094_ (
    .A(_1711_),
    .B(_1713_),
    .Y(\z2.z4.z1.z1.c )
);

INVX1 _5095_ (
    .A(\z2.z4.z1.z1.c ),
    .Y(_1715_)
);

NAND2X1 _5096_ (
    .A(\z2.z4.z1.z2.a ),
    .B(_1715_),
    .Y(_1716_)
);

INVX1 _5097_ (
    .A(\z2.z4.z1.z2.a ),
    .Y(_1717_)
);

NAND2X1 _5098_ (
    .A(\z2.z4.z1.z1.c ),
    .B(_1717_),
    .Y(_1718_)
);

NAND2X1 _5099_ (
    .A(_1716_),
    .B(_1718_),
    .Y(\z2.z4.z1.z2.s )
);

NOR2X1 _5100_ (
    .A(_1715_),
    .B(_1717_),
    .Y(\z2.z4.z1.z2.c )
);

AND2X2 _5101_ (
    .A(b[4]),
    .B(a[14]),
    .Y(\z2.z4.q1 [0])
);

AND2X2 _5102_ (
    .A(b[4]),
    .B(a[15]),
    .Y(\z2.z4.z2.z1.a )
);

AND2X2 _5103_ (
    .A(a[14]),
    .B(b[5]),
    .Y(\z2.z4.z2.z1.b )
);

AND2X2 _5104_ (
    .A(a[15]),
    .B(b[5]),
    .Y(\z2.z4.z2.z2.a )
);

INVX1 _5105_ (
    .A(\z2.z4.z2.z1.b ),
    .Y(_1719_)
);

NAND2X1 _5106_ (
    .A(\z2.z4.z2.z1.a ),
    .B(_1719_),
    .Y(_1720_)
);

INVX1 _5107_ (
    .A(\z2.z4.z2.z1.a ),
    .Y(_1721_)
);

NAND2X1 _5108_ (
    .A(\z2.z4.z2.z1.b ),
    .B(_1721_),
    .Y(_1722_)
);

NAND2X1 _5109_ (
    .A(_1720_),
    .B(_1722_),
    .Y(\z2.z4.z2.z1.s )
);

NOR2X1 _5110_ (
    .A(_1719_),
    .B(_1721_),
    .Y(\z2.z4.z2.z1.c )
);

INVX1 _5111_ (
    .A(\z2.z4.z2.z1.c ),
    .Y(_1723_)
);

NAND2X1 _5112_ (
    .A(\z2.z4.z2.z2.a ),
    .B(_1723_),
    .Y(_1724_)
);

INVX1 _5113_ (
    .A(\z2.z4.z2.z2.a ),
    .Y(_1725_)
);

NAND2X1 _5114_ (
    .A(\z2.z4.z2.z1.c ),
    .B(_1725_),
    .Y(_1726_)
);

NAND2X1 _5115_ (
    .A(_1724_),
    .B(_1726_),
    .Y(\z2.z4.z2.z2.s )
);

NOR2X1 _5116_ (
    .A(_1723_),
    .B(_1725_),
    .Y(\z2.z4.z2.z2.c )
);

AND2X2 _5117_ (
    .A(b[6]),
    .B(a[12]),
    .Y(\z2.z4.q2 [0])
);

AND2X2 _5118_ (
    .A(b[6]),
    .B(a[13]),
    .Y(\z2.z4.z3.z1.a )
);

AND2X2 _5119_ (
    .A(a[12]),
    .B(b[7]),
    .Y(\z2.z4.z3.z1.b )
);

AND2X2 _5120_ (
    .A(a[13]),
    .B(b[7]),
    .Y(\z2.z4.z3.z2.a )
);

INVX1 _5121_ (
    .A(\z2.z4.z3.z1.b ),
    .Y(_1727_)
);

NAND2X1 _5122_ (
    .A(\z2.z4.z3.z1.a ),
    .B(_1727_),
    .Y(_1728_)
);

INVX1 _5123_ (
    .A(\z2.z4.z3.z1.a ),
    .Y(_1729_)
);

NAND2X1 _5124_ (
    .A(\z2.z4.z3.z1.b ),
    .B(_1729_),
    .Y(_1730_)
);

NAND2X1 _5125_ (
    .A(_1728_),
    .B(_1730_),
    .Y(\z2.z4.z3.z1.s )
);

NOR2X1 _5126_ (
    .A(_1727_),
    .B(_1729_),
    .Y(\z2.z4.z3.z1.c )
);

INVX1 _5127_ (
    .A(\z2.z4.z3.z1.c ),
    .Y(_1731_)
);

NAND2X1 _5128_ (
    .A(\z2.z4.z3.z2.a ),
    .B(_1731_),
    .Y(_1732_)
);

INVX1 _5129_ (
    .A(\z2.z4.z3.z2.a ),
    .Y(_1733_)
);

NAND2X1 _5130_ (
    .A(\z2.z4.z3.z1.c ),
    .B(_1733_),
    .Y(_1734_)
);

NAND2X1 _5131_ (
    .A(_1732_),
    .B(_1734_),
    .Y(\z2.z4.z3.z2.s )
);

NOR2X1 _5132_ (
    .A(_1731_),
    .B(_1733_),
    .Y(\z2.z4.z3.z2.c )
);

AND2X2 _5133_ (
    .A(b[6]),
    .B(a[14]),
    .Y(\z2.z4.q3 [0])
);

AND2X2 _5134_ (
    .A(b[6]),
    .B(a[15]),
    .Y(\z2.z4.z4.z1.a )
);

AND2X2 _5135_ (
    .A(a[14]),
    .B(b[7]),
    .Y(\z2.z4.z4.z1.b )
);

AND2X2 _5136_ (
    .A(a[15]),
    .B(b[7]),
    .Y(\z2.z4.z4.z2.a )
);

INVX1 _5137_ (
    .A(\z2.z4.z4.z1.b ),
    .Y(_1735_)
);

NAND2X1 _5138_ (
    .A(\z2.z4.z4.z1.a ),
    .B(_1735_),
    .Y(_1736_)
);

INVX1 _5139_ (
    .A(\z2.z4.z4.z1.a ),
    .Y(_1737_)
);

NAND2X1 _5140_ (
    .A(\z2.z4.z4.z1.b ),
    .B(_1737_),
    .Y(_1738_)
);

NAND2X1 _5141_ (
    .A(_1736_),
    .B(_1738_),
    .Y(\z2.z4.z4.z1.s )
);

NOR2X1 _5142_ (
    .A(_1735_),
    .B(_1737_),
    .Y(\z2.z4.z4.z1.c )
);

INVX1 _5143_ (
    .A(\z2.z4.z4.z1.c ),
    .Y(_1739_)
);

NAND2X1 _5144_ (
    .A(\z2.z4.z4.z2.a ),
    .B(_1739_),
    .Y(_1740_)
);

INVX1 _5145_ (
    .A(\z2.z4.z4.z2.a ),
    .Y(_1741_)
);

NAND2X1 _5146_ (
    .A(\z2.z4.z4.z1.c ),
    .B(_1741_),
    .Y(_1742_)
);

NAND2X1 _5147_ (
    .A(_1740_),
    .B(_1742_),
    .Y(\z2.z4.z4.z2.s )
);

NOR2X1 _5148_ (
    .A(_1739_),
    .B(_1741_),
    .Y(\z2.z4.z4.z2.c )
);

OR2X2 _5149_ (
    .A(\z3.q1 [0]),
    .B(\z3.q0 [4]),
    .Y(_1885_)
);

NAND2X1 _5150_ (
    .A(\z3.q1 [0]),
    .B(\z3.q0 [4]),
    .Y(_1886_)
);

NAND2X1 _5151_ (
    .A(_1886_),
    .B(_1885_),
    .Y(_1887_)
);

INVX1 _5152_ (
    .A(_1887_),
    .Y(_1888_)
);

AND2X2 _5153_ (
    .A(_1888_),
    .B(\z3.q2 [0]),
    .Y(_1889_)
);

NOR2X1 _5154_ (
    .A(\z3.q2 [0]),
    .B(_1888_),
    .Y(_1890_)
);

NOR2X1 _5155_ (
    .A(_1890_),
    .B(_1889_),
    .Y(q2[4])
);

INVX1 _5156_ (
    .A(\z3.z3.z1.z1.s ),
    .Y(_1891_)
);

INVX1 _5157_ (
    .A(_1886_),
    .Y(_1892_)
);

NAND2X1 _5158_ (
    .A(\z3.z2.z1.z1.s ),
    .B(\z3.q0 [5]),
    .Y(_1893_)
);

OR2X2 _5159_ (
    .A(\z3.z2.z1.z1.s ),
    .B(\z3.q0 [5]),
    .Y(_1894_)
);

NAND3X1 _5160_ (
    .A(_1893_),
    .B(_1894_),
    .C(_1892_),
    .Y(_1895_)
);

AND2X2 _5161_ (
    .A(\z3.z2.z1.z1.s ),
    .B(\z3.q0 [5]),
    .Y(_1896_)
);

NOR2X1 _5162_ (
    .A(\z3.z2.z1.z1.s ),
    .B(\z3.q0 [5]),
    .Y(_1897_)
);

OAI21X1 _5163_ (
    .A(_1897_),
    .B(_1896_),
    .C(_1886_),
    .Y(_1898_)
);

NAND2X1 _5164_ (
    .A(_1898_),
    .B(_1895_),
    .Y(_1899_)
);

OR2X2 _5165_ (
    .A(_1899_),
    .B(_1891_),
    .Y(_1900_)
);

NAND2X1 _5166_ (
    .A(_1891_),
    .B(_1899_),
    .Y(_1901_)
);

AND2X2 _5167_ (
    .A(_1900_),
    .B(_1901_),
    .Y(_1902_)
);

NAND2X1 _5168_ (
    .A(_1889_),
    .B(_1902_),
    .Y(_1903_)
);

INVX1 _5169_ (
    .A(_1900_),
    .Y(_1904_)
);

OAI21X1 _5170_ (
    .A(_1886_),
    .B(_1897_),
    .C(_1893_),
    .Y(_1905_)
);

INVX1 _5171_ (
    .A(\z3.q0 [6]),
    .Y(_1906_)
);

NOR2X1 _5172_ (
    .A(\z3.q1 [2]),
    .B(_1906_),
    .Y(_1907_)
);

INVX1 _5173_ (
    .A(\z3.q1 [2]),
    .Y(_1908_)
);

NOR2X1 _5174_ (
    .A(\z3.q0 [6]),
    .B(_1908_),
    .Y(_1909_)
);

OAI21X1 _5175_ (
    .A(_1907_),
    .B(_1909_),
    .C(_1905_),
    .Y(_1910_)
);

NAND2X1 _5176_ (
    .A(\z3.q0 [6]),
    .B(_1908_),
    .Y(_1911_)
);

NAND2X1 _5177_ (
    .A(\z3.q1 [2]),
    .B(_1906_),
    .Y(_1912_)
);

NAND2X1 _5178_ (
    .A(_1911_),
    .B(_1912_),
    .Y(_1913_)
);

OR2X2 _5179_ (
    .A(_1913_),
    .B(_1905_),
    .Y(_1914_)
);

NAND3X1 _5180_ (
    .A(\z3.q2 [2]),
    .B(_1910_),
    .C(_1914_),
    .Y(_1915_)
);

INVX1 _5181_ (
    .A(\z3.q2 [2]),
    .Y(_1916_)
);

NAND2X1 _5182_ (
    .A(_1910_),
    .B(_1914_),
    .Y(_1917_)
);

NAND2X1 _5183_ (
    .A(_1916_),
    .B(_1917_),
    .Y(_1918_)
);

AOI21X1 _5184_ (
    .A(_1918_),
    .B(_1915_),
    .C(_1904_),
    .Y(_1919_)
);

INVX1 _5185_ (
    .A(_1919_),
    .Y(_1920_)
);

NAND3X1 _5186_ (
    .A(_1915_),
    .B(_1918_),
    .C(_1904_),
    .Y(_1921_)
);

NAND3X1 _5187_ (
    .A(_1903_),
    .B(_1921_),
    .C(_1920_),
    .Y(_1922_)
);

INVX1 _5188_ (
    .A(_1903_),
    .Y(_1923_)
);

INVX1 _5189_ (
    .A(_1921_),
    .Y(_1924_)
);

OAI21X1 _5190_ (
    .A(_1919_),
    .B(_1924_),
    .C(_1923_),
    .Y(_1925_)
);

NAND2X1 _5191_ (
    .A(_1922_),
    .B(_1925_),
    .Y(q2[6])
);

OAI21X1 _5192_ (
    .A(_1919_),
    .B(_1903_),
    .C(_1921_),
    .Y(_1926_)
);

INVX1 _5193_ (
    .A(_1915_),
    .Y(_1927_)
);

INVX1 _5194_ (
    .A(\z3.q2 [3]),
    .Y(_1928_)
);

INVX1 _5195_ (
    .A(\z3.q0 [7]),
    .Y(_1929_)
);

NOR2X1 _5196_ (
    .A(\z3.q1 [3]),
    .B(_1929_),
    .Y(_1930_)
);

INVX1 _5197_ (
    .A(\z3.q1 [3]),
    .Y(_1931_)
);

NOR2X1 _5198_ (
    .A(\z3.q0 [7]),
    .B(_1931_),
    .Y(_1932_)
);

NAND2X1 _5199_ (
    .A(\z3.q1 [2]),
    .B(\z3.q0 [6]),
    .Y(_1933_)
);

INVX1 _5200_ (
    .A(_1933_),
    .Y(_1934_)
);

AOI21X1 _5201_ (
    .A(_1913_),
    .B(_1905_),
    .C(_1934_),
    .Y(_1935_)
);

OAI21X1 _5202_ (
    .A(_1930_),
    .B(_1932_),
    .C(_1935_),
    .Y(_1936_)
);

NAND2X1 _5203_ (
    .A(\z3.q1 [3]),
    .B(\z3.q0 [7]),
    .Y(_1937_)
);

INVX1 _5204_ (
    .A(_1937_),
    .Y(_1938_)
);

NOR2X1 _5205_ (
    .A(\z3.q1 [3]),
    .B(\z3.q0 [7]),
    .Y(_1939_)
);

INVX1 _5206_ (
    .A(_1935_),
    .Y(_1940_)
);

OAI21X1 _5207_ (
    .A(_1938_),
    .B(_1939_),
    .C(_1940_),
    .Y(_1941_)
);

AOI21X1 _5208_ (
    .A(_1941_),
    .B(_1936_),
    .C(_1928_),
    .Y(_1743_)
);

INVX1 _5209_ (
    .A(_1743_),
    .Y(_1744_)
);

NAND3X1 _5210_ (
    .A(_1928_),
    .B(_1936_),
    .C(_1941_),
    .Y(_1745_)
);

AOI21X1 _5211_ (
    .A(_1744_),
    .B(_1745_),
    .C(_1927_),
    .Y(_1746_)
);

NAND3X1 _5212_ (
    .A(_1927_),
    .B(_1745_),
    .C(_1744_),
    .Y(_1747_)
);

INVX1 _5213_ (
    .A(_1747_),
    .Y(_1748_)
);

OAI21X1 _5214_ (
    .A(_1746_),
    .B(_1748_),
    .C(_1926_),
    .Y(_1749_)
);

INVX1 _5215_ (
    .A(_1926_),
    .Y(_1750_)
);

NAND2X1 _5216_ (
    .A(_1745_),
    .B(_1744_),
    .Y(_1751_)
);

OAI21X1 _5217_ (
    .A(_1916_),
    .B(_1917_),
    .C(_1751_),
    .Y(_1752_)
);

NAND3X1 _5218_ (
    .A(_1747_),
    .B(_1750_),
    .C(_1752_),
    .Y(_1753_)
);

NAND2X1 _5219_ (
    .A(_1753_),
    .B(_1749_),
    .Y(q2[7])
);

AOI21X1 _5220_ (
    .A(_1752_),
    .B(_1926_),
    .C(_1748_),
    .Y(_1754_)
);

AOI21X1 _5221_ (
    .A(_1892_),
    .B(_1894_),
    .C(_1896_),
    .Y(_1755_)
);

OAI22X1 _5222_ (
    .A(_1907_),
    .B(_1909_),
    .C(_1930_),
    .D(_1932_),
    .Y(_1756_)
);

OAI21X1 _5223_ (
    .A(_1933_),
    .B(_1939_),
    .C(_1937_),
    .Y(_1757_)
);

INVX1 _5224_ (
    .A(_1757_),
    .Y(_1758_)
);

OAI21X1 _5225_ (
    .A(_1755_),
    .B(_1756_),
    .C(_1758_),
    .Y(_1759_)
);

NAND2X1 _5226_ (
    .A(\z3.q1 [4]),
    .B(_1759_),
    .Y(_1760_)
);

INVX1 _5227_ (
    .A(\z3.q1 [4]),
    .Y(_1761_)
);

NAND2X1 _5228_ (
    .A(\z3.q0 [7]),
    .B(_1931_),
    .Y(_1762_)
);

NAND2X1 _5229_ (
    .A(\z3.q1 [3]),
    .B(_1929_),
    .Y(_1763_)
);

NAND2X1 _5230_ (
    .A(_1762_),
    .B(_1763_),
    .Y(_1764_)
);

NAND3X1 _5231_ (
    .A(_1905_),
    .B(_1913_),
    .C(_1764_),
    .Y(_1765_)
);

NAND3X1 _5232_ (
    .A(_1761_),
    .B(_1758_),
    .C(_1765_),
    .Y(_1766_)
);

NAND2X1 _5233_ (
    .A(\z3.q3 [0]),
    .B(\z3.q2 [4]),
    .Y(_1767_)
);

INVX1 _5234_ (
    .A(\z3.q3 [0]),
    .Y(_1768_)
);

INVX1 _5235_ (
    .A(\z3.q2 [4]),
    .Y(_1769_)
);

NAND2X1 _5236_ (
    .A(_1768_),
    .B(_1769_),
    .Y(_1770_)
);

NAND2X1 _5237_ (
    .A(_1767_),
    .B(_1770_),
    .Y(_1771_)
);

INVX1 _5238_ (
    .A(_1771_),
    .Y(_1772_)
);

NAND3X1 _5239_ (
    .A(_1766_),
    .B(_1772_),
    .C(_1760_),
    .Y(_1773_)
);

AOI21X1 _5240_ (
    .A(_1765_),
    .B(_1758_),
    .C(_1761_),
    .Y(_1774_)
);

INVX1 _5241_ (
    .A(_1766_),
    .Y(_1775_)
);

OAI21X1 _5242_ (
    .A(_1774_),
    .B(_1775_),
    .C(_1771_),
    .Y(_1776_)
);

NAND3X1 _5243_ (
    .A(_1773_),
    .B(_1776_),
    .C(_1743_),
    .Y(_1777_)
);

NAND2X1 _5244_ (
    .A(_1773_),
    .B(_1776_),
    .Y(_1778_)
);

NAND2X1 _5245_ (
    .A(_1778_),
    .B(_1744_),
    .Y(_1779_)
);

AND2X2 _5246_ (
    .A(_1779_),
    .B(_1777_),
    .Y(_1780_)
);

NAND2X1 _5247_ (
    .A(_1780_),
    .B(_1754_),
    .Y(_1781_)
);

OAI21X1 _5248_ (
    .A(_1746_),
    .B(_1750_),
    .C(_1747_),
    .Y(_1782_)
);

NAND2X1 _5249_ (
    .A(_1777_),
    .B(_1779_),
    .Y(_1783_)
);

NAND2X1 _5250_ (
    .A(_1783_),
    .B(_1782_),
    .Y(_1784_)
);

NAND2X1 _5251_ (
    .A(_1781_),
    .B(_1784_),
    .Y(q2[8])
);

OAI21X1 _5252_ (
    .A(_1783_),
    .B(_1754_),
    .C(_1777_),
    .Y(_1785_)
);

OAI21X1 _5253_ (
    .A(_1768_),
    .B(_1769_),
    .C(_1773_),
    .Y(_1786_)
);

NAND3X1 _5254_ (
    .A(\z3.q1 [4]),
    .B(\z3.q1 [5]),
    .C(_1759_),
    .Y(_1787_)
);

INVX1 _5255_ (
    .A(\z3.q1 [5]),
    .Y(_1788_)
);

AOI22X1 _5256_ (
    .A(_1911_),
    .B(_1912_),
    .C(_1762_),
    .D(_1763_),
    .Y(_1789_)
);

AOI21X1 _5257_ (
    .A(_1789_),
    .B(_1905_),
    .C(_1757_),
    .Y(_1790_)
);

OAI21X1 _5258_ (
    .A(_1761_),
    .B(_1790_),
    .C(_1788_),
    .Y(_1791_)
);

INVX1 _5259_ (
    .A(\z3.z4.z1.z1.s ),
    .Y(_1792_)
);

INVX1 _5260_ (
    .A(\z3.q2 [5]),
    .Y(_1793_)
);

NAND2X1 _5261_ (
    .A(_1792_),
    .B(_1793_),
    .Y(_1794_)
);

NAND2X1 _5262_ (
    .A(\z3.z4.z1.z1.s ),
    .B(\z3.q2 [5]),
    .Y(_1795_)
);

AND2X2 _5263_ (
    .A(_1794_),
    .B(_1795_),
    .Y(_1796_)
);

NAND3X1 _5264_ (
    .A(_1796_),
    .B(_1791_),
    .C(_1787_),
    .Y(_1797_)
);

AOI21X1 _5265_ (
    .A(_1787_),
    .B(_1791_),
    .C(_1796_),
    .Y(_1798_)
);

INVX1 _5266_ (
    .A(_1798_),
    .Y(_1799_)
);

NAND3X1 _5267_ (
    .A(_1797_),
    .B(_1786_),
    .C(_1799_),
    .Y(_1800_)
);

AND2X2 _5268_ (
    .A(_1773_),
    .B(_1767_),
    .Y(_1801_)
);

INVX1 _5269_ (
    .A(_1797_),
    .Y(_1802_)
);

OAI21X1 _5270_ (
    .A(_1802_),
    .B(_1798_),
    .C(_1801_),
    .Y(_1803_)
);

NAND2X1 _5271_ (
    .A(_1800_),
    .B(_1803_),
    .Y(_1804_)
);

OR2X2 _5272_ (
    .A(_1785_),
    .B(_1804_),
    .Y(_1805_)
);

NAND2X1 _5273_ (
    .A(_1804_),
    .B(_1785_),
    .Y(_1806_)
);

NAND2X1 _5274_ (
    .A(_1806_),
    .B(_1805_),
    .Y(q2[9])
);

NAND3X1 _5275_ (
    .A(_1800_),
    .B(_1803_),
    .C(_1780_),
    .Y(_1807_)
);

OAI21X1 _5276_ (
    .A(_1744_),
    .B(_1778_),
    .C(_1800_),
    .Y(_1808_)
);

NAND2X1 _5277_ (
    .A(_1803_),
    .B(_1808_),
    .Y(_1809_)
);

OAI21X1 _5278_ (
    .A(_1754_),
    .B(_1807_),
    .C(_1809_),
    .Y(_1810_)
);

OAI21X1 _5279_ (
    .A(_1792_),
    .B(_1793_),
    .C(_1797_),
    .Y(_1811_)
);

NAND3X1 _5280_ (
    .A(\z3.q1 [5]),
    .B(\z3.q1 [6]),
    .C(_1774_),
    .Y(_1812_)
);

INVX1 _5281_ (
    .A(\z3.q1 [6]),
    .Y(_1813_)
);

NAND2X1 _5282_ (
    .A(_1813_),
    .B(_1787_),
    .Y(_1814_)
);

INVX1 _5283_ (
    .A(\z3.q3 [2]),
    .Y(_1815_)
);

INVX1 _5284_ (
    .A(\z3.q2 [6]),
    .Y(_1816_)
);

NAND2X1 _5285_ (
    .A(_1815_),
    .B(_1816_),
    .Y(_1817_)
);

NAND2X1 _5286_ (
    .A(\z3.q3 [2]),
    .B(\z3.q2 [6]),
    .Y(_1818_)
);

NAND2X1 _5287_ (
    .A(_1818_),
    .B(_1817_),
    .Y(_1819_)
);

INVX1 _5288_ (
    .A(_1819_),
    .Y(_1820_)
);

NAND3X1 _5289_ (
    .A(_1812_),
    .B(_1820_),
    .C(_1814_),
    .Y(_1821_)
);

AOI21X1 _5290_ (
    .A(_1814_),
    .B(_1812_),
    .C(_1820_),
    .Y(_1822_)
);

INVX1 _5291_ (
    .A(_1822_),
    .Y(_1823_)
);

NAND3X1 _5292_ (
    .A(_1811_),
    .B(_1821_),
    .C(_1823_),
    .Y(_1824_)
);

INVX1 _5293_ (
    .A(_1811_),
    .Y(_1825_)
);

INVX1 _5294_ (
    .A(_1821_),
    .Y(_1826_)
);

OAI21X1 _5295_ (
    .A(_1822_),
    .B(_1826_),
    .C(_1825_),
    .Y(_1827_)
);

NAND2X1 _5296_ (
    .A(_1827_),
    .B(_1824_),
    .Y(_1828_)
);

NAND2X1 _5297_ (
    .A(_1828_),
    .B(_1810_),
    .Y(_1829_)
);

NOR2X1 _5298_ (
    .A(_1783_),
    .B(_1804_),
    .Y(_1830_)
);

AOI22X1 _5299_ (
    .A(_1803_),
    .B(_1808_),
    .C(_1830_),
    .D(_1782_),
    .Y(_1831_)
);

AND2X2 _5300_ (
    .A(_1824_),
    .B(_1827_),
    .Y(_1832_)
);

NAND2X1 _5301_ (
    .A(_1832_),
    .B(_1831_),
    .Y(_1833_)
);

NAND2X1 _5302_ (
    .A(_1829_),
    .B(_1833_),
    .Y(q2[10])
);

OAI21X1 _5303_ (
    .A(_1828_),
    .B(_1831_),
    .C(_1824_),
    .Y(_1834_)
);

OAI21X1 _5304_ (
    .A(_1815_),
    .B(_1816_),
    .C(_1821_),
    .Y(_1835_)
);

NOR2X1 _5305_ (
    .A(\z3.q3 [3]),
    .B(\z3.q2 [7]),
    .Y(_1836_)
);

INVX1 _5306_ (
    .A(\z3.q3 [3]),
    .Y(_1837_)
);

INVX1 _5307_ (
    .A(\z3.q2 [7]),
    .Y(_1838_)
);

NOR2X1 _5308_ (
    .A(_1837_),
    .B(_1838_),
    .Y(_1839_)
);

NOR2X1 _5309_ (
    .A(_1836_),
    .B(_1839_),
    .Y(_1840_)
);

INVX1 _5310_ (
    .A(\z3.q1 [7]),
    .Y(_1841_)
);

OAI21X1 _5311_ (
    .A(_1813_),
    .B(_1787_),
    .C(_1841_),
    .Y(_1842_)
);

AND2X2 _5312_ (
    .A(_1774_),
    .B(\z3.q1 [5]),
    .Y(_1843_)
);

NAND3X1 _5313_ (
    .A(\z3.q1 [6]),
    .B(\z3.q1 [7]),
    .C(_1843_),
    .Y(_1844_)
);

NAND3X1 _5314_ (
    .A(_1840_),
    .B(_1842_),
    .C(_1844_),
    .Y(_1845_)
);

INVX1 _5315_ (
    .A(_1840_),
    .Y(_1846_)
);

OAI21X1 _5316_ (
    .A(_1813_),
    .B(_1787_),
    .C(\z3.q1 [7]),
    .Y(_1847_)
);

NAND3X1 _5317_ (
    .A(\z3.q1 [6]),
    .B(_1841_),
    .C(_1843_),
    .Y(_1848_)
);

NAND3X1 _5318_ (
    .A(_1846_),
    .B(_1847_),
    .C(_1848_),
    .Y(_1849_)
);

NAND3X1 _5319_ (
    .A(_1845_),
    .B(_1849_),
    .C(_1835_),
    .Y(_1850_)
);

AND2X2 _5320_ (
    .A(_1821_),
    .B(_1818_),
    .Y(_1851_)
);

NAND2X1 _5321_ (
    .A(_1845_),
    .B(_1849_),
    .Y(_1852_)
);

NAND2X1 _5322_ (
    .A(_1851_),
    .B(_1852_),
    .Y(_1853_)
);

NAND2X1 _5323_ (
    .A(_1850_),
    .B(_1853_),
    .Y(_1854_)
);

OR2X2 _5324_ (
    .A(_1834_),
    .B(_1854_),
    .Y(_1855_)
);

NAND2X1 _5325_ (
    .A(_1854_),
    .B(_1834_),
    .Y(_1856_)
);

NAND2X1 _5326_ (
    .A(_1856_),
    .B(_1855_),
    .Y(q2[11])
);

OAI21X1 _5327_ (
    .A(_1851_),
    .B(_1852_),
    .C(_1824_),
    .Y(_1857_)
);

NAND2X1 _5328_ (
    .A(_1853_),
    .B(_1857_),
    .Y(_1858_)
);

NAND3X1 _5329_ (
    .A(_1850_),
    .B(_1853_),
    .C(_1832_),
    .Y(_1859_)
);

OAI21X1 _5330_ (
    .A(_1859_),
    .B(_1831_),
    .C(_1858_),
    .Y(_1860_)
);

OAI21X1 _5331_ (
    .A(_1837_),
    .B(_1838_),
    .C(_1845_),
    .Y(_1861_)
);

NAND2X1 _5332_ (
    .A(\z3.q3 [4]),
    .B(_1861_),
    .Y(_1862_)
);

OR2X2 _5333_ (
    .A(_1861_),
    .B(\z3.q3 [4]),
    .Y(_1863_)
);

NAND3X1 _5334_ (
    .A(_1862_),
    .B(_1863_),
    .C(_1860_),
    .Y(_1864_)
);

NOR2X1 _5335_ (
    .A(_1828_),
    .B(_1854_),
    .Y(_1865_)
);

AOI22X1 _5336_ (
    .A(_1853_),
    .B(_1857_),
    .C(_1865_),
    .D(_1810_),
    .Y(_1866_)
);

NAND2X1 _5337_ (
    .A(_1862_),
    .B(_1863_),
    .Y(_1867_)
);

NAND2X1 _5338_ (
    .A(_1867_),
    .B(_1866_),
    .Y(_1868_)
);

AND2X2 _5339_ (
    .A(_1864_),
    .B(_1868_),
    .Y(q2[12])
);

INVX1 _5340_ (
    .A(\z3.q3 [5]),
    .Y(_1869_)
);

OAI21X1 _5341_ (
    .A(_1867_),
    .B(_1866_),
    .C(_1862_),
    .Y(_1870_)
);

NAND2X1 _5342_ (
    .A(_1869_),
    .B(_1870_),
    .Y(_1871_)
);

NAND3X1 _5343_ (
    .A(\z3.q3 [5]),
    .B(_1862_),
    .C(_1864_),
    .Y(_1872_)
);

NAND2X1 _5344_ (
    .A(_1872_),
    .B(_1871_),
    .Y(q2[13])
);

INVX1 _5345_ (
    .A(\z3.q3 [6]),
    .Y(_1873_)
);

NAND3X1 _5346_ (
    .A(\z3.q3 [5]),
    .B(_1862_),
    .C(_1863_),
    .Y(_1874_)
);

OAI22X1 _5347_ (
    .A(_1869_),
    .B(_1862_),
    .C(_1874_),
    .D(_1866_),
    .Y(_1875_)
);

NAND2X1 _5348_ (
    .A(_1873_),
    .B(_1875_),
    .Y(_1876_)
);

INVX1 _5349_ (
    .A(_1862_),
    .Y(_1877_)
);

INVX1 _5350_ (
    .A(_1874_),
    .Y(_1878_)
);

AOI22X1 _5351_ (
    .A(\z3.q3 [5]),
    .B(_1877_),
    .C(_1860_),
    .D(_1878_),
    .Y(_1879_)
);

NAND2X1 _5352_ (
    .A(\z3.q3 [6]),
    .B(_1879_),
    .Y(_1880_)
);

NAND2X1 _5353_ (
    .A(_1880_),
    .B(_1876_),
    .Y(q2[14])
);

OAI21X1 _5354_ (
    .A(_1873_),
    .B(_1879_),
    .C(\z3.q3 [7]),
    .Y(_1881_)
);

INVX1 _5355_ (
    .A(\z3.q3 [7]),
    .Y(_1882_)
);

NAND3X1 _5356_ (
    .A(\z3.q3 [6]),
    .B(_1882_),
    .C(_1875_),
    .Y(_1883_)
);

NAND2X1 _5357_ (
    .A(_1883_),
    .B(_1881_),
    .Y(q2[15])
);

NOR2X1 _5358_ (
    .A(_1889_),
    .B(_1902_),
    .Y(_1884_)
);

NOR2X1 _5359_ (
    .A(_1884_),
    .B(_1923_),
    .Y(q2[5])
);

NOR2X1 _5360_ (
    .A(\z3.z1.q1 [0]),
    .B(\z3.z1.z1.z2.s ),
    .Y(_1949_)
);

AND2X2 _5361_ (
    .A(\z3.z1.q1 [0]),
    .B(\z3.z1.z1.z2.s ),
    .Y(_1950_)
);

NOR2X1 _5362_ (
    .A(_1949_),
    .B(_1950_),
    .Y(_1951_)
);

NAND2X1 _5363_ (
    .A(\z3.z1.q2 [0]),
    .B(_1951_),
    .Y(_1952_)
);

INVX1 _5364_ (
    .A(_1952_),
    .Y(_1953_)
);

NOR2X1 _5365_ (
    .A(\z3.z1.q2 [0]),
    .B(_1951_),
    .Y(_1954_)
);

NOR2X1 _5366_ (
    .A(_1954_),
    .B(_1953_),
    .Y(q2[2])
);

NAND2X1 _5367_ (
    .A(\z3.z1.q1 [0]),
    .B(\z3.z1.z1.z2.s ),
    .Y(_1955_)
);

NOR2X1 _5368_ (
    .A(\z3.z1.z2.z1.s ),
    .B(\z3.z1.z1.z2.c ),
    .Y(_1956_)
);

NAND2X1 _5369_ (
    .A(\z3.z1.z2.z1.s ),
    .B(\z3.z1.z1.z2.c ),
    .Y(_1957_)
);

INVX1 _5370_ (
    .A(_1957_),
    .Y(_1958_)
);

OAI21X1 _5371_ (
    .A(_1956_),
    .B(_1958_),
    .C(_1955_),
    .Y(_1959_)
);

INVX1 _5372_ (
    .A(\z3.z1.z2.z1.s ),
    .Y(_1960_)
);

INVX1 _5373_ (
    .A(\z3.z1.z1.z2.c ),
    .Y(_1961_)
);

NAND2X1 _5374_ (
    .A(_1960_),
    .B(_1961_),
    .Y(_1962_)
);

NAND3X1 _5375_ (
    .A(_1950_),
    .B(_1957_),
    .C(_1962_),
    .Y(_1963_)
);

NAND3X1 _5376_ (
    .A(\z3.z1.z3.z1.s ),
    .B(_1963_),
    .C(_1959_),
    .Y(_1964_)
);

INVX1 _5377_ (
    .A(\z3.z1.z3.z1.s ),
    .Y(_1965_)
);

NAND2X1 _5378_ (
    .A(_1963_),
    .B(_1959_),
    .Y(_1966_)
);

NAND2X1 _5379_ (
    .A(_1965_),
    .B(_1966_),
    .Y(_1967_)
);

NAND3X1 _5380_ (
    .A(_1953_),
    .B(_1964_),
    .C(_1967_),
    .Y(_1968_)
);

INVX1 _5381_ (
    .A(_1968_),
    .Y(_1969_)
);

INVX1 _5382_ (
    .A(_1964_),
    .Y(_1970_)
);

OAI21X1 _5383_ (
    .A(_1955_),
    .B(_1956_),
    .C(_1957_),
    .Y(_1971_)
);

NAND2X1 _5384_ (
    .A(\z3.z1.z2.z2.s ),
    .B(_1971_),
    .Y(_1972_)
);

INVX1 _5385_ (
    .A(\z3.z1.z2.z2.s ),
    .Y(_1973_)
);

NAND3X1 _5386_ (
    .A(_1973_),
    .B(_1957_),
    .C(_1963_),
    .Y(_1974_)
);

NAND2X1 _5387_ (
    .A(\z3.z1.q3 [0]),
    .B(\z3.z1.z3.z2.s ),
    .Y(_1975_)
);

INVX1 _5388_ (
    .A(\z3.z1.q3 [0]),
    .Y(_1976_)
);

INVX1 _5389_ (
    .A(\z3.z1.z3.z2.s ),
    .Y(_1977_)
);

NAND2X1 _5390_ (
    .A(_1976_),
    .B(_1977_),
    .Y(_1978_)
);

NAND2X1 _5391_ (
    .A(_1975_),
    .B(_1978_),
    .Y(_1979_)
);

INVX1 _5392_ (
    .A(_1979_),
    .Y(_1980_)
);

NAND3X1 _5393_ (
    .A(_1972_),
    .B(_1980_),
    .C(_1974_),
    .Y(_1981_)
);

AND2X2 _5394_ (
    .A(_1971_),
    .B(\z3.z1.z2.z2.s ),
    .Y(_1982_)
);

NOR2X1 _5395_ (
    .A(\z3.z1.z2.z2.s ),
    .B(_1971_),
    .Y(_1983_)
);

OAI21X1 _5396_ (
    .A(_1983_),
    .B(_1982_),
    .C(_1979_),
    .Y(_1984_)
);

NAND3X1 _5397_ (
    .A(_1970_),
    .B(_1981_),
    .C(_1984_),
    .Y(_1985_)
);

INVX1 _5398_ (
    .A(_1981_),
    .Y(_1986_)
);

AOI21X1 _5399_ (
    .A(_1974_),
    .B(_1972_),
    .C(_1980_),
    .Y(_1987_)
);

OAI21X1 _5400_ (
    .A(_1987_),
    .B(_1986_),
    .C(_1964_),
    .Y(_1988_)
);

NAND3X1 _5401_ (
    .A(_1969_),
    .B(_1985_),
    .C(_1988_),
    .Y(_1989_)
);

INVX1 _5402_ (
    .A(_1985_),
    .Y(_1990_)
);

INVX1 _5403_ (
    .A(_1966_),
    .Y(_1991_)
);

AOI22X1 _5404_ (
    .A(\z3.z1.z3.z1.s ),
    .B(_1991_),
    .C(_1984_),
    .D(_1981_),
    .Y(_1992_)
);

OAI21X1 _5405_ (
    .A(_1992_),
    .B(_1990_),
    .C(_1968_),
    .Y(_1993_)
);

AND2X2 _5406_ (
    .A(_1993_),
    .B(_1989_),
    .Y(\z3.q0 [4])
);

OAI21X1 _5407_ (
    .A(_1968_),
    .B(_1992_),
    .C(_1985_),
    .Y(_1994_)
);

OAI21X1 _5408_ (
    .A(_1976_),
    .B(_1977_),
    .C(_1981_),
    .Y(_1995_)
);

NAND2X1 _5409_ (
    .A(\z3.z1.z4.z1.s ),
    .B(\z3.z1.z3.z2.c ),
    .Y(_1996_)
);

OR2X2 _5410_ (
    .A(\z3.z1.z4.z1.s ),
    .B(\z3.z1.z3.z2.c ),
    .Y(_1997_)
);

NAND2X1 _5411_ (
    .A(_1996_),
    .B(_1997_),
    .Y(_1998_)
);

INVX1 _5412_ (
    .A(_1998_),
    .Y(_1999_)
);

NAND2X1 _5413_ (
    .A(\z3.z1.z2.z2.c ),
    .B(_1982_),
    .Y(_2000_)
);

INVX1 _5414_ (
    .A(\z3.z1.z2.z2.c ),
    .Y(_2001_)
);

NAND2X1 _5415_ (
    .A(_2001_),
    .B(_1972_),
    .Y(_2002_)
);

NAND3X1 _5416_ (
    .A(_1999_),
    .B(_2002_),
    .C(_2000_),
    .Y(_2003_)
);

NAND2X1 _5417_ (
    .A(\z3.z1.z2.z2.c ),
    .B(_1972_),
    .Y(_2004_)
);

NAND2X1 _5418_ (
    .A(_2001_),
    .B(_1982_),
    .Y(_2005_)
);

NAND3X1 _5419_ (
    .A(_1998_),
    .B(_2004_),
    .C(_2005_),
    .Y(_2006_)
);

NAND3X1 _5420_ (
    .A(_1995_),
    .B(_2003_),
    .C(_2006_),
    .Y(_2007_)
);

INVX1 _5421_ (
    .A(_1995_),
    .Y(_2008_)
);

AOI21X1 _5422_ (
    .A(_2005_),
    .B(_2004_),
    .C(_1998_),
    .Y(_2009_)
);

AOI21X1 _5423_ (
    .A(_2000_),
    .B(_2002_),
    .C(_1999_),
    .Y(_2010_)
);

OAI21X1 _5424_ (
    .A(_2009_),
    .B(_2010_),
    .C(_2008_),
    .Y(_2011_)
);

NAND2X1 _5425_ (
    .A(_2007_),
    .B(_2011_),
    .Y(_2012_)
);

NAND2X1 _5426_ (
    .A(_1994_),
    .B(_2012_),
    .Y(_2013_)
);

OR2X2 _5427_ (
    .A(_2012_),
    .B(_1994_),
    .Y(_2014_)
);

NAND2X1 _5428_ (
    .A(_2013_),
    .B(_2014_),
    .Y(\z3.q0 [5])
);

INVX1 _5429_ (
    .A(\z3.z1.z4.z2.s ),
    .Y(_2015_)
);

INVX1 _5430_ (
    .A(_1996_),
    .Y(_2016_)
);

OAI21X1 _5431_ (
    .A(_2016_),
    .B(_2009_),
    .C(_2015_),
    .Y(_2017_)
);

NAND3X1 _5432_ (
    .A(\z3.z1.z4.z2.s ),
    .B(_1996_),
    .C(_2003_),
    .Y(_2018_)
);

NAND2X1 _5433_ (
    .A(_2011_),
    .B(_1994_),
    .Y(_2019_)
);

AOI22X1 _5434_ (
    .A(_2017_),
    .B(_2018_),
    .C(_2019_),
    .D(_2007_),
    .Y(_2020_)
);

NAND2X1 _5435_ (
    .A(_2018_),
    .B(_2017_),
    .Y(_2021_)
);

NAND3X1 _5436_ (
    .A(_1985_),
    .B(_2007_),
    .C(_1989_),
    .Y(_2022_)
);

AOI21X1 _5437_ (
    .A(_2022_),
    .B(_2011_),
    .C(_2021_),
    .Y(_2023_)
);

NOR2X1 _5438_ (
    .A(_2020_),
    .B(_2023_),
    .Y(\z3.q0 [6])
);

OAI21X1 _5439_ (
    .A(_2016_),
    .B(_2009_),
    .C(\z3.z1.z4.z2.s ),
    .Y(_1942_)
);

NAND3X1 _5440_ (
    .A(_2011_),
    .B(_2021_),
    .C(_2022_),
    .Y(_1943_)
);

NAND3X1 _5441_ (
    .A(\z3.z1.z4.z2.c ),
    .B(_1942_),
    .C(_1943_),
    .Y(_1944_)
);

INVX1 _5442_ (
    .A(\z3.z1.z4.z2.c ),
    .Y(_1945_)
);

INVX1 _5443_ (
    .A(_1942_),
    .Y(_1946_)
);

OAI21X1 _5444_ (
    .A(_1946_),
    .B(_2020_),
    .C(_1945_),
    .Y(_1947_)
);

NAND2X1 _5445_ (
    .A(_1944_),
    .B(_1947_),
    .Y(\z3.q0 [7])
);

AOI21X1 _5446_ (
    .A(_1967_),
    .B(_1964_),
    .C(_1953_),
    .Y(_1948_)
);

NOR2X1 _5447_ (
    .A(_1948_),
    .B(_1969_),
    .Y(q2[3])
);

AND2X2 _5448_ (
    .A(b[8]),
    .B(a[0]),
    .Y(q2[0])
);

AND2X2 _5449_ (
    .A(b[8]),
    .B(a[1]),
    .Y(\z3.z1.z1.z1.a )
);

AND2X2 _5450_ (
    .A(a[0]),
    .B(b[9]),
    .Y(\z3.z1.z1.z1.b )
);

AND2X2 _5451_ (
    .A(a[1]),
    .B(b[9]),
    .Y(\z3.z1.z1.z2.a )
);

INVX1 _5452_ (
    .A(\z3.z1.z1.z1.b ),
    .Y(_2024_)
);

NAND2X1 _5453_ (
    .A(\z3.z1.z1.z1.a ),
    .B(_2024_),
    .Y(_2025_)
);

INVX1 _5454_ (
    .A(\z3.z1.z1.z1.a ),
    .Y(_2026_)
);

NAND2X1 _5455_ (
    .A(\z3.z1.z1.z1.b ),
    .B(_2026_),
    .Y(_2027_)
);

NAND2X1 _5456_ (
    .A(_2025_),
    .B(_2027_),
    .Y(\z3.z1.z1.z1.s )
);

NOR2X1 _5457_ (
    .A(_2024_),
    .B(_2026_),
    .Y(\z3.z1.z1.z1.c )
);

INVX1 _5458_ (
    .A(\z3.z1.z1.z1.c ),
    .Y(_2028_)
);

NAND2X1 _5459_ (
    .A(\z3.z1.z1.z2.a ),
    .B(_2028_),
    .Y(_2029_)
);

INVX1 _5460_ (
    .A(\z3.z1.z1.z2.a ),
    .Y(_2030_)
);

NAND2X1 _5461_ (
    .A(\z3.z1.z1.z1.c ),
    .B(_2030_),
    .Y(_2031_)
);

NAND2X1 _5462_ (
    .A(_2029_),
    .B(_2031_),
    .Y(\z3.z1.z1.z2.s )
);

NOR2X1 _5463_ (
    .A(_2028_),
    .B(_2030_),
    .Y(\z3.z1.z1.z2.c )
);

AND2X2 _5464_ (
    .A(b[8]),
    .B(a[2]),
    .Y(\z3.z1.q1 [0])
);

AND2X2 _5465_ (
    .A(b[8]),
    .B(a[3]),
    .Y(\z3.z1.z2.z1.a )
);

AND2X2 _5466_ (
    .A(a[2]),
    .B(b[9]),
    .Y(\z3.z1.z2.z1.b )
);

AND2X2 _5467_ (
    .A(a[3]),
    .B(b[9]),
    .Y(\z3.z1.z2.z2.a )
);

INVX1 _5468_ (
    .A(\z3.z1.z2.z1.b ),
    .Y(_2032_)
);

NAND2X1 _5469_ (
    .A(\z3.z1.z2.z1.a ),
    .B(_2032_),
    .Y(_2033_)
);

INVX1 _5470_ (
    .A(\z3.z1.z2.z1.a ),
    .Y(_2034_)
);

NAND2X1 _5471_ (
    .A(\z3.z1.z2.z1.b ),
    .B(_2034_),
    .Y(_2035_)
);

NAND2X1 _5472_ (
    .A(_2033_),
    .B(_2035_),
    .Y(\z3.z1.z2.z1.s )
);

NOR2X1 _5473_ (
    .A(_2032_),
    .B(_2034_),
    .Y(\z3.z1.z2.z1.c )
);

INVX1 _5474_ (
    .A(\z3.z1.z2.z1.c ),
    .Y(_2036_)
);

NAND2X1 _5475_ (
    .A(\z3.z1.z2.z2.a ),
    .B(_2036_),
    .Y(_2037_)
);

INVX1 _5476_ (
    .A(\z3.z1.z2.z2.a ),
    .Y(_2038_)
);

NAND2X1 _5477_ (
    .A(\z3.z1.z2.z1.c ),
    .B(_2038_),
    .Y(_2039_)
);

NAND2X1 _5478_ (
    .A(_2037_),
    .B(_2039_),
    .Y(\z3.z1.z2.z2.s )
);

NOR2X1 _5479_ (
    .A(_2036_),
    .B(_2038_),
    .Y(\z3.z1.z2.z2.c )
);

AND2X2 _5480_ (
    .A(b[10]),
    .B(a[0]),
    .Y(\z3.z1.q2 [0])
);

AND2X2 _5481_ (
    .A(b[10]),
    .B(a[1]),
    .Y(\z3.z1.z3.z1.a )
);

AND2X2 _5482_ (
    .A(a[0]),
    .B(b[11]),
    .Y(\z3.z1.z3.z1.b )
);

AND2X2 _5483_ (
    .A(a[1]),
    .B(b[11]),
    .Y(\z3.z1.z3.z2.a )
);

INVX1 _5484_ (
    .A(\z3.z1.z3.z1.b ),
    .Y(_2040_)
);

NAND2X1 _5485_ (
    .A(\z3.z1.z3.z1.a ),
    .B(_2040_),
    .Y(_2041_)
);

INVX1 _5486_ (
    .A(\z3.z1.z3.z1.a ),
    .Y(_2042_)
);

NAND2X1 _5487_ (
    .A(\z3.z1.z3.z1.b ),
    .B(_2042_),
    .Y(_2043_)
);

NAND2X1 _5488_ (
    .A(_2041_),
    .B(_2043_),
    .Y(\z3.z1.z3.z1.s )
);

NOR2X1 _5489_ (
    .A(_2040_),
    .B(_2042_),
    .Y(\z3.z1.z3.z1.c )
);

INVX1 _5490_ (
    .A(\z3.z1.z3.z1.c ),
    .Y(_2044_)
);

NAND2X1 _5491_ (
    .A(\z3.z1.z3.z2.a ),
    .B(_2044_),
    .Y(_2045_)
);

INVX1 _5492_ (
    .A(\z3.z1.z3.z2.a ),
    .Y(_2046_)
);

NAND2X1 _5493_ (
    .A(\z3.z1.z3.z1.c ),
    .B(_2046_),
    .Y(_2047_)
);

NAND2X1 _5494_ (
    .A(_2045_),
    .B(_2047_),
    .Y(\z3.z1.z3.z2.s )
);

NOR2X1 _5495_ (
    .A(_2044_),
    .B(_2046_),
    .Y(\z3.z1.z3.z2.c )
);

AND2X2 _5496_ (
    .A(b[10]),
    .B(a[2]),
    .Y(\z3.z1.q3 [0])
);

AND2X2 _5497_ (
    .A(b[10]),
    .B(a[3]),
    .Y(\z3.z1.z4.z1.a )
);

AND2X2 _5498_ (
    .A(a[2]),
    .B(b[11]),
    .Y(\z3.z1.z4.z1.b )
);

AND2X2 _5499_ (
    .A(a[3]),
    .B(b[11]),
    .Y(\z3.z1.z4.z2.a )
);

INVX1 _5500_ (
    .A(\z3.z1.z4.z1.b ),
    .Y(_2048_)
);

NAND2X1 _5501_ (
    .A(\z3.z1.z4.z1.a ),
    .B(_2048_),
    .Y(_2049_)
);

INVX1 _5502_ (
    .A(\z3.z1.z4.z1.a ),
    .Y(_2050_)
);

NAND2X1 _5503_ (
    .A(\z3.z1.z4.z1.b ),
    .B(_2050_),
    .Y(_2051_)
);

NAND2X1 _5504_ (
    .A(_2049_),
    .B(_2051_),
    .Y(\z3.z1.z4.z1.s )
);

NOR2X1 _5505_ (
    .A(_2048_),
    .B(_2050_),
    .Y(\z3.z1.z4.z1.c )
);

INVX1 _5506_ (
    .A(\z3.z1.z4.z1.c ),
    .Y(_2052_)
);

NAND2X1 _5507_ (
    .A(\z3.z1.z4.z2.a ),
    .B(_2052_),
    .Y(_2053_)
);

INVX1 _5508_ (
    .A(\z3.z1.z4.z2.a ),
    .Y(_2054_)
);

NAND2X1 _5509_ (
    .A(\z3.z1.z4.z1.c ),
    .B(_2054_),
    .Y(_2055_)
);

NAND2X1 _5510_ (
    .A(_2053_),
    .B(_2055_),
    .Y(\z3.z1.z4.z2.s )
);

NOR2X1 _5511_ (
    .A(_2052_),
    .B(_2054_),
    .Y(\z3.z1.z4.z2.c )
);

NOR2X1 _5512_ (
    .A(\z3.z2.q1 [0]),
    .B(\z3.z2.z1.z2.s ),
    .Y(_2063_)
);

AND2X2 _5513_ (
    .A(\z3.z2.q1 [0]),
    .B(\z3.z2.z1.z2.s ),
    .Y(_2064_)
);

NOR2X1 _5514_ (
    .A(_2063_),
    .B(_2064_),
    .Y(_2065_)
);

NAND2X1 _5515_ (
    .A(\z3.z2.q2 [0]),
    .B(_2065_),
    .Y(_2066_)
);

INVX1 _5516_ (
    .A(_2066_),
    .Y(_2067_)
);

NOR2X1 _5517_ (
    .A(\z3.z2.q2 [0]),
    .B(_2065_),
    .Y(_2068_)
);

NOR2X1 _5518_ (
    .A(_2068_),
    .B(_2067_),
    .Y(\z3.q1 [2])
);

NAND2X1 _5519_ (
    .A(\z3.z2.q1 [0]),
    .B(\z3.z2.z1.z2.s ),
    .Y(_2069_)
);

NOR2X1 _5520_ (
    .A(\z3.z2.z2.z1.s ),
    .B(\z3.z2.z1.z2.c ),
    .Y(_2070_)
);

NAND2X1 _5521_ (
    .A(\z3.z2.z2.z1.s ),
    .B(\z3.z2.z1.z2.c ),
    .Y(_2071_)
);

INVX1 _5522_ (
    .A(_2071_),
    .Y(_2072_)
);

OAI21X1 _5523_ (
    .A(_2070_),
    .B(_2072_),
    .C(_2069_),
    .Y(_2073_)
);

INVX1 _5524_ (
    .A(\z3.z2.z2.z1.s ),
    .Y(_2074_)
);

INVX1 _5525_ (
    .A(\z3.z2.z1.z2.c ),
    .Y(_2075_)
);

NAND2X1 _5526_ (
    .A(_2074_),
    .B(_2075_),
    .Y(_2076_)
);

NAND3X1 _5527_ (
    .A(_2064_),
    .B(_2071_),
    .C(_2076_),
    .Y(_2077_)
);

NAND3X1 _5528_ (
    .A(\z3.z2.z3.z1.s ),
    .B(_2077_),
    .C(_2073_),
    .Y(_2078_)
);

INVX1 _5529_ (
    .A(\z3.z2.z3.z1.s ),
    .Y(_2079_)
);

NAND2X1 _5530_ (
    .A(_2077_),
    .B(_2073_),
    .Y(_2080_)
);

NAND2X1 _5531_ (
    .A(_2079_),
    .B(_2080_),
    .Y(_2081_)
);

NAND3X1 _5532_ (
    .A(_2067_),
    .B(_2078_),
    .C(_2081_),
    .Y(_2082_)
);

INVX1 _5533_ (
    .A(_2082_),
    .Y(_2083_)
);

INVX1 _5534_ (
    .A(_2078_),
    .Y(_2084_)
);

OAI21X1 _5535_ (
    .A(_2069_),
    .B(_2070_),
    .C(_2071_),
    .Y(_2085_)
);

NAND2X1 _5536_ (
    .A(\z3.z2.z2.z2.s ),
    .B(_2085_),
    .Y(_2086_)
);

INVX1 _5537_ (
    .A(\z3.z2.z2.z2.s ),
    .Y(_2087_)
);

NAND3X1 _5538_ (
    .A(_2087_),
    .B(_2071_),
    .C(_2077_),
    .Y(_2088_)
);

NAND2X1 _5539_ (
    .A(\z3.z2.q3 [0]),
    .B(\z3.z2.z3.z2.s ),
    .Y(_2089_)
);

INVX1 _5540_ (
    .A(\z3.z2.q3 [0]),
    .Y(_2090_)
);

INVX1 _5541_ (
    .A(\z3.z2.z3.z2.s ),
    .Y(_2091_)
);

NAND2X1 _5542_ (
    .A(_2090_),
    .B(_2091_),
    .Y(_2092_)
);

NAND2X1 _5543_ (
    .A(_2089_),
    .B(_2092_),
    .Y(_2093_)
);

INVX1 _5544_ (
    .A(_2093_),
    .Y(_2094_)
);

NAND3X1 _5545_ (
    .A(_2086_),
    .B(_2094_),
    .C(_2088_),
    .Y(_2095_)
);

AND2X2 _5546_ (
    .A(_2085_),
    .B(\z3.z2.z2.z2.s ),
    .Y(_2096_)
);

NOR2X1 _5547_ (
    .A(\z3.z2.z2.z2.s ),
    .B(_2085_),
    .Y(_2097_)
);

OAI21X1 _5548_ (
    .A(_2097_),
    .B(_2096_),
    .C(_2093_),
    .Y(_2098_)
);

NAND3X1 _5549_ (
    .A(_2084_),
    .B(_2095_),
    .C(_2098_),
    .Y(_2099_)
);

INVX1 _5550_ (
    .A(_2095_),
    .Y(_2100_)
);

AOI21X1 _5551_ (
    .A(_2088_),
    .B(_2086_),
    .C(_2094_),
    .Y(_2101_)
);

OAI21X1 _5552_ (
    .A(_2101_),
    .B(_2100_),
    .C(_2078_),
    .Y(_2102_)
);

NAND3X1 _5553_ (
    .A(_2083_),
    .B(_2099_),
    .C(_2102_),
    .Y(_2103_)
);

INVX1 _5554_ (
    .A(_2099_),
    .Y(_2104_)
);

INVX1 _5555_ (
    .A(_2080_),
    .Y(_2105_)
);

AOI22X1 _5556_ (
    .A(\z3.z2.z3.z1.s ),
    .B(_2105_),
    .C(_2098_),
    .D(_2095_),
    .Y(_2106_)
);

OAI21X1 _5557_ (
    .A(_2106_),
    .B(_2104_),
    .C(_2082_),
    .Y(_2107_)
);

AND2X2 _5558_ (
    .A(_2107_),
    .B(_2103_),
    .Y(\z3.q1 [4])
);

OAI21X1 _5559_ (
    .A(_2082_),
    .B(_2106_),
    .C(_2099_),
    .Y(_2108_)
);

OAI21X1 _5560_ (
    .A(_2090_),
    .B(_2091_),
    .C(_2095_),
    .Y(_2109_)
);

NAND2X1 _5561_ (
    .A(\z3.z2.z4.z1.s ),
    .B(\z3.z2.z3.z2.c ),
    .Y(_2110_)
);

OR2X2 _5562_ (
    .A(\z3.z2.z4.z1.s ),
    .B(\z3.z2.z3.z2.c ),
    .Y(_2111_)
);

NAND2X1 _5563_ (
    .A(_2110_),
    .B(_2111_),
    .Y(_2112_)
);

INVX1 _5564_ (
    .A(_2112_),
    .Y(_2113_)
);

NAND2X1 _5565_ (
    .A(\z3.z2.z2.z2.c ),
    .B(_2096_),
    .Y(_2114_)
);

INVX1 _5566_ (
    .A(\z3.z2.z2.z2.c ),
    .Y(_2115_)
);

NAND2X1 _5567_ (
    .A(_2115_),
    .B(_2086_),
    .Y(_2116_)
);

NAND3X1 _5568_ (
    .A(_2113_),
    .B(_2116_),
    .C(_2114_),
    .Y(_2117_)
);

NAND2X1 _5569_ (
    .A(\z3.z2.z2.z2.c ),
    .B(_2086_),
    .Y(_2118_)
);

NAND2X1 _5570_ (
    .A(_2115_),
    .B(_2096_),
    .Y(_2119_)
);

NAND3X1 _5571_ (
    .A(_2112_),
    .B(_2118_),
    .C(_2119_),
    .Y(_2120_)
);

NAND3X1 _5572_ (
    .A(_2109_),
    .B(_2117_),
    .C(_2120_),
    .Y(_2121_)
);

INVX1 _5573_ (
    .A(_2109_),
    .Y(_2122_)
);

AOI21X1 _5574_ (
    .A(_2119_),
    .B(_2118_),
    .C(_2112_),
    .Y(_2123_)
);

AOI21X1 _5575_ (
    .A(_2114_),
    .B(_2116_),
    .C(_2113_),
    .Y(_2124_)
);

OAI21X1 _5576_ (
    .A(_2123_),
    .B(_2124_),
    .C(_2122_),
    .Y(_2125_)
);

NAND2X1 _5577_ (
    .A(_2121_),
    .B(_2125_),
    .Y(_2126_)
);

NAND2X1 _5578_ (
    .A(_2108_),
    .B(_2126_),
    .Y(_2127_)
);

OR2X2 _5579_ (
    .A(_2126_),
    .B(_2108_),
    .Y(_2128_)
);

NAND2X1 _5580_ (
    .A(_2127_),
    .B(_2128_),
    .Y(\z3.q1 [5])
);

INVX1 _5581_ (
    .A(\z3.z2.z4.z2.s ),
    .Y(_2129_)
);

INVX1 _5582_ (
    .A(_2110_),
    .Y(_2130_)
);

OAI21X1 _5583_ (
    .A(_2130_),
    .B(_2123_),
    .C(_2129_),
    .Y(_2131_)
);

NAND3X1 _5584_ (
    .A(\z3.z2.z4.z2.s ),
    .B(_2110_),
    .C(_2117_),
    .Y(_2132_)
);

NAND2X1 _5585_ (
    .A(_2125_),
    .B(_2108_),
    .Y(_2133_)
);

AOI22X1 _5586_ (
    .A(_2131_),
    .B(_2132_),
    .C(_2133_),
    .D(_2121_),
    .Y(_2134_)
);

NAND2X1 _5587_ (
    .A(_2132_),
    .B(_2131_),
    .Y(_2135_)
);

NAND3X1 _5588_ (
    .A(_2099_),
    .B(_2121_),
    .C(_2103_),
    .Y(_2136_)
);

AOI21X1 _5589_ (
    .A(_2136_),
    .B(_2125_),
    .C(_2135_),
    .Y(_2137_)
);

NOR2X1 _5590_ (
    .A(_2134_),
    .B(_2137_),
    .Y(\z3.q1 [6])
);

OAI21X1 _5591_ (
    .A(_2130_),
    .B(_2123_),
    .C(\z3.z2.z4.z2.s ),
    .Y(_2056_)
);

NAND3X1 _5592_ (
    .A(_2125_),
    .B(_2135_),
    .C(_2136_),
    .Y(_2057_)
);

NAND3X1 _5593_ (
    .A(\z3.z2.z4.z2.c ),
    .B(_2056_),
    .C(_2057_),
    .Y(_2058_)
);

INVX1 _5594_ (
    .A(\z3.z2.z4.z2.c ),
    .Y(_2059_)
);

INVX1 _5595_ (
    .A(_2056_),
    .Y(_2060_)
);

OAI21X1 _5596_ (
    .A(_2060_),
    .B(_2134_),
    .C(_2059_),
    .Y(_2061_)
);

NAND2X1 _5597_ (
    .A(_2058_),
    .B(_2061_),
    .Y(\z3.q1 [7])
);

AOI21X1 _5598_ (
    .A(_2081_),
    .B(_2078_),
    .C(_2067_),
    .Y(_2062_)
);

NOR2X1 _5599_ (
    .A(_2062_),
    .B(_2083_),
    .Y(\z3.q1 [3])
);

AND2X2 _5600_ (
    .A(b[8]),
    .B(a[4]),
    .Y(\z3.q1 [0])
);

AND2X2 _5601_ (
    .A(b[8]),
    .B(a[5]),
    .Y(\z3.z2.z1.z1.a )
);

AND2X2 _5602_ (
    .A(a[4]),
    .B(b[9]),
    .Y(\z3.z2.z1.z1.b )
);

AND2X2 _5603_ (
    .A(a[5]),
    .B(b[9]),
    .Y(\z3.z2.z1.z2.a )
);

INVX1 _5604_ (
    .A(\z3.z2.z1.z1.b ),
    .Y(_2138_)
);

NAND2X1 _5605_ (
    .A(\z3.z2.z1.z1.a ),
    .B(_2138_),
    .Y(_2139_)
);

INVX1 _5606_ (
    .A(\z3.z2.z1.z1.a ),
    .Y(_2140_)
);

NAND2X1 _5607_ (
    .A(\z3.z2.z1.z1.b ),
    .B(_2140_),
    .Y(_2141_)
);

NAND2X1 _5608_ (
    .A(_2139_),
    .B(_2141_),
    .Y(\z3.z2.z1.z1.s )
);

NOR2X1 _5609_ (
    .A(_2138_),
    .B(_2140_),
    .Y(\z3.z2.z1.z1.c )
);

INVX1 _5610_ (
    .A(\z3.z2.z1.z1.c ),
    .Y(_2142_)
);

NAND2X1 _5611_ (
    .A(\z3.z2.z1.z2.a ),
    .B(_2142_),
    .Y(_2143_)
);

INVX1 _5612_ (
    .A(\z3.z2.z1.z2.a ),
    .Y(_2144_)
);

NAND2X1 _5613_ (
    .A(\z3.z2.z1.z1.c ),
    .B(_2144_),
    .Y(_2145_)
);

NAND2X1 _5614_ (
    .A(_2143_),
    .B(_2145_),
    .Y(\z3.z2.z1.z2.s )
);

NOR2X1 _5615_ (
    .A(_2142_),
    .B(_2144_),
    .Y(\z3.z2.z1.z2.c )
);

AND2X2 _5616_ (
    .A(b[8]),
    .B(a[6]),
    .Y(\z3.z2.q1 [0])
);

AND2X2 _5617_ (
    .A(b[8]),
    .B(a[7]),
    .Y(\z3.z2.z2.z1.a )
);

AND2X2 _5618_ (
    .A(a[6]),
    .B(b[9]),
    .Y(\z3.z2.z2.z1.b )
);

AND2X2 _5619_ (
    .A(a[7]),
    .B(b[9]),
    .Y(\z3.z2.z2.z2.a )
);

INVX1 _5620_ (
    .A(\z3.z2.z2.z1.b ),
    .Y(_2146_)
);

NAND2X1 _5621_ (
    .A(\z3.z2.z2.z1.a ),
    .B(_2146_),
    .Y(_2147_)
);

INVX1 _5622_ (
    .A(\z3.z2.z2.z1.a ),
    .Y(_2148_)
);

NAND2X1 _5623_ (
    .A(\z3.z2.z2.z1.b ),
    .B(_2148_),
    .Y(_2149_)
);

NAND2X1 _5624_ (
    .A(_2147_),
    .B(_2149_),
    .Y(\z3.z2.z2.z1.s )
);

NOR2X1 _5625_ (
    .A(_2146_),
    .B(_2148_),
    .Y(\z3.z2.z2.z1.c )
);

INVX1 _5626_ (
    .A(\z3.z2.z2.z1.c ),
    .Y(_2150_)
);

NAND2X1 _5627_ (
    .A(\z3.z2.z2.z2.a ),
    .B(_2150_),
    .Y(_2151_)
);

INVX1 _5628_ (
    .A(\z3.z2.z2.z2.a ),
    .Y(_2152_)
);

NAND2X1 _5629_ (
    .A(\z3.z2.z2.z1.c ),
    .B(_2152_),
    .Y(_2153_)
);

NAND2X1 _5630_ (
    .A(_2151_),
    .B(_2153_),
    .Y(\z3.z2.z2.z2.s )
);

NOR2X1 _5631_ (
    .A(_2150_),
    .B(_2152_),
    .Y(\z3.z2.z2.z2.c )
);

AND2X2 _5632_ (
    .A(b[10]),
    .B(a[4]),
    .Y(\z3.z2.q2 [0])
);

AND2X2 _5633_ (
    .A(b[10]),
    .B(a[5]),
    .Y(\z3.z2.z3.z1.a )
);

AND2X2 _5634_ (
    .A(a[4]),
    .B(b[11]),
    .Y(\z3.z2.z3.z1.b )
);

AND2X2 _5635_ (
    .A(a[5]),
    .B(b[11]),
    .Y(\z3.z2.z3.z2.a )
);

INVX1 _5636_ (
    .A(\z3.z2.z3.z1.b ),
    .Y(_2154_)
);

NAND2X1 _5637_ (
    .A(\z3.z2.z3.z1.a ),
    .B(_2154_),
    .Y(_2155_)
);

INVX1 _5638_ (
    .A(\z3.z2.z3.z1.a ),
    .Y(_2156_)
);

NAND2X1 _5639_ (
    .A(\z3.z2.z3.z1.b ),
    .B(_2156_),
    .Y(_2157_)
);

NAND2X1 _5640_ (
    .A(_2155_),
    .B(_2157_),
    .Y(\z3.z2.z3.z1.s )
);

NOR2X1 _5641_ (
    .A(_2154_),
    .B(_2156_),
    .Y(\z3.z2.z3.z1.c )
);

INVX1 _5642_ (
    .A(\z3.z2.z3.z1.c ),
    .Y(_2158_)
);

NAND2X1 _5643_ (
    .A(\z3.z2.z3.z2.a ),
    .B(_2158_),
    .Y(_2159_)
);

INVX1 _5644_ (
    .A(\z3.z2.z3.z2.a ),
    .Y(_2160_)
);

NAND2X1 _5645_ (
    .A(\z3.z2.z3.z1.c ),
    .B(_2160_),
    .Y(_2161_)
);

NAND2X1 _5646_ (
    .A(_2159_),
    .B(_2161_),
    .Y(\z3.z2.z3.z2.s )
);

NOR2X1 _5647_ (
    .A(_2158_),
    .B(_2160_),
    .Y(\z3.z2.z3.z2.c )
);

AND2X2 _5648_ (
    .A(b[10]),
    .B(a[6]),
    .Y(\z3.z2.q3 [0])
);

AND2X2 _5649_ (
    .A(b[10]),
    .B(a[7]),
    .Y(\z3.z2.z4.z1.a )
);

AND2X2 _5650_ (
    .A(a[6]),
    .B(b[11]),
    .Y(\z3.z2.z4.z1.b )
);

AND2X2 _5651_ (
    .A(a[7]),
    .B(b[11]),
    .Y(\z3.z2.z4.z2.a )
);

INVX1 _5652_ (
    .A(\z3.z2.z4.z1.b ),
    .Y(_2162_)
);

NAND2X1 _5653_ (
    .A(\z3.z2.z4.z1.a ),
    .B(_2162_),
    .Y(_2163_)
);

INVX1 _5654_ (
    .A(\z3.z2.z4.z1.a ),
    .Y(_2164_)
);

NAND2X1 _5655_ (
    .A(\z3.z2.z4.z1.b ),
    .B(_2164_),
    .Y(_2165_)
);

NAND2X1 _5656_ (
    .A(_2163_),
    .B(_2165_),
    .Y(\z3.z2.z4.z1.s )
);

NOR2X1 _5657_ (
    .A(_2162_),
    .B(_2164_),
    .Y(\z3.z2.z4.z1.c )
);

INVX1 _5658_ (
    .A(\z3.z2.z4.z1.c ),
    .Y(_2166_)
);

NAND2X1 _5659_ (
    .A(\z3.z2.z4.z2.a ),
    .B(_2166_),
    .Y(_2167_)
);

INVX1 _5660_ (
    .A(\z3.z2.z4.z2.a ),
    .Y(_2168_)
);

NAND2X1 _5661_ (
    .A(\z3.z2.z4.z1.c ),
    .B(_2168_),
    .Y(_2169_)
);

NAND2X1 _5662_ (
    .A(_2167_),
    .B(_2169_),
    .Y(\z3.z2.z4.z2.s )
);

NOR2X1 _5663_ (
    .A(_2166_),
    .B(_2168_),
    .Y(\z3.z2.z4.z2.c )
);

NOR2X1 _5664_ (
    .A(\z3.z3.q1 [0]),
    .B(\z3.z3.z1.z2.s ),
    .Y(_2177_)
);

AND2X2 _5665_ (
    .A(\z3.z3.q1 [0]),
    .B(\z3.z3.z1.z2.s ),
    .Y(_2178_)
);

NOR2X1 _5666_ (
    .A(_2177_),
    .B(_2178_),
    .Y(_2179_)
);

NAND2X1 _5667_ (
    .A(\z3.z3.q2 [0]),
    .B(_2179_),
    .Y(_2180_)
);

INVX1 _5668_ (
    .A(_2180_),
    .Y(_2181_)
);

NOR2X1 _5669_ (
    .A(\z3.z3.q2 [0]),
    .B(_2179_),
    .Y(_2182_)
);

NOR2X1 _5670_ (
    .A(_2182_),
    .B(_2181_),
    .Y(\z3.q2 [2])
);

NAND2X1 _5671_ (
    .A(\z3.z3.q1 [0]),
    .B(\z3.z3.z1.z2.s ),
    .Y(_2183_)
);

NOR2X1 _5672_ (
    .A(\z3.z3.z2.z1.s ),
    .B(\z3.z3.z1.z2.c ),
    .Y(_2184_)
);

NAND2X1 _5673_ (
    .A(\z3.z3.z2.z1.s ),
    .B(\z3.z3.z1.z2.c ),
    .Y(_2185_)
);

INVX1 _5674_ (
    .A(_2185_),
    .Y(_2186_)
);

OAI21X1 _5675_ (
    .A(_2184_),
    .B(_2186_),
    .C(_2183_),
    .Y(_2187_)
);

INVX1 _5676_ (
    .A(\z3.z3.z2.z1.s ),
    .Y(_2188_)
);

INVX1 _5677_ (
    .A(\z3.z3.z1.z2.c ),
    .Y(_2189_)
);

NAND2X1 _5678_ (
    .A(_2188_),
    .B(_2189_),
    .Y(_2190_)
);

NAND3X1 _5679_ (
    .A(_2178_),
    .B(_2185_),
    .C(_2190_),
    .Y(_2191_)
);

NAND3X1 _5680_ (
    .A(\z3.z3.z3.z1.s ),
    .B(_2191_),
    .C(_2187_),
    .Y(_2192_)
);

INVX1 _5681_ (
    .A(\z3.z3.z3.z1.s ),
    .Y(_2193_)
);

NAND2X1 _5682_ (
    .A(_2191_),
    .B(_2187_),
    .Y(_2194_)
);

NAND2X1 _5683_ (
    .A(_2193_),
    .B(_2194_),
    .Y(_2195_)
);

NAND3X1 _5684_ (
    .A(_2181_),
    .B(_2192_),
    .C(_2195_),
    .Y(_2196_)
);

INVX1 _5685_ (
    .A(_2196_),
    .Y(_2197_)
);

INVX1 _5686_ (
    .A(_2192_),
    .Y(_2198_)
);

OAI21X1 _5687_ (
    .A(_2183_),
    .B(_2184_),
    .C(_2185_),
    .Y(_2199_)
);

NAND2X1 _5688_ (
    .A(\z3.z3.z2.z2.s ),
    .B(_2199_),
    .Y(_2200_)
);

INVX1 _5689_ (
    .A(\z3.z3.z2.z2.s ),
    .Y(_2201_)
);

NAND3X1 _5690_ (
    .A(_2201_),
    .B(_2185_),
    .C(_2191_),
    .Y(_2202_)
);

NAND2X1 _5691_ (
    .A(\z3.z3.q3 [0]),
    .B(\z3.z3.z3.z2.s ),
    .Y(_2203_)
);

INVX1 _5692_ (
    .A(\z3.z3.q3 [0]),
    .Y(_2204_)
);

INVX1 _5693_ (
    .A(\z3.z3.z3.z2.s ),
    .Y(_2205_)
);

NAND2X1 _5694_ (
    .A(_2204_),
    .B(_2205_),
    .Y(_2206_)
);

NAND2X1 _5695_ (
    .A(_2203_),
    .B(_2206_),
    .Y(_2207_)
);

INVX1 _5696_ (
    .A(_2207_),
    .Y(_2208_)
);

NAND3X1 _5697_ (
    .A(_2200_),
    .B(_2208_),
    .C(_2202_),
    .Y(_2209_)
);

AND2X2 _5698_ (
    .A(_2199_),
    .B(\z3.z3.z2.z2.s ),
    .Y(_2210_)
);

NOR2X1 _5699_ (
    .A(\z3.z3.z2.z2.s ),
    .B(_2199_),
    .Y(_2211_)
);

OAI21X1 _5700_ (
    .A(_2211_),
    .B(_2210_),
    .C(_2207_),
    .Y(_2212_)
);

NAND3X1 _5701_ (
    .A(_2198_),
    .B(_2209_),
    .C(_2212_),
    .Y(_2213_)
);

INVX1 _5702_ (
    .A(_2209_),
    .Y(_2214_)
);

AOI21X1 _5703_ (
    .A(_2202_),
    .B(_2200_),
    .C(_2208_),
    .Y(_2215_)
);

OAI21X1 _5704_ (
    .A(_2215_),
    .B(_2214_),
    .C(_2192_),
    .Y(_2216_)
);

NAND3X1 _5705_ (
    .A(_2197_),
    .B(_2213_),
    .C(_2216_),
    .Y(_2217_)
);

INVX1 _5706_ (
    .A(_2213_),
    .Y(_2218_)
);

INVX1 _5707_ (
    .A(_2194_),
    .Y(_2219_)
);

AOI22X1 _5708_ (
    .A(\z3.z3.z3.z1.s ),
    .B(_2219_),
    .C(_2212_),
    .D(_2209_),
    .Y(_2220_)
);

OAI21X1 _5709_ (
    .A(_2220_),
    .B(_2218_),
    .C(_2196_),
    .Y(_2221_)
);

AND2X2 _5710_ (
    .A(_2221_),
    .B(_2217_),
    .Y(\z3.q2 [4])
);

OAI21X1 _5711_ (
    .A(_2196_),
    .B(_2220_),
    .C(_2213_),
    .Y(_2222_)
);

OAI21X1 _5712_ (
    .A(_2204_),
    .B(_2205_),
    .C(_2209_),
    .Y(_2223_)
);

NAND2X1 _5713_ (
    .A(\z3.z3.z4.z1.s ),
    .B(\z3.z3.z3.z2.c ),
    .Y(_2224_)
);

OR2X2 _5714_ (
    .A(\z3.z3.z4.z1.s ),
    .B(\z3.z3.z3.z2.c ),
    .Y(_2225_)
);

NAND2X1 _5715_ (
    .A(_2224_),
    .B(_2225_),
    .Y(_2226_)
);

INVX1 _5716_ (
    .A(_2226_),
    .Y(_2227_)
);

NAND2X1 _5717_ (
    .A(\z3.z3.z2.z2.c ),
    .B(_2210_),
    .Y(_2228_)
);

INVX1 _5718_ (
    .A(\z3.z3.z2.z2.c ),
    .Y(_2229_)
);

NAND2X1 _5719_ (
    .A(_2229_),
    .B(_2200_),
    .Y(_2230_)
);

NAND3X1 _5720_ (
    .A(_2227_),
    .B(_2230_),
    .C(_2228_),
    .Y(_2231_)
);

NAND2X1 _5721_ (
    .A(\z3.z3.z2.z2.c ),
    .B(_2200_),
    .Y(_2232_)
);

NAND2X1 _5722_ (
    .A(_2229_),
    .B(_2210_),
    .Y(_2233_)
);

NAND3X1 _5723_ (
    .A(_2226_),
    .B(_2232_),
    .C(_2233_),
    .Y(_2234_)
);

NAND3X1 _5724_ (
    .A(_2223_),
    .B(_2231_),
    .C(_2234_),
    .Y(_2235_)
);

INVX1 _5725_ (
    .A(_2223_),
    .Y(_2236_)
);

AOI21X1 _5726_ (
    .A(_2233_),
    .B(_2232_),
    .C(_2226_),
    .Y(_2237_)
);

AOI21X1 _5727_ (
    .A(_2228_),
    .B(_2230_),
    .C(_2227_),
    .Y(_2238_)
);

OAI21X1 _5728_ (
    .A(_2237_),
    .B(_2238_),
    .C(_2236_),
    .Y(_2239_)
);

NAND2X1 _5729_ (
    .A(_2235_),
    .B(_2239_),
    .Y(_2240_)
);

NAND2X1 _5730_ (
    .A(_2222_),
    .B(_2240_),
    .Y(_2241_)
);

OR2X2 _5731_ (
    .A(_2240_),
    .B(_2222_),
    .Y(_2242_)
);

NAND2X1 _5732_ (
    .A(_2241_),
    .B(_2242_),
    .Y(\z3.q2 [5])
);

INVX1 _5733_ (
    .A(\z3.z3.z4.z2.s ),
    .Y(_2243_)
);

INVX1 _5734_ (
    .A(_2224_),
    .Y(_2244_)
);

OAI21X1 _5735_ (
    .A(_2244_),
    .B(_2237_),
    .C(_2243_),
    .Y(_2245_)
);

NAND3X1 _5736_ (
    .A(\z3.z3.z4.z2.s ),
    .B(_2224_),
    .C(_2231_),
    .Y(_2246_)
);

NAND2X1 _5737_ (
    .A(_2239_),
    .B(_2222_),
    .Y(_2247_)
);

AOI22X1 _5738_ (
    .A(_2245_),
    .B(_2246_),
    .C(_2247_),
    .D(_2235_),
    .Y(_2248_)
);

NAND2X1 _5739_ (
    .A(_2246_),
    .B(_2245_),
    .Y(_2249_)
);

NAND3X1 _5740_ (
    .A(_2213_),
    .B(_2235_),
    .C(_2217_),
    .Y(_2250_)
);

AOI21X1 _5741_ (
    .A(_2250_),
    .B(_2239_),
    .C(_2249_),
    .Y(_2251_)
);

NOR2X1 _5742_ (
    .A(_2248_),
    .B(_2251_),
    .Y(\z3.q2 [6])
);

OAI21X1 _5743_ (
    .A(_2244_),
    .B(_2237_),
    .C(\z3.z3.z4.z2.s ),
    .Y(_2170_)
);

NAND3X1 _5744_ (
    .A(_2239_),
    .B(_2249_),
    .C(_2250_),
    .Y(_2171_)
);

NAND3X1 _5745_ (
    .A(\z3.z3.z4.z2.c ),
    .B(_2170_),
    .C(_2171_),
    .Y(_2172_)
);

INVX1 _5746_ (
    .A(\z3.z3.z4.z2.c ),
    .Y(_2173_)
);

INVX1 _5747_ (
    .A(_2170_),
    .Y(_2174_)
);

OAI21X1 _5748_ (
    .A(_2174_),
    .B(_2248_),
    .C(_2173_),
    .Y(_2175_)
);

NAND2X1 _5749_ (
    .A(_2172_),
    .B(_2175_),
    .Y(\z3.q2 [7])
);

AOI21X1 _5750_ (
    .A(_2195_),
    .B(_2192_),
    .C(_2181_),
    .Y(_2176_)
);

NOR2X1 _5751_ (
    .A(_2176_),
    .B(_2197_),
    .Y(\z3.q2 [3])
);

AND2X2 _5752_ (
    .A(b[12]),
    .B(a[0]),
    .Y(\z3.q2 [0])
);

AND2X2 _5753_ (
    .A(b[12]),
    .B(a[1]),
    .Y(\z3.z3.z1.z1.a )
);

AND2X2 _5754_ (
    .A(a[0]),
    .B(b[13]),
    .Y(\z3.z3.z1.z1.b )
);

AND2X2 _5755_ (
    .A(a[1]),
    .B(b[13]),
    .Y(\z3.z3.z1.z2.a )
);

INVX1 _5756_ (
    .A(\z3.z3.z1.z1.b ),
    .Y(_2252_)
);

NAND2X1 _5757_ (
    .A(\z3.z3.z1.z1.a ),
    .B(_2252_),
    .Y(_2253_)
);

INVX1 _5758_ (
    .A(\z3.z3.z1.z1.a ),
    .Y(_2254_)
);

NAND2X1 _5759_ (
    .A(\z3.z3.z1.z1.b ),
    .B(_2254_),
    .Y(_2255_)
);

NAND2X1 _5760_ (
    .A(_2253_),
    .B(_2255_),
    .Y(\z3.z3.z1.z1.s )
);

NOR2X1 _5761_ (
    .A(_2252_),
    .B(_2254_),
    .Y(\z3.z3.z1.z1.c )
);

INVX1 _5762_ (
    .A(\z3.z3.z1.z1.c ),
    .Y(_2256_)
);

NAND2X1 _5763_ (
    .A(\z3.z3.z1.z2.a ),
    .B(_2256_),
    .Y(_2257_)
);

INVX1 _5764_ (
    .A(\z3.z3.z1.z2.a ),
    .Y(_2258_)
);

NAND2X1 _5765_ (
    .A(\z3.z3.z1.z1.c ),
    .B(_2258_),
    .Y(_2259_)
);

NAND2X1 _5766_ (
    .A(_2257_),
    .B(_2259_),
    .Y(\z3.z3.z1.z2.s )
);

NOR2X1 _5767_ (
    .A(_2256_),
    .B(_2258_),
    .Y(\z3.z3.z1.z2.c )
);

AND2X2 _5768_ (
    .A(b[12]),
    .B(a[2]),
    .Y(\z3.z3.q1 [0])
);

AND2X2 _5769_ (
    .A(b[12]),
    .B(a[3]),
    .Y(\z3.z3.z2.z1.a )
);

AND2X2 _5770_ (
    .A(a[2]),
    .B(b[13]),
    .Y(\z3.z3.z2.z1.b )
);

AND2X2 _5771_ (
    .A(a[3]),
    .B(b[13]),
    .Y(\z3.z3.z2.z2.a )
);

INVX1 _5772_ (
    .A(\z3.z3.z2.z1.b ),
    .Y(_2260_)
);

NAND2X1 _5773_ (
    .A(\z3.z3.z2.z1.a ),
    .B(_2260_),
    .Y(_2261_)
);

INVX1 _5774_ (
    .A(\z3.z3.z2.z1.a ),
    .Y(_2262_)
);

NAND2X1 _5775_ (
    .A(\z3.z3.z2.z1.b ),
    .B(_2262_),
    .Y(_2263_)
);

NAND2X1 _5776_ (
    .A(_2261_),
    .B(_2263_),
    .Y(\z3.z3.z2.z1.s )
);

NOR2X1 _5777_ (
    .A(_2260_),
    .B(_2262_),
    .Y(\z3.z3.z2.z1.c )
);

INVX1 _5778_ (
    .A(\z3.z3.z2.z1.c ),
    .Y(_2264_)
);

NAND2X1 _5779_ (
    .A(\z3.z3.z2.z2.a ),
    .B(_2264_),
    .Y(_2265_)
);

INVX1 _5780_ (
    .A(\z3.z3.z2.z2.a ),
    .Y(_2266_)
);

NAND2X1 _5781_ (
    .A(\z3.z3.z2.z1.c ),
    .B(_2266_),
    .Y(_2267_)
);

NAND2X1 _5782_ (
    .A(_2265_),
    .B(_2267_),
    .Y(\z3.z3.z2.z2.s )
);

NOR2X1 _5783_ (
    .A(_2264_),
    .B(_2266_),
    .Y(\z3.z3.z2.z2.c )
);

AND2X2 _5784_ (
    .A(b[14]),
    .B(a[0]),
    .Y(\z3.z3.q2 [0])
);

AND2X2 _5785_ (
    .A(b[14]),
    .B(a[1]),
    .Y(\z3.z3.z3.z1.a )
);

AND2X2 _5786_ (
    .A(a[0]),
    .B(b[15]),
    .Y(\z3.z3.z3.z1.b )
);

AND2X2 _5787_ (
    .A(a[1]),
    .B(b[15]),
    .Y(\z3.z3.z3.z2.a )
);

INVX1 _5788_ (
    .A(\z3.z3.z3.z1.b ),
    .Y(_2268_)
);

NAND2X1 _5789_ (
    .A(\z3.z3.z3.z1.a ),
    .B(_2268_),
    .Y(_2269_)
);

INVX1 _5790_ (
    .A(\z3.z3.z3.z1.a ),
    .Y(_2270_)
);

NAND2X1 _5791_ (
    .A(\z3.z3.z3.z1.b ),
    .B(_2270_),
    .Y(_2271_)
);

NAND2X1 _5792_ (
    .A(_2269_),
    .B(_2271_),
    .Y(\z3.z3.z3.z1.s )
);

NOR2X1 _5793_ (
    .A(_2268_),
    .B(_2270_),
    .Y(\z3.z3.z3.z1.c )
);

INVX1 _5794_ (
    .A(\z3.z3.z3.z1.c ),
    .Y(_2272_)
);

NAND2X1 _5795_ (
    .A(\z3.z3.z3.z2.a ),
    .B(_2272_),
    .Y(_2273_)
);

INVX1 _5796_ (
    .A(\z3.z3.z3.z2.a ),
    .Y(_2274_)
);

NAND2X1 _5797_ (
    .A(\z3.z3.z3.z1.c ),
    .B(_2274_),
    .Y(_2275_)
);

NAND2X1 _5798_ (
    .A(_2273_),
    .B(_2275_),
    .Y(\z3.z3.z3.z2.s )
);

NOR2X1 _5799_ (
    .A(_2272_),
    .B(_2274_),
    .Y(\z3.z3.z3.z2.c )
);

AND2X2 _5800_ (
    .A(b[14]),
    .B(a[2]),
    .Y(\z3.z3.q3 [0])
);

AND2X2 _5801_ (
    .A(b[14]),
    .B(a[3]),
    .Y(\z3.z3.z4.z1.a )
);

AND2X2 _5802_ (
    .A(a[2]),
    .B(b[15]),
    .Y(\z3.z3.z4.z1.b )
);

AND2X2 _5803_ (
    .A(a[3]),
    .B(b[15]),
    .Y(\z3.z3.z4.z2.a )
);

INVX1 _5804_ (
    .A(\z3.z3.z4.z1.b ),
    .Y(_2276_)
);

NAND2X1 _5805_ (
    .A(\z3.z3.z4.z1.a ),
    .B(_2276_),
    .Y(_2277_)
);

INVX1 _5806_ (
    .A(\z3.z3.z4.z1.a ),
    .Y(_2278_)
);

NAND2X1 _5807_ (
    .A(\z3.z3.z4.z1.b ),
    .B(_2278_),
    .Y(_2279_)
);

NAND2X1 _5808_ (
    .A(_2277_),
    .B(_2279_),
    .Y(\z3.z3.z4.z1.s )
);

NOR2X1 _5809_ (
    .A(_2276_),
    .B(_2278_),
    .Y(\z3.z3.z4.z1.c )
);

INVX1 _5810_ (
    .A(\z3.z3.z4.z1.c ),
    .Y(_2280_)
);

NAND2X1 _5811_ (
    .A(\z3.z3.z4.z2.a ),
    .B(_2280_),
    .Y(_2281_)
);

INVX1 _5812_ (
    .A(\z3.z3.z4.z2.a ),
    .Y(_2282_)
);

NAND2X1 _5813_ (
    .A(\z3.z3.z4.z1.c ),
    .B(_2282_),
    .Y(_2283_)
);

NAND2X1 _5814_ (
    .A(_2281_),
    .B(_2283_),
    .Y(\z3.z3.z4.z2.s )
);

NOR2X1 _5815_ (
    .A(_2280_),
    .B(_2282_),
    .Y(\z3.z3.z4.z2.c )
);

NOR2X1 _5816_ (
    .A(\z3.z4.q1 [0]),
    .B(\z3.z4.z1.z2.s ),
    .Y(_2291_)
);

AND2X2 _5817_ (
    .A(\z3.z4.q1 [0]),
    .B(\z3.z4.z1.z2.s ),
    .Y(_2292_)
);

NOR2X1 _5818_ (
    .A(_2291_),
    .B(_2292_),
    .Y(_2293_)
);

NAND2X1 _5819_ (
    .A(\z3.z4.q2 [0]),
    .B(_2293_),
    .Y(_2294_)
);

INVX1 _5820_ (
    .A(_2294_),
    .Y(_2295_)
);

NOR2X1 _5821_ (
    .A(\z3.z4.q2 [0]),
    .B(_2293_),
    .Y(_2296_)
);

NOR2X1 _5822_ (
    .A(_2296_),
    .B(_2295_),
    .Y(\z3.q3 [2])
);

NAND2X1 _5823_ (
    .A(\z3.z4.q1 [0]),
    .B(\z3.z4.z1.z2.s ),
    .Y(_2297_)
);

NOR2X1 _5824_ (
    .A(\z3.z4.z2.z1.s ),
    .B(\z3.z4.z1.z2.c ),
    .Y(_2298_)
);

NAND2X1 _5825_ (
    .A(\z3.z4.z2.z1.s ),
    .B(\z3.z4.z1.z2.c ),
    .Y(_2299_)
);

INVX1 _5826_ (
    .A(_2299_),
    .Y(_2300_)
);

OAI21X1 _5827_ (
    .A(_2298_),
    .B(_2300_),
    .C(_2297_),
    .Y(_2301_)
);

INVX1 _5828_ (
    .A(\z3.z4.z2.z1.s ),
    .Y(_2302_)
);

INVX1 _5829_ (
    .A(\z3.z4.z1.z2.c ),
    .Y(_2303_)
);

NAND2X1 _5830_ (
    .A(_2302_),
    .B(_2303_),
    .Y(_2304_)
);

NAND3X1 _5831_ (
    .A(_2292_),
    .B(_2299_),
    .C(_2304_),
    .Y(_2305_)
);

NAND3X1 _5832_ (
    .A(\z3.z4.z3.z1.s ),
    .B(_2305_),
    .C(_2301_),
    .Y(_2306_)
);

INVX1 _5833_ (
    .A(\z3.z4.z3.z1.s ),
    .Y(_2307_)
);

NAND2X1 _5834_ (
    .A(_2305_),
    .B(_2301_),
    .Y(_2308_)
);

NAND2X1 _5835_ (
    .A(_2307_),
    .B(_2308_),
    .Y(_2309_)
);

NAND3X1 _5836_ (
    .A(_2295_),
    .B(_2306_),
    .C(_2309_),
    .Y(_2310_)
);

INVX1 _5837_ (
    .A(_2310_),
    .Y(_2311_)
);

INVX1 _5838_ (
    .A(_2306_),
    .Y(_2312_)
);

OAI21X1 _5839_ (
    .A(_2297_),
    .B(_2298_),
    .C(_2299_),
    .Y(_2313_)
);

NAND2X1 _5840_ (
    .A(\z3.z4.z2.z2.s ),
    .B(_2313_),
    .Y(_2314_)
);

INVX1 _5841_ (
    .A(\z3.z4.z2.z2.s ),
    .Y(_2315_)
);

NAND3X1 _5842_ (
    .A(_2315_),
    .B(_2299_),
    .C(_2305_),
    .Y(_2316_)
);

NAND2X1 _5843_ (
    .A(\z3.z4.q3 [0]),
    .B(\z3.z4.z3.z2.s ),
    .Y(_2317_)
);

INVX1 _5844_ (
    .A(\z3.z4.q3 [0]),
    .Y(_2318_)
);

INVX1 _5845_ (
    .A(\z3.z4.z3.z2.s ),
    .Y(_2319_)
);

NAND2X1 _5846_ (
    .A(_2318_),
    .B(_2319_),
    .Y(_2320_)
);

NAND2X1 _5847_ (
    .A(_2317_),
    .B(_2320_),
    .Y(_2321_)
);

INVX1 _5848_ (
    .A(_2321_),
    .Y(_2322_)
);

NAND3X1 _5849_ (
    .A(_2314_),
    .B(_2322_),
    .C(_2316_),
    .Y(_2323_)
);

AND2X2 _5850_ (
    .A(_2313_),
    .B(\z3.z4.z2.z2.s ),
    .Y(_2324_)
);

NOR2X1 _5851_ (
    .A(\z3.z4.z2.z2.s ),
    .B(_2313_),
    .Y(_2325_)
);

OAI21X1 _5852_ (
    .A(_2325_),
    .B(_2324_),
    .C(_2321_),
    .Y(_2326_)
);

NAND3X1 _5853_ (
    .A(_2312_),
    .B(_2323_),
    .C(_2326_),
    .Y(_2327_)
);

INVX1 _5854_ (
    .A(_2323_),
    .Y(_2328_)
);

AOI21X1 _5855_ (
    .A(_2316_),
    .B(_2314_),
    .C(_2322_),
    .Y(_2329_)
);

OAI21X1 _5856_ (
    .A(_2329_),
    .B(_2328_),
    .C(_2306_),
    .Y(_2330_)
);

NAND3X1 _5857_ (
    .A(_2311_),
    .B(_2327_),
    .C(_2330_),
    .Y(_2331_)
);

INVX1 _5858_ (
    .A(_2327_),
    .Y(_2332_)
);

INVX1 _5859_ (
    .A(_2308_),
    .Y(_2333_)
);

AOI22X1 _5860_ (
    .A(\z3.z4.z3.z1.s ),
    .B(_2333_),
    .C(_2326_),
    .D(_2323_),
    .Y(_2334_)
);

OAI21X1 _5861_ (
    .A(_2334_),
    .B(_2332_),
    .C(_2310_),
    .Y(_2335_)
);

AND2X2 _5862_ (
    .A(_2335_),
    .B(_2331_),
    .Y(\z3.q3 [4])
);

OAI21X1 _5863_ (
    .A(_2310_),
    .B(_2334_),
    .C(_2327_),
    .Y(_2336_)
);

OAI21X1 _5864_ (
    .A(_2318_),
    .B(_2319_),
    .C(_2323_),
    .Y(_2337_)
);

NAND2X1 _5865_ (
    .A(\z3.z4.z4.z1.s ),
    .B(\z3.z4.z3.z2.c ),
    .Y(_2338_)
);

OR2X2 _5866_ (
    .A(\z3.z4.z4.z1.s ),
    .B(\z3.z4.z3.z2.c ),
    .Y(_2339_)
);

NAND2X1 _5867_ (
    .A(_2338_),
    .B(_2339_),
    .Y(_2340_)
);

INVX1 _5868_ (
    .A(_2340_),
    .Y(_2341_)
);

NAND2X1 _5869_ (
    .A(\z3.z4.z2.z2.c ),
    .B(_2324_),
    .Y(_2342_)
);

INVX1 _5870_ (
    .A(\z3.z4.z2.z2.c ),
    .Y(_2343_)
);

NAND2X1 _5871_ (
    .A(_2343_),
    .B(_2314_),
    .Y(_2344_)
);

NAND3X1 _5872_ (
    .A(_2341_),
    .B(_2344_),
    .C(_2342_),
    .Y(_2345_)
);

NAND2X1 _5873_ (
    .A(\z3.z4.z2.z2.c ),
    .B(_2314_),
    .Y(_2346_)
);

NAND2X1 _5874_ (
    .A(_2343_),
    .B(_2324_),
    .Y(_2347_)
);

NAND3X1 _5875_ (
    .A(_2340_),
    .B(_2346_),
    .C(_2347_),
    .Y(_2348_)
);

NAND3X1 _5876_ (
    .A(_2337_),
    .B(_2345_),
    .C(_2348_),
    .Y(_2349_)
);

INVX1 _5877_ (
    .A(_2337_),
    .Y(_2350_)
);

AOI21X1 _5878_ (
    .A(_2347_),
    .B(_2346_),
    .C(_2340_),
    .Y(_2351_)
);

AOI21X1 _5879_ (
    .A(_2342_),
    .B(_2344_),
    .C(_2341_),
    .Y(_2352_)
);

OAI21X1 _5880_ (
    .A(_2351_),
    .B(_2352_),
    .C(_2350_),
    .Y(_2353_)
);

NAND2X1 _5881_ (
    .A(_2349_),
    .B(_2353_),
    .Y(_2354_)
);

NAND2X1 _5882_ (
    .A(_2336_),
    .B(_2354_),
    .Y(_2355_)
);

OR2X2 _5883_ (
    .A(_2354_),
    .B(_2336_),
    .Y(_2356_)
);

NAND2X1 _5884_ (
    .A(_2355_),
    .B(_2356_),
    .Y(\z3.q3 [5])
);

INVX1 _5885_ (
    .A(\z3.z4.z4.z2.s ),
    .Y(_2357_)
);

INVX1 _5886_ (
    .A(_2338_),
    .Y(_2358_)
);

OAI21X1 _5887_ (
    .A(_2358_),
    .B(_2351_),
    .C(_2357_),
    .Y(_2359_)
);

NAND3X1 _5888_ (
    .A(\z3.z4.z4.z2.s ),
    .B(_2338_),
    .C(_2345_),
    .Y(_2360_)
);

NAND2X1 _5889_ (
    .A(_2353_),
    .B(_2336_),
    .Y(_2361_)
);

AOI22X1 _5890_ (
    .A(_2359_),
    .B(_2360_),
    .C(_2361_),
    .D(_2349_),
    .Y(_2362_)
);

NAND2X1 _5891_ (
    .A(_2360_),
    .B(_2359_),
    .Y(_2363_)
);

NAND3X1 _5892_ (
    .A(_2327_),
    .B(_2349_),
    .C(_2331_),
    .Y(_2364_)
);

AOI21X1 _5893_ (
    .A(_2364_),
    .B(_2353_),
    .C(_2363_),
    .Y(_2365_)
);

NOR2X1 _5894_ (
    .A(_2362_),
    .B(_2365_),
    .Y(\z3.q3 [6])
);

OAI21X1 _5895_ (
    .A(_2358_),
    .B(_2351_),
    .C(\z3.z4.z4.z2.s ),
    .Y(_2284_)
);

NAND3X1 _5896_ (
    .A(_2353_),
    .B(_2363_),
    .C(_2364_),
    .Y(_2285_)
);

NAND3X1 _5897_ (
    .A(\z3.z4.z4.z2.c ),
    .B(_2284_),
    .C(_2285_),
    .Y(_2286_)
);

INVX1 _5898_ (
    .A(\z3.z4.z4.z2.c ),
    .Y(_2287_)
);

INVX1 _5899_ (
    .A(_2284_),
    .Y(_2288_)
);

OAI21X1 _5900_ (
    .A(_2288_),
    .B(_2362_),
    .C(_2287_),
    .Y(_2289_)
);

NAND2X1 _5901_ (
    .A(_2286_),
    .B(_2289_),
    .Y(\z3.q3 [7])
);

AOI21X1 _5902_ (
    .A(_2309_),
    .B(_2306_),
    .C(_2295_),
    .Y(_2290_)
);

NOR2X1 _5903_ (
    .A(_2290_),
    .B(_2311_),
    .Y(\z3.q3 [3])
);

AND2X2 _5904_ (
    .A(b[12]),
    .B(a[4]),
    .Y(\z3.q3 [0])
);

AND2X2 _5905_ (
    .A(b[12]),
    .B(a[5]),
    .Y(\z3.z4.z1.z1.a )
);

AND2X2 _5906_ (
    .A(a[4]),
    .B(b[13]),
    .Y(\z3.z4.z1.z1.b )
);

AND2X2 _5907_ (
    .A(a[5]),
    .B(b[13]),
    .Y(\z3.z4.z1.z2.a )
);

INVX1 _5908_ (
    .A(\z3.z4.z1.z1.b ),
    .Y(_2366_)
);

NAND2X1 _5909_ (
    .A(\z3.z4.z1.z1.a ),
    .B(_2366_),
    .Y(_2367_)
);

INVX1 _5910_ (
    .A(\z3.z4.z1.z1.a ),
    .Y(_2368_)
);

NAND2X1 _5911_ (
    .A(\z3.z4.z1.z1.b ),
    .B(_2368_),
    .Y(_2369_)
);

NAND2X1 _5912_ (
    .A(_2367_),
    .B(_2369_),
    .Y(\z3.z4.z1.z1.s )
);

NOR2X1 _5913_ (
    .A(_2366_),
    .B(_2368_),
    .Y(\z3.z4.z1.z1.c )
);

INVX1 _5914_ (
    .A(\z3.z4.z1.z1.c ),
    .Y(_2370_)
);

NAND2X1 _5915_ (
    .A(\z3.z4.z1.z2.a ),
    .B(_2370_),
    .Y(_2371_)
);

INVX1 _5916_ (
    .A(\z3.z4.z1.z2.a ),
    .Y(_2372_)
);

NAND2X1 _5917_ (
    .A(\z3.z4.z1.z1.c ),
    .B(_2372_),
    .Y(_2373_)
);

NAND2X1 _5918_ (
    .A(_2371_),
    .B(_2373_),
    .Y(\z3.z4.z1.z2.s )
);

NOR2X1 _5919_ (
    .A(_2370_),
    .B(_2372_),
    .Y(\z3.z4.z1.z2.c )
);

AND2X2 _5920_ (
    .A(b[12]),
    .B(a[6]),
    .Y(\z3.z4.q1 [0])
);

AND2X2 _5921_ (
    .A(b[12]),
    .B(a[7]),
    .Y(\z3.z4.z2.z1.a )
);

AND2X2 _5922_ (
    .A(a[6]),
    .B(b[13]),
    .Y(\z3.z4.z2.z1.b )
);

AND2X2 _5923_ (
    .A(a[7]),
    .B(b[13]),
    .Y(\z3.z4.z2.z2.a )
);

INVX1 _5924_ (
    .A(\z3.z4.z2.z1.b ),
    .Y(_2374_)
);

NAND2X1 _5925_ (
    .A(\z3.z4.z2.z1.a ),
    .B(_2374_),
    .Y(_2375_)
);

INVX1 _5926_ (
    .A(\z3.z4.z2.z1.a ),
    .Y(_2376_)
);

NAND2X1 _5927_ (
    .A(\z3.z4.z2.z1.b ),
    .B(_2376_),
    .Y(_2377_)
);

NAND2X1 _5928_ (
    .A(_2375_),
    .B(_2377_),
    .Y(\z3.z4.z2.z1.s )
);

NOR2X1 _5929_ (
    .A(_2374_),
    .B(_2376_),
    .Y(\z3.z4.z2.z1.c )
);

INVX1 _5930_ (
    .A(\z3.z4.z2.z1.c ),
    .Y(_2378_)
);

NAND2X1 _5931_ (
    .A(\z3.z4.z2.z2.a ),
    .B(_2378_),
    .Y(_2379_)
);

INVX1 _5932_ (
    .A(\z3.z4.z2.z2.a ),
    .Y(_2380_)
);

NAND2X1 _5933_ (
    .A(\z3.z4.z2.z1.c ),
    .B(_2380_),
    .Y(_2381_)
);

NAND2X1 _5934_ (
    .A(_2379_),
    .B(_2381_),
    .Y(\z3.z4.z2.z2.s )
);

NOR2X1 _5935_ (
    .A(_2378_),
    .B(_2380_),
    .Y(\z3.z4.z2.z2.c )
);

AND2X2 _5936_ (
    .A(b[14]),
    .B(a[4]),
    .Y(\z3.z4.q2 [0])
);

AND2X2 _5937_ (
    .A(b[14]),
    .B(a[5]),
    .Y(\z3.z4.z3.z1.a )
);

AND2X2 _5938_ (
    .A(a[4]),
    .B(b[15]),
    .Y(\z3.z4.z3.z1.b )
);

AND2X2 _5939_ (
    .A(a[5]),
    .B(b[15]),
    .Y(\z3.z4.z3.z2.a )
);

INVX1 _5940_ (
    .A(\z3.z4.z3.z1.b ),
    .Y(_2382_)
);

NAND2X1 _5941_ (
    .A(\z3.z4.z3.z1.a ),
    .B(_2382_),
    .Y(_2383_)
);

INVX1 _5942_ (
    .A(\z3.z4.z3.z1.a ),
    .Y(_2384_)
);

NAND2X1 _5943_ (
    .A(\z3.z4.z3.z1.b ),
    .B(_2384_),
    .Y(_2385_)
);

NAND2X1 _5944_ (
    .A(_2383_),
    .B(_2385_),
    .Y(\z3.z4.z3.z1.s )
);

NOR2X1 _5945_ (
    .A(_2382_),
    .B(_2384_),
    .Y(\z3.z4.z3.z1.c )
);

INVX1 _5946_ (
    .A(\z3.z4.z3.z1.c ),
    .Y(_2386_)
);

NAND2X1 _5947_ (
    .A(\z3.z4.z3.z2.a ),
    .B(_2386_),
    .Y(_2387_)
);

INVX1 _5948_ (
    .A(\z3.z4.z3.z2.a ),
    .Y(_2388_)
);

NAND2X1 _5949_ (
    .A(\z3.z4.z3.z1.c ),
    .B(_2388_),
    .Y(_2389_)
);

NAND2X1 _5950_ (
    .A(_2387_),
    .B(_2389_),
    .Y(\z3.z4.z3.z2.s )
);

NOR2X1 _5951_ (
    .A(_2386_),
    .B(_2388_),
    .Y(\z3.z4.z3.z2.c )
);

AND2X2 _5952_ (
    .A(b[14]),
    .B(a[6]),
    .Y(\z3.z4.q3 [0])
);

AND2X2 _5953_ (
    .A(b[14]),
    .B(a[7]),
    .Y(\z3.z4.z4.z1.a )
);

AND2X2 _5954_ (
    .A(a[6]),
    .B(b[15]),
    .Y(\z3.z4.z4.z1.b )
);

AND2X2 _5955_ (
    .A(a[7]),
    .B(b[15]),
    .Y(\z3.z4.z4.z2.a )
);

INVX1 _5956_ (
    .A(\z3.z4.z4.z1.b ),
    .Y(_2390_)
);

NAND2X1 _5957_ (
    .A(\z3.z4.z4.z1.a ),
    .B(_2390_),
    .Y(_2391_)
);

INVX1 _5958_ (
    .A(\z3.z4.z4.z1.a ),
    .Y(_2392_)
);

NAND2X1 _5959_ (
    .A(\z3.z4.z4.z1.b ),
    .B(_2392_),
    .Y(_2393_)
);

NAND2X1 _5960_ (
    .A(_2391_),
    .B(_2393_),
    .Y(\z3.z4.z4.z1.s )
);

NOR2X1 _5961_ (
    .A(_2390_),
    .B(_2392_),
    .Y(\z3.z4.z4.z1.c )
);

INVX1 _5962_ (
    .A(\z3.z4.z4.z1.c ),
    .Y(_2394_)
);

NAND2X1 _5963_ (
    .A(\z3.z4.z4.z2.a ),
    .B(_2394_),
    .Y(_2395_)
);

INVX1 _5964_ (
    .A(\z3.z4.z4.z2.a ),
    .Y(_2396_)
);

NAND2X1 _5965_ (
    .A(\z3.z4.z4.z1.c ),
    .B(_2396_),
    .Y(_2397_)
);

NAND2X1 _5966_ (
    .A(_2395_),
    .B(_2397_),
    .Y(\z3.z4.z4.z2.s )
);

NOR2X1 _5967_ (
    .A(_2394_),
    .B(_2396_),
    .Y(\z3.z4.z4.z2.c )
);

OR2X2 _5968_ (
    .A(\z4.q1 [0]),
    .B(\z4.q0 [4]),
    .Y(_2540_)
);

NAND2X1 _5969_ (
    .A(\z4.q1 [0]),
    .B(\z4.q0 [4]),
    .Y(_2541_)
);

NAND2X1 _5970_ (
    .A(_2541_),
    .B(_2540_),
    .Y(_2542_)
);

INVX1 _5971_ (
    .A(_2542_),
    .Y(_2543_)
);

AND2X2 _5972_ (
    .A(_2543_),
    .B(\z4.q2 [0]),
    .Y(_2544_)
);

NOR2X1 _5973_ (
    .A(\z4.q2 [0]),
    .B(_2543_),
    .Y(_2545_)
);

NOR2X1 _5974_ (
    .A(_2545_),
    .B(_2544_),
    .Y(q3[4])
);

INVX1 _5975_ (
    .A(\z4.z3.z1.z1.s ),
    .Y(_2546_)
);

INVX1 _5976_ (
    .A(_2541_),
    .Y(_2547_)
);

NAND2X1 _5977_ (
    .A(\z4.z2.z1.z1.s ),
    .B(\z4.q0 [5]),
    .Y(_2548_)
);

OR2X2 _5978_ (
    .A(\z4.z2.z1.z1.s ),
    .B(\z4.q0 [5]),
    .Y(_2549_)
);

NAND3X1 _5979_ (
    .A(_2548_),
    .B(_2549_),
    .C(_2547_),
    .Y(_2550_)
);

AND2X2 _5980_ (
    .A(\z4.z2.z1.z1.s ),
    .B(\z4.q0 [5]),
    .Y(_2551_)
);

NOR2X1 _5981_ (
    .A(\z4.z2.z1.z1.s ),
    .B(\z4.q0 [5]),
    .Y(_2552_)
);

OAI21X1 _5982_ (
    .A(_2552_),
    .B(_2551_),
    .C(_2541_),
    .Y(_2553_)
);

NAND2X1 _5983_ (
    .A(_2553_),
    .B(_2550_),
    .Y(_2554_)
);

OR2X2 _5984_ (
    .A(_2554_),
    .B(_2546_),
    .Y(_2555_)
);

NAND2X1 _5985_ (
    .A(_2546_),
    .B(_2554_),
    .Y(_2556_)
);

AND2X2 _5986_ (
    .A(_2555_),
    .B(_2556_),
    .Y(_2557_)
);

NAND2X1 _5987_ (
    .A(_2544_),
    .B(_2557_),
    .Y(_2558_)
);

INVX1 _5988_ (
    .A(_2555_),
    .Y(_2559_)
);

OAI21X1 _5989_ (
    .A(_2541_),
    .B(_2552_),
    .C(_2548_),
    .Y(_2560_)
);

INVX1 _5990_ (
    .A(\z4.q0 [6]),
    .Y(_2561_)
);

NOR2X1 _5991_ (
    .A(\z4.q1 [2]),
    .B(_2561_),
    .Y(_2562_)
);

INVX1 _5992_ (
    .A(\z4.q1 [2]),
    .Y(_2563_)
);

NOR2X1 _5993_ (
    .A(\z4.q0 [6]),
    .B(_2563_),
    .Y(_2564_)
);

OAI21X1 _5994_ (
    .A(_2562_),
    .B(_2564_),
    .C(_2560_),
    .Y(_2565_)
);

NAND2X1 _5995_ (
    .A(\z4.q0 [6]),
    .B(_2563_),
    .Y(_2566_)
);

NAND2X1 _5996_ (
    .A(\z4.q1 [2]),
    .B(_2561_),
    .Y(_2567_)
);

NAND2X1 _5997_ (
    .A(_2566_),
    .B(_2567_),
    .Y(_2568_)
);

OR2X2 _5998_ (
    .A(_2568_),
    .B(_2560_),
    .Y(_2569_)
);

NAND3X1 _5999_ (
    .A(\z4.q2 [2]),
    .B(_2565_),
    .C(_2569_),
    .Y(_2570_)
);

INVX1 _6000_ (
    .A(\z4.q2 [2]),
    .Y(_2571_)
);

NAND2X1 _6001_ (
    .A(_2565_),
    .B(_2569_),
    .Y(_2572_)
);

NAND2X1 _6002_ (
    .A(_2571_),
    .B(_2572_),
    .Y(_2573_)
);

AOI21X1 _6003_ (
    .A(_2573_),
    .B(_2570_),
    .C(_2559_),
    .Y(_2574_)
);

INVX1 _6004_ (
    .A(_2574_),
    .Y(_2575_)
);

NAND3X1 _6005_ (
    .A(_2570_),
    .B(_2573_),
    .C(_2559_),
    .Y(_2576_)
);

NAND3X1 _6006_ (
    .A(_2558_),
    .B(_2576_),
    .C(_2575_),
    .Y(_2577_)
);

INVX1 _6007_ (
    .A(_2558_),
    .Y(_2578_)
);

INVX1 _6008_ (
    .A(_2576_),
    .Y(_2579_)
);

OAI21X1 _6009_ (
    .A(_2574_),
    .B(_2579_),
    .C(_2578_),
    .Y(_2580_)
);

NAND2X1 _6010_ (
    .A(_2577_),
    .B(_2580_),
    .Y(q3[6])
);

OAI21X1 _6011_ (
    .A(_2574_),
    .B(_2558_),
    .C(_2576_),
    .Y(_2581_)
);

INVX1 _6012_ (
    .A(_2570_),
    .Y(_2582_)
);

INVX1 _6013_ (
    .A(\z4.q2 [3]),
    .Y(_2583_)
);

INVX1 _6014_ (
    .A(\z4.q0 [7]),
    .Y(_2584_)
);

NOR2X1 _6015_ (
    .A(\z4.q1 [3]),
    .B(_2584_),
    .Y(_2585_)
);

INVX1 _6016_ (
    .A(\z4.q1 [3]),
    .Y(_2586_)
);

NOR2X1 _6017_ (
    .A(\z4.q0 [7]),
    .B(_2586_),
    .Y(_2587_)
);

NAND2X1 _6018_ (
    .A(\z4.q1 [2]),
    .B(\z4.q0 [6]),
    .Y(_2588_)
);

INVX1 _6019_ (
    .A(_2588_),
    .Y(_2589_)
);

AOI21X1 _6020_ (
    .A(_2568_),
    .B(_2560_),
    .C(_2589_),
    .Y(_2590_)
);

OAI21X1 _6021_ (
    .A(_2585_),
    .B(_2587_),
    .C(_2590_),
    .Y(_2591_)
);

NAND2X1 _6022_ (
    .A(\z4.q1 [3]),
    .B(\z4.q0 [7]),
    .Y(_2592_)
);

INVX1 _6023_ (
    .A(_2592_),
    .Y(_2593_)
);

NOR2X1 _6024_ (
    .A(\z4.q1 [3]),
    .B(\z4.q0 [7]),
    .Y(_2594_)
);

INVX1 _6025_ (
    .A(_2590_),
    .Y(_2595_)
);

OAI21X1 _6026_ (
    .A(_2593_),
    .B(_2594_),
    .C(_2595_),
    .Y(_2596_)
);

AOI21X1 _6027_ (
    .A(_2596_),
    .B(_2591_),
    .C(_2583_),
    .Y(_2398_)
);

INVX1 _6028_ (
    .A(_2398_),
    .Y(_2399_)
);

NAND3X1 _6029_ (
    .A(_2583_),
    .B(_2591_),
    .C(_2596_),
    .Y(_2400_)
);

AOI21X1 _6030_ (
    .A(_2399_),
    .B(_2400_),
    .C(_2582_),
    .Y(_2401_)
);

NAND3X1 _6031_ (
    .A(_2582_),
    .B(_2400_),
    .C(_2399_),
    .Y(_2402_)
);

INVX1 _6032_ (
    .A(_2402_),
    .Y(_2403_)
);

OAI21X1 _6033_ (
    .A(_2401_),
    .B(_2403_),
    .C(_2581_),
    .Y(_2404_)
);

INVX1 _6034_ (
    .A(_2581_),
    .Y(_2405_)
);

NAND2X1 _6035_ (
    .A(_2400_),
    .B(_2399_),
    .Y(_2406_)
);

OAI21X1 _6036_ (
    .A(_2571_),
    .B(_2572_),
    .C(_2406_),
    .Y(_2407_)
);

NAND3X1 _6037_ (
    .A(_2402_),
    .B(_2405_),
    .C(_2407_),
    .Y(_2408_)
);

NAND2X1 _6038_ (
    .A(_2408_),
    .B(_2404_),
    .Y(q3[7])
);

AOI21X1 _6039_ (
    .A(_2407_),
    .B(_2581_),
    .C(_2403_),
    .Y(_2409_)
);

AOI21X1 _6040_ (
    .A(_2547_),
    .B(_2549_),
    .C(_2551_),
    .Y(_2410_)
);

OAI22X1 _6041_ (
    .A(_2562_),
    .B(_2564_),
    .C(_2585_),
    .D(_2587_),
    .Y(_2411_)
);

OAI21X1 _6042_ (
    .A(_2588_),
    .B(_2594_),
    .C(_2592_),
    .Y(_2412_)
);

INVX1 _6043_ (
    .A(_2412_),
    .Y(_2413_)
);

OAI21X1 _6044_ (
    .A(_2410_),
    .B(_2411_),
    .C(_2413_),
    .Y(_2414_)
);

NAND2X1 _6045_ (
    .A(\z4.q1 [4]),
    .B(_2414_),
    .Y(_2415_)
);

INVX1 _6046_ (
    .A(\z4.q1 [4]),
    .Y(_2416_)
);

NAND2X1 _6047_ (
    .A(\z4.q0 [7]),
    .B(_2586_),
    .Y(_2417_)
);

NAND2X1 _6048_ (
    .A(\z4.q1 [3]),
    .B(_2584_),
    .Y(_2418_)
);

NAND2X1 _6049_ (
    .A(_2417_),
    .B(_2418_),
    .Y(_2419_)
);

NAND3X1 _6050_ (
    .A(_2560_),
    .B(_2568_),
    .C(_2419_),
    .Y(_2420_)
);

NAND3X1 _6051_ (
    .A(_2416_),
    .B(_2413_),
    .C(_2420_),
    .Y(_2421_)
);

NAND2X1 _6052_ (
    .A(\z4.q3 [0]),
    .B(\z4.q2 [4]),
    .Y(_2422_)
);

INVX1 _6053_ (
    .A(\z4.q3 [0]),
    .Y(_2423_)
);

INVX1 _6054_ (
    .A(\z4.q2 [4]),
    .Y(_2424_)
);

NAND2X1 _6055_ (
    .A(_2423_),
    .B(_2424_),
    .Y(_2425_)
);

NAND2X1 _6056_ (
    .A(_2422_),
    .B(_2425_),
    .Y(_2426_)
);

INVX1 _6057_ (
    .A(_2426_),
    .Y(_2427_)
);

NAND3X1 _6058_ (
    .A(_2421_),
    .B(_2427_),
    .C(_2415_),
    .Y(_2428_)
);

AOI21X1 _6059_ (
    .A(_2420_),
    .B(_2413_),
    .C(_2416_),
    .Y(_2429_)
);

INVX1 _6060_ (
    .A(_2421_),
    .Y(_2430_)
);

OAI21X1 _6061_ (
    .A(_2429_),
    .B(_2430_),
    .C(_2426_),
    .Y(_2431_)
);

NAND3X1 _6062_ (
    .A(_2428_),
    .B(_2431_),
    .C(_2398_),
    .Y(_2432_)
);

NAND2X1 _6063_ (
    .A(_2428_),
    .B(_2431_),
    .Y(_2433_)
);

NAND2X1 _6064_ (
    .A(_2433_),
    .B(_2399_),
    .Y(_2434_)
);

AND2X2 _6065_ (
    .A(_2434_),
    .B(_2432_),
    .Y(_2435_)
);

NAND2X1 _6066_ (
    .A(_2435_),
    .B(_2409_),
    .Y(_2436_)
);

OAI21X1 _6067_ (
    .A(_2401_),
    .B(_2405_),
    .C(_2402_),
    .Y(_2437_)
);

NAND2X1 _6068_ (
    .A(_2432_),
    .B(_2434_),
    .Y(_2438_)
);

NAND2X1 _6069_ (
    .A(_2438_),
    .B(_2437_),
    .Y(_2439_)
);

NAND2X1 _6070_ (
    .A(_2436_),
    .B(_2439_),
    .Y(q3[8])
);

OAI21X1 _6071_ (
    .A(_2438_),
    .B(_2409_),
    .C(_2432_),
    .Y(_2440_)
);

OAI21X1 _6072_ (
    .A(_2423_),
    .B(_2424_),
    .C(_2428_),
    .Y(_2441_)
);

NAND3X1 _6073_ (
    .A(\z4.q1 [4]),
    .B(\z4.q1 [5]),
    .C(_2414_),
    .Y(_2442_)
);

INVX1 _6074_ (
    .A(\z4.q1 [5]),
    .Y(_2443_)
);

AOI22X1 _6075_ (
    .A(_2566_),
    .B(_2567_),
    .C(_2417_),
    .D(_2418_),
    .Y(_2444_)
);

AOI21X1 _6076_ (
    .A(_2444_),
    .B(_2560_),
    .C(_2412_),
    .Y(_2445_)
);

OAI21X1 _6077_ (
    .A(_2416_),
    .B(_2445_),
    .C(_2443_),
    .Y(_2446_)
);

INVX1 _6078_ (
    .A(\z4.z4.z1.z1.s ),
    .Y(_2447_)
);

INVX1 _6079_ (
    .A(\z4.q2 [5]),
    .Y(_2448_)
);

NAND2X1 _6080_ (
    .A(_2447_),
    .B(_2448_),
    .Y(_2449_)
);

NAND2X1 _6081_ (
    .A(\z4.z4.z1.z1.s ),
    .B(\z4.q2 [5]),
    .Y(_2450_)
);

AND2X2 _6082_ (
    .A(_2449_),
    .B(_2450_),
    .Y(_2451_)
);

NAND3X1 _6083_ (
    .A(_2451_),
    .B(_2446_),
    .C(_2442_),
    .Y(_2452_)
);

AOI21X1 _6084_ (
    .A(_2442_),
    .B(_2446_),
    .C(_2451_),
    .Y(_2453_)
);

INVX1 _6085_ (
    .A(_2453_),
    .Y(_2454_)
);

NAND3X1 _6086_ (
    .A(_2452_),
    .B(_2441_),
    .C(_2454_),
    .Y(_2455_)
);

AND2X2 _6087_ (
    .A(_2428_),
    .B(_2422_),
    .Y(_2456_)
);

INVX1 _6088_ (
    .A(_2452_),
    .Y(_2457_)
);

OAI21X1 _6089_ (
    .A(_2457_),
    .B(_2453_),
    .C(_2456_),
    .Y(_2458_)
);

NAND2X1 _6090_ (
    .A(_2455_),
    .B(_2458_),
    .Y(_2459_)
);

OR2X2 _6091_ (
    .A(_2440_),
    .B(_2459_),
    .Y(_2460_)
);

NAND2X1 _6092_ (
    .A(_2459_),
    .B(_2440_),
    .Y(_2461_)
);

NAND2X1 _6093_ (
    .A(_2461_),
    .B(_2460_),
    .Y(q3[9])
);

NAND3X1 _6094_ (
    .A(_2455_),
    .B(_2458_),
    .C(_2435_),
    .Y(_2462_)
);

OAI21X1 _6095_ (
    .A(_2399_),
    .B(_2433_),
    .C(_2455_),
    .Y(_2463_)
);

NAND2X1 _6096_ (
    .A(_2458_),
    .B(_2463_),
    .Y(_2464_)
);

OAI21X1 _6097_ (
    .A(_2409_),
    .B(_2462_),
    .C(_2464_),
    .Y(_2465_)
);

OAI21X1 _6098_ (
    .A(_2447_),
    .B(_2448_),
    .C(_2452_),
    .Y(_2466_)
);

NAND3X1 _6099_ (
    .A(\z4.q1 [5]),
    .B(\z4.q1 [6]),
    .C(_2429_),
    .Y(_2467_)
);

INVX1 _6100_ (
    .A(\z4.q1 [6]),
    .Y(_2468_)
);

NAND2X1 _6101_ (
    .A(_2468_),
    .B(_2442_),
    .Y(_2469_)
);

INVX1 _6102_ (
    .A(\z4.q3 [2]),
    .Y(_2470_)
);

INVX1 _6103_ (
    .A(\z4.q2 [6]),
    .Y(_2471_)
);

NAND2X1 _6104_ (
    .A(_2470_),
    .B(_2471_),
    .Y(_2472_)
);

NAND2X1 _6105_ (
    .A(\z4.q3 [2]),
    .B(\z4.q2 [6]),
    .Y(_2473_)
);

NAND2X1 _6106_ (
    .A(_2473_),
    .B(_2472_),
    .Y(_2474_)
);

INVX1 _6107_ (
    .A(_2474_),
    .Y(_2475_)
);

NAND3X1 _6108_ (
    .A(_2467_),
    .B(_2475_),
    .C(_2469_),
    .Y(_2476_)
);

AOI21X1 _6109_ (
    .A(_2469_),
    .B(_2467_),
    .C(_2475_),
    .Y(_2477_)
);

INVX1 _6110_ (
    .A(_2477_),
    .Y(_2478_)
);

NAND3X1 _6111_ (
    .A(_2466_),
    .B(_2476_),
    .C(_2478_),
    .Y(_2479_)
);

INVX1 _6112_ (
    .A(_2466_),
    .Y(_2480_)
);

INVX1 _6113_ (
    .A(_2476_),
    .Y(_2481_)
);

OAI21X1 _6114_ (
    .A(_2477_),
    .B(_2481_),
    .C(_2480_),
    .Y(_2482_)
);

NAND2X1 _6115_ (
    .A(_2482_),
    .B(_2479_),
    .Y(_2483_)
);

NAND2X1 _6116_ (
    .A(_2483_),
    .B(_2465_),
    .Y(_2484_)
);

NOR2X1 _6117_ (
    .A(_2438_),
    .B(_2459_),
    .Y(_2485_)
);

AOI22X1 _6118_ (
    .A(_2458_),
    .B(_2463_),
    .C(_2485_),
    .D(_2437_),
    .Y(_2486_)
);

AND2X2 _6119_ (
    .A(_2479_),
    .B(_2482_),
    .Y(_2487_)
);

NAND2X1 _6120_ (
    .A(_2487_),
    .B(_2486_),
    .Y(_2488_)
);

NAND2X1 _6121_ (
    .A(_2484_),
    .B(_2488_),
    .Y(q3[10])
);

OAI21X1 _6122_ (
    .A(_2483_),
    .B(_2486_),
    .C(_2479_),
    .Y(_2489_)
);

OAI21X1 _6123_ (
    .A(_2470_),
    .B(_2471_),
    .C(_2476_),
    .Y(_2490_)
);

NOR2X1 _6124_ (
    .A(\z4.q3 [3]),
    .B(\z4.q2 [7]),
    .Y(_2491_)
);

INVX1 _6125_ (
    .A(\z4.q3 [3]),
    .Y(_2492_)
);

INVX1 _6126_ (
    .A(\z4.q2 [7]),
    .Y(_2493_)
);

NOR2X1 _6127_ (
    .A(_2492_),
    .B(_2493_),
    .Y(_2494_)
);

NOR2X1 _6128_ (
    .A(_2491_),
    .B(_2494_),
    .Y(_2495_)
);

INVX1 _6129_ (
    .A(\z4.q1 [7]),
    .Y(_2496_)
);

OAI21X1 _6130_ (
    .A(_2468_),
    .B(_2442_),
    .C(_2496_),
    .Y(_2497_)
);

AND2X2 _6131_ (
    .A(_2429_),
    .B(\z4.q1 [5]),
    .Y(_2498_)
);

NAND3X1 _6132_ (
    .A(\z4.q1 [6]),
    .B(\z4.q1 [7]),
    .C(_2498_),
    .Y(_2499_)
);

NAND3X1 _6133_ (
    .A(_2495_),
    .B(_2497_),
    .C(_2499_),
    .Y(_2500_)
);

INVX1 _6134_ (
    .A(_2495_),
    .Y(_2501_)
);

OAI21X1 _6135_ (
    .A(_2468_),
    .B(_2442_),
    .C(\z4.q1 [7]),
    .Y(_2502_)
);

NAND3X1 _6136_ (
    .A(\z4.q1 [6]),
    .B(_2496_),
    .C(_2498_),
    .Y(_2503_)
);

NAND3X1 _6137_ (
    .A(_2501_),
    .B(_2502_),
    .C(_2503_),
    .Y(_2504_)
);

NAND3X1 _6138_ (
    .A(_2500_),
    .B(_2504_),
    .C(_2490_),
    .Y(_2505_)
);

AND2X2 _6139_ (
    .A(_2476_),
    .B(_2473_),
    .Y(_2506_)
);

NAND2X1 _6140_ (
    .A(_2500_),
    .B(_2504_),
    .Y(_2507_)
);

NAND2X1 _6141_ (
    .A(_2506_),
    .B(_2507_),
    .Y(_2508_)
);

NAND2X1 _6142_ (
    .A(_2505_),
    .B(_2508_),
    .Y(_2509_)
);

OR2X2 _6143_ (
    .A(_2489_),
    .B(_2509_),
    .Y(_2510_)
);

NAND2X1 _6144_ (
    .A(_2509_),
    .B(_2489_),
    .Y(_2511_)
);

NAND2X1 _6145_ (
    .A(_2511_),
    .B(_2510_),
    .Y(q3[11])
);

OAI21X1 _6146_ (
    .A(_2506_),
    .B(_2507_),
    .C(_2479_),
    .Y(_2512_)
);

NAND2X1 _6147_ (
    .A(_2508_),
    .B(_2512_),
    .Y(_2513_)
);

NAND3X1 _6148_ (
    .A(_2505_),
    .B(_2508_),
    .C(_2487_),
    .Y(_2514_)
);

OAI21X1 _6149_ (
    .A(_2514_),
    .B(_2486_),
    .C(_2513_),
    .Y(_2515_)
);

OAI21X1 _6150_ (
    .A(_2492_),
    .B(_2493_),
    .C(_2500_),
    .Y(_2516_)
);

NAND2X1 _6151_ (
    .A(\z4.q3 [4]),
    .B(_2516_),
    .Y(_2517_)
);

OR2X2 _6152_ (
    .A(_2516_),
    .B(\z4.q3 [4]),
    .Y(_2518_)
);

NAND3X1 _6153_ (
    .A(_2517_),
    .B(_2518_),
    .C(_2515_),
    .Y(_2519_)
);

NOR2X1 _6154_ (
    .A(_2483_),
    .B(_2509_),
    .Y(_2520_)
);

AOI22X1 _6155_ (
    .A(_2508_),
    .B(_2512_),
    .C(_2520_),
    .D(_2465_),
    .Y(_2521_)
);

NAND2X1 _6156_ (
    .A(_2517_),
    .B(_2518_),
    .Y(_2522_)
);

NAND2X1 _6157_ (
    .A(_2522_),
    .B(_2521_),
    .Y(_2523_)
);

AND2X2 _6158_ (
    .A(_2519_),
    .B(_2523_),
    .Y(q3[12])
);

INVX1 _6159_ (
    .A(\z4.q3 [5]),
    .Y(_2524_)
);

OAI21X1 _6160_ (
    .A(_2522_),
    .B(_2521_),
    .C(_2517_),
    .Y(_2525_)
);

NAND2X1 _6161_ (
    .A(_2524_),
    .B(_2525_),
    .Y(_2526_)
);

NAND3X1 _6162_ (
    .A(\z4.q3 [5]),
    .B(_2517_),
    .C(_2519_),
    .Y(_2527_)
);

NAND2X1 _6163_ (
    .A(_2527_),
    .B(_2526_),
    .Y(q3[13])
);

INVX1 _6164_ (
    .A(\z4.q3 [6]),
    .Y(_2528_)
);

NAND3X1 _6165_ (
    .A(\z4.q3 [5]),
    .B(_2517_),
    .C(_2518_),
    .Y(_2529_)
);

OAI22X1 _6166_ (
    .A(_2524_),
    .B(_2517_),
    .C(_2529_),
    .D(_2521_),
    .Y(_2530_)
);

NAND2X1 _6167_ (
    .A(_2528_),
    .B(_2530_),
    .Y(_2531_)
);

INVX1 _6168_ (
    .A(_2517_),
    .Y(_2532_)
);

INVX1 _6169_ (
    .A(_2529_),
    .Y(_2533_)
);

AOI22X1 _6170_ (
    .A(\z4.q3 [5]),
    .B(_2532_),
    .C(_2515_),
    .D(_2533_),
    .Y(_2534_)
);

NAND2X1 _6171_ (
    .A(\z4.q3 [6]),
    .B(_2534_),
    .Y(_2535_)
);

NAND2X1 _6172_ (
    .A(_2535_),
    .B(_2531_),
    .Y(q3[14])
);

OAI21X1 _6173_ (
    .A(_2528_),
    .B(_2534_),
    .C(\z4.q3 [7]),
    .Y(_2536_)
);

INVX1 _6174_ (
    .A(\z4.q3 [7]),
    .Y(_2537_)
);

NAND3X1 _6175_ (
    .A(\z4.q3 [6]),
    .B(_2537_),
    .C(_2530_),
    .Y(_2538_)
);

NAND2X1 _6176_ (
    .A(_2538_),
    .B(_2536_),
    .Y(q3[15])
);

NOR2X1 _6177_ (
    .A(_2544_),
    .B(_2557_),
    .Y(_2539_)
);

NOR2X1 _6178_ (
    .A(_2539_),
    .B(_2578_),
    .Y(q3[5])
);

NOR2X1 _6179_ (
    .A(\z4.z1.q1 [0]),
    .B(\z4.z1.z1.z2.s ),
    .Y(_2604_)
);

AND2X2 _6180_ (
    .A(\z4.z1.q1 [0]),
    .B(\z4.z1.z1.z2.s ),
    .Y(_2605_)
);

NOR2X1 _6181_ (
    .A(_2604_),
    .B(_2605_),
    .Y(_2606_)
);

NAND2X1 _6182_ (
    .A(\z4.z1.q2 [0]),
    .B(_2606_),
    .Y(_2607_)
);

INVX1 _6183_ (
    .A(_2607_),
    .Y(_2608_)
);

NOR2X1 _6184_ (
    .A(\z4.z1.q2 [0]),
    .B(_2606_),
    .Y(_2609_)
);

NOR2X1 _6185_ (
    .A(_2609_),
    .B(_2608_),
    .Y(q3[2])
);

NAND2X1 _6186_ (
    .A(\z4.z1.q1 [0]),
    .B(\z4.z1.z1.z2.s ),
    .Y(_2610_)
);

NOR2X1 _6187_ (
    .A(\z4.z1.z2.z1.s ),
    .B(\z4.z1.z1.z2.c ),
    .Y(_2611_)
);

NAND2X1 _6188_ (
    .A(\z4.z1.z2.z1.s ),
    .B(\z4.z1.z1.z2.c ),
    .Y(_2612_)
);

INVX1 _6189_ (
    .A(_2612_),
    .Y(_2613_)
);

OAI21X1 _6190_ (
    .A(_2611_),
    .B(_2613_),
    .C(_2610_),
    .Y(_2614_)
);

INVX1 _6191_ (
    .A(\z4.z1.z2.z1.s ),
    .Y(_2615_)
);

INVX1 _6192_ (
    .A(\z4.z1.z1.z2.c ),
    .Y(_2616_)
);

NAND2X1 _6193_ (
    .A(_2615_),
    .B(_2616_),
    .Y(_2617_)
);

NAND3X1 _6194_ (
    .A(_2605_),
    .B(_2612_),
    .C(_2617_),
    .Y(_2618_)
);

NAND3X1 _6195_ (
    .A(\z4.z1.z3.z1.s ),
    .B(_2618_),
    .C(_2614_),
    .Y(_2619_)
);

INVX1 _6196_ (
    .A(\z4.z1.z3.z1.s ),
    .Y(_2620_)
);

NAND2X1 _6197_ (
    .A(_2618_),
    .B(_2614_),
    .Y(_2621_)
);

NAND2X1 _6198_ (
    .A(_2620_),
    .B(_2621_),
    .Y(_2622_)
);

NAND3X1 _6199_ (
    .A(_2608_),
    .B(_2619_),
    .C(_2622_),
    .Y(_2623_)
);

INVX1 _6200_ (
    .A(_2623_),
    .Y(_2624_)
);

INVX1 _6201_ (
    .A(_2619_),
    .Y(_2625_)
);

OAI21X1 _6202_ (
    .A(_2610_),
    .B(_2611_),
    .C(_2612_),
    .Y(_2626_)
);

NAND2X1 _6203_ (
    .A(\z4.z1.z2.z2.s ),
    .B(_2626_),
    .Y(_2627_)
);

INVX1 _6204_ (
    .A(\z4.z1.z2.z2.s ),
    .Y(_2628_)
);

NAND3X1 _6205_ (
    .A(_2628_),
    .B(_2612_),
    .C(_2618_),
    .Y(_2629_)
);

NAND2X1 _6206_ (
    .A(\z4.z1.q3 [0]),
    .B(\z4.z1.z3.z2.s ),
    .Y(_2630_)
);

INVX1 _6207_ (
    .A(\z4.z1.q3 [0]),
    .Y(_2631_)
);

INVX1 _6208_ (
    .A(\z4.z1.z3.z2.s ),
    .Y(_2632_)
);

NAND2X1 _6209_ (
    .A(_2631_),
    .B(_2632_),
    .Y(_2633_)
);

NAND2X1 _6210_ (
    .A(_2630_),
    .B(_2633_),
    .Y(_2634_)
);

INVX1 _6211_ (
    .A(_2634_),
    .Y(_2635_)
);

NAND3X1 _6212_ (
    .A(_2627_),
    .B(_2635_),
    .C(_2629_),
    .Y(_2636_)
);

AND2X2 _6213_ (
    .A(_2626_),
    .B(\z4.z1.z2.z2.s ),
    .Y(_2637_)
);

NOR2X1 _6214_ (
    .A(\z4.z1.z2.z2.s ),
    .B(_2626_),
    .Y(_2638_)
);

OAI21X1 _6215_ (
    .A(_2638_),
    .B(_2637_),
    .C(_2634_),
    .Y(_2639_)
);

NAND3X1 _6216_ (
    .A(_2625_),
    .B(_2636_),
    .C(_2639_),
    .Y(_2640_)
);

INVX1 _6217_ (
    .A(_2636_),
    .Y(_2641_)
);

AOI21X1 _6218_ (
    .A(_2629_),
    .B(_2627_),
    .C(_2635_),
    .Y(_2642_)
);

OAI21X1 _6219_ (
    .A(_2642_),
    .B(_2641_),
    .C(_2619_),
    .Y(_2643_)
);

NAND3X1 _6220_ (
    .A(_2624_),
    .B(_2640_),
    .C(_2643_),
    .Y(_2644_)
);

INVX1 _6221_ (
    .A(_2640_),
    .Y(_2645_)
);

INVX1 _6222_ (
    .A(_2621_),
    .Y(_2646_)
);

AOI22X1 _6223_ (
    .A(\z4.z1.z3.z1.s ),
    .B(_2646_),
    .C(_2639_),
    .D(_2636_),
    .Y(_2647_)
);

OAI21X1 _6224_ (
    .A(_2647_),
    .B(_2645_),
    .C(_2623_),
    .Y(_2648_)
);

AND2X2 _6225_ (
    .A(_2648_),
    .B(_2644_),
    .Y(\z4.q0 [4])
);

OAI21X1 _6226_ (
    .A(_2623_),
    .B(_2647_),
    .C(_2640_),
    .Y(_2649_)
);

OAI21X1 _6227_ (
    .A(_2631_),
    .B(_2632_),
    .C(_2636_),
    .Y(_2650_)
);

NAND2X1 _6228_ (
    .A(\z4.z1.z4.z1.s ),
    .B(\z4.z1.z3.z2.c ),
    .Y(_2651_)
);

OR2X2 _6229_ (
    .A(\z4.z1.z4.z1.s ),
    .B(\z4.z1.z3.z2.c ),
    .Y(_2652_)
);

NAND2X1 _6230_ (
    .A(_2651_),
    .B(_2652_),
    .Y(_2653_)
);

INVX1 _6231_ (
    .A(_2653_),
    .Y(_2654_)
);

NAND2X1 _6232_ (
    .A(\z4.z1.z2.z2.c ),
    .B(_2637_),
    .Y(_2655_)
);

INVX1 _6233_ (
    .A(\z4.z1.z2.z2.c ),
    .Y(_2656_)
);

NAND2X1 _6234_ (
    .A(_2656_),
    .B(_2627_),
    .Y(_2657_)
);

NAND3X1 _6235_ (
    .A(_2654_),
    .B(_2657_),
    .C(_2655_),
    .Y(_2658_)
);

NAND2X1 _6236_ (
    .A(\z4.z1.z2.z2.c ),
    .B(_2627_),
    .Y(_2659_)
);

NAND2X1 _6237_ (
    .A(_2656_),
    .B(_2637_),
    .Y(_2660_)
);

NAND3X1 _6238_ (
    .A(_2653_),
    .B(_2659_),
    .C(_2660_),
    .Y(_2661_)
);

NAND3X1 _6239_ (
    .A(_2650_),
    .B(_2658_),
    .C(_2661_),
    .Y(_2662_)
);

INVX1 _6240_ (
    .A(_2650_),
    .Y(_2663_)
);

AOI21X1 _6241_ (
    .A(_2660_),
    .B(_2659_),
    .C(_2653_),
    .Y(_2664_)
);

AOI21X1 _6242_ (
    .A(_2655_),
    .B(_2657_),
    .C(_2654_),
    .Y(_2665_)
);

OAI21X1 _6243_ (
    .A(_2664_),
    .B(_2665_),
    .C(_2663_),
    .Y(_2666_)
);

NAND2X1 _6244_ (
    .A(_2662_),
    .B(_2666_),
    .Y(_2667_)
);

NAND2X1 _6245_ (
    .A(_2649_),
    .B(_2667_),
    .Y(_2668_)
);

OR2X2 _6246_ (
    .A(_2667_),
    .B(_2649_),
    .Y(_2669_)
);

NAND2X1 _6247_ (
    .A(_2668_),
    .B(_2669_),
    .Y(\z4.q0 [5])
);

INVX1 _6248_ (
    .A(\z4.z1.z4.z2.s ),
    .Y(_2670_)
);

INVX1 _6249_ (
    .A(_2651_),
    .Y(_2671_)
);

OAI21X1 _6250_ (
    .A(_2671_),
    .B(_2664_),
    .C(_2670_),
    .Y(_2672_)
);

NAND3X1 _6251_ (
    .A(\z4.z1.z4.z2.s ),
    .B(_2651_),
    .C(_2658_),
    .Y(_2673_)
);

NAND2X1 _6252_ (
    .A(_2666_),
    .B(_2649_),
    .Y(_2674_)
);

AOI22X1 _6253_ (
    .A(_2672_),
    .B(_2673_),
    .C(_2674_),
    .D(_2662_),
    .Y(_2675_)
);

NAND2X1 _6254_ (
    .A(_2673_),
    .B(_2672_),
    .Y(_2676_)
);

NAND3X1 _6255_ (
    .A(_2640_),
    .B(_2662_),
    .C(_2644_),
    .Y(_2677_)
);

AOI21X1 _6256_ (
    .A(_2677_),
    .B(_2666_),
    .C(_2676_),
    .Y(_2678_)
);

NOR2X1 _6257_ (
    .A(_2675_),
    .B(_2678_),
    .Y(\z4.q0 [6])
);

OAI21X1 _6258_ (
    .A(_2671_),
    .B(_2664_),
    .C(\z4.z1.z4.z2.s ),
    .Y(_2597_)
);

NAND3X1 _6259_ (
    .A(_2666_),
    .B(_2676_),
    .C(_2677_),
    .Y(_2598_)
);

NAND3X1 _6260_ (
    .A(\z4.z1.z4.z2.c ),
    .B(_2597_),
    .C(_2598_),
    .Y(_2599_)
);

INVX1 _6261_ (
    .A(\z4.z1.z4.z2.c ),
    .Y(_2600_)
);

INVX1 _6262_ (
    .A(_2597_),
    .Y(_2601_)
);

OAI21X1 _6263_ (
    .A(_2601_),
    .B(_2675_),
    .C(_2600_),
    .Y(_2602_)
);

NAND2X1 _6264_ (
    .A(_2599_),
    .B(_2602_),
    .Y(\z4.q0 [7])
);

AOI21X1 _6265_ (
    .A(_2622_),
    .B(_2619_),
    .C(_2608_),
    .Y(_2603_)
);

NOR2X1 _6266_ (
    .A(_2603_),
    .B(_2624_),
    .Y(q3[3])
);

AND2X2 _6267_ (
    .A(b[8]),
    .B(a[8]),
    .Y(q3[0])
);

AND2X2 _6268_ (
    .A(b[8]),
    .B(a[9]),
    .Y(\z4.z1.z1.z1.a )
);

AND2X2 _6269_ (
    .A(a[8]),
    .B(b[9]),
    .Y(\z4.z1.z1.z1.b )
);

AND2X2 _6270_ (
    .A(a[9]),
    .B(b[9]),
    .Y(\z4.z1.z1.z2.a )
);

INVX1 _6271_ (
    .A(\z4.z1.z1.z1.b ),
    .Y(_2679_)
);

NAND2X1 _6272_ (
    .A(\z4.z1.z1.z1.a ),
    .B(_2679_),
    .Y(_2680_)
);

INVX1 _6273_ (
    .A(\z4.z1.z1.z1.a ),
    .Y(_2681_)
);

NAND2X1 _6274_ (
    .A(\z4.z1.z1.z1.b ),
    .B(_2681_),
    .Y(_2682_)
);

NAND2X1 _6275_ (
    .A(_2680_),
    .B(_2682_),
    .Y(\z4.z1.z1.z1.s )
);

NOR2X1 _6276_ (
    .A(_2679_),
    .B(_2681_),
    .Y(\z4.z1.z1.z1.c )
);

INVX1 _6277_ (
    .A(\z4.z1.z1.z1.c ),
    .Y(_2683_)
);

NAND2X1 _6278_ (
    .A(\z4.z1.z1.z2.a ),
    .B(_2683_),
    .Y(_2684_)
);

INVX1 _6279_ (
    .A(\z4.z1.z1.z2.a ),
    .Y(_2685_)
);

NAND2X1 _6280_ (
    .A(\z4.z1.z1.z1.c ),
    .B(_2685_),
    .Y(_2686_)
);

NAND2X1 _6281_ (
    .A(_2684_),
    .B(_2686_),
    .Y(\z4.z1.z1.z2.s )
);

NOR2X1 _6282_ (
    .A(_2683_),
    .B(_2685_),
    .Y(\z4.z1.z1.z2.c )
);

AND2X2 _6283_ (
    .A(b[8]),
    .B(a[10]),
    .Y(\z4.z1.q1 [0])
);

AND2X2 _6284_ (
    .A(b[8]),
    .B(a[11]),
    .Y(\z4.z1.z2.z1.a )
);

AND2X2 _6285_ (
    .A(a[10]),
    .B(b[9]),
    .Y(\z4.z1.z2.z1.b )
);

AND2X2 _6286_ (
    .A(a[11]),
    .B(b[9]),
    .Y(\z4.z1.z2.z2.a )
);

INVX1 _6287_ (
    .A(\z4.z1.z2.z1.b ),
    .Y(_2687_)
);

NAND2X1 _6288_ (
    .A(\z4.z1.z2.z1.a ),
    .B(_2687_),
    .Y(_2688_)
);

INVX1 _6289_ (
    .A(\z4.z1.z2.z1.a ),
    .Y(_2689_)
);

NAND2X1 _6290_ (
    .A(\z4.z1.z2.z1.b ),
    .B(_2689_),
    .Y(_2690_)
);

NAND2X1 _6291_ (
    .A(_2688_),
    .B(_2690_),
    .Y(\z4.z1.z2.z1.s )
);

NOR2X1 _6292_ (
    .A(_2687_),
    .B(_2689_),
    .Y(\z4.z1.z2.z1.c )
);

INVX1 _6293_ (
    .A(\z4.z1.z2.z1.c ),
    .Y(_2691_)
);

NAND2X1 _6294_ (
    .A(\z4.z1.z2.z2.a ),
    .B(_2691_),
    .Y(_2692_)
);

INVX1 _6295_ (
    .A(\z4.z1.z2.z2.a ),
    .Y(_2693_)
);

NAND2X1 _6296_ (
    .A(\z4.z1.z2.z1.c ),
    .B(_2693_),
    .Y(_2694_)
);

NAND2X1 _6297_ (
    .A(_2692_),
    .B(_2694_),
    .Y(\z4.z1.z2.z2.s )
);

NOR2X1 _6298_ (
    .A(_2691_),
    .B(_2693_),
    .Y(\z4.z1.z2.z2.c )
);

AND2X2 _6299_ (
    .A(b[10]),
    .B(a[8]),
    .Y(\z4.z1.q2 [0])
);

AND2X2 _6300_ (
    .A(b[10]),
    .B(a[9]),
    .Y(\z4.z1.z3.z1.a )
);

AND2X2 _6301_ (
    .A(a[8]),
    .B(b[11]),
    .Y(\z4.z1.z3.z1.b )
);

AND2X2 _6302_ (
    .A(a[9]),
    .B(b[11]),
    .Y(\z4.z1.z3.z2.a )
);

INVX1 _6303_ (
    .A(\z4.z1.z3.z1.b ),
    .Y(_2695_)
);

NAND2X1 _6304_ (
    .A(\z4.z1.z3.z1.a ),
    .B(_2695_),
    .Y(_2696_)
);

INVX1 _6305_ (
    .A(\z4.z1.z3.z1.a ),
    .Y(_2697_)
);

NAND2X1 _6306_ (
    .A(\z4.z1.z3.z1.b ),
    .B(_2697_),
    .Y(_2698_)
);

NAND2X1 _6307_ (
    .A(_2696_),
    .B(_2698_),
    .Y(\z4.z1.z3.z1.s )
);

NOR2X1 _6308_ (
    .A(_2695_),
    .B(_2697_),
    .Y(\z4.z1.z3.z1.c )
);

INVX1 _6309_ (
    .A(\z4.z1.z3.z1.c ),
    .Y(_2699_)
);

NAND2X1 _6310_ (
    .A(\z4.z1.z3.z2.a ),
    .B(_2699_),
    .Y(_2700_)
);

INVX1 _6311_ (
    .A(\z4.z1.z3.z2.a ),
    .Y(_2701_)
);

NAND2X1 _6312_ (
    .A(\z4.z1.z3.z1.c ),
    .B(_2701_),
    .Y(_2702_)
);

NAND2X1 _6313_ (
    .A(_2700_),
    .B(_2702_),
    .Y(\z4.z1.z3.z2.s )
);

NOR2X1 _6314_ (
    .A(_2699_),
    .B(_2701_),
    .Y(\z4.z1.z3.z2.c )
);

AND2X2 _6315_ (
    .A(b[10]),
    .B(a[10]),
    .Y(\z4.z1.q3 [0])
);

AND2X2 _6316_ (
    .A(b[10]),
    .B(a[11]),
    .Y(\z4.z1.z4.z1.a )
);

AND2X2 _6317_ (
    .A(a[10]),
    .B(b[11]),
    .Y(\z4.z1.z4.z1.b )
);

AND2X2 _6318_ (
    .A(a[11]),
    .B(b[11]),
    .Y(\z4.z1.z4.z2.a )
);

INVX1 _6319_ (
    .A(\z4.z1.z4.z1.b ),
    .Y(_2703_)
);

NAND2X1 _6320_ (
    .A(\z4.z1.z4.z1.a ),
    .B(_2703_),
    .Y(_2704_)
);

INVX1 _6321_ (
    .A(\z4.z1.z4.z1.a ),
    .Y(_2705_)
);

NAND2X1 _6322_ (
    .A(\z4.z1.z4.z1.b ),
    .B(_2705_),
    .Y(_2706_)
);

NAND2X1 _6323_ (
    .A(_2704_),
    .B(_2706_),
    .Y(\z4.z1.z4.z1.s )
);

NOR2X1 _6324_ (
    .A(_2703_),
    .B(_2705_),
    .Y(\z4.z1.z4.z1.c )
);

INVX1 _6325_ (
    .A(\z4.z1.z4.z1.c ),
    .Y(_2707_)
);

NAND2X1 _6326_ (
    .A(\z4.z1.z4.z2.a ),
    .B(_2707_),
    .Y(_2708_)
);

INVX1 _6327_ (
    .A(\z4.z1.z4.z2.a ),
    .Y(_2709_)
);

NAND2X1 _6328_ (
    .A(\z4.z1.z4.z1.c ),
    .B(_2709_),
    .Y(_2710_)
);

NAND2X1 _6329_ (
    .A(_2708_),
    .B(_2710_),
    .Y(\z4.z1.z4.z2.s )
);

NOR2X1 _6330_ (
    .A(_2707_),
    .B(_2709_),
    .Y(\z4.z1.z4.z2.c )
);

NOR2X1 _6331_ (
    .A(\z4.z2.q1 [0]),
    .B(\z4.z2.z1.z2.s ),
    .Y(_2718_)
);

AND2X2 _6332_ (
    .A(\z4.z2.q1 [0]),
    .B(\z4.z2.z1.z2.s ),
    .Y(_2719_)
);

NOR2X1 _6333_ (
    .A(_2718_),
    .B(_2719_),
    .Y(_2720_)
);

NAND2X1 _6334_ (
    .A(\z4.z2.q2 [0]),
    .B(_2720_),
    .Y(_2721_)
);

INVX1 _6335_ (
    .A(_2721_),
    .Y(_2722_)
);

NOR2X1 _6336_ (
    .A(\z4.z2.q2 [0]),
    .B(_2720_),
    .Y(_2723_)
);

NOR2X1 _6337_ (
    .A(_2723_),
    .B(_2722_),
    .Y(\z4.q1 [2])
);

NAND2X1 _6338_ (
    .A(\z4.z2.q1 [0]),
    .B(\z4.z2.z1.z2.s ),
    .Y(_2724_)
);

NOR2X1 _6339_ (
    .A(\z4.z2.z2.z1.s ),
    .B(\z4.z2.z1.z2.c ),
    .Y(_2725_)
);

NAND2X1 _6340_ (
    .A(\z4.z2.z2.z1.s ),
    .B(\z4.z2.z1.z2.c ),
    .Y(_2726_)
);

INVX1 _6341_ (
    .A(_2726_),
    .Y(_2727_)
);

OAI21X1 _6342_ (
    .A(_2725_),
    .B(_2727_),
    .C(_2724_),
    .Y(_2728_)
);

INVX1 _6343_ (
    .A(\z4.z2.z2.z1.s ),
    .Y(_2729_)
);

INVX1 _6344_ (
    .A(\z4.z2.z1.z2.c ),
    .Y(_2730_)
);

NAND2X1 _6345_ (
    .A(_2729_),
    .B(_2730_),
    .Y(_2731_)
);

NAND3X1 _6346_ (
    .A(_2719_),
    .B(_2726_),
    .C(_2731_),
    .Y(_2732_)
);

NAND3X1 _6347_ (
    .A(\z4.z2.z3.z1.s ),
    .B(_2732_),
    .C(_2728_),
    .Y(_2733_)
);

INVX1 _6348_ (
    .A(\z4.z2.z3.z1.s ),
    .Y(_2734_)
);

NAND2X1 _6349_ (
    .A(_2732_),
    .B(_2728_),
    .Y(_2735_)
);

NAND2X1 _6350_ (
    .A(_2734_),
    .B(_2735_),
    .Y(_2736_)
);

NAND3X1 _6351_ (
    .A(_2722_),
    .B(_2733_),
    .C(_2736_),
    .Y(_2737_)
);

INVX1 _6352_ (
    .A(_2737_),
    .Y(_2738_)
);

INVX1 _6353_ (
    .A(_2733_),
    .Y(_2739_)
);

OAI21X1 _6354_ (
    .A(_2724_),
    .B(_2725_),
    .C(_2726_),
    .Y(_2740_)
);

NAND2X1 _6355_ (
    .A(\z4.z2.z2.z2.s ),
    .B(_2740_),
    .Y(_2741_)
);

INVX1 _6356_ (
    .A(\z4.z2.z2.z2.s ),
    .Y(_2742_)
);

NAND3X1 _6357_ (
    .A(_2742_),
    .B(_2726_),
    .C(_2732_),
    .Y(_2743_)
);

NAND2X1 _6358_ (
    .A(\z4.z2.q3 [0]),
    .B(\z4.z2.z3.z2.s ),
    .Y(_2744_)
);

INVX1 _6359_ (
    .A(\z4.z2.q3 [0]),
    .Y(_2745_)
);

INVX1 _6360_ (
    .A(\z4.z2.z3.z2.s ),
    .Y(_2746_)
);

NAND2X1 _6361_ (
    .A(_2745_),
    .B(_2746_),
    .Y(_2747_)
);

NAND2X1 _6362_ (
    .A(_2744_),
    .B(_2747_),
    .Y(_2748_)
);

INVX1 _6363_ (
    .A(_2748_),
    .Y(_2749_)
);

NAND3X1 _6364_ (
    .A(_2741_),
    .B(_2749_),
    .C(_2743_),
    .Y(_2750_)
);

AND2X2 _6365_ (
    .A(_2740_),
    .B(\z4.z2.z2.z2.s ),
    .Y(_2751_)
);

NOR2X1 _6366_ (
    .A(\z4.z2.z2.z2.s ),
    .B(_2740_),
    .Y(_2752_)
);

OAI21X1 _6367_ (
    .A(_2752_),
    .B(_2751_),
    .C(_2748_),
    .Y(_2753_)
);

NAND3X1 _6368_ (
    .A(_2739_),
    .B(_2750_),
    .C(_2753_),
    .Y(_2754_)
);

INVX1 _6369_ (
    .A(_2750_),
    .Y(_2755_)
);

AOI21X1 _6370_ (
    .A(_2743_),
    .B(_2741_),
    .C(_2749_),
    .Y(_2756_)
);

OAI21X1 _6371_ (
    .A(_2756_),
    .B(_2755_),
    .C(_2733_),
    .Y(_2757_)
);

NAND3X1 _6372_ (
    .A(_2738_),
    .B(_2754_),
    .C(_2757_),
    .Y(_2758_)
);

INVX1 _6373_ (
    .A(_2754_),
    .Y(_2759_)
);

INVX1 _6374_ (
    .A(_2735_),
    .Y(_2760_)
);

AOI22X1 _6375_ (
    .A(\z4.z2.z3.z1.s ),
    .B(_2760_),
    .C(_2753_),
    .D(_2750_),
    .Y(_2761_)
);

OAI21X1 _6376_ (
    .A(_2761_),
    .B(_2759_),
    .C(_2737_),
    .Y(_2762_)
);

AND2X2 _6377_ (
    .A(_2762_),
    .B(_2758_),
    .Y(\z4.q1 [4])
);

OAI21X1 _6378_ (
    .A(_2737_),
    .B(_2761_),
    .C(_2754_),
    .Y(_2763_)
);

OAI21X1 _6379_ (
    .A(_2745_),
    .B(_2746_),
    .C(_2750_),
    .Y(_2764_)
);

NAND2X1 _6380_ (
    .A(\z4.z2.z4.z1.s ),
    .B(\z4.z2.z3.z2.c ),
    .Y(_2765_)
);

OR2X2 _6381_ (
    .A(\z4.z2.z4.z1.s ),
    .B(\z4.z2.z3.z2.c ),
    .Y(_2766_)
);

NAND2X1 _6382_ (
    .A(_2765_),
    .B(_2766_),
    .Y(_2767_)
);

INVX1 _6383_ (
    .A(_2767_),
    .Y(_2768_)
);

NAND2X1 _6384_ (
    .A(\z4.z2.z2.z2.c ),
    .B(_2751_),
    .Y(_2769_)
);

INVX1 _6385_ (
    .A(\z4.z2.z2.z2.c ),
    .Y(_2770_)
);

NAND2X1 _6386_ (
    .A(_2770_),
    .B(_2741_),
    .Y(_2771_)
);

NAND3X1 _6387_ (
    .A(_2768_),
    .B(_2771_),
    .C(_2769_),
    .Y(_2772_)
);

NAND2X1 _6388_ (
    .A(\z4.z2.z2.z2.c ),
    .B(_2741_),
    .Y(_2773_)
);

NAND2X1 _6389_ (
    .A(_2770_),
    .B(_2751_),
    .Y(_2774_)
);

NAND3X1 _6390_ (
    .A(_2767_),
    .B(_2773_),
    .C(_2774_),
    .Y(_2775_)
);

NAND3X1 _6391_ (
    .A(_2764_),
    .B(_2772_),
    .C(_2775_),
    .Y(_2776_)
);

INVX1 _6392_ (
    .A(_2764_),
    .Y(_2777_)
);

AOI21X1 _6393_ (
    .A(_2774_),
    .B(_2773_),
    .C(_2767_),
    .Y(_2778_)
);

AOI21X1 _6394_ (
    .A(_2769_),
    .B(_2771_),
    .C(_2768_),
    .Y(_2779_)
);

OAI21X1 _6395_ (
    .A(_2778_),
    .B(_2779_),
    .C(_2777_),
    .Y(_2780_)
);

NAND2X1 _6396_ (
    .A(_2776_),
    .B(_2780_),
    .Y(_2781_)
);

NAND2X1 _6397_ (
    .A(_2763_),
    .B(_2781_),
    .Y(_2782_)
);

OR2X2 _6398_ (
    .A(_2781_),
    .B(_2763_),
    .Y(_2783_)
);

NAND2X1 _6399_ (
    .A(_2782_),
    .B(_2783_),
    .Y(\z4.q1 [5])
);

INVX1 _6400_ (
    .A(\z4.z2.z4.z2.s ),
    .Y(_2784_)
);

INVX1 _6401_ (
    .A(_2765_),
    .Y(_2785_)
);

OAI21X1 _6402_ (
    .A(_2785_),
    .B(_2778_),
    .C(_2784_),
    .Y(_2786_)
);

NAND3X1 _6403_ (
    .A(\z4.z2.z4.z2.s ),
    .B(_2765_),
    .C(_2772_),
    .Y(_2787_)
);

NAND2X1 _6404_ (
    .A(_2780_),
    .B(_2763_),
    .Y(_2788_)
);

AOI22X1 _6405_ (
    .A(_2786_),
    .B(_2787_),
    .C(_2788_),
    .D(_2776_),
    .Y(_2789_)
);

NAND2X1 _6406_ (
    .A(_2787_),
    .B(_2786_),
    .Y(_2790_)
);

NAND3X1 _6407_ (
    .A(_2754_),
    .B(_2776_),
    .C(_2758_),
    .Y(_2791_)
);

AOI21X1 _6408_ (
    .A(_2791_),
    .B(_2780_),
    .C(_2790_),
    .Y(_2792_)
);

NOR2X1 _6409_ (
    .A(_2789_),
    .B(_2792_),
    .Y(\z4.q1 [6])
);

OAI21X1 _6410_ (
    .A(_2785_),
    .B(_2778_),
    .C(\z4.z2.z4.z2.s ),
    .Y(_2711_)
);

NAND3X1 _6411_ (
    .A(_2780_),
    .B(_2790_),
    .C(_2791_),
    .Y(_2712_)
);

NAND3X1 _6412_ (
    .A(\z4.z2.z4.z2.c ),
    .B(_2711_),
    .C(_2712_),
    .Y(_2713_)
);

INVX1 _6413_ (
    .A(\z4.z2.z4.z2.c ),
    .Y(_2714_)
);

INVX1 _6414_ (
    .A(_2711_),
    .Y(_2715_)
);

OAI21X1 _6415_ (
    .A(_2715_),
    .B(_2789_),
    .C(_2714_),
    .Y(_2716_)
);

NAND2X1 _6416_ (
    .A(_2713_),
    .B(_2716_),
    .Y(\z4.q1 [7])
);

AOI21X1 _6417_ (
    .A(_2736_),
    .B(_2733_),
    .C(_2722_),
    .Y(_2717_)
);

NOR2X1 _6418_ (
    .A(_2717_),
    .B(_2738_),
    .Y(\z4.q1 [3])
);

AND2X2 _6419_ (
    .A(b[8]),
    .B(a[12]),
    .Y(\z4.q1 [0])
);

AND2X2 _6420_ (
    .A(b[8]),
    .B(a[13]),
    .Y(\z4.z2.z1.z1.a )
);

AND2X2 _6421_ (
    .A(a[12]),
    .B(b[9]),
    .Y(\z4.z2.z1.z1.b )
);

AND2X2 _6422_ (
    .A(a[13]),
    .B(b[9]),
    .Y(\z4.z2.z1.z2.a )
);

INVX1 _6423_ (
    .A(\z4.z2.z1.z1.b ),
    .Y(_2793_)
);

NAND2X1 _6424_ (
    .A(\z4.z2.z1.z1.a ),
    .B(_2793_),
    .Y(_2794_)
);

INVX1 _6425_ (
    .A(\z4.z2.z1.z1.a ),
    .Y(_2795_)
);

NAND2X1 _6426_ (
    .A(\z4.z2.z1.z1.b ),
    .B(_2795_),
    .Y(_2796_)
);

NAND2X1 _6427_ (
    .A(_2794_),
    .B(_2796_),
    .Y(\z4.z2.z1.z1.s )
);

NOR2X1 _6428_ (
    .A(_2793_),
    .B(_2795_),
    .Y(\z4.z2.z1.z1.c )
);

INVX1 _6429_ (
    .A(\z4.z2.z1.z1.c ),
    .Y(_2797_)
);

NAND2X1 _6430_ (
    .A(\z4.z2.z1.z2.a ),
    .B(_2797_),
    .Y(_2798_)
);

INVX1 _6431_ (
    .A(\z4.z2.z1.z2.a ),
    .Y(_2799_)
);

NAND2X1 _6432_ (
    .A(\z4.z2.z1.z1.c ),
    .B(_2799_),
    .Y(_2800_)
);

NAND2X1 _6433_ (
    .A(_2798_),
    .B(_2800_),
    .Y(\z4.z2.z1.z2.s )
);

NOR2X1 _6434_ (
    .A(_2797_),
    .B(_2799_),
    .Y(\z4.z2.z1.z2.c )
);

AND2X2 _6435_ (
    .A(b[8]),
    .B(a[14]),
    .Y(\z4.z2.q1 [0])
);

AND2X2 _6436_ (
    .A(b[8]),
    .B(a[15]),
    .Y(\z4.z2.z2.z1.a )
);

AND2X2 _6437_ (
    .A(a[14]),
    .B(b[9]),
    .Y(\z4.z2.z2.z1.b )
);

AND2X2 _6438_ (
    .A(a[15]),
    .B(b[9]),
    .Y(\z4.z2.z2.z2.a )
);

INVX1 _6439_ (
    .A(\z4.z2.z2.z1.b ),
    .Y(_2801_)
);

NAND2X1 _6440_ (
    .A(\z4.z2.z2.z1.a ),
    .B(_2801_),
    .Y(_2802_)
);

INVX1 _6441_ (
    .A(\z4.z2.z2.z1.a ),
    .Y(_2803_)
);

NAND2X1 _6442_ (
    .A(\z4.z2.z2.z1.b ),
    .B(_2803_),
    .Y(_2804_)
);

NAND2X1 _6443_ (
    .A(_2802_),
    .B(_2804_),
    .Y(\z4.z2.z2.z1.s )
);

NOR2X1 _6444_ (
    .A(_2801_),
    .B(_2803_),
    .Y(\z4.z2.z2.z1.c )
);

INVX1 _6445_ (
    .A(\z4.z2.z2.z1.c ),
    .Y(_2805_)
);

NAND2X1 _6446_ (
    .A(\z4.z2.z2.z2.a ),
    .B(_2805_),
    .Y(_2806_)
);

INVX1 _6447_ (
    .A(\z4.z2.z2.z2.a ),
    .Y(_2807_)
);

NAND2X1 _6448_ (
    .A(\z4.z2.z2.z1.c ),
    .B(_2807_),
    .Y(_2808_)
);

NAND2X1 _6449_ (
    .A(_2806_),
    .B(_2808_),
    .Y(\z4.z2.z2.z2.s )
);

NOR2X1 _6450_ (
    .A(_2805_),
    .B(_2807_),
    .Y(\z4.z2.z2.z2.c )
);

AND2X2 _6451_ (
    .A(b[10]),
    .B(a[12]),
    .Y(\z4.z2.q2 [0])
);

AND2X2 _6452_ (
    .A(b[10]),
    .B(a[13]),
    .Y(\z4.z2.z3.z1.a )
);

AND2X2 _6453_ (
    .A(a[12]),
    .B(b[11]),
    .Y(\z4.z2.z3.z1.b )
);

AND2X2 _6454_ (
    .A(a[13]),
    .B(b[11]),
    .Y(\z4.z2.z3.z2.a )
);

INVX1 _6455_ (
    .A(\z4.z2.z3.z1.b ),
    .Y(_2809_)
);

NAND2X1 _6456_ (
    .A(\z4.z2.z3.z1.a ),
    .B(_2809_),
    .Y(_2810_)
);

INVX1 _6457_ (
    .A(\z4.z2.z3.z1.a ),
    .Y(_2811_)
);

NAND2X1 _6458_ (
    .A(\z4.z2.z3.z1.b ),
    .B(_2811_),
    .Y(_2812_)
);

NAND2X1 _6459_ (
    .A(_2810_),
    .B(_2812_),
    .Y(\z4.z2.z3.z1.s )
);

NOR2X1 _6460_ (
    .A(_2809_),
    .B(_2811_),
    .Y(\z4.z2.z3.z1.c )
);

INVX1 _6461_ (
    .A(\z4.z2.z3.z1.c ),
    .Y(_2813_)
);

NAND2X1 _6462_ (
    .A(\z4.z2.z3.z2.a ),
    .B(_2813_),
    .Y(_2814_)
);

INVX1 _6463_ (
    .A(\z4.z2.z3.z2.a ),
    .Y(_2815_)
);

NAND2X1 _6464_ (
    .A(\z4.z2.z3.z1.c ),
    .B(_2815_),
    .Y(_2816_)
);

NAND2X1 _6465_ (
    .A(_2814_),
    .B(_2816_),
    .Y(\z4.z2.z3.z2.s )
);

NOR2X1 _6466_ (
    .A(_2813_),
    .B(_2815_),
    .Y(\z4.z2.z3.z2.c )
);

AND2X2 _6467_ (
    .A(b[10]),
    .B(a[14]),
    .Y(\z4.z2.q3 [0])
);

AND2X2 _6468_ (
    .A(b[10]),
    .B(a[15]),
    .Y(\z4.z2.z4.z1.a )
);

AND2X2 _6469_ (
    .A(a[14]),
    .B(b[11]),
    .Y(\z4.z2.z4.z1.b )
);

AND2X2 _6470_ (
    .A(a[15]),
    .B(b[11]),
    .Y(\z4.z2.z4.z2.a )
);

INVX1 _6471_ (
    .A(\z4.z2.z4.z1.b ),
    .Y(_2817_)
);

NAND2X1 _6472_ (
    .A(\z4.z2.z4.z1.a ),
    .B(_2817_),
    .Y(_2818_)
);

INVX1 _6473_ (
    .A(\z4.z2.z4.z1.a ),
    .Y(_2819_)
);

NAND2X1 _6474_ (
    .A(\z4.z2.z4.z1.b ),
    .B(_2819_),
    .Y(_2820_)
);

NAND2X1 _6475_ (
    .A(_2818_),
    .B(_2820_),
    .Y(\z4.z2.z4.z1.s )
);

NOR2X1 _6476_ (
    .A(_2817_),
    .B(_2819_),
    .Y(\z4.z2.z4.z1.c )
);

INVX1 _6477_ (
    .A(\z4.z2.z4.z1.c ),
    .Y(_2821_)
);

NAND2X1 _6478_ (
    .A(\z4.z2.z4.z2.a ),
    .B(_2821_),
    .Y(_2822_)
);

INVX1 _6479_ (
    .A(\z4.z2.z4.z2.a ),
    .Y(_2823_)
);

NAND2X1 _6480_ (
    .A(\z4.z2.z4.z1.c ),
    .B(_2823_),
    .Y(_2824_)
);

NAND2X1 _6481_ (
    .A(_2822_),
    .B(_2824_),
    .Y(\z4.z2.z4.z2.s )
);

NOR2X1 _6482_ (
    .A(_2821_),
    .B(_2823_),
    .Y(\z4.z2.z4.z2.c )
);

NOR2X1 _6483_ (
    .A(\z4.z3.q1 [0]),
    .B(\z4.z3.z1.z2.s ),
    .Y(_2832_)
);

AND2X2 _6484_ (
    .A(\z4.z3.q1 [0]),
    .B(\z4.z3.z1.z2.s ),
    .Y(_2833_)
);

NOR2X1 _6485_ (
    .A(_2832_),
    .B(_2833_),
    .Y(_2834_)
);

NAND2X1 _6486_ (
    .A(\z4.z3.q2 [0]),
    .B(_2834_),
    .Y(_2835_)
);

INVX1 _6487_ (
    .A(_2835_),
    .Y(_2836_)
);

NOR2X1 _6488_ (
    .A(\z4.z3.q2 [0]),
    .B(_2834_),
    .Y(_2837_)
);

NOR2X1 _6489_ (
    .A(_2837_),
    .B(_2836_),
    .Y(\z4.q2 [2])
);

NAND2X1 _6490_ (
    .A(\z4.z3.q1 [0]),
    .B(\z4.z3.z1.z2.s ),
    .Y(_2838_)
);

NOR2X1 _6491_ (
    .A(\z4.z3.z2.z1.s ),
    .B(\z4.z3.z1.z2.c ),
    .Y(_2839_)
);

NAND2X1 _6492_ (
    .A(\z4.z3.z2.z1.s ),
    .B(\z4.z3.z1.z2.c ),
    .Y(_2840_)
);

INVX1 _6493_ (
    .A(_2840_),
    .Y(_2841_)
);

OAI21X1 _6494_ (
    .A(_2839_),
    .B(_2841_),
    .C(_2838_),
    .Y(_2842_)
);

INVX1 _6495_ (
    .A(\z4.z3.z2.z1.s ),
    .Y(_2843_)
);

INVX1 _6496_ (
    .A(\z4.z3.z1.z2.c ),
    .Y(_2844_)
);

NAND2X1 _6497_ (
    .A(_2843_),
    .B(_2844_),
    .Y(_2845_)
);

NAND3X1 _6498_ (
    .A(_2833_),
    .B(_2840_),
    .C(_2845_),
    .Y(_2846_)
);

NAND3X1 _6499_ (
    .A(\z4.z3.z3.z1.s ),
    .B(_2846_),
    .C(_2842_),
    .Y(_2847_)
);

INVX1 _6500_ (
    .A(\z4.z3.z3.z1.s ),
    .Y(_2848_)
);

NAND2X1 _6501_ (
    .A(_2846_),
    .B(_2842_),
    .Y(_2849_)
);

NAND2X1 _6502_ (
    .A(_2848_),
    .B(_2849_),
    .Y(_2850_)
);

NAND3X1 _6503_ (
    .A(_2836_),
    .B(_2847_),
    .C(_2850_),
    .Y(_2851_)
);

INVX1 _6504_ (
    .A(_2851_),
    .Y(_2852_)
);

INVX1 _6505_ (
    .A(_2847_),
    .Y(_2853_)
);

OAI21X1 _6506_ (
    .A(_2838_),
    .B(_2839_),
    .C(_2840_),
    .Y(_2854_)
);

NAND2X1 _6507_ (
    .A(\z4.z3.z2.z2.s ),
    .B(_2854_),
    .Y(_2855_)
);

INVX1 _6508_ (
    .A(\z4.z3.z2.z2.s ),
    .Y(_2856_)
);

NAND3X1 _6509_ (
    .A(_2856_),
    .B(_2840_),
    .C(_2846_),
    .Y(_2857_)
);

NAND2X1 _6510_ (
    .A(\z4.z3.q3 [0]),
    .B(\z4.z3.z3.z2.s ),
    .Y(_2858_)
);

INVX1 _6511_ (
    .A(\z4.z3.q3 [0]),
    .Y(_2859_)
);

INVX1 _6512_ (
    .A(\z4.z3.z3.z2.s ),
    .Y(_2860_)
);

NAND2X1 _6513_ (
    .A(_2859_),
    .B(_2860_),
    .Y(_2861_)
);

NAND2X1 _6514_ (
    .A(_2858_),
    .B(_2861_),
    .Y(_2862_)
);

INVX1 _6515_ (
    .A(_2862_),
    .Y(_2863_)
);

NAND3X1 _6516_ (
    .A(_2855_),
    .B(_2863_),
    .C(_2857_),
    .Y(_2864_)
);

AND2X2 _6517_ (
    .A(_2854_),
    .B(\z4.z3.z2.z2.s ),
    .Y(_2865_)
);

NOR2X1 _6518_ (
    .A(\z4.z3.z2.z2.s ),
    .B(_2854_),
    .Y(_2866_)
);

OAI21X1 _6519_ (
    .A(_2866_),
    .B(_2865_),
    .C(_2862_),
    .Y(_2867_)
);

NAND3X1 _6520_ (
    .A(_2853_),
    .B(_2864_),
    .C(_2867_),
    .Y(_2868_)
);

INVX1 _6521_ (
    .A(_2864_),
    .Y(_2869_)
);

AOI21X1 _6522_ (
    .A(_2857_),
    .B(_2855_),
    .C(_2863_),
    .Y(_2870_)
);

OAI21X1 _6523_ (
    .A(_2870_),
    .B(_2869_),
    .C(_2847_),
    .Y(_2871_)
);

NAND3X1 _6524_ (
    .A(_2852_),
    .B(_2868_),
    .C(_2871_),
    .Y(_2872_)
);

INVX1 _6525_ (
    .A(_2868_),
    .Y(_2873_)
);

INVX1 _6526_ (
    .A(_2849_),
    .Y(_2874_)
);

AOI22X1 _6527_ (
    .A(\z4.z3.z3.z1.s ),
    .B(_2874_),
    .C(_2867_),
    .D(_2864_),
    .Y(_2875_)
);

OAI21X1 _6528_ (
    .A(_2875_),
    .B(_2873_),
    .C(_2851_),
    .Y(_2876_)
);

AND2X2 _6529_ (
    .A(_2876_),
    .B(_2872_),
    .Y(\z4.q2 [4])
);

OAI21X1 _6530_ (
    .A(_2851_),
    .B(_2875_),
    .C(_2868_),
    .Y(_2877_)
);

OAI21X1 _6531_ (
    .A(_2859_),
    .B(_2860_),
    .C(_2864_),
    .Y(_2878_)
);

NAND2X1 _6532_ (
    .A(\z4.z3.z4.z1.s ),
    .B(\z4.z3.z3.z2.c ),
    .Y(_2879_)
);

OR2X2 _6533_ (
    .A(\z4.z3.z4.z1.s ),
    .B(\z4.z3.z3.z2.c ),
    .Y(_2880_)
);

NAND2X1 _6534_ (
    .A(_2879_),
    .B(_2880_),
    .Y(_2881_)
);

INVX1 _6535_ (
    .A(_2881_),
    .Y(_2882_)
);

NAND2X1 _6536_ (
    .A(\z4.z3.z2.z2.c ),
    .B(_2865_),
    .Y(_2883_)
);

INVX1 _6537_ (
    .A(\z4.z3.z2.z2.c ),
    .Y(_2884_)
);

NAND2X1 _6538_ (
    .A(_2884_),
    .B(_2855_),
    .Y(_2885_)
);

NAND3X1 _6539_ (
    .A(_2882_),
    .B(_2885_),
    .C(_2883_),
    .Y(_2886_)
);

NAND2X1 _6540_ (
    .A(\z4.z3.z2.z2.c ),
    .B(_2855_),
    .Y(_2887_)
);

NAND2X1 _6541_ (
    .A(_2884_),
    .B(_2865_),
    .Y(_2888_)
);

NAND3X1 _6542_ (
    .A(_2881_),
    .B(_2887_),
    .C(_2888_),
    .Y(_2889_)
);

NAND3X1 _6543_ (
    .A(_2878_),
    .B(_2886_),
    .C(_2889_),
    .Y(_2890_)
);

INVX1 _6544_ (
    .A(_2878_),
    .Y(_2891_)
);

AOI21X1 _6545_ (
    .A(_2888_),
    .B(_2887_),
    .C(_2881_),
    .Y(_2892_)
);

AOI21X1 _6546_ (
    .A(_2883_),
    .B(_2885_),
    .C(_2882_),
    .Y(_2893_)
);

OAI21X1 _6547_ (
    .A(_2892_),
    .B(_2893_),
    .C(_2891_),
    .Y(_2894_)
);

NAND2X1 _6548_ (
    .A(_2890_),
    .B(_2894_),
    .Y(_2895_)
);

NAND2X1 _6549_ (
    .A(_2877_),
    .B(_2895_),
    .Y(_2896_)
);

OR2X2 _6550_ (
    .A(_2895_),
    .B(_2877_),
    .Y(_2897_)
);

NAND2X1 _6551_ (
    .A(_2896_),
    .B(_2897_),
    .Y(\z4.q2 [5])
);

INVX1 _6552_ (
    .A(\z4.z3.z4.z2.s ),
    .Y(_2898_)
);

INVX1 _6553_ (
    .A(_2879_),
    .Y(_2899_)
);

OAI21X1 _6554_ (
    .A(_2899_),
    .B(_2892_),
    .C(_2898_),
    .Y(_2900_)
);

NAND3X1 _6555_ (
    .A(\z4.z3.z4.z2.s ),
    .B(_2879_),
    .C(_2886_),
    .Y(_2901_)
);

NAND2X1 _6556_ (
    .A(_2894_),
    .B(_2877_),
    .Y(_2902_)
);

AOI22X1 _6557_ (
    .A(_2900_),
    .B(_2901_),
    .C(_2902_),
    .D(_2890_),
    .Y(_2903_)
);

NAND2X1 _6558_ (
    .A(_2901_),
    .B(_2900_),
    .Y(_2904_)
);

NAND3X1 _6559_ (
    .A(_2868_),
    .B(_2890_),
    .C(_2872_),
    .Y(_2905_)
);

AOI21X1 _6560_ (
    .A(_2905_),
    .B(_2894_),
    .C(_2904_),
    .Y(_2906_)
);

NOR2X1 _6561_ (
    .A(_2903_),
    .B(_2906_),
    .Y(\z4.q2 [6])
);

OAI21X1 _6562_ (
    .A(_2899_),
    .B(_2892_),
    .C(\z4.z3.z4.z2.s ),
    .Y(_2825_)
);

NAND3X1 _6563_ (
    .A(_2894_),
    .B(_2904_),
    .C(_2905_),
    .Y(_2826_)
);

NAND3X1 _6564_ (
    .A(\z4.z3.z4.z2.c ),
    .B(_2825_),
    .C(_2826_),
    .Y(_2827_)
);

INVX1 _6565_ (
    .A(\z4.z3.z4.z2.c ),
    .Y(_2828_)
);

INVX1 _6566_ (
    .A(_2825_),
    .Y(_2829_)
);

OAI21X1 _6567_ (
    .A(_2829_),
    .B(_2903_),
    .C(_2828_),
    .Y(_2830_)
);

NAND2X1 _6568_ (
    .A(_2827_),
    .B(_2830_),
    .Y(\z4.q2 [7])
);

AOI21X1 _6569_ (
    .A(_2850_),
    .B(_2847_),
    .C(_2836_),
    .Y(_2831_)
);

NOR2X1 _6570_ (
    .A(_2831_),
    .B(_2852_),
    .Y(\z4.q2 [3])
);

AND2X2 _6571_ (
    .A(b[12]),
    .B(a[8]),
    .Y(\z4.q2 [0])
);

AND2X2 _6572_ (
    .A(b[12]),
    .B(a[9]),
    .Y(\z4.z3.z1.z1.a )
);

AND2X2 _6573_ (
    .A(a[8]),
    .B(b[13]),
    .Y(\z4.z3.z1.z1.b )
);

AND2X2 _6574_ (
    .A(a[9]),
    .B(b[13]),
    .Y(\z4.z3.z1.z2.a )
);

INVX1 _6575_ (
    .A(\z4.z3.z1.z1.b ),
    .Y(_2907_)
);

NAND2X1 _6576_ (
    .A(\z4.z3.z1.z1.a ),
    .B(_2907_),
    .Y(_2908_)
);

INVX1 _6577_ (
    .A(\z4.z3.z1.z1.a ),
    .Y(_2909_)
);

NAND2X1 _6578_ (
    .A(\z4.z3.z1.z1.b ),
    .B(_2909_),
    .Y(_2910_)
);

NAND2X1 _6579_ (
    .A(_2908_),
    .B(_2910_),
    .Y(\z4.z3.z1.z1.s )
);

NOR2X1 _6580_ (
    .A(_2907_),
    .B(_2909_),
    .Y(\z4.z3.z1.z1.c )
);

INVX1 _6581_ (
    .A(\z4.z3.z1.z1.c ),
    .Y(_2911_)
);

NAND2X1 _6582_ (
    .A(\z4.z3.z1.z2.a ),
    .B(_2911_),
    .Y(_2912_)
);

INVX1 _6583_ (
    .A(\z4.z3.z1.z2.a ),
    .Y(_2913_)
);

NAND2X1 _6584_ (
    .A(\z4.z3.z1.z1.c ),
    .B(_2913_),
    .Y(_2914_)
);

NAND2X1 _6585_ (
    .A(_2912_),
    .B(_2914_),
    .Y(\z4.z3.z1.z2.s )
);

NOR2X1 _6586_ (
    .A(_2911_),
    .B(_2913_),
    .Y(\z4.z3.z1.z2.c )
);

AND2X2 _6587_ (
    .A(b[12]),
    .B(a[10]),
    .Y(\z4.z3.q1 [0])
);

AND2X2 _6588_ (
    .A(b[12]),
    .B(a[11]),
    .Y(\z4.z3.z2.z1.a )
);

AND2X2 _6589_ (
    .A(a[10]),
    .B(b[13]),
    .Y(\z4.z3.z2.z1.b )
);

AND2X2 _6590_ (
    .A(a[11]),
    .B(b[13]),
    .Y(\z4.z3.z2.z2.a )
);

INVX1 _6591_ (
    .A(\z4.z3.z2.z1.b ),
    .Y(_2915_)
);

NAND2X1 _6592_ (
    .A(\z4.z3.z2.z1.a ),
    .B(_2915_),
    .Y(_2916_)
);

INVX1 _6593_ (
    .A(\z4.z3.z2.z1.a ),
    .Y(_2917_)
);

NAND2X1 _6594_ (
    .A(\z4.z3.z2.z1.b ),
    .B(_2917_),
    .Y(_2918_)
);

NAND2X1 _6595_ (
    .A(_2916_),
    .B(_2918_),
    .Y(\z4.z3.z2.z1.s )
);

NOR2X1 _6596_ (
    .A(_2915_),
    .B(_2917_),
    .Y(\z4.z3.z2.z1.c )
);

INVX1 _6597_ (
    .A(\z4.z3.z2.z1.c ),
    .Y(_2919_)
);

NAND2X1 _6598_ (
    .A(\z4.z3.z2.z2.a ),
    .B(_2919_),
    .Y(_2920_)
);

INVX1 _6599_ (
    .A(\z4.z3.z2.z2.a ),
    .Y(_2921_)
);

NAND2X1 _6600_ (
    .A(\z4.z3.z2.z1.c ),
    .B(_2921_),
    .Y(_2922_)
);

NAND2X1 _6601_ (
    .A(_2920_),
    .B(_2922_),
    .Y(\z4.z3.z2.z2.s )
);

NOR2X1 _6602_ (
    .A(_2919_),
    .B(_2921_),
    .Y(\z4.z3.z2.z2.c )
);

AND2X2 _6603_ (
    .A(b[14]),
    .B(a[8]),
    .Y(\z4.z3.q2 [0])
);

AND2X2 _6604_ (
    .A(b[14]),
    .B(a[9]),
    .Y(\z4.z3.z3.z1.a )
);

AND2X2 _6605_ (
    .A(a[8]),
    .B(b[15]),
    .Y(\z4.z3.z3.z1.b )
);

AND2X2 _6606_ (
    .A(a[9]),
    .B(b[15]),
    .Y(\z4.z3.z3.z2.a )
);

INVX1 _6607_ (
    .A(\z4.z3.z3.z1.b ),
    .Y(_2923_)
);

NAND2X1 _6608_ (
    .A(\z4.z3.z3.z1.a ),
    .B(_2923_),
    .Y(_2924_)
);

INVX1 _6609_ (
    .A(\z4.z3.z3.z1.a ),
    .Y(_2925_)
);

NAND2X1 _6610_ (
    .A(\z4.z3.z3.z1.b ),
    .B(_2925_),
    .Y(_2926_)
);

NAND2X1 _6611_ (
    .A(_2924_),
    .B(_2926_),
    .Y(\z4.z3.z3.z1.s )
);

NOR2X1 _6612_ (
    .A(_2923_),
    .B(_2925_),
    .Y(\z4.z3.z3.z1.c )
);

INVX1 _6613_ (
    .A(\z4.z3.z3.z1.c ),
    .Y(_2927_)
);

NAND2X1 _6614_ (
    .A(\z4.z3.z3.z2.a ),
    .B(_2927_),
    .Y(_2928_)
);

INVX1 _6615_ (
    .A(\z4.z3.z3.z2.a ),
    .Y(_2929_)
);

NAND2X1 _6616_ (
    .A(\z4.z3.z3.z1.c ),
    .B(_2929_),
    .Y(_2930_)
);

NAND2X1 _6617_ (
    .A(_2928_),
    .B(_2930_),
    .Y(\z4.z3.z3.z2.s )
);

NOR2X1 _6618_ (
    .A(_2927_),
    .B(_2929_),
    .Y(\z4.z3.z3.z2.c )
);

AND2X2 _6619_ (
    .A(b[14]),
    .B(a[10]),
    .Y(\z4.z3.q3 [0])
);

AND2X2 _6620_ (
    .A(b[14]),
    .B(a[11]),
    .Y(\z4.z3.z4.z1.a )
);

AND2X2 _6621_ (
    .A(a[10]),
    .B(b[15]),
    .Y(\z4.z3.z4.z1.b )
);

AND2X2 _6622_ (
    .A(a[11]),
    .B(b[15]),
    .Y(\z4.z3.z4.z2.a )
);

INVX1 _6623_ (
    .A(\z4.z3.z4.z1.b ),
    .Y(_2931_)
);

NAND2X1 _6624_ (
    .A(\z4.z3.z4.z1.a ),
    .B(_2931_),
    .Y(_2932_)
);

INVX1 _6625_ (
    .A(\z4.z3.z4.z1.a ),
    .Y(_2933_)
);

NAND2X1 _6626_ (
    .A(\z4.z3.z4.z1.b ),
    .B(_2933_),
    .Y(_2934_)
);

NAND2X1 _6627_ (
    .A(_2932_),
    .B(_2934_),
    .Y(\z4.z3.z4.z1.s )
);

NOR2X1 _6628_ (
    .A(_2931_),
    .B(_2933_),
    .Y(\z4.z3.z4.z1.c )
);

INVX1 _6629_ (
    .A(\z4.z3.z4.z1.c ),
    .Y(_2935_)
);

NAND2X1 _6630_ (
    .A(\z4.z3.z4.z2.a ),
    .B(_2935_),
    .Y(_2936_)
);

INVX1 _6631_ (
    .A(\z4.z3.z4.z2.a ),
    .Y(_2937_)
);

NAND2X1 _6632_ (
    .A(\z4.z3.z4.z1.c ),
    .B(_2937_),
    .Y(_2938_)
);

NAND2X1 _6633_ (
    .A(_2936_),
    .B(_2938_),
    .Y(\z4.z3.z4.z2.s )
);

NOR2X1 _6634_ (
    .A(_2935_),
    .B(_2937_),
    .Y(\z4.z3.z4.z2.c )
);

NOR2X1 _6635_ (
    .A(\z4.z4.q1 [0]),
    .B(\z4.z4.z1.z2.s ),
    .Y(_2946_)
);

AND2X2 _6636_ (
    .A(\z4.z4.q1 [0]),
    .B(\z4.z4.z1.z2.s ),
    .Y(_2947_)
);

NOR2X1 _6637_ (
    .A(_2946_),
    .B(_2947_),
    .Y(_2948_)
);

NAND2X1 _6638_ (
    .A(\z4.z4.q2 [0]),
    .B(_2948_),
    .Y(_2949_)
);

INVX1 _6639_ (
    .A(_2949_),
    .Y(_2950_)
);

NOR2X1 _6640_ (
    .A(\z4.z4.q2 [0]),
    .B(_2948_),
    .Y(_2951_)
);

NOR2X1 _6641_ (
    .A(_2951_),
    .B(_2950_),
    .Y(\z4.q3 [2])
);

NAND2X1 _6642_ (
    .A(\z4.z4.q1 [0]),
    .B(\z4.z4.z1.z2.s ),
    .Y(_2952_)
);

NOR2X1 _6643_ (
    .A(\z4.z4.z2.z1.s ),
    .B(\z4.z4.z1.z2.c ),
    .Y(_2953_)
);

NAND2X1 _6644_ (
    .A(\z4.z4.z2.z1.s ),
    .B(\z4.z4.z1.z2.c ),
    .Y(_2954_)
);

INVX1 _6645_ (
    .A(_2954_),
    .Y(_2955_)
);

OAI21X1 _6646_ (
    .A(_2953_),
    .B(_2955_),
    .C(_2952_),
    .Y(_2956_)
);

INVX1 _6647_ (
    .A(\z4.z4.z2.z1.s ),
    .Y(_2957_)
);

INVX1 _6648_ (
    .A(\z4.z4.z1.z2.c ),
    .Y(_2958_)
);

NAND2X1 _6649_ (
    .A(_2957_),
    .B(_2958_),
    .Y(_2959_)
);

NAND3X1 _6650_ (
    .A(_2947_),
    .B(_2954_),
    .C(_2959_),
    .Y(_2960_)
);

NAND3X1 _6651_ (
    .A(\z4.z4.z3.z1.s ),
    .B(_2960_),
    .C(_2956_),
    .Y(_2961_)
);

INVX1 _6652_ (
    .A(\z4.z4.z3.z1.s ),
    .Y(_2962_)
);

NAND2X1 _6653_ (
    .A(_2960_),
    .B(_2956_),
    .Y(_2963_)
);

NAND2X1 _6654_ (
    .A(_2962_),
    .B(_2963_),
    .Y(_2964_)
);

NAND3X1 _6655_ (
    .A(_2950_),
    .B(_2961_),
    .C(_2964_),
    .Y(_2965_)
);

INVX1 _6656_ (
    .A(_2965_),
    .Y(_2966_)
);

INVX1 _6657_ (
    .A(_2961_),
    .Y(_2967_)
);

OAI21X1 _6658_ (
    .A(_2952_),
    .B(_2953_),
    .C(_2954_),
    .Y(_2968_)
);

NAND2X1 _6659_ (
    .A(\z4.z4.z2.z2.s ),
    .B(_2968_),
    .Y(_2969_)
);

INVX1 _6660_ (
    .A(\z4.z4.z2.z2.s ),
    .Y(_2970_)
);

NAND3X1 _6661_ (
    .A(_2970_),
    .B(_2954_),
    .C(_2960_),
    .Y(_2971_)
);

NAND2X1 _6662_ (
    .A(\z4.z4.q3 [0]),
    .B(\z4.z4.z3.z2.s ),
    .Y(_2972_)
);

INVX1 _6663_ (
    .A(\z4.z4.q3 [0]),
    .Y(_2973_)
);

INVX1 _6664_ (
    .A(\z4.z4.z3.z2.s ),
    .Y(_2974_)
);

NAND2X1 _6665_ (
    .A(_2973_),
    .B(_2974_),
    .Y(_2975_)
);

NAND2X1 _6666_ (
    .A(_2972_),
    .B(_2975_),
    .Y(_2976_)
);

INVX1 _6667_ (
    .A(_2976_),
    .Y(_2977_)
);

NAND3X1 _6668_ (
    .A(_2969_),
    .B(_2977_),
    .C(_2971_),
    .Y(_2978_)
);

AND2X2 _6669_ (
    .A(_2968_),
    .B(\z4.z4.z2.z2.s ),
    .Y(_2979_)
);

NOR2X1 _6670_ (
    .A(\z4.z4.z2.z2.s ),
    .B(_2968_),
    .Y(_2980_)
);

OAI21X1 _6671_ (
    .A(_2980_),
    .B(_2979_),
    .C(_2976_),
    .Y(_2981_)
);

NAND3X1 _6672_ (
    .A(_2967_),
    .B(_2978_),
    .C(_2981_),
    .Y(_2982_)
);

INVX1 _6673_ (
    .A(_2978_),
    .Y(_2983_)
);

AOI21X1 _6674_ (
    .A(_2971_),
    .B(_2969_),
    .C(_2977_),
    .Y(_2984_)
);

OAI21X1 _6675_ (
    .A(_2984_),
    .B(_2983_),
    .C(_2961_),
    .Y(_2985_)
);

NAND3X1 _6676_ (
    .A(_2966_),
    .B(_2982_),
    .C(_2985_),
    .Y(_2986_)
);

INVX1 _6677_ (
    .A(_2982_),
    .Y(_2987_)
);

INVX1 _6678_ (
    .A(_2963_),
    .Y(_2988_)
);

AOI22X1 _6679_ (
    .A(\z4.z4.z3.z1.s ),
    .B(_2988_),
    .C(_2981_),
    .D(_2978_),
    .Y(_2989_)
);

OAI21X1 _6680_ (
    .A(_2989_),
    .B(_2987_),
    .C(_2965_),
    .Y(_2990_)
);

AND2X2 _6681_ (
    .A(_2990_),
    .B(_2986_),
    .Y(\z4.q3 [4])
);

OAI21X1 _6682_ (
    .A(_2965_),
    .B(_2989_),
    .C(_2982_),
    .Y(_2991_)
);

OAI21X1 _6683_ (
    .A(_2973_),
    .B(_2974_),
    .C(_2978_),
    .Y(_2992_)
);

NAND2X1 _6684_ (
    .A(\z4.z4.z4.z1.s ),
    .B(\z4.z4.z3.z2.c ),
    .Y(_2993_)
);

OR2X2 _6685_ (
    .A(\z4.z4.z4.z1.s ),
    .B(\z4.z4.z3.z2.c ),
    .Y(_2994_)
);

NAND2X1 _6686_ (
    .A(_2993_),
    .B(_2994_),
    .Y(_2995_)
);

INVX1 _6687_ (
    .A(_2995_),
    .Y(_2996_)
);

NAND2X1 _6688_ (
    .A(\z4.z4.z2.z2.c ),
    .B(_2979_),
    .Y(_2997_)
);

INVX1 _6689_ (
    .A(\z4.z4.z2.z2.c ),
    .Y(_2998_)
);

NAND2X1 _6690_ (
    .A(_2998_),
    .B(_2969_),
    .Y(_2999_)
);

NAND3X1 _6691_ (
    .A(_2996_),
    .B(_2999_),
    .C(_2997_),
    .Y(_3000_)
);

NAND2X1 _6692_ (
    .A(\z4.z4.z2.z2.c ),
    .B(_2969_),
    .Y(_3001_)
);

NAND2X1 _6693_ (
    .A(_2998_),
    .B(_2979_),
    .Y(_3002_)
);

NAND3X1 _6694_ (
    .A(_2995_),
    .B(_3001_),
    .C(_3002_),
    .Y(_3003_)
);

NAND3X1 _6695_ (
    .A(_2992_),
    .B(_3000_),
    .C(_3003_),
    .Y(_3004_)
);

INVX1 _6696_ (
    .A(_2992_),
    .Y(_3005_)
);

AOI21X1 _6697_ (
    .A(_3002_),
    .B(_3001_),
    .C(_2995_),
    .Y(_3006_)
);

AOI21X1 _6698_ (
    .A(_2997_),
    .B(_2999_),
    .C(_2996_),
    .Y(_3007_)
);

OAI21X1 _6699_ (
    .A(_3006_),
    .B(_3007_),
    .C(_3005_),
    .Y(_3008_)
);

NAND2X1 _6700_ (
    .A(_3004_),
    .B(_3008_),
    .Y(_3009_)
);

NAND2X1 _6701_ (
    .A(_2991_),
    .B(_3009_),
    .Y(_3010_)
);

OR2X2 _6702_ (
    .A(_3009_),
    .B(_2991_),
    .Y(_3011_)
);

NAND2X1 _6703_ (
    .A(_3010_),
    .B(_3011_),
    .Y(\z4.q3 [5])
);

INVX1 _6704_ (
    .A(\z4.z4.z4.z2.s ),
    .Y(_3012_)
);

INVX1 _6705_ (
    .A(_2993_),
    .Y(_3013_)
);

OAI21X1 _6706_ (
    .A(_3013_),
    .B(_3006_),
    .C(_3012_),
    .Y(_3014_)
);

NAND3X1 _6707_ (
    .A(\z4.z4.z4.z2.s ),
    .B(_2993_),
    .C(_3000_),
    .Y(_3015_)
);

NAND2X1 _6708_ (
    .A(_3008_),
    .B(_2991_),
    .Y(_3016_)
);

AOI22X1 _6709_ (
    .A(_3014_),
    .B(_3015_),
    .C(_3016_),
    .D(_3004_),
    .Y(_3017_)
);

NAND2X1 _6710_ (
    .A(_3015_),
    .B(_3014_),
    .Y(_3018_)
);

NAND3X1 _6711_ (
    .A(_2982_),
    .B(_3004_),
    .C(_2986_),
    .Y(_3019_)
);

AOI21X1 _6712_ (
    .A(_3019_),
    .B(_3008_),
    .C(_3018_),
    .Y(_3020_)
);

NOR2X1 _6713_ (
    .A(_3017_),
    .B(_3020_),
    .Y(\z4.q3 [6])
);

OAI21X1 _6714_ (
    .A(_3013_),
    .B(_3006_),
    .C(\z4.z4.z4.z2.s ),
    .Y(_2939_)
);

NAND3X1 _6715_ (
    .A(_3008_),
    .B(_3018_),
    .C(_3019_),
    .Y(_2940_)
);

NAND3X1 _6716_ (
    .A(\z4.z4.z4.z2.c ),
    .B(_2939_),
    .C(_2940_),
    .Y(_2941_)
);

INVX1 _6717_ (
    .A(\z4.z4.z4.z2.c ),
    .Y(_2942_)
);

INVX1 _6718_ (
    .A(_2939_),
    .Y(_2943_)
);

OAI21X1 _6719_ (
    .A(_2943_),
    .B(_3017_),
    .C(_2942_),
    .Y(_2944_)
);

NAND2X1 _6720_ (
    .A(_2941_),
    .B(_2944_),
    .Y(\z4.q3 [7])
);

AOI21X1 _6721_ (
    .A(_2964_),
    .B(_2961_),
    .C(_2950_),
    .Y(_2945_)
);

NOR2X1 _6722_ (
    .A(_2945_),
    .B(_2966_),
    .Y(\z4.q3 [3])
);

AND2X2 _6723_ (
    .A(b[12]),
    .B(a[12]),
    .Y(\z4.q3 [0])
);

AND2X2 _6724_ (
    .A(b[12]),
    .B(a[13]),
    .Y(\z4.z4.z1.z1.a )
);

AND2X2 _6725_ (
    .A(a[12]),
    .B(b[13]),
    .Y(\z4.z4.z1.z1.b )
);

AND2X2 _6726_ (
    .A(a[13]),
    .B(b[13]),
    .Y(\z4.z4.z1.z2.a )
);

INVX1 _6727_ (
    .A(\z4.z4.z1.z1.b ),
    .Y(_3021_)
);

NAND2X1 _6728_ (
    .A(\z4.z4.z1.z1.a ),
    .B(_3021_),
    .Y(_3022_)
);

INVX1 _6729_ (
    .A(\z4.z4.z1.z1.a ),
    .Y(_3023_)
);

NAND2X1 _6730_ (
    .A(\z4.z4.z1.z1.b ),
    .B(_3023_),
    .Y(_3024_)
);

NAND2X1 _6731_ (
    .A(_3022_),
    .B(_3024_),
    .Y(\z4.z4.z1.z1.s )
);

NOR2X1 _6732_ (
    .A(_3021_),
    .B(_3023_),
    .Y(\z4.z4.z1.z1.c )
);

INVX1 _6733_ (
    .A(\z4.z4.z1.z1.c ),
    .Y(_3025_)
);

NAND2X1 _6734_ (
    .A(\z4.z4.z1.z2.a ),
    .B(_3025_),
    .Y(_3026_)
);

INVX1 _6735_ (
    .A(\z4.z4.z1.z2.a ),
    .Y(_3027_)
);

NAND2X1 _6736_ (
    .A(\z4.z4.z1.z1.c ),
    .B(_3027_),
    .Y(_3028_)
);

NAND2X1 _6737_ (
    .A(_3026_),
    .B(_3028_),
    .Y(\z4.z4.z1.z2.s )
);

NOR2X1 _6738_ (
    .A(_3025_),
    .B(_3027_),
    .Y(\z4.z4.z1.z2.c )
);

AND2X2 _6739_ (
    .A(b[12]),
    .B(a[14]),
    .Y(\z4.z4.q1 [0])
);

AND2X2 _6740_ (
    .A(b[12]),
    .B(a[15]),
    .Y(\z4.z4.z2.z1.a )
);

AND2X2 _6741_ (
    .A(a[14]),
    .B(b[13]),
    .Y(\z4.z4.z2.z1.b )
);

AND2X2 _6742_ (
    .A(a[15]),
    .B(b[13]),
    .Y(\z4.z4.z2.z2.a )
);

INVX1 _6743_ (
    .A(\z4.z4.z2.z1.b ),
    .Y(_3029_)
);

NAND2X1 _6744_ (
    .A(\z4.z4.z2.z1.a ),
    .B(_3029_),
    .Y(_3030_)
);

INVX1 _6745_ (
    .A(\z4.z4.z2.z1.a ),
    .Y(_3031_)
);

NAND2X1 _6746_ (
    .A(\z4.z4.z2.z1.b ),
    .B(_3031_),
    .Y(_3032_)
);

NAND2X1 _6747_ (
    .A(_3030_),
    .B(_3032_),
    .Y(\z4.z4.z2.z1.s )
);

NOR2X1 _6748_ (
    .A(_3029_),
    .B(_3031_),
    .Y(\z4.z4.z2.z1.c )
);

INVX1 _6749_ (
    .A(\z4.z4.z2.z1.c ),
    .Y(_3033_)
);

NAND2X1 _6750_ (
    .A(\z4.z4.z2.z2.a ),
    .B(_3033_),
    .Y(_3034_)
);

INVX1 _6751_ (
    .A(\z4.z4.z2.z2.a ),
    .Y(_3035_)
);

NAND2X1 _6752_ (
    .A(\z4.z4.z2.z1.c ),
    .B(_3035_),
    .Y(_3036_)
);

NAND2X1 _6753_ (
    .A(_3034_),
    .B(_3036_),
    .Y(\z4.z4.z2.z2.s )
);

NOR2X1 _6754_ (
    .A(_3033_),
    .B(_3035_),
    .Y(\z4.z4.z2.z2.c )
);

AND2X2 _6755_ (
    .A(b[14]),
    .B(a[12]),
    .Y(\z4.z4.q2 [0])
);

AND2X2 _6756_ (
    .A(b[14]),
    .B(a[13]),
    .Y(\z4.z4.z3.z1.a )
);

AND2X2 _6757_ (
    .A(a[12]),
    .B(b[15]),
    .Y(\z4.z4.z3.z1.b )
);

AND2X2 _6758_ (
    .A(a[13]),
    .B(b[15]),
    .Y(\z4.z4.z3.z2.a )
);

INVX1 _6759_ (
    .A(\z4.z4.z3.z1.b ),
    .Y(_3037_)
);

NAND2X1 _6760_ (
    .A(\z4.z4.z3.z1.a ),
    .B(_3037_),
    .Y(_3038_)
);

INVX1 _6761_ (
    .A(\z4.z4.z3.z1.a ),
    .Y(_3039_)
);

NAND2X1 _6762_ (
    .A(\z4.z4.z3.z1.b ),
    .B(_3039_),
    .Y(_3040_)
);

NAND2X1 _6763_ (
    .A(_3038_),
    .B(_3040_),
    .Y(\z4.z4.z3.z1.s )
);

NOR2X1 _6764_ (
    .A(_3037_),
    .B(_3039_),
    .Y(\z4.z4.z3.z1.c )
);

INVX1 _6765_ (
    .A(\z4.z4.z3.z1.c ),
    .Y(_3041_)
);

NAND2X1 _6766_ (
    .A(\z4.z4.z3.z2.a ),
    .B(_3041_),
    .Y(_3042_)
);

INVX1 _6767_ (
    .A(\z4.z4.z3.z2.a ),
    .Y(_3043_)
);

NAND2X1 _6768_ (
    .A(\z4.z4.z3.z1.c ),
    .B(_3043_),
    .Y(_3044_)
);

NAND2X1 _6769_ (
    .A(_3042_),
    .B(_3044_),
    .Y(\z4.z4.z3.z2.s )
);

NOR2X1 _6770_ (
    .A(_3041_),
    .B(_3043_),
    .Y(\z4.z4.z3.z2.c )
);

AND2X2 _6771_ (
    .A(b[14]),
    .B(a[14]),
    .Y(\z4.z4.q3 [0])
);

AND2X2 _6772_ (
    .A(b[14]),
    .B(a[15]),
    .Y(\z4.z4.z4.z1.a )
);

AND2X2 _6773_ (
    .A(a[14]),
    .B(b[15]),
    .Y(\z4.z4.z4.z1.b )
);

AND2X2 _6774_ (
    .A(a[15]),
    .B(b[15]),
    .Y(\z4.z4.z4.z2.a )
);

INVX1 _6775_ (
    .A(\z4.z4.z4.z1.b ),
    .Y(_3045_)
);

NAND2X1 _6776_ (
    .A(\z4.z4.z4.z1.a ),
    .B(_3045_),
    .Y(_3046_)
);

INVX1 _6777_ (
    .A(\z4.z4.z4.z1.a ),
    .Y(_3047_)
);

NAND2X1 _6778_ (
    .A(\z4.z4.z4.z1.b ),
    .B(_3047_),
    .Y(_3048_)
);

NAND2X1 _6779_ (
    .A(_3046_),
    .B(_3048_),
    .Y(\z4.z4.z4.z1.s )
);

NOR2X1 _6780_ (
    .A(_3045_),
    .B(_3047_),
    .Y(\z4.z4.z4.z1.c )
);

INVX1 _6781_ (
    .A(\z4.z4.z4.z1.c ),
    .Y(_3049_)
);

NAND2X1 _6782_ (
    .A(\z4.z4.z4.z2.a ),
    .B(_3049_),
    .Y(_3050_)
);

INVX1 _6783_ (
    .A(\z4.z4.z4.z2.a ),
    .Y(_3051_)
);

NAND2X1 _6784_ (
    .A(\z4.z4.z4.z1.c ),
    .B(_3051_),
    .Y(_3052_)
);

NAND2X1 _6785_ (
    .A(_3050_),
    .B(_3052_),
    .Y(\z4.z4.z4.z2.s )
);

NOR2X1 _6786_ (
    .A(_3049_),
    .B(_3051_),
    .Y(\z4.z4.z4.z2.c )
);

BUFX2 _6787_ (
    .A(q0[0]),
    .Y(c[0])
);

BUFX2 _6788_ (
    .A(\z1.z1.z1.z1.s ),
    .Y(c[1])
);

BUFX2 _6789_ (
    .A(_3053_[10]),
    .Y(c[10])
);

BUFX2 _6790_ (
    .A(_3053_[11]),
    .Y(c[11])
);

BUFX2 _6791_ (
    .A(_3053_[12]),
    .Y(c[12])
);

BUFX2 _6792_ (
    .A(_3053_[13]),
    .Y(c[13])
);

BUFX2 _6793_ (
    .A(_3053_[14]),
    .Y(c[14])
);

BUFX2 _6794_ (
    .A(_3053_[15]),
    .Y(c[15])
);

BUFX2 _6795_ (
    .A(_3053_[16]),
    .Y(c[16])
);

BUFX2 _6796_ (
    .A(_3053_[17]),
    .Y(c[17])
);

BUFX2 _6797_ (
    .A(_3053_[18]),
    .Y(c[18])
);

BUFX2 _6798_ (
    .A(_3053_[19]),
    .Y(c[19])
);

BUFX2 _6799_ (
    .A(q0[2]),
    .Y(c[2])
);

BUFX2 _6800_ (
    .A(_3053_[20]),
    .Y(c[20])
);

BUFX2 _6801_ (
    .A(_3053_[21]),
    .Y(c[21])
);

BUFX2 _6802_ (
    .A(_3053_[22]),
    .Y(c[22])
);

BUFX2 _6803_ (
    .A(_3053_[23]),
    .Y(c[23])
);

BUFX2 _6804_ (
    .A(_3053_[24]),
    .Y(c[24])
);

BUFX2 _6805_ (
    .A(_3053_[25]),
    .Y(c[25])
);

BUFX2 _6806_ (
    .A(_3053_[26]),
    .Y(c[26])
);

BUFX2 _6807_ (
    .A(_3053_[27]),
    .Y(c[27])
);

BUFX2 _6808_ (
    .A(_3053_[28]),
    .Y(c[28])
);

BUFX2 _6809_ (
    .A(_3053_[29]),
    .Y(c[29])
);

BUFX2 _6810_ (
    .A(q0[3]),
    .Y(c[3])
);

BUFX2 _6811_ (
    .A(_3053_[30]),
    .Y(c[30])
);

BUFX2 _6812_ (
    .A(_3053_[31]),
    .Y(c[31])
);

BUFX2 _6813_ (
    .A(q0[4]),
    .Y(c[4])
);

BUFX2 _6814_ (
    .A(q0[5]),
    .Y(c[5])
);

BUFX2 _6815_ (
    .A(q0[6]),
    .Y(c[6])
);

BUFX2 _6816_ (
    .A(q0[7]),
    .Y(c[7])
);

BUFX2 _6817_ (
    .A(_3053_[8]),
    .Y(c[8])
);

BUFX2 _6818_ (
    .A(_3053_[9]),
    .Y(c[9])
);

endmodule
