magic
tech scmos
magscale 1 3
timestamp 1555596690
<< checkpaint >>
rect -56 -56 84 354
<< genericcontact >>
rect 11 272 17 278
rect 11 244 17 250
rect 11 216 17 222
rect 11 188 17 194
rect 11 160 17 166
rect 11 132 17 138
rect 11 104 17 110
rect 11 76 17 82
rect 11 48 17 54
rect 11 20 17 26
<< metal1 >>
rect 4 4 24 294
<< end >>
