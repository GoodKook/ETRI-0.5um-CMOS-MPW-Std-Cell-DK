//
// Apple-1 KBD & DSP IO Address
//

`define PIA_KBD_REG     16'hD010
`define PIA_KBD_CTL     16'hD011

`define PIA_DSP_REG     16'hD012
`define PIA_DSP_CTL     16'hD013
