magic
tech scmos
magscale 1 2
timestamp 1726842657
<< nwell >>
rect -13 154 213 272
<< ntransistor >>
rect 20 14 24 54
rect 28 14 32 54
rect 72 14 76 34
rect 92 14 96 54
rect 112 14 116 54
rect 132 14 136 54
rect 176 14 180 34
<< ptransistor >>
rect 20 206 24 246
rect 40 206 44 246
rect 84 206 88 246
rect 104 206 108 246
rect 124 166 128 246
rect 132 166 136 246
rect 152 206 156 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 14 28 54
rect 32 14 34 54
rect 81 34 92 54
rect 62 33 72 34
rect 70 14 72 33
rect 76 14 78 34
rect 90 14 92 34
rect 96 14 98 54
rect 110 14 112 54
rect 116 26 118 54
rect 130 26 132 54
rect 116 14 132 26
rect 136 50 150 54
rect 136 18 138 50
rect 136 14 150 18
rect 174 14 176 34
rect 180 14 182 34
<< pdiffusion >>
rect 18 206 20 246
rect 24 214 26 246
rect 38 214 40 246
rect 24 206 40 214
rect 44 206 46 246
rect 82 206 84 246
rect 88 206 90 246
rect 102 206 104 246
rect 108 206 110 246
rect 122 166 124 246
rect 128 166 132 246
rect 136 206 138 246
rect 150 206 152 246
rect 156 206 158 246
rect 136 166 145 206
<< ndcontact >>
rect 6 14 18 54
rect 34 14 46 54
rect 58 14 70 33
rect 78 14 90 34
rect 98 14 110 54
rect 118 26 130 54
rect 138 18 150 50
rect 162 14 174 34
rect 182 14 194 34
<< pdcontact >>
rect 6 206 18 246
rect 26 214 38 246
rect 46 206 58 246
rect 70 206 82 246
rect 90 206 102 246
rect 110 166 122 246
rect 138 206 150 246
rect 158 206 170 246
<< psubstratepcontact >>
rect -6 -6 206 6
<< nsubstratencontact >>
rect -6 254 206 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 84 246 88 250
rect 104 246 108 250
rect 124 246 128 250
rect 132 246 136 250
rect 152 246 156 250
rect 20 116 24 206
rect 20 54 24 103
rect 40 99 44 206
rect 84 202 88 206
rect 104 202 108 206
rect 84 198 108 202
rect 40 68 44 87
rect 28 63 44 68
rect 84 66 88 198
rect 124 162 128 166
rect 112 158 128 162
rect 112 103 116 158
rect 28 54 32 63
rect 77 60 96 66
rect 92 54 96 60
rect 112 54 116 91
rect 132 83 136 166
rect 152 71 156 206
rect 132 54 136 71
rect 156 59 180 63
rect 72 34 76 54
rect 176 34 180 59
rect 20 10 24 14
rect 28 10 32 14
rect 72 10 76 14
rect 92 10 96 14
rect 112 10 116 14
rect 132 10 136 14
rect 176 10 180 14
<< polycontact >>
rect 17 103 29 116
rect 40 87 52 99
rect 104 91 116 103
rect 65 54 77 66
rect 124 71 136 83
rect 144 59 156 71
<< metal1 >>
rect -6 266 206 268
rect -6 252 206 254
rect 26 246 38 252
rect 90 246 102 252
rect 138 246 150 252
rect 26 210 38 214
rect 8 204 18 206
rect 46 204 54 206
rect 8 198 54 204
rect 47 119 54 198
rect 70 117 77 206
rect 111 153 117 166
rect 111 147 133 153
rect 19 81 28 103
rect 52 91 104 97
rect 124 95 133 147
rect 158 117 164 206
rect 157 103 164 117
rect 124 89 148 95
rect 19 74 124 81
rect 142 71 148 89
rect 158 83 164 103
rect 158 77 188 83
rect 34 54 43 68
rect 57 54 65 66
rect 142 65 144 71
rect 119 59 144 65
rect 119 54 131 59
rect 58 33 72 34
rect 110 18 138 20
rect 182 34 188 77
rect 110 14 150 18
rect 6 8 18 14
rect 78 8 90 14
rect 162 8 174 14
rect -6 6 206 8
rect -6 -8 206 -6
<< m2contact >>
rect 3 103 17 117
rect 43 105 57 119
rect 63 103 77 117
rect 103 103 117 117
rect 143 103 157 117
rect 43 54 57 68
rect 58 34 72 48
<< metal2 >>
rect 66 117 74 134
rect 106 117 114 134
rect 6 86 14 103
rect 46 68 53 105
rect 68 48 76 103
rect 146 86 154 103
rect 72 34 76 48
<< m1p >>
rect -6 252 206 268
rect -6 -8 206 8
<< m2p >>
rect 66 119 74 134
rect 106 119 114 134
rect 6 86 14 101
rect 146 86 154 101
<< labels >>
rlabel metal2 10 90 10 90 7 A
port 1 n signal input
rlabel metal2 110 131 110 131 3 B
port 2 n signal input
rlabel metal2 150 90 150 90 3 YS
port 3 n signal output
rlabel metal2 70 131 70 131 7 YC
port 4 n signal output
rlabel metal1 -6 252 206 268 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -6 -8 206 8 0 gnd
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 200 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
