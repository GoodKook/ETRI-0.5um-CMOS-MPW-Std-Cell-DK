magic
tech scmos
magscale 1 2
timestamp 1701862152
<< checkpaint >>
rect -34 157 54 159
rect -34 78 94 157
rect -14 46 94 78
<< nwell >>
rect -12 154 72 272
<< ntransistor >>
rect 18 14 22 54
rect 38 14 42 54
<< ptransistor >>
rect 18 166 22 246
rect 38 166 42 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 14 24 54
rect 36 14 38 54
rect 42 14 44 54
<< pdiffusion >>
rect 4 244 18 246
rect 16 166 18 244
rect 22 166 24 246
rect 36 166 38 246
rect 42 166 44 246
<< ndcontact >>
rect 4 14 16 54
rect 24 14 36 54
rect 44 14 56 54
<< pdcontact >>
rect 4 166 16 244
rect 24 166 36 246
rect 44 166 56 246
<< psubstratepcontact >>
rect -6 -6 66 6
<< nsubstratencontact >>
rect -6 254 66 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 18 164 22 166
rect 38 164 42 166
rect 18 160 42 164
rect 18 62 22 160
rect 18 58 42 62
rect 18 54 22 58
rect 38 54 42 58
rect 18 10 22 14
rect 38 10 42 14
<< polycontact >>
rect 6 91 18 103
<< metal1 >>
rect -6 266 66 268
rect -6 252 66 254
rect 4 244 16 252
rect 44 246 56 252
rect 26 117 33 166
rect 26 103 40 117
rect 26 54 33 103
rect 4 8 16 14
rect 44 8 56 14
rect -6 6 66 8
rect -6 -8 66 -6
<< m2contact >>
rect 6 103 20 117
rect 40 103 54 117
<< metal2 >>
rect 6 117 14 134
rect 46 86 54 103
<< m1p >>
rect -6 252 66 268
rect -6 -8 66 8
<< m2p >>
rect 6 119 14 134
rect 46 86 54 101
<< labels >>
rlabel metal2 10 130 10 130 1 A
port 1 n signal input
rlabel metal2 50 88 50 88 1 Y
port 2 n signal output
rlabel metal1 -6 252 66 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -6 -8 66 8 0 gnd
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 60 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
