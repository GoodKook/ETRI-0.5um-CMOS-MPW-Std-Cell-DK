magic
tech scmos
magscale 1 30
timestamp 1725865881
<< checkpaint >>
rect -510 34810 5760 34880
rect 10530 34810 12360 35120
rect -1035 34705 12735 34810
rect -1035 19580 13695 34705
rect -1085 16505 13695 19580
rect -1035 8550 13695 16505
rect -510 8460 13695 8550
rect 1250 8445 13695 8460
rect 1250 8350 12430 8445
rect 1250 7900 10953 8350
<< nwell >>
rect 0 30150 12195 32010
rect 0 20350 12200 28350
rect 100 9150 12100 16950
<< psubstratepdiff >>
rect 100 32550 12100 34210
<< nsubstratendiff >>
rect 100 30250 12100 31910
rect 100 20450 12100 28250
rect 100 9150 12100 16950
<< metal1 >>
rect 100 32550 12100 34210
rect 100 30250 12100 31910
rect 100 20450 12100 28250
rect 100 9150 12100 16950
rect 1850 8250 10350 8500
rect 1850 250 2100 8250
rect 2200 8090 2400 8150
rect 2200 8010 2260 8090
rect 2340 8010 2400 8090
rect 2200 7950 2400 8010
rect 2600 8090 2800 8150
rect 2600 8010 2660 8090
rect 2740 8010 2800 8090
rect 2600 7950 2800 8010
rect 3000 8090 3200 8150
rect 3000 8010 3060 8090
rect 3140 8010 3200 8090
rect 3000 7950 3200 8010
rect 3400 8090 3600 8150
rect 3400 8010 3460 8090
rect 3540 8010 3600 8090
rect 3400 7950 3600 8010
rect 3800 8090 4000 8150
rect 3800 8010 3860 8090
rect 3940 8010 4000 8090
rect 3800 7950 4000 8010
rect 4200 8090 4400 8150
rect 4200 8010 4260 8090
rect 4340 8010 4400 8090
rect 4200 7950 4400 8010
rect 4600 8090 4800 8150
rect 4600 8010 4660 8090
rect 4740 8010 4800 8090
rect 4600 7950 4800 8010
rect 5000 8090 5200 8150
rect 5000 8010 5060 8090
rect 5140 8010 5200 8090
rect 5000 7950 5200 8010
rect 5400 8090 5600 8150
rect 5400 8010 5460 8090
rect 5540 8010 5600 8090
rect 5400 7950 5600 8010
rect 5800 8090 6000 8150
rect 5800 8010 5860 8090
rect 5940 8010 6000 8090
rect 5800 7950 6000 8010
rect 6200 8090 6400 8150
rect 6200 8010 6260 8090
rect 6340 8010 6400 8090
rect 6200 7950 6400 8010
rect 6600 8090 6800 8150
rect 6600 8010 6660 8090
rect 6740 8010 6800 8090
rect 6600 7950 6800 8010
rect 7000 8090 7200 8150
rect 7000 8010 7060 8090
rect 7140 8010 7200 8090
rect 7000 7950 7200 8010
rect 7400 8090 7600 8150
rect 7400 8010 7460 8090
rect 7540 8010 7600 8090
rect 7400 7950 7600 8010
rect 7800 8090 8000 8150
rect 7800 8010 7860 8090
rect 7940 8010 8000 8090
rect 7800 7950 8000 8010
rect 8200 8090 8400 8150
rect 8200 8010 8260 8090
rect 8340 8010 8400 8090
rect 8200 7950 8400 8010
rect 8600 8090 8800 8150
rect 8600 8010 8660 8090
rect 8740 8010 8800 8090
rect 8600 7950 8800 8010
rect 9000 8090 9200 8150
rect 9000 8010 9060 8090
rect 9140 8010 9200 8090
rect 9000 7950 9200 8010
rect 9400 8090 9600 8150
rect 9400 8010 9460 8090
rect 9540 8010 9600 8090
rect 9400 7950 9600 8010
rect 9800 8090 10000 8150
rect 9800 8010 9860 8090
rect 9940 8010 10000 8090
rect 9800 7950 10000 8010
rect 2200 7690 2400 7750
rect 2200 7610 2260 7690
rect 2340 7610 2400 7690
rect 2200 7550 2400 7610
rect 2600 7690 2800 7750
rect 2600 7610 2660 7690
rect 2740 7610 2800 7690
rect 2600 7550 2800 7610
rect 3000 7690 3200 7750
rect 3000 7610 3060 7690
rect 3140 7610 3200 7690
rect 3000 7550 3200 7610
rect 3400 7690 3600 7750
rect 3400 7610 3460 7690
rect 3540 7610 3600 7690
rect 3400 7550 3600 7610
rect 3800 7690 4000 7750
rect 3800 7610 3860 7690
rect 3940 7610 4000 7690
rect 3800 7550 4000 7610
rect 4200 7690 4400 7750
rect 4200 7610 4260 7690
rect 4340 7610 4400 7690
rect 4200 7550 4400 7610
rect 4600 7690 4800 7750
rect 4600 7610 4660 7690
rect 4740 7610 4800 7690
rect 4600 7550 4800 7610
rect 5000 7690 5200 7750
rect 5000 7610 5060 7690
rect 5140 7610 5200 7690
rect 5000 7550 5200 7610
rect 5400 7690 5600 7750
rect 5400 7610 5460 7690
rect 5540 7610 5600 7690
rect 5400 7550 5600 7610
rect 5800 7690 6000 7750
rect 5800 7610 5860 7690
rect 5940 7610 6000 7690
rect 5800 7550 6000 7610
rect 6200 7690 6400 7750
rect 6200 7610 6260 7690
rect 6340 7610 6400 7690
rect 6200 7550 6400 7610
rect 6600 7690 6800 7750
rect 6600 7610 6660 7690
rect 6740 7610 6800 7690
rect 6600 7550 6800 7610
rect 7000 7690 7200 7750
rect 7000 7610 7060 7690
rect 7140 7610 7200 7690
rect 7000 7550 7200 7610
rect 7400 7690 7600 7750
rect 7400 7610 7460 7690
rect 7540 7610 7600 7690
rect 7400 7550 7600 7610
rect 7800 7690 8000 7750
rect 7800 7610 7860 7690
rect 7940 7610 8000 7690
rect 7800 7550 8000 7610
rect 8200 7690 8400 7750
rect 8200 7610 8260 7690
rect 8340 7610 8400 7690
rect 8200 7550 8400 7610
rect 8600 7690 8800 7750
rect 8600 7610 8660 7690
rect 8740 7610 8800 7690
rect 8600 7550 8800 7610
rect 9000 7690 9200 7750
rect 9000 7610 9060 7690
rect 9140 7610 9200 7690
rect 9000 7550 9200 7610
rect 9400 7690 9600 7750
rect 9400 7610 9460 7690
rect 9540 7610 9600 7690
rect 9400 7550 9600 7610
rect 9800 7690 10000 7750
rect 9800 7610 9860 7690
rect 9940 7610 10000 7690
rect 9800 7550 10000 7610
rect 2200 7290 2400 7350
rect 2200 7210 2260 7290
rect 2340 7210 2400 7290
rect 2200 7150 2400 7210
rect 2600 7290 2800 7350
rect 2600 7210 2660 7290
rect 2740 7210 2800 7290
rect 2600 7150 2800 7210
rect 3000 7290 3200 7350
rect 3000 7210 3060 7290
rect 3140 7210 3200 7290
rect 3000 7150 3200 7210
rect 3400 7290 3600 7350
rect 3400 7210 3460 7290
rect 3540 7210 3600 7290
rect 3400 7150 3600 7210
rect 3800 7290 4000 7350
rect 3800 7210 3860 7290
rect 3940 7210 4000 7290
rect 3800 7150 4000 7210
rect 4200 7290 4400 7350
rect 4200 7210 4260 7290
rect 4340 7210 4400 7290
rect 4200 7150 4400 7210
rect 4600 7290 4800 7350
rect 4600 7210 4660 7290
rect 4740 7210 4800 7290
rect 4600 7150 4800 7210
rect 5000 7290 5200 7350
rect 5000 7210 5060 7290
rect 5140 7210 5200 7290
rect 5000 7150 5200 7210
rect 5400 7290 5600 7350
rect 5400 7210 5460 7290
rect 5540 7210 5600 7290
rect 5400 7150 5600 7210
rect 5800 7290 6000 7350
rect 5800 7210 5860 7290
rect 5940 7210 6000 7290
rect 5800 7150 6000 7210
rect 6200 7290 6400 7350
rect 6200 7210 6260 7290
rect 6340 7210 6400 7290
rect 6200 7150 6400 7210
rect 6600 7290 6800 7350
rect 6600 7210 6660 7290
rect 6740 7210 6800 7290
rect 6600 7150 6800 7210
rect 7000 7290 7200 7350
rect 7000 7210 7060 7290
rect 7140 7210 7200 7290
rect 7000 7150 7200 7210
rect 7400 7290 7600 7350
rect 7400 7210 7460 7290
rect 7540 7210 7600 7290
rect 7400 7150 7600 7210
rect 7800 7290 8000 7350
rect 7800 7210 7860 7290
rect 7940 7210 8000 7290
rect 7800 7150 8000 7210
rect 8200 7290 8400 7350
rect 8200 7210 8260 7290
rect 8340 7210 8400 7290
rect 8200 7150 8400 7210
rect 8600 7290 8800 7350
rect 8600 7210 8660 7290
rect 8740 7210 8800 7290
rect 8600 7150 8800 7210
rect 9000 7290 9200 7350
rect 9000 7210 9060 7290
rect 9140 7210 9200 7290
rect 9000 7150 9200 7210
rect 9400 7290 9600 7350
rect 9400 7210 9460 7290
rect 9540 7210 9600 7290
rect 9400 7150 9600 7210
rect 9800 7290 10000 7350
rect 9800 7210 9860 7290
rect 9940 7210 10000 7290
rect 9800 7150 10000 7210
rect 2200 6890 2400 6950
rect 2200 6810 2260 6890
rect 2340 6810 2400 6890
rect 2200 6750 2400 6810
rect 2600 6890 2800 6950
rect 2600 6810 2660 6890
rect 2740 6810 2800 6890
rect 2600 6750 2800 6810
rect 3000 6890 3200 6950
rect 3000 6810 3060 6890
rect 3140 6810 3200 6890
rect 3000 6750 3200 6810
rect 3400 6890 3600 6950
rect 3400 6810 3460 6890
rect 3540 6810 3600 6890
rect 3400 6750 3600 6810
rect 3800 6890 4000 6950
rect 3800 6810 3860 6890
rect 3940 6810 4000 6890
rect 3800 6750 4000 6810
rect 4200 6890 4400 6950
rect 4200 6810 4260 6890
rect 4340 6810 4400 6890
rect 4200 6750 4400 6810
rect 4600 6890 4800 6950
rect 4600 6810 4660 6890
rect 4740 6810 4800 6890
rect 4600 6750 4800 6810
rect 5000 6890 5200 6950
rect 5000 6810 5060 6890
rect 5140 6810 5200 6890
rect 5000 6750 5200 6810
rect 5400 6890 5600 6950
rect 5400 6810 5460 6890
rect 5540 6810 5600 6890
rect 5400 6750 5600 6810
rect 5800 6890 6000 6950
rect 5800 6810 5860 6890
rect 5940 6810 6000 6890
rect 5800 6750 6000 6810
rect 6200 6890 6400 6950
rect 6200 6810 6260 6890
rect 6340 6810 6400 6890
rect 6200 6750 6400 6810
rect 6600 6890 6800 6950
rect 6600 6810 6660 6890
rect 6740 6810 6800 6890
rect 6600 6750 6800 6810
rect 7000 6890 7200 6950
rect 7000 6810 7060 6890
rect 7140 6810 7200 6890
rect 7000 6750 7200 6810
rect 7400 6890 7600 6950
rect 7400 6810 7460 6890
rect 7540 6810 7600 6890
rect 7400 6750 7600 6810
rect 7800 6890 8000 6950
rect 7800 6810 7860 6890
rect 7940 6810 8000 6890
rect 7800 6750 8000 6810
rect 8200 6890 8400 6950
rect 8200 6810 8260 6890
rect 8340 6810 8400 6890
rect 8200 6750 8400 6810
rect 8600 6890 8800 6950
rect 8600 6810 8660 6890
rect 8740 6810 8800 6890
rect 8600 6750 8800 6810
rect 9000 6890 9200 6950
rect 9000 6810 9060 6890
rect 9140 6810 9200 6890
rect 9000 6750 9200 6810
rect 9400 6890 9600 6950
rect 9400 6810 9460 6890
rect 9540 6810 9600 6890
rect 9400 6750 9600 6810
rect 9800 6890 10000 6950
rect 9800 6810 9860 6890
rect 9940 6810 10000 6890
rect 9800 6750 10000 6810
rect 2200 6490 2400 6550
rect 2200 6410 2260 6490
rect 2340 6410 2400 6490
rect 2200 6350 2400 6410
rect 2600 6490 2800 6550
rect 2600 6410 2660 6490
rect 2740 6410 2800 6490
rect 2600 6350 2800 6410
rect 3000 6490 3200 6550
rect 3000 6410 3060 6490
rect 3140 6410 3200 6490
rect 3000 6350 3200 6410
rect 3400 6490 3600 6550
rect 3400 6410 3460 6490
rect 3540 6410 3600 6490
rect 3400 6350 3600 6410
rect 3800 6490 4000 6550
rect 3800 6410 3860 6490
rect 3940 6410 4000 6490
rect 3800 6350 4000 6410
rect 4200 6490 4400 6550
rect 4200 6410 4260 6490
rect 4340 6410 4400 6490
rect 4200 6350 4400 6410
rect 4600 6490 4800 6550
rect 4600 6410 4660 6490
rect 4740 6410 4800 6490
rect 4600 6350 4800 6410
rect 5000 6490 5200 6550
rect 5000 6410 5060 6490
rect 5140 6410 5200 6490
rect 5000 6350 5200 6410
rect 5400 6490 5600 6550
rect 5400 6410 5460 6490
rect 5540 6410 5600 6490
rect 5400 6350 5600 6410
rect 5800 6490 6000 6550
rect 5800 6410 5860 6490
rect 5940 6410 6000 6490
rect 5800 6350 6000 6410
rect 6200 6490 6400 6550
rect 6200 6410 6260 6490
rect 6340 6410 6400 6490
rect 6200 6350 6400 6410
rect 6600 6490 6800 6550
rect 6600 6410 6660 6490
rect 6740 6410 6800 6490
rect 6600 6350 6800 6410
rect 7000 6490 7200 6550
rect 7000 6410 7060 6490
rect 7140 6410 7200 6490
rect 7000 6350 7200 6410
rect 7400 6490 7600 6550
rect 7400 6410 7460 6490
rect 7540 6410 7600 6490
rect 7400 6350 7600 6410
rect 7800 6490 8000 6550
rect 7800 6410 7860 6490
rect 7940 6410 8000 6490
rect 7800 6350 8000 6410
rect 8200 6490 8400 6550
rect 8200 6410 8260 6490
rect 8340 6410 8400 6490
rect 8200 6350 8400 6410
rect 8600 6490 8800 6550
rect 8600 6410 8660 6490
rect 8740 6410 8800 6490
rect 8600 6350 8800 6410
rect 9000 6490 9200 6550
rect 9000 6410 9060 6490
rect 9140 6410 9200 6490
rect 9000 6350 9200 6410
rect 9400 6490 9600 6550
rect 9400 6410 9460 6490
rect 9540 6410 9600 6490
rect 9400 6350 9600 6410
rect 9800 6490 10000 6550
rect 9800 6410 9860 6490
rect 9940 6410 10000 6490
rect 9800 6350 10000 6410
rect 2200 6090 2400 6150
rect 2200 6010 2260 6090
rect 2340 6010 2400 6090
rect 2200 5950 2400 6010
rect 2600 6090 2800 6150
rect 2600 6010 2660 6090
rect 2740 6010 2800 6090
rect 2600 5950 2800 6010
rect 3000 6090 3200 6150
rect 3000 6010 3060 6090
rect 3140 6010 3200 6090
rect 3000 5950 3200 6010
rect 3400 6090 3600 6150
rect 3400 6010 3460 6090
rect 3540 6010 3600 6090
rect 3400 5950 3600 6010
rect 3800 6090 4000 6150
rect 3800 6010 3860 6090
rect 3940 6010 4000 6090
rect 3800 5950 4000 6010
rect 4200 6090 4400 6150
rect 4200 6010 4260 6090
rect 4340 6010 4400 6090
rect 4200 5950 4400 6010
rect 4600 6090 4800 6150
rect 4600 6010 4660 6090
rect 4740 6010 4800 6090
rect 4600 5950 4800 6010
rect 5000 6090 5200 6150
rect 5000 6010 5060 6090
rect 5140 6010 5200 6090
rect 5000 5950 5200 6010
rect 5400 6090 5600 6150
rect 5400 6010 5460 6090
rect 5540 6010 5600 6090
rect 5400 5950 5600 6010
rect 5800 6090 6000 6150
rect 5800 6010 5860 6090
rect 5940 6010 6000 6090
rect 5800 5950 6000 6010
rect 6200 6090 6400 6150
rect 6200 6010 6260 6090
rect 6340 6010 6400 6090
rect 6200 5950 6400 6010
rect 6600 6090 6800 6150
rect 6600 6010 6660 6090
rect 6740 6010 6800 6090
rect 6600 5950 6800 6010
rect 7000 6090 7200 6150
rect 7000 6010 7060 6090
rect 7140 6010 7200 6090
rect 7000 5950 7200 6010
rect 7400 6090 7600 6150
rect 7400 6010 7460 6090
rect 7540 6010 7600 6090
rect 7400 5950 7600 6010
rect 7800 6090 8000 6150
rect 7800 6010 7860 6090
rect 7940 6010 8000 6090
rect 7800 5950 8000 6010
rect 8200 6090 8400 6150
rect 8200 6010 8260 6090
rect 8340 6010 8400 6090
rect 8200 5950 8400 6010
rect 8600 6090 8800 6150
rect 8600 6010 8660 6090
rect 8740 6010 8800 6090
rect 8600 5950 8800 6010
rect 9000 6090 9200 6150
rect 9000 6010 9060 6090
rect 9140 6010 9200 6090
rect 9000 5950 9200 6010
rect 9400 6090 9600 6150
rect 9400 6010 9460 6090
rect 9540 6010 9600 6090
rect 9400 5950 9600 6010
rect 9800 6090 10000 6150
rect 9800 6010 9860 6090
rect 9940 6010 10000 6090
rect 9800 5950 10000 6010
rect 2200 5690 2400 5750
rect 2200 5610 2260 5690
rect 2340 5610 2400 5690
rect 2200 5550 2400 5610
rect 2600 5690 2800 5750
rect 2600 5610 2660 5690
rect 2740 5610 2800 5690
rect 2600 5550 2800 5610
rect 3000 5690 3200 5750
rect 3000 5610 3060 5690
rect 3140 5610 3200 5690
rect 3000 5550 3200 5610
rect 3400 5690 3600 5750
rect 3400 5610 3460 5690
rect 3540 5610 3600 5690
rect 3400 5550 3600 5610
rect 3800 5690 4000 5750
rect 3800 5610 3860 5690
rect 3940 5610 4000 5690
rect 3800 5550 4000 5610
rect 4200 5690 4400 5750
rect 4200 5610 4260 5690
rect 4340 5610 4400 5690
rect 4200 5550 4400 5610
rect 4600 5690 4800 5750
rect 4600 5610 4660 5690
rect 4740 5610 4800 5690
rect 4600 5550 4800 5610
rect 5000 5690 5200 5750
rect 5000 5610 5060 5690
rect 5140 5610 5200 5690
rect 5000 5550 5200 5610
rect 5400 5690 5600 5750
rect 5400 5610 5460 5690
rect 5540 5610 5600 5690
rect 5400 5550 5600 5610
rect 5800 5690 6000 5750
rect 5800 5610 5860 5690
rect 5940 5610 6000 5690
rect 5800 5550 6000 5610
rect 6200 5690 6400 5750
rect 6200 5610 6260 5690
rect 6340 5610 6400 5690
rect 6200 5550 6400 5610
rect 6600 5690 6800 5750
rect 6600 5610 6660 5690
rect 6740 5610 6800 5690
rect 6600 5550 6800 5610
rect 7000 5690 7200 5750
rect 7000 5610 7060 5690
rect 7140 5610 7200 5690
rect 7000 5550 7200 5610
rect 7400 5690 7600 5750
rect 7400 5610 7460 5690
rect 7540 5610 7600 5690
rect 7400 5550 7600 5610
rect 7800 5690 8000 5750
rect 7800 5610 7860 5690
rect 7940 5610 8000 5690
rect 7800 5550 8000 5610
rect 8200 5690 8400 5750
rect 8200 5610 8260 5690
rect 8340 5610 8400 5690
rect 8200 5550 8400 5610
rect 8600 5690 8800 5750
rect 8600 5610 8660 5690
rect 8740 5610 8800 5690
rect 8600 5550 8800 5610
rect 9000 5690 9200 5750
rect 9000 5610 9060 5690
rect 9140 5610 9200 5690
rect 9000 5550 9200 5610
rect 9400 5690 9600 5750
rect 9400 5610 9460 5690
rect 9540 5610 9600 5690
rect 9400 5550 9600 5610
rect 9800 5690 10000 5750
rect 9800 5610 9860 5690
rect 9940 5610 10000 5690
rect 9800 5550 10000 5610
rect 2200 5290 2400 5350
rect 2200 5210 2260 5290
rect 2340 5210 2400 5290
rect 2200 5150 2400 5210
rect 2600 5290 2800 5350
rect 2600 5210 2660 5290
rect 2740 5210 2800 5290
rect 2600 5150 2800 5210
rect 3000 5290 3200 5350
rect 3000 5210 3060 5290
rect 3140 5210 3200 5290
rect 3000 5150 3200 5210
rect 3400 5290 3600 5350
rect 3400 5210 3460 5290
rect 3540 5210 3600 5290
rect 3400 5150 3600 5210
rect 3800 5290 4000 5350
rect 3800 5210 3860 5290
rect 3940 5210 4000 5290
rect 3800 5150 4000 5210
rect 4200 5290 4400 5350
rect 4200 5210 4260 5290
rect 4340 5210 4400 5290
rect 4200 5150 4400 5210
rect 4600 5290 4800 5350
rect 4600 5210 4660 5290
rect 4740 5210 4800 5290
rect 4600 5150 4800 5210
rect 5000 5290 5200 5350
rect 5000 5210 5060 5290
rect 5140 5210 5200 5290
rect 5000 5150 5200 5210
rect 5400 5290 5600 5350
rect 5400 5210 5460 5290
rect 5540 5210 5600 5290
rect 5400 5150 5600 5210
rect 5800 5290 6000 5350
rect 5800 5210 5860 5290
rect 5940 5210 6000 5290
rect 5800 5150 6000 5210
rect 6200 5290 6400 5350
rect 6200 5210 6260 5290
rect 6340 5210 6400 5290
rect 6200 5150 6400 5210
rect 6600 5290 6800 5350
rect 6600 5210 6660 5290
rect 6740 5210 6800 5290
rect 6600 5150 6800 5210
rect 7000 5290 7200 5350
rect 7000 5210 7060 5290
rect 7140 5210 7200 5290
rect 7000 5150 7200 5210
rect 7400 5290 7600 5350
rect 7400 5210 7460 5290
rect 7540 5210 7600 5290
rect 7400 5150 7600 5210
rect 7800 5290 8000 5350
rect 7800 5210 7860 5290
rect 7940 5210 8000 5290
rect 7800 5150 8000 5210
rect 8200 5290 8400 5350
rect 8200 5210 8260 5290
rect 8340 5210 8400 5290
rect 8200 5150 8400 5210
rect 8600 5290 8800 5350
rect 8600 5210 8660 5290
rect 8740 5210 8800 5290
rect 8600 5150 8800 5210
rect 9000 5290 9200 5350
rect 9000 5210 9060 5290
rect 9140 5210 9200 5290
rect 9000 5150 9200 5210
rect 9400 5290 9600 5350
rect 9400 5210 9460 5290
rect 9540 5210 9600 5290
rect 9400 5150 9600 5210
rect 9800 5290 10000 5350
rect 9800 5210 9860 5290
rect 9940 5210 10000 5290
rect 9800 5150 10000 5210
rect 2200 4890 2400 4950
rect 2200 4810 2260 4890
rect 2340 4810 2400 4890
rect 2200 4750 2400 4810
rect 2600 4890 2800 4950
rect 2600 4810 2660 4890
rect 2740 4810 2800 4890
rect 2600 4750 2800 4810
rect 3000 4890 3200 4950
rect 3000 4810 3060 4890
rect 3140 4810 3200 4890
rect 3000 4750 3200 4810
rect 3400 4890 3600 4950
rect 3400 4810 3460 4890
rect 3540 4810 3600 4890
rect 3400 4750 3600 4810
rect 3800 4890 4000 4950
rect 3800 4810 3860 4890
rect 3940 4810 4000 4890
rect 3800 4750 4000 4810
rect 4200 4890 4400 4950
rect 4200 4810 4260 4890
rect 4340 4810 4400 4890
rect 4200 4750 4400 4810
rect 4600 4890 4800 4950
rect 4600 4810 4660 4890
rect 4740 4810 4800 4890
rect 4600 4750 4800 4810
rect 5000 4890 5200 4950
rect 5000 4810 5060 4890
rect 5140 4810 5200 4890
rect 5000 4750 5200 4810
rect 5400 4890 5600 4950
rect 5400 4810 5460 4890
rect 5540 4810 5600 4890
rect 5400 4750 5600 4810
rect 5800 4890 6000 4950
rect 5800 4810 5860 4890
rect 5940 4810 6000 4890
rect 5800 4750 6000 4810
rect 6200 4890 6400 4950
rect 6200 4810 6260 4890
rect 6340 4810 6400 4890
rect 6200 4750 6400 4810
rect 6600 4890 6800 4950
rect 6600 4810 6660 4890
rect 6740 4810 6800 4890
rect 6600 4750 6800 4810
rect 7000 4890 7200 4950
rect 7000 4810 7060 4890
rect 7140 4810 7200 4890
rect 7000 4750 7200 4810
rect 7400 4890 7600 4950
rect 7400 4810 7460 4890
rect 7540 4810 7600 4890
rect 7400 4750 7600 4810
rect 7800 4890 8000 4950
rect 7800 4810 7860 4890
rect 7940 4810 8000 4890
rect 7800 4750 8000 4810
rect 8200 4890 8400 4950
rect 8200 4810 8260 4890
rect 8340 4810 8400 4890
rect 8200 4750 8400 4810
rect 8600 4890 8800 4950
rect 8600 4810 8660 4890
rect 8740 4810 8800 4890
rect 8600 4750 8800 4810
rect 9000 4890 9200 4950
rect 9000 4810 9060 4890
rect 9140 4810 9200 4890
rect 9000 4750 9200 4810
rect 9400 4890 9600 4950
rect 9400 4810 9460 4890
rect 9540 4810 9600 4890
rect 9400 4750 9600 4810
rect 9800 4890 10000 4950
rect 9800 4810 9860 4890
rect 9940 4810 10000 4890
rect 9800 4750 10000 4810
rect 2200 4490 2400 4550
rect 2200 4410 2260 4490
rect 2340 4410 2400 4490
rect 2200 4350 2400 4410
rect 2600 4490 2800 4550
rect 2600 4410 2660 4490
rect 2740 4410 2800 4490
rect 2600 4350 2800 4410
rect 3000 4490 3200 4550
rect 3000 4410 3060 4490
rect 3140 4410 3200 4490
rect 3000 4350 3200 4410
rect 3400 4490 3600 4550
rect 3400 4410 3460 4490
rect 3540 4410 3600 4490
rect 3400 4350 3600 4410
rect 3800 4490 4000 4550
rect 3800 4410 3860 4490
rect 3940 4410 4000 4490
rect 3800 4350 4000 4410
rect 4200 4490 4400 4550
rect 4200 4410 4260 4490
rect 4340 4410 4400 4490
rect 4200 4350 4400 4410
rect 4600 4490 4800 4550
rect 4600 4410 4660 4490
rect 4740 4410 4800 4490
rect 4600 4350 4800 4410
rect 5000 4490 5200 4550
rect 5000 4410 5060 4490
rect 5140 4410 5200 4490
rect 5000 4350 5200 4410
rect 5400 4490 5600 4550
rect 5400 4410 5460 4490
rect 5540 4410 5600 4490
rect 5400 4350 5600 4410
rect 5800 4490 6000 4550
rect 5800 4410 5860 4490
rect 5940 4410 6000 4490
rect 5800 4350 6000 4410
rect 6200 4490 6400 4550
rect 6200 4410 6260 4490
rect 6340 4410 6400 4490
rect 6200 4350 6400 4410
rect 6600 4490 6800 4550
rect 6600 4410 6660 4490
rect 6740 4410 6800 4490
rect 6600 4350 6800 4410
rect 7000 4490 7200 4550
rect 7000 4410 7060 4490
rect 7140 4410 7200 4490
rect 7000 4350 7200 4410
rect 7400 4490 7600 4550
rect 7400 4410 7460 4490
rect 7540 4410 7600 4490
rect 7400 4350 7600 4410
rect 7800 4490 8000 4550
rect 7800 4410 7860 4490
rect 7940 4410 8000 4490
rect 7800 4350 8000 4410
rect 8200 4490 8400 4550
rect 8200 4410 8260 4490
rect 8340 4410 8400 4490
rect 8200 4350 8400 4410
rect 8600 4490 8800 4550
rect 8600 4410 8660 4490
rect 8740 4410 8800 4490
rect 8600 4350 8800 4410
rect 9000 4490 9200 4550
rect 9000 4410 9060 4490
rect 9140 4410 9200 4490
rect 9000 4350 9200 4410
rect 9400 4490 9600 4550
rect 9400 4410 9460 4490
rect 9540 4410 9600 4490
rect 9400 4350 9600 4410
rect 9800 4490 10000 4550
rect 9800 4410 9860 4490
rect 9940 4410 10000 4490
rect 9800 4350 10000 4410
rect 2200 4090 2400 4150
rect 2200 4010 2260 4090
rect 2340 4010 2400 4090
rect 2200 3950 2400 4010
rect 2600 4090 2800 4150
rect 2600 4010 2660 4090
rect 2740 4010 2800 4090
rect 2600 3950 2800 4010
rect 3000 4090 3200 4150
rect 3000 4010 3060 4090
rect 3140 4010 3200 4090
rect 3000 3950 3200 4010
rect 3400 4090 3600 4150
rect 3400 4010 3460 4090
rect 3540 4010 3600 4090
rect 3400 3950 3600 4010
rect 3800 4090 4000 4150
rect 3800 4010 3860 4090
rect 3940 4010 4000 4090
rect 3800 3950 4000 4010
rect 4200 4090 4400 4150
rect 4200 4010 4260 4090
rect 4340 4010 4400 4090
rect 4200 3950 4400 4010
rect 4600 4090 4800 4150
rect 4600 4010 4660 4090
rect 4740 4010 4800 4090
rect 4600 3950 4800 4010
rect 5000 4090 5200 4150
rect 5000 4010 5060 4090
rect 5140 4010 5200 4090
rect 5000 3950 5200 4010
rect 5400 4090 5600 4150
rect 5400 4010 5460 4090
rect 5540 4010 5600 4090
rect 5400 3950 5600 4010
rect 5800 4090 6000 4150
rect 5800 4010 5860 4090
rect 5940 4010 6000 4090
rect 5800 3950 6000 4010
rect 6200 4090 6400 4150
rect 6200 4010 6260 4090
rect 6340 4010 6400 4090
rect 6200 3950 6400 4010
rect 6600 4090 6800 4150
rect 6600 4010 6660 4090
rect 6740 4010 6800 4090
rect 6600 3950 6800 4010
rect 7000 4090 7200 4150
rect 7000 4010 7060 4090
rect 7140 4010 7200 4090
rect 7000 3950 7200 4010
rect 7400 4090 7600 4150
rect 7400 4010 7460 4090
rect 7540 4010 7600 4090
rect 7400 3950 7600 4010
rect 7800 4090 8000 4150
rect 7800 4010 7860 4090
rect 7940 4010 8000 4090
rect 7800 3950 8000 4010
rect 8200 4090 8400 4150
rect 8200 4010 8260 4090
rect 8340 4010 8400 4090
rect 8200 3950 8400 4010
rect 8600 4090 8800 4150
rect 8600 4010 8660 4090
rect 8740 4010 8800 4090
rect 8600 3950 8800 4010
rect 9000 4090 9200 4150
rect 9000 4010 9060 4090
rect 9140 4010 9200 4090
rect 9000 3950 9200 4010
rect 9400 4090 9600 4150
rect 9400 4010 9460 4090
rect 9540 4010 9600 4090
rect 9400 3950 9600 4010
rect 9800 4090 10000 4150
rect 9800 4010 9860 4090
rect 9940 4010 10000 4090
rect 9800 3950 10000 4010
rect 2200 3690 2400 3750
rect 2200 3610 2260 3690
rect 2340 3610 2400 3690
rect 2200 3550 2400 3610
rect 2600 3690 2800 3750
rect 2600 3610 2660 3690
rect 2740 3610 2800 3690
rect 2600 3550 2800 3610
rect 3000 3690 3200 3750
rect 3000 3610 3060 3690
rect 3140 3610 3200 3690
rect 3000 3550 3200 3610
rect 3400 3690 3600 3750
rect 3400 3610 3460 3690
rect 3540 3610 3600 3690
rect 3400 3550 3600 3610
rect 3800 3690 4000 3750
rect 3800 3610 3860 3690
rect 3940 3610 4000 3690
rect 3800 3550 4000 3610
rect 4200 3690 4400 3750
rect 4200 3610 4260 3690
rect 4340 3610 4400 3690
rect 4200 3550 4400 3610
rect 4600 3690 4800 3750
rect 4600 3610 4660 3690
rect 4740 3610 4800 3690
rect 4600 3550 4800 3610
rect 5000 3690 5200 3750
rect 5000 3610 5060 3690
rect 5140 3610 5200 3690
rect 5000 3550 5200 3610
rect 5400 3690 5600 3750
rect 5400 3610 5460 3690
rect 5540 3610 5600 3690
rect 5400 3550 5600 3610
rect 5800 3690 6000 3750
rect 5800 3610 5860 3690
rect 5940 3610 6000 3690
rect 5800 3550 6000 3610
rect 6200 3690 6400 3750
rect 6200 3610 6260 3690
rect 6340 3610 6400 3690
rect 6200 3550 6400 3610
rect 6600 3690 6800 3750
rect 6600 3610 6660 3690
rect 6740 3610 6800 3690
rect 6600 3550 6800 3610
rect 7000 3690 7200 3750
rect 7000 3610 7060 3690
rect 7140 3610 7200 3690
rect 7000 3550 7200 3610
rect 7400 3690 7600 3750
rect 7400 3610 7460 3690
rect 7540 3610 7600 3690
rect 7400 3550 7600 3610
rect 7800 3690 8000 3750
rect 7800 3610 7860 3690
rect 7940 3610 8000 3690
rect 7800 3550 8000 3610
rect 8200 3690 8400 3750
rect 8200 3610 8260 3690
rect 8340 3610 8400 3690
rect 8200 3550 8400 3610
rect 8600 3690 8800 3750
rect 8600 3610 8660 3690
rect 8740 3610 8800 3690
rect 8600 3550 8800 3610
rect 9000 3690 9200 3750
rect 9000 3610 9060 3690
rect 9140 3610 9200 3690
rect 9000 3550 9200 3610
rect 9400 3690 9600 3750
rect 9400 3610 9460 3690
rect 9540 3610 9600 3690
rect 9400 3550 9600 3610
rect 9800 3690 10000 3750
rect 9800 3610 9860 3690
rect 9940 3610 10000 3690
rect 9800 3550 10000 3610
rect 2200 3290 2400 3350
rect 2200 3210 2260 3290
rect 2340 3210 2400 3290
rect 2200 3150 2400 3210
rect 2600 3290 2800 3350
rect 2600 3210 2660 3290
rect 2740 3210 2800 3290
rect 2600 3150 2800 3210
rect 3000 3290 3200 3350
rect 3000 3210 3060 3290
rect 3140 3210 3200 3290
rect 3000 3150 3200 3210
rect 3400 3290 3600 3350
rect 3400 3210 3460 3290
rect 3540 3210 3600 3290
rect 3400 3150 3600 3210
rect 3800 3290 4000 3350
rect 3800 3210 3860 3290
rect 3940 3210 4000 3290
rect 3800 3150 4000 3210
rect 4200 3290 4400 3350
rect 4200 3210 4260 3290
rect 4340 3210 4400 3290
rect 4200 3150 4400 3210
rect 4600 3290 4800 3350
rect 4600 3210 4660 3290
rect 4740 3210 4800 3290
rect 4600 3150 4800 3210
rect 5000 3290 5200 3350
rect 5000 3210 5060 3290
rect 5140 3210 5200 3290
rect 5000 3150 5200 3210
rect 5400 3290 5600 3350
rect 5400 3210 5460 3290
rect 5540 3210 5600 3290
rect 5400 3150 5600 3210
rect 5800 3290 6000 3350
rect 5800 3210 5860 3290
rect 5940 3210 6000 3290
rect 5800 3150 6000 3210
rect 6200 3290 6400 3350
rect 6200 3210 6260 3290
rect 6340 3210 6400 3290
rect 6200 3150 6400 3210
rect 6600 3290 6800 3350
rect 6600 3210 6660 3290
rect 6740 3210 6800 3290
rect 6600 3150 6800 3210
rect 7000 3290 7200 3350
rect 7000 3210 7060 3290
rect 7140 3210 7200 3290
rect 7000 3150 7200 3210
rect 7400 3290 7600 3350
rect 7400 3210 7460 3290
rect 7540 3210 7600 3290
rect 7400 3150 7600 3210
rect 7800 3290 8000 3350
rect 7800 3210 7860 3290
rect 7940 3210 8000 3290
rect 7800 3150 8000 3210
rect 8200 3290 8400 3350
rect 8200 3210 8260 3290
rect 8340 3210 8400 3290
rect 8200 3150 8400 3210
rect 8600 3290 8800 3350
rect 8600 3210 8660 3290
rect 8740 3210 8800 3290
rect 8600 3150 8800 3210
rect 9000 3290 9200 3350
rect 9000 3210 9060 3290
rect 9140 3210 9200 3290
rect 9000 3150 9200 3210
rect 9400 3290 9600 3350
rect 9400 3210 9460 3290
rect 9540 3210 9600 3290
rect 9400 3150 9600 3210
rect 9800 3290 10000 3350
rect 9800 3210 9860 3290
rect 9940 3210 10000 3290
rect 9800 3150 10000 3210
rect 2200 2890 2400 2950
rect 2200 2810 2260 2890
rect 2340 2810 2400 2890
rect 2200 2750 2400 2810
rect 2600 2890 2800 2950
rect 2600 2810 2660 2890
rect 2740 2810 2800 2890
rect 2600 2750 2800 2810
rect 3000 2890 3200 2950
rect 3000 2810 3060 2890
rect 3140 2810 3200 2890
rect 3000 2750 3200 2810
rect 3400 2890 3600 2950
rect 3400 2810 3460 2890
rect 3540 2810 3600 2890
rect 3400 2750 3600 2810
rect 3800 2890 4000 2950
rect 3800 2810 3860 2890
rect 3940 2810 4000 2890
rect 3800 2750 4000 2810
rect 4200 2890 4400 2950
rect 4200 2810 4260 2890
rect 4340 2810 4400 2890
rect 4200 2750 4400 2810
rect 4600 2890 4800 2950
rect 4600 2810 4660 2890
rect 4740 2810 4800 2890
rect 4600 2750 4800 2810
rect 5000 2890 5200 2950
rect 5000 2810 5060 2890
rect 5140 2810 5200 2890
rect 5000 2750 5200 2810
rect 5400 2890 5600 2950
rect 5400 2810 5460 2890
rect 5540 2810 5600 2890
rect 5400 2750 5600 2810
rect 5800 2890 6000 2950
rect 5800 2810 5860 2890
rect 5940 2810 6000 2890
rect 5800 2750 6000 2810
rect 6200 2890 6400 2950
rect 6200 2810 6260 2890
rect 6340 2810 6400 2890
rect 6200 2750 6400 2810
rect 6600 2890 6800 2950
rect 6600 2810 6660 2890
rect 6740 2810 6800 2890
rect 6600 2750 6800 2810
rect 7000 2890 7200 2950
rect 7000 2810 7060 2890
rect 7140 2810 7200 2890
rect 7000 2750 7200 2810
rect 7400 2890 7600 2950
rect 7400 2810 7460 2890
rect 7540 2810 7600 2890
rect 7400 2750 7600 2810
rect 7800 2890 8000 2950
rect 7800 2810 7860 2890
rect 7940 2810 8000 2890
rect 7800 2750 8000 2810
rect 8200 2890 8400 2950
rect 8200 2810 8260 2890
rect 8340 2810 8400 2890
rect 8200 2750 8400 2810
rect 8600 2890 8800 2950
rect 8600 2810 8660 2890
rect 8740 2810 8800 2890
rect 8600 2750 8800 2810
rect 9000 2890 9200 2950
rect 9000 2810 9060 2890
rect 9140 2810 9200 2890
rect 9000 2750 9200 2810
rect 9400 2890 9600 2950
rect 9400 2810 9460 2890
rect 9540 2810 9600 2890
rect 9400 2750 9600 2810
rect 9800 2890 10000 2950
rect 9800 2810 9860 2890
rect 9940 2810 10000 2890
rect 9800 2750 10000 2810
rect 2200 2490 2400 2550
rect 2200 2410 2260 2490
rect 2340 2410 2400 2490
rect 2200 2350 2400 2410
rect 2600 2490 2800 2550
rect 2600 2410 2660 2490
rect 2740 2410 2800 2490
rect 2600 2350 2800 2410
rect 3000 2490 3200 2550
rect 3000 2410 3060 2490
rect 3140 2410 3200 2490
rect 3000 2350 3200 2410
rect 3400 2490 3600 2550
rect 3400 2410 3460 2490
rect 3540 2410 3600 2490
rect 3400 2350 3600 2410
rect 3800 2490 4000 2550
rect 3800 2410 3860 2490
rect 3940 2410 4000 2490
rect 3800 2350 4000 2410
rect 4200 2490 4400 2550
rect 4200 2410 4260 2490
rect 4340 2410 4400 2490
rect 4200 2350 4400 2410
rect 4600 2490 4800 2550
rect 4600 2410 4660 2490
rect 4740 2410 4800 2490
rect 4600 2350 4800 2410
rect 5000 2490 5200 2550
rect 5000 2410 5060 2490
rect 5140 2410 5200 2490
rect 5000 2350 5200 2410
rect 5400 2490 5600 2550
rect 5400 2410 5460 2490
rect 5540 2410 5600 2490
rect 5400 2350 5600 2410
rect 5800 2490 6000 2550
rect 5800 2410 5860 2490
rect 5940 2410 6000 2490
rect 5800 2350 6000 2410
rect 6200 2490 6400 2550
rect 6200 2410 6260 2490
rect 6340 2410 6400 2490
rect 6200 2350 6400 2410
rect 6600 2490 6800 2550
rect 6600 2410 6660 2490
rect 6740 2410 6800 2490
rect 6600 2350 6800 2410
rect 7000 2490 7200 2550
rect 7000 2410 7060 2490
rect 7140 2410 7200 2490
rect 7000 2350 7200 2410
rect 7400 2490 7600 2550
rect 7400 2410 7460 2490
rect 7540 2410 7600 2490
rect 7400 2350 7600 2410
rect 7800 2490 8000 2550
rect 7800 2410 7860 2490
rect 7940 2410 8000 2490
rect 7800 2350 8000 2410
rect 8200 2490 8400 2550
rect 8200 2410 8260 2490
rect 8340 2410 8400 2490
rect 8200 2350 8400 2410
rect 8600 2490 8800 2550
rect 8600 2410 8660 2490
rect 8740 2410 8800 2490
rect 8600 2350 8800 2410
rect 9000 2490 9200 2550
rect 9000 2410 9060 2490
rect 9140 2410 9200 2490
rect 9000 2350 9200 2410
rect 9400 2490 9600 2550
rect 9400 2410 9460 2490
rect 9540 2410 9600 2490
rect 9400 2350 9600 2410
rect 9800 2490 10000 2550
rect 9800 2410 9860 2490
rect 9940 2410 10000 2490
rect 9800 2350 10000 2410
rect 2200 2090 2400 2150
rect 2200 2010 2260 2090
rect 2340 2010 2400 2090
rect 2200 1950 2400 2010
rect 2600 2090 2800 2150
rect 2600 2010 2660 2090
rect 2740 2010 2800 2090
rect 2600 1950 2800 2010
rect 3000 2090 3200 2150
rect 3000 2010 3060 2090
rect 3140 2010 3200 2090
rect 3000 1950 3200 2010
rect 3400 2090 3600 2150
rect 3400 2010 3460 2090
rect 3540 2010 3600 2090
rect 3400 1950 3600 2010
rect 3800 2090 4000 2150
rect 3800 2010 3860 2090
rect 3940 2010 4000 2090
rect 3800 1950 4000 2010
rect 4200 2090 4400 2150
rect 4200 2010 4260 2090
rect 4340 2010 4400 2090
rect 4200 1950 4400 2010
rect 4600 2090 4800 2150
rect 4600 2010 4660 2090
rect 4740 2010 4800 2090
rect 4600 1950 4800 2010
rect 5000 2090 5200 2150
rect 5000 2010 5060 2090
rect 5140 2010 5200 2090
rect 5000 1950 5200 2010
rect 5400 2090 5600 2150
rect 5400 2010 5460 2090
rect 5540 2010 5600 2090
rect 5400 1950 5600 2010
rect 5800 2090 6000 2150
rect 5800 2010 5860 2090
rect 5940 2010 6000 2090
rect 5800 1950 6000 2010
rect 6200 2090 6400 2150
rect 6200 2010 6260 2090
rect 6340 2010 6400 2090
rect 6200 1950 6400 2010
rect 6600 2090 6800 2150
rect 6600 2010 6660 2090
rect 6740 2010 6800 2090
rect 6600 1950 6800 2010
rect 7000 2090 7200 2150
rect 7000 2010 7060 2090
rect 7140 2010 7200 2090
rect 7000 1950 7200 2010
rect 7400 2090 7600 2150
rect 7400 2010 7460 2090
rect 7540 2010 7600 2090
rect 7400 1950 7600 2010
rect 7800 2090 8000 2150
rect 7800 2010 7860 2090
rect 7940 2010 8000 2090
rect 7800 1950 8000 2010
rect 8200 2090 8400 2150
rect 8200 2010 8260 2090
rect 8340 2010 8400 2090
rect 8200 1950 8400 2010
rect 8600 2090 8800 2150
rect 8600 2010 8660 2090
rect 8740 2010 8800 2090
rect 8600 1950 8800 2010
rect 9000 2090 9200 2150
rect 9000 2010 9060 2090
rect 9140 2010 9200 2090
rect 9000 1950 9200 2010
rect 9400 2090 9600 2150
rect 9400 2010 9460 2090
rect 9540 2010 9600 2090
rect 9400 1950 9600 2010
rect 9800 2090 10000 2150
rect 9800 2010 9860 2090
rect 9940 2010 10000 2090
rect 9800 1950 10000 2010
rect 2200 1690 2400 1750
rect 2200 1610 2260 1690
rect 2340 1610 2400 1690
rect 2200 1550 2400 1610
rect 2600 1690 2800 1750
rect 2600 1610 2660 1690
rect 2740 1610 2800 1690
rect 2600 1550 2800 1610
rect 3000 1690 3200 1750
rect 3000 1610 3060 1690
rect 3140 1610 3200 1690
rect 3000 1550 3200 1610
rect 3400 1690 3600 1750
rect 3400 1610 3460 1690
rect 3540 1610 3600 1690
rect 3400 1550 3600 1610
rect 3800 1690 4000 1750
rect 3800 1610 3860 1690
rect 3940 1610 4000 1690
rect 3800 1550 4000 1610
rect 4200 1690 4400 1750
rect 4200 1610 4260 1690
rect 4340 1610 4400 1690
rect 4200 1550 4400 1610
rect 4600 1690 4800 1750
rect 4600 1610 4660 1690
rect 4740 1610 4800 1690
rect 4600 1550 4800 1610
rect 5000 1690 5200 1750
rect 5000 1610 5060 1690
rect 5140 1610 5200 1690
rect 5000 1550 5200 1610
rect 5400 1690 5600 1750
rect 5400 1610 5460 1690
rect 5540 1610 5600 1690
rect 5400 1550 5600 1610
rect 5800 1690 6000 1750
rect 5800 1610 5860 1690
rect 5940 1610 6000 1690
rect 5800 1550 6000 1610
rect 6200 1690 6400 1750
rect 6200 1610 6260 1690
rect 6340 1610 6400 1690
rect 6200 1550 6400 1610
rect 6600 1690 6800 1750
rect 6600 1610 6660 1690
rect 6740 1610 6800 1690
rect 6600 1550 6800 1610
rect 7000 1690 7200 1750
rect 7000 1610 7060 1690
rect 7140 1610 7200 1690
rect 7000 1550 7200 1610
rect 7400 1690 7600 1750
rect 7400 1610 7460 1690
rect 7540 1610 7600 1690
rect 7400 1550 7600 1610
rect 7800 1690 8000 1750
rect 7800 1610 7860 1690
rect 7940 1610 8000 1690
rect 7800 1550 8000 1610
rect 8200 1690 8400 1750
rect 8200 1610 8260 1690
rect 8340 1610 8400 1690
rect 8200 1550 8400 1610
rect 8600 1690 8800 1750
rect 8600 1610 8660 1690
rect 8740 1610 8800 1690
rect 8600 1550 8800 1610
rect 9000 1690 9200 1750
rect 9000 1610 9060 1690
rect 9140 1610 9200 1690
rect 9000 1550 9200 1610
rect 9400 1690 9600 1750
rect 9400 1610 9460 1690
rect 9540 1610 9600 1690
rect 9400 1550 9600 1610
rect 9800 1690 10000 1750
rect 9800 1610 9860 1690
rect 9940 1610 10000 1690
rect 9800 1550 10000 1610
rect 2200 1290 2400 1350
rect 2200 1210 2260 1290
rect 2340 1210 2400 1290
rect 2200 1150 2400 1210
rect 2600 1290 2800 1350
rect 2600 1210 2660 1290
rect 2740 1210 2800 1290
rect 2600 1150 2800 1210
rect 3000 1290 3200 1350
rect 3000 1210 3060 1290
rect 3140 1210 3200 1290
rect 3000 1150 3200 1210
rect 3400 1290 3600 1350
rect 3400 1210 3460 1290
rect 3540 1210 3600 1290
rect 3400 1150 3600 1210
rect 3800 1290 4000 1350
rect 3800 1210 3860 1290
rect 3940 1210 4000 1290
rect 3800 1150 4000 1210
rect 4200 1290 4400 1350
rect 4200 1210 4260 1290
rect 4340 1210 4400 1290
rect 4200 1150 4400 1210
rect 4600 1290 4800 1350
rect 4600 1210 4660 1290
rect 4740 1210 4800 1290
rect 4600 1150 4800 1210
rect 5000 1290 5200 1350
rect 5000 1210 5060 1290
rect 5140 1210 5200 1290
rect 5000 1150 5200 1210
rect 5400 1290 5600 1350
rect 5400 1210 5460 1290
rect 5540 1210 5600 1290
rect 5400 1150 5600 1210
rect 5800 1290 6000 1350
rect 5800 1210 5860 1290
rect 5940 1210 6000 1290
rect 5800 1150 6000 1210
rect 6200 1290 6400 1350
rect 6200 1210 6260 1290
rect 6340 1210 6400 1290
rect 6200 1150 6400 1210
rect 6600 1290 6800 1350
rect 6600 1210 6660 1290
rect 6740 1210 6800 1290
rect 6600 1150 6800 1210
rect 7000 1290 7200 1350
rect 7000 1210 7060 1290
rect 7140 1210 7200 1290
rect 7000 1150 7200 1210
rect 7400 1290 7600 1350
rect 7400 1210 7460 1290
rect 7540 1210 7600 1290
rect 7400 1150 7600 1210
rect 7800 1290 8000 1350
rect 7800 1210 7860 1290
rect 7940 1210 8000 1290
rect 7800 1150 8000 1210
rect 8200 1290 8400 1350
rect 8200 1210 8260 1290
rect 8340 1210 8400 1290
rect 8200 1150 8400 1210
rect 8600 1290 8800 1350
rect 8600 1210 8660 1290
rect 8740 1210 8800 1290
rect 8600 1150 8800 1210
rect 9000 1290 9200 1350
rect 9000 1210 9060 1290
rect 9140 1210 9200 1290
rect 9000 1150 9200 1210
rect 9400 1290 9600 1350
rect 9400 1210 9460 1290
rect 9540 1210 9600 1290
rect 9400 1150 9600 1210
rect 9800 1290 10000 1350
rect 9800 1210 9860 1290
rect 9940 1210 10000 1290
rect 9800 1150 10000 1210
rect 2200 890 2400 950
rect 2200 810 2260 890
rect 2340 810 2400 890
rect 2200 750 2400 810
rect 2600 890 2800 950
rect 2600 810 2660 890
rect 2740 810 2800 890
rect 2600 750 2800 810
rect 3000 890 3200 950
rect 3000 810 3060 890
rect 3140 810 3200 890
rect 3000 750 3200 810
rect 3400 890 3600 950
rect 3400 810 3460 890
rect 3540 810 3600 890
rect 3400 750 3600 810
rect 3800 890 4000 950
rect 3800 810 3860 890
rect 3940 810 4000 890
rect 3800 750 4000 810
rect 4200 890 4400 950
rect 4200 810 4260 890
rect 4340 810 4400 890
rect 4200 750 4400 810
rect 4600 890 4800 950
rect 4600 810 4660 890
rect 4740 810 4800 890
rect 4600 750 4800 810
rect 5000 890 5200 950
rect 5000 810 5060 890
rect 5140 810 5200 890
rect 5000 750 5200 810
rect 5400 890 5600 950
rect 5400 810 5460 890
rect 5540 810 5600 890
rect 5400 750 5600 810
rect 5800 890 6000 950
rect 5800 810 5860 890
rect 5940 810 6000 890
rect 5800 750 6000 810
rect 6200 890 6400 950
rect 6200 810 6260 890
rect 6340 810 6400 890
rect 6200 750 6400 810
rect 6600 890 6800 950
rect 6600 810 6660 890
rect 6740 810 6800 890
rect 6600 750 6800 810
rect 7000 890 7200 950
rect 7000 810 7060 890
rect 7140 810 7200 890
rect 7000 750 7200 810
rect 7400 890 7600 950
rect 7400 810 7460 890
rect 7540 810 7600 890
rect 7400 750 7600 810
rect 7800 890 8000 950
rect 7800 810 7860 890
rect 7940 810 8000 890
rect 7800 750 8000 810
rect 8200 890 8400 950
rect 8200 810 8260 890
rect 8340 810 8400 890
rect 8200 750 8400 810
rect 8600 890 8800 950
rect 8600 810 8660 890
rect 8740 810 8800 890
rect 8600 750 8800 810
rect 9000 890 9200 950
rect 9000 810 9060 890
rect 9140 810 9200 890
rect 9000 750 9200 810
rect 9400 890 9600 950
rect 9400 810 9460 890
rect 9540 810 9600 890
rect 9400 750 9600 810
rect 9800 890 10000 950
rect 9800 810 9860 890
rect 9940 810 10000 890
rect 9800 750 10000 810
rect 2200 490 2400 550
rect 2200 410 2260 490
rect 2340 410 2400 490
rect 2200 350 2400 410
rect 2600 490 2800 550
rect 2600 410 2660 490
rect 2740 410 2800 490
rect 2600 350 2800 410
rect 3000 490 3200 550
rect 3000 410 3060 490
rect 3140 410 3200 490
rect 3000 350 3200 410
rect 3400 490 3600 550
rect 3400 410 3460 490
rect 3540 410 3600 490
rect 3400 350 3600 410
rect 3800 490 4000 550
rect 3800 410 3860 490
rect 3940 410 4000 490
rect 3800 350 4000 410
rect 4200 490 4400 550
rect 4200 410 4260 490
rect 4340 410 4400 490
rect 4200 350 4400 410
rect 4600 490 4800 550
rect 4600 410 4660 490
rect 4740 410 4800 490
rect 4600 350 4800 410
rect 5000 490 5200 550
rect 5000 410 5060 490
rect 5140 410 5200 490
rect 5000 350 5200 410
rect 5400 490 5600 550
rect 5400 410 5460 490
rect 5540 410 5600 490
rect 5400 350 5600 410
rect 5800 490 6000 550
rect 5800 410 5860 490
rect 5940 410 6000 490
rect 5800 350 6000 410
rect 6200 490 6400 550
rect 6200 410 6260 490
rect 6340 410 6400 490
rect 6200 350 6400 410
rect 6600 490 6800 550
rect 6600 410 6660 490
rect 6740 410 6800 490
rect 6600 350 6800 410
rect 7000 490 7200 550
rect 7000 410 7060 490
rect 7140 410 7200 490
rect 7000 350 7200 410
rect 7400 490 7600 550
rect 7400 410 7460 490
rect 7540 410 7600 490
rect 7400 350 7600 410
rect 7800 490 8000 550
rect 7800 410 7860 490
rect 7940 410 8000 490
rect 7800 350 8000 410
rect 8200 490 8400 550
rect 8200 410 8260 490
rect 8340 410 8400 490
rect 8200 350 8400 410
rect 8600 490 8800 550
rect 8600 410 8660 490
rect 8740 410 8800 490
rect 8600 350 8800 410
rect 9000 490 9200 550
rect 9000 410 9060 490
rect 9140 410 9200 490
rect 9000 350 9200 410
rect 9400 490 9600 550
rect 9400 410 9460 490
rect 9540 410 9600 490
rect 9400 350 9600 410
rect 9800 490 10000 550
rect 9800 410 9860 490
rect 9940 410 10000 490
rect 9800 350 10000 410
rect 10100 250 10350 8250
rect 1850 0 10350 250
<< m2contact >>
rect 2260 8010 2340 8090
rect 2660 8010 2740 8090
rect 3060 8010 3140 8090
rect 3460 8010 3540 8090
rect 3860 8010 3940 8090
rect 4260 8010 4340 8090
rect 4660 8010 4740 8090
rect 5060 8010 5140 8090
rect 5460 8010 5540 8090
rect 5860 8010 5940 8090
rect 6260 8010 6340 8090
rect 6660 8010 6740 8090
rect 7060 8010 7140 8090
rect 7460 8010 7540 8090
rect 7860 8010 7940 8090
rect 8260 8010 8340 8090
rect 8660 8010 8740 8090
rect 9060 8010 9140 8090
rect 9460 8010 9540 8090
rect 9860 8010 9940 8090
rect 2260 7610 2340 7690
rect 2660 7610 2740 7690
rect 3060 7610 3140 7690
rect 3460 7610 3540 7690
rect 3860 7610 3940 7690
rect 4260 7610 4340 7690
rect 4660 7610 4740 7690
rect 5060 7610 5140 7690
rect 5460 7610 5540 7690
rect 5860 7610 5940 7690
rect 6260 7610 6340 7690
rect 6660 7610 6740 7690
rect 7060 7610 7140 7690
rect 7460 7610 7540 7690
rect 7860 7610 7940 7690
rect 8260 7610 8340 7690
rect 8660 7610 8740 7690
rect 9060 7610 9140 7690
rect 9460 7610 9540 7690
rect 9860 7610 9940 7690
rect 2260 7210 2340 7290
rect 2660 7210 2740 7290
rect 3060 7210 3140 7290
rect 3460 7210 3540 7290
rect 3860 7210 3940 7290
rect 4260 7210 4340 7290
rect 4660 7210 4740 7290
rect 5060 7210 5140 7290
rect 5460 7210 5540 7290
rect 5860 7210 5940 7290
rect 6260 7210 6340 7290
rect 6660 7210 6740 7290
rect 7060 7210 7140 7290
rect 7460 7210 7540 7290
rect 7860 7210 7940 7290
rect 8260 7210 8340 7290
rect 8660 7210 8740 7290
rect 9060 7210 9140 7290
rect 9460 7210 9540 7290
rect 9860 7210 9940 7290
rect 2260 6810 2340 6890
rect 2660 6810 2740 6890
rect 3060 6810 3140 6890
rect 3460 6810 3540 6890
rect 3860 6810 3940 6890
rect 4260 6810 4340 6890
rect 4660 6810 4740 6890
rect 5060 6810 5140 6890
rect 5460 6810 5540 6890
rect 5860 6810 5940 6890
rect 6260 6810 6340 6890
rect 6660 6810 6740 6890
rect 7060 6810 7140 6890
rect 7460 6810 7540 6890
rect 7860 6810 7940 6890
rect 8260 6810 8340 6890
rect 8660 6810 8740 6890
rect 9060 6810 9140 6890
rect 9460 6810 9540 6890
rect 9860 6810 9940 6890
rect 2260 6410 2340 6490
rect 2660 6410 2740 6490
rect 3060 6410 3140 6490
rect 3460 6410 3540 6490
rect 3860 6410 3940 6490
rect 4260 6410 4340 6490
rect 4660 6410 4740 6490
rect 5060 6410 5140 6490
rect 5460 6410 5540 6490
rect 5860 6410 5940 6490
rect 6260 6410 6340 6490
rect 6660 6410 6740 6490
rect 7060 6410 7140 6490
rect 7460 6410 7540 6490
rect 7860 6410 7940 6490
rect 8260 6410 8340 6490
rect 8660 6410 8740 6490
rect 9060 6410 9140 6490
rect 9460 6410 9540 6490
rect 9860 6410 9940 6490
rect 2260 6010 2340 6090
rect 2660 6010 2740 6090
rect 3060 6010 3140 6090
rect 3460 6010 3540 6090
rect 3860 6010 3940 6090
rect 4260 6010 4340 6090
rect 4660 6010 4740 6090
rect 5060 6010 5140 6090
rect 5460 6010 5540 6090
rect 5860 6010 5940 6090
rect 6260 6010 6340 6090
rect 6660 6010 6740 6090
rect 7060 6010 7140 6090
rect 7460 6010 7540 6090
rect 7860 6010 7940 6090
rect 8260 6010 8340 6090
rect 8660 6010 8740 6090
rect 9060 6010 9140 6090
rect 9460 6010 9540 6090
rect 9860 6010 9940 6090
rect 2260 5610 2340 5690
rect 2660 5610 2740 5690
rect 3060 5610 3140 5690
rect 3460 5610 3540 5690
rect 3860 5610 3940 5690
rect 4260 5610 4340 5690
rect 4660 5610 4740 5690
rect 5060 5610 5140 5690
rect 5460 5610 5540 5690
rect 5860 5610 5940 5690
rect 6260 5610 6340 5690
rect 6660 5610 6740 5690
rect 7060 5610 7140 5690
rect 7460 5610 7540 5690
rect 7860 5610 7940 5690
rect 8260 5610 8340 5690
rect 8660 5610 8740 5690
rect 9060 5610 9140 5690
rect 9460 5610 9540 5690
rect 9860 5610 9940 5690
rect 2260 5210 2340 5290
rect 2660 5210 2740 5290
rect 3060 5210 3140 5290
rect 3460 5210 3540 5290
rect 3860 5210 3940 5290
rect 4260 5210 4340 5290
rect 4660 5210 4740 5290
rect 5060 5210 5140 5290
rect 5460 5210 5540 5290
rect 5860 5210 5940 5290
rect 6260 5210 6340 5290
rect 6660 5210 6740 5290
rect 7060 5210 7140 5290
rect 7460 5210 7540 5290
rect 7860 5210 7940 5290
rect 8260 5210 8340 5290
rect 8660 5210 8740 5290
rect 9060 5210 9140 5290
rect 9460 5210 9540 5290
rect 9860 5210 9940 5290
rect 2260 4810 2340 4890
rect 2660 4810 2740 4890
rect 3060 4810 3140 4890
rect 3460 4810 3540 4890
rect 3860 4810 3940 4890
rect 4260 4810 4340 4890
rect 4660 4810 4740 4890
rect 5060 4810 5140 4890
rect 5460 4810 5540 4890
rect 5860 4810 5940 4890
rect 6260 4810 6340 4890
rect 6660 4810 6740 4890
rect 7060 4810 7140 4890
rect 7460 4810 7540 4890
rect 7860 4810 7940 4890
rect 8260 4810 8340 4890
rect 8660 4810 8740 4890
rect 9060 4810 9140 4890
rect 9460 4810 9540 4890
rect 9860 4810 9940 4890
rect 2260 4410 2340 4490
rect 2660 4410 2740 4490
rect 3060 4410 3140 4490
rect 3460 4410 3540 4490
rect 3860 4410 3940 4490
rect 4260 4410 4340 4490
rect 4660 4410 4740 4490
rect 5060 4410 5140 4490
rect 5460 4410 5540 4490
rect 5860 4410 5940 4490
rect 6260 4410 6340 4490
rect 6660 4410 6740 4490
rect 7060 4410 7140 4490
rect 7460 4410 7540 4490
rect 7860 4410 7940 4490
rect 8260 4410 8340 4490
rect 8660 4410 8740 4490
rect 9060 4410 9140 4490
rect 9460 4410 9540 4490
rect 9860 4410 9940 4490
rect 2260 4010 2340 4090
rect 2660 4010 2740 4090
rect 3060 4010 3140 4090
rect 3460 4010 3540 4090
rect 3860 4010 3940 4090
rect 4260 4010 4340 4090
rect 4660 4010 4740 4090
rect 5060 4010 5140 4090
rect 5460 4010 5540 4090
rect 5860 4010 5940 4090
rect 6260 4010 6340 4090
rect 6660 4010 6740 4090
rect 7060 4010 7140 4090
rect 7460 4010 7540 4090
rect 7860 4010 7940 4090
rect 8260 4010 8340 4090
rect 8660 4010 8740 4090
rect 9060 4010 9140 4090
rect 9460 4010 9540 4090
rect 9860 4010 9940 4090
rect 2260 3610 2340 3690
rect 2660 3610 2740 3690
rect 3060 3610 3140 3690
rect 3460 3610 3540 3690
rect 3860 3610 3940 3690
rect 4260 3610 4340 3690
rect 4660 3610 4740 3690
rect 5060 3610 5140 3690
rect 5460 3610 5540 3690
rect 5860 3610 5940 3690
rect 6260 3610 6340 3690
rect 6660 3610 6740 3690
rect 7060 3610 7140 3690
rect 7460 3610 7540 3690
rect 7860 3610 7940 3690
rect 8260 3610 8340 3690
rect 8660 3610 8740 3690
rect 9060 3610 9140 3690
rect 9460 3610 9540 3690
rect 9860 3610 9940 3690
rect 2260 3210 2340 3290
rect 2660 3210 2740 3290
rect 3060 3210 3140 3290
rect 3460 3210 3540 3290
rect 3860 3210 3940 3290
rect 4260 3210 4340 3290
rect 4660 3210 4740 3290
rect 5060 3210 5140 3290
rect 5460 3210 5540 3290
rect 5860 3210 5940 3290
rect 6260 3210 6340 3290
rect 6660 3210 6740 3290
rect 7060 3210 7140 3290
rect 7460 3210 7540 3290
rect 7860 3210 7940 3290
rect 8260 3210 8340 3290
rect 8660 3210 8740 3290
rect 9060 3210 9140 3290
rect 9460 3210 9540 3290
rect 9860 3210 9940 3290
rect 2260 2810 2340 2890
rect 2660 2810 2740 2890
rect 3060 2810 3140 2890
rect 3460 2810 3540 2890
rect 3860 2810 3940 2890
rect 4260 2810 4340 2890
rect 4660 2810 4740 2890
rect 5060 2810 5140 2890
rect 5460 2810 5540 2890
rect 5860 2810 5940 2890
rect 6260 2810 6340 2890
rect 6660 2810 6740 2890
rect 7060 2810 7140 2890
rect 7460 2810 7540 2890
rect 7860 2810 7940 2890
rect 8260 2810 8340 2890
rect 8660 2810 8740 2890
rect 9060 2810 9140 2890
rect 9460 2810 9540 2890
rect 9860 2810 9940 2890
rect 2260 2410 2340 2490
rect 2660 2410 2740 2490
rect 3060 2410 3140 2490
rect 3460 2410 3540 2490
rect 3860 2410 3940 2490
rect 4260 2410 4340 2490
rect 4660 2410 4740 2490
rect 5060 2410 5140 2490
rect 5460 2410 5540 2490
rect 5860 2410 5940 2490
rect 6260 2410 6340 2490
rect 6660 2410 6740 2490
rect 7060 2410 7140 2490
rect 7460 2410 7540 2490
rect 7860 2410 7940 2490
rect 8260 2410 8340 2490
rect 8660 2410 8740 2490
rect 9060 2410 9140 2490
rect 9460 2410 9540 2490
rect 9860 2410 9940 2490
rect 2260 2010 2340 2090
rect 2660 2010 2740 2090
rect 3060 2010 3140 2090
rect 3460 2010 3540 2090
rect 3860 2010 3940 2090
rect 4260 2010 4340 2090
rect 4660 2010 4740 2090
rect 5060 2010 5140 2090
rect 5460 2010 5540 2090
rect 5860 2010 5940 2090
rect 6260 2010 6340 2090
rect 6660 2010 6740 2090
rect 7060 2010 7140 2090
rect 7460 2010 7540 2090
rect 7860 2010 7940 2090
rect 8260 2010 8340 2090
rect 8660 2010 8740 2090
rect 9060 2010 9140 2090
rect 9460 2010 9540 2090
rect 9860 2010 9940 2090
rect 2260 1610 2340 1690
rect 2660 1610 2740 1690
rect 3060 1610 3140 1690
rect 3460 1610 3540 1690
rect 3860 1610 3940 1690
rect 4260 1610 4340 1690
rect 4660 1610 4740 1690
rect 5060 1610 5140 1690
rect 5460 1610 5540 1690
rect 5860 1610 5940 1690
rect 6260 1610 6340 1690
rect 6660 1610 6740 1690
rect 7060 1610 7140 1690
rect 7460 1610 7540 1690
rect 7860 1610 7940 1690
rect 8260 1610 8340 1690
rect 8660 1610 8740 1690
rect 9060 1610 9140 1690
rect 9460 1610 9540 1690
rect 9860 1610 9940 1690
rect 2260 1210 2340 1290
rect 2660 1210 2740 1290
rect 3060 1210 3140 1290
rect 3460 1210 3540 1290
rect 3860 1210 3940 1290
rect 4260 1210 4340 1290
rect 4660 1210 4740 1290
rect 5060 1210 5140 1290
rect 5460 1210 5540 1290
rect 5860 1210 5940 1290
rect 6260 1210 6340 1290
rect 6660 1210 6740 1290
rect 7060 1210 7140 1290
rect 7460 1210 7540 1290
rect 7860 1210 7940 1290
rect 8260 1210 8340 1290
rect 8660 1210 8740 1290
rect 9060 1210 9140 1290
rect 9460 1210 9540 1290
rect 9860 1210 9940 1290
rect 2260 810 2340 890
rect 2660 810 2740 890
rect 3060 810 3140 890
rect 3460 810 3540 890
rect 3860 810 3940 890
rect 4260 810 4340 890
rect 4660 810 4740 890
rect 5060 810 5140 890
rect 5460 810 5540 890
rect 5860 810 5940 890
rect 6260 810 6340 890
rect 6660 810 6740 890
rect 7060 810 7140 890
rect 7460 810 7540 890
rect 7860 810 7940 890
rect 8260 810 8340 890
rect 8660 810 8740 890
rect 9060 810 9140 890
rect 9460 810 9540 890
rect 9860 810 9940 890
rect 2260 410 2340 490
rect 2660 410 2740 490
rect 3060 410 3140 490
rect 3460 410 3540 490
rect 3860 410 3940 490
rect 4260 410 4340 490
rect 4660 410 4740 490
rect 5060 410 5140 490
rect 5460 410 5540 490
rect 5860 410 5940 490
rect 6260 410 6340 490
rect 6660 410 6740 490
rect 7060 410 7140 490
rect 7460 410 7540 490
rect 7860 410 7940 490
rect 8260 410 8340 490
rect 8660 410 8740 490
rect 9060 410 9140 490
rect 9460 410 9540 490
rect 9860 410 9940 490
<< metal2 >>
rect 100 32550 12100 34210
rect 100 30250 12100 31910
rect 100 20450 12100 28250
rect 100 9150 12100 16950
rect 1850 8250 10350 8500
rect 1850 250 2100 8250
rect 2200 8090 2400 8150
rect 2200 8010 2260 8090
rect 2340 8010 2400 8090
rect 2200 7950 2400 8010
rect 2600 8090 2800 8150
rect 2600 8010 2660 8090
rect 2740 8010 2800 8090
rect 2600 7950 2800 8010
rect 3000 8090 3200 8150
rect 3000 8010 3060 8090
rect 3140 8010 3200 8090
rect 3000 7950 3200 8010
rect 3400 8090 3600 8150
rect 3400 8010 3460 8090
rect 3540 8010 3600 8090
rect 3400 7950 3600 8010
rect 3800 8090 4000 8150
rect 3800 8010 3860 8090
rect 3940 8010 4000 8090
rect 3800 7950 4000 8010
rect 4200 8090 4400 8150
rect 4200 8010 4260 8090
rect 4340 8010 4400 8090
rect 4200 7950 4400 8010
rect 4600 8090 4800 8150
rect 4600 8010 4660 8090
rect 4740 8010 4800 8090
rect 4600 7950 4800 8010
rect 5000 8090 5200 8150
rect 5000 8010 5060 8090
rect 5140 8010 5200 8090
rect 5000 7950 5200 8010
rect 5400 8090 5600 8150
rect 5400 8010 5460 8090
rect 5540 8010 5600 8090
rect 5400 7950 5600 8010
rect 5800 8090 6000 8150
rect 5800 8010 5860 8090
rect 5940 8010 6000 8090
rect 5800 7950 6000 8010
rect 6200 8090 6400 8150
rect 6200 8010 6260 8090
rect 6340 8010 6400 8090
rect 6200 7950 6400 8010
rect 6600 8090 6800 8150
rect 6600 8010 6660 8090
rect 6740 8010 6800 8090
rect 6600 7950 6800 8010
rect 7000 8090 7200 8150
rect 7000 8010 7060 8090
rect 7140 8010 7200 8090
rect 7000 7950 7200 8010
rect 7400 8090 7600 8150
rect 7400 8010 7460 8090
rect 7540 8010 7600 8090
rect 7400 7950 7600 8010
rect 7800 8090 8000 8150
rect 7800 8010 7860 8090
rect 7940 8010 8000 8090
rect 7800 7950 8000 8010
rect 8200 8090 8400 8150
rect 8200 8010 8260 8090
rect 8340 8010 8400 8090
rect 8200 7950 8400 8010
rect 8600 8090 8800 8150
rect 8600 8010 8660 8090
rect 8740 8010 8800 8090
rect 8600 7950 8800 8010
rect 9000 8090 9200 8150
rect 9000 8010 9060 8090
rect 9140 8010 9200 8090
rect 9000 7950 9200 8010
rect 9400 8090 9600 8150
rect 9400 8010 9460 8090
rect 9540 8010 9600 8090
rect 9400 7950 9600 8010
rect 9800 8090 10000 8150
rect 9800 8010 9860 8090
rect 9940 8010 10000 8090
rect 9800 7950 10000 8010
rect 2400 7890 2600 7950
rect 2400 7810 2460 7890
rect 2540 7810 2600 7890
rect 2400 7750 2600 7810
rect 2800 7890 3000 7950
rect 2800 7810 2860 7890
rect 2940 7810 3000 7890
rect 2800 7750 3000 7810
rect 3200 7890 3400 7950
rect 3200 7810 3260 7890
rect 3340 7810 3400 7890
rect 3200 7750 3400 7810
rect 3600 7890 3800 7950
rect 3600 7810 3660 7890
rect 3740 7810 3800 7890
rect 3600 7750 3800 7810
rect 4000 7890 4200 7950
rect 4000 7810 4060 7890
rect 4140 7810 4200 7890
rect 4000 7750 4200 7810
rect 4400 7890 4600 7950
rect 4400 7810 4460 7890
rect 4540 7810 4600 7890
rect 4400 7750 4600 7810
rect 4800 7890 5000 7950
rect 4800 7810 4860 7890
rect 4940 7810 5000 7890
rect 4800 7750 5000 7810
rect 5200 7890 5400 7950
rect 5200 7810 5260 7890
rect 5340 7810 5400 7890
rect 5200 7750 5400 7810
rect 5600 7890 5800 7950
rect 5600 7810 5660 7890
rect 5740 7810 5800 7890
rect 5600 7750 5800 7810
rect 6000 7890 6200 7950
rect 6000 7810 6060 7890
rect 6140 7810 6200 7890
rect 6000 7750 6200 7810
rect 6400 7890 6600 7950
rect 6400 7810 6460 7890
rect 6540 7810 6600 7890
rect 6400 7750 6600 7810
rect 6800 7890 7000 7950
rect 6800 7810 6860 7890
rect 6940 7810 7000 7890
rect 6800 7750 7000 7810
rect 7200 7890 7400 7950
rect 7200 7810 7260 7890
rect 7340 7810 7400 7890
rect 7200 7750 7400 7810
rect 7600 7890 7800 7950
rect 7600 7810 7660 7890
rect 7740 7810 7800 7890
rect 7600 7750 7800 7810
rect 8000 7890 8200 7950
rect 8000 7810 8060 7890
rect 8140 7810 8200 7890
rect 8000 7750 8200 7810
rect 8400 7890 8600 7950
rect 8400 7810 8460 7890
rect 8540 7810 8600 7890
rect 8400 7750 8600 7810
rect 8800 7890 9000 7950
rect 8800 7810 8860 7890
rect 8940 7810 9000 7890
rect 8800 7750 9000 7810
rect 9200 7890 9400 7950
rect 9200 7810 9260 7890
rect 9340 7810 9400 7890
rect 9200 7750 9400 7810
rect 9600 7890 9800 7950
rect 9600 7810 9660 7890
rect 9740 7810 9800 7890
rect 9600 7750 9800 7810
rect 2200 7690 2400 7750
rect 2200 7610 2260 7690
rect 2340 7610 2400 7690
rect 2200 7550 2400 7610
rect 2600 7690 2800 7750
rect 2600 7610 2660 7690
rect 2740 7610 2800 7690
rect 2600 7550 2800 7610
rect 3000 7690 3200 7750
rect 3000 7610 3060 7690
rect 3140 7610 3200 7690
rect 3000 7550 3200 7610
rect 3400 7690 3600 7750
rect 3400 7610 3460 7690
rect 3540 7610 3600 7690
rect 3400 7550 3600 7610
rect 3800 7690 4000 7750
rect 3800 7610 3860 7690
rect 3940 7610 4000 7690
rect 3800 7550 4000 7610
rect 4200 7690 4400 7750
rect 4200 7610 4260 7690
rect 4340 7610 4400 7690
rect 4200 7550 4400 7610
rect 4600 7690 4800 7750
rect 4600 7610 4660 7690
rect 4740 7610 4800 7690
rect 4600 7550 4800 7610
rect 5000 7690 5200 7750
rect 5000 7610 5060 7690
rect 5140 7610 5200 7690
rect 5000 7550 5200 7610
rect 5400 7690 5600 7750
rect 5400 7610 5460 7690
rect 5540 7610 5600 7690
rect 5400 7550 5600 7610
rect 5800 7690 6000 7750
rect 5800 7610 5860 7690
rect 5940 7610 6000 7690
rect 5800 7550 6000 7610
rect 6200 7690 6400 7750
rect 6200 7610 6260 7690
rect 6340 7610 6400 7690
rect 6200 7550 6400 7610
rect 6600 7690 6800 7750
rect 6600 7610 6660 7690
rect 6740 7610 6800 7690
rect 6600 7550 6800 7610
rect 7000 7690 7200 7750
rect 7000 7610 7060 7690
rect 7140 7610 7200 7690
rect 7000 7550 7200 7610
rect 7400 7690 7600 7750
rect 7400 7610 7460 7690
rect 7540 7610 7600 7690
rect 7400 7550 7600 7610
rect 7800 7690 8000 7750
rect 7800 7610 7860 7690
rect 7940 7610 8000 7690
rect 7800 7550 8000 7610
rect 8200 7690 8400 7750
rect 8200 7610 8260 7690
rect 8340 7610 8400 7690
rect 8200 7550 8400 7610
rect 8600 7690 8800 7750
rect 8600 7610 8660 7690
rect 8740 7610 8800 7690
rect 8600 7550 8800 7610
rect 9000 7690 9200 7750
rect 9000 7610 9060 7690
rect 9140 7610 9200 7690
rect 9000 7550 9200 7610
rect 9400 7690 9600 7750
rect 9400 7610 9460 7690
rect 9540 7610 9600 7690
rect 9400 7550 9600 7610
rect 9800 7690 10000 7750
rect 9800 7610 9860 7690
rect 9940 7610 10000 7690
rect 9800 7550 10000 7610
rect 2400 7490 2600 7550
rect 2400 7410 2460 7490
rect 2540 7410 2600 7490
rect 2400 7350 2600 7410
rect 2800 7490 3000 7550
rect 2800 7410 2860 7490
rect 2940 7410 3000 7490
rect 2800 7350 3000 7410
rect 3200 7490 3400 7550
rect 3200 7410 3260 7490
rect 3340 7410 3400 7490
rect 3200 7350 3400 7410
rect 3600 7490 3800 7550
rect 3600 7410 3660 7490
rect 3740 7410 3800 7490
rect 3600 7350 3800 7410
rect 4000 7490 4200 7550
rect 4000 7410 4060 7490
rect 4140 7410 4200 7490
rect 4000 7350 4200 7410
rect 4400 7490 4600 7550
rect 4400 7410 4460 7490
rect 4540 7410 4600 7490
rect 4400 7350 4600 7410
rect 4800 7490 5000 7550
rect 4800 7410 4860 7490
rect 4940 7410 5000 7490
rect 4800 7350 5000 7410
rect 5200 7490 5400 7550
rect 5200 7410 5260 7490
rect 5340 7410 5400 7490
rect 5200 7350 5400 7410
rect 5600 7490 5800 7550
rect 5600 7410 5660 7490
rect 5740 7410 5800 7490
rect 5600 7350 5800 7410
rect 6000 7490 6200 7550
rect 6000 7410 6060 7490
rect 6140 7410 6200 7490
rect 6000 7350 6200 7410
rect 6400 7490 6600 7550
rect 6400 7410 6460 7490
rect 6540 7410 6600 7490
rect 6400 7350 6600 7410
rect 6800 7490 7000 7550
rect 6800 7410 6860 7490
rect 6940 7410 7000 7490
rect 6800 7350 7000 7410
rect 7200 7490 7400 7550
rect 7200 7410 7260 7490
rect 7340 7410 7400 7490
rect 7200 7350 7400 7410
rect 7600 7490 7800 7550
rect 7600 7410 7660 7490
rect 7740 7410 7800 7490
rect 7600 7350 7800 7410
rect 8000 7490 8200 7550
rect 8000 7410 8060 7490
rect 8140 7410 8200 7490
rect 8000 7350 8200 7410
rect 8400 7490 8600 7550
rect 8400 7410 8460 7490
rect 8540 7410 8600 7490
rect 8400 7350 8600 7410
rect 8800 7490 9000 7550
rect 8800 7410 8860 7490
rect 8940 7410 9000 7490
rect 8800 7350 9000 7410
rect 9200 7490 9400 7550
rect 9200 7410 9260 7490
rect 9340 7410 9400 7490
rect 9200 7350 9400 7410
rect 9600 7490 9800 7550
rect 9600 7410 9660 7490
rect 9740 7410 9800 7490
rect 9600 7350 9800 7410
rect 2200 7290 2400 7350
rect 2200 7210 2260 7290
rect 2340 7210 2400 7290
rect 2200 7150 2400 7210
rect 2600 7290 2800 7350
rect 2600 7210 2660 7290
rect 2740 7210 2800 7290
rect 2600 7150 2800 7210
rect 3000 7290 3200 7350
rect 3000 7210 3060 7290
rect 3140 7210 3200 7290
rect 3000 7150 3200 7210
rect 3400 7290 3600 7350
rect 3400 7210 3460 7290
rect 3540 7210 3600 7290
rect 3400 7150 3600 7210
rect 3800 7290 4000 7350
rect 3800 7210 3860 7290
rect 3940 7210 4000 7290
rect 3800 7150 4000 7210
rect 4200 7290 4400 7350
rect 4200 7210 4260 7290
rect 4340 7210 4400 7290
rect 4200 7150 4400 7210
rect 4600 7290 4800 7350
rect 4600 7210 4660 7290
rect 4740 7210 4800 7290
rect 4600 7150 4800 7210
rect 5000 7290 5200 7350
rect 5000 7210 5060 7290
rect 5140 7210 5200 7290
rect 5000 7150 5200 7210
rect 5400 7290 5600 7350
rect 5400 7210 5460 7290
rect 5540 7210 5600 7290
rect 5400 7150 5600 7210
rect 5800 7290 6000 7350
rect 5800 7210 5860 7290
rect 5940 7210 6000 7290
rect 5800 7150 6000 7210
rect 6200 7290 6400 7350
rect 6200 7210 6260 7290
rect 6340 7210 6400 7290
rect 6200 7150 6400 7210
rect 6600 7290 6800 7350
rect 6600 7210 6660 7290
rect 6740 7210 6800 7290
rect 6600 7150 6800 7210
rect 7000 7290 7200 7350
rect 7000 7210 7060 7290
rect 7140 7210 7200 7290
rect 7000 7150 7200 7210
rect 7400 7290 7600 7350
rect 7400 7210 7460 7290
rect 7540 7210 7600 7290
rect 7400 7150 7600 7210
rect 7800 7290 8000 7350
rect 7800 7210 7860 7290
rect 7940 7210 8000 7290
rect 7800 7150 8000 7210
rect 8200 7290 8400 7350
rect 8200 7210 8260 7290
rect 8340 7210 8400 7290
rect 8200 7150 8400 7210
rect 8600 7290 8800 7350
rect 8600 7210 8660 7290
rect 8740 7210 8800 7290
rect 8600 7150 8800 7210
rect 9000 7290 9200 7350
rect 9000 7210 9060 7290
rect 9140 7210 9200 7290
rect 9000 7150 9200 7210
rect 9400 7290 9600 7350
rect 9400 7210 9460 7290
rect 9540 7210 9600 7290
rect 9400 7150 9600 7210
rect 9800 7290 10000 7350
rect 9800 7210 9860 7290
rect 9940 7210 10000 7290
rect 9800 7150 10000 7210
rect 2400 7090 2600 7150
rect 2400 7010 2460 7090
rect 2540 7010 2600 7090
rect 2400 6950 2600 7010
rect 2800 7090 3000 7150
rect 2800 7010 2860 7090
rect 2940 7010 3000 7090
rect 2800 6950 3000 7010
rect 3200 7090 3400 7150
rect 3200 7010 3260 7090
rect 3340 7010 3400 7090
rect 3200 6950 3400 7010
rect 3600 7090 3800 7150
rect 3600 7010 3660 7090
rect 3740 7010 3800 7090
rect 3600 6950 3800 7010
rect 4000 7090 4200 7150
rect 4000 7010 4060 7090
rect 4140 7010 4200 7090
rect 4000 6950 4200 7010
rect 4400 7090 4600 7150
rect 4400 7010 4460 7090
rect 4540 7010 4600 7090
rect 4400 6950 4600 7010
rect 4800 7090 5000 7150
rect 4800 7010 4860 7090
rect 4940 7010 5000 7090
rect 4800 6950 5000 7010
rect 5200 7090 5400 7150
rect 5200 7010 5260 7090
rect 5340 7010 5400 7090
rect 5200 6950 5400 7010
rect 5600 7090 5800 7150
rect 5600 7010 5660 7090
rect 5740 7010 5800 7090
rect 5600 6950 5800 7010
rect 6000 7090 6200 7150
rect 6000 7010 6060 7090
rect 6140 7010 6200 7090
rect 6000 6950 6200 7010
rect 6400 7090 6600 7150
rect 6400 7010 6460 7090
rect 6540 7010 6600 7090
rect 6400 6950 6600 7010
rect 6800 7090 7000 7150
rect 6800 7010 6860 7090
rect 6940 7010 7000 7090
rect 6800 6950 7000 7010
rect 7200 7090 7400 7150
rect 7200 7010 7260 7090
rect 7340 7010 7400 7090
rect 7200 6950 7400 7010
rect 7600 7090 7800 7150
rect 7600 7010 7660 7090
rect 7740 7010 7800 7090
rect 7600 6950 7800 7010
rect 8000 7090 8200 7150
rect 8000 7010 8060 7090
rect 8140 7010 8200 7090
rect 8000 6950 8200 7010
rect 8400 7090 8600 7150
rect 8400 7010 8460 7090
rect 8540 7010 8600 7090
rect 8400 6950 8600 7010
rect 8800 7090 9000 7150
rect 8800 7010 8860 7090
rect 8940 7010 9000 7090
rect 8800 6950 9000 7010
rect 9200 7090 9400 7150
rect 9200 7010 9260 7090
rect 9340 7010 9400 7090
rect 9200 6950 9400 7010
rect 9600 7090 9800 7150
rect 9600 7010 9660 7090
rect 9740 7010 9800 7090
rect 9600 6950 9800 7010
rect 2200 6890 2400 6950
rect 2200 6810 2260 6890
rect 2340 6810 2400 6890
rect 2200 6750 2400 6810
rect 2600 6890 2800 6950
rect 2600 6810 2660 6890
rect 2740 6810 2800 6890
rect 2600 6750 2800 6810
rect 3000 6890 3200 6950
rect 3000 6810 3060 6890
rect 3140 6810 3200 6890
rect 3000 6750 3200 6810
rect 3400 6890 3600 6950
rect 3400 6810 3460 6890
rect 3540 6810 3600 6890
rect 3400 6750 3600 6810
rect 3800 6890 4000 6950
rect 3800 6810 3860 6890
rect 3940 6810 4000 6890
rect 3800 6750 4000 6810
rect 4200 6890 4400 6950
rect 4200 6810 4260 6890
rect 4340 6810 4400 6890
rect 4200 6750 4400 6810
rect 4600 6890 4800 6950
rect 4600 6810 4660 6890
rect 4740 6810 4800 6890
rect 4600 6750 4800 6810
rect 5000 6890 5200 6950
rect 5000 6810 5060 6890
rect 5140 6810 5200 6890
rect 5000 6750 5200 6810
rect 5400 6890 5600 6950
rect 5400 6810 5460 6890
rect 5540 6810 5600 6890
rect 5400 6750 5600 6810
rect 5800 6890 6000 6950
rect 5800 6810 5860 6890
rect 5940 6810 6000 6890
rect 5800 6750 6000 6810
rect 6200 6890 6400 6950
rect 6200 6810 6260 6890
rect 6340 6810 6400 6890
rect 6200 6750 6400 6810
rect 6600 6890 6800 6950
rect 6600 6810 6660 6890
rect 6740 6810 6800 6890
rect 6600 6750 6800 6810
rect 7000 6890 7200 6950
rect 7000 6810 7060 6890
rect 7140 6810 7200 6890
rect 7000 6750 7200 6810
rect 7400 6890 7600 6950
rect 7400 6810 7460 6890
rect 7540 6810 7600 6890
rect 7400 6750 7600 6810
rect 7800 6890 8000 6950
rect 7800 6810 7860 6890
rect 7940 6810 8000 6890
rect 7800 6750 8000 6810
rect 8200 6890 8400 6950
rect 8200 6810 8260 6890
rect 8340 6810 8400 6890
rect 8200 6750 8400 6810
rect 8600 6890 8800 6950
rect 8600 6810 8660 6890
rect 8740 6810 8800 6890
rect 8600 6750 8800 6810
rect 9000 6890 9200 6950
rect 9000 6810 9060 6890
rect 9140 6810 9200 6890
rect 9000 6750 9200 6810
rect 9400 6890 9600 6950
rect 9400 6810 9460 6890
rect 9540 6810 9600 6890
rect 9400 6750 9600 6810
rect 9800 6890 10000 6950
rect 9800 6810 9860 6890
rect 9940 6810 10000 6890
rect 9800 6750 10000 6810
rect 2400 6690 2600 6750
rect 2400 6610 2460 6690
rect 2540 6610 2600 6690
rect 2400 6550 2600 6610
rect 2800 6690 3000 6750
rect 2800 6610 2860 6690
rect 2940 6610 3000 6690
rect 2800 6550 3000 6610
rect 3200 6690 3400 6750
rect 3200 6610 3260 6690
rect 3340 6610 3400 6690
rect 3200 6550 3400 6610
rect 3600 6690 3800 6750
rect 3600 6610 3660 6690
rect 3740 6610 3800 6690
rect 3600 6550 3800 6610
rect 4000 6690 4200 6750
rect 4000 6610 4060 6690
rect 4140 6610 4200 6690
rect 4000 6550 4200 6610
rect 4400 6690 4600 6750
rect 4400 6610 4460 6690
rect 4540 6610 4600 6690
rect 4400 6550 4600 6610
rect 4800 6690 5000 6750
rect 4800 6610 4860 6690
rect 4940 6610 5000 6690
rect 4800 6550 5000 6610
rect 5200 6690 5400 6750
rect 5200 6610 5260 6690
rect 5340 6610 5400 6690
rect 5200 6550 5400 6610
rect 5600 6690 5800 6750
rect 5600 6610 5660 6690
rect 5740 6610 5800 6690
rect 5600 6550 5800 6610
rect 6000 6690 6200 6750
rect 6000 6610 6060 6690
rect 6140 6610 6200 6690
rect 6000 6550 6200 6610
rect 6400 6690 6600 6750
rect 6400 6610 6460 6690
rect 6540 6610 6600 6690
rect 6400 6550 6600 6610
rect 6800 6690 7000 6750
rect 6800 6610 6860 6690
rect 6940 6610 7000 6690
rect 6800 6550 7000 6610
rect 7200 6690 7400 6750
rect 7200 6610 7260 6690
rect 7340 6610 7400 6690
rect 7200 6550 7400 6610
rect 7600 6690 7800 6750
rect 7600 6610 7660 6690
rect 7740 6610 7800 6690
rect 7600 6550 7800 6610
rect 8000 6690 8200 6750
rect 8000 6610 8060 6690
rect 8140 6610 8200 6690
rect 8000 6550 8200 6610
rect 8400 6690 8600 6750
rect 8400 6610 8460 6690
rect 8540 6610 8600 6690
rect 8400 6550 8600 6610
rect 8800 6690 9000 6750
rect 8800 6610 8860 6690
rect 8940 6610 9000 6690
rect 8800 6550 9000 6610
rect 9200 6690 9400 6750
rect 9200 6610 9260 6690
rect 9340 6610 9400 6690
rect 9200 6550 9400 6610
rect 9600 6690 9800 6750
rect 9600 6610 9660 6690
rect 9740 6610 9800 6690
rect 9600 6550 9800 6610
rect 2200 6490 2400 6550
rect 2200 6410 2260 6490
rect 2340 6410 2400 6490
rect 2200 6350 2400 6410
rect 2600 6490 2800 6550
rect 2600 6410 2660 6490
rect 2740 6410 2800 6490
rect 2600 6350 2800 6410
rect 3000 6490 3200 6550
rect 3000 6410 3060 6490
rect 3140 6410 3200 6490
rect 3000 6350 3200 6410
rect 3400 6490 3600 6550
rect 3400 6410 3460 6490
rect 3540 6410 3600 6490
rect 3400 6350 3600 6410
rect 3800 6490 4000 6550
rect 3800 6410 3860 6490
rect 3940 6410 4000 6490
rect 3800 6350 4000 6410
rect 4200 6490 4400 6550
rect 4200 6410 4260 6490
rect 4340 6410 4400 6490
rect 4200 6350 4400 6410
rect 4600 6490 4800 6550
rect 4600 6410 4660 6490
rect 4740 6410 4800 6490
rect 4600 6350 4800 6410
rect 5000 6490 5200 6550
rect 5000 6410 5060 6490
rect 5140 6410 5200 6490
rect 5000 6350 5200 6410
rect 5400 6490 5600 6550
rect 5400 6410 5460 6490
rect 5540 6410 5600 6490
rect 5400 6350 5600 6410
rect 5800 6490 6000 6550
rect 5800 6410 5860 6490
rect 5940 6410 6000 6490
rect 5800 6350 6000 6410
rect 6200 6490 6400 6550
rect 6200 6410 6260 6490
rect 6340 6410 6400 6490
rect 6200 6350 6400 6410
rect 6600 6490 6800 6550
rect 6600 6410 6660 6490
rect 6740 6410 6800 6490
rect 6600 6350 6800 6410
rect 7000 6490 7200 6550
rect 7000 6410 7060 6490
rect 7140 6410 7200 6490
rect 7000 6350 7200 6410
rect 7400 6490 7600 6550
rect 7400 6410 7460 6490
rect 7540 6410 7600 6490
rect 7400 6350 7600 6410
rect 7800 6490 8000 6550
rect 7800 6410 7860 6490
rect 7940 6410 8000 6490
rect 7800 6350 8000 6410
rect 8200 6490 8400 6550
rect 8200 6410 8260 6490
rect 8340 6410 8400 6490
rect 8200 6350 8400 6410
rect 8600 6490 8800 6550
rect 8600 6410 8660 6490
rect 8740 6410 8800 6490
rect 8600 6350 8800 6410
rect 9000 6490 9200 6550
rect 9000 6410 9060 6490
rect 9140 6410 9200 6490
rect 9000 6350 9200 6410
rect 9400 6490 9600 6550
rect 9400 6410 9460 6490
rect 9540 6410 9600 6490
rect 9400 6350 9600 6410
rect 9800 6490 10000 6550
rect 9800 6410 9860 6490
rect 9940 6410 10000 6490
rect 9800 6350 10000 6410
rect 2400 6290 2600 6350
rect 2400 6210 2460 6290
rect 2540 6210 2600 6290
rect 2400 6150 2600 6210
rect 2800 6290 3000 6350
rect 2800 6210 2860 6290
rect 2940 6210 3000 6290
rect 2800 6150 3000 6210
rect 3200 6290 3400 6350
rect 3200 6210 3260 6290
rect 3340 6210 3400 6290
rect 3200 6150 3400 6210
rect 3600 6290 3800 6350
rect 3600 6210 3660 6290
rect 3740 6210 3800 6290
rect 3600 6150 3800 6210
rect 4000 6290 4200 6350
rect 4000 6210 4060 6290
rect 4140 6210 4200 6290
rect 4000 6150 4200 6210
rect 4400 6290 4600 6350
rect 4400 6210 4460 6290
rect 4540 6210 4600 6290
rect 4400 6150 4600 6210
rect 4800 6290 5000 6350
rect 4800 6210 4860 6290
rect 4940 6210 5000 6290
rect 4800 6150 5000 6210
rect 5200 6290 5400 6350
rect 5200 6210 5260 6290
rect 5340 6210 5400 6290
rect 5200 6150 5400 6210
rect 5600 6290 5800 6350
rect 5600 6210 5660 6290
rect 5740 6210 5800 6290
rect 5600 6150 5800 6210
rect 6000 6290 6200 6350
rect 6000 6210 6060 6290
rect 6140 6210 6200 6290
rect 6000 6150 6200 6210
rect 6400 6290 6600 6350
rect 6400 6210 6460 6290
rect 6540 6210 6600 6290
rect 6400 6150 6600 6210
rect 6800 6290 7000 6350
rect 6800 6210 6860 6290
rect 6940 6210 7000 6290
rect 6800 6150 7000 6210
rect 7200 6290 7400 6350
rect 7200 6210 7260 6290
rect 7340 6210 7400 6290
rect 7200 6150 7400 6210
rect 7600 6290 7800 6350
rect 7600 6210 7660 6290
rect 7740 6210 7800 6290
rect 7600 6150 7800 6210
rect 8000 6290 8200 6350
rect 8000 6210 8060 6290
rect 8140 6210 8200 6290
rect 8000 6150 8200 6210
rect 8400 6290 8600 6350
rect 8400 6210 8460 6290
rect 8540 6210 8600 6290
rect 8400 6150 8600 6210
rect 8800 6290 9000 6350
rect 8800 6210 8860 6290
rect 8940 6210 9000 6290
rect 8800 6150 9000 6210
rect 9200 6290 9400 6350
rect 9200 6210 9260 6290
rect 9340 6210 9400 6290
rect 9200 6150 9400 6210
rect 9600 6290 9800 6350
rect 9600 6210 9660 6290
rect 9740 6210 9800 6290
rect 9600 6150 9800 6210
rect 2200 6090 2400 6150
rect 2200 6010 2260 6090
rect 2340 6010 2400 6090
rect 2200 5950 2400 6010
rect 2600 6090 2800 6150
rect 2600 6010 2660 6090
rect 2740 6010 2800 6090
rect 2600 5950 2800 6010
rect 3000 6090 3200 6150
rect 3000 6010 3060 6090
rect 3140 6010 3200 6090
rect 3000 5950 3200 6010
rect 3400 6090 3600 6150
rect 3400 6010 3460 6090
rect 3540 6010 3600 6090
rect 3400 5950 3600 6010
rect 3800 6090 4000 6150
rect 3800 6010 3860 6090
rect 3940 6010 4000 6090
rect 3800 5950 4000 6010
rect 4200 6090 4400 6150
rect 4200 6010 4260 6090
rect 4340 6010 4400 6090
rect 4200 5950 4400 6010
rect 4600 6090 4800 6150
rect 4600 6010 4660 6090
rect 4740 6010 4800 6090
rect 4600 5950 4800 6010
rect 5000 6090 5200 6150
rect 5000 6010 5060 6090
rect 5140 6010 5200 6090
rect 5000 5950 5200 6010
rect 5400 6090 5600 6150
rect 5400 6010 5460 6090
rect 5540 6010 5600 6090
rect 5400 5950 5600 6010
rect 5800 6090 6000 6150
rect 5800 6010 5860 6090
rect 5940 6010 6000 6090
rect 5800 5950 6000 6010
rect 6200 6090 6400 6150
rect 6200 6010 6260 6090
rect 6340 6010 6400 6090
rect 6200 5950 6400 6010
rect 6600 6090 6800 6150
rect 6600 6010 6660 6090
rect 6740 6010 6800 6090
rect 6600 5950 6800 6010
rect 7000 6090 7200 6150
rect 7000 6010 7060 6090
rect 7140 6010 7200 6090
rect 7000 5950 7200 6010
rect 7400 6090 7600 6150
rect 7400 6010 7460 6090
rect 7540 6010 7600 6090
rect 7400 5950 7600 6010
rect 7800 6090 8000 6150
rect 7800 6010 7860 6090
rect 7940 6010 8000 6090
rect 7800 5950 8000 6010
rect 8200 6090 8400 6150
rect 8200 6010 8260 6090
rect 8340 6010 8400 6090
rect 8200 5950 8400 6010
rect 8600 6090 8800 6150
rect 8600 6010 8660 6090
rect 8740 6010 8800 6090
rect 8600 5950 8800 6010
rect 9000 6090 9200 6150
rect 9000 6010 9060 6090
rect 9140 6010 9200 6090
rect 9000 5950 9200 6010
rect 9400 6090 9600 6150
rect 9400 6010 9460 6090
rect 9540 6010 9600 6090
rect 9400 5950 9600 6010
rect 9800 6090 10000 6150
rect 9800 6010 9860 6090
rect 9940 6010 10000 6090
rect 9800 5950 10000 6010
rect 2400 5890 2600 5950
rect 2400 5810 2460 5890
rect 2540 5810 2600 5890
rect 2400 5750 2600 5810
rect 2800 5890 3000 5950
rect 2800 5810 2860 5890
rect 2940 5810 3000 5890
rect 2800 5750 3000 5810
rect 3200 5890 3400 5950
rect 3200 5810 3260 5890
rect 3340 5810 3400 5890
rect 3200 5750 3400 5810
rect 3600 5890 3800 5950
rect 3600 5810 3660 5890
rect 3740 5810 3800 5890
rect 3600 5750 3800 5810
rect 4000 5890 4200 5950
rect 4000 5810 4060 5890
rect 4140 5810 4200 5890
rect 4000 5750 4200 5810
rect 4400 5890 4600 5950
rect 4400 5810 4460 5890
rect 4540 5810 4600 5890
rect 4400 5750 4600 5810
rect 4800 5890 5000 5950
rect 4800 5810 4860 5890
rect 4940 5810 5000 5890
rect 4800 5750 5000 5810
rect 5200 5890 5400 5950
rect 5200 5810 5260 5890
rect 5340 5810 5400 5890
rect 5200 5750 5400 5810
rect 5600 5890 5800 5950
rect 5600 5810 5660 5890
rect 5740 5810 5800 5890
rect 5600 5750 5800 5810
rect 6000 5890 6200 5950
rect 6000 5810 6060 5890
rect 6140 5810 6200 5890
rect 6000 5750 6200 5810
rect 6400 5890 6600 5950
rect 6400 5810 6460 5890
rect 6540 5810 6600 5890
rect 6400 5750 6600 5810
rect 6800 5890 7000 5950
rect 6800 5810 6860 5890
rect 6940 5810 7000 5890
rect 6800 5750 7000 5810
rect 7200 5890 7400 5950
rect 7200 5810 7260 5890
rect 7340 5810 7400 5890
rect 7200 5750 7400 5810
rect 7600 5890 7800 5950
rect 7600 5810 7660 5890
rect 7740 5810 7800 5890
rect 7600 5750 7800 5810
rect 8000 5890 8200 5950
rect 8000 5810 8060 5890
rect 8140 5810 8200 5890
rect 8000 5750 8200 5810
rect 8400 5890 8600 5950
rect 8400 5810 8460 5890
rect 8540 5810 8600 5890
rect 8400 5750 8600 5810
rect 8800 5890 9000 5950
rect 8800 5810 8860 5890
rect 8940 5810 9000 5890
rect 8800 5750 9000 5810
rect 9200 5890 9400 5950
rect 9200 5810 9260 5890
rect 9340 5810 9400 5890
rect 9200 5750 9400 5810
rect 9600 5890 9800 5950
rect 9600 5810 9660 5890
rect 9740 5810 9800 5890
rect 9600 5750 9800 5810
rect 2200 5690 2400 5750
rect 2200 5610 2260 5690
rect 2340 5610 2400 5690
rect 2200 5550 2400 5610
rect 2600 5690 2800 5750
rect 2600 5610 2660 5690
rect 2740 5610 2800 5690
rect 2600 5550 2800 5610
rect 3000 5690 3200 5750
rect 3000 5610 3060 5690
rect 3140 5610 3200 5690
rect 3000 5550 3200 5610
rect 3400 5690 3600 5750
rect 3400 5610 3460 5690
rect 3540 5610 3600 5690
rect 3400 5550 3600 5610
rect 3800 5690 4000 5750
rect 3800 5610 3860 5690
rect 3940 5610 4000 5690
rect 3800 5550 4000 5610
rect 4200 5690 4400 5750
rect 4200 5610 4260 5690
rect 4340 5610 4400 5690
rect 4200 5550 4400 5610
rect 4600 5690 4800 5750
rect 4600 5610 4660 5690
rect 4740 5610 4800 5690
rect 4600 5550 4800 5610
rect 5000 5690 5200 5750
rect 5000 5610 5060 5690
rect 5140 5610 5200 5690
rect 5000 5550 5200 5610
rect 5400 5690 5600 5750
rect 5400 5610 5460 5690
rect 5540 5610 5600 5690
rect 5400 5550 5600 5610
rect 5800 5690 6000 5750
rect 5800 5610 5860 5690
rect 5940 5610 6000 5690
rect 5800 5550 6000 5610
rect 6200 5690 6400 5750
rect 6200 5610 6260 5690
rect 6340 5610 6400 5690
rect 6200 5550 6400 5610
rect 6600 5690 6800 5750
rect 6600 5610 6660 5690
rect 6740 5610 6800 5690
rect 6600 5550 6800 5610
rect 7000 5690 7200 5750
rect 7000 5610 7060 5690
rect 7140 5610 7200 5690
rect 7000 5550 7200 5610
rect 7400 5690 7600 5750
rect 7400 5610 7460 5690
rect 7540 5610 7600 5690
rect 7400 5550 7600 5610
rect 7800 5690 8000 5750
rect 7800 5610 7860 5690
rect 7940 5610 8000 5690
rect 7800 5550 8000 5610
rect 8200 5690 8400 5750
rect 8200 5610 8260 5690
rect 8340 5610 8400 5690
rect 8200 5550 8400 5610
rect 8600 5690 8800 5750
rect 8600 5610 8660 5690
rect 8740 5610 8800 5690
rect 8600 5550 8800 5610
rect 9000 5690 9200 5750
rect 9000 5610 9060 5690
rect 9140 5610 9200 5690
rect 9000 5550 9200 5610
rect 9400 5690 9600 5750
rect 9400 5610 9460 5690
rect 9540 5610 9600 5690
rect 9400 5550 9600 5610
rect 9800 5690 10000 5750
rect 9800 5610 9860 5690
rect 9940 5610 10000 5690
rect 9800 5550 10000 5610
rect 2400 5490 2600 5550
rect 2400 5410 2460 5490
rect 2540 5410 2600 5490
rect 2400 5350 2600 5410
rect 2800 5490 3000 5550
rect 2800 5410 2860 5490
rect 2940 5410 3000 5490
rect 2800 5350 3000 5410
rect 3200 5490 3400 5550
rect 3200 5410 3260 5490
rect 3340 5410 3400 5490
rect 3200 5350 3400 5410
rect 3600 5490 3800 5550
rect 3600 5410 3660 5490
rect 3740 5410 3800 5490
rect 3600 5350 3800 5410
rect 4000 5490 4200 5550
rect 4000 5410 4060 5490
rect 4140 5410 4200 5490
rect 4000 5350 4200 5410
rect 4400 5490 4600 5550
rect 4400 5410 4460 5490
rect 4540 5410 4600 5490
rect 4400 5350 4600 5410
rect 4800 5490 5000 5550
rect 4800 5410 4860 5490
rect 4940 5410 5000 5490
rect 4800 5350 5000 5410
rect 5200 5490 5400 5550
rect 5200 5410 5260 5490
rect 5340 5410 5400 5490
rect 5200 5350 5400 5410
rect 5600 5490 5800 5550
rect 5600 5410 5660 5490
rect 5740 5410 5800 5490
rect 5600 5350 5800 5410
rect 6000 5490 6200 5550
rect 6000 5410 6060 5490
rect 6140 5410 6200 5490
rect 6000 5350 6200 5410
rect 6400 5490 6600 5550
rect 6400 5410 6460 5490
rect 6540 5410 6600 5490
rect 6400 5350 6600 5410
rect 6800 5490 7000 5550
rect 6800 5410 6860 5490
rect 6940 5410 7000 5490
rect 6800 5350 7000 5410
rect 7200 5490 7400 5550
rect 7200 5410 7260 5490
rect 7340 5410 7400 5490
rect 7200 5350 7400 5410
rect 7600 5490 7800 5550
rect 7600 5410 7660 5490
rect 7740 5410 7800 5490
rect 7600 5350 7800 5410
rect 8000 5490 8200 5550
rect 8000 5410 8060 5490
rect 8140 5410 8200 5490
rect 8000 5350 8200 5410
rect 8400 5490 8600 5550
rect 8400 5410 8460 5490
rect 8540 5410 8600 5490
rect 8400 5350 8600 5410
rect 8800 5490 9000 5550
rect 8800 5410 8860 5490
rect 8940 5410 9000 5490
rect 8800 5350 9000 5410
rect 9200 5490 9400 5550
rect 9200 5410 9260 5490
rect 9340 5410 9400 5490
rect 9200 5350 9400 5410
rect 9600 5490 9800 5550
rect 9600 5410 9660 5490
rect 9740 5410 9800 5490
rect 9600 5350 9800 5410
rect 2200 5290 2400 5350
rect 2200 5210 2260 5290
rect 2340 5210 2400 5290
rect 2200 5150 2400 5210
rect 2600 5290 2800 5350
rect 2600 5210 2660 5290
rect 2740 5210 2800 5290
rect 2600 5150 2800 5210
rect 3000 5290 3200 5350
rect 3000 5210 3060 5290
rect 3140 5210 3200 5290
rect 3000 5150 3200 5210
rect 3400 5290 3600 5350
rect 3400 5210 3460 5290
rect 3540 5210 3600 5290
rect 3400 5150 3600 5210
rect 3800 5290 4000 5350
rect 3800 5210 3860 5290
rect 3940 5210 4000 5290
rect 3800 5150 4000 5210
rect 4200 5290 4400 5350
rect 4200 5210 4260 5290
rect 4340 5210 4400 5290
rect 4200 5150 4400 5210
rect 4600 5290 4800 5350
rect 4600 5210 4660 5290
rect 4740 5210 4800 5290
rect 4600 5150 4800 5210
rect 5000 5290 5200 5350
rect 5000 5210 5060 5290
rect 5140 5210 5200 5290
rect 5000 5150 5200 5210
rect 5400 5290 5600 5350
rect 5400 5210 5460 5290
rect 5540 5210 5600 5290
rect 5400 5150 5600 5210
rect 5800 5290 6000 5350
rect 5800 5210 5860 5290
rect 5940 5210 6000 5290
rect 5800 5150 6000 5210
rect 6200 5290 6400 5350
rect 6200 5210 6260 5290
rect 6340 5210 6400 5290
rect 6200 5150 6400 5210
rect 6600 5290 6800 5350
rect 6600 5210 6660 5290
rect 6740 5210 6800 5290
rect 6600 5150 6800 5210
rect 7000 5290 7200 5350
rect 7000 5210 7060 5290
rect 7140 5210 7200 5290
rect 7000 5150 7200 5210
rect 7400 5290 7600 5350
rect 7400 5210 7460 5290
rect 7540 5210 7600 5290
rect 7400 5150 7600 5210
rect 7800 5290 8000 5350
rect 7800 5210 7860 5290
rect 7940 5210 8000 5290
rect 7800 5150 8000 5210
rect 8200 5290 8400 5350
rect 8200 5210 8260 5290
rect 8340 5210 8400 5290
rect 8200 5150 8400 5210
rect 8600 5290 8800 5350
rect 8600 5210 8660 5290
rect 8740 5210 8800 5290
rect 8600 5150 8800 5210
rect 9000 5290 9200 5350
rect 9000 5210 9060 5290
rect 9140 5210 9200 5290
rect 9000 5150 9200 5210
rect 9400 5290 9600 5350
rect 9400 5210 9460 5290
rect 9540 5210 9600 5290
rect 9400 5150 9600 5210
rect 9800 5290 10000 5350
rect 9800 5210 9860 5290
rect 9940 5210 10000 5290
rect 9800 5150 10000 5210
rect 2400 5090 2600 5150
rect 2400 5010 2460 5090
rect 2540 5010 2600 5090
rect 2400 4950 2600 5010
rect 2800 5090 3000 5150
rect 2800 5010 2860 5090
rect 2940 5010 3000 5090
rect 2800 4950 3000 5010
rect 3200 5090 3400 5150
rect 3200 5010 3260 5090
rect 3340 5010 3400 5090
rect 3200 4950 3400 5010
rect 3600 5090 3800 5150
rect 3600 5010 3660 5090
rect 3740 5010 3800 5090
rect 3600 4950 3800 5010
rect 4000 5090 4200 5150
rect 4000 5010 4060 5090
rect 4140 5010 4200 5090
rect 4000 4950 4200 5010
rect 4400 5090 4600 5150
rect 4400 5010 4460 5090
rect 4540 5010 4600 5090
rect 4400 4950 4600 5010
rect 4800 5090 5000 5150
rect 4800 5010 4860 5090
rect 4940 5010 5000 5090
rect 4800 4950 5000 5010
rect 5200 5090 5400 5150
rect 5200 5010 5260 5090
rect 5340 5010 5400 5090
rect 5200 4950 5400 5010
rect 5600 5090 5800 5150
rect 5600 5010 5660 5090
rect 5740 5010 5800 5090
rect 5600 4950 5800 5010
rect 6000 5090 6200 5150
rect 6000 5010 6060 5090
rect 6140 5010 6200 5090
rect 6000 4950 6200 5010
rect 6400 5090 6600 5150
rect 6400 5010 6460 5090
rect 6540 5010 6600 5090
rect 6400 4950 6600 5010
rect 6800 5090 7000 5150
rect 6800 5010 6860 5090
rect 6940 5010 7000 5090
rect 6800 4950 7000 5010
rect 7200 5090 7400 5150
rect 7200 5010 7260 5090
rect 7340 5010 7400 5090
rect 7200 4950 7400 5010
rect 7600 5090 7800 5150
rect 7600 5010 7660 5090
rect 7740 5010 7800 5090
rect 7600 4950 7800 5010
rect 8000 5090 8200 5150
rect 8000 5010 8060 5090
rect 8140 5010 8200 5090
rect 8000 4950 8200 5010
rect 8400 5090 8600 5150
rect 8400 5010 8460 5090
rect 8540 5010 8600 5090
rect 8400 4950 8600 5010
rect 8800 5090 9000 5150
rect 8800 5010 8860 5090
rect 8940 5010 9000 5090
rect 8800 4950 9000 5010
rect 9200 5090 9400 5150
rect 9200 5010 9260 5090
rect 9340 5010 9400 5090
rect 9200 4950 9400 5010
rect 9600 5090 9800 5150
rect 9600 5010 9660 5090
rect 9740 5010 9800 5090
rect 9600 4950 9800 5010
rect 2200 4890 2400 4950
rect 2200 4810 2260 4890
rect 2340 4810 2400 4890
rect 2200 4750 2400 4810
rect 2600 4890 2800 4950
rect 2600 4810 2660 4890
rect 2740 4810 2800 4890
rect 2600 4750 2800 4810
rect 3000 4890 3200 4950
rect 3000 4810 3060 4890
rect 3140 4810 3200 4890
rect 3000 4750 3200 4810
rect 3400 4890 3600 4950
rect 3400 4810 3460 4890
rect 3540 4810 3600 4890
rect 3400 4750 3600 4810
rect 3800 4890 4000 4950
rect 3800 4810 3860 4890
rect 3940 4810 4000 4890
rect 3800 4750 4000 4810
rect 4200 4890 4400 4950
rect 4200 4810 4260 4890
rect 4340 4810 4400 4890
rect 4200 4750 4400 4810
rect 4600 4890 4800 4950
rect 4600 4810 4660 4890
rect 4740 4810 4800 4890
rect 4600 4750 4800 4810
rect 5000 4890 5200 4950
rect 5000 4810 5060 4890
rect 5140 4810 5200 4890
rect 5000 4750 5200 4810
rect 5400 4890 5600 4950
rect 5400 4810 5460 4890
rect 5540 4810 5600 4890
rect 5400 4750 5600 4810
rect 5800 4890 6000 4950
rect 5800 4810 5860 4890
rect 5940 4810 6000 4890
rect 5800 4750 6000 4810
rect 6200 4890 6400 4950
rect 6200 4810 6260 4890
rect 6340 4810 6400 4890
rect 6200 4750 6400 4810
rect 6600 4890 6800 4950
rect 6600 4810 6660 4890
rect 6740 4810 6800 4890
rect 6600 4750 6800 4810
rect 7000 4890 7200 4950
rect 7000 4810 7060 4890
rect 7140 4810 7200 4890
rect 7000 4750 7200 4810
rect 7400 4890 7600 4950
rect 7400 4810 7460 4890
rect 7540 4810 7600 4890
rect 7400 4750 7600 4810
rect 7800 4890 8000 4950
rect 7800 4810 7860 4890
rect 7940 4810 8000 4890
rect 7800 4750 8000 4810
rect 8200 4890 8400 4950
rect 8200 4810 8260 4890
rect 8340 4810 8400 4890
rect 8200 4750 8400 4810
rect 8600 4890 8800 4950
rect 8600 4810 8660 4890
rect 8740 4810 8800 4890
rect 8600 4750 8800 4810
rect 9000 4890 9200 4950
rect 9000 4810 9060 4890
rect 9140 4810 9200 4890
rect 9000 4750 9200 4810
rect 9400 4890 9600 4950
rect 9400 4810 9460 4890
rect 9540 4810 9600 4890
rect 9400 4750 9600 4810
rect 9800 4890 10000 4950
rect 9800 4810 9860 4890
rect 9940 4810 10000 4890
rect 9800 4750 10000 4810
rect 2400 4690 2600 4750
rect 2400 4610 2460 4690
rect 2540 4610 2600 4690
rect 2400 4550 2600 4610
rect 2800 4690 3000 4750
rect 2800 4610 2860 4690
rect 2940 4610 3000 4690
rect 2800 4550 3000 4610
rect 3200 4690 3400 4750
rect 3200 4610 3260 4690
rect 3340 4610 3400 4690
rect 3200 4550 3400 4610
rect 3600 4690 3800 4750
rect 3600 4610 3660 4690
rect 3740 4610 3800 4690
rect 3600 4550 3800 4610
rect 4000 4690 4200 4750
rect 4000 4610 4060 4690
rect 4140 4610 4200 4690
rect 4000 4550 4200 4610
rect 4400 4690 4600 4750
rect 4400 4610 4460 4690
rect 4540 4610 4600 4690
rect 4400 4550 4600 4610
rect 4800 4690 5000 4750
rect 4800 4610 4860 4690
rect 4940 4610 5000 4690
rect 4800 4550 5000 4610
rect 5200 4690 5400 4750
rect 5200 4610 5260 4690
rect 5340 4610 5400 4690
rect 5200 4550 5400 4610
rect 5600 4690 5800 4750
rect 5600 4610 5660 4690
rect 5740 4610 5800 4690
rect 5600 4550 5800 4610
rect 6000 4690 6200 4750
rect 6000 4610 6060 4690
rect 6140 4610 6200 4690
rect 6000 4550 6200 4610
rect 6400 4690 6600 4750
rect 6400 4610 6460 4690
rect 6540 4610 6600 4690
rect 6400 4550 6600 4610
rect 6800 4690 7000 4750
rect 6800 4610 6860 4690
rect 6940 4610 7000 4690
rect 6800 4550 7000 4610
rect 7200 4690 7400 4750
rect 7200 4610 7260 4690
rect 7340 4610 7400 4690
rect 7200 4550 7400 4610
rect 7600 4690 7800 4750
rect 7600 4610 7660 4690
rect 7740 4610 7800 4690
rect 7600 4550 7800 4610
rect 8000 4690 8200 4750
rect 8000 4610 8060 4690
rect 8140 4610 8200 4690
rect 8000 4550 8200 4610
rect 8400 4690 8600 4750
rect 8400 4610 8460 4690
rect 8540 4610 8600 4690
rect 8400 4550 8600 4610
rect 8800 4690 9000 4750
rect 8800 4610 8860 4690
rect 8940 4610 9000 4690
rect 8800 4550 9000 4610
rect 9200 4690 9400 4750
rect 9200 4610 9260 4690
rect 9340 4610 9400 4690
rect 9200 4550 9400 4610
rect 9600 4690 9800 4750
rect 9600 4610 9660 4690
rect 9740 4610 9800 4690
rect 9600 4550 9800 4610
rect 2200 4490 2400 4550
rect 2200 4410 2260 4490
rect 2340 4410 2400 4490
rect 2200 4350 2400 4410
rect 2600 4490 2800 4550
rect 2600 4410 2660 4490
rect 2740 4410 2800 4490
rect 2600 4350 2800 4410
rect 3000 4490 3200 4550
rect 3000 4410 3060 4490
rect 3140 4410 3200 4490
rect 3000 4350 3200 4410
rect 3400 4490 3600 4550
rect 3400 4410 3460 4490
rect 3540 4410 3600 4490
rect 3400 4350 3600 4410
rect 3800 4490 4000 4550
rect 3800 4410 3860 4490
rect 3940 4410 4000 4490
rect 3800 4350 4000 4410
rect 4200 4490 4400 4550
rect 4200 4410 4260 4490
rect 4340 4410 4400 4490
rect 4200 4350 4400 4410
rect 4600 4490 4800 4550
rect 4600 4410 4660 4490
rect 4740 4410 4800 4490
rect 4600 4350 4800 4410
rect 5000 4490 5200 4550
rect 5000 4410 5060 4490
rect 5140 4410 5200 4490
rect 5000 4350 5200 4410
rect 5400 4490 5600 4550
rect 5400 4410 5460 4490
rect 5540 4410 5600 4490
rect 5400 4350 5600 4410
rect 5800 4490 6000 4550
rect 5800 4410 5860 4490
rect 5940 4410 6000 4490
rect 5800 4350 6000 4410
rect 6200 4490 6400 4550
rect 6200 4410 6260 4490
rect 6340 4410 6400 4490
rect 6200 4350 6400 4410
rect 6600 4490 6800 4550
rect 6600 4410 6660 4490
rect 6740 4410 6800 4490
rect 6600 4350 6800 4410
rect 7000 4490 7200 4550
rect 7000 4410 7060 4490
rect 7140 4410 7200 4490
rect 7000 4350 7200 4410
rect 7400 4490 7600 4550
rect 7400 4410 7460 4490
rect 7540 4410 7600 4490
rect 7400 4350 7600 4410
rect 7800 4490 8000 4550
rect 7800 4410 7860 4490
rect 7940 4410 8000 4490
rect 7800 4350 8000 4410
rect 8200 4490 8400 4550
rect 8200 4410 8260 4490
rect 8340 4410 8400 4490
rect 8200 4350 8400 4410
rect 8600 4490 8800 4550
rect 8600 4410 8660 4490
rect 8740 4410 8800 4490
rect 8600 4350 8800 4410
rect 9000 4490 9200 4550
rect 9000 4410 9060 4490
rect 9140 4410 9200 4490
rect 9000 4350 9200 4410
rect 9400 4490 9600 4550
rect 9400 4410 9460 4490
rect 9540 4410 9600 4490
rect 9400 4350 9600 4410
rect 9800 4490 10000 4550
rect 9800 4410 9860 4490
rect 9940 4410 10000 4490
rect 9800 4350 10000 4410
rect 2400 4290 2600 4350
rect 2400 4210 2460 4290
rect 2540 4210 2600 4290
rect 2400 4150 2600 4210
rect 2800 4290 3000 4350
rect 2800 4210 2860 4290
rect 2940 4210 3000 4290
rect 2800 4150 3000 4210
rect 3200 4290 3400 4350
rect 3200 4210 3260 4290
rect 3340 4210 3400 4290
rect 3200 4150 3400 4210
rect 3600 4290 3800 4350
rect 3600 4210 3660 4290
rect 3740 4210 3800 4290
rect 3600 4150 3800 4210
rect 4000 4290 4200 4350
rect 4000 4210 4060 4290
rect 4140 4210 4200 4290
rect 4000 4150 4200 4210
rect 4400 4290 4600 4350
rect 4400 4210 4460 4290
rect 4540 4210 4600 4290
rect 4400 4150 4600 4210
rect 4800 4290 5000 4350
rect 4800 4210 4860 4290
rect 4940 4210 5000 4290
rect 4800 4150 5000 4210
rect 5200 4290 5400 4350
rect 5200 4210 5260 4290
rect 5340 4210 5400 4290
rect 5200 4150 5400 4210
rect 5600 4290 5800 4350
rect 5600 4210 5660 4290
rect 5740 4210 5800 4290
rect 5600 4150 5800 4210
rect 6000 4290 6200 4350
rect 6000 4210 6060 4290
rect 6140 4210 6200 4290
rect 6000 4150 6200 4210
rect 6400 4290 6600 4350
rect 6400 4210 6460 4290
rect 6540 4210 6600 4290
rect 6400 4150 6600 4210
rect 6800 4290 7000 4350
rect 6800 4210 6860 4290
rect 6940 4210 7000 4290
rect 6800 4150 7000 4210
rect 7200 4290 7400 4350
rect 7200 4210 7260 4290
rect 7340 4210 7400 4290
rect 7200 4150 7400 4210
rect 7600 4290 7800 4350
rect 7600 4210 7660 4290
rect 7740 4210 7800 4290
rect 7600 4150 7800 4210
rect 8000 4290 8200 4350
rect 8000 4210 8060 4290
rect 8140 4210 8200 4290
rect 8000 4150 8200 4210
rect 8400 4290 8600 4350
rect 8400 4210 8460 4290
rect 8540 4210 8600 4290
rect 8400 4150 8600 4210
rect 8800 4290 9000 4350
rect 8800 4210 8860 4290
rect 8940 4210 9000 4290
rect 8800 4150 9000 4210
rect 9200 4290 9400 4350
rect 9200 4210 9260 4290
rect 9340 4210 9400 4290
rect 9200 4150 9400 4210
rect 9600 4290 9800 4350
rect 9600 4210 9660 4290
rect 9740 4210 9800 4290
rect 9600 4150 9800 4210
rect 2200 4090 2400 4150
rect 2200 4010 2260 4090
rect 2340 4010 2400 4090
rect 2200 3950 2400 4010
rect 2600 4090 2800 4150
rect 2600 4010 2660 4090
rect 2740 4010 2800 4090
rect 2600 3950 2800 4010
rect 3000 4090 3200 4150
rect 3000 4010 3060 4090
rect 3140 4010 3200 4090
rect 3000 3950 3200 4010
rect 3400 4090 3600 4150
rect 3400 4010 3460 4090
rect 3540 4010 3600 4090
rect 3400 3950 3600 4010
rect 3800 4090 4000 4150
rect 3800 4010 3860 4090
rect 3940 4010 4000 4090
rect 3800 3950 4000 4010
rect 4200 4090 4400 4150
rect 4200 4010 4260 4090
rect 4340 4010 4400 4090
rect 4200 3950 4400 4010
rect 4600 4090 4800 4150
rect 4600 4010 4660 4090
rect 4740 4010 4800 4090
rect 4600 3950 4800 4010
rect 5000 4090 5200 4150
rect 5000 4010 5060 4090
rect 5140 4010 5200 4090
rect 5000 3950 5200 4010
rect 5400 4090 5600 4150
rect 5400 4010 5460 4090
rect 5540 4010 5600 4090
rect 5400 3950 5600 4010
rect 5800 4090 6000 4150
rect 5800 4010 5860 4090
rect 5940 4010 6000 4090
rect 5800 3950 6000 4010
rect 6200 4090 6400 4150
rect 6200 4010 6260 4090
rect 6340 4010 6400 4090
rect 6200 3950 6400 4010
rect 6600 4090 6800 4150
rect 6600 4010 6660 4090
rect 6740 4010 6800 4090
rect 6600 3950 6800 4010
rect 7000 4090 7200 4150
rect 7000 4010 7060 4090
rect 7140 4010 7200 4090
rect 7000 3950 7200 4010
rect 7400 4090 7600 4150
rect 7400 4010 7460 4090
rect 7540 4010 7600 4090
rect 7400 3950 7600 4010
rect 7800 4090 8000 4150
rect 7800 4010 7860 4090
rect 7940 4010 8000 4090
rect 7800 3950 8000 4010
rect 8200 4090 8400 4150
rect 8200 4010 8260 4090
rect 8340 4010 8400 4090
rect 8200 3950 8400 4010
rect 8600 4090 8800 4150
rect 8600 4010 8660 4090
rect 8740 4010 8800 4090
rect 8600 3950 8800 4010
rect 9000 4090 9200 4150
rect 9000 4010 9060 4090
rect 9140 4010 9200 4090
rect 9000 3950 9200 4010
rect 9400 4090 9600 4150
rect 9400 4010 9460 4090
rect 9540 4010 9600 4090
rect 9400 3950 9600 4010
rect 9800 4090 10000 4150
rect 9800 4010 9860 4090
rect 9940 4010 10000 4090
rect 9800 3950 10000 4010
rect 2400 3890 2600 3950
rect 2400 3810 2460 3890
rect 2540 3810 2600 3890
rect 2400 3750 2600 3810
rect 2800 3890 3000 3950
rect 2800 3810 2860 3890
rect 2940 3810 3000 3890
rect 2800 3750 3000 3810
rect 3200 3890 3400 3950
rect 3200 3810 3260 3890
rect 3340 3810 3400 3890
rect 3200 3750 3400 3810
rect 3600 3890 3800 3950
rect 3600 3810 3660 3890
rect 3740 3810 3800 3890
rect 3600 3750 3800 3810
rect 4000 3890 4200 3950
rect 4000 3810 4060 3890
rect 4140 3810 4200 3890
rect 4000 3750 4200 3810
rect 4400 3890 4600 3950
rect 4400 3810 4460 3890
rect 4540 3810 4600 3890
rect 4400 3750 4600 3810
rect 4800 3890 5000 3950
rect 4800 3810 4860 3890
rect 4940 3810 5000 3890
rect 4800 3750 5000 3810
rect 5200 3890 5400 3950
rect 5200 3810 5260 3890
rect 5340 3810 5400 3890
rect 5200 3750 5400 3810
rect 5600 3890 5800 3950
rect 5600 3810 5660 3890
rect 5740 3810 5800 3890
rect 5600 3750 5800 3810
rect 6000 3890 6200 3950
rect 6000 3810 6060 3890
rect 6140 3810 6200 3890
rect 6000 3750 6200 3810
rect 6400 3890 6600 3950
rect 6400 3810 6460 3890
rect 6540 3810 6600 3890
rect 6400 3750 6600 3810
rect 6800 3890 7000 3950
rect 6800 3810 6860 3890
rect 6940 3810 7000 3890
rect 6800 3750 7000 3810
rect 7200 3890 7400 3950
rect 7200 3810 7260 3890
rect 7340 3810 7400 3890
rect 7200 3750 7400 3810
rect 7600 3890 7800 3950
rect 7600 3810 7660 3890
rect 7740 3810 7800 3890
rect 7600 3750 7800 3810
rect 8000 3890 8200 3950
rect 8000 3810 8060 3890
rect 8140 3810 8200 3890
rect 8000 3750 8200 3810
rect 8400 3890 8600 3950
rect 8400 3810 8460 3890
rect 8540 3810 8600 3890
rect 8400 3750 8600 3810
rect 8800 3890 9000 3950
rect 8800 3810 8860 3890
rect 8940 3810 9000 3890
rect 8800 3750 9000 3810
rect 9200 3890 9400 3950
rect 9200 3810 9260 3890
rect 9340 3810 9400 3890
rect 9200 3750 9400 3810
rect 9600 3890 9800 3950
rect 9600 3810 9660 3890
rect 9740 3810 9800 3890
rect 9600 3750 9800 3810
rect 2200 3690 2400 3750
rect 2200 3610 2260 3690
rect 2340 3610 2400 3690
rect 2200 3550 2400 3610
rect 2600 3690 2800 3750
rect 2600 3610 2660 3690
rect 2740 3610 2800 3690
rect 2600 3550 2800 3610
rect 3000 3690 3200 3750
rect 3000 3610 3060 3690
rect 3140 3610 3200 3690
rect 3000 3550 3200 3610
rect 3400 3690 3600 3750
rect 3400 3610 3460 3690
rect 3540 3610 3600 3690
rect 3400 3550 3600 3610
rect 3800 3690 4000 3750
rect 3800 3610 3860 3690
rect 3940 3610 4000 3690
rect 3800 3550 4000 3610
rect 4200 3690 4400 3750
rect 4200 3610 4260 3690
rect 4340 3610 4400 3690
rect 4200 3550 4400 3610
rect 4600 3690 4800 3750
rect 4600 3610 4660 3690
rect 4740 3610 4800 3690
rect 4600 3550 4800 3610
rect 5000 3690 5200 3750
rect 5000 3610 5060 3690
rect 5140 3610 5200 3690
rect 5000 3550 5200 3610
rect 5400 3690 5600 3750
rect 5400 3610 5460 3690
rect 5540 3610 5600 3690
rect 5400 3550 5600 3610
rect 5800 3690 6000 3750
rect 5800 3610 5860 3690
rect 5940 3610 6000 3690
rect 5800 3550 6000 3610
rect 6200 3690 6400 3750
rect 6200 3610 6260 3690
rect 6340 3610 6400 3690
rect 6200 3550 6400 3610
rect 6600 3690 6800 3750
rect 6600 3610 6660 3690
rect 6740 3610 6800 3690
rect 6600 3550 6800 3610
rect 7000 3690 7200 3750
rect 7000 3610 7060 3690
rect 7140 3610 7200 3690
rect 7000 3550 7200 3610
rect 7400 3690 7600 3750
rect 7400 3610 7460 3690
rect 7540 3610 7600 3690
rect 7400 3550 7600 3610
rect 7800 3690 8000 3750
rect 7800 3610 7860 3690
rect 7940 3610 8000 3690
rect 7800 3550 8000 3610
rect 8200 3690 8400 3750
rect 8200 3610 8260 3690
rect 8340 3610 8400 3690
rect 8200 3550 8400 3610
rect 8600 3690 8800 3750
rect 8600 3610 8660 3690
rect 8740 3610 8800 3690
rect 8600 3550 8800 3610
rect 9000 3690 9200 3750
rect 9000 3610 9060 3690
rect 9140 3610 9200 3690
rect 9000 3550 9200 3610
rect 9400 3690 9600 3750
rect 9400 3610 9460 3690
rect 9540 3610 9600 3690
rect 9400 3550 9600 3610
rect 9800 3690 10000 3750
rect 9800 3610 9860 3690
rect 9940 3610 10000 3690
rect 9800 3550 10000 3610
rect 2400 3490 2600 3550
rect 2400 3410 2460 3490
rect 2540 3410 2600 3490
rect 2400 3350 2600 3410
rect 2800 3490 3000 3550
rect 2800 3410 2860 3490
rect 2940 3410 3000 3490
rect 2800 3350 3000 3410
rect 3200 3490 3400 3550
rect 3200 3410 3260 3490
rect 3340 3410 3400 3490
rect 3200 3350 3400 3410
rect 3600 3490 3800 3550
rect 3600 3410 3660 3490
rect 3740 3410 3800 3490
rect 3600 3350 3800 3410
rect 4000 3490 4200 3550
rect 4000 3410 4060 3490
rect 4140 3410 4200 3490
rect 4000 3350 4200 3410
rect 4400 3490 4600 3550
rect 4400 3410 4460 3490
rect 4540 3410 4600 3490
rect 4400 3350 4600 3410
rect 4800 3490 5000 3550
rect 4800 3410 4860 3490
rect 4940 3410 5000 3490
rect 4800 3350 5000 3410
rect 5200 3490 5400 3550
rect 5200 3410 5260 3490
rect 5340 3410 5400 3490
rect 5200 3350 5400 3410
rect 5600 3490 5800 3550
rect 5600 3410 5660 3490
rect 5740 3410 5800 3490
rect 5600 3350 5800 3410
rect 6000 3490 6200 3550
rect 6000 3410 6060 3490
rect 6140 3410 6200 3490
rect 6000 3350 6200 3410
rect 6400 3490 6600 3550
rect 6400 3410 6460 3490
rect 6540 3410 6600 3490
rect 6400 3350 6600 3410
rect 6800 3490 7000 3550
rect 6800 3410 6860 3490
rect 6940 3410 7000 3490
rect 6800 3350 7000 3410
rect 7200 3490 7400 3550
rect 7200 3410 7260 3490
rect 7340 3410 7400 3490
rect 7200 3350 7400 3410
rect 7600 3490 7800 3550
rect 7600 3410 7660 3490
rect 7740 3410 7800 3490
rect 7600 3350 7800 3410
rect 8000 3490 8200 3550
rect 8000 3410 8060 3490
rect 8140 3410 8200 3490
rect 8000 3350 8200 3410
rect 8400 3490 8600 3550
rect 8400 3410 8460 3490
rect 8540 3410 8600 3490
rect 8400 3350 8600 3410
rect 8800 3490 9000 3550
rect 8800 3410 8860 3490
rect 8940 3410 9000 3490
rect 8800 3350 9000 3410
rect 9200 3490 9400 3550
rect 9200 3410 9260 3490
rect 9340 3410 9400 3490
rect 9200 3350 9400 3410
rect 9600 3490 9800 3550
rect 9600 3410 9660 3490
rect 9740 3410 9800 3490
rect 9600 3350 9800 3410
rect 2200 3290 2400 3350
rect 2200 3210 2260 3290
rect 2340 3210 2400 3290
rect 2200 3150 2400 3210
rect 2600 3290 2800 3350
rect 2600 3210 2660 3290
rect 2740 3210 2800 3290
rect 2600 3150 2800 3210
rect 3000 3290 3200 3350
rect 3000 3210 3060 3290
rect 3140 3210 3200 3290
rect 3000 3150 3200 3210
rect 3400 3290 3600 3350
rect 3400 3210 3460 3290
rect 3540 3210 3600 3290
rect 3400 3150 3600 3210
rect 3800 3290 4000 3350
rect 3800 3210 3860 3290
rect 3940 3210 4000 3290
rect 3800 3150 4000 3210
rect 4200 3290 4400 3350
rect 4200 3210 4260 3290
rect 4340 3210 4400 3290
rect 4200 3150 4400 3210
rect 4600 3290 4800 3350
rect 4600 3210 4660 3290
rect 4740 3210 4800 3290
rect 4600 3150 4800 3210
rect 5000 3290 5200 3350
rect 5000 3210 5060 3290
rect 5140 3210 5200 3290
rect 5000 3150 5200 3210
rect 5400 3290 5600 3350
rect 5400 3210 5460 3290
rect 5540 3210 5600 3290
rect 5400 3150 5600 3210
rect 5800 3290 6000 3350
rect 5800 3210 5860 3290
rect 5940 3210 6000 3290
rect 5800 3150 6000 3210
rect 6200 3290 6400 3350
rect 6200 3210 6260 3290
rect 6340 3210 6400 3290
rect 6200 3150 6400 3210
rect 6600 3290 6800 3350
rect 6600 3210 6660 3290
rect 6740 3210 6800 3290
rect 6600 3150 6800 3210
rect 7000 3290 7200 3350
rect 7000 3210 7060 3290
rect 7140 3210 7200 3290
rect 7000 3150 7200 3210
rect 7400 3290 7600 3350
rect 7400 3210 7460 3290
rect 7540 3210 7600 3290
rect 7400 3150 7600 3210
rect 7800 3290 8000 3350
rect 7800 3210 7860 3290
rect 7940 3210 8000 3290
rect 7800 3150 8000 3210
rect 8200 3290 8400 3350
rect 8200 3210 8260 3290
rect 8340 3210 8400 3290
rect 8200 3150 8400 3210
rect 8600 3290 8800 3350
rect 8600 3210 8660 3290
rect 8740 3210 8800 3290
rect 8600 3150 8800 3210
rect 9000 3290 9200 3350
rect 9000 3210 9060 3290
rect 9140 3210 9200 3290
rect 9000 3150 9200 3210
rect 9400 3290 9600 3350
rect 9400 3210 9460 3290
rect 9540 3210 9600 3290
rect 9400 3150 9600 3210
rect 9800 3290 10000 3350
rect 9800 3210 9860 3290
rect 9940 3210 10000 3290
rect 9800 3150 10000 3210
rect 2400 3090 2600 3150
rect 2400 3010 2460 3090
rect 2540 3010 2600 3090
rect 2400 2950 2600 3010
rect 2800 3090 3000 3150
rect 2800 3010 2860 3090
rect 2940 3010 3000 3090
rect 2800 2950 3000 3010
rect 3200 3090 3400 3150
rect 3200 3010 3260 3090
rect 3340 3010 3400 3090
rect 3200 2950 3400 3010
rect 3600 3090 3800 3150
rect 3600 3010 3660 3090
rect 3740 3010 3800 3090
rect 3600 2950 3800 3010
rect 4000 3090 4200 3150
rect 4000 3010 4060 3090
rect 4140 3010 4200 3090
rect 4000 2950 4200 3010
rect 4400 3090 4600 3150
rect 4400 3010 4460 3090
rect 4540 3010 4600 3090
rect 4400 2950 4600 3010
rect 4800 3090 5000 3150
rect 4800 3010 4860 3090
rect 4940 3010 5000 3090
rect 4800 2950 5000 3010
rect 5200 3090 5400 3150
rect 5200 3010 5260 3090
rect 5340 3010 5400 3090
rect 5200 2950 5400 3010
rect 5600 3090 5800 3150
rect 5600 3010 5660 3090
rect 5740 3010 5800 3090
rect 5600 2950 5800 3010
rect 6000 3090 6200 3150
rect 6000 3010 6060 3090
rect 6140 3010 6200 3090
rect 6000 2950 6200 3010
rect 6400 3090 6600 3150
rect 6400 3010 6460 3090
rect 6540 3010 6600 3090
rect 6400 2950 6600 3010
rect 6800 3090 7000 3150
rect 6800 3010 6860 3090
rect 6940 3010 7000 3090
rect 6800 2950 7000 3010
rect 7200 3090 7400 3150
rect 7200 3010 7260 3090
rect 7340 3010 7400 3090
rect 7200 2950 7400 3010
rect 7600 3090 7800 3150
rect 7600 3010 7660 3090
rect 7740 3010 7800 3090
rect 7600 2950 7800 3010
rect 8000 3090 8200 3150
rect 8000 3010 8060 3090
rect 8140 3010 8200 3090
rect 8000 2950 8200 3010
rect 8400 3090 8600 3150
rect 8400 3010 8460 3090
rect 8540 3010 8600 3090
rect 8400 2950 8600 3010
rect 8800 3090 9000 3150
rect 8800 3010 8860 3090
rect 8940 3010 9000 3090
rect 8800 2950 9000 3010
rect 9200 3090 9400 3150
rect 9200 3010 9260 3090
rect 9340 3010 9400 3090
rect 9200 2950 9400 3010
rect 9600 3090 9800 3150
rect 9600 3010 9660 3090
rect 9740 3010 9800 3090
rect 9600 2950 9800 3010
rect 2200 2890 2400 2950
rect 2200 2810 2260 2890
rect 2340 2810 2400 2890
rect 2200 2750 2400 2810
rect 2600 2890 2800 2950
rect 2600 2810 2660 2890
rect 2740 2810 2800 2890
rect 2600 2750 2800 2810
rect 3000 2890 3200 2950
rect 3000 2810 3060 2890
rect 3140 2810 3200 2890
rect 3000 2750 3200 2810
rect 3400 2890 3600 2950
rect 3400 2810 3460 2890
rect 3540 2810 3600 2890
rect 3400 2750 3600 2810
rect 3800 2890 4000 2950
rect 3800 2810 3860 2890
rect 3940 2810 4000 2890
rect 3800 2750 4000 2810
rect 4200 2890 4400 2950
rect 4200 2810 4260 2890
rect 4340 2810 4400 2890
rect 4200 2750 4400 2810
rect 4600 2890 4800 2950
rect 4600 2810 4660 2890
rect 4740 2810 4800 2890
rect 4600 2750 4800 2810
rect 5000 2890 5200 2950
rect 5000 2810 5060 2890
rect 5140 2810 5200 2890
rect 5000 2750 5200 2810
rect 5400 2890 5600 2950
rect 5400 2810 5460 2890
rect 5540 2810 5600 2890
rect 5400 2750 5600 2810
rect 5800 2890 6000 2950
rect 5800 2810 5860 2890
rect 5940 2810 6000 2890
rect 5800 2750 6000 2810
rect 6200 2890 6400 2950
rect 6200 2810 6260 2890
rect 6340 2810 6400 2890
rect 6200 2750 6400 2810
rect 6600 2890 6800 2950
rect 6600 2810 6660 2890
rect 6740 2810 6800 2890
rect 6600 2750 6800 2810
rect 7000 2890 7200 2950
rect 7000 2810 7060 2890
rect 7140 2810 7200 2890
rect 7000 2750 7200 2810
rect 7400 2890 7600 2950
rect 7400 2810 7460 2890
rect 7540 2810 7600 2890
rect 7400 2750 7600 2810
rect 7800 2890 8000 2950
rect 7800 2810 7860 2890
rect 7940 2810 8000 2890
rect 7800 2750 8000 2810
rect 8200 2890 8400 2950
rect 8200 2810 8260 2890
rect 8340 2810 8400 2890
rect 8200 2750 8400 2810
rect 8600 2890 8800 2950
rect 8600 2810 8660 2890
rect 8740 2810 8800 2890
rect 8600 2750 8800 2810
rect 9000 2890 9200 2950
rect 9000 2810 9060 2890
rect 9140 2810 9200 2890
rect 9000 2750 9200 2810
rect 9400 2890 9600 2950
rect 9400 2810 9460 2890
rect 9540 2810 9600 2890
rect 9400 2750 9600 2810
rect 9800 2890 10000 2950
rect 9800 2810 9860 2890
rect 9940 2810 10000 2890
rect 9800 2750 10000 2810
rect 2400 2690 2600 2750
rect 2400 2610 2460 2690
rect 2540 2610 2600 2690
rect 2400 2550 2600 2610
rect 2800 2690 3000 2750
rect 2800 2610 2860 2690
rect 2940 2610 3000 2690
rect 2800 2550 3000 2610
rect 3200 2690 3400 2750
rect 3200 2610 3260 2690
rect 3340 2610 3400 2690
rect 3200 2550 3400 2610
rect 3600 2690 3800 2750
rect 3600 2610 3660 2690
rect 3740 2610 3800 2690
rect 3600 2550 3800 2610
rect 4000 2690 4200 2750
rect 4000 2610 4060 2690
rect 4140 2610 4200 2690
rect 4000 2550 4200 2610
rect 4400 2690 4600 2750
rect 4400 2610 4460 2690
rect 4540 2610 4600 2690
rect 4400 2550 4600 2610
rect 4800 2690 5000 2750
rect 4800 2610 4860 2690
rect 4940 2610 5000 2690
rect 4800 2550 5000 2610
rect 5200 2690 5400 2750
rect 5200 2610 5260 2690
rect 5340 2610 5400 2690
rect 5200 2550 5400 2610
rect 5600 2690 5800 2750
rect 5600 2610 5660 2690
rect 5740 2610 5800 2690
rect 5600 2550 5800 2610
rect 6000 2690 6200 2750
rect 6000 2610 6060 2690
rect 6140 2610 6200 2690
rect 6000 2550 6200 2610
rect 6400 2690 6600 2750
rect 6400 2610 6460 2690
rect 6540 2610 6600 2690
rect 6400 2550 6600 2610
rect 6800 2690 7000 2750
rect 6800 2610 6860 2690
rect 6940 2610 7000 2690
rect 6800 2550 7000 2610
rect 7200 2690 7400 2750
rect 7200 2610 7260 2690
rect 7340 2610 7400 2690
rect 7200 2550 7400 2610
rect 7600 2690 7800 2750
rect 7600 2610 7660 2690
rect 7740 2610 7800 2690
rect 7600 2550 7800 2610
rect 8000 2690 8200 2750
rect 8000 2610 8060 2690
rect 8140 2610 8200 2690
rect 8000 2550 8200 2610
rect 8400 2690 8600 2750
rect 8400 2610 8460 2690
rect 8540 2610 8600 2690
rect 8400 2550 8600 2610
rect 8800 2690 9000 2750
rect 8800 2610 8860 2690
rect 8940 2610 9000 2690
rect 8800 2550 9000 2610
rect 9200 2690 9400 2750
rect 9200 2610 9260 2690
rect 9340 2610 9400 2690
rect 9200 2550 9400 2610
rect 9600 2690 9800 2750
rect 9600 2610 9660 2690
rect 9740 2610 9800 2690
rect 9600 2550 9800 2610
rect 2200 2490 2400 2550
rect 2200 2410 2260 2490
rect 2340 2410 2400 2490
rect 2200 2350 2400 2410
rect 2600 2490 2800 2550
rect 2600 2410 2660 2490
rect 2740 2410 2800 2490
rect 2600 2350 2800 2410
rect 3000 2490 3200 2550
rect 3000 2410 3060 2490
rect 3140 2410 3200 2490
rect 3000 2350 3200 2410
rect 3400 2490 3600 2550
rect 3400 2410 3460 2490
rect 3540 2410 3600 2490
rect 3400 2350 3600 2410
rect 3800 2490 4000 2550
rect 3800 2410 3860 2490
rect 3940 2410 4000 2490
rect 3800 2350 4000 2410
rect 4200 2490 4400 2550
rect 4200 2410 4260 2490
rect 4340 2410 4400 2490
rect 4200 2350 4400 2410
rect 4600 2490 4800 2550
rect 4600 2410 4660 2490
rect 4740 2410 4800 2490
rect 4600 2350 4800 2410
rect 5000 2490 5200 2550
rect 5000 2410 5060 2490
rect 5140 2410 5200 2490
rect 5000 2350 5200 2410
rect 5400 2490 5600 2550
rect 5400 2410 5460 2490
rect 5540 2410 5600 2490
rect 5400 2350 5600 2410
rect 5800 2490 6000 2550
rect 5800 2410 5860 2490
rect 5940 2410 6000 2490
rect 5800 2350 6000 2410
rect 6200 2490 6400 2550
rect 6200 2410 6260 2490
rect 6340 2410 6400 2490
rect 6200 2350 6400 2410
rect 6600 2490 6800 2550
rect 6600 2410 6660 2490
rect 6740 2410 6800 2490
rect 6600 2350 6800 2410
rect 7000 2490 7200 2550
rect 7000 2410 7060 2490
rect 7140 2410 7200 2490
rect 7000 2350 7200 2410
rect 7400 2490 7600 2550
rect 7400 2410 7460 2490
rect 7540 2410 7600 2490
rect 7400 2350 7600 2410
rect 7800 2490 8000 2550
rect 7800 2410 7860 2490
rect 7940 2410 8000 2490
rect 7800 2350 8000 2410
rect 8200 2490 8400 2550
rect 8200 2410 8260 2490
rect 8340 2410 8400 2490
rect 8200 2350 8400 2410
rect 8600 2490 8800 2550
rect 8600 2410 8660 2490
rect 8740 2410 8800 2490
rect 8600 2350 8800 2410
rect 9000 2490 9200 2550
rect 9000 2410 9060 2490
rect 9140 2410 9200 2490
rect 9000 2350 9200 2410
rect 9400 2490 9600 2550
rect 9400 2410 9460 2490
rect 9540 2410 9600 2490
rect 9400 2350 9600 2410
rect 9800 2490 10000 2550
rect 9800 2410 9860 2490
rect 9940 2410 10000 2490
rect 9800 2350 10000 2410
rect 2400 2290 2600 2350
rect 2400 2210 2460 2290
rect 2540 2210 2600 2290
rect 2400 2150 2600 2210
rect 2800 2290 3000 2350
rect 2800 2210 2860 2290
rect 2940 2210 3000 2290
rect 2800 2150 3000 2210
rect 3200 2290 3400 2350
rect 3200 2210 3260 2290
rect 3340 2210 3400 2290
rect 3200 2150 3400 2210
rect 3600 2290 3800 2350
rect 3600 2210 3660 2290
rect 3740 2210 3800 2290
rect 3600 2150 3800 2210
rect 4000 2290 4200 2350
rect 4000 2210 4060 2290
rect 4140 2210 4200 2290
rect 4000 2150 4200 2210
rect 4400 2290 4600 2350
rect 4400 2210 4460 2290
rect 4540 2210 4600 2290
rect 4400 2150 4600 2210
rect 4800 2290 5000 2350
rect 4800 2210 4860 2290
rect 4940 2210 5000 2290
rect 4800 2150 5000 2210
rect 5200 2290 5400 2350
rect 5200 2210 5260 2290
rect 5340 2210 5400 2290
rect 5200 2150 5400 2210
rect 5600 2290 5800 2350
rect 5600 2210 5660 2290
rect 5740 2210 5800 2290
rect 5600 2150 5800 2210
rect 6000 2290 6200 2350
rect 6000 2210 6060 2290
rect 6140 2210 6200 2290
rect 6000 2150 6200 2210
rect 6400 2290 6600 2350
rect 6400 2210 6460 2290
rect 6540 2210 6600 2290
rect 6400 2150 6600 2210
rect 6800 2290 7000 2350
rect 6800 2210 6860 2290
rect 6940 2210 7000 2290
rect 6800 2150 7000 2210
rect 7200 2290 7400 2350
rect 7200 2210 7260 2290
rect 7340 2210 7400 2290
rect 7200 2150 7400 2210
rect 7600 2290 7800 2350
rect 7600 2210 7660 2290
rect 7740 2210 7800 2290
rect 7600 2150 7800 2210
rect 8000 2290 8200 2350
rect 8000 2210 8060 2290
rect 8140 2210 8200 2290
rect 8000 2150 8200 2210
rect 8400 2290 8600 2350
rect 8400 2210 8460 2290
rect 8540 2210 8600 2290
rect 8400 2150 8600 2210
rect 8800 2290 9000 2350
rect 8800 2210 8860 2290
rect 8940 2210 9000 2290
rect 8800 2150 9000 2210
rect 9200 2290 9400 2350
rect 9200 2210 9260 2290
rect 9340 2210 9400 2290
rect 9200 2150 9400 2210
rect 9600 2290 9800 2350
rect 9600 2210 9660 2290
rect 9740 2210 9800 2290
rect 9600 2150 9800 2210
rect 2200 2090 2400 2150
rect 2200 2010 2260 2090
rect 2340 2010 2400 2090
rect 2200 1950 2400 2010
rect 2600 2090 2800 2150
rect 2600 2010 2660 2090
rect 2740 2010 2800 2090
rect 2600 1950 2800 2010
rect 3000 2090 3200 2150
rect 3000 2010 3060 2090
rect 3140 2010 3200 2090
rect 3000 1950 3200 2010
rect 3400 2090 3600 2150
rect 3400 2010 3460 2090
rect 3540 2010 3600 2090
rect 3400 1950 3600 2010
rect 3800 2090 4000 2150
rect 3800 2010 3860 2090
rect 3940 2010 4000 2090
rect 3800 1950 4000 2010
rect 4200 2090 4400 2150
rect 4200 2010 4260 2090
rect 4340 2010 4400 2090
rect 4200 1950 4400 2010
rect 4600 2090 4800 2150
rect 4600 2010 4660 2090
rect 4740 2010 4800 2090
rect 4600 1950 4800 2010
rect 5000 2090 5200 2150
rect 5000 2010 5060 2090
rect 5140 2010 5200 2090
rect 5000 1950 5200 2010
rect 5400 2090 5600 2150
rect 5400 2010 5460 2090
rect 5540 2010 5600 2090
rect 5400 1950 5600 2010
rect 5800 2090 6000 2150
rect 5800 2010 5860 2090
rect 5940 2010 6000 2090
rect 5800 1950 6000 2010
rect 6200 2090 6400 2150
rect 6200 2010 6260 2090
rect 6340 2010 6400 2090
rect 6200 1950 6400 2010
rect 6600 2090 6800 2150
rect 6600 2010 6660 2090
rect 6740 2010 6800 2090
rect 6600 1950 6800 2010
rect 7000 2090 7200 2150
rect 7000 2010 7060 2090
rect 7140 2010 7200 2090
rect 7000 1950 7200 2010
rect 7400 2090 7600 2150
rect 7400 2010 7460 2090
rect 7540 2010 7600 2090
rect 7400 1950 7600 2010
rect 7800 2090 8000 2150
rect 7800 2010 7860 2090
rect 7940 2010 8000 2090
rect 7800 1950 8000 2010
rect 8200 2090 8400 2150
rect 8200 2010 8260 2090
rect 8340 2010 8400 2090
rect 8200 1950 8400 2010
rect 8600 2090 8800 2150
rect 8600 2010 8660 2090
rect 8740 2010 8800 2090
rect 8600 1950 8800 2010
rect 9000 2090 9200 2150
rect 9000 2010 9060 2090
rect 9140 2010 9200 2090
rect 9000 1950 9200 2010
rect 9400 2090 9600 2150
rect 9400 2010 9460 2090
rect 9540 2010 9600 2090
rect 9400 1950 9600 2010
rect 9800 2090 10000 2150
rect 9800 2010 9860 2090
rect 9940 2010 10000 2090
rect 9800 1950 10000 2010
rect 2400 1890 2600 1950
rect 2400 1810 2460 1890
rect 2540 1810 2600 1890
rect 2400 1750 2600 1810
rect 2800 1890 3000 1950
rect 2800 1810 2860 1890
rect 2940 1810 3000 1890
rect 2800 1750 3000 1810
rect 3200 1890 3400 1950
rect 3200 1810 3260 1890
rect 3340 1810 3400 1890
rect 3200 1750 3400 1810
rect 3600 1890 3800 1950
rect 3600 1810 3660 1890
rect 3740 1810 3800 1890
rect 3600 1750 3800 1810
rect 4000 1890 4200 1950
rect 4000 1810 4060 1890
rect 4140 1810 4200 1890
rect 4000 1750 4200 1810
rect 4400 1890 4600 1950
rect 4400 1810 4460 1890
rect 4540 1810 4600 1890
rect 4400 1750 4600 1810
rect 4800 1890 5000 1950
rect 4800 1810 4860 1890
rect 4940 1810 5000 1890
rect 4800 1750 5000 1810
rect 5200 1890 5400 1950
rect 5200 1810 5260 1890
rect 5340 1810 5400 1890
rect 5200 1750 5400 1810
rect 5600 1890 5800 1950
rect 5600 1810 5660 1890
rect 5740 1810 5800 1890
rect 5600 1750 5800 1810
rect 6000 1890 6200 1950
rect 6000 1810 6060 1890
rect 6140 1810 6200 1890
rect 6000 1750 6200 1810
rect 6400 1890 6600 1950
rect 6400 1810 6460 1890
rect 6540 1810 6600 1890
rect 6400 1750 6600 1810
rect 6800 1890 7000 1950
rect 6800 1810 6860 1890
rect 6940 1810 7000 1890
rect 6800 1750 7000 1810
rect 7200 1890 7400 1950
rect 7200 1810 7260 1890
rect 7340 1810 7400 1890
rect 7200 1750 7400 1810
rect 7600 1890 7800 1950
rect 7600 1810 7660 1890
rect 7740 1810 7800 1890
rect 7600 1750 7800 1810
rect 8000 1890 8200 1950
rect 8000 1810 8060 1890
rect 8140 1810 8200 1890
rect 8000 1750 8200 1810
rect 8400 1890 8600 1950
rect 8400 1810 8460 1890
rect 8540 1810 8600 1890
rect 8400 1750 8600 1810
rect 8800 1890 9000 1950
rect 8800 1810 8860 1890
rect 8940 1810 9000 1890
rect 8800 1750 9000 1810
rect 9200 1890 9400 1950
rect 9200 1810 9260 1890
rect 9340 1810 9400 1890
rect 9200 1750 9400 1810
rect 9600 1890 9800 1950
rect 9600 1810 9660 1890
rect 9740 1810 9800 1890
rect 9600 1750 9800 1810
rect 2200 1690 2400 1750
rect 2200 1610 2260 1690
rect 2340 1610 2400 1690
rect 2200 1550 2400 1610
rect 2600 1690 2800 1750
rect 2600 1610 2660 1690
rect 2740 1610 2800 1690
rect 2600 1550 2800 1610
rect 3000 1690 3200 1750
rect 3000 1610 3060 1690
rect 3140 1610 3200 1690
rect 3000 1550 3200 1610
rect 3400 1690 3600 1750
rect 3400 1610 3460 1690
rect 3540 1610 3600 1690
rect 3400 1550 3600 1610
rect 3800 1690 4000 1750
rect 3800 1610 3860 1690
rect 3940 1610 4000 1690
rect 3800 1550 4000 1610
rect 4200 1690 4400 1750
rect 4200 1610 4260 1690
rect 4340 1610 4400 1690
rect 4200 1550 4400 1610
rect 4600 1690 4800 1750
rect 4600 1610 4660 1690
rect 4740 1610 4800 1690
rect 4600 1550 4800 1610
rect 5000 1690 5200 1750
rect 5000 1610 5060 1690
rect 5140 1610 5200 1690
rect 5000 1550 5200 1610
rect 5400 1690 5600 1750
rect 5400 1610 5460 1690
rect 5540 1610 5600 1690
rect 5400 1550 5600 1610
rect 5800 1690 6000 1750
rect 5800 1610 5860 1690
rect 5940 1610 6000 1690
rect 5800 1550 6000 1610
rect 6200 1690 6400 1750
rect 6200 1610 6260 1690
rect 6340 1610 6400 1690
rect 6200 1550 6400 1610
rect 6600 1690 6800 1750
rect 6600 1610 6660 1690
rect 6740 1610 6800 1690
rect 6600 1550 6800 1610
rect 7000 1690 7200 1750
rect 7000 1610 7060 1690
rect 7140 1610 7200 1690
rect 7000 1550 7200 1610
rect 7400 1690 7600 1750
rect 7400 1610 7460 1690
rect 7540 1610 7600 1690
rect 7400 1550 7600 1610
rect 7800 1690 8000 1750
rect 7800 1610 7860 1690
rect 7940 1610 8000 1690
rect 7800 1550 8000 1610
rect 8200 1690 8400 1750
rect 8200 1610 8260 1690
rect 8340 1610 8400 1690
rect 8200 1550 8400 1610
rect 8600 1690 8800 1750
rect 8600 1610 8660 1690
rect 8740 1610 8800 1690
rect 8600 1550 8800 1610
rect 9000 1690 9200 1750
rect 9000 1610 9060 1690
rect 9140 1610 9200 1690
rect 9000 1550 9200 1610
rect 9400 1690 9600 1750
rect 9400 1610 9460 1690
rect 9540 1610 9600 1690
rect 9400 1550 9600 1610
rect 9800 1690 10000 1750
rect 9800 1610 9860 1690
rect 9940 1610 10000 1690
rect 9800 1550 10000 1610
rect 2400 1490 2600 1550
rect 2400 1410 2460 1490
rect 2540 1410 2600 1490
rect 2400 1350 2600 1410
rect 2800 1490 3000 1550
rect 2800 1410 2860 1490
rect 2940 1410 3000 1490
rect 2800 1350 3000 1410
rect 3200 1490 3400 1550
rect 3200 1410 3260 1490
rect 3340 1410 3400 1490
rect 3200 1350 3400 1410
rect 3600 1490 3800 1550
rect 3600 1410 3660 1490
rect 3740 1410 3800 1490
rect 3600 1350 3800 1410
rect 4000 1490 4200 1550
rect 4000 1410 4060 1490
rect 4140 1410 4200 1490
rect 4000 1350 4200 1410
rect 4400 1490 4600 1550
rect 4400 1410 4460 1490
rect 4540 1410 4600 1490
rect 4400 1350 4600 1410
rect 4800 1490 5000 1550
rect 4800 1410 4860 1490
rect 4940 1410 5000 1490
rect 4800 1350 5000 1410
rect 5200 1490 5400 1550
rect 5200 1410 5260 1490
rect 5340 1410 5400 1490
rect 5200 1350 5400 1410
rect 5600 1490 5800 1550
rect 5600 1410 5660 1490
rect 5740 1410 5800 1490
rect 5600 1350 5800 1410
rect 6000 1490 6200 1550
rect 6000 1410 6060 1490
rect 6140 1410 6200 1490
rect 6000 1350 6200 1410
rect 6400 1490 6600 1550
rect 6400 1410 6460 1490
rect 6540 1410 6600 1490
rect 6400 1350 6600 1410
rect 6800 1490 7000 1550
rect 6800 1410 6860 1490
rect 6940 1410 7000 1490
rect 6800 1350 7000 1410
rect 7200 1490 7400 1550
rect 7200 1410 7260 1490
rect 7340 1410 7400 1490
rect 7200 1350 7400 1410
rect 7600 1490 7800 1550
rect 7600 1410 7660 1490
rect 7740 1410 7800 1490
rect 7600 1350 7800 1410
rect 8000 1490 8200 1550
rect 8000 1410 8060 1490
rect 8140 1410 8200 1490
rect 8000 1350 8200 1410
rect 8400 1490 8600 1550
rect 8400 1410 8460 1490
rect 8540 1410 8600 1490
rect 8400 1350 8600 1410
rect 8800 1490 9000 1550
rect 8800 1410 8860 1490
rect 8940 1410 9000 1490
rect 8800 1350 9000 1410
rect 9200 1490 9400 1550
rect 9200 1410 9260 1490
rect 9340 1410 9400 1490
rect 9200 1350 9400 1410
rect 9600 1490 9800 1550
rect 9600 1410 9660 1490
rect 9740 1410 9800 1490
rect 9600 1350 9800 1410
rect 2200 1290 2400 1350
rect 2200 1210 2260 1290
rect 2340 1210 2400 1290
rect 2200 1150 2400 1210
rect 2600 1290 2800 1350
rect 2600 1210 2660 1290
rect 2740 1210 2800 1290
rect 2600 1150 2800 1210
rect 3000 1290 3200 1350
rect 3000 1210 3060 1290
rect 3140 1210 3200 1290
rect 3000 1150 3200 1210
rect 3400 1290 3600 1350
rect 3400 1210 3460 1290
rect 3540 1210 3600 1290
rect 3400 1150 3600 1210
rect 3800 1290 4000 1350
rect 3800 1210 3860 1290
rect 3940 1210 4000 1290
rect 3800 1150 4000 1210
rect 4200 1290 4400 1350
rect 4200 1210 4260 1290
rect 4340 1210 4400 1290
rect 4200 1150 4400 1210
rect 4600 1290 4800 1350
rect 4600 1210 4660 1290
rect 4740 1210 4800 1290
rect 4600 1150 4800 1210
rect 5000 1290 5200 1350
rect 5000 1210 5060 1290
rect 5140 1210 5200 1290
rect 5000 1150 5200 1210
rect 5400 1290 5600 1350
rect 5400 1210 5460 1290
rect 5540 1210 5600 1290
rect 5400 1150 5600 1210
rect 5800 1290 6000 1350
rect 5800 1210 5860 1290
rect 5940 1210 6000 1290
rect 5800 1150 6000 1210
rect 6200 1290 6400 1350
rect 6200 1210 6260 1290
rect 6340 1210 6400 1290
rect 6200 1150 6400 1210
rect 6600 1290 6800 1350
rect 6600 1210 6660 1290
rect 6740 1210 6800 1290
rect 6600 1150 6800 1210
rect 7000 1290 7200 1350
rect 7000 1210 7060 1290
rect 7140 1210 7200 1290
rect 7000 1150 7200 1210
rect 7400 1290 7600 1350
rect 7400 1210 7460 1290
rect 7540 1210 7600 1290
rect 7400 1150 7600 1210
rect 7800 1290 8000 1350
rect 7800 1210 7860 1290
rect 7940 1210 8000 1290
rect 7800 1150 8000 1210
rect 8200 1290 8400 1350
rect 8200 1210 8260 1290
rect 8340 1210 8400 1290
rect 8200 1150 8400 1210
rect 8600 1290 8800 1350
rect 8600 1210 8660 1290
rect 8740 1210 8800 1290
rect 8600 1150 8800 1210
rect 9000 1290 9200 1350
rect 9000 1210 9060 1290
rect 9140 1210 9200 1290
rect 9000 1150 9200 1210
rect 9400 1290 9600 1350
rect 9400 1210 9460 1290
rect 9540 1210 9600 1290
rect 9400 1150 9600 1210
rect 9800 1290 10000 1350
rect 9800 1210 9860 1290
rect 9940 1210 10000 1290
rect 9800 1150 10000 1210
rect 2400 1090 2600 1150
rect 2400 1010 2460 1090
rect 2540 1010 2600 1090
rect 2400 950 2600 1010
rect 2800 1090 3000 1150
rect 2800 1010 2860 1090
rect 2940 1010 3000 1090
rect 2800 950 3000 1010
rect 3200 1090 3400 1150
rect 3200 1010 3260 1090
rect 3340 1010 3400 1090
rect 3200 950 3400 1010
rect 3600 1090 3800 1150
rect 3600 1010 3660 1090
rect 3740 1010 3800 1090
rect 3600 950 3800 1010
rect 4000 1090 4200 1150
rect 4000 1010 4060 1090
rect 4140 1010 4200 1090
rect 4000 950 4200 1010
rect 4400 1090 4600 1150
rect 4400 1010 4460 1090
rect 4540 1010 4600 1090
rect 4400 950 4600 1010
rect 4800 1090 5000 1150
rect 4800 1010 4860 1090
rect 4940 1010 5000 1090
rect 4800 950 5000 1010
rect 5200 1090 5400 1150
rect 5200 1010 5260 1090
rect 5340 1010 5400 1090
rect 5200 950 5400 1010
rect 5600 1090 5800 1150
rect 5600 1010 5660 1090
rect 5740 1010 5800 1090
rect 5600 950 5800 1010
rect 6000 1090 6200 1150
rect 6000 1010 6060 1090
rect 6140 1010 6200 1090
rect 6000 950 6200 1010
rect 6400 1090 6600 1150
rect 6400 1010 6460 1090
rect 6540 1010 6600 1090
rect 6400 950 6600 1010
rect 6800 1090 7000 1150
rect 6800 1010 6860 1090
rect 6940 1010 7000 1090
rect 6800 950 7000 1010
rect 7200 1090 7400 1150
rect 7200 1010 7260 1090
rect 7340 1010 7400 1090
rect 7200 950 7400 1010
rect 7600 1090 7800 1150
rect 7600 1010 7660 1090
rect 7740 1010 7800 1090
rect 7600 950 7800 1010
rect 8000 1090 8200 1150
rect 8000 1010 8060 1090
rect 8140 1010 8200 1090
rect 8000 950 8200 1010
rect 8400 1090 8600 1150
rect 8400 1010 8460 1090
rect 8540 1010 8600 1090
rect 8400 950 8600 1010
rect 8800 1090 9000 1150
rect 8800 1010 8860 1090
rect 8940 1010 9000 1090
rect 8800 950 9000 1010
rect 9200 1090 9400 1150
rect 9200 1010 9260 1090
rect 9340 1010 9400 1090
rect 9200 950 9400 1010
rect 9600 1090 9800 1150
rect 9600 1010 9660 1090
rect 9740 1010 9800 1090
rect 9600 950 9800 1010
rect 2200 890 2400 950
rect 2200 810 2260 890
rect 2340 810 2400 890
rect 2200 750 2400 810
rect 2600 890 2800 950
rect 2600 810 2660 890
rect 2740 810 2800 890
rect 2600 750 2800 810
rect 3000 890 3200 950
rect 3000 810 3060 890
rect 3140 810 3200 890
rect 3000 750 3200 810
rect 3400 890 3600 950
rect 3400 810 3460 890
rect 3540 810 3600 890
rect 3400 750 3600 810
rect 3800 890 4000 950
rect 3800 810 3860 890
rect 3940 810 4000 890
rect 3800 750 4000 810
rect 4200 890 4400 950
rect 4200 810 4260 890
rect 4340 810 4400 890
rect 4200 750 4400 810
rect 4600 890 4800 950
rect 4600 810 4660 890
rect 4740 810 4800 890
rect 4600 750 4800 810
rect 5000 890 5200 950
rect 5000 810 5060 890
rect 5140 810 5200 890
rect 5000 750 5200 810
rect 5400 890 5600 950
rect 5400 810 5460 890
rect 5540 810 5600 890
rect 5400 750 5600 810
rect 5800 890 6000 950
rect 5800 810 5860 890
rect 5940 810 6000 890
rect 5800 750 6000 810
rect 6200 890 6400 950
rect 6200 810 6260 890
rect 6340 810 6400 890
rect 6200 750 6400 810
rect 6600 890 6800 950
rect 6600 810 6660 890
rect 6740 810 6800 890
rect 6600 750 6800 810
rect 7000 890 7200 950
rect 7000 810 7060 890
rect 7140 810 7200 890
rect 7000 750 7200 810
rect 7400 890 7600 950
rect 7400 810 7460 890
rect 7540 810 7600 890
rect 7400 750 7600 810
rect 7800 890 8000 950
rect 7800 810 7860 890
rect 7940 810 8000 890
rect 7800 750 8000 810
rect 8200 890 8400 950
rect 8200 810 8260 890
rect 8340 810 8400 890
rect 8200 750 8400 810
rect 8600 890 8800 950
rect 8600 810 8660 890
rect 8740 810 8800 890
rect 8600 750 8800 810
rect 9000 890 9200 950
rect 9000 810 9060 890
rect 9140 810 9200 890
rect 9000 750 9200 810
rect 9400 890 9600 950
rect 9400 810 9460 890
rect 9540 810 9600 890
rect 9400 750 9600 810
rect 9800 890 10000 950
rect 9800 810 9860 890
rect 9940 810 10000 890
rect 9800 750 10000 810
rect 2400 690 2600 750
rect 2400 610 2460 690
rect 2540 610 2600 690
rect 2400 550 2600 610
rect 2800 690 3000 750
rect 2800 610 2860 690
rect 2940 610 3000 690
rect 2800 550 3000 610
rect 3200 690 3400 750
rect 3200 610 3260 690
rect 3340 610 3400 690
rect 3200 550 3400 610
rect 3600 690 3800 750
rect 3600 610 3660 690
rect 3740 610 3800 690
rect 3600 550 3800 610
rect 4000 690 4200 750
rect 4000 610 4060 690
rect 4140 610 4200 690
rect 4000 550 4200 610
rect 4400 690 4600 750
rect 4400 610 4460 690
rect 4540 610 4600 690
rect 4400 550 4600 610
rect 4800 690 5000 750
rect 4800 610 4860 690
rect 4940 610 5000 690
rect 4800 550 5000 610
rect 5200 690 5400 750
rect 5200 610 5260 690
rect 5340 610 5400 690
rect 5200 550 5400 610
rect 5600 690 5800 750
rect 5600 610 5660 690
rect 5740 610 5800 690
rect 5600 550 5800 610
rect 6000 690 6200 750
rect 6000 610 6060 690
rect 6140 610 6200 690
rect 6000 550 6200 610
rect 6400 690 6600 750
rect 6400 610 6460 690
rect 6540 610 6600 690
rect 6400 550 6600 610
rect 6800 690 7000 750
rect 6800 610 6860 690
rect 6940 610 7000 690
rect 6800 550 7000 610
rect 7200 690 7400 750
rect 7200 610 7260 690
rect 7340 610 7400 690
rect 7200 550 7400 610
rect 7600 690 7800 750
rect 7600 610 7660 690
rect 7740 610 7800 690
rect 7600 550 7800 610
rect 8000 690 8200 750
rect 8000 610 8060 690
rect 8140 610 8200 690
rect 8000 550 8200 610
rect 8400 690 8600 750
rect 8400 610 8460 690
rect 8540 610 8600 690
rect 8400 550 8600 610
rect 8800 690 9000 750
rect 8800 610 8860 690
rect 8940 610 9000 690
rect 8800 550 9000 610
rect 9200 690 9400 750
rect 9200 610 9260 690
rect 9340 610 9400 690
rect 9200 550 9400 610
rect 9600 690 9800 750
rect 9600 610 9660 690
rect 9740 610 9800 690
rect 9600 550 9800 610
rect 2200 490 2400 550
rect 2200 410 2260 490
rect 2340 410 2400 490
rect 2200 350 2400 410
rect 2600 490 2800 550
rect 2600 410 2660 490
rect 2740 410 2800 490
rect 2600 350 2800 410
rect 3000 490 3200 550
rect 3000 410 3060 490
rect 3140 410 3200 490
rect 3000 350 3200 410
rect 3400 490 3600 550
rect 3400 410 3460 490
rect 3540 410 3600 490
rect 3400 350 3600 410
rect 3800 490 4000 550
rect 3800 410 3860 490
rect 3940 410 4000 490
rect 3800 350 4000 410
rect 4200 490 4400 550
rect 4200 410 4260 490
rect 4340 410 4400 490
rect 4200 350 4400 410
rect 4600 490 4800 550
rect 4600 410 4660 490
rect 4740 410 4800 490
rect 4600 350 4800 410
rect 5000 490 5200 550
rect 5000 410 5060 490
rect 5140 410 5200 490
rect 5000 350 5200 410
rect 5400 490 5600 550
rect 5400 410 5460 490
rect 5540 410 5600 490
rect 5400 350 5600 410
rect 5800 490 6000 550
rect 5800 410 5860 490
rect 5940 410 6000 490
rect 5800 350 6000 410
rect 6200 490 6400 550
rect 6200 410 6260 490
rect 6340 410 6400 490
rect 6200 350 6400 410
rect 6600 490 6800 550
rect 6600 410 6660 490
rect 6740 410 6800 490
rect 6600 350 6800 410
rect 7000 490 7200 550
rect 7000 410 7060 490
rect 7140 410 7200 490
rect 7000 350 7200 410
rect 7400 490 7600 550
rect 7400 410 7460 490
rect 7540 410 7600 490
rect 7400 350 7600 410
rect 7800 490 8000 550
rect 7800 410 7860 490
rect 7940 410 8000 490
rect 7800 350 8000 410
rect 8200 490 8400 550
rect 8200 410 8260 490
rect 8340 410 8400 490
rect 8200 350 8400 410
rect 8600 490 8800 550
rect 8600 410 8660 490
rect 8740 410 8800 490
rect 8600 350 8800 410
rect 9000 490 9200 550
rect 9000 410 9060 490
rect 9140 410 9200 490
rect 9000 350 9200 410
rect 9400 490 9600 550
rect 9400 410 9460 490
rect 9540 410 9600 490
rect 9400 350 9600 410
rect 9800 490 10000 550
rect 9800 410 9860 490
rect 9940 410 10000 490
rect 9800 350 10000 410
rect 10100 250 10350 8250
rect 1850 0 10350 250
<< m3contact >>
rect 2460 7810 2540 7890
rect 2860 7810 2940 7890
rect 3260 7810 3340 7890
rect 3660 7810 3740 7890
rect 4060 7810 4140 7890
rect 4460 7810 4540 7890
rect 4860 7810 4940 7890
rect 5260 7810 5340 7890
rect 5660 7810 5740 7890
rect 6060 7810 6140 7890
rect 6460 7810 6540 7890
rect 6860 7810 6940 7890
rect 7260 7810 7340 7890
rect 7660 7810 7740 7890
rect 8060 7810 8140 7890
rect 8460 7810 8540 7890
rect 8860 7810 8940 7890
rect 9260 7810 9340 7890
rect 9660 7810 9740 7890
rect 2460 7410 2540 7490
rect 2860 7410 2940 7490
rect 3260 7410 3340 7490
rect 3660 7410 3740 7490
rect 4060 7410 4140 7490
rect 4460 7410 4540 7490
rect 4860 7410 4940 7490
rect 5260 7410 5340 7490
rect 5660 7410 5740 7490
rect 6060 7410 6140 7490
rect 6460 7410 6540 7490
rect 6860 7410 6940 7490
rect 7260 7410 7340 7490
rect 7660 7410 7740 7490
rect 8060 7410 8140 7490
rect 8460 7410 8540 7490
rect 8860 7410 8940 7490
rect 9260 7410 9340 7490
rect 9660 7410 9740 7490
rect 2460 7010 2540 7090
rect 2860 7010 2940 7090
rect 3260 7010 3340 7090
rect 3660 7010 3740 7090
rect 4060 7010 4140 7090
rect 4460 7010 4540 7090
rect 4860 7010 4940 7090
rect 5260 7010 5340 7090
rect 5660 7010 5740 7090
rect 6060 7010 6140 7090
rect 6460 7010 6540 7090
rect 6860 7010 6940 7090
rect 7260 7010 7340 7090
rect 7660 7010 7740 7090
rect 8060 7010 8140 7090
rect 8460 7010 8540 7090
rect 8860 7010 8940 7090
rect 9260 7010 9340 7090
rect 9660 7010 9740 7090
rect 2460 6610 2540 6690
rect 2860 6610 2940 6690
rect 3260 6610 3340 6690
rect 3660 6610 3740 6690
rect 4060 6610 4140 6690
rect 4460 6610 4540 6690
rect 4860 6610 4940 6690
rect 5260 6610 5340 6690
rect 5660 6610 5740 6690
rect 6060 6610 6140 6690
rect 6460 6610 6540 6690
rect 6860 6610 6940 6690
rect 7260 6610 7340 6690
rect 7660 6610 7740 6690
rect 8060 6610 8140 6690
rect 8460 6610 8540 6690
rect 8860 6610 8940 6690
rect 9260 6610 9340 6690
rect 9660 6610 9740 6690
rect 2460 6210 2540 6290
rect 2860 6210 2940 6290
rect 3260 6210 3340 6290
rect 3660 6210 3740 6290
rect 4060 6210 4140 6290
rect 4460 6210 4540 6290
rect 4860 6210 4940 6290
rect 5260 6210 5340 6290
rect 5660 6210 5740 6290
rect 6060 6210 6140 6290
rect 6460 6210 6540 6290
rect 6860 6210 6940 6290
rect 7260 6210 7340 6290
rect 7660 6210 7740 6290
rect 8060 6210 8140 6290
rect 8460 6210 8540 6290
rect 8860 6210 8940 6290
rect 9260 6210 9340 6290
rect 9660 6210 9740 6290
rect 2460 5810 2540 5890
rect 2860 5810 2940 5890
rect 3260 5810 3340 5890
rect 3660 5810 3740 5890
rect 4060 5810 4140 5890
rect 4460 5810 4540 5890
rect 4860 5810 4940 5890
rect 5260 5810 5340 5890
rect 5660 5810 5740 5890
rect 6060 5810 6140 5890
rect 6460 5810 6540 5890
rect 6860 5810 6940 5890
rect 7260 5810 7340 5890
rect 7660 5810 7740 5890
rect 8060 5810 8140 5890
rect 8460 5810 8540 5890
rect 8860 5810 8940 5890
rect 9260 5810 9340 5890
rect 9660 5810 9740 5890
rect 2460 5410 2540 5490
rect 2860 5410 2940 5490
rect 3260 5410 3340 5490
rect 3660 5410 3740 5490
rect 4060 5410 4140 5490
rect 4460 5410 4540 5490
rect 4860 5410 4940 5490
rect 5260 5410 5340 5490
rect 5660 5410 5740 5490
rect 6060 5410 6140 5490
rect 6460 5410 6540 5490
rect 6860 5410 6940 5490
rect 7260 5410 7340 5490
rect 7660 5410 7740 5490
rect 8060 5410 8140 5490
rect 8460 5410 8540 5490
rect 8860 5410 8940 5490
rect 9260 5410 9340 5490
rect 9660 5410 9740 5490
rect 2460 5010 2540 5090
rect 2860 5010 2940 5090
rect 3260 5010 3340 5090
rect 3660 5010 3740 5090
rect 4060 5010 4140 5090
rect 4460 5010 4540 5090
rect 4860 5010 4940 5090
rect 5260 5010 5340 5090
rect 5660 5010 5740 5090
rect 6060 5010 6140 5090
rect 6460 5010 6540 5090
rect 6860 5010 6940 5090
rect 7260 5010 7340 5090
rect 7660 5010 7740 5090
rect 8060 5010 8140 5090
rect 8460 5010 8540 5090
rect 8860 5010 8940 5090
rect 9260 5010 9340 5090
rect 9660 5010 9740 5090
rect 2460 4610 2540 4690
rect 2860 4610 2940 4690
rect 3260 4610 3340 4690
rect 3660 4610 3740 4690
rect 4060 4610 4140 4690
rect 4460 4610 4540 4690
rect 4860 4610 4940 4690
rect 5260 4610 5340 4690
rect 5660 4610 5740 4690
rect 6060 4610 6140 4690
rect 6460 4610 6540 4690
rect 6860 4610 6940 4690
rect 7260 4610 7340 4690
rect 7660 4610 7740 4690
rect 8060 4610 8140 4690
rect 8460 4610 8540 4690
rect 8860 4610 8940 4690
rect 9260 4610 9340 4690
rect 9660 4610 9740 4690
rect 2460 4210 2540 4290
rect 2860 4210 2940 4290
rect 3260 4210 3340 4290
rect 3660 4210 3740 4290
rect 4060 4210 4140 4290
rect 4460 4210 4540 4290
rect 4860 4210 4940 4290
rect 5260 4210 5340 4290
rect 5660 4210 5740 4290
rect 6060 4210 6140 4290
rect 6460 4210 6540 4290
rect 6860 4210 6940 4290
rect 7260 4210 7340 4290
rect 7660 4210 7740 4290
rect 8060 4210 8140 4290
rect 8460 4210 8540 4290
rect 8860 4210 8940 4290
rect 9260 4210 9340 4290
rect 9660 4210 9740 4290
rect 2460 3810 2540 3890
rect 2860 3810 2940 3890
rect 3260 3810 3340 3890
rect 3660 3810 3740 3890
rect 4060 3810 4140 3890
rect 4460 3810 4540 3890
rect 4860 3810 4940 3890
rect 5260 3810 5340 3890
rect 5660 3810 5740 3890
rect 6060 3810 6140 3890
rect 6460 3810 6540 3890
rect 6860 3810 6940 3890
rect 7260 3810 7340 3890
rect 7660 3810 7740 3890
rect 8060 3810 8140 3890
rect 8460 3810 8540 3890
rect 8860 3810 8940 3890
rect 9260 3810 9340 3890
rect 9660 3810 9740 3890
rect 2460 3410 2540 3490
rect 2860 3410 2940 3490
rect 3260 3410 3340 3490
rect 3660 3410 3740 3490
rect 4060 3410 4140 3490
rect 4460 3410 4540 3490
rect 4860 3410 4940 3490
rect 5260 3410 5340 3490
rect 5660 3410 5740 3490
rect 6060 3410 6140 3490
rect 6460 3410 6540 3490
rect 6860 3410 6940 3490
rect 7260 3410 7340 3490
rect 7660 3410 7740 3490
rect 8060 3410 8140 3490
rect 8460 3410 8540 3490
rect 8860 3410 8940 3490
rect 9260 3410 9340 3490
rect 9660 3410 9740 3490
rect 2460 3010 2540 3090
rect 2860 3010 2940 3090
rect 3260 3010 3340 3090
rect 3660 3010 3740 3090
rect 4060 3010 4140 3090
rect 4460 3010 4540 3090
rect 4860 3010 4940 3090
rect 5260 3010 5340 3090
rect 5660 3010 5740 3090
rect 6060 3010 6140 3090
rect 6460 3010 6540 3090
rect 6860 3010 6940 3090
rect 7260 3010 7340 3090
rect 7660 3010 7740 3090
rect 8060 3010 8140 3090
rect 8460 3010 8540 3090
rect 8860 3010 8940 3090
rect 9260 3010 9340 3090
rect 9660 3010 9740 3090
rect 2460 2610 2540 2690
rect 2860 2610 2940 2690
rect 3260 2610 3340 2690
rect 3660 2610 3740 2690
rect 4060 2610 4140 2690
rect 4460 2610 4540 2690
rect 4860 2610 4940 2690
rect 5260 2610 5340 2690
rect 5660 2610 5740 2690
rect 6060 2610 6140 2690
rect 6460 2610 6540 2690
rect 6860 2610 6940 2690
rect 7260 2610 7340 2690
rect 7660 2610 7740 2690
rect 8060 2610 8140 2690
rect 8460 2610 8540 2690
rect 8860 2610 8940 2690
rect 9260 2610 9340 2690
rect 9660 2610 9740 2690
rect 2460 2210 2540 2290
rect 2860 2210 2940 2290
rect 3260 2210 3340 2290
rect 3660 2210 3740 2290
rect 4060 2210 4140 2290
rect 4460 2210 4540 2290
rect 4860 2210 4940 2290
rect 5260 2210 5340 2290
rect 5660 2210 5740 2290
rect 6060 2210 6140 2290
rect 6460 2210 6540 2290
rect 6860 2210 6940 2290
rect 7260 2210 7340 2290
rect 7660 2210 7740 2290
rect 8060 2210 8140 2290
rect 8460 2210 8540 2290
rect 8860 2210 8940 2290
rect 9260 2210 9340 2290
rect 9660 2210 9740 2290
rect 2460 1810 2540 1890
rect 2860 1810 2940 1890
rect 3260 1810 3340 1890
rect 3660 1810 3740 1890
rect 4060 1810 4140 1890
rect 4460 1810 4540 1890
rect 4860 1810 4940 1890
rect 5260 1810 5340 1890
rect 5660 1810 5740 1890
rect 6060 1810 6140 1890
rect 6460 1810 6540 1890
rect 6860 1810 6940 1890
rect 7260 1810 7340 1890
rect 7660 1810 7740 1890
rect 8060 1810 8140 1890
rect 8460 1810 8540 1890
rect 8860 1810 8940 1890
rect 9260 1810 9340 1890
rect 9660 1810 9740 1890
rect 2460 1410 2540 1490
rect 2860 1410 2940 1490
rect 3260 1410 3340 1490
rect 3660 1410 3740 1490
rect 4060 1410 4140 1490
rect 4460 1410 4540 1490
rect 4860 1410 4940 1490
rect 5260 1410 5340 1490
rect 5660 1410 5740 1490
rect 6060 1410 6140 1490
rect 6460 1410 6540 1490
rect 6860 1410 6940 1490
rect 7260 1410 7340 1490
rect 7660 1410 7740 1490
rect 8060 1410 8140 1490
rect 8460 1410 8540 1490
rect 8860 1410 8940 1490
rect 9260 1410 9340 1490
rect 9660 1410 9740 1490
rect 2460 1010 2540 1090
rect 2860 1010 2940 1090
rect 3260 1010 3340 1090
rect 3660 1010 3740 1090
rect 4060 1010 4140 1090
rect 4460 1010 4540 1090
rect 4860 1010 4940 1090
rect 5260 1010 5340 1090
rect 5660 1010 5740 1090
rect 6060 1010 6140 1090
rect 6460 1010 6540 1090
rect 6860 1010 6940 1090
rect 7260 1010 7340 1090
rect 7660 1010 7740 1090
rect 8060 1010 8140 1090
rect 8460 1010 8540 1090
rect 8860 1010 8940 1090
rect 9260 1010 9340 1090
rect 9660 1010 9740 1090
rect 2460 610 2540 690
rect 2860 610 2940 690
rect 3260 610 3340 690
rect 3660 610 3740 690
rect 4060 610 4140 690
rect 4460 610 4540 690
rect 4860 610 4940 690
rect 5260 610 5340 690
rect 5660 610 5740 690
rect 6060 610 6140 690
rect 6460 610 6540 690
rect 6860 610 6940 690
rect 7260 610 7340 690
rect 7660 610 7740 690
rect 8060 610 8140 690
rect 8460 610 8540 690
rect 8860 610 8940 690
rect 9260 610 9340 690
rect 9660 610 9740 690
<< metal3 >>
rect 100 32550 12100 34210
rect 100 30250 12100 31910
rect 100 20450 12100 28250
rect 100 9150 12100 16950
rect 1850 8250 10350 8500
rect 1850 250 2100 8250
rect 10100 250 10350 8250
rect 1850 0 10350 250
<< pad >>
rect 2100 7890 10100 8250
rect 2100 7810 2460 7890
rect 2540 7810 2860 7890
rect 2940 7810 3260 7890
rect 3340 7810 3660 7890
rect 3740 7810 4060 7890
rect 4140 7810 4460 7890
rect 4540 7810 4860 7890
rect 4940 7810 5260 7890
rect 5340 7810 5660 7890
rect 5740 7810 6060 7890
rect 6140 7810 6460 7890
rect 6540 7810 6860 7890
rect 6940 7810 7260 7890
rect 7340 7810 7660 7890
rect 7740 7810 8060 7890
rect 8140 7810 8460 7890
rect 8540 7810 8860 7890
rect 8940 7810 9260 7890
rect 9340 7810 9660 7890
rect 9740 7810 10100 7890
rect 2100 7490 10100 7810
rect 2100 7410 2460 7490
rect 2540 7410 2860 7490
rect 2940 7410 3260 7490
rect 3340 7410 3660 7490
rect 3740 7410 4060 7490
rect 4140 7410 4460 7490
rect 4540 7410 4860 7490
rect 4940 7410 5260 7490
rect 5340 7410 5660 7490
rect 5740 7410 6060 7490
rect 6140 7410 6460 7490
rect 6540 7410 6860 7490
rect 6940 7410 7260 7490
rect 7340 7410 7660 7490
rect 7740 7410 8060 7490
rect 8140 7410 8460 7490
rect 8540 7410 8860 7490
rect 8940 7410 9260 7490
rect 9340 7410 9660 7490
rect 9740 7410 10100 7490
rect 2100 7090 10100 7410
rect 2100 7010 2460 7090
rect 2540 7010 2860 7090
rect 2940 7010 3260 7090
rect 3340 7010 3660 7090
rect 3740 7010 4060 7090
rect 4140 7010 4460 7090
rect 4540 7010 4860 7090
rect 4940 7010 5260 7090
rect 5340 7010 5660 7090
rect 5740 7010 6060 7090
rect 6140 7010 6460 7090
rect 6540 7010 6860 7090
rect 6940 7010 7260 7090
rect 7340 7010 7660 7090
rect 7740 7010 8060 7090
rect 8140 7010 8460 7090
rect 8540 7010 8860 7090
rect 8940 7010 9260 7090
rect 9340 7010 9660 7090
rect 9740 7010 10100 7090
rect 2100 6690 10100 7010
rect 2100 6610 2460 6690
rect 2540 6610 2860 6690
rect 2940 6610 3260 6690
rect 3340 6610 3660 6690
rect 3740 6610 4060 6690
rect 4140 6610 4460 6690
rect 4540 6610 4860 6690
rect 4940 6610 5260 6690
rect 5340 6610 5660 6690
rect 5740 6610 6060 6690
rect 6140 6610 6460 6690
rect 6540 6610 6860 6690
rect 6940 6610 7260 6690
rect 7340 6610 7660 6690
rect 7740 6610 8060 6690
rect 8140 6610 8460 6690
rect 8540 6610 8860 6690
rect 8940 6610 9260 6690
rect 9340 6610 9660 6690
rect 9740 6610 10100 6690
rect 2100 6290 10100 6610
rect 2100 6210 2460 6290
rect 2540 6210 2860 6290
rect 2940 6210 3260 6290
rect 3340 6210 3660 6290
rect 3740 6210 4060 6290
rect 4140 6210 4460 6290
rect 4540 6210 4860 6290
rect 4940 6210 5260 6290
rect 5340 6210 5660 6290
rect 5740 6210 6060 6290
rect 6140 6210 6460 6290
rect 6540 6210 6860 6290
rect 6940 6210 7260 6290
rect 7340 6210 7660 6290
rect 7740 6210 8060 6290
rect 8140 6210 8460 6290
rect 8540 6210 8860 6290
rect 8940 6210 9260 6290
rect 9340 6210 9660 6290
rect 9740 6210 10100 6290
rect 2100 5890 10100 6210
rect 2100 5810 2460 5890
rect 2540 5810 2860 5890
rect 2940 5810 3260 5890
rect 3340 5810 3660 5890
rect 3740 5810 4060 5890
rect 4140 5810 4460 5890
rect 4540 5810 4860 5890
rect 4940 5810 5260 5890
rect 5340 5810 5660 5890
rect 5740 5810 6060 5890
rect 6140 5810 6460 5890
rect 6540 5810 6860 5890
rect 6940 5810 7260 5890
rect 7340 5810 7660 5890
rect 7740 5810 8060 5890
rect 8140 5810 8460 5890
rect 8540 5810 8860 5890
rect 8940 5810 9260 5890
rect 9340 5810 9660 5890
rect 9740 5810 10100 5890
rect 2100 5490 10100 5810
rect 2100 5410 2460 5490
rect 2540 5410 2860 5490
rect 2940 5410 3260 5490
rect 3340 5410 3660 5490
rect 3740 5410 4060 5490
rect 4140 5410 4460 5490
rect 4540 5410 4860 5490
rect 4940 5410 5260 5490
rect 5340 5410 5660 5490
rect 5740 5410 6060 5490
rect 6140 5410 6460 5490
rect 6540 5410 6860 5490
rect 6940 5410 7260 5490
rect 7340 5410 7660 5490
rect 7740 5410 8060 5490
rect 8140 5410 8460 5490
rect 8540 5410 8860 5490
rect 8940 5410 9260 5490
rect 9340 5410 9660 5490
rect 9740 5410 10100 5490
rect 2100 5090 10100 5410
rect 2100 5010 2460 5090
rect 2540 5010 2860 5090
rect 2940 5010 3260 5090
rect 3340 5010 3660 5090
rect 3740 5010 4060 5090
rect 4140 5010 4460 5090
rect 4540 5010 4860 5090
rect 4940 5010 5260 5090
rect 5340 5010 5660 5090
rect 5740 5010 6060 5090
rect 6140 5010 6460 5090
rect 6540 5010 6860 5090
rect 6940 5010 7260 5090
rect 7340 5010 7660 5090
rect 7740 5010 8060 5090
rect 8140 5010 8460 5090
rect 8540 5010 8860 5090
rect 8940 5010 9260 5090
rect 9340 5010 9660 5090
rect 9740 5010 10100 5090
rect 2100 4690 10100 5010
rect 2100 4610 2460 4690
rect 2540 4610 2860 4690
rect 2940 4610 3260 4690
rect 3340 4610 3660 4690
rect 3740 4610 4060 4690
rect 4140 4610 4460 4690
rect 4540 4610 4860 4690
rect 4940 4610 5260 4690
rect 5340 4610 5660 4690
rect 5740 4610 6060 4690
rect 6140 4610 6460 4690
rect 6540 4610 6860 4690
rect 6940 4610 7260 4690
rect 7340 4610 7660 4690
rect 7740 4610 8060 4690
rect 8140 4610 8460 4690
rect 8540 4610 8860 4690
rect 8940 4610 9260 4690
rect 9340 4610 9660 4690
rect 9740 4610 10100 4690
rect 2100 4290 10100 4610
rect 2100 4210 2460 4290
rect 2540 4210 2860 4290
rect 2940 4210 3260 4290
rect 3340 4210 3660 4290
rect 3740 4210 4060 4290
rect 4140 4210 4460 4290
rect 4540 4210 4860 4290
rect 4940 4210 5260 4290
rect 5340 4210 5660 4290
rect 5740 4210 6060 4290
rect 6140 4210 6460 4290
rect 6540 4210 6860 4290
rect 6940 4210 7260 4290
rect 7340 4210 7660 4290
rect 7740 4210 8060 4290
rect 8140 4210 8460 4290
rect 8540 4210 8860 4290
rect 8940 4210 9260 4290
rect 9340 4210 9660 4290
rect 9740 4210 10100 4290
rect 2100 3890 10100 4210
rect 2100 3810 2460 3890
rect 2540 3810 2860 3890
rect 2940 3810 3260 3890
rect 3340 3810 3660 3890
rect 3740 3810 4060 3890
rect 4140 3810 4460 3890
rect 4540 3810 4860 3890
rect 4940 3810 5260 3890
rect 5340 3810 5660 3890
rect 5740 3810 6060 3890
rect 6140 3810 6460 3890
rect 6540 3810 6860 3890
rect 6940 3810 7260 3890
rect 7340 3810 7660 3890
rect 7740 3810 8060 3890
rect 8140 3810 8460 3890
rect 8540 3810 8860 3890
rect 8940 3810 9260 3890
rect 9340 3810 9660 3890
rect 9740 3810 10100 3890
rect 2100 3490 10100 3810
rect 2100 3410 2460 3490
rect 2540 3410 2860 3490
rect 2940 3410 3260 3490
rect 3340 3410 3660 3490
rect 3740 3410 4060 3490
rect 4140 3410 4460 3490
rect 4540 3410 4860 3490
rect 4940 3410 5260 3490
rect 5340 3410 5660 3490
rect 5740 3410 6060 3490
rect 6140 3410 6460 3490
rect 6540 3410 6860 3490
rect 6940 3410 7260 3490
rect 7340 3410 7660 3490
rect 7740 3410 8060 3490
rect 8140 3410 8460 3490
rect 8540 3410 8860 3490
rect 8940 3410 9260 3490
rect 9340 3410 9660 3490
rect 9740 3410 10100 3490
rect 2100 3090 10100 3410
rect 2100 3010 2460 3090
rect 2540 3010 2860 3090
rect 2940 3010 3260 3090
rect 3340 3010 3660 3090
rect 3740 3010 4060 3090
rect 4140 3010 4460 3090
rect 4540 3010 4860 3090
rect 4940 3010 5260 3090
rect 5340 3010 5660 3090
rect 5740 3010 6060 3090
rect 6140 3010 6460 3090
rect 6540 3010 6860 3090
rect 6940 3010 7260 3090
rect 7340 3010 7660 3090
rect 7740 3010 8060 3090
rect 8140 3010 8460 3090
rect 8540 3010 8860 3090
rect 8940 3010 9260 3090
rect 9340 3010 9660 3090
rect 9740 3010 10100 3090
rect 2100 2690 10100 3010
rect 2100 2610 2460 2690
rect 2540 2610 2860 2690
rect 2940 2610 3260 2690
rect 3340 2610 3660 2690
rect 3740 2610 4060 2690
rect 4140 2610 4460 2690
rect 4540 2610 4860 2690
rect 4940 2610 5260 2690
rect 5340 2610 5660 2690
rect 5740 2610 6060 2690
rect 6140 2610 6460 2690
rect 6540 2610 6860 2690
rect 6940 2610 7260 2690
rect 7340 2610 7660 2690
rect 7740 2610 8060 2690
rect 8140 2610 8460 2690
rect 8540 2610 8860 2690
rect 8940 2610 9260 2690
rect 9340 2610 9660 2690
rect 9740 2610 10100 2690
rect 2100 2290 10100 2610
rect 2100 2210 2460 2290
rect 2540 2210 2860 2290
rect 2940 2210 3260 2290
rect 3340 2210 3660 2290
rect 3740 2210 4060 2290
rect 4140 2210 4460 2290
rect 4540 2210 4860 2290
rect 4940 2210 5260 2290
rect 5340 2210 5660 2290
rect 5740 2210 6060 2290
rect 6140 2210 6460 2290
rect 6540 2210 6860 2290
rect 6940 2210 7260 2290
rect 7340 2210 7660 2290
rect 7740 2210 8060 2290
rect 8140 2210 8460 2290
rect 8540 2210 8860 2290
rect 8940 2210 9260 2290
rect 9340 2210 9660 2290
rect 9740 2210 10100 2290
rect 2100 1890 10100 2210
rect 2100 1810 2460 1890
rect 2540 1810 2860 1890
rect 2940 1810 3260 1890
rect 3340 1810 3660 1890
rect 3740 1810 4060 1890
rect 4140 1810 4460 1890
rect 4540 1810 4860 1890
rect 4940 1810 5260 1890
rect 5340 1810 5660 1890
rect 5740 1810 6060 1890
rect 6140 1810 6460 1890
rect 6540 1810 6860 1890
rect 6940 1810 7260 1890
rect 7340 1810 7660 1890
rect 7740 1810 8060 1890
rect 8140 1810 8460 1890
rect 8540 1810 8860 1890
rect 8940 1810 9260 1890
rect 9340 1810 9660 1890
rect 9740 1810 10100 1890
rect 2100 1490 10100 1810
rect 2100 1410 2460 1490
rect 2540 1410 2860 1490
rect 2940 1410 3260 1490
rect 3340 1410 3660 1490
rect 3740 1410 4060 1490
rect 4140 1410 4460 1490
rect 4540 1410 4860 1490
rect 4940 1410 5260 1490
rect 5340 1410 5660 1490
rect 5740 1410 6060 1490
rect 6140 1410 6460 1490
rect 6540 1410 6860 1490
rect 6940 1410 7260 1490
rect 7340 1410 7660 1490
rect 7740 1410 8060 1490
rect 8140 1410 8460 1490
rect 8540 1410 8860 1490
rect 8940 1410 9260 1490
rect 9340 1410 9660 1490
rect 9740 1410 10100 1490
rect 2100 1090 10100 1410
rect 2100 1010 2460 1090
rect 2540 1010 2860 1090
rect 2940 1010 3260 1090
rect 3340 1010 3660 1090
rect 3740 1010 4060 1090
rect 4140 1010 4460 1090
rect 4540 1010 4860 1090
rect 4940 1010 5260 1090
rect 5340 1010 5660 1090
rect 5740 1010 6060 1090
rect 6140 1010 6460 1090
rect 6540 1010 6860 1090
rect 6940 1010 7260 1090
rect 7340 1010 7660 1090
rect 7740 1010 8060 1090
rect 8140 1010 8460 1090
rect 8540 1010 8860 1090
rect 8940 1010 9260 1090
rect 9340 1010 9660 1090
rect 9740 1010 10100 1090
rect 2100 690 10100 1010
rect 2100 610 2460 690
rect 2540 610 2860 690
rect 2940 610 3260 690
rect 3340 610 3660 690
rect 3740 610 4060 690
rect 4140 610 4460 690
rect 4540 610 4860 690
rect 4940 610 5260 690
rect 5340 610 5660 690
rect 5740 610 6060 690
rect 6140 610 6460 690
rect 6540 610 6860 690
rect 6940 610 7260 690
rect 7340 610 7660 690
rect 7740 610 8060 690
rect 8140 610 8460 690
rect 8540 610 8860 690
rect 8940 610 9260 690
rect 9340 610 9660 690
rect 9740 610 10100 690
rect 2100 250 10100 610
use IOFILLER50  IOFILLER50_0
timestamp 1537935238
transform 1 0 6600 0 1 9150
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1537935238
transform 1 0 600 0 1 9150
box -35 0 5035 25060
<< end >>
