magic
tech scmos
magscale 1 2
timestamp 1726842831
<< nwell >>
rect -12 154 133 272
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 60 14 64 54
rect 80 14 84 54
<< ptransistor >>
rect 20 166 24 246
rect 40 166 44 246
rect 60 166 64 246
rect 80 166 84 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 14 26 54
rect 38 14 40 54
rect 44 14 46 54
rect 58 14 60 54
rect 64 14 66 54
rect 78 14 80 54
rect 84 14 86 54
<< pdiffusion >>
rect 18 166 20 246
rect 24 166 26 246
rect 38 166 40 246
rect 44 166 46 246
rect 58 166 60 246
rect 64 166 66 246
rect 78 166 80 246
rect 84 166 86 246
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 54
rect 46 14 58 54
rect 66 14 78 54
rect 86 14 98 54
<< pdcontact >>
rect 6 166 18 246
rect 26 166 38 246
rect 46 166 58 246
rect 66 166 78 246
rect 86 166 98 246
<< psubstratepcontact >>
rect -6 -6 126 6
<< nsubstratencontact >>
rect -6 254 126 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 80 246 84 250
rect 20 162 24 166
rect 40 162 44 166
rect 60 162 64 166
rect 80 162 84 166
rect 20 158 84 162
rect 20 62 24 158
rect 20 58 84 62
rect 20 54 24 58
rect 40 54 44 58
rect 60 54 64 58
rect 80 54 84 58
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
rect 80 10 84 14
<< polycontact >>
rect 24 117 36 129
<< metal1 >>
rect -6 266 126 268
rect -6 252 126 254
rect 6 246 18 252
rect 46 246 58 252
rect 86 246 98 252
rect 26 160 38 166
rect 66 160 74 166
rect 26 154 74 160
rect 66 117 74 154
rect 66 68 74 103
rect 26 60 74 68
rect 26 54 34 60
rect 66 54 74 60
rect 6 8 18 14
rect 46 8 58 14
rect 86 8 98 14
rect -6 6 126 8
rect -6 -8 126 -6
<< m2contact >>
rect 23 103 37 117
rect 63 103 77 117
<< metal2 >>
rect 66 117 74 135
rect 26 87 34 103
<< m1p >>
rect -6 252 126 268
rect -6 -8 126 8
<< m2p >>
rect 66 119 74 135
rect 26 87 34 101
<< labels >>
rlabel metal1 -6 252 106 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -6 -8 106 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal2 30 89 30 89 1 A
port 1 n signal input
rlabel metal2 70 131 70 131 1 Y
port 2 n signal output
<< properties >>
string FIXED_BBOX 0 0 120 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
