magic
tech scmos
magscale 1 6
timestamp 1554524574
<< checkpaint >>
rect -136 -136 280 388
<< nwell >>
rect -16 -16 160 244
<< ptransistor >>
rect 49 14 59 214
<< pdiffusion >>
rect 12 204 49 214
rect 12 192 22 204
rect 34 192 49 204
rect 12 180 49 192
rect 12 168 22 180
rect 34 168 49 180
rect 12 156 49 168
rect 12 144 22 156
rect 34 144 49 156
rect 12 132 49 144
rect 12 120 22 132
rect 34 120 49 132
rect 12 108 49 120
rect 12 96 22 108
rect 34 96 49 108
rect 12 84 49 96
rect 12 72 22 84
rect 34 72 49 84
rect 12 60 49 72
rect 12 48 22 60
rect 34 48 49 60
rect 12 36 49 48
rect 12 24 22 36
rect 34 24 49 36
rect 12 14 49 24
rect 59 204 96 214
rect 59 192 74 204
rect 86 192 96 204
rect 59 180 96 192
rect 59 168 74 180
rect 86 168 96 180
rect 59 156 96 168
rect 59 144 74 156
rect 86 144 96 156
rect 59 132 96 144
rect 59 120 74 132
rect 86 120 96 132
rect 59 108 96 120
rect 59 96 74 108
rect 86 96 96 108
rect 59 84 96 96
rect 59 72 74 84
rect 86 72 96 84
rect 59 60 96 72
rect 59 48 74 60
rect 86 48 96 60
rect 59 36 96 48
rect 59 24 74 36
rect 86 24 96 36
rect 59 14 96 24
<< pdcontact >>
rect 22 192 34 204
rect 22 168 34 180
rect 22 144 34 156
rect 22 120 34 132
rect 22 96 34 108
rect 22 72 34 84
rect 22 48 34 60
rect 22 24 34 36
rect 74 192 86 204
rect 74 168 86 180
rect 74 144 86 156
rect 74 120 86 132
rect 74 96 86 108
rect 74 72 86 84
rect 74 48 86 60
rect 74 24 86 36
<< polysilicon >>
rect 49 214 59 234
rect 49 4 59 14
<< metal1 >>
rect 10 204 46 216
rect 10 192 22 204
rect 34 192 46 204
rect 10 180 46 192
rect 10 168 22 180
rect 34 168 46 180
rect 10 156 46 168
rect 10 144 22 156
rect 34 144 46 156
rect 10 132 46 144
rect 10 120 22 132
rect 34 120 46 132
rect 10 108 46 120
rect 10 96 22 108
rect 34 96 46 108
rect 10 84 46 96
rect 10 72 22 84
rect 34 72 46 84
rect 10 60 46 72
rect 10 48 22 60
rect 34 48 46 60
rect 10 36 46 48
rect 10 24 22 36
rect 34 24 46 36
rect 10 12 46 24
rect 62 204 98 216
rect 62 192 74 204
rect 86 192 98 204
rect 62 180 98 192
rect 62 168 74 180
rect 86 168 98 180
rect 62 156 98 168
rect 62 144 74 156
rect 86 144 98 156
rect 62 132 98 144
rect 62 120 74 132
rect 86 120 98 132
rect 62 108 98 120
rect 62 96 74 108
rect 86 96 98 108
rect 62 84 98 96
rect 62 72 74 84
rect 86 72 98 84
rect 62 60 98 72
rect 62 48 74 60
rect 86 48 98 60
rect 62 36 98 48
rect 62 24 74 36
rect 86 24 98 36
rect 62 12 98 24
use ntap_CDNS_7230122529111  ntap_CDNS_7230122529111_0
timestamp 1554524574
transform 1 0 108 0 1 4
box 8 8 44 208
use poly1cont_CDNS_723012252918  poly1cont_CDNS_723012252918_0
timestamp 1554524574
transform 1 0 36 0 1 232
box 0 0 36 36
<< end >>
