magic
tech scmos
timestamp 1701862152
<< checkpaint >>
rect -17 71 27 79
rect -17 39 37 71
rect -7 30 37 39
<< nwell >>
rect -6 77 26 136
<< ntransistor >>
rect 9 7 11 27
<< ptransistor >>
rect 9 83 11 123
<< ndiffusion >>
rect 8 7 9 27
rect 11 7 12 27
<< pdiffusion >>
rect 8 83 9 123
rect 11 83 12 123
<< ndcontact >>
rect 2 7 8 27
rect 12 7 18 27
<< pdcontact >>
rect 2 83 8 123
rect 12 83 18 123
<< psubstratepcontact >>
rect -3 -3 23 3
<< nsubstratencontact >>
rect -3 127 23 133
<< polysilicon >>
rect 9 123 11 125
rect 9 51 11 83
rect 8 45 11 51
rect 9 27 11 45
rect 9 5 11 7
<< polycontact >>
rect 2 45 8 51
<< metal1 >>
rect -3 133 23 134
rect -3 126 23 127
rect 2 123 8 126
rect 12 58 16 83
rect 12 27 16 51
rect 2 4 8 7
rect -3 3 23 4
rect -3 -4 23 -3
<< m2contact >>
rect 1 51 8 58
rect 11 51 18 58
<< metal2 >>
rect 3 58 7 67
rect 13 43 17 51
<< m1p >>
rect -3 126 23 134
rect -3 -4 23 4
<< m2p >>
rect 3 59 7 67
rect 13 43 17 50
<< labels >>
rlabel metal2 5 65 5 65 1 A
port 1 n signal input
rlabel metal2 15 44 15 44 5 Y
port 2 n signal output
rlabel metal1 -3 126 23 134 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -3 -4 23 4 0 gnd
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 20 130
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
