magic
tech scmos
timestamp 1702508443
<< nwell >>
rect -6 77 46 136
<< ntransistor >>
rect 12 7 14 27
rect 17 7 19 27
rect 27 7 29 17
<< ptransistor >>
rect 9 83 11 123
rect 19 83 21 123
rect 29 83 31 123
<< ndiffusion >>
rect 11 7 12 27
rect 14 7 17 27
rect 19 7 20 27
rect 26 7 27 17
rect 29 7 30 17
<< pdiffusion >>
rect 8 87 9 123
rect 2 83 9 87
rect 11 89 12 123
rect 18 89 19 123
rect 11 83 19 89
rect 21 83 22 123
rect 28 83 29 123
rect 31 83 32 123
<< ndcontact >>
rect 5 7 11 27
rect 20 7 26 27
rect 30 7 36 17
<< pdcontact >>
rect 2 87 8 123
rect 12 89 18 123
rect 22 83 28 123
rect 32 83 38 123
<< psubstratepcontact >>
rect -3 -3 43 3
<< nsubstratencontact >>
rect -3 127 43 133
<< polysilicon >>
rect 9 123 11 125
rect 19 123 21 125
rect 29 123 31 125
rect 9 76 11 83
rect 19 76 21 83
rect 5 73 11 76
rect 15 73 21 76
rect 5 51 8 73
rect 15 64 18 73
rect 5 30 8 45
rect 15 41 18 58
rect 29 51 31 83
rect 15 36 19 41
rect 5 28 14 30
rect 12 27 14 28
rect 17 27 19 36
rect 28 32 31 51
rect 27 29 31 32
rect 27 17 29 29
rect 12 5 14 7
rect 17 5 19 7
rect 27 5 29 7
<< polycontact >>
rect 12 58 18 64
rect 2 45 8 51
rect 22 45 28 51
<< metal1 >>
rect -3 133 43 134
rect -3 126 43 127
rect 12 123 18 126
rect 2 86 8 87
rect 2 83 22 86
rect 34 58 37 83
rect 34 27 37 51
rect 26 23 37 27
rect 5 4 11 7
rect 30 4 36 7
rect -3 3 43 4
rect -3 -4 43 -3
<< m2contact >>
rect 1 51 8 58
rect 11 51 18 58
rect 21 51 28 58
rect 31 51 38 58
<< metal2 >>
rect 3 58 7 67
rect 23 58 27 67
rect 13 43 17 51
rect 33 43 37 51
<< m1p >>
rect -3 126 43 134
rect -3 -4 43 4
<< m2p >>
rect 3 59 7 67
rect 23 59 27 67
rect 13 43 17 50
rect 33 43 37 50
<< labels >>
rlabel metal2 15 45 15 45 1 B
port 2 n signal input
rlabel metal2 25 65 25 65 1 C
port 3 n signal input
rlabel metal2 35 44 35 44 1 Y
port 4 n signal output
rlabel metal1 -3 126 43 134 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -3 -4 43 4 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal2 5 65 5 65 1 A
port 1 n signal input
<< properties >>
string FIXED_BBOX 0 0 40 130
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
