magic
tech scmos
magscale 1 2
timestamp 1727732147
<< nwell >>
rect -12 134 212 252
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 60 14 64 54
rect 80 14 84 54
rect 100 14 104 54
rect 120 14 124 54
rect 140 14 144 54
rect 160 14 164 54
<< ptransistor >>
rect 20 146 24 226
rect 40 146 44 226
rect 60 146 64 226
rect 80 146 84 226
rect 100 146 104 226
rect 120 146 124 226
rect 140 146 144 226
rect 160 146 164 226
<< ndiffusion >>
rect 18 14 20 54
rect 24 14 26 54
rect 38 14 40 54
rect 44 14 46 54
rect 58 14 60 54
rect 64 14 66 54
rect 78 14 80 54
rect 84 14 86 54
rect 98 14 100 54
rect 104 14 106 54
rect 118 14 120 54
rect 124 14 126 54
rect 138 14 140 54
rect 144 14 146 54
rect 158 14 160 54
rect 164 14 166 54
<< pdiffusion >>
rect 18 146 20 226
rect 24 146 26 226
rect 38 146 40 226
rect 44 146 46 226
rect 58 146 60 226
rect 64 146 66 226
rect 78 146 80 226
rect 84 146 86 226
rect 98 146 100 226
rect 104 146 106 226
rect 118 146 120 226
rect 124 146 126 226
rect 138 146 140 226
rect 144 146 146 226
rect 158 146 160 226
rect 164 146 166 226
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 54
rect 46 14 58 54
rect 66 14 78 54
rect 86 14 98 54
rect 106 14 118 54
rect 126 14 138 54
rect 146 14 158 54
rect 166 14 178 54
<< pdcontact >>
rect 6 146 18 226
rect 26 146 38 226
rect 46 146 58 226
rect 66 146 78 226
rect 86 146 98 226
rect 106 146 118 226
rect 126 146 138 226
rect 146 146 158 226
rect 166 146 178 226
<< psubstratepcontact >>
rect -6 -6 206 6
<< nsubstratencontact >>
rect -6 234 206 246
<< polysilicon >>
rect 20 226 24 230
rect 40 226 44 230
rect 60 226 64 230
rect 80 226 84 230
rect 100 226 104 230
rect 120 226 124 230
rect 140 226 144 230
rect 160 226 164 230
rect 20 54 24 146
rect 40 103 44 146
rect 36 91 44 103
rect 40 54 44 91
rect 60 86 64 146
rect 80 86 84 146
rect 72 74 84 86
rect 60 54 64 74
rect 80 54 84 74
rect 100 86 104 146
rect 120 86 124 146
rect 112 74 124 86
rect 100 54 104 74
rect 120 54 124 74
rect 140 86 144 146
rect 160 86 164 146
rect 152 74 164 86
rect 140 54 144 74
rect 160 54 164 74
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
rect 80 10 84 14
rect 100 10 104 14
rect 120 10 124 14
rect 140 10 144 14
rect 160 10 164 14
<< polycontact >>
rect 24 91 36 103
rect 60 74 72 86
rect 100 74 112 86
rect 140 74 152 86
<< metal1 >>
rect -6 246 206 248
rect -6 232 206 234
rect 6 226 18 232
rect 46 226 58 232
rect 86 226 98 232
rect 126 226 138 232
rect 166 226 178 232
rect 26 140 38 146
rect 66 140 78 146
rect 106 140 118 146
rect 146 140 158 146
rect 26 132 52 140
rect 66 132 92 140
rect 106 132 132 140
rect 146 132 164 140
rect 23 103 37 117
rect 44 82 52 132
rect 44 74 60 82
rect 84 82 92 132
rect 84 74 100 82
rect 124 82 132 132
rect 158 117 164 132
rect 158 103 177 117
rect 124 74 140 82
rect 44 68 52 74
rect 84 68 92 74
rect 124 68 132 74
rect 158 68 164 103
rect 26 60 52 68
rect 66 60 92 68
rect 106 60 132 68
rect 146 60 164 68
rect 26 54 38 60
rect 66 54 78 60
rect 106 54 118 60
rect 146 54 158 60
rect 6 8 18 14
rect 46 8 58 14
rect 86 8 98 14
rect 126 8 138 14
rect 166 8 178 14
rect -6 6 206 8
rect -6 -8 206 -6
<< m1p >>
rect 23 103 37 117
rect 163 103 177 117
<< labels >>
rlabel metal1 23 103 37 117 0 A
port 0 nsew signal input
rlabel metal1 163 103 177 117 0 Y
port 1 nsew signal output
rlabel metal1 -6 -8 206 8 0 gnd
port 3 nsew ground bidirectional abutment
rlabel metal1 -6 232 206 248 0 vdd
port 2 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 200 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
