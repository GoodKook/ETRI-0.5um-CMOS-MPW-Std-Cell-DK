magic
tech scmos
magscale 1 2
timestamp 1740356047
<< metal1 >>
rect -62 5762 30 5778
rect -62 5298 -2 5762
rect 5822 5538 5882 5778
rect 5790 5522 5882 5538
rect 5697 5457 5713 5463
rect 1127 5397 1193 5403
rect 5697 5383 5703 5457
rect 5697 5377 5713 5383
rect -62 5282 30 5298
rect -62 4818 -2 5282
rect 3967 5197 3983 5203
rect 3977 5143 3983 5197
rect 3977 5137 4013 5143
rect 5757 5127 5763 5193
rect 1587 5097 1613 5103
rect 5822 5058 5882 5522
rect 5790 5042 5882 5058
rect 5577 4977 5593 4983
rect 4127 4957 4173 4963
rect 2807 4897 2833 4903
rect 5557 4903 5563 4973
rect 5547 4897 5563 4903
rect 5577 4903 5583 4977
rect 5577 4897 5603 4903
rect 5597 4887 5603 4897
rect -62 4802 30 4818
rect -62 4338 -2 4802
rect 5327 4717 5343 4723
rect 5337 4703 5343 4717
rect 5387 4717 5403 4723
rect 3807 4697 3823 4703
rect 5337 4697 5373 4703
rect 3817 4663 3823 4697
rect 3817 4657 3853 4663
rect 5397 4643 5403 4717
rect 5507 4717 5533 4723
rect 5607 4717 5653 4723
rect 5397 4637 5413 4643
rect 5822 4578 5882 5042
rect 5790 4562 5882 4578
rect 167 4517 193 4523
rect 1967 4497 2013 4503
rect 287 4477 313 4483
rect -62 4322 30 4338
rect -62 3858 -2 4322
rect 5067 4217 5133 4223
rect 507 4137 533 4143
rect 5822 4098 5882 4562
rect 5790 4082 5882 4098
rect 1667 4037 1693 4043
rect 2607 4017 2623 4023
rect 107 3937 133 3943
rect 157 3923 163 4013
rect 2617 3967 2623 4017
rect 2637 3943 2643 3973
rect 2607 3937 2643 3943
rect 107 3917 163 3923
rect -62 3842 30 3858
rect -62 3378 -2 3842
rect 3367 3777 3393 3783
rect 3087 3757 3193 3763
rect 1367 3737 1413 3743
rect 4847 3737 4873 3743
rect 5822 3618 5882 4082
rect 5790 3602 5882 3618
rect 2167 3537 2193 3543
rect 4347 3537 4393 3543
rect 57 3517 73 3523
rect 57 3443 63 3517
rect 3407 3517 3433 3523
rect 1217 3463 1223 3513
rect 1217 3457 1253 3463
rect 57 3437 73 3443
rect -62 3362 30 3378
rect -62 2898 -2 3362
rect 1867 3297 1893 3303
rect 107 3257 123 3263
rect 117 3183 123 3257
rect 2807 3217 2833 3223
rect 2947 3217 2973 3223
rect 107 3177 123 3183
rect 2887 3177 2933 3183
rect 5822 3138 5882 3602
rect 5790 3122 5882 3138
rect 987 3037 1013 3043
rect 2547 2997 2593 3003
rect 3127 2977 3153 2983
rect -62 2882 30 2898
rect -62 2418 -2 2882
rect 3207 2797 3233 2803
rect 2407 2717 2453 2723
rect 1607 2697 1633 2703
rect 5822 2658 5882 3122
rect 5790 2642 5882 2658
rect 1797 2503 1803 2553
rect 2817 2527 2823 2593
rect 3187 2577 3213 2583
rect 3717 2577 3733 2583
rect 3127 2557 3143 2563
rect 3137 2543 3143 2557
rect 3717 2547 3723 2577
rect 3137 2537 3193 2543
rect 1797 2497 1843 2503
rect 1767 2477 1813 2483
rect 1837 2463 1843 2497
rect 1827 2457 1843 2463
rect -62 2402 30 2418
rect -62 1938 -2 2402
rect 3467 2377 3513 2383
rect 5167 2317 5193 2323
rect 3377 2303 3383 2313
rect 3307 2297 3383 2303
rect 5267 2297 5313 2303
rect 3257 2243 3263 2293
rect 3227 2237 3263 2243
rect 5822 2178 5882 2642
rect 5790 2162 5882 2178
rect 287 2077 333 2083
rect 857 2043 863 2073
rect 827 2037 863 2043
rect 3727 2037 3773 2043
rect 2927 1997 2993 2003
rect -62 1922 30 1938
rect -62 1458 -2 1922
rect 4357 1837 4373 1843
rect 737 1817 793 1823
rect 737 1763 743 1817
rect 4357 1823 4363 1837
rect 4337 1817 4363 1823
rect 707 1757 743 1763
rect 3917 1763 3923 1813
rect 3887 1757 3923 1763
rect 4337 1727 4343 1817
rect 5357 1743 5363 1833
rect 5327 1737 5363 1743
rect 5822 1698 5882 2162
rect 5790 1682 5882 1698
rect 5227 1637 5253 1643
rect 4507 1617 4563 1623
rect 2787 1597 2833 1603
rect 4557 1567 4563 1617
rect 5257 1617 5273 1623
rect 5137 1597 5153 1603
rect 5137 1523 5143 1597
rect 5257 1527 5263 1617
rect 5517 1617 5533 1623
rect 5517 1543 5523 1617
rect 5507 1537 5523 1543
rect 5137 1517 5153 1523
rect -62 1442 30 1458
rect -62 978 -2 1442
rect 2857 1283 2863 1373
rect 3667 1337 3713 1343
rect 2847 1277 2863 1283
rect 5822 1218 5882 1682
rect 5790 1202 5882 1218
rect 1827 1117 1853 1123
rect 1127 1077 1153 1083
rect 3797 1067 3803 1133
rect 5687 1117 5703 1123
rect 5697 1087 5703 1117
rect 4647 1077 4713 1083
rect -62 962 30 978
rect -62 498 -2 962
rect 1607 877 1653 883
rect 3817 877 3853 883
rect 1147 797 1173 803
rect 3817 783 3823 877
rect 5047 857 5093 863
rect 3807 777 3823 783
rect 5822 738 5882 1202
rect 5790 722 5882 738
rect 3857 657 3873 663
rect 3287 637 3313 643
rect 3707 637 3733 643
rect 3857 627 3863 657
rect -62 482 30 498
rect -62 18 -2 482
rect 3167 377 3293 383
rect 1427 337 1473 343
rect 5822 258 5882 722
rect 5790 242 5882 258
rect 4587 157 4613 163
rect 2987 97 3033 103
rect -62 2 30 18
rect 5822 2 5882 242
<< m2contact >>
rect 1113 5393 1127 5407
rect 1193 5393 1207 5407
rect 5713 5453 5727 5467
rect 5713 5373 5727 5387
rect 3953 5193 3967 5207
rect 5753 5193 5767 5207
rect 4013 5133 4027 5147
rect 5753 5113 5767 5127
rect 1573 5093 1587 5107
rect 1613 5093 1627 5107
rect 5553 4973 5567 4987
rect 4113 4953 4127 4967
rect 4173 4953 4187 4967
rect 2793 4893 2807 4907
rect 2833 4893 2847 4907
rect 5533 4893 5547 4907
rect 5593 4973 5607 4987
rect 5593 4873 5607 4887
rect 5313 4713 5327 4727
rect 3793 4693 3807 4707
rect 5373 4713 5387 4727
rect 5373 4693 5387 4707
rect 3853 4653 3867 4667
rect 5493 4713 5507 4727
rect 5533 4713 5547 4727
rect 5593 4713 5607 4727
rect 5653 4713 5667 4727
rect 5413 4633 5427 4647
rect 153 4513 167 4527
rect 193 4513 207 4527
rect 1953 4493 1967 4507
rect 2013 4493 2027 4507
rect 273 4473 287 4487
rect 313 4473 327 4487
rect 5053 4213 5067 4227
rect 5133 4213 5147 4227
rect 493 4133 507 4147
rect 533 4133 547 4147
rect 1653 4033 1667 4047
rect 1693 4033 1707 4047
rect 153 4013 167 4027
rect 2593 4013 2607 4027
rect 93 3933 107 3947
rect 133 3933 147 3947
rect 93 3913 107 3927
rect 2633 3973 2647 3987
rect 2613 3953 2627 3967
rect 2593 3933 2607 3947
rect 3353 3773 3367 3787
rect 3393 3773 3407 3787
rect 3073 3753 3087 3767
rect 3193 3753 3207 3767
rect 1353 3733 1367 3747
rect 1413 3733 1427 3747
rect 4833 3733 4847 3747
rect 4873 3733 4887 3747
rect 2153 3533 2167 3547
rect 2193 3533 2207 3547
rect 4333 3533 4347 3547
rect 4393 3533 4407 3547
rect 73 3513 87 3527
rect 1213 3513 1227 3527
rect 3393 3513 3407 3527
rect 3433 3513 3447 3527
rect 1253 3453 1267 3467
rect 73 3433 87 3447
rect 1853 3293 1867 3307
rect 1893 3293 1907 3307
rect 93 3253 107 3267
rect 93 3173 107 3187
rect 2793 3213 2807 3227
rect 2833 3213 2847 3227
rect 2933 3213 2947 3227
rect 2973 3213 2987 3227
rect 2873 3173 2887 3187
rect 2933 3173 2947 3187
rect 973 3033 987 3047
rect 1013 3033 1027 3047
rect 2533 2993 2547 3007
rect 2593 2993 2607 3007
rect 3113 2973 3127 2987
rect 3153 2973 3167 2987
rect 4373 2873 4387 2887
rect 3193 2793 3207 2807
rect 3233 2793 3247 2807
rect 2393 2713 2407 2727
rect 2453 2713 2467 2727
rect 1593 2693 1607 2707
rect 1633 2693 1647 2707
rect 2813 2593 2827 2607
rect 1793 2553 1807 2567
rect 3173 2573 3187 2587
rect 3213 2573 3227 2587
rect 3113 2553 3127 2567
rect 3733 2573 3747 2587
rect 3193 2533 3207 2547
rect 3713 2533 3727 2547
rect 2813 2513 2827 2527
rect 1753 2473 1767 2487
rect 1813 2473 1827 2487
rect 1813 2453 1827 2467
rect 2533 2393 2547 2407
rect 4353 2393 4367 2407
rect 4493 2393 4507 2407
rect 3453 2373 3467 2387
rect 3513 2373 3527 2387
rect 3373 2313 3387 2327
rect 5153 2313 5167 2327
rect 5193 2313 5207 2327
rect 3253 2293 3267 2307
rect 3293 2293 3307 2307
rect 5253 2293 5267 2307
rect 5313 2293 5327 2307
rect 3213 2233 3227 2247
rect 273 2073 287 2087
rect 333 2073 347 2087
rect 853 2073 867 2087
rect 813 2033 827 2047
rect 3713 2033 3727 2047
rect 3773 2033 3787 2047
rect 2913 1993 2927 2007
rect 2993 1993 3007 2007
rect 2653 1913 2667 1927
rect 2773 1913 2787 1927
rect 693 1753 707 1767
rect 793 1813 807 1827
rect 3913 1813 3927 1827
rect 4373 1833 4387 1847
rect 5353 1833 5367 1847
rect 3873 1753 3887 1767
rect 5313 1733 5327 1747
rect 4333 1713 4347 1727
rect 5213 1633 5227 1647
rect 5253 1633 5267 1647
rect 4493 1613 4507 1627
rect 2773 1593 2787 1607
rect 2833 1593 2847 1607
rect 4553 1553 4567 1567
rect 5153 1593 5167 1607
rect 5273 1613 5287 1627
rect 5493 1533 5507 1547
rect 5533 1613 5547 1627
rect 5153 1513 5167 1527
rect 5253 1513 5267 1527
rect 2133 1433 2147 1447
rect 3233 1433 3247 1447
rect 2853 1373 2867 1387
rect 2833 1273 2847 1287
rect 3653 1333 3667 1347
rect 3713 1333 3727 1347
rect 3793 1133 3807 1147
rect 1813 1113 1827 1127
rect 1853 1113 1867 1127
rect 1113 1073 1127 1087
rect 1153 1073 1167 1087
rect 5673 1113 5687 1127
rect 4633 1073 4647 1087
rect 4713 1073 4727 1087
rect 5693 1073 5707 1087
rect 3793 1053 3807 1067
rect 1593 873 1607 887
rect 1653 873 1667 887
rect 1133 793 1147 807
rect 1173 793 1187 807
rect 3793 773 3807 787
rect 3853 873 3867 887
rect 5033 853 5047 867
rect 5093 853 5107 867
rect 3273 633 3287 647
rect 3313 633 3327 647
rect 3693 633 3707 647
rect 3733 633 3747 647
rect 3873 653 3887 667
rect 3853 613 3867 627
rect 3153 373 3167 387
rect 3293 373 3307 387
rect 1413 333 1427 347
rect 1473 333 1487 347
rect 4573 153 4587 167
rect 4613 153 4627 167
rect 2973 93 2987 107
rect 3033 93 3047 107
<< metal2 >>
rect 4716 5667 4723 5823
rect 5196 5816 5223 5823
rect 556 5656 583 5663
rect 76 5467 83 5643
rect 96 5487 103 5623
rect 136 5436 143 5453
rect 196 5427 203 5613
rect 236 5443 243 5623
rect 256 5547 263 5643
rect 456 5643 463 5653
rect 436 5636 463 5643
rect 236 5436 263 5443
rect 56 5416 83 5423
rect 56 5387 63 5416
rect 256 5416 263 5436
rect 36 4787 43 5013
rect 36 4187 43 4673
rect 56 4507 63 5313
rect 76 5176 83 5373
rect 96 5327 103 5393
rect 156 5187 163 5213
rect 116 5167 123 5183
rect 116 4983 123 5153
rect 136 5127 143 5163
rect 96 4976 123 4983
rect 76 4936 83 4973
rect 96 4956 103 4976
rect 136 4956 163 4963
rect 116 4887 123 4943
rect 96 4676 103 4753
rect 116 4707 123 4773
rect 136 4676 143 4833
rect 156 4767 163 4956
rect 176 4803 183 5233
rect 196 5187 203 5413
rect 236 5247 243 5403
rect 276 5396 283 5433
rect 296 5416 323 5423
rect 396 5416 403 5473
rect 236 5156 243 5213
rect 316 5187 323 5416
rect 276 5143 283 5173
rect 256 5136 283 5143
rect 316 5123 323 5173
rect 356 5167 363 5393
rect 316 5116 343 5123
rect 216 4967 223 5113
rect 376 5027 383 5403
rect 456 5367 463 5636
rect 496 5607 503 5643
rect 536 5607 543 5633
rect 496 5443 503 5593
rect 576 5487 583 5656
rect 776 5656 803 5663
rect 656 5567 663 5643
rect 476 5436 503 5443
rect 276 4936 293 4943
rect 376 4936 383 4973
rect 396 4967 403 5333
rect 416 5147 423 5353
rect 476 5347 483 5436
rect 536 5416 543 5473
rect 576 5416 583 5453
rect 496 5367 503 5413
rect 196 4847 203 4933
rect 296 4907 303 4933
rect 176 4796 203 4803
rect 76 4483 83 4663
rect 56 4476 83 4483
rect 96 4476 103 4493
rect 136 4476 143 4573
rect 156 4527 163 4713
rect 56 4127 63 4476
rect 156 4423 163 4493
rect 176 4447 183 4773
rect 196 4727 203 4796
rect 216 4703 223 4893
rect 196 4696 223 4703
rect 196 4647 203 4696
rect 236 4647 243 4673
rect 256 4627 263 4703
rect 156 4416 183 4423
rect 56 3983 63 4093
rect 76 4027 83 4413
rect 96 4107 103 4203
rect 176 4187 183 4416
rect 56 3976 83 3983
rect 96 3947 103 3973
rect 16 3027 23 3133
rect 16 1507 23 1553
rect 36 1147 43 1573
rect 36 607 43 1133
rect 56 627 63 3773
rect 96 3763 103 3913
rect 116 3787 123 4113
rect 136 3967 143 4153
rect 156 4087 163 4183
rect 156 4027 163 4033
rect 176 4027 183 4153
rect 196 4047 203 4513
rect 236 4456 243 4553
rect 256 4447 263 4493
rect 276 4487 283 4653
rect 296 4487 303 4873
rect 316 4787 323 4913
rect 416 4783 423 4973
rect 396 4776 423 4783
rect 376 4687 383 4713
rect 396 4707 403 4776
rect 316 4676 343 4683
rect 316 4647 323 4676
rect 416 4663 423 4753
rect 396 4656 423 4663
rect 356 4627 363 4633
rect 216 4147 223 4193
rect 236 4167 243 4203
rect 176 3996 183 4013
rect 76 3756 103 3763
rect 76 3747 83 3756
rect 116 3736 123 3753
rect 76 3527 83 3693
rect 96 3607 103 3723
rect 136 3707 143 3933
rect 96 3516 103 3573
rect 136 3527 143 3553
rect 87 3436 93 3443
rect 76 3236 83 3253
rect 96 3247 103 3253
rect 116 3187 123 3433
rect 136 3227 143 3453
rect 76 2987 83 3173
rect 96 3036 103 3173
rect 156 3063 163 3993
rect 236 3976 243 4113
rect 256 3987 263 4133
rect 296 4087 303 4183
rect 296 4047 303 4073
rect 176 3467 183 3953
rect 316 3747 323 4473
rect 416 4467 423 4553
rect 336 4447 343 4453
rect 336 4187 343 4413
rect 356 4016 363 4053
rect 216 3707 223 3723
rect 256 3707 263 3723
rect 216 3547 223 3593
rect 296 3587 303 3713
rect 276 3507 283 3573
rect 136 3056 163 3063
rect 76 2776 83 2793
rect 116 2787 123 2973
rect 96 2576 103 2733
rect 76 2307 83 2543
rect 116 2527 123 2733
rect 76 1816 83 2113
rect 96 2076 103 2273
rect 116 2167 123 2263
rect 136 2103 143 3056
rect 176 3003 183 3213
rect 156 2996 183 3003
rect 156 2747 163 2996
rect 196 2756 203 3223
rect 256 3207 263 3273
rect 276 3227 283 3253
rect 216 3016 243 3023
rect 216 3007 223 3016
rect 256 3007 263 3033
rect 276 3016 283 3213
rect 296 3047 303 3513
rect 316 3287 323 3733
rect 336 3716 363 3723
rect 336 3707 343 3716
rect 376 3703 383 4253
rect 396 4216 403 4433
rect 436 4267 443 5153
rect 496 5107 503 5173
rect 536 5163 543 5193
rect 516 5156 543 5163
rect 456 4956 483 4963
rect 516 4956 523 5133
rect 536 5127 543 5156
rect 596 5163 603 5413
rect 616 5227 623 5433
rect 656 5416 663 5533
rect 676 5427 683 5623
rect 716 5587 723 5623
rect 696 5416 703 5473
rect 736 5427 743 5633
rect 776 5627 783 5656
rect 1376 5656 1403 5663
rect 776 5467 783 5613
rect 816 5567 823 5643
rect 976 5636 1003 5643
rect 896 5587 903 5633
rect 916 5607 923 5623
rect 996 5607 1003 5636
rect 796 5436 803 5553
rect 956 5447 963 5603
rect 1056 5547 1063 5623
rect 1096 5603 1103 5623
rect 1096 5596 1123 5603
rect 716 5367 723 5403
rect 587 5156 603 5163
rect 616 5156 623 5173
rect 796 5156 803 5173
rect 816 5147 823 5413
rect 876 5167 883 5183
rect 916 5176 923 5413
rect 956 5396 963 5433
rect 1076 5427 1083 5593
rect 1116 5587 1123 5596
rect 1096 5436 1103 5573
rect 1116 5407 1123 5423
rect 996 5207 1003 5403
rect 856 5147 863 5163
rect 636 4967 643 5143
rect 856 5127 863 5133
rect 456 4767 463 4956
rect 496 4887 503 4943
rect 536 4936 553 4943
rect 556 4847 563 4933
rect 456 4696 483 4703
rect 456 4667 463 4696
rect 456 4447 463 4633
rect 496 4587 503 4673
rect 416 4127 423 4203
rect 436 4107 443 4223
rect 496 4147 503 4533
rect 516 4456 523 4593
rect 536 4476 543 4653
rect 576 4547 583 4953
rect 636 4907 643 4923
rect 576 4476 583 4513
rect 596 4487 603 4893
rect 656 4687 663 4703
rect 636 4547 643 4683
rect 656 4456 663 4533
rect 676 4507 683 4683
rect 696 4567 703 4953
rect 716 4487 723 4513
rect 536 4216 543 4433
rect 416 3983 423 4053
rect 456 4016 463 4093
rect 496 3996 523 4003
rect 416 3976 443 3983
rect 376 3696 403 3703
rect 336 3536 343 3693
rect 376 3547 383 3553
rect 376 3503 383 3533
rect 396 3507 403 3696
rect 356 3496 383 3503
rect 416 3307 423 3573
rect 436 3516 443 3693
rect 496 3567 503 3713
rect 496 3496 503 3553
rect 516 3463 523 3996
rect 536 3707 543 4133
rect 556 4127 563 4203
rect 576 4167 583 4223
rect 736 4207 743 5093
rect 756 4936 763 5093
rect 776 4696 783 4913
rect 816 4507 823 4703
rect 836 4607 843 4683
rect 876 4667 883 5153
rect 896 4967 903 5113
rect 916 4956 923 5133
rect 1036 5107 1043 5163
rect 1056 4983 1063 5173
rect 1116 5087 1123 5393
rect 1156 5387 1163 5413
rect 1176 5407 1183 5453
rect 1196 5416 1223 5423
rect 1196 5407 1203 5416
rect 1296 5403 1303 5433
rect 1276 5396 1303 5403
rect 1176 5383 1183 5393
rect 1176 5376 1203 5383
rect 1167 5156 1183 5163
rect 1056 4976 1083 4983
rect 956 4956 963 4973
rect 896 4936 903 4953
rect 996 4947 1003 4973
rect 1016 4956 1043 4963
rect 1016 4727 1023 4956
rect 1116 4943 1123 4953
rect 1096 4936 1123 4943
rect 916 4676 943 4683
rect 896 4607 903 4643
rect 936 4547 943 4676
rect 1056 4647 1063 4933
rect 996 4567 1003 4643
rect 856 4463 863 4533
rect 896 4507 903 4513
rect 996 4467 1003 4553
rect 1056 4496 1083 4503
rect 856 4456 883 4463
rect 656 4196 683 4203
rect 576 4147 583 4153
rect 596 4067 603 4193
rect 656 4127 663 4196
rect 556 3987 563 4033
rect 616 4016 623 4033
rect 636 3996 643 4093
rect 716 4007 723 4183
rect 736 4107 743 4163
rect 756 4016 763 4193
rect 816 3996 823 4153
rect 876 4047 883 4183
rect 716 3967 723 3993
rect 876 3976 883 4033
rect 676 3736 703 3743
rect 556 3707 563 3723
rect 576 3667 583 3703
rect 616 3687 623 3703
rect 556 3496 583 3503
rect 556 3487 563 3496
rect 596 3476 603 3513
rect 616 3496 623 3533
rect 496 3456 523 3463
rect 316 3247 323 3253
rect 356 3203 363 3293
rect 396 3256 403 3273
rect 436 3256 463 3263
rect 456 3227 463 3256
rect 336 3196 363 3203
rect 356 3067 363 3196
rect 396 3087 403 3213
rect 396 3016 403 3073
rect 316 3003 323 3013
rect 296 2996 323 3003
rect 216 2987 223 2993
rect 376 2987 383 3003
rect 176 2667 183 2743
rect 156 2576 163 2593
rect 156 2267 163 2433
rect 136 2096 163 2103
rect 116 2076 143 2083
rect 116 2007 123 2076
rect 116 1767 123 1813
rect 136 1787 143 1803
rect 136 1707 143 1773
rect 76 1576 83 1633
rect 76 1336 83 1513
rect 116 1427 123 1533
rect 116 1247 123 1343
rect 136 1227 143 1323
rect 96 1136 103 1173
rect 156 1143 163 2096
rect 176 1267 183 2513
rect 196 2296 203 2713
rect 236 2587 243 2763
rect 256 2447 263 2793
rect 376 2787 383 2973
rect 416 2863 423 2993
rect 476 2907 483 3033
rect 496 2883 503 3456
rect 556 3447 563 3473
rect 556 3236 563 3253
rect 516 3196 543 3203
rect 516 3027 523 3196
rect 576 3127 583 3223
rect 576 3036 583 3053
rect 596 2947 603 3433
rect 636 3187 643 3483
rect 656 3307 663 3733
rect 676 3587 683 3736
rect 716 3707 723 3723
rect 896 3707 903 4293
rect 956 4196 983 4203
rect 916 4167 923 4193
rect 956 4016 963 4033
rect 976 4027 983 4196
rect 776 3696 803 3703
rect 716 3647 723 3693
rect 676 3223 683 3293
rect 656 3216 683 3223
rect 636 3036 643 3053
rect 676 3036 683 3053
rect 496 2876 523 2883
rect 396 2856 423 2863
rect 356 2667 363 2723
rect 276 2556 283 2653
rect 376 2607 383 2773
rect 396 2727 403 2856
rect 496 2747 503 2813
rect 476 2727 483 2743
rect 436 2707 443 2723
rect 316 2576 363 2583
rect 356 2527 363 2576
rect 396 2536 403 2553
rect 236 2263 243 2293
rect 256 2267 263 2283
rect 216 2256 243 2263
rect 196 2047 203 2093
rect 216 2023 223 2256
rect 276 2107 283 2513
rect 296 2267 303 2313
rect 356 2296 363 2313
rect 276 2036 283 2073
rect 296 2067 303 2093
rect 216 2016 243 2023
rect 196 1807 203 1833
rect 216 1827 223 1853
rect 236 1827 243 2016
rect 196 1547 203 1673
rect 216 1567 223 1733
rect 256 1727 263 1783
rect 276 1607 283 1953
rect 296 1687 303 2013
rect 316 1783 323 2253
rect 376 2247 383 2533
rect 476 2523 483 2573
rect 456 2516 483 2523
rect 336 2087 343 2193
rect 416 2187 423 2273
rect 336 1967 343 2073
rect 356 2027 363 2063
rect 336 1803 343 1833
rect 376 1827 383 1933
rect 336 1796 363 1803
rect 396 1796 403 1873
rect 416 1827 423 2013
rect 316 1776 343 1783
rect 316 1583 323 1613
rect 296 1576 323 1583
rect 236 1547 243 1563
rect 276 1556 283 1573
rect 196 1327 203 1333
rect 216 1227 223 1283
rect 136 1136 163 1143
rect 76 856 83 1073
rect 136 887 143 1136
rect 216 1116 223 1153
rect 116 807 123 863
rect 136 727 143 833
rect 116 596 123 633
rect 156 623 163 653
rect 136 616 163 623
rect 156 587 163 616
rect 76 376 83 573
rect 116 347 123 383
rect 156 363 163 533
rect 136 356 163 363
rect 96 136 103 153
rect 116 147 123 333
rect 156 127 163 173
rect 176 167 183 873
rect 236 867 243 1253
rect 276 1247 283 1313
rect 296 1167 303 1473
rect 316 1467 323 1576
rect 316 1267 323 1413
rect 276 1116 303 1123
rect 336 1116 343 1776
rect 356 1727 363 1773
rect 416 1767 423 1783
rect 416 1596 423 1733
rect 356 1547 363 1573
rect 376 1527 383 1573
rect 396 1567 403 1583
rect 396 1487 403 1553
rect 356 1336 363 1453
rect 396 1327 403 1343
rect 376 1287 383 1323
rect 276 1107 283 1116
rect 236 836 243 853
rect 276 807 283 1093
rect 316 1087 323 1103
rect 356 1096 363 1113
rect 376 1107 383 1253
rect 396 1127 403 1313
rect 316 827 323 1073
rect 396 1027 403 1113
rect 416 1027 423 1323
rect 436 1307 443 2253
rect 476 2247 483 2263
rect 496 2247 503 2283
rect 516 2227 523 2876
rect 616 2803 623 3033
rect 736 3027 743 3693
rect 776 3687 783 3696
rect 776 3496 783 3673
rect 896 3496 903 3573
rect 916 3527 923 3993
rect 976 3967 983 3983
rect 1016 3767 1023 4473
rect 1076 4447 1083 4496
rect 1096 4427 1103 4873
rect 1136 4683 1143 5093
rect 1156 4903 1163 5073
rect 1176 4967 1183 5156
rect 1196 4956 1203 5376
rect 1256 5176 1263 5373
rect 1276 5107 1283 5163
rect 1296 4987 1303 5173
rect 1316 5127 1323 5163
rect 1336 5147 1343 5653
rect 1396 5627 1403 5656
rect 1356 5587 1363 5623
rect 1376 5507 1383 5613
rect 1416 5607 1423 5623
rect 1536 5607 1543 5663
rect 1776 5656 1803 5663
rect 1556 5627 1563 5643
rect 1376 5436 1383 5493
rect 1396 5456 1403 5533
rect 1416 5447 1423 5593
rect 1636 5487 1643 5653
rect 1716 5636 1743 5643
rect 1736 5627 1743 5636
rect 1356 5167 1363 5433
rect 1516 5183 1523 5403
rect 1556 5396 1563 5433
rect 1596 5423 1603 5433
rect 1576 5416 1603 5423
rect 1496 5176 1523 5183
rect 1236 4956 1243 4973
rect 1176 4936 1183 4953
rect 1156 4896 1183 4903
rect 1116 4676 1143 4683
rect 1156 4467 1163 4673
rect 1176 4507 1183 4896
rect 1296 4787 1303 4973
rect 1356 4747 1363 5113
rect 1416 5027 1423 5153
rect 1396 4723 1403 4933
rect 1416 4907 1423 4923
rect 1476 4887 1483 5143
rect 1496 4927 1503 5176
rect 1396 4716 1423 4723
rect 1036 3983 1043 4213
rect 1136 4207 1143 4443
rect 1176 4436 1183 4473
rect 1116 4196 1133 4203
rect 1056 4167 1063 4183
rect 1096 4127 1103 4163
rect 1036 3976 1063 3983
rect 1096 3976 1103 4013
rect 956 3547 963 3753
rect 996 3716 1003 3733
rect 1036 3716 1043 3793
rect 976 3587 983 3703
rect 1076 3703 1083 3813
rect 1056 3696 1083 3703
rect 1096 3687 1103 3853
rect 1116 3767 1123 3963
rect 1156 3947 1163 4413
rect 1216 4243 1223 4633
rect 1256 4267 1263 4633
rect 1276 4547 1283 4663
rect 1336 4643 1343 4663
rect 1376 4647 1383 4663
rect 1336 4636 1363 4643
rect 1316 4507 1323 4613
rect 1276 4476 1283 4493
rect 1296 4447 1303 4463
rect 1356 4447 1363 4636
rect 1356 4367 1363 4433
rect 1196 4236 1223 4243
rect 1176 4003 1183 4233
rect 1196 4167 1203 4236
rect 1296 4227 1303 4253
rect 1256 4127 1263 4213
rect 1276 4196 1303 4203
rect 1276 4187 1283 4196
rect 1176 3996 1203 4003
rect 1236 3996 1243 4073
rect 1276 3996 1283 4013
rect 1176 3827 1183 3996
rect 1216 3967 1223 3983
rect 1216 3807 1223 3953
rect 1256 3867 1263 3983
rect 1296 3907 1303 4196
rect 1316 3967 1323 4253
rect 1376 4247 1383 4573
rect 1396 4547 1403 4683
rect 1416 4503 1423 4716
rect 1436 4587 1443 4713
rect 1516 4647 1523 5153
rect 1536 5147 1543 5373
rect 1596 5287 1603 5416
rect 1556 5156 1563 5273
rect 1616 5163 1623 5473
rect 1656 5467 1663 5623
rect 1696 5416 1703 5473
rect 1736 5467 1743 5613
rect 1596 5156 1623 5163
rect 1576 5107 1583 5123
rect 1576 4936 1583 4973
rect 1536 4687 1543 4913
rect 1556 4907 1563 4923
rect 1596 4916 1603 5156
rect 1696 5156 1703 5173
rect 1756 5167 1763 5633
rect 1776 5607 1783 5656
rect 1816 5567 1823 5643
rect 1836 5623 1843 5663
rect 2496 5656 2523 5663
rect 1856 5636 1883 5643
rect 1936 5636 1943 5653
rect 1876 5627 1883 5636
rect 2076 5636 2083 5653
rect 1836 5616 1863 5623
rect 1856 5607 1863 5616
rect 1616 4943 1623 5093
rect 1616 4936 1643 4943
rect 1636 4927 1643 4936
rect 1556 4707 1563 4893
rect 1596 4676 1623 4683
rect 1596 4663 1603 4676
rect 1576 4656 1603 4663
rect 1476 4627 1483 4643
rect 1396 4496 1423 4503
rect 1436 4496 1443 4533
rect 1396 4263 1403 4496
rect 1396 4256 1423 4263
rect 1387 4236 1403 4243
rect 1396 4216 1403 4236
rect 1136 3707 1143 3723
rect 956 3516 983 3523
rect 1016 3516 1023 3673
rect 756 3227 763 3483
rect 796 3467 803 3483
rect 876 3447 883 3483
rect 816 3223 823 3433
rect 836 3256 843 3293
rect 816 3216 843 3223
rect 836 3027 843 3216
rect 856 3167 863 3243
rect 696 3016 723 3023
rect 656 2967 663 2993
rect 616 2796 643 2803
rect 556 2776 583 2783
rect 536 2687 543 2753
rect 556 2747 563 2776
rect 456 1267 463 2213
rect 476 2067 483 2173
rect 536 2096 543 2233
rect 576 2227 583 2733
rect 636 2707 643 2796
rect 656 2767 663 2953
rect 716 2947 723 3016
rect 756 2987 763 3013
rect 756 2727 763 2973
rect 776 2747 783 2793
rect 796 2787 803 2993
rect 856 2827 863 3093
rect 816 2776 823 2793
rect 856 2776 863 2813
rect 636 2556 643 2653
rect 676 2567 683 2673
rect 596 2207 603 2283
rect 676 2263 683 2293
rect 616 2207 623 2263
rect 656 2256 683 2263
rect 656 2247 663 2256
rect 476 1747 483 2053
rect 516 2047 523 2063
rect 516 1847 523 1873
rect 496 1816 503 1833
rect 516 1747 523 1803
rect 496 1736 513 1743
rect 496 1587 503 1736
rect 516 1596 523 1713
rect 536 1623 543 1813
rect 556 1727 563 1773
rect 576 1647 583 2133
rect 636 2076 643 2213
rect 616 2056 623 2073
rect 656 1947 663 2063
rect 716 2027 723 2673
rect 736 2547 743 2693
rect 876 2687 883 3193
rect 896 2807 903 3453
rect 916 3267 923 3473
rect 916 3036 923 3213
rect 936 3167 943 3493
rect 956 3447 963 3516
rect 976 3207 983 3243
rect 976 3047 983 3173
rect 996 2883 1003 3153
rect 1016 3087 1023 3243
rect 1036 3147 1043 3353
rect 976 2876 1003 2883
rect 896 2727 903 2773
rect 936 2767 943 2773
rect 976 2756 983 2876
rect 756 2556 763 2573
rect 796 2556 803 2593
rect 816 2536 823 2553
rect 876 2547 883 2573
rect 896 2447 903 2713
rect 936 2576 943 2693
rect 756 2296 763 2433
rect 776 2207 783 2283
rect 796 2127 803 2303
rect 936 2296 943 2533
rect 856 2087 863 2273
rect 916 2147 923 2283
rect 956 2267 963 2543
rect 776 2047 783 2063
rect 816 2027 823 2033
rect 716 1847 723 1853
rect 536 1616 553 1623
rect 596 1583 603 1793
rect 576 1576 603 1583
rect 536 1347 543 1573
rect 596 1567 603 1576
rect 476 1303 483 1333
rect 476 1296 503 1303
rect 496 1283 503 1296
rect 556 1287 563 1293
rect 496 1276 543 1283
rect 536 1267 543 1276
rect 436 1147 443 1173
rect 436 1116 443 1133
rect 476 1116 483 1233
rect 456 1087 463 1103
rect 356 856 363 1013
rect 516 967 523 1253
rect 536 1087 543 1213
rect 376 807 383 833
rect 396 807 403 863
rect 436 843 443 853
rect 416 836 443 843
rect 216 463 223 793
rect 236 636 243 793
rect 196 456 223 463
rect 196 343 203 456
rect 296 367 303 413
rect 196 336 243 343
rect 256 156 263 313
rect 276 267 283 343
rect 296 327 303 353
rect 316 347 323 613
rect 336 307 343 793
rect 356 603 363 713
rect 456 623 463 653
rect 436 616 463 623
rect 356 596 383 603
rect 456 547 463 616
rect 416 367 423 373
rect 376 347 383 363
rect 396 307 403 343
rect 436 327 443 343
rect 376 156 383 253
rect 416 176 423 193
rect 176 127 183 153
rect 196 107 203 133
rect 236 127 243 143
rect 456 143 463 353
rect 476 247 483 953
rect 576 907 583 1313
rect 616 1147 623 1633
rect 656 1576 663 1783
rect 716 1767 723 1833
rect 736 1796 763 1803
rect 796 1796 803 1813
rect 836 1807 843 2073
rect 856 2056 883 2063
rect 856 2047 863 2056
rect 896 2047 903 2093
rect 916 2067 923 2113
rect 676 1756 693 1763
rect 736 1707 743 1796
rect 856 1747 863 2033
rect 936 2027 943 2043
rect 956 1827 963 2013
rect 976 1787 983 2513
rect 996 2427 1003 2593
rect 1016 2323 1023 3033
rect 1036 3027 1043 3133
rect 1036 2527 1043 2913
rect 1056 2543 1063 3533
rect 1096 3467 1103 3513
rect 1116 3483 1123 3553
rect 1156 3496 1163 3513
rect 1176 3487 1183 3753
rect 1296 3736 1303 3833
rect 1196 3627 1203 3733
rect 1216 3527 1223 3613
rect 1196 3496 1223 3503
rect 1116 3476 1143 3483
rect 1216 3463 1223 3496
rect 1196 3456 1223 3463
rect 1076 3107 1083 3313
rect 1136 3187 1143 3263
rect 1176 3243 1183 3273
rect 1156 3236 1183 3243
rect 1176 3147 1183 3213
rect 1076 2987 1083 3003
rect 1096 2803 1103 2973
rect 1116 2967 1123 3003
rect 1096 2796 1123 2803
rect 1116 2776 1123 2796
rect 1096 2587 1103 2763
rect 1136 2556 1143 3113
rect 1156 3007 1163 3073
rect 1156 2847 1163 2933
rect 1056 2536 1083 2543
rect 996 2316 1023 2323
rect 996 2083 1003 2316
rect 1056 2303 1063 2536
rect 1156 2523 1163 2833
rect 1176 2607 1183 3053
rect 1196 2687 1203 3456
rect 1236 3327 1243 3713
rect 1276 3627 1283 3723
rect 1316 3647 1323 3933
rect 1336 3767 1343 4013
rect 1356 3747 1363 4173
rect 1416 4003 1423 4256
rect 1436 4207 1443 4453
rect 1456 4183 1463 4473
rect 1476 4347 1483 4613
rect 1536 4476 1543 4513
rect 1516 4427 1523 4463
rect 1556 4456 1563 4473
rect 1516 4216 1523 4233
rect 1456 4176 1483 4183
rect 1416 3996 1443 4003
rect 1396 3976 1403 3993
rect 1376 3947 1383 3963
rect 1336 3527 1343 3733
rect 1296 3467 1303 3483
rect 1256 3303 1263 3453
rect 1236 3296 1263 3303
rect 1216 3247 1223 3253
rect 1236 3247 1243 3296
rect 1256 3247 1263 3273
rect 1236 3187 1243 3203
rect 1216 3036 1223 3153
rect 1236 3056 1243 3133
rect 1276 3067 1283 3223
rect 1296 3127 1303 3433
rect 1336 3147 1343 3493
rect 1356 3487 1363 3733
rect 1396 3727 1403 3753
rect 1416 3747 1423 3963
rect 1436 3747 1443 3996
rect 1456 3727 1463 3993
rect 1396 3667 1403 3683
rect 1376 3607 1383 3633
rect 1376 3447 1383 3593
rect 1416 3496 1423 3513
rect 1256 3036 1283 3043
rect 1276 2967 1283 3036
rect 1316 3036 1323 3053
rect 1356 3036 1363 3293
rect 1396 3127 1403 3203
rect 1296 2827 1303 3033
rect 1376 3016 1403 3023
rect 1396 2927 1403 3016
rect 1416 3007 1423 3453
rect 1476 3407 1483 4176
rect 1496 4047 1503 4203
rect 1536 4047 1543 4193
rect 1556 4127 1563 4413
rect 1576 4163 1583 4656
rect 1596 4627 1603 4633
rect 1596 4427 1603 4613
rect 1616 4207 1623 4653
rect 1656 4527 1663 5153
rect 1696 4943 1703 5113
rect 1716 4956 1723 4973
rect 1756 4956 1763 5133
rect 1776 5127 1783 5413
rect 1836 5396 1843 5593
rect 1916 5587 1923 5593
rect 1856 5416 1863 5453
rect 1916 5187 1923 5573
rect 1956 5416 1963 5433
rect 1976 5407 1983 5473
rect 2056 5467 2063 5623
rect 2096 5467 2103 5623
rect 2116 5607 2123 5653
rect 1996 5416 2023 5423
rect 1936 5183 1943 5403
rect 2016 5387 2023 5416
rect 1936 5176 1963 5183
rect 1896 5163 1903 5173
rect 1896 5156 1923 5163
rect 1776 4947 1783 5033
rect 1796 4947 1803 5153
rect 1876 5127 1883 5143
rect 1916 5047 1923 5156
rect 1956 4963 1963 5176
rect 1996 4983 2003 5193
rect 2016 5143 2023 5213
rect 2036 5207 2043 5413
rect 2096 5387 2103 5393
rect 2056 5156 2063 5173
rect 2096 5156 2103 5193
rect 2136 5167 2143 5633
rect 2216 5627 2223 5643
rect 2276 5636 2303 5643
rect 2156 5607 2163 5623
rect 2196 5607 2203 5623
rect 2216 5563 2223 5613
rect 2276 5567 2283 5636
rect 2376 5623 2383 5653
rect 2356 5616 2383 5623
rect 2316 5587 2323 5603
rect 2196 5556 2223 5563
rect 2196 5423 2203 5556
rect 2316 5436 2323 5553
rect 2376 5547 2383 5616
rect 2416 5467 2423 5633
rect 2516 5467 2523 5656
rect 2556 5656 2583 5663
rect 2556 5487 2563 5656
rect 2816 5656 2843 5663
rect 2416 5443 2423 5453
rect 2376 5436 2403 5443
rect 2196 5416 2223 5423
rect 2176 5183 2183 5293
rect 2196 5227 2203 5416
rect 2336 5307 2343 5403
rect 2396 5207 2403 5436
rect 2416 5436 2443 5443
rect 2156 5176 2183 5183
rect 2216 5176 2223 5193
rect 2016 5136 2043 5143
rect 2116 5107 2123 5143
rect 2156 5107 2163 5176
rect 1996 4976 2023 4983
rect 1936 4956 1963 4963
rect 1676 4936 1703 4943
rect 1676 4907 1683 4936
rect 1816 4927 1823 4943
rect 1816 4807 1823 4913
rect 1716 4683 1723 4693
rect 1716 4676 1743 4683
rect 1716 4667 1723 4676
rect 1676 4456 1683 4593
rect 1716 4467 1723 4633
rect 1756 4563 1763 4663
rect 1736 4556 1763 4563
rect 1656 4227 1663 4443
rect 1696 4407 1703 4443
rect 1576 4156 1603 4163
rect 1536 4016 1543 4033
rect 1516 3747 1523 3983
rect 1556 3947 1563 4033
rect 1536 3716 1543 3753
rect 1496 3687 1503 3713
rect 1596 3647 1603 4156
rect 1636 4127 1643 4183
rect 1656 4163 1663 4213
rect 1676 4187 1683 4273
rect 1736 4267 1743 4556
rect 1756 4443 1763 4533
rect 1796 4456 1803 4493
rect 1816 4447 1823 4533
rect 1836 4467 1843 4573
rect 1756 4436 1783 4443
rect 1796 4227 1803 4413
rect 1856 4387 1863 4893
rect 1896 4723 1903 4933
rect 1916 4927 1923 4953
rect 1887 4716 1903 4723
rect 1876 4696 1883 4713
rect 1936 4703 1943 4956
rect 2016 4923 2023 4976
rect 2096 4956 2103 5033
rect 2196 4947 2203 5153
rect 2276 4976 2283 5153
rect 2356 5067 2363 5173
rect 2376 5127 2383 5163
rect 2416 5147 2423 5436
rect 2456 5403 2463 5423
rect 2496 5416 2503 5453
rect 2436 5396 2463 5403
rect 2156 4927 2163 4943
rect 2356 4936 2363 5053
rect 2436 5047 2443 5396
rect 2556 5387 2563 5433
rect 2476 5156 2483 5173
rect 2527 5156 2543 5163
rect 2376 4956 2383 4973
rect 1996 4916 2023 4923
rect 1916 4696 1943 4703
rect 1696 4216 1723 4223
rect 1656 4156 1683 4163
rect 1616 4103 1623 4113
rect 1616 4096 1663 4103
rect 1656 4047 1663 4096
rect 1656 3996 1663 4013
rect 1496 3516 1523 3523
rect 1556 3516 1563 3633
rect 1496 3287 1503 3516
rect 1236 2667 1243 2763
rect 1316 2747 1323 2773
rect 1136 2516 1163 2523
rect 1036 2296 1063 2303
rect 1016 2276 1023 2293
rect 1036 2247 1043 2296
rect 1056 2227 1063 2263
rect 1096 2227 1103 2393
rect 1116 2087 1123 2293
rect 1136 2276 1143 2516
rect 996 2076 1023 2083
rect 996 1767 1003 2053
rect 1016 1887 1023 2076
rect 1116 2056 1123 2073
rect 1136 1847 1143 2073
rect 1036 1767 1043 1793
rect 956 1747 963 1763
rect 736 1627 743 1693
rect 696 1563 703 1613
rect 856 1587 863 1733
rect 896 1596 903 1613
rect 936 1596 943 1653
rect 876 1576 883 1593
rect 676 1556 703 1563
rect 636 1307 643 1323
rect 656 1267 663 1303
rect 616 1096 623 1113
rect 656 1096 663 1153
rect 676 1087 683 1133
rect 696 1123 703 1303
rect 696 1116 723 1123
rect 756 1116 763 1533
rect 956 1527 963 1733
rect 976 1587 983 1613
rect 816 1336 823 1353
rect 916 1336 923 1353
rect 876 1303 883 1333
rect 856 1296 883 1303
rect 936 1167 943 1323
rect 696 1087 703 1116
rect 776 1107 783 1153
rect 996 1147 1003 1753
rect 1056 1747 1063 1803
rect 1076 1603 1083 1783
rect 1136 1687 1143 1753
rect 1056 1596 1083 1603
rect 1036 1587 1043 1593
rect 1016 1367 1023 1563
rect 1056 1556 1063 1596
rect 1096 1583 1103 1653
rect 1076 1576 1103 1583
rect 1096 1283 1103 1576
rect 1136 1563 1143 1673
rect 1156 1607 1163 2253
rect 1176 2227 1183 2573
rect 1256 2563 1263 2743
rect 1296 2707 1303 2743
rect 1336 2727 1343 2753
rect 1356 2667 1363 2743
rect 1256 2556 1283 2563
rect 1316 2556 1343 2563
rect 1376 2556 1403 2563
rect 1196 2447 1203 2533
rect 1276 2527 1283 2556
rect 1216 2507 1223 2523
rect 1256 2516 1273 2523
rect 1336 2507 1343 2556
rect 1196 2203 1203 2433
rect 1396 2347 1403 2556
rect 1416 2547 1423 2553
rect 1416 2307 1423 2533
rect 1436 2307 1443 3233
rect 1496 3207 1503 3243
rect 1516 3227 1523 3263
rect 1556 3243 1563 3273
rect 1536 3236 1563 3243
rect 1496 3016 1503 3073
rect 1516 2996 1523 3053
rect 1536 3027 1543 3113
rect 1556 2987 1563 3193
rect 1576 3067 1583 3253
rect 1596 3247 1603 3613
rect 1616 3487 1623 3493
rect 1616 3267 1623 3473
rect 1636 3467 1643 3973
rect 1676 3867 1683 4156
rect 1696 4147 1703 4216
rect 1736 4187 1743 4203
rect 1816 4167 1823 4373
rect 1696 3987 1703 4033
rect 1676 3716 1683 3733
rect 1716 3567 1723 4153
rect 1736 3727 1743 3983
rect 1816 3976 1823 4033
rect 1836 4027 1843 4253
rect 1856 4216 1863 4273
rect 1896 4267 1903 4683
rect 1956 4667 1963 4913
rect 1996 4687 2003 4916
rect 1967 4656 1983 4663
rect 1936 4496 1943 4553
rect 2016 4527 2023 4663
rect 2036 4647 2043 4683
rect 1956 4476 1963 4493
rect 1936 4267 1943 4453
rect 1976 4363 1983 4513
rect 2027 4496 2043 4503
rect 2036 4487 2043 4496
rect 2016 4443 2023 4473
rect 2076 4447 2083 4673
rect 2096 4587 2103 4653
rect 2096 4456 2103 4573
rect 2016 4436 2043 4443
rect 1956 4356 1983 4363
rect 1876 4187 1883 4203
rect 1836 3956 1843 4013
rect 1876 4007 1883 4173
rect 1896 4167 1903 4223
rect 1936 4207 1943 4253
rect 1916 4196 1933 4203
rect 1876 3767 1883 3963
rect 1896 3767 1903 3973
rect 1756 3736 1783 3743
rect 1816 3736 1823 3753
rect 1756 3707 1763 3736
rect 1916 3736 1943 3743
rect 1656 3487 1663 3533
rect 1756 3503 1763 3573
rect 1696 3496 1723 3503
rect 1696 3243 1703 3473
rect 1716 3247 1723 3496
rect 1736 3496 1763 3503
rect 1736 3287 1743 3496
rect 1756 3263 1763 3453
rect 1776 3307 1783 3493
rect 1736 3256 1763 3263
rect 1676 3236 1703 3243
rect 1676 3227 1683 3236
rect 1476 2563 1483 2753
rect 1496 2747 1503 2953
rect 1576 2647 1583 2723
rect 1596 2707 1603 3093
rect 1616 2887 1623 3133
rect 1716 3027 1723 3233
rect 1736 3123 1743 3256
rect 1776 3236 1783 3293
rect 1796 3247 1803 3723
rect 1936 3667 1943 3736
rect 1956 3707 1963 4356
rect 2056 4247 2063 4413
rect 2116 4267 2123 4773
rect 2136 4696 2143 4733
rect 2156 4467 2163 4683
rect 2176 4647 2183 4703
rect 2196 4667 2203 4683
rect 2176 4547 2183 4633
rect 2216 4487 2223 4493
rect 2156 4287 2163 4453
rect 2176 4443 2183 4473
rect 2216 4456 2223 4473
rect 2176 4436 2203 4443
rect 2236 4436 2243 4713
rect 2356 4696 2383 4703
rect 2416 4696 2423 4733
rect 2356 4687 2363 4696
rect 2436 4687 2443 5013
rect 2256 4456 2263 4653
rect 2316 4627 2323 4663
rect 1996 4167 2003 4223
rect 2056 4187 2063 4233
rect 1976 3987 1983 4093
rect 1996 3996 2003 4053
rect 2036 3996 2043 4053
rect 2016 3947 2023 3983
rect 1976 3687 1983 3933
rect 2056 3807 2063 4093
rect 2076 3987 2083 4213
rect 2096 4203 2103 4253
rect 2176 4216 2183 4233
rect 2096 4196 2123 4203
rect 1996 3727 2003 3753
rect 2036 3703 2043 3733
rect 2056 3716 2063 3733
rect 2016 3696 2043 3703
rect 1996 3667 2003 3683
rect 1836 3496 1843 3513
rect 1856 3476 1863 3493
rect 1896 3307 1903 3633
rect 1916 3507 1923 3533
rect 1996 3516 2003 3553
rect 2016 3507 2023 3513
rect 1816 3236 1823 3273
rect 1756 3167 1763 3223
rect 1736 3116 1763 3123
rect 1656 2967 1663 3013
rect 1696 3007 1703 3023
rect 1716 2983 1723 3013
rect 1736 3007 1743 3073
rect 1716 2976 1743 2983
rect 1676 2727 1683 2743
rect 1656 2707 1663 2723
rect 1476 2556 1503 2563
rect 1496 2536 1503 2556
rect 1476 2507 1483 2523
rect 1296 2247 1303 2303
rect 1336 2283 1343 2293
rect 1316 2276 1343 2283
rect 1416 2276 1423 2293
rect 1456 2287 1463 2373
rect 1176 2196 1203 2203
rect 1176 1807 1183 2196
rect 1276 2067 1283 2093
rect 1236 1807 1243 1833
rect 1196 1767 1203 1803
rect 1136 1556 1163 1563
rect 1156 1307 1163 1343
rect 1216 1327 1223 1783
rect 1276 1603 1283 1793
rect 1296 1647 1303 2213
rect 1356 2076 1363 2113
rect 1396 2107 1403 2263
rect 1316 2056 1343 2063
rect 1316 1727 1323 2056
rect 1396 1787 1403 1933
rect 1356 1756 1383 1763
rect 1256 1596 1283 1603
rect 1316 1596 1323 1673
rect 1256 1567 1263 1596
rect 1256 1343 1263 1513
rect 1256 1336 1283 1343
rect 1316 1336 1323 1553
rect 1256 1287 1263 1336
rect 1296 1307 1303 1323
rect 1076 1276 1103 1283
rect 936 1116 943 1133
rect 1096 1116 1123 1123
rect 676 1027 683 1073
rect 556 847 563 853
rect 616 827 623 893
rect 636 856 643 1013
rect 736 907 743 1103
rect 656 787 663 843
rect 676 836 703 843
rect 676 767 683 836
rect 716 823 723 853
rect 696 816 723 823
rect 736 836 763 843
rect 796 836 803 853
rect 576 636 603 643
rect 696 636 703 816
rect 736 787 743 836
rect 776 767 783 803
rect 596 627 603 636
rect 516 376 523 533
rect 556 427 563 623
rect 476 147 483 233
rect 436 136 463 143
rect 516 136 523 213
rect 556 207 563 383
rect 576 247 583 363
rect 596 267 603 613
rect 636 607 643 623
rect 836 603 843 1113
rect 1116 1107 1123 1116
rect 896 1096 923 1103
rect 896 1087 903 1096
rect 1076 1083 1083 1103
rect 1076 1076 1113 1083
rect 856 607 863 833
rect 776 587 783 603
rect 816 596 843 603
rect 676 376 683 573
rect 816 407 823 596
rect 736 343 743 393
rect 716 336 743 343
rect 816 287 823 363
rect 536 156 543 173
rect 576 156 583 173
rect 636 156 643 173
rect 676 156 683 193
rect 816 136 823 273
rect 836 227 843 383
rect 876 363 883 873
rect 896 827 903 1073
rect 1136 867 1143 1153
rect 1316 1116 1323 1273
rect 1336 1147 1343 1613
rect 1176 1083 1183 1103
rect 1167 1076 1183 1083
rect 1216 887 1223 1113
rect 1256 1087 1263 1103
rect 1036 856 1063 863
rect 1016 827 1023 833
rect 936 807 943 823
rect 936 616 943 673
rect 956 636 963 773
rect 976 667 983 823
rect 996 636 1003 653
rect 1016 627 1023 813
rect 1036 767 1043 856
rect 1096 807 1103 863
rect 1136 847 1143 853
rect 1096 647 1103 793
rect 1116 783 1123 843
rect 1136 807 1143 833
rect 1176 807 1183 823
rect 1236 807 1243 843
rect 1116 776 1143 783
rect 1096 616 1103 633
rect 856 356 883 363
rect 956 356 963 373
rect 976 367 983 613
rect 1116 596 1123 673
rect 1136 627 1143 776
rect 1216 656 1223 673
rect 1256 636 1263 1053
rect 1296 827 1303 1033
rect 1336 887 1343 1133
rect 1356 1047 1363 1733
rect 1376 1727 1383 1756
rect 1416 1747 1423 2213
rect 1476 2147 1483 2293
rect 1496 2267 1503 2453
rect 1516 2227 1523 2273
rect 1536 2263 1543 2493
rect 1556 2487 1563 2513
rect 1576 2507 1583 2613
rect 1596 2576 1603 2653
rect 1636 2527 1643 2693
rect 1676 2643 1683 2713
rect 1667 2636 1683 2643
rect 1696 2607 1703 2973
rect 1656 2563 1663 2593
rect 1656 2556 1683 2563
rect 1596 2276 1603 2313
rect 1536 2256 1563 2263
rect 1436 1767 1443 1803
rect 1476 1796 1483 1973
rect 1556 1943 1563 2256
rect 1576 2247 1583 2263
rect 1616 2227 1623 2263
rect 1576 1947 1583 2113
rect 1536 1936 1563 1943
rect 1536 1787 1543 1936
rect 1596 1823 1603 2133
rect 1636 2067 1643 2353
rect 1656 2087 1663 2333
rect 1676 2087 1683 2556
rect 1736 2556 1743 2976
rect 1756 2707 1763 3116
rect 1796 3036 1803 3173
rect 1836 3047 1843 3133
rect 1796 2776 1823 2783
rect 1816 2767 1823 2776
rect 1836 2727 1843 2743
rect 1716 2523 1723 2543
rect 1696 2516 1723 2523
rect 1696 2467 1703 2516
rect 1716 2347 1723 2493
rect 1747 2476 1753 2483
rect 1716 2287 1723 2293
rect 1736 2287 1743 2453
rect 1756 2276 1763 2353
rect 1756 2227 1763 2233
rect 1656 2063 1663 2073
rect 1656 2056 1673 2063
rect 1696 2047 1703 2093
rect 1616 2027 1623 2043
rect 1576 1816 1603 1823
rect 1576 1796 1583 1816
rect 1616 1787 1623 1803
rect 1396 1596 1423 1603
rect 1376 1427 1383 1593
rect 1396 1507 1403 1596
rect 1436 1363 1443 1673
rect 1456 1627 1463 1783
rect 1456 1596 1483 1603
rect 1476 1567 1483 1596
rect 1416 1356 1443 1363
rect 1416 1336 1423 1356
rect 1436 1167 1443 1323
rect 1436 1136 1463 1143
rect 1376 1107 1383 1133
rect 1416 1087 1423 1103
rect 1456 1087 1463 1136
rect 1316 856 1343 863
rect 1156 547 1163 633
rect 1196 607 1203 613
rect 1316 587 1323 856
rect 1416 843 1423 853
rect 1396 836 1423 843
rect 856 207 863 356
rect 976 307 983 323
rect 1016 227 1023 413
rect 1116 376 1123 533
rect 1036 283 1043 373
rect 1056 307 1063 363
rect 1196 356 1223 363
rect 1196 287 1203 356
rect 1236 323 1243 553
rect 1336 347 1343 733
rect 1376 567 1383 623
rect 1416 587 1423 613
rect 1416 347 1423 363
rect 1216 316 1243 323
rect 1036 276 1063 283
rect 856 136 863 193
rect 916 176 923 213
rect 876 147 883 173
rect 836 127 843 133
rect 896 127 903 173
rect 1016 156 1023 213
rect 1056 156 1063 276
rect 936 127 943 143
rect 956 127 963 153
rect 1036 127 1043 143
rect 1076 136 1083 273
rect 1136 143 1143 193
rect 1216 156 1223 316
rect 1236 147 1243 173
rect 1276 167 1283 323
rect 1336 187 1343 333
rect 1436 203 1443 873
rect 1456 867 1463 1073
rect 1496 1067 1503 1733
rect 1516 1167 1523 1753
rect 1596 1687 1603 1783
rect 1636 1627 1643 1793
rect 1676 1596 1683 2013
rect 1716 1987 1723 2193
rect 1756 2103 1763 2213
rect 1776 2127 1783 2653
rect 1796 2567 1803 2693
rect 1796 2507 1803 2533
rect 1816 2487 1823 2553
rect 1836 2543 1843 2713
rect 1856 2607 1863 3293
rect 1916 3283 1923 3493
rect 1936 3467 1943 3503
rect 1976 3487 1983 3503
rect 1936 3307 1943 3453
rect 1896 3276 1923 3283
rect 1896 3207 1903 3276
rect 1956 3256 1983 3263
rect 1936 3207 1943 3243
rect 1896 3043 1903 3153
rect 1876 3036 1903 3043
rect 1936 3036 1943 3073
rect 1976 3067 1983 3256
rect 1876 3027 1883 3036
rect 1956 3016 1983 3023
rect 1976 2987 1983 3016
rect 1916 2667 1923 2853
rect 1936 2776 1943 2793
rect 1976 2776 1983 2933
rect 1996 2807 2003 3373
rect 2016 3287 2023 3493
rect 2036 3447 2043 3673
rect 2016 3047 2023 3273
rect 2056 3236 2063 3513
rect 2076 3307 2083 3793
rect 2096 3727 2103 4173
rect 2116 3707 2123 4173
rect 2136 4167 2143 4213
rect 2196 4207 2203 4273
rect 2156 4047 2163 4193
rect 2176 3956 2183 4013
rect 2136 3736 2143 3753
rect 2096 3683 2103 3693
rect 2096 3676 2123 3683
rect 2116 3516 2123 3676
rect 2156 3547 2163 3723
rect 2216 3627 2223 4313
rect 2236 4187 2243 4233
rect 2276 4223 2283 4553
rect 2396 4443 2403 4653
rect 2456 4587 2463 4953
rect 2536 4927 2543 5156
rect 2556 5147 2563 5193
rect 2596 5156 2603 5433
rect 2676 5416 2683 5433
rect 2696 5363 2703 5633
rect 2736 5607 2743 5643
rect 2776 5567 2783 5643
rect 2776 5416 2783 5533
rect 2796 5396 2803 5653
rect 2816 5567 2823 5656
rect 2816 5416 2823 5553
rect 2856 5467 2863 5643
rect 2996 5547 3003 5603
rect 2856 5427 2863 5453
rect 2876 5436 2883 5533
rect 2916 5436 2923 5453
rect 2936 5416 2943 5473
rect 3096 5447 3103 5623
rect 3136 5607 3143 5623
rect 3436 5623 3443 5653
rect 3416 5616 3443 5623
rect 3396 5527 3403 5593
rect 3036 5407 3043 5423
rect 3256 5416 3263 5453
rect 3436 5447 3443 5616
rect 3496 5463 3503 5613
rect 3496 5456 3523 5463
rect 3156 5387 3163 5403
rect 2676 5356 2703 5363
rect 2676 5127 2683 5356
rect 3016 5176 3043 5183
rect 2556 4943 2563 5113
rect 2656 4976 2663 5053
rect 2696 5027 2703 5163
rect 2716 5127 2723 5143
rect 2756 4987 2763 5143
rect 2556 4936 2583 4943
rect 2576 4903 2583 4936
rect 2776 4936 2783 4973
rect 2556 4896 2583 4903
rect 2536 4727 2543 4873
rect 2536 4696 2543 4713
rect 2516 4607 2523 4673
rect 2476 4467 2483 4493
rect 2336 4427 2343 4443
rect 2376 4436 2403 4443
rect 2336 4407 2343 4413
rect 2256 4216 2283 4223
rect 2256 4107 2263 4216
rect 2316 4107 2323 4183
rect 2336 4167 2343 4353
rect 2356 4187 2363 4253
rect 2247 3976 2263 3983
rect 2236 3723 2243 3973
rect 2276 3956 2283 4013
rect 2376 4007 2383 4333
rect 2396 4227 2403 4436
rect 2416 4327 2423 4453
rect 2436 4307 2443 4453
rect 2456 4347 2463 4443
rect 2496 4436 2503 4513
rect 2556 4463 2563 4896
rect 2596 4867 2603 4913
rect 2796 4907 2803 4923
rect 2576 4667 2583 4693
rect 2596 4567 2603 4853
rect 2536 4456 2563 4463
rect 2576 4456 2583 4513
rect 2616 4456 2623 4493
rect 2416 4147 2423 4203
rect 2456 4196 2463 4253
rect 2476 4167 2483 4183
rect 2296 3976 2303 3993
rect 2336 3767 2343 3993
rect 2396 3887 2403 4113
rect 2416 3987 2423 4093
rect 2496 4083 2503 4233
rect 2516 4127 2523 4253
rect 2496 4076 2523 4083
rect 2496 3987 2503 4013
rect 2456 3927 2463 3983
rect 2516 3967 2523 4076
rect 2276 3727 2283 3743
rect 2236 3716 2263 3723
rect 2256 3667 2263 3716
rect 2256 3543 2263 3573
rect 2276 3567 2283 3713
rect 2296 3707 2303 3723
rect 2336 3703 2343 3753
rect 2316 3696 2343 3703
rect 2256 3536 2283 3543
rect 2176 3507 2183 3533
rect 2036 3147 2043 3223
rect 2076 3196 2103 3203
rect 2036 2867 2043 3073
rect 2076 3016 2083 3053
rect 2096 3036 2103 3196
rect 2116 3087 2123 3393
rect 2196 3287 2203 3533
rect 2216 3516 2243 3523
rect 2276 3516 2283 3536
rect 2216 3487 2223 3516
rect 2296 3496 2303 3513
rect 2316 3483 2323 3696
rect 2336 3507 2343 3533
rect 2316 3476 2343 3483
rect 2147 3256 2163 3263
rect 2136 3107 2143 3253
rect 2136 3036 2163 3043
rect 2156 3007 2163 3036
rect 1996 2747 2003 2793
rect 2016 2743 2023 2773
rect 2056 2756 2063 2813
rect 2016 2736 2043 2743
rect 1916 2556 1923 2613
rect 1836 2536 1863 2543
rect 1836 2487 1843 2536
rect 1896 2523 1903 2543
rect 1876 2516 1903 2523
rect 1796 2267 1803 2473
rect 1876 2467 1883 2516
rect 1816 2227 1823 2453
rect 1876 2447 1883 2453
rect 1836 2296 1843 2333
rect 1896 2323 1903 2473
rect 1896 2316 1923 2323
rect 1916 2307 1923 2316
rect 1896 2276 1923 2283
rect 1736 2096 1763 2103
rect 1736 2076 1743 2096
rect 1776 2076 1783 2093
rect 1816 2063 1823 2193
rect 1756 2047 1763 2063
rect 1796 2056 1823 2063
rect 1696 1803 1703 1853
rect 1756 1807 1763 1933
rect 1696 1796 1723 1803
rect 1716 1603 1723 1796
rect 1736 1627 1743 1773
rect 1776 1767 1783 1783
rect 1816 1747 1823 2056
rect 1836 2027 1843 2173
rect 1876 2167 1883 2273
rect 1916 2267 1923 2276
rect 1896 2187 1903 2253
rect 1936 2127 1943 2593
rect 1836 1767 1843 1953
rect 1856 1867 1863 2113
rect 1916 1823 1923 1913
rect 1896 1816 1923 1823
rect 1876 1727 1883 1803
rect 1716 1596 1743 1603
rect 1556 1363 1563 1573
rect 1536 1356 1563 1363
rect 1536 1336 1543 1356
rect 1596 1343 1603 1593
rect 1696 1387 1703 1583
rect 1736 1367 1743 1596
rect 1776 1567 1783 1583
rect 1796 1523 1803 1673
rect 1776 1516 1803 1523
rect 1576 1336 1603 1343
rect 1516 1116 1523 1153
rect 1556 1116 1563 1173
rect 1476 836 1483 853
rect 1456 367 1463 693
rect 1536 687 1543 1093
rect 1596 887 1603 1336
rect 1756 1323 1763 1373
rect 1736 1316 1763 1323
rect 1596 856 1603 873
rect 1616 807 1623 1173
rect 1636 1136 1643 1153
rect 1656 887 1663 1103
rect 1776 1096 1783 1516
rect 1796 1336 1803 1373
rect 1836 1336 1843 1613
rect 1856 1576 1863 1693
rect 1916 1687 1923 1816
rect 1936 1747 1943 1873
rect 1956 1827 1963 2733
rect 1976 2556 1983 2573
rect 1996 2527 2003 2543
rect 1976 2296 1983 2373
rect 2056 2327 2063 2573
rect 1996 2207 2003 2283
rect 2036 2267 2043 2283
rect 1976 1947 1983 2113
rect 1996 2087 2003 2193
rect 2056 2103 2063 2313
rect 2076 2303 2083 2743
rect 2096 2667 2103 2763
rect 2116 2547 2123 2813
rect 2136 2567 2143 2893
rect 2156 2747 2163 2993
rect 2176 2827 2183 3113
rect 2196 2967 2203 3213
rect 2216 3207 2223 3473
rect 2236 3227 2243 3253
rect 2236 3063 2243 3213
rect 2256 3127 2263 3273
rect 2276 3203 2283 3433
rect 2316 3256 2323 3293
rect 2276 3196 2303 3203
rect 2216 3056 2243 3063
rect 2216 3016 2223 3056
rect 2256 2943 2263 3013
rect 2256 2936 2283 2943
rect 2096 2427 2103 2533
rect 2176 2527 2183 2793
rect 2196 2787 2203 2893
rect 2196 2536 2203 2593
rect 2116 2347 2123 2513
rect 2136 2367 2143 2523
rect 2136 2323 2143 2353
rect 2156 2327 2163 2493
rect 2216 2467 2223 2733
rect 2236 2603 2243 2913
rect 2256 2707 2263 2743
rect 2236 2596 2263 2603
rect 2236 2467 2243 2553
rect 2256 2487 2263 2596
rect 2276 2587 2283 2936
rect 2296 2727 2303 3196
rect 2316 2807 2323 3153
rect 2336 3147 2343 3476
rect 2356 3467 2363 3513
rect 2376 3507 2383 3813
rect 2396 3587 2403 3793
rect 2456 3727 2463 3873
rect 2476 3807 2483 3873
rect 2436 3647 2443 3703
rect 2436 3536 2443 3573
rect 2396 3516 2403 3533
rect 2376 3223 2383 3493
rect 2416 3383 2423 3503
rect 2396 3376 2423 3383
rect 2396 3227 2403 3376
rect 2416 3256 2423 3293
rect 2456 3256 2463 3493
rect 2356 3216 2383 3223
rect 2356 3067 2363 3113
rect 2356 3027 2363 3053
rect 2376 3036 2383 3193
rect 2436 3127 2443 3243
rect 2476 3223 2483 3253
rect 2456 3216 2483 3223
rect 2316 2776 2343 2783
rect 2316 2707 2323 2776
rect 2387 2776 2403 2783
rect 2396 2727 2403 2776
rect 2416 2767 2423 3013
rect 2436 2927 2443 3023
rect 2316 2576 2323 2593
rect 2276 2556 2283 2573
rect 2296 2527 2303 2543
rect 2336 2487 2343 2533
rect 2356 2527 2363 2573
rect 2116 2316 2143 2323
rect 2076 2296 2103 2303
rect 2096 2227 2103 2296
rect 2116 2267 2123 2316
rect 2056 2096 2083 2103
rect 2076 2067 2083 2096
rect 2076 2047 2083 2053
rect 1976 1816 1983 1873
rect 2016 1816 2023 1973
rect 1996 1687 2003 1803
rect 2036 1487 2043 1573
rect 1796 1076 1803 1233
rect 1816 1127 1823 1323
rect 1836 1103 1843 1133
rect 1816 1096 1843 1103
rect 1516 647 1523 653
rect 1476 616 1503 623
rect 1476 567 1483 616
rect 1516 596 1523 633
rect 1476 347 1483 393
rect 1596 387 1603 613
rect 1636 427 1643 853
rect 1736 827 1743 843
rect 1756 787 1763 863
rect 1816 827 1823 993
rect 1836 847 1843 1096
rect 1856 1067 1863 1113
rect 1876 1087 1883 1333
rect 1996 1287 2003 1323
rect 2016 1187 2023 1333
rect 2056 1327 2063 1933
rect 2116 1796 2123 1833
rect 2136 1607 2143 2293
rect 2156 2167 2163 2283
rect 2176 2247 2183 2373
rect 2176 2083 2183 2233
rect 2196 2087 2203 2313
rect 2156 2076 2183 2083
rect 2156 1796 2163 1813
rect 2196 1796 2203 1813
rect 2136 1576 2163 1583
rect 2076 1316 2083 1373
rect 2076 1116 2083 1173
rect 1896 1067 1903 1083
rect 1856 856 1863 873
rect 1876 827 1883 843
rect 1656 627 1663 653
rect 1696 387 1703 613
rect 1516 356 1523 373
rect 1656 356 1663 373
rect 1716 367 1723 593
rect 1616 327 1623 353
rect 1736 347 1743 633
rect 1776 627 1783 793
rect 1956 747 1963 1073
rect 1996 787 2003 863
rect 2016 827 2023 843
rect 1816 687 1823 693
rect 1816 616 1823 673
rect 1856 627 1863 693
rect 1976 636 1983 753
rect 1996 747 2003 773
rect 1996 647 2003 653
rect 1996 627 2003 633
rect 1796 587 1803 603
rect 1636 307 1643 343
rect 1416 196 1443 203
rect 1336 156 1343 173
rect 1416 167 1423 196
rect 1596 176 1603 193
rect 1136 136 1163 143
rect 796 107 803 123
rect 1436 123 1443 173
rect 1476 156 1503 163
rect 1496 127 1503 156
rect 1736 156 1743 173
rect 1756 147 1763 343
rect 1436 116 1463 123
rect 1796 123 1803 153
rect 1836 136 1843 553
rect 1916 407 1923 613
rect 2056 607 2063 853
rect 2076 827 2083 1053
rect 2096 767 2103 1253
rect 2116 1107 2123 1473
rect 2136 1447 2143 1576
rect 2136 907 2143 1373
rect 2176 1303 2183 1773
rect 2216 1563 2223 1833
rect 2236 1807 2243 2153
rect 2276 2056 2283 2173
rect 2336 2063 2343 2213
rect 2356 2203 2363 2513
rect 2376 2387 2383 2553
rect 2416 2536 2423 2593
rect 2436 2567 2443 2793
rect 2456 2787 2463 3216
rect 2476 3007 2483 3053
rect 2496 3003 2503 3953
rect 2516 3887 2523 3953
rect 2536 3887 2543 4456
rect 2636 4387 2643 4443
rect 2656 4407 2663 4733
rect 2676 4627 2683 4663
rect 2676 4607 2683 4613
rect 2556 4216 2583 4223
rect 2556 4147 2563 4216
rect 2596 4187 2603 4193
rect 2596 4003 2603 4013
rect 2576 3996 2603 4003
rect 2576 3976 2583 3996
rect 2616 3987 2623 4223
rect 2676 4147 2683 4573
rect 2696 4307 2703 4693
rect 2816 4687 2823 5173
rect 2836 4907 2843 5033
rect 2856 4987 2863 5163
rect 3036 5147 3043 5176
rect 2916 5127 2923 5143
rect 2976 4916 2983 4953
rect 2996 4936 3003 5013
rect 3036 4923 3043 5093
rect 3056 5007 3063 5143
rect 3156 5007 3163 5143
rect 3116 4936 3123 4993
rect 3176 4987 3183 5413
rect 3276 5396 3283 5433
rect 3256 5156 3283 5163
rect 3176 4956 3203 4963
rect 3156 4923 3163 4943
rect 3016 4916 3043 4923
rect 3136 4916 3163 4923
rect 2736 4667 2743 4683
rect 2776 4667 2783 4683
rect 2776 4647 2783 4653
rect 2756 4496 2763 4553
rect 2716 4447 2723 4493
rect 2836 4483 2843 4553
rect 2876 4527 2883 4913
rect 3136 4847 3143 4916
rect 3176 4903 3183 4913
rect 3156 4896 3183 4903
rect 2956 4663 2963 4693
rect 3036 4676 3043 4693
rect 2896 4587 2903 4663
rect 2936 4656 2963 4663
rect 2916 4627 2923 4643
rect 3016 4587 3023 4663
rect 3056 4643 3063 4663
rect 3036 4636 3063 4643
rect 2816 4476 2843 4483
rect 2716 4227 2723 4253
rect 2696 4127 2703 4163
rect 2636 3987 2643 3993
rect 2676 3976 2683 3993
rect 2647 3956 2663 3963
rect 2516 3736 2543 3743
rect 2576 3736 2583 3753
rect 2516 3667 2523 3736
rect 2596 3687 2603 3933
rect 2616 3927 2623 3953
rect 2516 3127 2523 3633
rect 2596 3516 2603 3613
rect 2556 3367 2563 3413
rect 2576 3287 2583 3513
rect 2616 3327 2623 3873
rect 2636 3667 2643 3953
rect 2656 3807 2663 3873
rect 2676 3727 2683 3913
rect 2716 3803 2723 4133
rect 2736 3827 2743 4353
rect 2756 4127 2763 4453
rect 2816 4243 2823 4476
rect 2796 4236 2823 4243
rect 2776 3987 2783 4213
rect 2796 4203 2803 4236
rect 2796 4196 2823 4203
rect 2836 4196 2863 4203
rect 2836 4107 2843 4196
rect 2896 4167 2903 4233
rect 2916 4207 2923 4513
rect 2936 4347 2943 4453
rect 2996 4447 3003 4473
rect 3016 4456 3023 4493
rect 2956 4287 2963 4443
rect 3036 4367 3043 4636
rect 3116 4456 3123 4513
rect 3136 4507 3143 4713
rect 3156 4707 3163 4896
rect 2996 4216 3003 4333
rect 2836 4087 2843 4093
rect 2816 4007 2823 4033
rect 2816 3976 2823 3993
rect 2756 3967 2763 3973
rect 2756 3943 2763 3953
rect 2756 3936 2783 3943
rect 2716 3796 2743 3803
rect 2696 3747 2703 3773
rect 2656 3643 2663 3703
rect 2696 3687 2703 3703
rect 2636 3636 2663 3643
rect 2556 3187 2563 3243
rect 2616 3167 2623 3223
rect 2516 3036 2523 3093
rect 2576 3067 2583 3113
rect 2496 2996 2523 3003
rect 2456 2507 2463 2713
rect 2476 2707 2483 2723
rect 2496 2707 2503 2743
rect 2476 2527 2483 2693
rect 2496 2547 2503 2693
rect 2516 2627 2523 2996
rect 2536 2603 2543 2993
rect 2576 2827 2583 3023
rect 2596 3007 2603 3133
rect 2636 3107 2643 3636
rect 2716 3487 2723 3693
rect 2736 3647 2743 3796
rect 2736 3507 2743 3613
rect 2656 3367 2663 3473
rect 2756 3347 2763 3853
rect 2656 3207 2663 3273
rect 2636 3087 2643 3093
rect 2656 3047 2663 3173
rect 2676 3087 2683 3293
rect 2716 3236 2723 3253
rect 2756 3247 2763 3313
rect 2776 3287 2783 3936
rect 2796 3687 2803 3733
rect 2816 3716 2823 3793
rect 2836 3767 2843 3963
rect 2836 3727 2843 3753
rect 2856 3516 2863 4133
rect 2876 4047 2883 4153
rect 2876 3947 2883 4013
rect 2916 4003 2923 4193
rect 2896 3996 2923 4003
rect 2896 3843 2903 3996
rect 2956 3987 2963 4113
rect 2976 4067 2983 4203
rect 3016 4043 3023 4233
rect 3036 4187 3043 4333
rect 3096 4203 3103 4443
rect 3136 4436 3143 4493
rect 3156 4456 3163 4693
rect 3176 4667 3183 4873
rect 3196 4747 3203 4956
rect 3236 4727 3243 4973
rect 3256 4936 3263 5156
rect 3276 4956 3283 5013
rect 3316 4987 3323 5403
rect 3336 5387 3343 5413
rect 3376 5403 3383 5433
rect 3376 5396 3403 5403
rect 3496 5267 3503 5456
rect 3536 5447 3543 5473
rect 3556 5467 3563 5643
rect 3736 5636 3763 5643
rect 3556 5187 3563 5213
rect 3376 5127 3383 5143
rect 3396 5023 3403 5123
rect 3376 5016 3403 5023
rect 3376 4967 3383 5016
rect 3416 5007 3423 5143
rect 3516 5127 3523 5163
rect 3556 5156 3563 5173
rect 3596 5143 3603 5433
rect 3396 4956 3403 4993
rect 3516 4976 3523 4993
rect 3536 4987 3543 5143
rect 3576 5136 3603 5143
rect 3376 4947 3383 4953
rect 3296 4887 3303 4943
rect 3436 4907 3443 4933
rect 3236 4696 3243 4713
rect 3316 4696 3323 4853
rect 3056 4196 3083 4203
rect 3096 4196 3123 4203
rect 3056 4107 3063 4196
rect 3096 4156 3113 4163
rect 2996 4036 3023 4043
rect 2996 4027 3003 4036
rect 3076 4023 3083 4113
rect 3056 4016 3083 4023
rect 2956 3887 2963 3933
rect 2996 3927 3003 3973
rect 3036 3967 3043 4013
rect 3056 3947 3063 4016
rect 2876 3836 2903 3843
rect 2876 3527 2883 3836
rect 2956 3716 2963 3793
rect 2996 3707 3003 3893
rect 2976 3687 2983 3703
rect 2836 3487 2843 3503
rect 2856 3387 2863 3473
rect 2796 3263 2803 3333
rect 2876 3307 2883 3493
rect 2776 3256 2803 3263
rect 2776 3203 2783 3256
rect 2836 3247 2843 3263
rect 2876 3256 2883 3293
rect 2796 3227 2803 3233
rect 2776 3196 2803 3203
rect 2696 3036 2703 3113
rect 2676 3007 2683 3023
rect 2576 2743 2583 2813
rect 2596 2776 2603 2913
rect 2676 2787 2683 2993
rect 2616 2743 2623 2763
rect 2576 2736 2623 2743
rect 2636 2623 2643 2773
rect 2696 2747 2703 2993
rect 2716 2987 2723 3023
rect 2616 2616 2643 2623
rect 2616 2607 2623 2616
rect 2516 2596 2543 2603
rect 2436 2263 2443 2493
rect 2496 2487 2503 2513
rect 2516 2367 2523 2596
rect 2556 2536 2563 2573
rect 2576 2556 2583 2593
rect 2596 2487 2603 2533
rect 2476 2296 2503 2303
rect 2436 2256 2463 2263
rect 2356 2196 2383 2203
rect 2316 2056 2343 2063
rect 2256 1967 2263 2043
rect 2236 1707 2243 1793
rect 2256 1663 2263 1813
rect 2296 1763 2303 1993
rect 2336 1947 2343 2056
rect 2356 2027 2363 2063
rect 2376 2007 2383 2196
rect 2416 1907 2423 2093
rect 2436 2056 2443 2153
rect 2456 1963 2463 2256
rect 2476 2067 2483 2296
rect 2516 2187 2523 2353
rect 2536 2287 2543 2393
rect 2556 2187 2563 2413
rect 2636 2403 2643 2593
rect 2616 2396 2643 2403
rect 2596 2227 2603 2263
rect 2616 2243 2623 2396
rect 2656 2307 2663 2713
rect 2696 2583 2703 2733
rect 2716 2587 2723 2953
rect 2756 2807 2763 3113
rect 2776 3047 2783 3073
rect 2796 3003 2803 3196
rect 2836 3023 2843 3213
rect 2856 3207 2863 3243
rect 2856 3176 2873 3183
rect 2856 3147 2863 3176
rect 2876 3056 2883 3073
rect 2816 3016 2843 3023
rect 2796 2996 2823 3003
rect 2776 2743 2783 2853
rect 2736 2707 2743 2743
rect 2776 2736 2803 2743
rect 2816 2723 2823 2996
rect 2836 2767 2843 2793
rect 2796 2716 2823 2723
rect 2676 2576 2703 2583
rect 2676 2567 2683 2576
rect 2696 2487 2703 2543
rect 2736 2536 2763 2543
rect 2716 2303 2723 2513
rect 2756 2507 2763 2536
rect 2776 2447 2783 2573
rect 2796 2307 2803 2716
rect 2816 2607 2823 2693
rect 2836 2583 2843 2733
rect 2816 2576 2843 2583
rect 2856 2583 2863 2873
rect 2876 2867 2883 3013
rect 2896 2967 2903 3573
rect 2936 3523 2943 3653
rect 2936 3516 2963 3523
rect 2996 3516 3003 3533
rect 2916 3387 2923 3413
rect 2916 3247 2923 3293
rect 2936 3267 2943 3516
rect 3016 3467 3023 3893
rect 3076 3767 3083 3983
rect 3116 3847 3123 4153
rect 3136 4127 3143 4183
rect 3156 4127 3163 4373
rect 3136 3847 3143 4033
rect 3036 3547 3043 3693
rect 3056 3547 3063 3723
rect 3116 3707 3123 3793
rect 3076 3607 3083 3653
rect 3036 3327 3043 3533
rect 3056 3507 3063 3513
rect 3096 3496 3103 3593
rect 3056 3483 3063 3493
rect 3056 3476 3083 3483
rect 3116 3467 3123 3483
rect 2936 3243 2943 3253
rect 2936 3236 2963 3243
rect 2976 3227 2983 3263
rect 3016 3256 3043 3263
rect 2936 3187 2943 3213
rect 2996 3203 3003 3243
rect 2976 3196 3003 3203
rect 2896 2756 2903 2873
rect 2916 2807 2923 3173
rect 2936 3036 2943 3073
rect 2976 3067 2983 3196
rect 2987 3036 3003 3043
rect 2956 2763 2963 2833
rect 2936 2756 2963 2763
rect 2876 2727 2883 2743
rect 2856 2576 2883 2583
rect 2816 2547 2823 2576
rect 2916 2543 2923 2713
rect 2936 2547 2943 2673
rect 2896 2536 2923 2543
rect 2716 2296 2743 2303
rect 2736 2276 2743 2296
rect 2716 2247 2723 2263
rect 2616 2236 2643 2243
rect 2616 2096 2623 2113
rect 2616 1967 2623 2053
rect 2456 1956 2483 1963
rect 2196 1556 2223 1563
rect 2236 1656 2263 1663
rect 2276 1756 2303 1763
rect 2236 1387 2243 1656
rect 2256 1587 2263 1633
rect 2216 1307 2223 1323
rect 2176 1296 2203 1303
rect 2176 1096 2183 1113
rect 2196 1087 2203 1296
rect 2256 1147 2263 1313
rect 2276 1267 2283 1756
rect 2476 1707 2483 1956
rect 2556 1767 2563 1893
rect 2336 1596 2343 1613
rect 2396 1543 2403 1693
rect 2416 1563 2423 1593
rect 2496 1563 2503 1633
rect 2416 1556 2443 1563
rect 2476 1556 2503 1563
rect 2436 1547 2443 1556
rect 2396 1536 2423 1543
rect 2296 1347 2303 1433
rect 2316 1336 2343 1343
rect 2316 1287 2323 1336
rect 2356 1307 2363 1323
rect 2216 1096 2223 1133
rect 2316 1127 2323 1193
rect 2316 1096 2323 1113
rect 2336 1107 2343 1273
rect 2356 1267 2363 1293
rect 2376 1247 2383 1333
rect 2136 836 2143 853
rect 2116 807 2123 823
rect 2176 687 2183 843
rect 2116 636 2123 653
rect 2176 623 2183 673
rect 2176 616 2203 623
rect 1856 343 1863 373
rect 1856 336 1883 343
rect 1996 323 2003 373
rect 1896 187 1903 323
rect 1996 316 2023 323
rect 1916 136 1923 153
rect 2076 127 2083 493
rect 2176 356 2183 573
rect 2216 383 2223 893
rect 2236 823 2243 913
rect 2276 887 2283 1093
rect 2296 927 2303 1083
rect 2336 1076 2343 1093
rect 2296 863 2303 893
rect 2276 856 2303 863
rect 2236 816 2263 823
rect 2256 667 2263 816
rect 2276 647 2283 856
rect 2316 807 2323 823
rect 2376 707 2383 1113
rect 2396 1107 2403 1313
rect 2416 1063 2423 1536
rect 2516 1543 2523 1673
rect 2496 1536 2523 1543
rect 2496 1323 2503 1536
rect 2536 1483 2543 1613
rect 2576 1576 2583 1733
rect 2596 1727 2603 1933
rect 2616 1847 2623 1953
rect 2616 1816 2623 1833
rect 2636 1787 2643 2236
rect 2716 1947 2723 2213
rect 2756 2107 2763 2263
rect 2776 2207 2783 2253
rect 2736 2056 2763 2063
rect 2756 1923 2763 2056
rect 2776 1967 2783 2043
rect 2756 1916 2773 1923
rect 2656 1807 2663 1913
rect 2696 1823 2703 1893
rect 2796 1887 2803 2293
rect 2816 1887 2823 2513
rect 2836 2287 2843 2393
rect 2876 2276 2883 2533
rect 2856 2227 2863 2263
rect 2916 2247 2923 2283
rect 2856 2083 2863 2093
rect 2836 2076 2863 2083
rect 2896 2076 2903 2113
rect 2916 2107 2923 2233
rect 2836 2027 2843 2076
rect 2756 1823 2763 1833
rect 2676 1816 2703 1823
rect 2736 1816 2763 1823
rect 2636 1596 2663 1603
rect 2476 1316 2503 1323
rect 2496 1187 2503 1316
rect 2516 1476 2543 1483
rect 2516 1243 2523 1476
rect 2536 1287 2543 1453
rect 2556 1307 2563 1393
rect 2596 1363 2603 1413
rect 2616 1407 2623 1583
rect 2656 1527 2663 1596
rect 2576 1356 2603 1363
rect 2576 1323 2583 1356
rect 2576 1316 2603 1323
rect 2636 1316 2643 1353
rect 2676 1327 2683 1816
rect 2516 1236 2543 1243
rect 2436 1096 2443 1133
rect 2496 1116 2503 1173
rect 2416 1056 2443 1063
rect 2416 836 2423 1033
rect 2436 827 2443 1056
rect 2516 1047 2523 1213
rect 2536 1107 2543 1236
rect 2556 1083 2563 1133
rect 2596 1096 2603 1113
rect 2556 1076 2583 1083
rect 2556 907 2563 1076
rect 2556 856 2583 863
rect 2576 847 2583 856
rect 2396 643 2403 803
rect 2296 636 2323 643
rect 2376 636 2403 643
rect 2296 507 2303 636
rect 2436 603 2443 753
rect 2436 596 2463 603
rect 2216 376 2243 383
rect 2216 343 2223 353
rect 2156 167 2163 343
rect 2196 336 2223 343
rect 2176 187 2183 193
rect 2116 136 2123 153
rect 2176 143 2183 173
rect 2236 163 2243 376
rect 2256 187 2263 413
rect 2336 356 2343 533
rect 2356 327 2363 393
rect 2456 347 2463 596
rect 2496 567 2503 603
rect 2536 427 2543 843
rect 2636 836 2643 853
rect 2656 767 2663 1303
rect 2676 1107 2683 1313
rect 2696 1207 2703 1753
rect 2716 1747 2723 1803
rect 2756 1767 2763 1816
rect 2716 1627 2723 1733
rect 2776 1607 2783 1813
rect 2796 1807 2803 1873
rect 2816 1767 2823 1853
rect 2896 1787 2903 1803
rect 2916 1747 2923 1993
rect 2756 1547 2763 1563
rect 2796 1547 2803 1613
rect 2736 1327 2743 1413
rect 2756 1336 2803 1343
rect 2756 1316 2763 1336
rect 2716 1187 2723 1273
rect 2736 1227 2743 1283
rect 2716 1136 2723 1173
rect 2756 1127 2763 1193
rect 2756 863 2763 1113
rect 2776 1107 2783 1273
rect 2796 1227 2803 1336
rect 2816 1307 2823 1713
rect 2856 1596 2863 1633
rect 2896 1596 2903 1653
rect 2836 1576 2843 1593
rect 2836 1307 2843 1393
rect 2856 1387 2863 1513
rect 2876 1407 2883 1583
rect 2916 1547 2923 1713
rect 2936 1427 2943 2213
rect 2956 2127 2963 2756
rect 2976 2607 2983 2913
rect 2996 2787 3003 3036
rect 2996 2607 3003 2713
rect 2996 2576 3003 2593
rect 3016 2543 3023 3213
rect 3036 3207 3043 3256
rect 3056 3227 3063 3453
rect 3036 2827 3043 3113
rect 3076 3047 3083 3273
rect 3096 3187 3103 3393
rect 3136 3347 3143 3673
rect 3156 3407 3163 4053
rect 3176 4027 3183 4633
rect 3216 4567 3223 4683
rect 3256 4647 3263 4673
rect 3356 4627 3363 4703
rect 3396 4683 3403 4773
rect 3416 4687 3423 4713
rect 3376 4676 3403 4683
rect 3216 4547 3223 4553
rect 3236 4207 3243 4463
rect 3196 4196 3223 4203
rect 3196 4107 3203 4196
rect 3256 4196 3263 4533
rect 3216 4083 3223 4113
rect 3196 4076 3223 4083
rect 3196 3976 3203 4076
rect 3176 3587 3183 3963
rect 3216 3956 3223 4053
rect 3236 3976 3243 4113
rect 3276 4003 3283 4093
rect 3296 4047 3303 4593
rect 3316 4476 3323 4493
rect 3336 4447 3343 4463
rect 3376 4456 3383 4473
rect 3316 4103 3323 4273
rect 3336 4167 3343 4393
rect 3316 4096 3343 4103
rect 3336 4087 3343 4096
rect 3316 4027 3323 4073
rect 3336 4016 3343 4053
rect 3276 3996 3303 4003
rect 3256 3967 3263 3993
rect 3236 3847 3243 3873
rect 3196 3736 3203 3753
rect 3256 3647 3263 3833
rect 3276 3663 3283 3973
rect 3296 3827 3303 3996
rect 3296 3687 3303 3753
rect 3316 3716 3323 3733
rect 3336 3727 3343 3813
rect 3356 3807 3363 4033
rect 3376 3847 3383 4153
rect 3396 4107 3403 4183
rect 3436 4107 3443 4793
rect 3456 4767 3463 4943
rect 3476 4707 3483 4753
rect 3476 4676 3483 4693
rect 3496 4687 3503 4973
rect 3556 4963 3563 5113
rect 3536 4956 3563 4963
rect 3516 4683 3523 4913
rect 3556 4867 3563 4956
rect 3576 4927 3583 4943
rect 3616 4907 3623 5573
rect 3736 5547 3743 5636
rect 3936 5607 3943 5623
rect 3776 5587 3783 5603
rect 3716 5427 3723 5533
rect 3736 5447 3743 5533
rect 3636 5176 3643 5193
rect 3676 5176 3693 5183
rect 3656 5147 3663 5163
rect 3696 4976 3703 5173
rect 3656 4956 3683 4963
rect 3716 4956 3723 5093
rect 3516 4676 3543 4683
rect 3536 4667 3543 4676
rect 3456 4647 3463 4663
rect 3456 4207 3463 4513
rect 3476 4476 3483 4513
rect 3516 4443 3523 4493
rect 3496 4436 3523 4443
rect 3516 4407 3523 4436
rect 3396 3787 3403 4073
rect 3476 3996 3483 4153
rect 3496 4127 3503 4193
rect 3556 4167 3563 4453
rect 3576 4247 3583 4893
rect 3656 4747 3663 4956
rect 3596 4696 3603 4713
rect 3636 4687 3643 4703
rect 3616 4667 3623 4683
rect 3636 4647 3643 4673
rect 3656 4527 3663 4593
rect 3596 4447 3603 4473
rect 3636 4456 3643 4473
rect 3616 4407 3623 4443
rect 3636 4387 3643 4413
rect 3456 3947 3463 3983
rect 3496 3963 3503 4093
rect 3556 3976 3563 4053
rect 3576 4047 3583 4233
rect 3596 4203 3603 4253
rect 3676 4227 3683 4853
rect 3696 4487 3703 4813
rect 3716 4663 3723 4873
rect 3756 4707 3763 5493
rect 3776 5387 3783 5493
rect 3796 5427 3803 5513
rect 3836 5467 3843 5603
rect 3947 5596 3963 5603
rect 3956 5527 3963 5596
rect 3976 5567 3983 5623
rect 3996 5607 4003 5643
rect 4096 5636 4103 5653
rect 4576 5636 4603 5643
rect 4736 5636 4743 5653
rect 4836 5636 4843 5673
rect 4136 5616 4163 5623
rect 3976 5507 3983 5533
rect 3856 5456 3863 5493
rect 3896 5423 3903 5433
rect 3876 5416 3903 5423
rect 3816 5176 3843 5183
rect 3836 5047 3843 5176
rect 3836 5007 3843 5033
rect 3856 5003 3863 5413
rect 3876 5407 3883 5416
rect 3916 5403 3923 5473
rect 3956 5416 3963 5493
rect 3916 5396 3943 5403
rect 3896 5167 3903 5393
rect 3976 5267 3983 5403
rect 3996 5387 4003 5593
rect 4136 5587 4143 5616
rect 4236 5607 4243 5623
rect 4516 5567 4523 5623
rect 4136 5436 4153 5443
rect 4056 5416 4083 5423
rect 4056 5367 4063 5416
rect 4156 5407 4163 5433
rect 3956 5176 3963 5193
rect 3856 4996 3883 5003
rect 3776 4923 3783 4993
rect 3856 4936 3863 4973
rect 3776 4916 3803 4923
rect 3796 4807 3803 4916
rect 3876 4827 3883 4996
rect 3916 4943 3923 5093
rect 3936 5067 3943 5163
rect 3916 4936 3943 4943
rect 3796 4676 3803 4693
rect 3716 4656 3743 4663
rect 3816 4647 3823 4713
rect 3696 4447 3703 4473
rect 3596 4196 3623 4203
rect 3636 4187 3643 4223
rect 3476 3956 3503 3963
rect 3356 3747 3363 3773
rect 3276 3656 3303 3663
rect 3196 3487 3203 3513
rect 3256 3467 3263 3493
rect 3276 3443 3283 3633
rect 3256 3436 3283 3443
rect 3116 3256 3123 3333
rect 3156 3283 3163 3313
rect 3156 3276 3183 3283
rect 3136 3167 3143 3243
rect 3096 3016 3103 3153
rect 3116 2987 3123 3003
rect 3136 2927 3143 3033
rect 3156 2987 3163 3073
rect 3116 2787 3123 2813
rect 3036 2547 3043 2733
rect 3056 2687 3063 2763
rect 3096 2747 3103 2763
rect 3136 2747 3143 2873
rect 3176 2807 3183 3276
rect 3196 3167 3203 3333
rect 3236 3267 3243 3333
rect 3256 3256 3263 3436
rect 3296 3347 3303 3656
rect 3316 3407 3323 3573
rect 3376 3503 3383 3753
rect 3396 3587 3403 3723
rect 3396 3527 3403 3533
rect 3376 3496 3403 3503
rect 3416 3467 3423 3533
rect 3476 3523 3483 3956
rect 3496 3547 3503 3913
rect 3516 3547 3523 3813
rect 3556 3716 3563 3753
rect 3536 3587 3543 3683
rect 3476 3516 3503 3523
rect 3536 3516 3543 3573
rect 3556 3567 3563 3673
rect 3296 3256 3303 3273
rect 3276 3147 3283 3243
rect 3216 3036 3223 3113
rect 3256 3003 3263 3053
rect 3276 3036 3283 3073
rect 3247 2996 3263 3003
rect 3296 2847 3303 2933
rect 3196 2776 3203 2793
rect 3176 2667 3183 2763
rect 3056 2576 3123 2583
rect 3056 2556 3063 2576
rect 3116 2567 3123 2576
rect 2996 2536 3023 2543
rect 2976 2327 2983 2533
rect 2956 2007 2963 2113
rect 2996 2007 3003 2536
rect 3076 2467 3083 2543
rect 3116 2536 3143 2543
rect 3016 2307 3023 2413
rect 3056 2296 3063 2313
rect 3036 2147 3043 2253
rect 3016 1983 3023 2043
rect 3056 2027 3063 2043
rect 3056 2007 3063 2013
rect 2996 1976 3023 1983
rect 2996 1867 3003 1976
rect 3016 1796 3023 1933
rect 3036 1827 3043 1993
rect 2916 1367 2923 1373
rect 2856 1287 2863 1353
rect 2916 1316 2923 1353
rect 2816 1116 2823 1173
rect 2836 1136 2843 1273
rect 2936 1143 2943 1303
rect 2956 1187 2963 1773
rect 2996 1767 3003 1783
rect 3036 1767 3043 1783
rect 2996 1596 3003 1633
rect 3056 1627 3063 1993
rect 3076 1763 3083 1953
rect 3096 1827 3103 2373
rect 3136 2303 3143 2536
rect 3156 2527 3163 2553
rect 3176 2507 3183 2573
rect 3196 2567 3203 2593
rect 3216 2587 3223 2773
rect 3236 2747 3243 2793
rect 3256 2727 3263 2793
rect 3276 2763 3283 2833
rect 3316 2787 3323 3313
rect 3336 3227 3343 3453
rect 3356 3367 3363 3453
rect 3416 3367 3423 3433
rect 3336 3056 3343 3113
rect 3356 3036 3363 3153
rect 3396 3087 3403 3253
rect 3376 2947 3383 3033
rect 3276 2756 3303 2763
rect 3356 2727 3363 2743
rect 3236 2536 3243 2593
rect 3196 2487 3203 2533
rect 3276 2527 3283 2553
rect 3196 2367 3203 2413
rect 3116 2296 3143 2303
rect 3176 2296 3183 2333
rect 3116 2247 3123 2296
rect 3156 2247 3163 2283
rect 3196 2267 3203 2333
rect 3216 2267 3223 2493
rect 3296 2467 3303 2673
rect 3207 2236 3213 2243
rect 3136 2056 3143 2173
rect 3176 2043 3183 2093
rect 3116 1827 3123 2043
rect 3156 2036 3183 2043
rect 3076 1756 3103 1763
rect 3036 1596 3043 1613
rect 3076 1603 3083 1733
rect 3056 1596 3083 1603
rect 2976 1307 2983 1533
rect 3016 1527 3023 1583
rect 2996 1203 3003 1353
rect 3036 1343 3043 1373
rect 3056 1367 3063 1596
rect 3096 1563 3103 1756
rect 3136 1683 3143 1783
rect 3116 1676 3143 1683
rect 3116 1607 3123 1676
rect 3156 1663 3163 1873
rect 3176 1727 3183 1933
rect 3196 1687 3203 2033
rect 3216 1807 3223 2073
rect 3236 2067 3243 2353
rect 3256 2307 3263 2393
rect 3316 2307 3323 2673
rect 3376 2667 3383 2773
rect 3396 2687 3403 2993
rect 3416 2787 3423 3353
rect 3436 3187 3443 3513
rect 3456 3427 3463 3473
rect 3496 3447 3503 3473
rect 3556 3387 3563 3553
rect 3576 3327 3583 3733
rect 3596 3463 3603 4173
rect 3656 4167 3663 4203
rect 3616 3687 3623 4153
rect 3716 4087 3723 4593
rect 3736 4187 3743 4633
rect 3776 4627 3783 4643
rect 3816 4496 3823 4553
rect 3816 4216 3823 4453
rect 3836 4207 3843 4693
rect 3876 4663 3883 4703
rect 3916 4696 3923 4773
rect 3867 4656 3883 4663
rect 3856 4467 3863 4653
rect 3896 4647 3903 4683
rect 3896 4627 3903 4633
rect 3936 4607 3943 4936
rect 3976 4867 3983 5193
rect 4076 5176 4083 5353
rect 4016 5156 4043 5163
rect 3996 5087 4003 5153
rect 4016 5127 4023 5133
rect 4016 4936 4023 4973
rect 4036 4927 4043 5156
rect 4056 4936 4063 4953
rect 3956 4707 3963 4793
rect 3896 4456 3903 4493
rect 3936 4443 3943 4553
rect 3916 4436 3943 4443
rect 3916 4227 3923 4253
rect 3976 4247 3983 4853
rect 4056 4696 4083 4703
rect 3996 4667 4003 4683
rect 3956 4216 3983 4223
rect 3756 4196 3783 4203
rect 3636 3807 3643 4073
rect 3716 3996 3723 4053
rect 3736 4016 3743 4073
rect 3776 4047 3783 4196
rect 3976 4187 3983 4216
rect 3996 4167 4003 4653
rect 4036 4607 4043 4683
rect 4076 4647 4083 4696
rect 4016 4476 4023 4493
rect 4036 4447 4043 4593
rect 4096 4527 4103 5053
rect 4136 5027 4143 5373
rect 4216 5367 4223 5403
rect 4316 5403 4323 5453
rect 4376 5407 4383 5453
rect 4396 5416 4423 5423
rect 4416 5407 4423 5416
rect 4316 5396 4343 5403
rect 4176 5127 4183 5163
rect 4256 5147 4263 5173
rect 4116 4927 4123 4953
rect 4136 4943 4143 4973
rect 4176 4967 4183 5113
rect 4236 5047 4243 5143
rect 4136 4936 4163 4943
rect 4136 4903 4143 4936
rect 4116 4896 4143 4903
rect 4116 4547 4123 4896
rect 4156 4676 4163 4753
rect 4176 4687 4183 4693
rect 4176 4647 4183 4673
rect 4236 4607 4243 5013
rect 4276 4967 4283 5333
rect 4296 5103 4303 5153
rect 4376 5147 4383 5163
rect 4316 5127 4323 5143
rect 4296 5096 4323 5103
rect 4316 4956 4323 5096
rect 4376 4963 4383 4973
rect 4356 4956 4383 4963
rect 4276 4887 4283 4893
rect 4276 4727 4283 4873
rect 4276 4696 4283 4713
rect 4296 4687 4303 4953
rect 4356 4927 4363 4956
rect 4336 4827 4343 4923
rect 4256 4627 4263 4663
rect 4056 4476 4063 4513
rect 4116 4507 4123 4533
rect 4116 4476 4123 4493
rect 4176 4476 4203 4483
rect 4036 4263 4043 4433
rect 4156 4427 4163 4443
rect 4036 4256 4063 4263
rect 3676 3967 3683 3983
rect 3636 3707 3643 3793
rect 3716 3747 3723 3933
rect 3616 3496 3623 3573
rect 3636 3516 3643 3613
rect 3656 3567 3663 3703
rect 3676 3647 3683 3683
rect 3676 3516 3683 3613
rect 3596 3456 3623 3463
rect 3596 3303 3603 3393
rect 3576 3296 3603 3303
rect 3436 3127 3443 3173
rect 3456 3007 3463 3273
rect 3436 2787 3443 2953
rect 3476 2807 3483 3133
rect 3496 3047 3503 3243
rect 3516 3167 3523 3263
rect 3536 3143 3543 3213
rect 3516 3136 3543 3143
rect 3516 3036 3523 3136
rect 3556 3047 3563 3193
rect 3576 3147 3583 3296
rect 3616 3287 3623 3456
rect 3676 3267 3683 3453
rect 3696 3427 3703 3533
rect 3696 3227 3703 3393
rect 3616 3167 3623 3203
rect 3496 3016 3503 3033
rect 3536 3007 3543 3023
rect 3516 2823 3523 2993
rect 3516 2816 3543 2823
rect 3456 2776 3483 2783
rect 3336 2487 3343 2653
rect 3376 2536 3383 2553
rect 3416 2536 3423 2713
rect 3287 2296 3293 2303
rect 3336 2276 3343 2353
rect 3256 2187 3263 2273
rect 3316 2227 3323 2243
rect 3356 2187 3363 2493
rect 3436 2467 3443 2513
rect 3376 2327 3383 2353
rect 3396 2307 3403 2433
rect 3296 2076 3303 2113
rect 3236 1667 3243 1783
rect 3256 1727 3263 1973
rect 3276 1796 3283 2053
rect 3316 2047 3323 2113
rect 3336 2047 3343 2173
rect 3296 1747 3303 1773
rect 3316 1687 3323 1813
rect 3356 1787 3363 2093
rect 3376 1847 3383 2293
rect 3416 2287 3423 2433
rect 3456 2387 3463 2693
rect 3476 2687 3483 2776
rect 3516 2747 3523 2793
rect 3496 2736 3513 2743
rect 3476 2567 3483 2653
rect 3456 2263 3463 2353
rect 3476 2327 3483 2473
rect 3396 2227 3403 2263
rect 3436 2256 3463 2263
rect 3416 2187 3423 2243
rect 3396 2076 3403 2173
rect 3416 1827 3423 2043
rect 3136 1656 3163 1663
rect 3076 1556 3103 1563
rect 3116 1407 3123 1533
rect 3136 1527 3143 1656
rect 3216 1423 3223 1653
rect 3236 1616 3243 1633
rect 3236 1447 3243 1573
rect 3376 1523 3383 1813
rect 3396 1543 3403 1753
rect 3416 1707 3423 1763
rect 3436 1583 3443 2153
rect 3476 2127 3483 2313
rect 3496 2267 3503 2713
rect 3536 2667 3543 2816
rect 3616 2747 3623 3133
rect 3696 3127 3703 3193
rect 3656 3036 3663 3053
rect 3696 3036 3703 3113
rect 3636 3016 3643 3033
rect 3676 3007 3683 3023
rect 3716 2847 3723 3733
rect 3736 3667 3743 3713
rect 3756 3543 3763 3993
rect 3776 3927 3783 4033
rect 3796 3963 3803 4053
rect 3876 3963 3883 4073
rect 3796 3956 3823 3963
rect 3856 3956 3883 3963
rect 3816 3736 3823 3833
rect 3796 3683 3803 3723
rect 3776 3676 3803 3683
rect 3776 3587 3783 3676
rect 3836 3667 3843 3753
rect 3736 3536 3763 3543
rect 3736 2823 3743 3536
rect 3796 3467 3803 3653
rect 3816 3516 3843 3523
rect 3836 3507 3843 3516
rect 3756 3067 3763 3243
rect 3796 3236 3803 3453
rect 3836 3407 3843 3493
rect 3836 3227 3843 3233
rect 3776 3167 3783 3223
rect 3816 3216 3833 3223
rect 3736 2816 3763 2823
rect 3556 2687 3563 2743
rect 3536 2556 3563 2563
rect 3516 2507 3523 2523
rect 3416 1576 3443 1583
rect 3396 1536 3423 1543
rect 3376 1516 3403 1523
rect 3216 1416 3243 1423
rect 3036 1336 3063 1343
rect 3056 1316 3063 1336
rect 3196 1316 3203 1353
rect 2976 1196 3023 1203
rect 2916 1136 2943 1143
rect 2856 1116 2883 1123
rect 2876 1047 2883 1116
rect 2896 867 2903 1113
rect 2916 987 2923 1136
rect 2976 1116 2983 1196
rect 2976 947 2983 1073
rect 2736 856 2763 863
rect 2796 856 2823 863
rect 2736 827 2743 856
rect 2696 787 2703 803
rect 2816 787 2823 856
rect 2936 856 2943 873
rect 2696 636 2723 643
rect 2756 636 2783 643
rect 2596 547 2603 603
rect 2636 527 2643 603
rect 2696 547 2703 636
rect 2496 376 2523 383
rect 2216 156 2243 163
rect 2256 156 2283 163
rect 2156 136 2183 143
rect 1796 116 1823 123
rect 1856 107 1863 123
rect 2096 107 2103 123
rect 2276 47 2283 156
rect 2336 123 2343 153
rect 2376 136 2383 293
rect 2496 163 2503 376
rect 2596 363 2603 433
rect 2636 407 2643 513
rect 2576 356 2603 363
rect 2656 356 2663 453
rect 2576 327 2583 356
rect 2696 347 2703 363
rect 2636 307 2643 343
rect 2716 207 2723 393
rect 2736 367 2743 613
rect 2776 527 2783 636
rect 2796 636 2823 643
rect 2856 636 2863 853
rect 2796 587 2803 636
rect 2876 616 2883 653
rect 2796 356 2803 513
rect 2916 467 2923 843
rect 2996 807 3003 1173
rect 3016 847 3023 1196
rect 3036 836 3043 1273
rect 3056 1116 3063 1133
rect 3076 1127 3083 1303
rect 3136 1067 3143 1293
rect 3176 1227 3183 1303
rect 3156 1087 3163 1153
rect 2476 156 2503 163
rect 2516 156 2523 193
rect 2476 127 2483 156
rect 2716 147 2723 193
rect 2756 156 2763 333
rect 2836 327 2843 413
rect 2876 347 2883 373
rect 2896 327 2903 343
rect 2816 316 2833 323
rect 2816 156 2843 163
rect 2836 147 2843 156
rect 2916 136 2923 153
rect 2336 116 2363 123
rect 2487 116 2503 123
rect 2776 107 2783 123
rect 2896 107 2903 123
rect 2636 -24 2643 13
rect 2676 -24 2683 33
rect 2956 27 2963 793
rect 3016 783 3023 803
rect 2996 776 3023 783
rect 2996 627 3003 776
rect 2976 107 2983 533
rect 2996 127 3003 313
rect 3036 187 3043 633
rect 3056 407 3063 833
rect 3116 807 3123 873
rect 3096 343 3103 573
rect 3156 547 3163 633
rect 3176 627 3183 833
rect 3196 667 3203 1233
rect 3216 1187 3223 1303
rect 3216 1116 3223 1173
rect 3236 1136 3243 1416
rect 3256 1147 3263 1473
rect 3276 1287 3283 1473
rect 3296 1316 3303 1393
rect 3396 1316 3403 1516
rect 3416 1307 3423 1536
rect 3436 1507 3443 1553
rect 3376 1247 3383 1283
rect 3376 1136 3383 1153
rect 3256 1116 3283 1123
rect 3236 643 3243 1093
rect 3276 1067 3283 1116
rect 3336 1116 3363 1123
rect 3396 1116 3403 1133
rect 3256 856 3263 913
rect 3276 787 3283 843
rect 3316 647 3323 1113
rect 3336 1047 3343 1116
rect 3336 807 3343 1033
rect 3416 847 3423 1213
rect 3436 1207 3443 1493
rect 3456 1467 3463 1973
rect 3496 1927 3503 2233
rect 3516 2207 3523 2373
rect 3556 2276 3563 2556
rect 3576 2487 3583 2653
rect 3596 2503 3603 2693
rect 3636 2536 3643 2673
rect 3656 2567 3663 2793
rect 3736 2776 3743 2793
rect 3756 2767 3763 2816
rect 3676 2747 3683 2763
rect 3596 2496 3623 2503
rect 3576 2307 3583 2473
rect 3596 2187 3603 2283
rect 3576 2076 3583 2093
rect 3556 2047 3563 2053
rect 3616 2047 3623 2496
rect 3656 2487 3663 2523
rect 3676 2507 3683 2713
rect 3636 2267 3643 2373
rect 3656 2247 3663 2373
rect 3676 2296 3683 2393
rect 3696 2387 3703 2673
rect 3736 2587 3743 2733
rect 3756 2587 3763 2753
rect 3716 2563 3723 2573
rect 3716 2556 3743 2563
rect 3776 2556 3783 2733
rect 3796 2707 3803 3153
rect 3836 3003 3843 3013
rect 3816 2996 3843 3003
rect 3816 2947 3823 2996
rect 3836 2803 3843 2893
rect 3856 2827 3863 3933
rect 3896 3827 3903 4033
rect 3916 3716 3923 3773
rect 3896 3647 3903 3683
rect 3876 3527 3883 3593
rect 3896 3536 3903 3613
rect 3916 3207 3923 3373
rect 3876 3087 3883 3193
rect 3876 2987 3883 3033
rect 3896 3007 3903 3033
rect 3836 2796 3863 2803
rect 3856 2776 3863 2796
rect 3836 2647 3843 2763
rect 3816 2556 3823 2573
rect 3716 2447 3723 2533
rect 3756 2527 3763 2543
rect 3736 2303 3743 2513
rect 3716 2296 3743 2303
rect 3696 2267 3703 2283
rect 3496 1867 3503 1913
rect 3536 1796 3543 1913
rect 3476 1747 3483 1783
rect 3476 1567 3483 1693
rect 3456 1307 3463 1373
rect 3436 1027 3443 1133
rect 3436 787 3443 823
rect 3216 636 3243 643
rect 3176 467 3183 613
rect 3136 356 3143 413
rect 3216 407 3223 636
rect 3276 596 3283 633
rect 3156 367 3163 373
rect 3256 367 3263 553
rect 3316 427 3323 633
rect 3376 616 3383 653
rect 3296 356 3303 373
rect 3096 336 3123 343
rect 3316 223 3323 343
rect 3336 327 3343 613
rect 3416 603 3423 653
rect 3396 596 3423 603
rect 3356 567 3363 593
rect 3416 356 3423 393
rect 3456 367 3463 1273
rect 3476 1207 3483 1533
rect 3496 1387 3503 1583
rect 3516 1547 3523 1783
rect 3556 1687 3563 1783
rect 3536 1547 3543 1593
rect 3496 1227 3503 1303
rect 3496 1136 3503 1173
rect 3476 867 3483 1103
rect 3516 1007 3523 1513
rect 3536 1447 3543 1473
rect 3556 1167 3563 1613
rect 3576 1267 3583 1813
rect 3596 1627 3603 2013
rect 3636 1963 3643 2073
rect 3656 2027 3663 2213
rect 3676 2107 3683 2253
rect 3676 2076 3703 2083
rect 3676 2007 3683 2076
rect 3716 1987 3723 2033
rect 3616 1956 3643 1963
rect 3616 1907 3623 1956
rect 3616 1787 3623 1833
rect 3636 1767 3643 1933
rect 3656 1767 3663 1803
rect 3696 1796 3703 1893
rect 3656 1747 3663 1753
rect 3636 1616 3643 1713
rect 3676 1687 3683 1783
rect 3616 1567 3623 1583
rect 3596 1187 3603 1533
rect 3656 1407 3663 1573
rect 3676 1567 3683 1613
rect 3696 1587 3703 1713
rect 3736 1667 3743 2273
rect 3756 1647 3763 2353
rect 3776 2247 3783 2473
rect 3796 2307 3803 2513
rect 3816 2427 3823 2493
rect 3796 2207 3803 2263
rect 3816 2187 3823 2413
rect 3836 2307 3843 2613
rect 3856 2547 3863 2573
rect 3856 2347 3863 2513
rect 3836 2247 3843 2263
rect 3776 2047 3783 2173
rect 3836 2087 3843 2233
rect 3856 2223 3863 2333
rect 3876 2243 3883 2813
rect 3916 2707 3923 3173
rect 3936 3147 3943 3993
rect 4036 3967 4043 4233
rect 4056 4227 4063 4256
rect 4096 4216 4103 4233
rect 3996 3683 4003 3953
rect 4056 3683 4063 4173
rect 4076 4007 4083 4203
rect 4136 4067 4143 4213
rect 4156 4107 4163 4413
rect 4196 4267 4203 4476
rect 4236 4307 4243 4573
rect 4316 4547 4323 4663
rect 4176 4216 4183 4253
rect 4236 4223 4243 4293
rect 4216 4216 4243 4223
rect 4236 4187 4243 4216
rect 4096 3996 4103 4053
rect 4136 4016 4143 4033
rect 4176 3983 4183 4053
rect 4156 3976 4183 3983
rect 4196 3947 4203 4173
rect 4256 4047 4263 4473
rect 4316 4407 4323 4443
rect 4336 4407 4343 4673
rect 4276 4387 4283 4393
rect 4216 3947 4223 3963
rect 4256 3847 4263 3963
rect 3996 3676 4023 3683
rect 3976 3487 3983 3613
rect 3996 3527 4003 3633
rect 3956 3247 3963 3253
rect 3956 3216 3963 3233
rect 3996 3167 4003 3373
rect 4016 3367 4023 3676
rect 4036 3676 4063 3683
rect 4036 3627 4043 3676
rect 4136 3667 4143 3713
rect 4156 3607 4163 3703
rect 4196 3587 4203 3703
rect 4056 3516 4063 3533
rect 4096 3516 4123 3523
rect 4116 3507 4123 3516
rect 4076 3483 4083 3503
rect 4056 3476 4083 3483
rect 3956 2987 3963 3003
rect 3976 2807 3983 3133
rect 3996 3047 4003 3053
rect 4016 2907 4023 3253
rect 4036 3167 4043 3223
rect 4056 3067 4063 3476
rect 4076 3467 4083 3476
rect 4076 3187 4083 3223
rect 4076 3056 4083 3113
rect 4096 3067 4103 3233
rect 4047 3036 4063 3043
rect 4096 3036 4123 3043
rect 3936 2556 3943 2793
rect 3996 2787 4003 2793
rect 4016 2787 4023 2873
rect 3956 2647 3963 2743
rect 3996 2687 4003 2773
rect 3876 2236 3903 2243
rect 3856 2216 3883 2223
rect 3796 2056 3803 2073
rect 3876 2043 3883 2216
rect 3856 2036 3883 2043
rect 3776 1787 3783 2013
rect 3776 1747 3783 1773
rect 3756 1596 3763 1613
rect 3736 1547 3743 1573
rect 3796 1427 3803 1873
rect 3816 1767 3823 1803
rect 3856 1796 3863 1833
rect 3876 1767 3883 1783
rect 3856 1756 3873 1763
rect 3836 1443 3843 1593
rect 3856 1527 3863 1756
rect 3896 1707 3903 2236
rect 3916 2007 3923 2533
rect 3936 2063 3943 2493
rect 3976 2343 3983 2653
rect 3996 2367 4003 2543
rect 4016 2487 4023 2773
rect 4036 2527 4043 3033
rect 4116 2987 4123 3036
rect 4056 2707 4063 2763
rect 4076 2727 4083 2743
rect 4116 2727 4123 2743
rect 4136 2707 4143 3313
rect 4156 3047 4163 3333
rect 4176 3127 4183 3473
rect 4196 3247 4203 3553
rect 4216 3547 4223 3693
rect 4256 3563 4263 3833
rect 4276 3567 4283 4373
rect 4356 4223 4363 4453
rect 4376 4427 4383 4913
rect 4396 4487 4403 5073
rect 4416 4947 4423 5213
rect 4416 4727 4423 4933
rect 4436 4887 4443 5473
rect 4536 5436 4543 5513
rect 4556 5507 4563 5633
rect 4576 5607 4583 5636
rect 4576 5527 4583 5593
rect 4596 5456 4623 5463
rect 4596 5447 4603 5456
rect 4716 5436 4723 5493
rect 4756 5436 4763 5453
rect 4816 5443 4823 5593
rect 4816 5436 4843 5443
rect 4476 5367 4483 5413
rect 4516 5407 4523 5413
rect 4736 5407 4743 5423
rect 4776 5416 4803 5423
rect 4476 4956 4493 4963
rect 4496 4827 4503 4953
rect 4536 4943 4543 5133
rect 4516 4936 4543 4943
rect 4556 4927 4563 5393
rect 4796 5383 4803 5416
rect 4776 5376 4803 5383
rect 4576 5176 4583 5193
rect 4596 5147 4603 5163
rect 4616 5127 4623 5183
rect 4656 5047 4663 5133
rect 4616 4976 4623 5033
rect 4596 4956 4603 4973
rect 4676 4943 4683 5253
rect 4776 5143 4783 5376
rect 4756 5136 4783 5143
rect 4656 4936 4683 4943
rect 4616 4847 4623 4913
rect 4456 4647 4463 4703
rect 4476 4547 4483 4673
rect 4476 4483 4483 4513
rect 4456 4476 4483 4483
rect 4436 4447 4443 4463
rect 4476 4323 4483 4476
rect 4496 4447 4503 4713
rect 4536 4456 4543 4593
rect 4556 4587 4563 4703
rect 4596 4696 4603 4813
rect 4576 4667 4583 4683
rect 4476 4316 4503 4323
rect 4356 4216 4383 4223
rect 4296 4127 4303 4203
rect 4376 4183 4383 4216
rect 4356 4176 4383 4183
rect 4376 4167 4383 4176
rect 4396 4127 4403 4173
rect 4496 4147 4503 4316
rect 4556 4307 4563 4443
rect 4596 4347 4603 4633
rect 4616 4367 4623 4833
rect 4656 4623 4663 4936
rect 4696 4687 4703 4733
rect 4656 4616 4683 4623
rect 4676 4456 4683 4616
rect 4656 4403 4663 4443
rect 4696 4407 4703 4443
rect 4656 4396 4683 4403
rect 4596 4227 4603 4333
rect 4296 3603 4303 4093
rect 4336 4007 4343 4113
rect 4376 3996 4383 4033
rect 4456 3996 4483 4003
rect 4296 3596 4323 3603
rect 4236 3556 4263 3563
rect 4216 3327 4223 3533
rect 4236 3267 4243 3556
rect 4256 3516 4263 3533
rect 4296 3516 4303 3573
rect 4316 3527 4323 3596
rect 4336 3563 4343 3873
rect 4376 3727 4383 3873
rect 4416 3716 4423 3893
rect 4436 3747 4443 3973
rect 4456 3707 4463 3996
rect 4476 3743 4483 3913
rect 4496 3767 4503 3983
rect 4536 3976 4543 3993
rect 4556 3923 4563 4213
rect 4616 4207 4623 4293
rect 4576 4127 4583 4203
rect 4596 4023 4603 4183
rect 4636 4167 4643 4183
rect 4656 4167 4663 4353
rect 4676 4187 4683 4396
rect 4716 4243 4723 5033
rect 4756 4956 4763 5113
rect 4796 4956 4803 5353
rect 4836 5347 4843 5436
rect 4876 5347 4883 5653
rect 4836 5107 4843 5133
rect 4856 5087 4863 5123
rect 4896 5047 4903 5653
rect 4936 5607 4943 5643
rect 4976 5636 4983 5673
rect 5076 5663 5083 5773
rect 5136 5663 5143 5673
rect 5056 5656 5083 5663
rect 5116 5656 5143 5663
rect 5056 5627 5063 5656
rect 4916 5436 4923 5513
rect 4956 5436 4963 5623
rect 4996 5603 5003 5613
rect 5096 5607 5103 5643
rect 5136 5627 5143 5656
rect 4976 5596 5003 5603
rect 4916 5136 4943 5143
rect 4916 5067 4923 5136
rect 4816 4956 4843 4963
rect 4736 4936 4743 4953
rect 4736 4656 4763 4663
rect 4736 4647 4743 4656
rect 4816 4643 4823 4956
rect 4836 4656 4863 4663
rect 4816 4636 4843 4643
rect 4736 4496 4763 4503
rect 4736 4327 4743 4496
rect 4776 4447 4783 4463
rect 4696 4236 4723 4243
rect 4596 4016 4623 4023
rect 4596 4007 4603 4016
rect 4636 3996 4653 4003
rect 4556 3916 4583 3923
rect 4536 3743 4543 3833
rect 4476 3736 4503 3743
rect 4536 3736 4563 3743
rect 4356 3587 4363 3703
rect 4476 3687 4483 3736
rect 4556 3687 4563 3736
rect 4576 3683 4583 3916
rect 4656 3823 4663 3993
rect 4676 3967 4683 3983
rect 4696 3827 4703 4236
rect 4736 4196 4743 4313
rect 4796 4203 4803 4413
rect 4776 4196 4803 4203
rect 4716 4147 4723 4183
rect 4716 4103 4723 4133
rect 4716 4096 4743 4103
rect 4716 3927 4723 4013
rect 4736 3907 4743 4096
rect 4756 3967 4763 4013
rect 4796 3976 4803 4196
rect 4816 4147 4823 4613
rect 4836 4587 4843 4636
rect 4836 4443 4843 4573
rect 4856 4507 4863 4656
rect 4876 4647 4883 4663
rect 4896 4607 4903 4993
rect 4936 4627 4943 5093
rect 4956 4956 4963 4973
rect 4976 4927 4983 5596
rect 5036 5143 5043 5513
rect 5096 5456 5103 5473
rect 5136 5447 5143 5473
rect 5156 5423 5163 5753
rect 5176 5656 5183 5673
rect 5216 5663 5223 5816
rect 5236 5787 5243 5823
rect 5216 5656 5243 5663
rect 5116 5367 5123 5423
rect 5136 5416 5163 5423
rect 5016 5136 5043 5143
rect 5016 5007 5023 5136
rect 5056 5087 5063 5143
rect 5076 5127 5083 5173
rect 5016 4967 5023 4993
rect 5056 4887 5063 4953
rect 5056 4727 5063 4873
rect 5076 4807 5083 5113
rect 5136 5107 5143 5416
rect 5136 4956 5143 4973
rect 5156 4967 5163 5393
rect 5116 4823 5123 4943
rect 5096 4816 5123 4823
rect 4956 4667 4963 4713
rect 4876 4456 4883 4473
rect 4936 4447 4943 4473
rect 4836 4436 4863 4443
rect 4636 3816 4663 3823
rect 4596 3703 4603 3793
rect 4636 3727 4643 3816
rect 4596 3696 4623 3703
rect 4676 3703 4683 3793
rect 4756 3716 4763 3773
rect 4667 3696 4683 3703
rect 4576 3676 4603 3683
rect 4336 3556 4363 3563
rect 4296 3243 4303 3253
rect 4276 3236 4303 3243
rect 4196 3107 4203 3233
rect 4216 3207 4223 3223
rect 4256 3187 4263 3223
rect 4336 3187 4343 3533
rect 4356 3427 4363 3556
rect 4376 3467 4383 3673
rect 4416 3603 4423 3673
rect 4396 3596 4423 3603
rect 4396 3547 4403 3596
rect 4396 3516 4503 3523
rect 4396 3507 4403 3516
rect 4496 3507 4503 3516
rect 4416 3363 4423 3483
rect 4416 3356 4443 3363
rect 4216 3047 4223 3073
rect 4156 3016 4183 3023
rect 4216 3016 4223 3033
rect 4156 2787 4163 3016
rect 4236 2987 4243 3003
rect 4256 2827 4263 3113
rect 4256 2787 4263 2813
rect 4236 2727 4243 2753
rect 4096 2407 4103 2693
rect 4256 2576 4263 2733
rect 4256 2347 4263 2533
rect 3976 2336 4003 2343
rect 3956 2283 3963 2333
rect 3956 2276 3983 2283
rect 3956 2167 3963 2276
rect 3996 2067 4003 2336
rect 4276 2323 4283 3133
rect 4356 3107 4363 3223
rect 4296 2807 4303 3053
rect 4296 2756 4303 2793
rect 4336 2743 4343 3093
rect 4356 3036 4363 3053
rect 4376 3007 4383 3173
rect 4396 3067 4403 3223
rect 4416 3167 4423 3173
rect 4416 3043 4423 3153
rect 4436 3107 4443 3356
rect 4476 3243 4483 3493
rect 4576 3483 4583 3533
rect 4556 3476 4583 3483
rect 4467 3236 4483 3243
rect 4456 3216 4483 3223
rect 4456 3127 4463 3216
rect 4396 3036 4423 3043
rect 4316 2736 4343 2743
rect 4356 2443 4363 2993
rect 4376 2536 4383 2873
rect 4416 2767 4423 2933
rect 4416 2447 4423 2523
rect 4336 2436 4363 2443
rect 4256 2316 4283 2323
rect 4016 2087 4023 2293
rect 3936 2056 3963 2063
rect 3936 2007 3943 2033
rect 3936 1983 3943 1993
rect 3916 1976 3943 1983
rect 3916 1827 3923 1976
rect 3956 1827 3963 2056
rect 4016 1863 4023 2053
rect 4036 1887 4043 2153
rect 4056 2047 4063 2113
rect 4016 1856 4043 1863
rect 3916 1596 3923 1653
rect 3836 1436 3863 1443
rect 3656 1316 3663 1333
rect 3696 1327 3703 1393
rect 3636 1223 3643 1303
rect 3716 1267 3723 1333
rect 3736 1287 3743 1373
rect 3776 1316 3783 1373
rect 3796 1267 3803 1303
rect 3816 1227 3823 1323
rect 3636 1216 3663 1223
rect 3436 307 3443 323
rect 3316 216 3343 223
rect 3316 176 3323 193
rect 3036 107 3043 123
rect 3156 107 3163 123
rect 3196 116 3203 173
rect 3336 147 3343 216
rect 3376 156 3383 193
rect 3476 -17 3483 833
rect 3496 823 3503 973
rect 3536 927 3543 1133
rect 3636 1116 3643 1193
rect 3656 1107 3663 1216
rect 3496 816 3513 823
rect 3556 807 3563 823
rect 3556 647 3563 673
rect 3596 663 3603 1073
rect 3656 1047 3663 1093
rect 3656 836 3663 913
rect 3676 847 3683 1173
rect 3696 1087 3703 1113
rect 3716 1096 3723 1193
rect 3776 1123 3783 1193
rect 3796 1147 3803 1173
rect 3836 1123 3843 1413
rect 3856 1187 3863 1436
rect 3896 1227 3903 1573
rect 3956 1427 3963 1733
rect 3976 1707 3983 1783
rect 3996 1667 4003 1773
rect 3916 1316 3923 1353
rect 3776 1116 3803 1123
rect 3756 1047 3763 1103
rect 3796 1087 3803 1116
rect 3816 1116 3843 1123
rect 3696 836 3703 973
rect 3796 947 3803 1053
rect 3816 923 3823 1116
rect 3856 1096 3863 1133
rect 3796 916 3823 923
rect 3636 683 3643 823
rect 3576 656 3603 663
rect 3616 676 3643 683
rect 3496 407 3503 433
rect 3576 407 3583 656
rect 3616 647 3623 676
rect 3596 603 3603 633
rect 3636 616 3643 653
rect 3596 596 3623 603
rect 3496 343 3503 393
rect 3536 356 3543 373
rect 3596 363 3603 393
rect 3676 387 3683 633
rect 3696 627 3703 633
rect 3576 356 3603 363
rect 3647 356 3663 363
rect 3696 356 3703 453
rect 3716 383 3723 853
rect 3796 847 3803 916
rect 3756 836 3783 843
rect 3736 647 3743 833
rect 3756 807 3763 836
rect 3796 727 3803 773
rect 3816 667 3823 893
rect 3836 863 3843 1073
rect 3856 887 3863 933
rect 3876 907 3883 1073
rect 3896 867 3903 1113
rect 3916 1027 3923 1093
rect 3936 1083 3943 1283
rect 3976 1127 3983 1613
rect 4016 1607 4023 1833
rect 4036 1563 4043 1856
rect 4056 1596 4063 1873
rect 4076 1687 4083 2093
rect 4176 2083 4183 2253
rect 4256 2107 4263 2316
rect 4316 2303 4323 2433
rect 4296 2296 4323 2303
rect 4156 2076 4183 2083
rect 4096 1816 4103 1933
rect 4116 1847 4123 2033
rect 4136 1907 4143 2073
rect 4156 1787 4163 1913
rect 4176 1887 4183 2076
rect 4016 1556 4043 1563
rect 4016 1487 4023 1556
rect 4076 1367 4083 1633
rect 4096 1327 4103 1693
rect 4136 1576 4143 1593
rect 4116 1527 4123 1563
rect 4176 1387 4183 1833
rect 4196 1783 4203 2053
rect 4216 2043 4223 2073
rect 4216 2036 4243 2043
rect 4276 2027 4283 2043
rect 4296 1987 4303 2296
rect 4336 2163 4343 2436
rect 4356 2287 4363 2393
rect 4376 2227 4383 2313
rect 4316 2156 4343 2163
rect 4296 1967 4303 1973
rect 4316 1927 4323 2156
rect 4416 2076 4423 2393
rect 4436 2327 4443 3033
rect 4456 2743 4463 2833
rect 4456 2736 4483 2743
rect 4456 2507 4463 2736
rect 4516 2667 4523 3453
rect 4556 3287 4563 3476
rect 4596 3387 4603 3676
rect 4616 3467 4623 3513
rect 4556 3187 4563 3223
rect 4576 3207 4583 3273
rect 4656 3207 4663 3553
rect 4676 3547 4683 3593
rect 4576 3036 4583 3193
rect 4676 3187 4683 3533
rect 4696 3516 4703 3533
rect 4736 3516 4743 3593
rect 4716 3223 4723 3273
rect 4756 3236 4763 3653
rect 4776 3607 4783 3703
rect 4816 3447 4823 3853
rect 4836 3747 4843 4436
rect 4916 4183 4923 4293
rect 4856 4167 4863 4183
rect 4896 4176 4923 4183
rect 4856 3887 4863 4153
rect 4936 4107 4943 4393
rect 4916 3976 4923 4013
rect 4896 3956 4903 3973
rect 4836 3427 4843 3453
rect 4796 3227 4803 3243
rect 4716 3216 4743 3223
rect 4716 3067 4723 3093
rect 4716 3036 4723 3053
rect 4536 2727 4543 3013
rect 4596 3003 4603 3023
rect 4576 2996 4603 3003
rect 4556 2687 4563 2743
rect 4576 2627 4583 2996
rect 4616 2843 4623 2993
rect 4596 2836 4623 2843
rect 4596 2787 4603 2836
rect 4496 2536 4523 2543
rect 4456 2487 4463 2493
rect 4476 2447 4483 2523
rect 4496 2407 4503 2536
rect 4436 2296 4443 2313
rect 4476 2263 4483 2293
rect 4456 2256 4483 2263
rect 4456 2143 4463 2256
rect 4516 2147 4523 2453
rect 4616 2387 4623 2813
rect 4696 2747 4703 3033
rect 4736 2947 4743 3023
rect 4776 3016 4783 3033
rect 4796 2967 4803 3193
rect 4816 3007 4823 3273
rect 4636 2576 4643 2593
rect 4796 2443 4803 2953
rect 4816 2687 4823 2743
rect 4816 2536 4823 2673
rect 4836 2467 4843 3413
rect 4776 2436 4803 2443
rect 4556 2276 4563 2313
rect 4536 2207 4543 2263
rect 4576 2223 4583 2263
rect 4556 2216 4583 2223
rect 4436 2136 4463 2143
rect 4436 2067 4443 2136
rect 4336 2056 4363 2063
rect 4216 1867 4223 1893
rect 4276 1796 4283 1833
rect 4196 1776 4223 1783
rect 4296 1723 4303 1783
rect 4336 1767 4343 2056
rect 4336 1747 4343 1753
rect 4296 1716 4323 1723
rect 4316 1683 4323 1716
rect 4336 1707 4343 1713
rect 4356 1683 4363 1833
rect 4376 1816 4383 1833
rect 4416 1823 4423 1913
rect 4456 1847 4463 2093
rect 4516 2076 4523 2093
rect 4556 2087 4563 2216
rect 4416 1816 4443 1823
rect 4316 1676 4343 1683
rect 4356 1676 4383 1683
rect 4016 1287 4023 1323
rect 4096 1303 4103 1313
rect 4016 1083 4023 1133
rect 3936 1076 3963 1083
rect 3996 1076 4023 1083
rect 3836 856 3863 863
rect 3816 636 3823 653
rect 3736 616 3763 623
rect 3736 607 3743 616
rect 3736 407 3743 593
rect 3716 376 3743 383
rect 3496 336 3523 343
rect 3556 207 3563 343
rect 3636 323 3643 353
rect 3636 316 3663 323
rect 3656 136 3663 316
rect 3676 307 3683 323
rect 3736 187 3743 376
rect 3756 156 3783 163
rect 3796 156 3803 393
rect 3816 376 3823 513
rect 3836 407 3843 833
rect 3856 767 3863 856
rect 3856 643 3863 753
rect 3876 707 3883 843
rect 3956 823 3963 1076
rect 3996 856 4003 893
rect 4036 883 4043 1303
rect 4076 1296 4103 1303
rect 4056 1116 4083 1123
rect 4056 1067 4063 1116
rect 4136 887 4143 1353
rect 4176 1287 4183 1303
rect 4176 1143 4183 1273
rect 4216 1247 4223 1303
rect 4216 1207 4223 1233
rect 4176 1136 4203 1143
rect 4036 876 4063 883
rect 3936 816 3963 823
rect 3896 663 3903 713
rect 3887 656 3903 663
rect 3856 636 3883 643
rect 3936 616 3943 653
rect 3856 427 3863 613
rect 3956 547 3963 816
rect 4056 807 4063 876
rect 3996 627 4003 793
rect 4036 656 4043 693
rect 4076 647 4083 773
rect 3836 347 3843 363
rect 3876 347 3883 363
rect 3896 183 3903 413
rect 3916 367 3923 533
rect 4016 527 4023 623
rect 4096 403 4103 873
rect 4156 867 4163 1113
rect 4116 447 4123 853
rect 4176 847 4183 1113
rect 4216 927 4223 1103
rect 4136 807 4143 843
rect 4156 407 4163 823
rect 4216 667 4223 913
rect 4236 907 4243 1673
rect 4296 1596 4303 1653
rect 4336 1607 4343 1676
rect 4316 1487 4323 1583
rect 4276 1287 4283 1473
rect 4356 1407 4363 1653
rect 4356 1316 4363 1393
rect 4376 1187 4383 1676
rect 4396 1643 4403 1803
rect 4436 1787 4443 1816
rect 4496 1796 4503 1833
rect 4456 1707 4463 1793
rect 4396 1636 4423 1643
rect 4416 1596 4423 1636
rect 4487 1616 4493 1623
rect 4456 1596 4463 1613
rect 4476 1563 4483 1583
rect 4476 1556 4503 1563
rect 4436 1267 4443 1323
rect 4476 1316 4483 1473
rect 4496 1347 4503 1556
rect 4516 1307 4523 1783
rect 4536 1747 4543 1803
rect 4556 1787 4563 1833
rect 4556 1727 4563 1773
rect 4536 1387 4543 1613
rect 4556 1587 4563 1693
rect 4576 1607 4583 2193
rect 4596 1807 4603 2233
rect 4636 2167 4643 2313
rect 4616 1707 4623 2013
rect 4656 2007 4663 2043
rect 4676 1847 4683 2353
rect 4696 2296 4703 2393
rect 4716 2267 4723 2283
rect 4696 1823 4703 2093
rect 4716 2027 4723 2173
rect 4776 2107 4783 2436
rect 4796 2043 4803 2393
rect 4856 2367 4863 3813
rect 4876 3716 4883 3733
rect 4916 3703 4923 3893
rect 4896 3696 4923 3703
rect 4876 3227 4883 3673
rect 4896 3587 4903 3696
rect 4936 3367 4943 3483
rect 4956 3287 4963 4653
rect 5056 4647 5063 4663
rect 5016 4476 5023 4613
rect 5076 4483 5083 4593
rect 5096 4527 5103 4816
rect 5116 4667 5123 4693
rect 5136 4547 5143 4913
rect 5176 4847 5183 5333
rect 5216 5327 5223 5613
rect 5236 5567 5243 5656
rect 5316 5636 5323 5653
rect 5236 5487 5243 5553
rect 5236 5407 5243 5473
rect 5256 5436 5263 5513
rect 5236 5387 5243 5393
rect 5276 5163 5283 5413
rect 5256 5156 5283 5163
rect 5196 5127 5203 5143
rect 5196 4963 5203 5093
rect 5236 5087 5243 5143
rect 5296 5023 5303 5193
rect 5276 5016 5303 5023
rect 5196 4956 5223 4963
rect 5216 4867 5223 4956
rect 5196 4696 5203 4713
rect 5076 4476 5103 4483
rect 4996 4427 5003 4463
rect 5036 4456 5063 4463
rect 4976 4007 4983 4163
rect 4976 3383 4983 3493
rect 4996 3487 5003 4133
rect 5016 4016 5023 4433
rect 5056 4427 5063 4456
rect 5056 4167 5063 4213
rect 5027 3976 5043 3983
rect 5016 3736 5023 3753
rect 5076 3687 5083 4476
rect 5136 4407 5143 4453
rect 5156 4227 5163 4513
rect 5176 4476 5183 4493
rect 5196 4443 5203 4633
rect 5216 4527 5223 4733
rect 5236 4443 5243 4833
rect 5276 4747 5283 5016
rect 5296 4956 5303 4993
rect 5316 4727 5323 5593
rect 5336 5523 5343 5623
rect 5356 5607 5363 5643
rect 5336 5516 5363 5523
rect 5356 5207 5363 5516
rect 5376 5123 5383 5613
rect 5336 5107 5343 5123
rect 5356 5116 5383 5123
rect 5336 4956 5343 5053
rect 5256 4563 5263 4713
rect 5276 4696 5283 4713
rect 5296 4567 5303 4683
rect 5316 4607 5323 4653
rect 5336 4647 5343 4693
rect 5356 4647 5363 5116
rect 5376 4727 5383 4773
rect 5376 4667 5383 4693
rect 5396 4607 5403 5773
rect 5456 5636 5463 5693
rect 5516 5663 5523 5823
rect 5556 5767 5563 5823
rect 5596 5787 5603 5823
rect 5636 5687 5643 5823
rect 5516 5656 5543 5663
rect 5516 5627 5523 5656
rect 5416 4707 5423 5573
rect 5436 5436 5443 5473
rect 5456 5367 5463 5423
rect 5496 5416 5503 5433
rect 5436 4927 5443 5143
rect 5456 5067 5463 5113
rect 5436 4907 5443 4913
rect 5456 4787 5463 4973
rect 5256 4556 5283 4563
rect 5176 4436 5203 4443
rect 5216 4436 5243 4443
rect 5136 4196 5143 4213
rect 5176 4183 5183 4436
rect 5196 4407 5203 4413
rect 5196 4207 5203 4393
rect 5156 4176 5183 4183
rect 5116 4127 5123 4163
rect 5116 3987 5123 4093
rect 5176 4003 5183 4153
rect 5196 4047 5203 4193
rect 5216 4147 5223 4436
rect 5276 4227 5283 4556
rect 5296 4527 5303 4533
rect 5296 4247 5303 4513
rect 5316 4183 5323 4593
rect 5236 4107 5243 4183
rect 5276 4087 5283 4183
rect 5296 4176 5323 4183
rect 5296 4067 5303 4176
rect 5176 3996 5203 4003
rect 5136 3967 5143 3983
rect 5036 3516 5043 3553
rect 5056 3467 5063 3503
rect 4976 3376 5003 3383
rect 4896 3256 4903 3273
rect 4976 3227 4983 3353
rect 4996 3243 5003 3376
rect 4996 3236 5023 3243
rect 4916 2987 4923 3003
rect 4896 2736 4923 2743
rect 4916 2727 4923 2736
rect 4816 2107 4823 2273
rect 4836 2247 4843 2263
rect 4776 2036 4803 2043
rect 4716 1867 4723 1873
rect 4656 1816 4703 1823
rect 4616 1596 4623 1613
rect 4556 1327 4563 1553
rect 4596 1547 4603 1583
rect 4676 1347 4683 1816
rect 4716 1783 4723 1853
rect 4736 1827 4743 2033
rect 4816 2027 4823 2093
rect 4696 1776 4723 1783
rect 4436 1227 4443 1253
rect 4256 843 4263 1173
rect 4356 1147 4363 1153
rect 4396 1103 4403 1153
rect 4376 1096 4403 1103
rect 4416 1087 4423 1193
rect 4456 1107 4463 1133
rect 4476 1096 4483 1253
rect 4496 1167 4503 1303
rect 4536 1116 4543 1153
rect 4576 847 4583 1273
rect 4616 1147 4623 1303
rect 4656 1187 4663 1333
rect 4696 1287 4703 1753
rect 4736 1703 4743 1813
rect 4756 1767 4763 2013
rect 4796 1807 4803 1873
rect 4776 1747 4783 1783
rect 4716 1696 4743 1703
rect 4716 1347 4723 1696
rect 4776 1607 4783 1673
rect 4796 1647 4803 1763
rect 4756 1576 4763 1593
rect 4736 1507 4743 1553
rect 4776 1527 4783 1563
rect 4756 1336 4763 1413
rect 4796 1287 4803 1613
rect 4816 1547 4823 1693
rect 4836 1667 4843 2233
rect 4856 2047 4863 2333
rect 4896 2327 4903 2543
rect 4896 2187 4903 2293
rect 4916 2287 4923 2713
rect 4936 2307 4943 3213
rect 4956 2787 4963 3213
rect 5036 3047 5043 3223
rect 5096 3203 5103 3933
rect 5136 3927 5143 3953
rect 5136 3716 5143 3793
rect 5156 3707 5163 3753
rect 5156 3527 5163 3693
rect 5176 3587 5183 3996
rect 5136 3467 5143 3513
rect 5076 3196 5103 3203
rect 4996 3016 5003 3033
rect 4976 2987 4983 3003
rect 4956 2747 4963 2773
rect 4976 2723 4983 2753
rect 4996 2727 5003 2733
rect 4956 2716 4983 2723
rect 4956 2276 4963 2716
rect 5036 2563 5043 2743
rect 5016 2556 5043 2563
rect 5056 2556 5063 2673
rect 4976 2267 4983 2433
rect 5076 2347 5083 3196
rect 5116 3067 5123 3453
rect 5156 3267 5163 3473
rect 5196 3467 5203 3483
rect 5176 3067 5183 3203
rect 5116 3007 5123 3053
rect 5176 3036 5203 3043
rect 5196 3027 5203 3036
rect 5176 2787 5183 2973
rect 5136 2447 5143 2563
rect 4956 2076 4963 2133
rect 4856 1627 4863 1833
rect 4876 1627 4883 2073
rect 4976 1883 4983 2253
rect 5036 2207 5043 2263
rect 5036 2187 5043 2193
rect 4956 1876 4983 1883
rect 4896 1816 4903 1853
rect 4836 1596 4863 1603
rect 4836 1567 4843 1596
rect 4856 1407 4863 1553
rect 4876 1527 4883 1583
rect 4916 1576 4923 1733
rect 4816 1303 4823 1393
rect 4856 1316 4863 1373
rect 4816 1296 4843 1303
rect 4796 1267 4803 1273
rect 4656 1136 4663 1173
rect 4596 1116 4623 1123
rect 4596 887 4603 1116
rect 4636 1087 4643 1103
rect 4656 883 4663 1093
rect 4696 1087 4703 1173
rect 4716 1147 4723 1153
rect 4716 1107 4723 1133
rect 4736 1116 4743 1133
rect 4756 1087 4763 1103
rect 4796 1096 4803 1253
rect 4876 1207 4883 1303
rect 4856 1116 4883 1123
rect 4816 1087 4823 1113
rect 4856 1087 4863 1116
rect 4727 1076 4743 1083
rect 4736 1063 4743 1076
rect 4776 1063 4783 1073
rect 4736 1056 4783 1063
rect 4636 876 4663 883
rect 4256 836 4283 843
rect 4256 827 4263 836
rect 4296 807 4303 823
rect 4336 767 4343 823
rect 4356 656 4363 673
rect 4176 636 4183 653
rect 4216 567 4223 593
rect 4076 396 4103 403
rect 3976 376 4003 383
rect 3996 347 4003 376
rect 4016 267 4023 353
rect 3876 176 3903 183
rect 3636 107 3643 123
rect 3776 -17 3783 156
rect 3876 -17 3883 176
rect 3896 156 3923 163
rect 3916 -17 3923 156
rect 4016 147 4023 253
rect 4056 123 4063 193
rect 4076 167 4083 396
rect 4176 363 4183 393
rect 4196 367 4203 433
rect 4216 396 4323 403
rect 4156 356 4183 363
rect 4216 347 4223 396
rect 4176 287 4183 313
rect 4236 307 4243 363
rect 4296 303 4303 343
rect 4316 327 4323 396
rect 4376 367 4383 653
rect 4396 627 4403 833
rect 4516 747 4523 833
rect 4536 827 4543 843
rect 4616 823 4623 853
rect 4556 807 4563 823
rect 4596 816 4623 823
rect 4436 636 4443 693
rect 4596 636 4603 673
rect 4636 647 4643 876
rect 4656 836 4663 853
rect 4676 747 4683 803
rect 4716 687 4723 823
rect 4736 807 4743 833
rect 4776 807 4783 853
rect 4656 627 4663 653
rect 4776 647 4783 753
rect 4796 667 4803 873
rect 4816 807 4823 823
rect 4856 787 4863 823
rect 4496 467 4503 623
rect 4716 616 4723 633
rect 4796 627 4803 653
rect 4836 627 4843 673
rect 4856 647 4863 693
rect 4876 667 4883 873
rect 4896 867 4903 1273
rect 4916 1116 4923 1133
rect 4896 847 4903 853
rect 4916 787 4923 1073
rect 4936 887 4943 1613
rect 4956 1087 4963 1876
rect 4976 1807 4983 1833
rect 4996 1827 5003 2153
rect 5016 2087 5023 2113
rect 5056 2076 5063 2133
rect 5076 2127 5083 2263
rect 5136 2247 5143 2273
rect 5096 2076 5103 2113
rect 5016 2056 5043 2063
rect 5016 2027 5023 2056
rect 5076 2047 5083 2063
rect 4996 1767 5003 1813
rect 5036 1796 5043 1833
rect 5076 1796 5083 1913
rect 5016 1687 5023 1773
rect 5096 1767 5103 1783
rect 5016 1627 5023 1673
rect 4996 1596 5023 1603
rect 4996 1527 5003 1596
rect 5036 1547 5043 1563
rect 4976 1147 4983 1303
rect 5016 1287 5023 1293
rect 4996 1247 5003 1283
rect 5016 1067 5023 1103
rect 5016 823 5023 953
rect 5036 907 5043 1453
rect 5056 967 5063 1753
rect 5116 1663 5123 2113
rect 5136 1807 5143 2233
rect 5156 2127 5163 2313
rect 5176 2107 5183 2733
rect 5196 2687 5203 3013
rect 5216 2707 5223 3873
rect 5236 3747 5243 4053
rect 5256 3807 5263 4033
rect 5276 3996 5293 4003
rect 5316 3996 5323 4053
rect 5336 4007 5343 4493
rect 5356 4476 5363 4513
rect 5356 4127 5363 4433
rect 5376 4427 5383 4463
rect 5416 4456 5423 4633
rect 5296 3727 5303 3993
rect 5376 3723 5383 4133
rect 5396 3887 5403 4153
rect 5416 4047 5423 4413
rect 5436 4167 5443 4653
rect 5456 4087 5463 4633
rect 5476 4447 5483 5113
rect 5496 5107 5503 5163
rect 5516 5127 5523 5593
rect 5556 4987 5563 5643
rect 5576 5367 5583 5613
rect 5636 5483 5643 5653
rect 5656 5587 5663 5603
rect 5636 5476 5663 5483
rect 5596 5367 5603 5403
rect 5576 4967 5583 5193
rect 5596 5176 5603 5313
rect 5636 5187 5643 5353
rect 5616 4983 5623 5163
rect 5607 4976 5623 4983
rect 5556 4956 5573 4963
rect 5556 4923 5563 4956
rect 5496 4887 5503 4923
rect 5536 4916 5563 4923
rect 5536 4727 5543 4893
rect 5576 4747 5583 4933
rect 5596 4903 5603 4923
rect 5596 4896 5623 4903
rect 5596 4727 5603 4873
rect 5616 4807 5623 4896
rect 5656 4743 5663 5476
rect 5676 5407 5683 5533
rect 5696 5403 5703 5823
rect 5716 5467 5723 5633
rect 5736 5547 5743 5823
rect 5736 5416 5743 5433
rect 5696 5396 5723 5403
rect 5676 5207 5683 5393
rect 5696 5183 5703 5396
rect 5756 5387 5763 5403
rect 5716 5207 5723 5373
rect 5747 5196 5753 5203
rect 5676 5176 5703 5183
rect 5736 5176 5763 5183
rect 5676 4927 5683 5176
rect 5756 5147 5763 5176
rect 5636 4736 5663 4743
rect 5496 4527 5503 4713
rect 5516 4696 5543 4703
rect 5576 4696 5603 4703
rect 5516 4627 5523 4696
rect 5596 4667 5603 4696
rect 5516 4476 5543 4483
rect 5536 4407 5543 4476
rect 5576 4463 5583 4653
rect 5556 4456 5583 4463
rect 5556 4203 5563 4293
rect 5536 4196 5563 4203
rect 5576 4187 5583 4413
rect 5416 4003 5423 4013
rect 5416 3996 5443 4003
rect 5416 3763 5423 3973
rect 5436 3827 5443 3996
rect 5356 3716 5383 3723
rect 5396 3756 5423 3763
rect 5356 3627 5363 3716
rect 5236 3147 5243 3573
rect 5316 3516 5323 3553
rect 5336 3523 5343 3533
rect 5336 3516 5363 3523
rect 5296 3283 5303 3513
rect 5296 3276 5323 3283
rect 5256 3256 5263 3273
rect 5276 3207 5283 3243
rect 5256 2756 5263 3033
rect 5316 2767 5323 3276
rect 5336 3023 5343 3516
rect 5376 3487 5383 3533
rect 5356 3067 5363 3203
rect 5336 3016 5363 3023
rect 5276 2756 5303 2763
rect 5196 2327 5203 2473
rect 5276 2367 5283 2756
rect 5316 2347 5323 2733
rect 5196 2296 5203 2313
rect 5316 2307 5323 2333
rect 5216 2267 5223 2283
rect 5096 1656 5123 1663
rect 5076 1596 5083 1653
rect 5076 1467 5083 1553
rect 5096 1427 5103 1656
rect 5116 1527 5123 1633
rect 5136 1387 5143 1773
rect 5156 1607 5163 2053
rect 5196 2047 5203 2093
rect 5176 1583 5183 1713
rect 5196 1687 5203 1763
rect 5156 1576 5183 1583
rect 5196 1576 5203 1653
rect 5216 1647 5223 2193
rect 5236 2043 5243 2113
rect 5256 2087 5263 2293
rect 5276 2107 5283 2293
rect 5316 2276 5323 2293
rect 5296 2076 5323 2083
rect 5316 2067 5323 2076
rect 5236 2036 5263 2043
rect 5236 1747 5243 2013
rect 5256 1927 5263 2036
rect 5136 1336 5143 1353
rect 5076 1136 5103 1143
rect 5036 827 5043 853
rect 5056 836 5063 953
rect 5076 847 5083 1136
rect 5136 1103 5143 1173
rect 5116 1096 5143 1103
rect 5096 836 5103 853
rect 4996 816 5023 823
rect 5116 807 5123 823
rect 4996 656 5003 673
rect 4916 616 4923 653
rect 4516 387 4523 393
rect 4456 376 4483 383
rect 4416 323 4423 373
rect 4396 316 4423 323
rect 4296 296 4323 303
rect 4096 127 4103 153
rect 4036 116 4063 123
rect 4136 123 4143 193
rect 4176 156 4183 273
rect 4316 176 4323 296
rect 4336 156 4343 193
rect 4416 136 4423 293
rect 4456 267 4463 376
rect 4536 367 4543 453
rect 4576 287 4583 353
rect 4596 347 4603 363
rect 4676 343 4683 353
rect 4616 327 4623 343
rect 4656 336 4683 343
rect 4516 156 4573 163
rect 4136 116 4163 123
rect 4456 123 4463 133
rect 4516 127 4523 156
rect 4596 136 4603 213
rect 4616 147 4623 153
rect 4436 116 4463 123
rect 4536 107 4543 123
rect 4636 107 4643 233
rect 4696 136 4703 213
rect 4756 156 4763 173
rect 4736 123 4743 143
rect 4796 123 4803 493
rect 4816 387 4823 593
rect 4816 363 4823 373
rect 4816 356 4843 363
rect 4876 356 4883 613
rect 4956 367 4963 653
rect 5016 387 5023 623
rect 5096 487 5103 653
rect 5116 636 5123 773
rect 5136 667 5143 893
rect 5156 687 5163 1513
rect 5156 636 5163 653
rect 5136 427 5143 633
rect 4816 327 4823 356
rect 4996 356 5023 363
rect 4856 247 4863 343
rect 4976 327 4983 343
rect 4876 123 4883 153
rect 4956 136 4963 213
rect 4996 207 5003 356
rect 5076 187 5083 393
rect 5156 387 5163 433
rect 5176 387 5183 1433
rect 5196 403 5203 1533
rect 5216 1527 5223 1563
rect 5236 1447 5243 1713
rect 5256 1667 5263 1853
rect 5296 1807 5303 1893
rect 5336 1867 5343 2263
rect 5356 2207 5363 2693
rect 5376 2107 5383 2313
rect 5396 2267 5403 3756
rect 5436 3696 5443 3713
rect 5436 3447 5443 3523
rect 5436 3403 5443 3433
rect 5416 3396 5443 3403
rect 5416 2427 5423 3396
rect 5436 2847 5443 3373
rect 5456 2927 5463 3613
rect 5476 3387 5483 4113
rect 5496 3987 5503 4073
rect 5516 4067 5523 4183
rect 5516 4007 5523 4033
rect 5496 3487 5503 3733
rect 5536 3527 5543 4153
rect 5556 3667 5563 3703
rect 5576 3527 5583 4173
rect 5596 4083 5603 4513
rect 5616 4307 5623 4733
rect 5596 4076 5623 4083
rect 5616 3787 5623 4076
rect 5516 3287 5523 3493
rect 5596 3483 5603 3513
rect 5576 3476 5603 3483
rect 5576 3447 5583 3476
rect 5556 3243 5563 3273
rect 5536 3236 5563 3243
rect 5516 3047 5523 3223
rect 5536 3043 5543 3053
rect 5536 3036 5563 3043
rect 5496 2927 5503 3023
rect 5436 2687 5443 2743
rect 5456 2547 5463 2913
rect 5496 2723 5503 2833
rect 5476 2716 5503 2723
rect 5416 2296 5423 2373
rect 5356 2043 5363 2073
rect 5396 2056 5403 2233
rect 5436 2127 5443 2283
rect 5356 2036 5383 2043
rect 5356 1847 5363 1853
rect 5316 1767 5323 1783
rect 5296 1743 5303 1763
rect 5296 1736 5313 1743
rect 5336 1687 5343 1833
rect 5376 1823 5383 2036
rect 5416 2027 5423 2043
rect 5356 1816 5383 1823
rect 5356 1767 5363 1816
rect 5396 1796 5403 1853
rect 5436 1847 5443 2093
rect 5376 1727 5383 1773
rect 5256 1547 5263 1633
rect 5276 1627 5283 1673
rect 5296 1596 5303 1653
rect 5376 1596 5383 1633
rect 5216 1287 5223 1373
rect 5236 1336 5243 1413
rect 5256 1367 5263 1513
rect 5276 1363 5283 1593
rect 5276 1356 5303 1363
rect 5296 1267 5303 1356
rect 5316 1347 5323 1513
rect 5336 1467 5343 1553
rect 5396 1547 5403 1713
rect 5416 1507 5423 1753
rect 5436 1747 5443 1803
rect 5456 1727 5463 2253
rect 5476 2047 5483 2716
rect 5536 2707 5543 2733
rect 5496 2096 5503 2373
rect 5556 2327 5563 3036
rect 5576 2523 5583 2913
rect 5596 2547 5603 3453
rect 5616 3267 5623 3733
rect 5636 3547 5643 4736
rect 5696 4727 5703 5133
rect 5716 4907 5723 5133
rect 5756 5107 5763 5113
rect 5756 4936 5763 4973
rect 5776 4907 5783 4923
rect 5656 4456 5663 4713
rect 5676 4696 5683 4713
rect 5696 4667 5703 4683
rect 5716 4627 5723 4703
rect 5756 4683 5763 4713
rect 5736 4676 5763 4683
rect 5776 4667 5783 4793
rect 5736 4483 5743 4653
rect 5716 4476 5743 4483
rect 5696 4443 5703 4463
rect 5696 4436 5723 4443
rect 5676 4227 5683 4433
rect 5656 3947 5663 4153
rect 5676 4003 5683 4193
rect 5696 4047 5703 4183
rect 5716 4147 5723 4436
rect 5736 4427 5743 4476
rect 5676 3996 5703 4003
rect 5676 3927 5683 3996
rect 5716 3967 5723 3983
rect 5676 3516 5683 3653
rect 5696 3496 5703 3773
rect 5716 3767 5723 3913
rect 5736 3767 5743 3953
rect 5716 3736 5723 3753
rect 5756 3747 5763 3933
rect 5716 3467 5723 3693
rect 5656 3263 5663 3433
rect 5636 3256 5663 3263
rect 5636 3227 5643 3256
rect 5676 3063 5683 3243
rect 5676 3056 5703 3063
rect 5616 3036 5643 3043
rect 5616 3027 5623 3036
rect 5696 2763 5703 3056
rect 5736 2927 5743 3493
rect 5676 2756 5703 2763
rect 5616 2727 5623 2743
rect 5656 2707 5663 2743
rect 5616 2543 5623 2673
rect 5616 2536 5643 2543
rect 5576 2516 5603 2523
rect 5516 2247 5523 2293
rect 5536 2167 5543 2243
rect 5536 2147 5543 2153
rect 5496 2056 5513 2063
rect 5436 1567 5443 1693
rect 5476 1667 5483 2013
rect 5496 1887 5503 2056
rect 5496 1807 5503 1873
rect 5476 1576 5483 1593
rect 5316 1147 5323 1333
rect 5396 1316 5403 1333
rect 5376 1167 5383 1303
rect 5416 1267 5423 1303
rect 5236 1096 5243 1133
rect 5276 1083 5283 1113
rect 5216 836 5223 1083
rect 5256 1076 5283 1083
rect 5216 527 5223 673
rect 5196 396 5223 403
rect 5136 327 5143 353
rect 5096 176 5103 193
rect 5036 147 5043 173
rect 5076 156 5083 173
rect 4736 116 4823 123
rect 4856 116 4883 123
rect 5196 123 5203 233
rect 5216 207 5223 396
rect 5236 367 5243 873
rect 5256 747 5263 793
rect 5276 687 5283 793
rect 5296 787 5303 1133
rect 5336 1123 5343 1153
rect 5316 1116 5343 1123
rect 5316 887 5323 1116
rect 5416 1116 5423 1133
rect 5336 1096 5363 1103
rect 5316 827 5323 833
rect 5316 636 5323 813
rect 5336 807 5343 1096
rect 5416 827 5423 893
rect 5436 747 5443 1473
rect 5296 607 5303 623
rect 5336 607 5343 713
rect 5356 467 5363 693
rect 5376 636 5383 693
rect 5436 616 5443 693
rect 5456 667 5463 1533
rect 5496 1347 5503 1533
rect 5516 1487 5523 2033
rect 5576 1796 5583 2273
rect 5596 2063 5603 2516
rect 5636 2276 5643 2333
rect 5676 2243 5683 2733
rect 5736 2556 5763 2563
rect 5716 2307 5723 2533
rect 5716 2247 5723 2263
rect 5656 2236 5683 2243
rect 5636 2096 5643 2233
rect 5596 2056 5623 2063
rect 5536 1627 5543 1773
rect 5536 1387 5543 1593
rect 5556 1567 5563 1783
rect 5596 1767 5603 1783
rect 5576 1647 5583 1733
rect 5576 1587 5583 1633
rect 5636 1627 5643 2053
rect 5656 2023 5663 2236
rect 5736 2207 5743 2273
rect 5676 2107 5683 2193
rect 5736 2163 5743 2173
rect 5756 2163 5763 2556
rect 5736 2156 5763 2163
rect 5736 2107 5743 2156
rect 5676 2076 5703 2083
rect 5676 2047 5683 2076
rect 5756 2056 5763 2133
rect 5656 2016 5683 2023
rect 5556 1323 5563 1353
rect 5536 1316 5563 1323
rect 5476 1187 5483 1303
rect 5476 1116 5483 1133
rect 5516 1127 5523 1303
rect 5536 927 5543 1133
rect 5576 1087 5583 1393
rect 5596 1207 5603 1333
rect 5496 847 5503 913
rect 5536 836 5543 873
rect 5576 847 5583 1073
rect 5596 827 5603 1173
rect 5616 1127 5623 1533
rect 5636 1347 5643 1563
rect 5656 1407 5663 1593
rect 5676 1547 5683 2016
rect 5696 2003 5703 2033
rect 5716 2027 5723 2053
rect 5776 2047 5783 4133
rect 5696 1996 5723 2003
rect 5696 1796 5703 1973
rect 5716 1643 5723 1996
rect 5696 1636 5723 1643
rect 5656 1316 5663 1373
rect 5696 1367 5703 1636
rect 5636 1287 5643 1303
rect 5636 1096 5643 1193
rect 5676 1187 5683 1303
rect 5676 1127 5683 1153
rect 5696 1107 5703 1323
rect 5716 1147 5723 1613
rect 5616 907 5623 1083
rect 5696 887 5703 1073
rect 5476 627 5483 733
rect 5496 547 5503 773
rect 5236 167 5243 353
rect 5256 343 5263 453
rect 5296 356 5303 393
rect 5256 336 5283 343
rect 5316 227 5323 343
rect 5356 247 5363 413
rect 5376 347 5383 393
rect 5336 163 5343 193
rect 5336 156 5363 163
rect 5396 156 5403 513
rect 5516 507 5523 823
rect 5596 707 5603 813
rect 5556 636 5563 673
rect 5596 647 5603 693
rect 5536 616 5543 633
rect 5416 327 5423 473
rect 5296 143 5303 153
rect 5356 147 5363 156
rect 5296 136 5323 143
rect 5376 127 5383 143
rect 5436 127 5443 373
rect 5516 356 5523 393
rect 5556 343 5563 393
rect 5596 356 5603 473
rect 5616 447 5623 853
rect 5656 836 5663 853
rect 5636 667 5643 823
rect 5616 387 5623 433
rect 5636 407 5643 653
rect 5656 636 5663 733
rect 5676 656 5683 713
rect 5716 603 5723 1093
rect 5736 607 5743 2033
rect 5756 1596 5763 1633
rect 5796 1607 5803 5693
rect 5816 3947 5823 5673
rect 5816 2147 5823 3813
rect 5776 1527 5783 1583
rect 5756 1167 5763 1353
rect 5776 1136 5783 1493
rect 5696 596 5723 603
rect 5456 187 5463 343
rect 5556 336 5583 343
rect 5467 176 5483 183
rect 5656 147 5663 593
rect 5676 187 5683 533
rect 5696 136 5703 596
rect 5756 407 5763 873
rect 5716 376 5723 393
rect 5776 383 5783 1093
rect 5756 376 5783 383
rect 5796 367 5803 1573
rect 5196 116 5223 123
rect 5736 123 5743 173
rect 5716 116 5743 123
rect 3476 -24 3503 -17
rect 3756 -24 3783 -17
rect 3856 -24 3883 -17
rect 3896 -24 3923 -17
<< m3contact >>
rect 5073 5773 5087 5787
rect 4833 5673 4847 5687
rect 4973 5673 4987 5687
rect 453 5653 467 5667
rect 513 5653 527 5667
rect 113 5633 127 5647
rect 213 5633 227 5647
rect 133 5613 147 5627
rect 193 5613 207 5627
rect 93 5473 107 5487
rect 73 5453 87 5467
rect 133 5453 147 5467
rect 93 5433 107 5447
rect 393 5633 407 5647
rect 373 5613 387 5627
rect 413 5593 427 5607
rect 253 5533 267 5547
rect 393 5473 407 5487
rect 113 5413 127 5427
rect 193 5413 207 5427
rect 273 5433 287 5447
rect 93 5393 107 5407
rect 53 5373 67 5387
rect 73 5373 87 5387
rect 53 5313 67 5327
rect 33 5013 47 5027
rect 33 4773 47 4787
rect 33 4673 47 4687
rect 93 5313 107 5327
rect 173 5233 187 5247
rect 153 5213 167 5227
rect 153 5173 167 5187
rect 93 5153 107 5167
rect 113 5153 127 5167
rect 73 4973 87 4987
rect 133 5113 147 5127
rect 113 4873 127 4887
rect 133 4833 147 4847
rect 113 4773 127 4787
rect 93 4753 107 4767
rect 113 4693 127 4707
rect 233 5233 247 5247
rect 233 5213 247 5227
rect 193 5173 207 5187
rect 193 5153 207 5167
rect 433 5413 447 5427
rect 353 5393 367 5407
rect 273 5173 287 5187
rect 313 5173 327 5187
rect 213 5113 227 5127
rect 353 5153 367 5167
rect 413 5393 427 5407
rect 533 5633 547 5647
rect 493 5593 507 5607
rect 533 5593 547 5607
rect 693 5633 707 5647
rect 733 5633 747 5647
rect 653 5553 667 5567
rect 653 5533 667 5547
rect 533 5473 547 5487
rect 573 5473 587 5487
rect 413 5353 427 5367
rect 453 5353 467 5367
rect 393 5333 407 5347
rect 373 5013 387 5027
rect 373 4973 387 4987
rect 213 4953 227 4967
rect 193 4933 207 4947
rect 233 4933 247 4947
rect 293 4933 307 4947
rect 333 4933 347 4947
rect 493 5413 507 5427
rect 573 5453 587 5467
rect 613 5433 627 5447
rect 593 5413 607 5427
rect 513 5393 527 5407
rect 553 5393 567 5407
rect 493 5353 507 5367
rect 473 5333 487 5347
rect 533 5193 547 5207
rect 453 5173 467 5187
rect 493 5173 507 5187
rect 433 5153 447 5167
rect 473 5153 487 5167
rect 413 5133 427 5147
rect 413 4973 427 4987
rect 393 4953 407 4967
rect 213 4913 227 4927
rect 253 4913 267 4927
rect 313 4913 327 4927
rect 353 4913 367 4927
rect 393 4913 407 4927
rect 213 4893 227 4907
rect 293 4893 307 4907
rect 193 4833 207 4847
rect 173 4773 187 4787
rect 153 4753 167 4767
rect 153 4713 167 4727
rect 53 4493 67 4507
rect 113 4633 127 4647
rect 133 4573 147 4587
rect 93 4493 107 4507
rect 153 4493 167 4507
rect 33 4173 47 4187
rect 73 4453 87 4467
rect 113 4453 127 4467
rect 73 4413 87 4427
rect 193 4713 207 4727
rect 293 4873 307 4887
rect 233 4673 247 4687
rect 193 4633 207 4647
rect 233 4633 247 4647
rect 273 4673 287 4687
rect 273 4653 287 4667
rect 253 4613 267 4627
rect 233 4553 247 4567
rect 173 4433 187 4447
rect 53 4113 67 4127
rect 53 4093 67 4107
rect 133 4193 147 4207
rect 113 4173 127 4187
rect 133 4153 147 4167
rect 113 4113 127 4127
rect 93 4093 107 4107
rect 73 4013 87 4027
rect 93 4013 107 4027
rect 93 3973 107 3987
rect 53 3773 67 3787
rect 13 3133 27 3147
rect 13 3013 27 3027
rect 33 1573 47 1587
rect 13 1553 27 1567
rect 13 1493 27 1507
rect 33 1133 47 1147
rect 173 4173 187 4187
rect 173 4153 187 4167
rect 153 4073 167 4087
rect 153 4033 167 4047
rect 253 4493 267 4507
rect 313 4773 327 4787
rect 373 4713 387 4727
rect 413 4753 427 4767
rect 393 4693 407 4707
rect 373 4673 387 4687
rect 313 4633 327 4647
rect 353 4633 367 4647
rect 353 4613 367 4627
rect 413 4553 427 4567
rect 353 4493 367 4507
rect 293 4473 307 4487
rect 393 4473 407 4487
rect 273 4453 287 4467
rect 213 4433 227 4447
rect 253 4433 267 4447
rect 213 4193 227 4207
rect 273 4193 287 4207
rect 253 4173 267 4187
rect 233 4153 247 4167
rect 213 4133 227 4147
rect 253 4133 267 4147
rect 233 4113 247 4127
rect 193 4033 207 4047
rect 173 4013 187 4027
rect 153 3993 167 4007
rect 213 3993 227 4007
rect 133 3953 147 3967
rect 113 3773 127 3787
rect 113 3753 127 3767
rect 73 3733 87 3747
rect 73 3693 87 3707
rect 133 3693 147 3707
rect 93 3593 107 3607
rect 93 3573 107 3587
rect 133 3553 147 3567
rect 133 3513 147 3527
rect 73 3493 87 3507
rect 113 3493 127 3507
rect 133 3453 147 3467
rect 93 3433 107 3447
rect 113 3433 127 3447
rect 73 3253 87 3267
rect 93 3233 107 3247
rect 93 3193 107 3207
rect 133 3213 147 3227
rect 73 3173 87 3187
rect 113 3173 127 3187
rect 193 3973 207 3987
rect 293 4073 307 4087
rect 293 4033 307 4047
rect 253 3973 267 3987
rect 173 3953 187 3967
rect 333 4453 347 4467
rect 373 4453 387 4467
rect 413 4453 427 4467
rect 333 4433 347 4447
rect 393 4433 407 4447
rect 333 4413 347 4427
rect 373 4253 387 4267
rect 333 4173 347 4187
rect 353 4053 367 4067
rect 333 3973 347 3987
rect 193 3733 207 3747
rect 233 3733 247 3747
rect 313 3733 327 3747
rect 293 3713 307 3727
rect 213 3693 227 3707
rect 253 3693 267 3707
rect 213 3593 227 3607
rect 273 3573 287 3587
rect 293 3573 307 3587
rect 213 3533 227 3547
rect 253 3513 267 3527
rect 293 3513 307 3527
rect 193 3493 207 3507
rect 233 3493 247 3507
rect 273 3493 287 3507
rect 173 3453 187 3467
rect 253 3273 267 3287
rect 173 3233 187 3247
rect 213 3233 227 3247
rect 173 3213 187 3227
rect 113 2993 127 3007
rect 73 2973 87 2987
rect 113 2973 127 2987
rect 73 2793 87 2807
rect 113 2773 127 2787
rect 93 2753 107 2767
rect 93 2733 107 2747
rect 113 2733 127 2747
rect 113 2513 127 2527
rect 73 2293 87 2307
rect 93 2273 107 2287
rect 73 2253 87 2267
rect 73 2113 87 2127
rect 113 2153 127 2167
rect 153 3033 167 3047
rect 233 3213 247 3227
rect 273 3253 287 3267
rect 273 3213 287 3227
rect 253 3193 267 3207
rect 253 3033 267 3047
rect 333 3693 347 3707
rect 513 5133 527 5147
rect 493 5093 507 5107
rect 573 5153 587 5167
rect 713 5573 727 5587
rect 693 5473 707 5487
rect 673 5413 687 5427
rect 833 5653 847 5667
rect 1333 5653 1347 5667
rect 773 5613 787 5627
rect 893 5633 907 5647
rect 933 5633 947 5647
rect 1213 5633 1227 5647
rect 913 5593 927 5607
rect 893 5573 907 5587
rect 793 5553 807 5567
rect 813 5553 827 5567
rect 773 5453 787 5467
rect 993 5593 1007 5607
rect 1073 5593 1087 5607
rect 1253 5613 1267 5627
rect 1053 5533 1067 5547
rect 833 5433 847 5447
rect 953 5433 967 5447
rect 733 5413 747 5427
rect 813 5413 827 5427
rect 853 5413 867 5427
rect 913 5413 927 5427
rect 933 5413 947 5427
rect 673 5393 687 5407
rect 713 5353 727 5367
rect 613 5213 627 5227
rect 613 5173 627 5187
rect 793 5173 807 5187
rect 753 5153 767 5167
rect 1273 5593 1287 5607
rect 1093 5573 1107 5587
rect 1113 5573 1127 5587
rect 1133 5453 1147 5467
rect 1173 5453 1187 5467
rect 973 5413 987 5427
rect 1073 5413 1087 5427
rect 1153 5413 1167 5427
rect 993 5193 1007 5207
rect 1013 5173 1027 5187
rect 1053 5173 1067 5187
rect 873 5153 887 5167
rect 893 5153 907 5167
rect 533 5113 547 5127
rect 593 5113 607 5127
rect 733 5133 747 5147
rect 813 5133 827 5147
rect 853 5133 867 5147
rect 773 5113 787 5127
rect 853 5113 867 5127
rect 733 5093 747 5107
rect 753 5093 767 5107
rect 573 4953 587 4967
rect 633 4953 647 4967
rect 693 4953 707 4967
rect 553 4933 567 4947
rect 493 4873 507 4887
rect 553 4833 567 4847
rect 453 4753 467 4767
rect 513 4693 527 4707
rect 493 4673 507 4687
rect 453 4653 467 4667
rect 453 4633 467 4647
rect 533 4653 547 4667
rect 513 4593 527 4607
rect 493 4573 507 4587
rect 493 4533 507 4547
rect 453 4433 467 4447
rect 433 4253 447 4267
rect 413 4113 427 4127
rect 453 4193 467 4207
rect 653 4933 667 4947
rect 673 4913 687 4927
rect 593 4893 607 4907
rect 633 4893 647 4907
rect 573 4533 587 4547
rect 573 4513 587 4527
rect 613 4693 627 4707
rect 653 4673 667 4687
rect 633 4533 647 4547
rect 653 4533 667 4547
rect 593 4473 607 4487
rect 553 4453 567 4467
rect 693 4553 707 4567
rect 713 4513 727 4527
rect 673 4493 687 4507
rect 673 4473 687 4487
rect 713 4473 727 4487
rect 693 4453 707 4467
rect 533 4433 547 4447
rect 433 4093 447 4107
rect 453 4093 467 4107
rect 413 4053 427 4067
rect 473 3973 487 3987
rect 413 3713 427 3727
rect 493 3713 507 3727
rect 373 3553 387 3567
rect 373 3533 387 3547
rect 433 3693 447 3707
rect 453 3693 467 3707
rect 413 3573 427 3587
rect 393 3493 407 3507
rect 493 3553 507 3567
rect 473 3513 487 3527
rect 453 3493 467 3507
rect 773 4953 787 4967
rect 813 4953 827 4967
rect 793 4933 807 4947
rect 773 4913 787 4927
rect 793 4673 807 4687
rect 913 5133 927 5147
rect 893 5113 907 5127
rect 893 4953 907 4967
rect 1033 5093 1047 5107
rect 953 4973 967 4987
rect 993 4973 1007 4987
rect 1073 5153 1087 5167
rect 1293 5433 1307 5447
rect 1253 5413 1267 5427
rect 1173 5393 1187 5407
rect 1233 5393 1247 5407
rect 1153 5373 1167 5387
rect 1153 5153 1167 5167
rect 1133 5113 1147 5127
rect 1133 5093 1147 5107
rect 1113 5073 1127 5087
rect 933 4933 947 4947
rect 993 4933 1007 4947
rect 1113 4953 1127 4967
rect 1053 4933 1067 4947
rect 1013 4713 1027 4727
rect 873 4653 887 4667
rect 833 4593 847 4607
rect 893 4593 907 4607
rect 1013 4673 1027 4687
rect 1093 4873 1107 4887
rect 1053 4633 1067 4647
rect 993 4553 1007 4567
rect 853 4533 867 4547
rect 933 4533 947 4547
rect 773 4493 787 4507
rect 813 4493 827 4507
rect 793 4453 807 4467
rect 893 4513 907 4527
rect 893 4493 907 4507
rect 933 4473 947 4487
rect 1013 4473 1027 4487
rect 913 4453 927 4467
rect 993 4453 1007 4467
rect 893 4293 907 4307
rect 593 4193 607 4207
rect 573 4153 587 4167
rect 573 4133 587 4147
rect 553 4113 567 4127
rect 733 4193 747 4207
rect 753 4193 767 4207
rect 813 4193 827 4207
rect 853 4193 867 4207
rect 653 4113 667 4127
rect 633 4093 647 4107
rect 593 4053 607 4067
rect 553 4033 567 4047
rect 613 4033 627 4047
rect 593 3993 607 4007
rect 733 4093 747 4107
rect 833 4173 847 4187
rect 813 4153 827 4167
rect 713 3993 727 4007
rect 873 4033 887 4047
rect 853 3993 867 4007
rect 553 3973 567 3987
rect 733 3973 747 3987
rect 833 3973 847 3987
rect 713 3953 727 3967
rect 653 3733 667 3747
rect 593 3713 607 3727
rect 533 3693 547 3707
rect 553 3693 567 3707
rect 613 3673 627 3687
rect 573 3653 587 3667
rect 613 3533 627 3547
rect 593 3513 607 3527
rect 553 3473 567 3487
rect 353 3293 367 3307
rect 413 3293 427 3307
rect 313 3273 327 3287
rect 313 3253 327 3267
rect 313 3233 327 3247
rect 393 3273 407 3287
rect 413 3233 427 3247
rect 393 3213 407 3227
rect 453 3213 467 3227
rect 393 3073 407 3087
rect 353 3053 367 3067
rect 293 3033 307 3047
rect 313 3013 327 3027
rect 473 3033 487 3047
rect 213 2993 227 3007
rect 253 2993 267 3007
rect 413 2993 427 3007
rect 213 2973 227 2987
rect 373 2973 387 2987
rect 253 2793 267 2807
rect 153 2733 167 2747
rect 213 2733 227 2747
rect 193 2713 207 2727
rect 173 2653 187 2667
rect 153 2593 167 2607
rect 173 2533 187 2547
rect 173 2513 187 2527
rect 153 2433 167 2447
rect 153 2253 167 2267
rect 113 1993 127 2007
rect 113 1813 127 1827
rect 93 1793 107 1807
rect 133 1773 147 1787
rect 113 1753 127 1767
rect 133 1693 147 1707
rect 73 1633 87 1647
rect 113 1573 127 1587
rect 93 1553 107 1567
rect 133 1553 147 1567
rect 113 1533 127 1547
rect 73 1513 87 1527
rect 113 1413 127 1427
rect 93 1313 107 1327
rect 113 1233 127 1247
rect 133 1213 147 1227
rect 93 1173 107 1187
rect 233 2573 247 2587
rect 473 2893 487 2907
rect 553 3433 567 3447
rect 593 3433 607 3447
rect 553 3253 567 3267
rect 513 3233 527 3247
rect 573 3113 587 3127
rect 573 3053 587 3067
rect 533 3033 547 3047
rect 513 3013 527 3027
rect 553 3013 567 3027
rect 733 3733 747 3747
rect 813 3713 827 3727
rect 853 3713 867 3727
rect 913 4193 927 4207
rect 913 4153 927 4167
rect 933 4153 947 4167
rect 953 4033 967 4047
rect 973 4013 987 4027
rect 913 3993 927 4007
rect 713 3693 727 3707
rect 733 3693 747 3707
rect 713 3633 727 3647
rect 673 3573 687 3587
rect 653 3293 667 3307
rect 673 3293 687 3307
rect 693 3253 707 3267
rect 713 3213 727 3227
rect 633 3173 647 3187
rect 633 3053 647 3067
rect 673 3053 687 3067
rect 613 3033 627 3047
rect 593 2933 607 2947
rect 373 2773 387 2787
rect 333 2753 347 2767
rect 273 2653 287 2667
rect 353 2653 367 2667
rect 493 2813 507 2827
rect 413 2753 427 2767
rect 453 2753 467 2767
rect 493 2733 507 2747
rect 393 2713 407 2727
rect 473 2713 487 2727
rect 433 2693 447 2707
rect 373 2593 387 2607
rect 293 2533 307 2547
rect 333 2533 347 2547
rect 473 2573 487 2587
rect 393 2553 407 2567
rect 373 2533 387 2547
rect 433 2533 447 2547
rect 273 2513 287 2527
rect 353 2513 367 2527
rect 253 2433 267 2447
rect 233 2293 247 2307
rect 213 2273 227 2287
rect 193 2093 207 2107
rect 193 2033 207 2047
rect 253 2253 267 2267
rect 293 2313 307 2327
rect 353 2313 367 2327
rect 313 2293 327 2307
rect 333 2273 347 2287
rect 293 2253 307 2267
rect 313 2253 327 2267
rect 273 2093 287 2107
rect 293 2093 307 2107
rect 253 2053 267 2067
rect 233 2033 247 2047
rect 293 2053 307 2067
rect 213 1853 227 1867
rect 193 1833 207 1847
rect 293 2013 307 2027
rect 273 1953 287 1967
rect 213 1813 227 1827
rect 233 1813 247 1827
rect 193 1793 207 1807
rect 233 1793 247 1807
rect 213 1753 227 1767
rect 213 1733 227 1747
rect 193 1673 207 1687
rect 253 1713 267 1727
rect 413 2513 427 2527
rect 413 2273 427 2287
rect 453 2273 467 2287
rect 373 2233 387 2247
rect 333 2193 347 2207
rect 433 2253 447 2267
rect 413 2173 427 2187
rect 373 2093 387 2107
rect 413 2073 427 2087
rect 393 2053 407 2067
rect 353 2013 367 2027
rect 413 2013 427 2027
rect 333 1953 347 1967
rect 373 1933 387 1947
rect 333 1833 347 1847
rect 393 1873 407 1887
rect 373 1813 387 1827
rect 413 1813 427 1827
rect 293 1673 307 1687
rect 313 1613 327 1627
rect 273 1593 287 1607
rect 253 1573 267 1587
rect 273 1573 287 1587
rect 213 1553 227 1567
rect 193 1533 207 1547
rect 233 1533 247 1547
rect 293 1473 307 1487
rect 193 1333 207 1347
rect 193 1313 207 1327
rect 233 1313 247 1327
rect 273 1313 287 1327
rect 253 1293 267 1307
rect 173 1253 187 1267
rect 233 1253 247 1267
rect 213 1213 227 1227
rect 213 1153 227 1167
rect 73 1093 87 1107
rect 73 1073 87 1087
rect 173 1133 187 1147
rect 153 1093 167 1107
rect 193 1093 207 1107
rect 133 873 147 887
rect 173 873 187 887
rect 93 833 107 847
rect 133 833 147 847
rect 113 793 127 807
rect 133 713 147 727
rect 153 653 167 667
rect 113 633 127 647
rect 53 613 67 627
rect 93 613 107 627
rect 33 593 47 607
rect 73 593 87 607
rect 73 573 87 587
rect 153 573 167 587
rect 153 533 167 547
rect 93 353 107 367
rect 113 333 127 347
rect 93 153 107 167
rect 153 173 167 187
rect 113 133 127 147
rect 133 133 147 147
rect 273 1233 287 1247
rect 313 1453 327 1467
rect 313 1413 327 1427
rect 313 1253 327 1267
rect 293 1153 307 1167
rect 353 1773 367 1787
rect 373 1773 387 1787
rect 413 1753 427 1767
rect 413 1733 427 1747
rect 353 1713 367 1727
rect 373 1613 387 1627
rect 353 1573 367 1587
rect 373 1573 387 1587
rect 353 1533 367 1547
rect 393 1553 407 1567
rect 373 1513 387 1527
rect 393 1473 407 1487
rect 353 1453 367 1467
rect 393 1313 407 1327
rect 373 1273 387 1287
rect 373 1253 387 1267
rect 353 1113 367 1127
rect 273 1093 287 1107
rect 233 853 247 867
rect 193 833 207 847
rect 253 813 267 827
rect 393 1113 407 1127
rect 373 1093 387 1107
rect 313 1073 327 1087
rect 473 2233 487 2247
rect 493 2233 507 2247
rect 833 3693 847 3707
rect 893 3693 907 3707
rect 773 3673 787 3687
rect 893 3573 907 3587
rect 973 3953 987 3967
rect 1033 4453 1047 4467
rect 1073 4433 1087 4447
rect 1153 5073 1167 5087
rect 1173 4953 1187 4967
rect 1253 5373 1267 5387
rect 1293 5173 1307 5187
rect 1273 5093 1287 5107
rect 1493 5653 1507 5667
rect 1513 5633 1527 5647
rect 1373 5613 1387 5627
rect 1393 5613 1407 5627
rect 1353 5573 1367 5587
rect 1633 5653 1647 5667
rect 1553 5613 1567 5627
rect 1413 5593 1427 5607
rect 1533 5593 1547 5607
rect 1393 5533 1407 5547
rect 1373 5493 1387 5507
rect 1353 5433 1367 5447
rect 1673 5633 1687 5647
rect 1753 5633 1767 5647
rect 1613 5473 1627 5487
rect 1633 5473 1647 5487
rect 1413 5433 1427 5447
rect 1553 5433 1567 5447
rect 1593 5433 1607 5447
rect 1533 5413 1547 5427
rect 1533 5373 1547 5387
rect 1353 5153 1367 5167
rect 1413 5153 1427 5167
rect 1453 5153 1467 5167
rect 1333 5133 1347 5147
rect 1313 5113 1327 5127
rect 1353 5113 1367 5127
rect 1233 4973 1247 4987
rect 1293 4973 1307 4987
rect 1333 4973 1347 4987
rect 1213 4933 1227 4947
rect 1153 4673 1167 4687
rect 1133 4633 1147 4647
rect 1313 4933 1327 4947
rect 1293 4773 1307 4787
rect 1433 5133 1447 5147
rect 1413 5013 1427 5027
rect 1393 4933 1407 4947
rect 1433 4933 1447 4947
rect 1353 4733 1367 4747
rect 1453 4913 1467 4927
rect 1413 4893 1427 4907
rect 1513 5153 1527 5167
rect 1493 4913 1507 4927
rect 1473 4873 1487 4887
rect 1213 4673 1227 4687
rect 1253 4673 1267 4687
rect 1353 4673 1367 4687
rect 1233 4653 1247 4667
rect 1213 4633 1227 4647
rect 1253 4633 1267 4647
rect 1173 4493 1187 4507
rect 1173 4473 1187 4487
rect 1153 4453 1167 4467
rect 1093 4413 1107 4427
rect 1033 4213 1047 4227
rect 1193 4453 1207 4467
rect 1153 4413 1167 4427
rect 1073 4193 1087 4207
rect 1133 4193 1147 4207
rect 1053 4153 1067 4167
rect 1093 4113 1107 4127
rect 1093 4013 1107 4027
rect 1073 3953 1087 3967
rect 1093 3853 1107 3867
rect 1073 3813 1087 3827
rect 1033 3793 1047 3807
rect 953 3753 967 3767
rect 1013 3753 1027 3767
rect 993 3733 1007 3747
rect 1013 3693 1027 3707
rect 1173 4233 1187 4247
rect 1313 4613 1327 4627
rect 1273 4533 1287 4547
rect 1273 4493 1287 4507
rect 1313 4493 1327 4507
rect 1333 4453 1347 4467
rect 1373 4633 1387 4647
rect 1373 4573 1387 4587
rect 1293 4433 1307 4447
rect 1353 4433 1367 4447
rect 1353 4353 1367 4367
rect 1253 4253 1267 4267
rect 1293 4253 1307 4267
rect 1313 4253 1327 4267
rect 1213 4213 1227 4227
rect 1253 4213 1267 4227
rect 1293 4213 1307 4227
rect 1233 4193 1247 4207
rect 1193 4153 1207 4167
rect 1273 4173 1287 4187
rect 1253 4113 1267 4127
rect 1233 4073 1247 4087
rect 1273 4013 1287 4027
rect 1153 3933 1167 3947
rect 1213 3953 1227 3967
rect 1173 3813 1187 3827
rect 1393 4533 1407 4547
rect 1433 4713 1447 4727
rect 1493 4673 1507 4687
rect 1553 5273 1567 5287
rect 1593 5273 1607 5287
rect 1733 5613 1747 5627
rect 1693 5593 1707 5607
rect 1693 5473 1707 5487
rect 1653 5453 1667 5467
rect 1633 5433 1647 5447
rect 1673 5433 1687 5447
rect 1653 5413 1667 5427
rect 1733 5453 1747 5467
rect 1693 5173 1707 5187
rect 1533 5133 1547 5147
rect 1573 4973 1587 4987
rect 1533 4913 1547 4927
rect 1653 5153 1667 5167
rect 1773 5593 1787 5607
rect 1933 5653 1947 5667
rect 2073 5653 2087 5667
rect 2113 5653 2127 5667
rect 2373 5653 2387 5667
rect 2453 5653 2467 5667
rect 2033 5633 2047 5647
rect 1873 5613 1887 5627
rect 1833 5593 1847 5607
rect 1853 5593 1867 5607
rect 1913 5593 1927 5607
rect 1813 5553 1827 5567
rect 1773 5413 1787 5427
rect 1813 5413 1827 5427
rect 1753 5153 1767 5167
rect 1633 4913 1647 4927
rect 1553 4893 1567 4907
rect 1553 4693 1567 4707
rect 1593 4693 1607 4707
rect 1633 4693 1647 4707
rect 1533 4673 1547 4687
rect 1573 4673 1587 4687
rect 1513 4633 1527 4647
rect 1473 4613 1487 4627
rect 1433 4573 1447 4587
rect 1433 4533 1447 4547
rect 1453 4473 1467 4487
rect 1413 4453 1427 4467
rect 1433 4453 1447 4467
rect 1373 4233 1387 4247
rect 1353 4213 1367 4227
rect 1373 4193 1387 4207
rect 1353 4173 1367 4187
rect 1333 4013 1347 4027
rect 1313 3953 1327 3967
rect 1313 3933 1327 3947
rect 1293 3893 1307 3907
rect 1253 3853 1267 3867
rect 1293 3833 1307 3847
rect 1213 3793 1227 3807
rect 1113 3753 1127 3767
rect 1173 3753 1187 3767
rect 1113 3733 1127 3747
rect 1153 3733 1167 3747
rect 1133 3693 1147 3707
rect 1013 3673 1027 3687
rect 1093 3673 1107 3687
rect 973 3573 987 3587
rect 953 3533 967 3547
rect 913 3513 927 3527
rect 1113 3553 1127 3567
rect 1053 3533 1067 3547
rect 933 3493 947 3507
rect 793 3453 807 3467
rect 913 3473 927 3487
rect 893 3453 907 3467
rect 813 3433 827 3447
rect 873 3433 887 3447
rect 753 3213 767 3227
rect 833 3293 847 3307
rect 873 3253 887 3267
rect 773 3033 787 3047
rect 813 3033 827 3047
rect 873 3193 887 3207
rect 853 3153 867 3167
rect 853 3093 867 3107
rect 653 3013 667 3027
rect 653 2993 667 3007
rect 653 2953 667 2967
rect 533 2753 547 2767
rect 613 2773 627 2787
rect 593 2753 607 2767
rect 553 2733 567 2747
rect 573 2733 587 2747
rect 533 2673 547 2687
rect 533 2573 547 2587
rect 553 2533 567 2547
rect 533 2233 547 2247
rect 453 2213 467 2227
rect 513 2213 527 2227
rect 433 1293 447 1307
rect 473 2173 487 2187
rect 733 3013 747 3027
rect 753 3013 767 3027
rect 793 3013 807 3027
rect 833 3013 847 3027
rect 793 2993 807 3007
rect 753 2973 767 2987
rect 713 2933 727 2947
rect 713 2773 727 2787
rect 653 2753 667 2767
rect 673 2733 687 2747
rect 733 2733 747 2747
rect 773 2793 787 2807
rect 853 2813 867 2827
rect 813 2793 827 2807
rect 793 2773 807 2787
rect 833 2753 847 2767
rect 773 2733 787 2747
rect 753 2713 767 2727
rect 633 2693 647 2707
rect 733 2693 747 2707
rect 673 2673 687 2687
rect 713 2673 727 2687
rect 633 2653 647 2667
rect 653 2573 667 2587
rect 673 2553 687 2567
rect 673 2293 687 2307
rect 573 2213 587 2227
rect 633 2273 647 2287
rect 653 2233 667 2247
rect 633 2213 647 2227
rect 593 2193 607 2207
rect 613 2193 627 2207
rect 573 2133 587 2147
rect 473 2053 487 2067
rect 513 2033 527 2047
rect 513 1873 527 1887
rect 493 1833 507 1847
rect 513 1833 527 1847
rect 533 1813 547 1827
rect 473 1733 487 1747
rect 513 1733 527 1747
rect 513 1713 527 1727
rect 553 1793 567 1807
rect 553 1773 567 1787
rect 553 1713 567 1727
rect 613 2073 627 2087
rect 673 2073 687 2087
rect 913 3253 927 3267
rect 913 3213 927 3227
rect 993 3493 1007 3507
rect 1033 3493 1047 3507
rect 953 3433 967 3447
rect 1033 3353 1047 3367
rect 953 3253 967 3267
rect 993 3253 1007 3267
rect 973 3193 987 3207
rect 973 3173 987 3187
rect 933 3153 947 3167
rect 993 3153 1007 3167
rect 953 3033 967 3047
rect 933 3013 947 3027
rect 973 3013 987 3027
rect 1033 3133 1047 3147
rect 1013 3073 1027 3087
rect 893 2793 907 2807
rect 893 2773 907 2787
rect 933 2773 947 2787
rect 933 2753 947 2767
rect 993 2733 1007 2747
rect 893 2713 907 2727
rect 953 2713 967 2727
rect 873 2673 887 2687
rect 793 2593 807 2607
rect 753 2573 767 2587
rect 873 2573 887 2587
rect 813 2553 827 2567
rect 733 2533 747 2547
rect 773 2533 787 2547
rect 873 2533 887 2547
rect 933 2693 947 2707
rect 993 2593 1007 2607
rect 973 2553 987 2567
rect 913 2533 927 2547
rect 933 2533 947 2547
rect 753 2433 767 2447
rect 893 2433 907 2447
rect 773 2193 787 2207
rect 893 2293 907 2307
rect 813 2273 827 2287
rect 853 2273 867 2287
rect 793 2113 807 2127
rect 793 2093 807 2107
rect 973 2513 987 2527
rect 953 2253 967 2267
rect 913 2133 927 2147
rect 913 2113 927 2127
rect 893 2093 907 2107
rect 753 2073 767 2087
rect 833 2073 847 2087
rect 813 2053 827 2067
rect 773 2033 787 2047
rect 713 2013 727 2027
rect 813 2013 827 2027
rect 653 1933 667 1947
rect 713 1853 727 1867
rect 713 1833 727 1847
rect 593 1793 607 1807
rect 573 1633 587 1647
rect 553 1613 567 1627
rect 493 1573 507 1587
rect 533 1573 547 1587
rect 613 1633 627 1647
rect 593 1553 607 1567
rect 473 1333 487 1347
rect 533 1333 547 1347
rect 493 1313 507 1327
rect 533 1313 547 1327
rect 573 1313 587 1327
rect 513 1293 527 1307
rect 553 1293 567 1307
rect 553 1273 567 1287
rect 453 1253 467 1267
rect 513 1253 527 1267
rect 533 1253 547 1267
rect 473 1233 487 1247
rect 433 1173 447 1187
rect 433 1133 447 1147
rect 493 1093 507 1107
rect 453 1073 467 1087
rect 353 1013 367 1027
rect 393 1013 407 1027
rect 413 1013 427 1027
rect 533 1213 547 1227
rect 533 1073 547 1087
rect 473 953 487 967
rect 513 953 527 967
rect 373 833 387 847
rect 313 813 327 827
rect 433 853 447 867
rect 213 793 227 807
rect 233 793 247 807
rect 273 793 287 807
rect 333 793 347 807
rect 373 793 387 807
rect 393 793 407 807
rect 273 653 287 667
rect 253 613 267 627
rect 293 613 307 627
rect 313 613 327 627
rect 293 413 307 427
rect 213 353 227 367
rect 253 353 267 367
rect 293 353 307 367
rect 253 313 267 327
rect 213 173 227 187
rect 173 153 187 167
rect 313 333 327 347
rect 293 313 307 327
rect 353 713 367 727
rect 453 653 467 667
rect 393 613 407 627
rect 413 593 427 607
rect 453 533 467 547
rect 413 373 427 387
rect 413 353 427 367
rect 453 353 467 367
rect 373 333 387 347
rect 433 313 447 327
rect 333 293 347 307
rect 393 293 407 307
rect 273 253 287 267
rect 373 253 387 267
rect 413 193 427 207
rect 193 133 207 147
rect 73 113 87 127
rect 113 113 127 127
rect 153 113 167 127
rect 173 113 187 127
rect 393 133 407 147
rect 693 1773 707 1787
rect 913 2053 927 2067
rect 853 2033 867 2047
rect 893 2033 907 2047
rect 713 1753 727 1767
rect 833 1793 847 1807
rect 813 1773 827 1787
rect 773 1753 787 1767
rect 933 2013 947 2027
rect 953 2013 967 2027
rect 953 1813 967 1827
rect 933 1793 947 1807
rect 993 2413 1007 2427
rect 1033 3013 1047 3027
rect 1033 2913 1047 2927
rect 1093 3513 1107 3527
rect 1153 3513 1167 3527
rect 1193 3733 1207 3747
rect 1253 3733 1267 3747
rect 1233 3713 1247 3727
rect 1193 3613 1207 3627
rect 1213 3613 1227 3627
rect 1173 3473 1187 3487
rect 1093 3453 1107 3467
rect 1073 3313 1087 3327
rect 1173 3273 1187 3287
rect 1093 3253 1107 3267
rect 1113 3233 1127 3247
rect 1173 3213 1187 3227
rect 1133 3173 1147 3187
rect 1173 3133 1187 3147
rect 1133 3113 1147 3127
rect 1073 3093 1087 3107
rect 1093 3013 1107 3027
rect 1073 2973 1087 2987
rect 1093 2973 1107 2987
rect 1113 2953 1127 2967
rect 1073 2773 1087 2787
rect 1093 2573 1107 2587
rect 1093 2553 1107 2567
rect 1153 3073 1167 3087
rect 1173 3053 1187 3067
rect 1153 2993 1167 3007
rect 1153 2933 1167 2947
rect 1153 2833 1167 2847
rect 1033 2513 1047 2527
rect 1013 2293 1027 2307
rect 1113 2533 1127 2547
rect 1333 3753 1347 3767
rect 1393 3993 1407 4007
rect 1433 4193 1447 4207
rect 1533 4513 1547 4527
rect 1493 4473 1507 4487
rect 1553 4473 1567 4487
rect 1513 4413 1527 4427
rect 1553 4413 1567 4427
rect 1473 4333 1487 4347
rect 1513 4233 1527 4247
rect 1473 4213 1487 4227
rect 1373 3933 1387 3947
rect 1393 3753 1407 3767
rect 1333 3733 1347 3747
rect 1313 3633 1327 3647
rect 1273 3613 1287 3627
rect 1333 3513 1347 3527
rect 1273 3493 1287 3507
rect 1333 3493 1347 3507
rect 1253 3473 1267 3487
rect 1293 3453 1307 3467
rect 1233 3313 1247 3327
rect 1293 3433 1307 3447
rect 1213 3253 1227 3267
rect 1253 3273 1267 3287
rect 1213 3233 1227 3247
rect 1233 3233 1247 3247
rect 1253 3233 1267 3247
rect 1233 3173 1247 3187
rect 1213 3153 1227 3167
rect 1233 3133 1247 3147
rect 1453 3993 1467 4007
rect 1433 3733 1447 3747
rect 1373 3713 1387 3727
rect 1393 3713 1407 3727
rect 1413 3713 1427 3727
rect 1453 3713 1467 3727
rect 1433 3693 1447 3707
rect 1393 3653 1407 3667
rect 1373 3633 1387 3647
rect 1373 3593 1387 3607
rect 1353 3473 1367 3487
rect 1413 3513 1427 3527
rect 1453 3493 1467 3507
rect 1393 3473 1407 3487
rect 1433 3473 1447 3487
rect 1413 3453 1427 3467
rect 1373 3433 1387 3447
rect 1353 3293 1367 3307
rect 1333 3133 1347 3147
rect 1293 3113 1307 3127
rect 1273 3053 1287 3067
rect 1313 3053 1327 3067
rect 1293 3033 1307 3047
rect 1373 3233 1387 3247
rect 1393 3113 1407 3127
rect 1273 2953 1287 2967
rect 1333 3013 1347 3027
rect 1533 4193 1547 4207
rect 1613 4653 1627 4667
rect 1593 4633 1607 4647
rect 1593 4613 1607 4627
rect 1593 4413 1607 4427
rect 1673 5133 1687 5147
rect 1713 5133 1727 5147
rect 1753 5133 1767 5147
rect 1693 5113 1707 5127
rect 1713 4973 1727 4987
rect 1793 5393 1807 5407
rect 1913 5573 1927 5587
rect 1853 5453 1867 5467
rect 1973 5473 1987 5487
rect 1953 5433 1967 5447
rect 2133 5633 2147 5647
rect 2173 5633 2187 5647
rect 2113 5593 2127 5607
rect 2053 5453 2067 5467
rect 2093 5453 2107 5467
rect 1893 5173 1907 5187
rect 1913 5173 1927 5187
rect 1973 5393 1987 5407
rect 2033 5413 2047 5427
rect 2073 5413 2087 5427
rect 2013 5373 2027 5387
rect 2013 5213 2027 5227
rect 1993 5193 2007 5207
rect 1793 5153 1807 5167
rect 1833 5153 1847 5167
rect 1773 5113 1787 5127
rect 1773 5033 1787 5047
rect 1873 5113 1887 5127
rect 1933 5133 1947 5147
rect 1913 5033 1927 5047
rect 1833 4973 1847 4987
rect 1873 4953 1887 4967
rect 1913 4953 1927 4967
rect 2053 5393 2067 5407
rect 2093 5393 2107 5407
rect 2093 5373 2107 5387
rect 2033 5193 2047 5207
rect 2093 5193 2107 5207
rect 2053 5173 2067 5187
rect 2213 5613 2227 5627
rect 2153 5593 2167 5607
rect 2193 5593 2207 5607
rect 2333 5633 2347 5647
rect 2413 5633 2427 5647
rect 2473 5633 2487 5647
rect 2313 5573 2327 5587
rect 2273 5553 2287 5567
rect 2313 5553 2327 5567
rect 2233 5453 2247 5467
rect 2373 5533 2387 5547
rect 2613 5653 2627 5667
rect 2713 5653 2727 5667
rect 2753 5653 2767 5667
rect 2793 5653 2807 5667
rect 2593 5633 2607 5647
rect 2633 5633 2647 5647
rect 2693 5633 2707 5647
rect 2553 5473 2567 5487
rect 2413 5453 2427 5467
rect 2493 5453 2507 5467
rect 2513 5453 2527 5467
rect 2173 5293 2187 5307
rect 2333 5293 2347 5307
rect 2193 5213 2207 5227
rect 2213 5193 2227 5207
rect 2393 5193 2407 5207
rect 2133 5153 2147 5167
rect 2073 5133 2087 5147
rect 2313 5173 2327 5187
rect 2353 5173 2367 5187
rect 2193 5153 2207 5167
rect 2273 5153 2287 5167
rect 2333 5153 2347 5167
rect 2113 5093 2127 5107
rect 2153 5093 2167 5107
rect 2093 5033 2107 5047
rect 1733 4933 1747 4947
rect 1773 4933 1787 4947
rect 1793 4933 1807 4947
rect 1853 4933 1867 4947
rect 1893 4933 1907 4947
rect 1813 4913 1827 4927
rect 1673 4893 1687 4907
rect 1853 4893 1867 4907
rect 1813 4793 1827 4807
rect 1713 4693 1727 4707
rect 1773 4673 1787 4687
rect 1713 4653 1727 4667
rect 1713 4633 1727 4647
rect 1673 4593 1687 4607
rect 1653 4513 1667 4527
rect 1793 4653 1807 4667
rect 1833 4573 1847 4587
rect 1713 4453 1727 4467
rect 1693 4393 1707 4407
rect 1673 4273 1687 4287
rect 1653 4213 1667 4227
rect 1613 4193 1627 4207
rect 1593 4173 1607 4187
rect 1553 4113 1567 4127
rect 1493 4033 1507 4047
rect 1533 4033 1547 4047
rect 1553 4033 1567 4047
rect 1553 3933 1567 3947
rect 1533 3753 1547 3767
rect 1513 3733 1527 3747
rect 1493 3713 1507 3727
rect 1573 3713 1587 3727
rect 1513 3693 1527 3707
rect 1553 3693 1567 3707
rect 1493 3673 1507 3687
rect 1613 4153 1627 4167
rect 1753 4533 1767 4547
rect 1813 4533 1827 4547
rect 1793 4493 1807 4507
rect 1833 4453 1847 4467
rect 1813 4433 1827 4447
rect 1793 4413 1807 4427
rect 1733 4253 1747 4267
rect 1873 4713 1887 4727
rect 1913 4913 1927 4927
rect 1973 4933 1987 4947
rect 1953 4913 1967 4927
rect 2133 4973 2147 4987
rect 2473 5433 2487 5447
rect 2553 5433 2567 5447
rect 2593 5433 2607 5447
rect 2673 5433 2687 5447
rect 2413 5133 2427 5147
rect 2373 5113 2387 5127
rect 2353 5053 2367 5067
rect 2113 4933 2127 4947
rect 2193 4933 2207 4947
rect 2253 4933 2267 4947
rect 2553 5373 2567 5387
rect 2553 5193 2567 5207
rect 2473 5173 2487 5187
rect 2513 5153 2527 5167
rect 2453 5133 2467 5147
rect 2493 5113 2507 5127
rect 2433 5033 2447 5047
rect 2433 5013 2447 5027
rect 2373 4973 2387 4987
rect 2413 4953 2427 4967
rect 2393 4933 2407 4947
rect 1813 4373 1827 4387
rect 1853 4373 1867 4387
rect 1673 4173 1687 4187
rect 1613 4113 1627 4127
rect 1633 4113 1647 4127
rect 1633 4013 1647 4027
rect 1653 4013 1667 4027
rect 1613 3993 1627 4007
rect 1633 3973 1647 3987
rect 1553 3633 1567 3647
rect 1593 3633 1607 3647
rect 1593 3613 1607 3627
rect 1473 3393 1487 3407
rect 1533 3493 1547 3507
rect 1573 3493 1587 3507
rect 1493 3273 1507 3287
rect 1553 3273 1567 3287
rect 1473 3253 1487 3267
rect 1433 3233 1447 3247
rect 1413 2993 1427 3007
rect 1393 2913 1407 2927
rect 1293 2813 1307 2827
rect 1313 2773 1327 2787
rect 1193 2673 1207 2687
rect 1273 2753 1287 2767
rect 1333 2753 1347 2767
rect 1373 2753 1387 2767
rect 1413 2753 1427 2767
rect 1233 2653 1247 2667
rect 1173 2593 1187 2607
rect 1173 2573 1187 2587
rect 1093 2393 1107 2407
rect 1033 2233 1047 2247
rect 1073 2233 1087 2247
rect 1113 2293 1127 2307
rect 1053 2213 1067 2227
rect 1093 2213 1107 2227
rect 1153 2253 1167 2267
rect 993 2053 1007 2067
rect 973 1773 987 1787
rect 1113 2073 1127 2087
rect 1133 2073 1147 2087
rect 1073 2053 1087 2067
rect 1053 2033 1067 2047
rect 1093 2033 1107 2047
rect 1013 1873 1027 1887
rect 1133 1833 1147 1847
rect 1033 1793 1047 1807
rect 993 1753 1007 1767
rect 1033 1753 1047 1767
rect 853 1733 867 1747
rect 953 1733 967 1747
rect 733 1693 747 1707
rect 693 1613 707 1627
rect 733 1613 747 1627
rect 753 1613 767 1627
rect 633 1553 647 1567
rect 933 1653 947 1667
rect 893 1613 907 1627
rect 873 1593 887 1607
rect 773 1573 787 1587
rect 853 1573 867 1587
rect 913 1573 927 1587
rect 753 1533 767 1547
rect 673 1313 687 1327
rect 633 1293 647 1307
rect 653 1253 667 1267
rect 653 1153 667 1167
rect 613 1133 627 1147
rect 613 1113 627 1127
rect 673 1133 687 1147
rect 973 1613 987 1627
rect 973 1573 987 1587
rect 953 1513 967 1527
rect 813 1353 827 1367
rect 913 1353 927 1367
rect 873 1333 887 1347
rect 953 1333 967 1347
rect 793 1293 807 1307
rect 773 1153 787 1167
rect 933 1153 947 1167
rect 1093 1793 1107 1807
rect 1053 1733 1067 1747
rect 1033 1593 1047 1607
rect 1113 1773 1127 1787
rect 1133 1753 1147 1767
rect 1133 1673 1147 1687
rect 1093 1653 1107 1667
rect 1033 1573 1047 1587
rect 1013 1353 1027 1367
rect 1053 1313 1067 1327
rect 1313 2733 1327 2747
rect 1333 2713 1347 2727
rect 1293 2693 1307 2707
rect 1393 2733 1407 2747
rect 1353 2653 1367 2667
rect 1193 2533 1207 2547
rect 1233 2533 1247 2547
rect 1273 2513 1287 2527
rect 1353 2513 1367 2527
rect 1213 2493 1227 2507
rect 1333 2493 1347 2507
rect 1193 2433 1207 2447
rect 1173 2213 1187 2227
rect 1413 2553 1427 2567
rect 1413 2533 1427 2547
rect 1393 2333 1407 2347
rect 1573 3253 1587 3267
rect 1513 3213 1527 3227
rect 1493 3193 1507 3207
rect 1553 3193 1567 3207
rect 1533 3113 1547 3127
rect 1493 3073 1507 3087
rect 1513 3053 1527 3067
rect 1473 2993 1487 3007
rect 1533 3013 1547 3027
rect 1613 3493 1627 3507
rect 1613 3473 1627 3487
rect 1753 4213 1767 4227
rect 1793 4213 1807 4227
rect 1773 4193 1787 4207
rect 1733 4173 1747 4187
rect 1853 4273 1867 4287
rect 1833 4253 1847 4267
rect 1713 4153 1727 4167
rect 1813 4153 1827 4167
rect 1693 4133 1707 4147
rect 1693 3973 1707 3987
rect 1673 3853 1687 3867
rect 1673 3733 1687 3747
rect 1653 3673 1667 3687
rect 1813 4033 1827 4047
rect 1753 4013 1767 4027
rect 2153 4913 2167 4927
rect 2113 4773 2127 4787
rect 1993 4673 2007 4687
rect 1953 4653 1967 4667
rect 1933 4553 1947 4567
rect 2073 4673 2087 4687
rect 2033 4633 2047 4647
rect 1973 4513 1987 4527
rect 2013 4513 2027 4527
rect 1913 4473 1927 4487
rect 1933 4453 1947 4467
rect 2013 4473 2027 4487
rect 2033 4473 2047 4487
rect 2053 4453 2067 4467
rect 2093 4653 2107 4667
rect 2093 4573 2107 4587
rect 2073 4433 2087 4447
rect 2053 4413 2067 4427
rect 1893 4253 1907 4267
rect 1933 4253 1947 4267
rect 1873 4173 1887 4187
rect 1833 4013 1847 4027
rect 1933 4193 1947 4207
rect 1893 4153 1907 4167
rect 1873 3993 1887 4007
rect 1853 3973 1867 3987
rect 1893 3973 1907 3987
rect 1813 3753 1827 3767
rect 1873 3753 1887 3767
rect 1893 3753 1907 3767
rect 1733 3713 1747 3727
rect 1873 3733 1887 3747
rect 1753 3693 1767 3707
rect 1753 3573 1767 3587
rect 1713 3553 1727 3567
rect 1653 3533 1667 3547
rect 1713 3533 1727 3547
rect 1673 3513 1687 3527
rect 1653 3473 1667 3487
rect 1693 3473 1707 3487
rect 1633 3453 1647 3467
rect 1613 3253 1627 3267
rect 1653 3253 1667 3267
rect 1593 3233 1607 3247
rect 1633 3233 1647 3247
rect 1773 3493 1787 3507
rect 1753 3453 1767 3467
rect 1733 3273 1747 3287
rect 1773 3293 1787 3307
rect 1713 3233 1727 3247
rect 1673 3213 1687 3227
rect 1613 3133 1627 3147
rect 1593 3093 1607 3107
rect 1573 3053 1587 3067
rect 1553 2973 1567 2987
rect 1493 2953 1507 2967
rect 1473 2753 1487 2767
rect 1513 2753 1527 2767
rect 1493 2733 1507 2747
rect 1553 2733 1567 2747
rect 1673 3053 1687 3067
rect 1633 3033 1647 3047
rect 1893 3713 1907 3727
rect 2133 4733 2147 4747
rect 2413 4733 2427 4747
rect 2233 4713 2247 4727
rect 2193 4653 2207 4667
rect 2173 4633 2187 4647
rect 2173 4533 2187 4547
rect 2213 4493 2227 4507
rect 2173 4473 2187 4487
rect 2213 4473 2227 4487
rect 2153 4453 2167 4467
rect 2453 4953 2467 4967
rect 2353 4673 2367 4687
rect 2393 4673 2407 4687
rect 2433 4673 2447 4687
rect 2253 4653 2267 4667
rect 2273 4653 2287 4667
rect 2393 4653 2407 4667
rect 2313 4613 2327 4627
rect 2273 4553 2287 4567
rect 2213 4313 2227 4327
rect 2153 4273 2167 4287
rect 2193 4273 2207 4287
rect 2093 4253 2107 4267
rect 2113 4253 2127 4267
rect 2053 4233 2067 4247
rect 1973 4193 1987 4207
rect 2033 4213 2047 4227
rect 2013 4193 2027 4207
rect 2073 4213 2087 4227
rect 2053 4173 2067 4187
rect 1993 4153 2007 4167
rect 1973 4093 1987 4107
rect 2053 4093 2067 4107
rect 1993 4053 2007 4067
rect 2033 4053 2047 4067
rect 1973 3973 1987 3987
rect 1973 3933 1987 3947
rect 2013 3933 2027 3947
rect 1953 3693 1967 3707
rect 2173 4233 2187 4247
rect 2133 4213 2147 4227
rect 2093 4173 2107 4187
rect 2113 4173 2127 4187
rect 2073 3973 2087 3987
rect 2053 3793 2067 3807
rect 2073 3793 2087 3807
rect 1993 3753 2007 3767
rect 2033 3733 2047 3747
rect 2053 3733 2067 3747
rect 1993 3713 2007 3727
rect 1973 3673 1987 3687
rect 2033 3673 2047 3687
rect 1933 3653 1947 3667
rect 1993 3653 2007 3667
rect 1893 3633 1907 3647
rect 1833 3513 1847 3527
rect 1853 3493 1867 3507
rect 1873 3493 1887 3507
rect 1813 3473 1827 3487
rect 1993 3553 2007 3567
rect 1913 3533 1927 3547
rect 1953 3533 1967 3547
rect 2013 3513 2027 3527
rect 1913 3493 1927 3507
rect 1813 3273 1827 3287
rect 1793 3233 1807 3247
rect 1793 3193 1807 3207
rect 1793 3173 1807 3187
rect 1753 3153 1767 3167
rect 1733 3073 1747 3087
rect 1653 3013 1667 3027
rect 1713 3013 1727 3027
rect 1693 2993 1707 3007
rect 1693 2973 1707 2987
rect 1733 2993 1747 3007
rect 1653 2953 1667 2967
rect 1613 2873 1627 2887
rect 1633 2733 1647 2747
rect 1673 2713 1687 2727
rect 1653 2693 1667 2707
rect 1593 2653 1607 2667
rect 1573 2633 1587 2647
rect 1573 2613 1587 2627
rect 1533 2533 1547 2547
rect 1513 2513 1527 2527
rect 1553 2513 1567 2527
rect 1473 2493 1487 2507
rect 1533 2493 1547 2507
rect 1493 2453 1507 2467
rect 1453 2373 1467 2387
rect 1253 2293 1267 2307
rect 1273 2273 1287 2287
rect 1333 2293 1347 2307
rect 1413 2293 1427 2307
rect 1433 2293 1447 2307
rect 1473 2293 1487 2307
rect 1453 2273 1467 2287
rect 1293 2233 1307 2247
rect 1293 2213 1307 2227
rect 1273 2093 1287 2107
rect 1213 2073 1227 2087
rect 1253 2073 1267 2087
rect 1193 2053 1207 2067
rect 1233 2053 1247 2067
rect 1273 2053 1287 2067
rect 1233 1833 1247 1847
rect 1173 1793 1187 1807
rect 1233 1793 1247 1807
rect 1273 1793 1287 1807
rect 1193 1753 1207 1767
rect 1153 1593 1167 1607
rect 1173 1573 1187 1587
rect 1193 1553 1207 1567
rect 1133 1313 1147 1327
rect 1193 1333 1207 1347
rect 1253 1773 1267 1787
rect 1353 2113 1367 2127
rect 1433 2233 1447 2247
rect 1413 2213 1427 2227
rect 1393 2093 1407 2107
rect 1393 2073 1407 2087
rect 1373 2053 1387 2067
rect 1393 1933 1407 1947
rect 1333 1793 1347 1807
rect 1393 1773 1407 1787
rect 1353 1733 1367 1747
rect 1313 1713 1327 1727
rect 1313 1673 1327 1687
rect 1293 1633 1307 1647
rect 1293 1613 1307 1627
rect 1333 1613 1347 1627
rect 1253 1553 1267 1567
rect 1313 1553 1327 1567
rect 1253 1513 1267 1527
rect 1173 1313 1187 1327
rect 1213 1313 1227 1327
rect 1153 1293 1167 1307
rect 1293 1293 1307 1307
rect 1253 1273 1267 1287
rect 1313 1273 1327 1287
rect 1133 1153 1147 1167
rect 893 1133 907 1147
rect 933 1133 947 1147
rect 993 1133 1007 1147
rect 833 1113 847 1127
rect 1053 1113 1067 1127
rect 593 1073 607 1087
rect 633 1073 647 1087
rect 673 1073 687 1087
rect 693 1073 707 1087
rect 633 1013 647 1027
rect 673 1013 687 1027
rect 573 893 587 907
rect 613 893 627 907
rect 553 853 567 867
rect 513 833 527 847
rect 553 833 567 847
rect 773 1093 787 1107
rect 733 893 747 907
rect 673 853 687 867
rect 713 853 727 867
rect 793 853 807 867
rect 493 813 507 827
rect 613 813 627 827
rect 533 793 547 807
rect 653 773 667 787
rect 673 753 687 767
rect 653 653 667 667
rect 533 633 547 647
rect 813 813 827 827
rect 733 773 747 787
rect 773 753 787 767
rect 513 613 527 627
rect 513 533 527 547
rect 593 613 607 627
rect 553 413 567 427
rect 533 353 547 367
rect 473 233 487 247
rect 513 213 527 227
rect 473 133 487 147
rect 673 613 687 627
rect 793 613 807 627
rect 633 593 647 607
rect 873 1093 887 1107
rect 1033 1093 1047 1107
rect 893 1073 907 1087
rect 1113 1093 1127 1107
rect 873 873 887 887
rect 853 833 867 847
rect 673 573 687 587
rect 773 573 787 587
rect 853 593 867 607
rect 733 393 747 407
rect 813 393 827 407
rect 653 333 667 347
rect 793 373 807 387
rect 813 273 827 287
rect 593 253 607 267
rect 573 233 587 247
rect 553 193 567 207
rect 673 193 687 207
rect 533 173 547 187
rect 573 173 587 187
rect 633 173 647 187
rect 553 133 567 147
rect 653 133 667 147
rect 693 133 707 147
rect 1193 1133 1207 1147
rect 1273 1133 1287 1147
rect 1213 1113 1227 1127
rect 1333 1133 1347 1147
rect 1293 1093 1307 1107
rect 1253 1073 1267 1087
rect 1253 1053 1267 1067
rect 1213 873 1227 887
rect 913 833 927 847
rect 953 833 967 847
rect 1013 833 1027 847
rect 893 813 907 827
rect 933 793 947 807
rect 953 773 967 787
rect 933 673 947 687
rect 1013 813 1027 827
rect 973 653 987 667
rect 993 653 1007 667
rect 1073 833 1087 847
rect 1133 853 1147 867
rect 1093 793 1107 807
rect 1033 753 1047 767
rect 1133 833 1147 847
rect 1193 833 1207 847
rect 1213 813 1227 827
rect 1233 793 1247 807
rect 1113 673 1127 687
rect 1093 633 1107 647
rect 973 613 987 627
rect 1013 613 1027 627
rect 953 373 967 387
rect 1073 593 1087 607
rect 1213 673 1227 687
rect 1153 633 1167 647
rect 1293 1033 1307 1047
rect 1513 2273 1527 2287
rect 1493 2253 1507 2267
rect 1613 2533 1627 2547
rect 1653 2633 1667 2647
rect 1653 2593 1667 2607
rect 1693 2593 1707 2607
rect 1633 2513 1647 2527
rect 1573 2493 1587 2507
rect 1553 2473 1567 2487
rect 1633 2353 1647 2367
rect 1593 2313 1607 2327
rect 1553 2273 1567 2287
rect 1513 2213 1527 2227
rect 1473 2133 1487 2147
rect 1513 2093 1527 2107
rect 1473 2073 1487 2087
rect 1493 2053 1507 2067
rect 1533 2053 1547 2067
rect 1473 1973 1487 1987
rect 1573 2233 1587 2247
rect 1613 2213 1627 2227
rect 1593 2133 1607 2147
rect 1573 2113 1587 2127
rect 1573 1933 1587 1947
rect 1653 2333 1667 2347
rect 1693 2553 1707 2567
rect 1833 3133 1847 3147
rect 1833 3033 1847 3047
rect 1773 3013 1787 3027
rect 1813 3013 1827 3027
rect 1813 2753 1827 2767
rect 1773 2733 1787 2747
rect 1833 2713 1847 2727
rect 1753 2693 1767 2707
rect 1793 2693 1807 2707
rect 1773 2653 1787 2667
rect 1753 2533 1767 2547
rect 1713 2493 1727 2507
rect 1693 2453 1707 2467
rect 1733 2473 1747 2487
rect 1733 2453 1747 2467
rect 1713 2333 1727 2347
rect 1713 2293 1727 2307
rect 1753 2353 1767 2367
rect 1713 2273 1727 2287
rect 1733 2273 1747 2287
rect 1693 2253 1707 2267
rect 1733 2233 1747 2247
rect 1753 2233 1767 2247
rect 1753 2213 1767 2227
rect 1713 2193 1727 2207
rect 1693 2093 1707 2107
rect 1653 2073 1667 2087
rect 1673 2073 1687 2087
rect 1633 2053 1647 2067
rect 1673 2053 1687 2067
rect 1653 2033 1667 2047
rect 1693 2033 1707 2047
rect 1613 2013 1627 2027
rect 1673 2013 1687 2027
rect 1633 1793 1647 1807
rect 1433 1753 1447 1767
rect 1413 1733 1427 1747
rect 1373 1713 1387 1727
rect 1433 1673 1447 1687
rect 1373 1593 1387 1607
rect 1393 1493 1407 1507
rect 1373 1413 1387 1427
rect 1493 1773 1507 1787
rect 1533 1773 1547 1787
rect 1553 1773 1567 1787
rect 1513 1753 1527 1767
rect 1493 1733 1507 1747
rect 1453 1613 1467 1627
rect 1473 1553 1487 1567
rect 1453 1333 1467 1347
rect 1433 1153 1447 1167
rect 1373 1133 1387 1147
rect 1373 1093 1387 1107
rect 1413 1073 1427 1087
rect 1453 1073 1467 1087
rect 1353 1033 1367 1047
rect 1333 873 1347 887
rect 1433 873 1447 887
rect 1293 813 1307 827
rect 1133 613 1147 627
rect 1193 613 1207 627
rect 1233 613 1247 627
rect 1193 593 1207 607
rect 1373 853 1387 867
rect 1413 853 1427 867
rect 1353 833 1367 847
rect 1333 733 1347 747
rect 1313 573 1327 587
rect 1233 553 1247 567
rect 1113 533 1127 547
rect 1153 533 1167 547
rect 1013 413 1027 427
rect 833 213 847 227
rect 973 353 987 367
rect 993 353 1007 367
rect 933 333 947 347
rect 973 293 987 307
rect 1033 373 1047 387
rect 1073 373 1087 387
rect 1093 353 1107 367
rect 1053 293 1067 307
rect 1393 653 1407 667
rect 1353 633 1367 647
rect 1413 613 1427 627
rect 1413 573 1427 587
rect 1373 553 1387 567
rect 1353 373 1367 387
rect 1393 373 1407 387
rect 1373 353 1387 367
rect 1253 333 1267 347
rect 1333 333 1347 347
rect 913 213 927 227
rect 1013 213 1027 227
rect 853 193 867 207
rect 833 133 847 147
rect 873 173 887 187
rect 893 173 907 187
rect 873 133 887 147
rect 953 153 967 167
rect 1073 273 1087 287
rect 1193 273 1207 287
rect 1133 193 1147 207
rect 1173 173 1187 187
rect 1233 173 1247 187
rect 1613 1773 1627 1787
rect 1593 1673 1607 1687
rect 1573 1613 1587 1627
rect 1633 1613 1647 1627
rect 1593 1593 1607 1607
rect 1633 1593 1647 1607
rect 1813 2553 1827 2567
rect 1793 2533 1807 2547
rect 1793 2493 1807 2507
rect 2013 3493 2027 3507
rect 1973 3473 1987 3487
rect 1933 3453 1947 3467
rect 1993 3373 2007 3387
rect 1933 3293 1947 3307
rect 1913 3253 1927 3267
rect 1893 3193 1907 3207
rect 1933 3193 1947 3207
rect 1893 3153 1907 3167
rect 1933 3073 1947 3087
rect 1973 3053 1987 3067
rect 1873 3013 1887 3027
rect 1913 3013 1927 3027
rect 1973 2973 1987 2987
rect 1973 2933 1987 2947
rect 1913 2853 1927 2867
rect 1933 2793 1947 2807
rect 2053 3513 2067 3527
rect 2033 3433 2047 3447
rect 2013 3273 2027 3287
rect 2093 3713 2107 3727
rect 2153 4193 2167 4207
rect 2193 4193 2207 4207
rect 2133 4153 2147 4167
rect 2153 4033 2167 4047
rect 2173 4013 2187 4027
rect 2153 3973 2167 3987
rect 2133 3953 2147 3967
rect 2193 3973 2207 3987
rect 2133 3753 2147 3767
rect 2173 3733 2187 3747
rect 2093 3693 2107 3707
rect 2113 3693 2127 3707
rect 2233 4233 2247 4247
rect 2353 4453 2367 4467
rect 2513 4933 2527 4947
rect 2633 5413 2647 5427
rect 2613 5393 2627 5407
rect 2653 5393 2667 5407
rect 2733 5593 2747 5607
rect 2773 5553 2787 5567
rect 2773 5533 2787 5547
rect 2753 5393 2767 5407
rect 2873 5653 2887 5667
rect 3253 5653 3267 5667
rect 3433 5653 3447 5667
rect 3493 5653 3507 5667
rect 3533 5653 3547 5667
rect 4093 5653 4107 5667
rect 4713 5653 4727 5667
rect 4733 5653 4747 5667
rect 2813 5553 2827 5567
rect 2973 5633 2987 5647
rect 3073 5633 3087 5647
rect 3113 5633 3127 5647
rect 2873 5533 2887 5547
rect 2993 5533 3007 5547
rect 2853 5453 2867 5467
rect 2933 5473 2947 5487
rect 2913 5453 2927 5467
rect 2853 5413 2867 5427
rect 2893 5413 2907 5427
rect 3013 5453 3027 5467
rect 3233 5613 3247 5627
rect 3293 5613 3307 5627
rect 3373 5613 3387 5627
rect 3513 5633 3527 5647
rect 3133 5593 3147 5607
rect 3393 5593 3407 5607
rect 3393 5513 3407 5527
rect 3253 5453 3267 5467
rect 3093 5433 3107 5447
rect 3133 5413 3147 5427
rect 3173 5413 3187 5427
rect 3493 5613 3507 5627
rect 3533 5473 3547 5487
rect 3273 5433 3287 5447
rect 3373 5433 3387 5447
rect 3433 5433 3447 5447
rect 3033 5393 3047 5407
rect 3113 5393 3127 5407
rect 3153 5373 3167 5387
rect 2553 5133 2567 5147
rect 2813 5173 2827 5187
rect 2553 5113 2567 5127
rect 2613 5113 2627 5127
rect 2673 5113 2687 5127
rect 2653 5053 2667 5067
rect 2733 5153 2747 5167
rect 2713 5113 2727 5127
rect 2693 5013 2707 5027
rect 2753 4973 2767 4987
rect 2773 4973 2787 4987
rect 2493 4913 2507 4927
rect 2533 4913 2547 4927
rect 2633 4933 2647 4947
rect 2593 4913 2607 4927
rect 2753 4913 2767 4927
rect 2533 4873 2547 4887
rect 2533 4713 2547 4727
rect 2493 4693 2507 4707
rect 2513 4673 2527 4687
rect 2513 4593 2527 4607
rect 2453 4573 2467 4587
rect 2493 4513 2507 4527
rect 2473 4493 2487 4507
rect 2413 4453 2427 4467
rect 2433 4453 2447 4467
rect 2473 4453 2487 4467
rect 2333 4413 2347 4427
rect 2333 4393 2347 4407
rect 2333 4353 2347 4367
rect 2233 4173 2247 4187
rect 2273 4173 2287 4187
rect 2293 4153 2307 4167
rect 2373 4333 2387 4347
rect 2353 4253 2367 4267
rect 2353 4173 2367 4187
rect 2333 4153 2347 4167
rect 2253 4093 2267 4107
rect 2313 4093 2327 4107
rect 2273 4013 2287 4027
rect 2233 3973 2247 3987
rect 2413 4313 2427 4327
rect 2513 4453 2527 4467
rect 2593 4853 2607 4867
rect 2573 4693 2587 4707
rect 2573 4653 2587 4667
rect 2653 4733 2667 4747
rect 2633 4653 2647 4667
rect 2593 4553 2607 4567
rect 2573 4513 2587 4527
rect 2613 4493 2627 4507
rect 2453 4333 2467 4347
rect 2433 4293 2447 4307
rect 2453 4253 2467 4267
rect 2513 4253 2527 4267
rect 2393 4213 2407 4227
rect 2493 4233 2507 4247
rect 2433 4173 2447 4187
rect 2473 4153 2487 4167
rect 2413 4133 2427 4147
rect 2393 4113 2407 4127
rect 2293 3993 2307 4007
rect 2333 3993 2347 4007
rect 2373 3993 2387 4007
rect 2313 3953 2327 3967
rect 2413 4093 2427 4107
rect 2513 4113 2527 4127
rect 2493 4013 2507 4027
rect 2433 3993 2447 4007
rect 2473 3993 2487 4007
rect 2413 3973 2427 3987
rect 2493 3973 2507 3987
rect 2493 3953 2507 3967
rect 2513 3953 2527 3967
rect 2453 3913 2467 3927
rect 2393 3873 2407 3887
rect 2453 3873 2467 3887
rect 2473 3873 2487 3887
rect 2373 3813 2387 3827
rect 2333 3753 2347 3767
rect 2313 3733 2327 3747
rect 2273 3713 2287 3727
rect 2253 3653 2267 3667
rect 2213 3613 2227 3627
rect 2253 3573 2267 3587
rect 2173 3533 2187 3547
rect 2293 3693 2307 3707
rect 2273 3553 2287 3567
rect 2153 3513 2167 3527
rect 2093 3493 2107 3507
rect 2133 3493 2147 3507
rect 2173 3493 2187 3507
rect 2113 3393 2127 3407
rect 2073 3293 2087 3307
rect 2093 3233 2107 3247
rect 2033 3133 2047 3147
rect 2033 3073 2047 3087
rect 2013 3033 2027 3047
rect 2073 3053 2087 3067
rect 2293 3513 2307 3527
rect 2253 3493 2267 3507
rect 2213 3473 2227 3487
rect 2333 3533 2347 3547
rect 2353 3513 2367 3527
rect 2333 3493 2347 3507
rect 2193 3273 2207 3287
rect 2133 3253 2147 3267
rect 2193 3253 2207 3267
rect 2173 3233 2187 3247
rect 2193 3213 2207 3227
rect 2173 3113 2187 3127
rect 2133 3093 2147 3107
rect 2113 3073 2127 3087
rect 2113 3013 2127 3027
rect 2153 2993 2167 3007
rect 2133 2893 2147 2907
rect 2033 2853 2047 2867
rect 2053 2813 2067 2827
rect 2113 2813 2127 2827
rect 1993 2793 2007 2807
rect 1953 2753 1967 2767
rect 2013 2773 2027 2787
rect 1953 2733 1967 2747
rect 1993 2733 2007 2747
rect 1913 2653 1927 2667
rect 1913 2613 1927 2627
rect 1853 2593 1867 2607
rect 1873 2553 1887 2567
rect 1933 2593 1947 2607
rect 1793 2473 1807 2487
rect 1833 2473 1847 2487
rect 1893 2473 1907 2487
rect 1873 2453 1887 2467
rect 1793 2253 1807 2267
rect 1873 2433 1887 2447
rect 1833 2333 1847 2347
rect 1873 2293 1887 2307
rect 1913 2293 1927 2307
rect 1853 2273 1867 2287
rect 1873 2273 1887 2287
rect 1813 2213 1827 2227
rect 1813 2193 1827 2207
rect 1773 2113 1787 2127
rect 1773 2093 1787 2107
rect 1833 2173 1847 2187
rect 1753 2033 1767 2047
rect 1713 1973 1727 1987
rect 1753 1933 1767 1947
rect 1693 1853 1707 1867
rect 1753 1793 1767 1807
rect 1733 1773 1747 1787
rect 1773 1753 1787 1767
rect 1893 2253 1907 2267
rect 1913 2253 1927 2267
rect 1893 2173 1907 2187
rect 1873 2153 1887 2167
rect 1853 2113 1867 2127
rect 1933 2113 1947 2127
rect 1833 2013 1847 2027
rect 1833 1953 1847 1967
rect 1893 2093 1907 2107
rect 1933 2073 1947 2087
rect 1873 2053 1887 2067
rect 1913 2053 1927 2067
rect 1913 1913 1927 1927
rect 1853 1853 1867 1867
rect 1853 1813 1867 1827
rect 1933 1873 1947 1887
rect 1833 1753 1847 1767
rect 1813 1733 1827 1747
rect 1873 1713 1887 1727
rect 1853 1693 1867 1707
rect 1793 1673 1807 1687
rect 1733 1613 1747 1627
rect 1553 1573 1567 1587
rect 1653 1573 1667 1587
rect 1693 1373 1707 1387
rect 1773 1553 1787 1567
rect 1833 1613 1847 1627
rect 1753 1373 1767 1387
rect 1733 1353 1747 1367
rect 1553 1313 1567 1327
rect 1553 1173 1567 1187
rect 1513 1153 1527 1167
rect 1533 1133 1547 1147
rect 1533 1093 1547 1107
rect 1493 1053 1507 1067
rect 1453 853 1467 867
rect 1473 853 1487 867
rect 1453 793 1467 807
rect 1453 693 1467 707
rect 1673 1333 1687 1347
rect 1713 1333 1727 1347
rect 1693 1313 1707 1327
rect 1613 1173 1627 1187
rect 1553 853 1567 867
rect 1573 833 1587 847
rect 1633 1153 1647 1167
rect 1793 1373 1807 1387
rect 1973 2573 1987 2587
rect 2053 2573 2067 2587
rect 2013 2553 2027 2567
rect 2033 2533 2047 2547
rect 1993 2513 2007 2527
rect 1973 2373 1987 2387
rect 2053 2313 2067 2327
rect 2013 2293 2027 2307
rect 2033 2253 2047 2267
rect 1993 2193 2007 2207
rect 1973 2113 1987 2127
rect 2093 2653 2107 2667
rect 2273 3433 2287 3447
rect 2253 3273 2267 3287
rect 2233 3253 2247 3267
rect 2233 3213 2247 3227
rect 2213 3193 2227 3207
rect 2313 3293 2327 3307
rect 2293 3213 2307 3227
rect 2253 3113 2267 3127
rect 2233 3033 2247 3047
rect 2273 3033 2287 3047
rect 2253 3013 2267 3027
rect 2193 2953 2207 2967
rect 2233 2913 2247 2927
rect 2193 2893 2207 2907
rect 2173 2813 2187 2827
rect 2173 2793 2187 2807
rect 2153 2733 2167 2747
rect 2133 2553 2147 2567
rect 2093 2533 2107 2547
rect 2113 2533 2127 2547
rect 2153 2533 2167 2547
rect 2193 2773 2207 2787
rect 2213 2773 2227 2787
rect 2193 2733 2207 2747
rect 2213 2733 2227 2747
rect 2193 2593 2207 2607
rect 2113 2513 2127 2527
rect 2093 2413 2107 2427
rect 2173 2513 2187 2527
rect 2153 2493 2167 2507
rect 2133 2353 2147 2367
rect 2113 2333 2127 2347
rect 2253 2693 2267 2707
rect 2233 2553 2247 2567
rect 2313 3153 2327 3167
rect 2393 3793 2407 3807
rect 2473 3793 2487 3807
rect 2413 3713 2427 3727
rect 2453 3713 2467 3727
rect 2473 3693 2487 3707
rect 2433 3633 2447 3647
rect 2393 3573 2407 3587
rect 2433 3573 2447 3587
rect 2393 3533 2407 3547
rect 2373 3493 2387 3507
rect 2353 3453 2367 3467
rect 2453 3493 2467 3507
rect 2413 3293 2427 3307
rect 2473 3253 2487 3267
rect 2393 3213 2407 3227
rect 2373 3193 2387 3207
rect 2333 3133 2347 3147
rect 2353 3113 2367 3127
rect 2353 3053 2367 3067
rect 2433 3113 2447 3127
rect 2413 3053 2427 3067
rect 2353 3013 2367 3027
rect 2393 3013 2407 3027
rect 2413 3013 2427 3027
rect 2313 2793 2327 2807
rect 2293 2713 2307 2727
rect 2373 2773 2387 2787
rect 2353 2753 2367 2767
rect 2433 2913 2447 2927
rect 2433 2793 2447 2807
rect 2413 2753 2427 2767
rect 2313 2693 2327 2707
rect 2313 2593 2327 2607
rect 2413 2593 2427 2607
rect 2273 2573 2287 2587
rect 2353 2573 2367 2587
rect 2333 2533 2347 2547
rect 2293 2513 2307 2527
rect 2373 2553 2387 2567
rect 2353 2513 2367 2527
rect 2253 2473 2267 2487
rect 2333 2473 2347 2487
rect 2213 2453 2227 2467
rect 2233 2453 2247 2467
rect 2173 2373 2187 2387
rect 2073 2273 2087 2287
rect 2153 2313 2167 2327
rect 2133 2293 2147 2307
rect 2113 2253 2127 2267
rect 2093 2213 2107 2227
rect 1993 2073 2007 2087
rect 2093 2073 2107 2087
rect 2053 2053 2067 2067
rect 2073 2053 2087 2067
rect 2113 2053 2127 2067
rect 2073 2033 2087 2047
rect 2013 1973 2027 1987
rect 1973 1933 1987 1947
rect 1973 1873 1987 1887
rect 1953 1813 1967 1827
rect 2053 1933 2067 1947
rect 1933 1733 1947 1747
rect 1913 1673 1927 1687
rect 1993 1673 2007 1687
rect 2033 1613 2047 1627
rect 2033 1573 2047 1587
rect 2033 1473 2047 1487
rect 1873 1333 1887 1347
rect 1933 1333 1947 1347
rect 1973 1333 1987 1347
rect 2013 1333 2027 1347
rect 1793 1233 1807 1247
rect 1753 1073 1767 1087
rect 1833 1133 1847 1147
rect 1813 993 1827 1007
rect 1633 853 1647 867
rect 1713 853 1727 867
rect 1613 793 1627 807
rect 1533 673 1547 687
rect 1513 653 1527 667
rect 1513 633 1527 647
rect 1533 613 1547 627
rect 1593 613 1607 627
rect 1553 593 1567 607
rect 1473 553 1487 567
rect 1473 393 1487 407
rect 1453 353 1467 367
rect 1733 813 1747 827
rect 1773 833 1787 847
rect 1953 1313 1967 1327
rect 1993 1273 2007 1287
rect 2113 1833 2127 1847
rect 2193 2313 2207 2327
rect 2173 2233 2187 2247
rect 2153 2153 2167 2167
rect 2333 2233 2347 2247
rect 2333 2213 2347 2227
rect 2273 2173 2287 2187
rect 2233 2153 2247 2167
rect 2193 2073 2207 2087
rect 2213 1833 2227 1847
rect 2153 1813 2167 1827
rect 2193 1813 2207 1827
rect 2173 1773 2187 1787
rect 2133 1593 2147 1607
rect 2113 1473 2127 1487
rect 2073 1373 2087 1387
rect 2053 1313 2067 1327
rect 2093 1273 2107 1287
rect 2093 1253 2107 1267
rect 2013 1173 2027 1187
rect 2073 1173 2087 1187
rect 2033 1113 2047 1127
rect 1913 1093 1927 1107
rect 2013 1093 2027 1107
rect 2053 1093 2067 1107
rect 1873 1073 1887 1087
rect 1933 1073 1947 1087
rect 1953 1073 1967 1087
rect 1853 1053 1867 1067
rect 1893 1053 1907 1067
rect 1853 873 1867 887
rect 1893 853 1907 867
rect 1833 833 1847 847
rect 1913 833 1927 847
rect 1813 813 1827 827
rect 1873 813 1887 827
rect 1773 793 1787 807
rect 1753 773 1767 787
rect 1653 653 1667 667
rect 1673 633 1687 647
rect 1713 633 1727 647
rect 1733 633 1747 647
rect 1653 613 1667 627
rect 1693 613 1707 627
rect 1633 413 1647 427
rect 1713 593 1727 607
rect 1513 373 1527 387
rect 1593 373 1607 387
rect 1653 373 1667 387
rect 1693 373 1707 387
rect 1613 353 1627 367
rect 1713 353 1727 367
rect 2073 1053 2087 1067
rect 1973 833 1987 847
rect 2033 853 2047 867
rect 2053 853 2067 867
rect 2013 813 2027 827
rect 1993 773 2007 787
rect 1973 753 1987 767
rect 1953 733 1967 747
rect 1813 693 1827 707
rect 1853 693 1867 707
rect 1813 673 1827 687
rect 1773 613 1787 627
rect 1933 653 1947 667
rect 1993 733 2007 747
rect 1993 653 2007 667
rect 1993 633 2007 647
rect 1853 613 1867 627
rect 1913 613 1927 627
rect 1953 613 1967 627
rect 1993 613 2007 627
rect 1833 593 1847 607
rect 1793 573 1807 587
rect 1833 553 1847 567
rect 1773 373 1787 387
rect 1533 313 1547 327
rect 1613 313 1627 327
rect 1673 333 1687 347
rect 1733 333 1747 347
rect 1633 293 1647 307
rect 1313 173 1327 187
rect 1333 173 1347 187
rect 1273 153 1287 167
rect 1293 153 1307 167
rect 1593 193 1607 207
rect 1433 173 1447 187
rect 1733 173 1747 187
rect 1413 153 1427 167
rect 1193 133 1207 147
rect 1233 133 1247 147
rect 233 113 247 127
rect 833 113 847 127
rect 893 113 907 127
rect 933 113 947 127
rect 953 113 967 127
rect 1033 113 1047 127
rect 1693 153 1707 167
rect 1813 333 1827 347
rect 1793 153 1807 167
rect 1573 133 1587 147
rect 1673 133 1687 147
rect 1713 133 1727 147
rect 1753 133 1767 147
rect 1493 113 1507 127
rect 2073 813 2087 827
rect 2133 1373 2147 1387
rect 2113 1093 2127 1107
rect 2473 3053 2487 3067
rect 2473 2993 2487 3007
rect 2593 4433 2607 4447
rect 2693 4693 2707 4707
rect 2753 4693 2767 4707
rect 2793 4693 2807 4707
rect 2673 4613 2687 4627
rect 2673 4593 2687 4607
rect 2673 4573 2687 4587
rect 2653 4393 2667 4407
rect 2633 4373 2647 4387
rect 2593 4193 2607 4207
rect 2593 4173 2607 4187
rect 2553 4133 2567 4147
rect 2633 4193 2647 4207
rect 2833 5033 2847 5047
rect 2893 5153 2907 5167
rect 2873 5133 2887 5147
rect 2993 5133 3007 5147
rect 3033 5133 3047 5147
rect 2913 5113 2927 5127
rect 3033 5093 3047 5107
rect 2993 5013 3007 5027
rect 2853 4973 2867 4987
rect 2973 4953 2987 4967
rect 2873 4933 2887 4947
rect 2953 4933 2967 4947
rect 2873 4913 2887 4927
rect 3113 5133 3127 5147
rect 3133 5113 3147 5127
rect 3053 4993 3067 5007
rect 3113 4993 3127 5007
rect 3153 4993 3167 5007
rect 3293 5413 3307 5427
rect 3333 5413 3347 5427
rect 3173 4973 3187 4987
rect 3233 4973 3247 4987
rect 3133 4953 3147 4967
rect 2813 4673 2827 4687
rect 2733 4653 2747 4667
rect 2773 4653 2787 4667
rect 2773 4633 2787 4647
rect 2753 4553 2767 4567
rect 2833 4553 2847 4567
rect 2713 4493 2727 4507
rect 3173 4913 3187 4927
rect 3133 4833 3147 4847
rect 3133 4713 3147 4727
rect 2953 4693 2967 4707
rect 3033 4693 3047 4707
rect 3073 4673 3087 4687
rect 2913 4613 2927 4627
rect 3093 4653 3107 4667
rect 2893 4573 2907 4587
rect 3013 4573 3027 4587
rect 2873 4513 2887 4527
rect 2913 4513 2927 4527
rect 2853 4493 2867 4507
rect 2733 4453 2747 4467
rect 2753 4453 2767 4467
rect 2713 4433 2727 4447
rect 2733 4353 2747 4367
rect 2693 4293 2707 4307
rect 2713 4253 2727 4267
rect 2713 4213 2727 4227
rect 2713 4193 2727 4207
rect 2673 4133 2687 4147
rect 2713 4133 2727 4147
rect 2693 4113 2707 4127
rect 2633 3993 2647 4007
rect 2673 3993 2687 4007
rect 2613 3973 2627 3987
rect 2553 3953 2567 3967
rect 2593 3953 2607 3967
rect 2633 3953 2647 3967
rect 2693 3953 2707 3967
rect 2513 3873 2527 3887
rect 2533 3873 2547 3887
rect 2573 3753 2587 3767
rect 2553 3713 2567 3727
rect 2613 3913 2627 3927
rect 2613 3873 2627 3887
rect 2593 3673 2607 3687
rect 2513 3653 2527 3667
rect 2513 3633 2527 3647
rect 2593 3613 2607 3627
rect 2533 3513 2547 3527
rect 2573 3513 2587 3527
rect 2553 3473 2567 3487
rect 2553 3413 2567 3427
rect 2553 3353 2567 3367
rect 2673 3913 2687 3927
rect 2653 3873 2667 3887
rect 2653 3793 2667 3807
rect 2873 4473 2887 4487
rect 2773 4213 2787 4227
rect 2753 4113 2767 4127
rect 2893 4233 2907 4247
rect 2833 4213 2847 4227
rect 2873 4213 2887 4227
rect 3013 4493 3027 4507
rect 2993 4473 3007 4487
rect 2933 4453 2947 4467
rect 2973 4453 2987 4467
rect 2933 4333 2947 4347
rect 2993 4433 3007 4447
rect 3113 4513 3127 4527
rect 3173 4873 3187 4887
rect 3153 4693 3167 4707
rect 3133 4493 3147 4507
rect 3033 4353 3047 4367
rect 2993 4333 3007 4347
rect 3033 4333 3047 4347
rect 2953 4273 2967 4287
rect 2953 4213 2967 4227
rect 3013 4233 3027 4247
rect 2913 4193 2927 4207
rect 2873 4153 2887 4167
rect 2893 4153 2907 4167
rect 2853 4133 2867 4147
rect 2833 4093 2847 4107
rect 2833 4073 2847 4087
rect 2813 4033 2827 4047
rect 2813 3993 2827 4007
rect 2753 3973 2767 3987
rect 2773 3973 2787 3987
rect 2753 3953 2767 3967
rect 2793 3953 2807 3967
rect 2753 3853 2767 3867
rect 2733 3813 2747 3827
rect 2693 3773 2707 3787
rect 2693 3733 2707 3747
rect 2673 3713 2687 3727
rect 2713 3713 2727 3727
rect 2633 3653 2647 3667
rect 2713 3693 2727 3707
rect 2693 3673 2707 3687
rect 2613 3313 2627 3327
rect 2573 3273 2587 3287
rect 2593 3233 2607 3247
rect 2573 3213 2587 3227
rect 2553 3173 2567 3187
rect 2613 3153 2627 3167
rect 2593 3133 2607 3147
rect 2513 3113 2527 3127
rect 2573 3113 2587 3127
rect 2513 3093 2527 3107
rect 2553 3053 2567 3067
rect 2573 3053 2587 3067
rect 2533 3013 2547 3027
rect 2453 2773 2467 2787
rect 2453 2733 2467 2747
rect 2433 2553 2447 2567
rect 2393 2513 2407 2527
rect 2433 2513 2447 2527
rect 2473 2693 2487 2707
rect 2493 2693 2507 2707
rect 2513 2613 2527 2627
rect 2673 3493 2687 3507
rect 2733 3633 2747 3647
rect 2733 3613 2747 3627
rect 2733 3493 2747 3507
rect 2653 3473 2667 3487
rect 2693 3473 2707 3487
rect 2713 3473 2727 3487
rect 2653 3353 2667 3367
rect 2753 3333 2767 3347
rect 2753 3313 2767 3327
rect 2673 3293 2687 3307
rect 2653 3273 2667 3287
rect 2653 3193 2667 3207
rect 2653 3173 2667 3187
rect 2633 3093 2647 3107
rect 2633 3073 2647 3087
rect 2713 3253 2727 3267
rect 2813 3793 2827 3807
rect 2793 3733 2807 3747
rect 2833 3753 2847 3767
rect 2833 3713 2847 3727
rect 2793 3673 2807 3687
rect 2833 3673 2847 3687
rect 2813 3513 2827 3527
rect 2873 4033 2887 4047
rect 2873 4013 2887 4027
rect 2953 4113 2967 4127
rect 2873 3933 2887 3947
rect 2973 4053 2987 4067
rect 3193 4733 3207 4747
rect 3293 5113 3307 5127
rect 3273 5013 3287 5027
rect 3413 5413 3427 5427
rect 3433 5393 3447 5407
rect 3333 5373 3347 5387
rect 3653 5633 3667 5647
rect 3673 5593 3687 5607
rect 3613 5573 3627 5587
rect 3553 5453 3567 5467
rect 3533 5433 3547 5447
rect 3593 5433 3607 5447
rect 3573 5413 3587 5427
rect 3493 5253 3507 5267
rect 3553 5213 3567 5227
rect 3553 5173 3567 5187
rect 3373 5113 3387 5127
rect 3313 4973 3327 4987
rect 3513 5113 3527 5127
rect 3393 4993 3407 5007
rect 3413 4993 3427 5007
rect 3513 4993 3527 5007
rect 3313 4953 3327 4967
rect 3373 4953 3387 4967
rect 3433 4973 3447 4987
rect 3493 4973 3507 4987
rect 3553 5113 3567 5127
rect 3533 4973 3547 4987
rect 3373 4933 3387 4947
rect 3413 4933 3427 4947
rect 3433 4933 3447 4947
rect 3433 4893 3447 4907
rect 3293 4873 3307 4887
rect 3313 4853 3327 4867
rect 3233 4713 3247 4727
rect 3193 4693 3207 4707
rect 3433 4793 3447 4807
rect 3393 4773 3407 4787
rect 3173 4653 3187 4667
rect 3173 4633 3187 4647
rect 3153 4373 3167 4387
rect 3033 4173 3047 4187
rect 3113 4153 3127 4167
rect 3073 4113 3087 4127
rect 3053 4093 3067 4107
rect 2993 4013 3007 4027
rect 3033 4013 3047 4027
rect 2913 3973 2927 3987
rect 2953 3973 2967 3987
rect 2993 3973 3007 3987
rect 2933 3953 2947 3967
rect 2973 3953 2987 3967
rect 2953 3933 2967 3947
rect 3033 3953 3047 3967
rect 3093 4013 3107 4027
rect 3053 3933 3067 3947
rect 2993 3913 3007 3927
rect 2993 3893 3007 3907
rect 3013 3893 3027 3907
rect 2953 3873 2967 3887
rect 2953 3793 2967 3807
rect 2913 3713 2927 3727
rect 2933 3693 2947 3707
rect 2993 3693 3007 3707
rect 2973 3673 2987 3687
rect 2933 3653 2947 3667
rect 2893 3573 2907 3587
rect 2873 3513 2887 3527
rect 2793 3493 2807 3507
rect 2873 3493 2887 3507
rect 2833 3473 2847 3487
rect 2853 3473 2867 3487
rect 2853 3373 2867 3387
rect 2793 3333 2807 3347
rect 2773 3273 2787 3287
rect 2873 3293 2887 3307
rect 2753 3233 2767 3247
rect 2693 3213 2707 3227
rect 2733 3193 2747 3207
rect 2793 3233 2807 3247
rect 2813 3233 2827 3247
rect 2833 3233 2847 3247
rect 2693 3113 2707 3127
rect 2753 3113 2767 3127
rect 2673 3073 2687 3087
rect 2653 3033 2667 3047
rect 2733 3033 2747 3047
rect 2673 2993 2687 3007
rect 2693 2993 2707 3007
rect 2593 2913 2607 2927
rect 2573 2813 2587 2827
rect 2633 2773 2647 2787
rect 2673 2773 2687 2787
rect 2653 2753 2667 2767
rect 2713 2973 2727 2987
rect 2713 2953 2727 2967
rect 2693 2733 2707 2747
rect 2653 2713 2667 2727
rect 2493 2533 2507 2547
rect 2473 2513 2487 2527
rect 2493 2513 2507 2527
rect 2433 2493 2447 2507
rect 2453 2493 2467 2507
rect 2373 2373 2387 2387
rect 2493 2473 2507 2487
rect 2573 2593 2587 2607
rect 2613 2593 2627 2607
rect 2633 2593 2647 2607
rect 2553 2573 2567 2587
rect 2613 2553 2627 2567
rect 2593 2533 2607 2547
rect 2593 2473 2607 2487
rect 2553 2413 2567 2427
rect 2513 2353 2527 2367
rect 2453 2273 2467 2287
rect 2293 2033 2307 2047
rect 2293 1993 2307 2007
rect 2253 1953 2267 1967
rect 2253 1813 2267 1827
rect 2233 1793 2247 1807
rect 2233 1693 2247 1707
rect 2273 1793 2287 1807
rect 2353 2013 2367 2027
rect 2433 2153 2447 2167
rect 2413 2093 2427 2107
rect 2373 1993 2387 2007
rect 2333 1933 2347 1947
rect 2533 2273 2547 2287
rect 2773 3073 2787 3087
rect 2773 3033 2787 3047
rect 2853 3193 2867 3207
rect 2853 3133 2867 3147
rect 2873 3073 2887 3087
rect 2853 3033 2867 3047
rect 2873 3013 2887 3027
rect 2773 2853 2787 2867
rect 2753 2793 2767 2807
rect 2753 2773 2767 2787
rect 2853 2873 2867 2887
rect 2833 2793 2847 2807
rect 2833 2753 2847 2767
rect 2833 2733 2847 2747
rect 2733 2693 2747 2707
rect 2713 2573 2727 2587
rect 2773 2573 2787 2587
rect 2673 2553 2687 2567
rect 2713 2553 2727 2567
rect 2713 2513 2727 2527
rect 2693 2473 2707 2487
rect 2653 2293 2667 2307
rect 2753 2493 2767 2507
rect 2773 2433 2787 2447
rect 2813 2693 2827 2707
rect 2993 3533 3007 3547
rect 2913 3413 2927 3427
rect 2913 3373 2927 3387
rect 2913 3293 2927 3307
rect 3133 4113 3147 4127
rect 3153 4113 3167 4127
rect 3153 4053 3167 4067
rect 3133 4033 3147 4047
rect 3113 3833 3127 3847
rect 3133 3833 3147 3847
rect 3113 3793 3127 3807
rect 3033 3733 3047 3747
rect 3073 3733 3087 3747
rect 3033 3693 3047 3707
rect 3113 3693 3127 3707
rect 3133 3673 3147 3687
rect 3073 3653 3087 3667
rect 3073 3593 3087 3607
rect 3093 3593 3107 3607
rect 3033 3533 3047 3547
rect 3053 3533 3067 3547
rect 3013 3453 3027 3467
rect 3053 3513 3067 3527
rect 3053 3493 3067 3507
rect 3053 3453 3067 3467
rect 3113 3453 3127 3467
rect 3033 3313 3047 3327
rect 2933 3253 2947 3267
rect 2913 3233 2927 3247
rect 3013 3213 3027 3227
rect 2913 3173 2927 3187
rect 2893 2953 2907 2967
rect 2893 2873 2907 2887
rect 2873 2853 2887 2867
rect 2933 3073 2947 3087
rect 2953 3053 2967 3067
rect 2973 3053 2987 3067
rect 2973 3033 2987 3047
rect 2973 2913 2987 2927
rect 2953 2833 2967 2847
rect 2913 2793 2927 2807
rect 2913 2733 2927 2747
rect 2873 2713 2887 2727
rect 2913 2713 2927 2727
rect 2833 2553 2847 2567
rect 2813 2533 2827 2547
rect 2853 2533 2867 2547
rect 2873 2533 2887 2547
rect 2933 2673 2947 2687
rect 2933 2533 2947 2547
rect 2793 2293 2807 2307
rect 2773 2273 2787 2287
rect 2633 2253 2647 2267
rect 2593 2213 2607 2227
rect 2513 2173 2527 2187
rect 2553 2173 2567 2187
rect 2613 2113 2627 2127
rect 2473 2053 2487 2067
rect 2613 2053 2627 2067
rect 2413 1893 2427 1907
rect 2253 1633 2267 1647
rect 2253 1573 2267 1587
rect 2233 1373 2247 1387
rect 2193 1333 2207 1347
rect 2233 1333 2247 1347
rect 2253 1313 2267 1327
rect 2173 1113 2187 1127
rect 2213 1293 2227 1307
rect 2453 1753 2467 1767
rect 2613 1953 2627 1967
rect 2593 1933 2607 1947
rect 2553 1893 2567 1907
rect 2573 1793 2587 1807
rect 2553 1753 2567 1767
rect 2573 1733 2587 1747
rect 2393 1693 2407 1707
rect 2473 1693 2487 1707
rect 2333 1613 2347 1627
rect 2293 1593 2307 1607
rect 2313 1573 2327 1587
rect 2353 1573 2367 1587
rect 2513 1673 2527 1687
rect 2493 1633 2507 1647
rect 2413 1593 2427 1607
rect 2453 1573 2467 1587
rect 2293 1433 2307 1447
rect 2293 1333 2307 1347
rect 2373 1333 2387 1347
rect 2353 1293 2367 1307
rect 2313 1273 2327 1287
rect 2333 1273 2347 1287
rect 2273 1253 2287 1267
rect 2313 1193 2327 1207
rect 2213 1133 2227 1147
rect 2253 1133 2267 1147
rect 2313 1113 2327 1127
rect 2273 1093 2287 1107
rect 2353 1253 2367 1267
rect 2393 1313 2407 1327
rect 2373 1233 2387 1247
rect 2373 1113 2387 1127
rect 2333 1093 2347 1107
rect 2353 1093 2367 1107
rect 2153 1073 2167 1087
rect 2193 1073 2207 1087
rect 2233 913 2247 927
rect 2133 893 2147 907
rect 2213 893 2227 907
rect 2133 853 2147 867
rect 2153 813 2167 827
rect 2113 793 2127 807
rect 2093 753 2107 767
rect 2173 673 2187 687
rect 2093 653 2107 667
rect 2113 653 2127 667
rect 2073 633 2087 647
rect 2053 593 2067 607
rect 2173 573 2187 587
rect 2073 493 2087 507
rect 1913 393 1927 407
rect 1853 373 1867 387
rect 1993 373 2007 387
rect 1913 333 1927 347
rect 2033 353 2047 367
rect 1893 173 1907 187
rect 1913 153 1927 167
rect 1953 133 1967 147
rect 2133 353 2147 367
rect 2293 913 2307 927
rect 2293 893 2307 907
rect 2273 873 2287 887
rect 2253 653 2267 667
rect 2313 793 2327 807
rect 2393 1093 2407 1107
rect 2433 1533 2447 1547
rect 2533 1613 2547 1627
rect 2613 1833 2627 1847
rect 2713 2233 2727 2247
rect 2713 2213 2727 2227
rect 2773 2253 2787 2267
rect 2773 2193 2787 2207
rect 2753 2093 2767 2107
rect 2713 1933 2727 1947
rect 2773 1953 2787 1967
rect 2693 1893 2707 1907
rect 2833 2393 2847 2407
rect 2833 2273 2847 2287
rect 2893 2253 2907 2267
rect 2913 2233 2927 2247
rect 2853 2213 2867 2227
rect 2893 2113 2907 2127
rect 2853 2093 2867 2107
rect 2933 2213 2947 2227
rect 2913 2093 2927 2107
rect 2873 2053 2887 2067
rect 2913 2053 2927 2067
rect 2833 2013 2847 2027
rect 2793 1873 2807 1887
rect 2813 1873 2827 1887
rect 2753 1833 2767 1847
rect 2653 1793 2667 1807
rect 2633 1773 2647 1787
rect 2593 1713 2607 1727
rect 2593 1593 2607 1607
rect 2453 1273 2467 1287
rect 2533 1453 2547 1467
rect 2593 1413 2607 1427
rect 2553 1393 2567 1407
rect 2653 1513 2667 1527
rect 2613 1393 2627 1407
rect 2633 1353 2647 1367
rect 2693 1753 2707 1767
rect 2673 1313 2687 1327
rect 2553 1293 2567 1307
rect 2613 1293 2627 1307
rect 2533 1273 2547 1287
rect 2513 1213 2527 1227
rect 2493 1173 2507 1187
rect 2433 1133 2447 1147
rect 2453 1113 2467 1127
rect 2473 1093 2487 1107
rect 2413 1033 2427 1047
rect 2553 1133 2567 1147
rect 2533 1093 2547 1107
rect 2593 1113 2607 1127
rect 2633 1093 2647 1107
rect 2513 1033 2527 1047
rect 2613 1073 2627 1087
rect 2553 893 2567 907
rect 2513 853 2527 867
rect 2633 853 2647 867
rect 2433 813 2447 827
rect 2373 693 2387 707
rect 2233 633 2247 647
rect 2273 633 2287 647
rect 2433 753 2447 767
rect 2353 593 2367 607
rect 2473 613 2487 627
rect 2333 533 2347 547
rect 2293 493 2307 507
rect 2253 413 2267 427
rect 2213 353 2227 367
rect 2173 193 2187 207
rect 2173 173 2187 187
rect 2113 153 2127 167
rect 2153 153 2167 167
rect 2293 353 2307 367
rect 2353 393 2367 407
rect 2273 333 2287 347
rect 2413 353 2427 367
rect 2493 553 2507 567
rect 2573 833 2587 847
rect 2773 1813 2787 1827
rect 2753 1753 2767 1767
rect 2713 1733 2727 1747
rect 2713 1613 2727 1627
rect 2813 1853 2827 1867
rect 2793 1793 2807 1807
rect 2833 1813 2847 1827
rect 2873 1813 2887 1827
rect 2853 1793 2867 1807
rect 2893 1773 2907 1787
rect 2813 1753 2827 1767
rect 2913 1733 2927 1747
rect 2813 1713 2827 1727
rect 2913 1713 2927 1727
rect 2793 1613 2807 1627
rect 2733 1573 2747 1587
rect 2713 1553 2727 1567
rect 2753 1533 2767 1547
rect 2793 1533 2807 1547
rect 2733 1413 2747 1427
rect 2713 1313 2727 1327
rect 2733 1313 2747 1327
rect 2773 1293 2787 1307
rect 2713 1273 2727 1287
rect 2693 1193 2707 1207
rect 2773 1273 2787 1287
rect 2733 1213 2747 1227
rect 2753 1193 2767 1207
rect 2713 1173 2727 1187
rect 2753 1113 2767 1127
rect 2673 1093 2687 1107
rect 2733 1093 2747 1107
rect 2893 1653 2907 1667
rect 2853 1633 2867 1647
rect 2853 1513 2867 1527
rect 2833 1393 2847 1407
rect 2913 1533 2927 1547
rect 2993 2773 3007 2787
rect 2993 2713 3007 2727
rect 2973 2593 2987 2607
rect 2993 2593 3007 2607
rect 2973 2533 2987 2547
rect 3093 3393 3107 3407
rect 3073 3273 3087 3287
rect 3053 3213 3067 3227
rect 3033 3193 3047 3207
rect 3033 3113 3047 3127
rect 3253 4673 3267 4687
rect 3333 4673 3347 4687
rect 3253 4633 3267 4647
rect 3413 4713 3427 4727
rect 3413 4673 3427 4687
rect 3353 4613 3367 4627
rect 3293 4593 3307 4607
rect 3213 4553 3227 4567
rect 3213 4533 3227 4547
rect 3253 4533 3267 4547
rect 3213 4493 3227 4507
rect 3233 4193 3247 4207
rect 3273 4173 3287 4187
rect 3233 4153 3247 4167
rect 3213 4113 3227 4127
rect 3233 4113 3247 4127
rect 3193 4093 3207 4107
rect 3173 4013 3187 4027
rect 3213 4053 3227 4067
rect 3273 4093 3287 4107
rect 3253 3993 3267 4007
rect 3313 4493 3327 4507
rect 3353 4473 3367 4487
rect 3373 4473 3387 4487
rect 3333 4433 3347 4447
rect 3333 4393 3347 4407
rect 3313 4273 3327 4287
rect 3373 4193 3387 4207
rect 3413 4193 3427 4207
rect 3353 4173 3367 4187
rect 3333 4153 3347 4167
rect 3373 4153 3387 4167
rect 3313 4073 3327 4087
rect 3333 4073 3347 4087
rect 3293 4033 3307 4047
rect 3333 4053 3347 4067
rect 3313 4013 3327 4027
rect 3353 4033 3367 4047
rect 3273 3973 3287 3987
rect 3253 3953 3267 3967
rect 3233 3873 3247 3887
rect 3233 3833 3247 3847
rect 3253 3833 3267 3847
rect 3233 3733 3247 3747
rect 3213 3713 3227 3727
rect 3313 3973 3327 3987
rect 3293 3813 3307 3827
rect 3333 3813 3347 3827
rect 3293 3753 3307 3767
rect 3313 3733 3327 3747
rect 3453 4753 3467 4767
rect 3473 4753 3487 4767
rect 3473 4693 3487 4707
rect 3513 4913 3527 4927
rect 3493 4673 3507 4687
rect 3573 4913 3587 4927
rect 3853 5633 3867 5647
rect 3953 5633 3967 5647
rect 3773 5573 3787 5587
rect 3713 5533 3727 5547
rect 3733 5533 3747 5547
rect 3793 5513 3807 5527
rect 3753 5493 3767 5507
rect 3773 5493 3787 5507
rect 3733 5433 3747 5447
rect 3693 5413 3707 5427
rect 3713 5413 3727 5427
rect 3733 5413 3747 5427
rect 3673 5393 3687 5407
rect 3713 5393 3727 5407
rect 3633 5193 3647 5207
rect 3693 5173 3707 5187
rect 3653 5133 3667 5147
rect 3713 5093 3727 5107
rect 3573 4893 3587 4907
rect 3613 4893 3627 4907
rect 3553 4853 3567 4867
rect 3533 4653 3547 4667
rect 3453 4633 3467 4647
rect 3493 4633 3507 4647
rect 3453 4513 3467 4527
rect 3473 4513 3487 4527
rect 3513 4493 3527 4507
rect 3533 4473 3547 4487
rect 3553 4453 3567 4467
rect 3513 4393 3527 4407
rect 3453 4193 3467 4207
rect 3493 4193 3507 4207
rect 3533 4193 3547 4207
rect 3473 4153 3487 4167
rect 3393 4093 3407 4107
rect 3433 4093 3447 4107
rect 3393 4073 3407 4087
rect 3373 3833 3387 3847
rect 3353 3793 3367 3807
rect 3433 3993 3447 4007
rect 3713 4873 3727 4887
rect 3673 4853 3687 4867
rect 3653 4733 3667 4747
rect 3593 4713 3607 4727
rect 3633 4673 3647 4687
rect 3653 4673 3667 4687
rect 3613 4653 3627 4667
rect 3633 4633 3647 4647
rect 3653 4593 3667 4607
rect 3653 4513 3667 4527
rect 3593 4473 3607 4487
rect 3633 4473 3647 4487
rect 3593 4433 3607 4447
rect 3653 4433 3667 4447
rect 3633 4413 3647 4427
rect 3613 4393 3627 4407
rect 3633 4373 3647 4387
rect 3593 4253 3607 4267
rect 3573 4233 3587 4247
rect 3513 4153 3527 4167
rect 3553 4153 3567 4167
rect 3493 4113 3507 4127
rect 3493 4093 3507 4107
rect 3413 3973 3427 3987
rect 3553 4053 3567 4067
rect 3693 4813 3707 4827
rect 3933 5593 3947 5607
rect 4453 5633 4467 5647
rect 4493 5633 4507 5647
rect 4553 5633 4567 5647
rect 4873 5653 4887 5667
rect 4893 5653 4907 5667
rect 3993 5593 4007 5607
rect 4073 5593 4087 5607
rect 3973 5553 3987 5567
rect 3973 5533 3987 5547
rect 3953 5513 3967 5527
rect 3853 5493 3867 5507
rect 3953 5493 3967 5507
rect 3973 5493 3987 5507
rect 3833 5453 3847 5467
rect 3913 5473 3927 5487
rect 3813 5433 3827 5447
rect 3893 5433 3907 5447
rect 3793 5413 3807 5427
rect 3833 5413 3847 5427
rect 3853 5413 3867 5427
rect 3773 5373 3787 5387
rect 3773 5173 3787 5187
rect 3793 5153 3807 5167
rect 3833 5033 3847 5047
rect 3773 4993 3787 5007
rect 3833 4993 3847 5007
rect 3873 5393 3887 5407
rect 3893 5393 3907 5407
rect 4273 5613 4287 5627
rect 4473 5613 4487 5627
rect 4233 5593 4247 5607
rect 4133 5573 4147 5587
rect 4513 5553 4527 5567
rect 4533 5513 4547 5527
rect 4433 5473 4447 5487
rect 4313 5453 4327 5467
rect 4373 5453 4387 5467
rect 4093 5433 4107 5447
rect 4153 5433 4167 5447
rect 3993 5373 4007 5387
rect 4113 5413 4127 5427
rect 4233 5413 4247 5427
rect 4153 5393 4167 5407
rect 4133 5373 4147 5387
rect 4053 5353 4067 5367
rect 4073 5353 4087 5367
rect 3973 5253 3987 5267
rect 3973 5193 3987 5207
rect 3913 5173 3927 5187
rect 3893 5153 3907 5167
rect 3913 5093 3927 5107
rect 3853 4973 3867 4987
rect 3813 4933 3827 4947
rect 3833 4913 3847 4927
rect 3933 5053 3947 5067
rect 3953 4973 3967 4987
rect 3873 4813 3887 4827
rect 3793 4793 3807 4807
rect 3913 4773 3927 4787
rect 3813 4713 3827 4727
rect 3753 4693 3767 4707
rect 3753 4673 3767 4687
rect 3833 4693 3847 4707
rect 3733 4633 3747 4647
rect 3713 4593 3727 4607
rect 3693 4473 3707 4487
rect 3693 4433 3707 4447
rect 3673 4213 3687 4227
rect 3593 4173 3607 4187
rect 3633 4173 3647 4187
rect 3573 4033 3587 4047
rect 3453 3933 3467 3947
rect 3373 3753 3387 3767
rect 3353 3733 3367 3747
rect 3333 3713 3347 3727
rect 3293 3673 3307 3687
rect 3333 3673 3347 3687
rect 3253 3633 3267 3647
rect 3273 3633 3287 3647
rect 3173 3573 3187 3587
rect 3193 3513 3207 3527
rect 3173 3493 3187 3507
rect 3213 3493 3227 3507
rect 3253 3493 3267 3507
rect 3193 3473 3207 3487
rect 3233 3473 3247 3487
rect 3253 3453 3267 3467
rect 3153 3393 3167 3407
rect 3113 3333 3127 3347
rect 3133 3333 3147 3347
rect 3193 3333 3207 3347
rect 3233 3333 3247 3347
rect 3153 3313 3167 3327
rect 3153 3253 3167 3267
rect 3093 3173 3107 3187
rect 3093 3153 3107 3167
rect 3133 3153 3147 3167
rect 3073 3033 3087 3047
rect 3153 3073 3167 3087
rect 3133 3033 3147 3047
rect 3073 2993 3087 3007
rect 3113 2973 3127 2987
rect 3133 2913 3147 2927
rect 3133 2873 3147 2887
rect 3033 2813 3047 2827
rect 3113 2813 3127 2827
rect 3033 2773 3047 2787
rect 3073 2773 3087 2787
rect 3113 2773 3127 2787
rect 3033 2733 3047 2747
rect 3233 3253 3247 3267
rect 3313 3573 3327 3587
rect 3353 3493 3367 3507
rect 3413 3733 3427 3747
rect 3453 3733 3467 3747
rect 3433 3713 3447 3727
rect 3393 3573 3407 3587
rect 3393 3533 3407 3547
rect 3413 3533 3427 3547
rect 3333 3473 3347 3487
rect 3373 3473 3387 3487
rect 3533 3953 3547 3967
rect 3573 3953 3587 3967
rect 3493 3913 3507 3927
rect 3513 3813 3527 3827
rect 3553 3753 3567 3767
rect 3573 3733 3587 3747
rect 3553 3673 3567 3687
rect 3533 3573 3547 3587
rect 3493 3533 3507 3547
rect 3513 3533 3527 3547
rect 3553 3553 3567 3567
rect 3333 3453 3347 3467
rect 3353 3453 3367 3467
rect 3413 3453 3427 3467
rect 3313 3393 3327 3407
rect 3293 3333 3307 3347
rect 3313 3313 3327 3327
rect 3293 3273 3307 3287
rect 3193 3153 3207 3167
rect 3273 3133 3287 3147
rect 3213 3113 3227 3127
rect 3273 3073 3287 3087
rect 3253 3053 3267 3067
rect 3233 2993 3247 3007
rect 3293 2933 3307 2947
rect 3273 2833 3287 2847
rect 3293 2833 3307 2847
rect 3173 2793 3187 2807
rect 3253 2793 3267 2807
rect 3153 2773 3167 2787
rect 3213 2773 3227 2787
rect 3093 2733 3107 2747
rect 3133 2733 3147 2747
rect 3053 2673 3067 2687
rect 3173 2653 3187 2667
rect 3193 2593 3207 2607
rect 3093 2553 3107 2567
rect 3153 2553 3167 2567
rect 2973 2313 2987 2327
rect 2953 2113 2967 2127
rect 3033 2533 3047 2547
rect 3073 2453 3087 2467
rect 3013 2413 3027 2427
rect 3093 2373 3107 2387
rect 3053 2313 3067 2327
rect 3013 2293 3027 2307
rect 3033 2273 3047 2287
rect 3033 2253 3047 2267
rect 3033 2133 3047 2147
rect 3033 2053 3047 2067
rect 2953 1993 2967 2007
rect 3053 2013 3067 2027
rect 3033 1993 3047 2007
rect 3053 1993 3067 2007
rect 3013 1933 3027 1947
rect 2993 1853 3007 1867
rect 2973 1793 2987 1807
rect 3033 1813 3047 1827
rect 2953 1773 2967 1787
rect 2933 1413 2947 1427
rect 2873 1393 2887 1407
rect 2913 1373 2927 1387
rect 2853 1353 2867 1367
rect 2913 1353 2927 1367
rect 2813 1293 2827 1307
rect 2833 1293 2847 1307
rect 2873 1313 2887 1327
rect 2893 1293 2907 1307
rect 2853 1273 2867 1287
rect 2793 1213 2807 1227
rect 2813 1173 2827 1187
rect 2993 1753 3007 1767
rect 3033 1753 3047 1767
rect 2993 1633 3007 1647
rect 3073 1953 3087 1967
rect 3153 2513 3167 2527
rect 3233 2733 3247 2747
rect 3413 3433 3427 3447
rect 3353 3353 3367 3367
rect 3413 3353 3427 3367
rect 3393 3253 3407 3267
rect 3373 3233 3387 3247
rect 3333 3213 3347 3227
rect 3353 3193 3367 3207
rect 3353 3153 3367 3167
rect 3333 3113 3347 3127
rect 3393 3073 3407 3087
rect 3373 3033 3387 3047
rect 3393 3013 3407 3027
rect 3393 2993 3407 3007
rect 3373 2933 3387 2947
rect 3313 2773 3327 2787
rect 3373 2773 3387 2787
rect 3333 2753 3347 2767
rect 3313 2733 3327 2747
rect 3253 2713 3267 2727
rect 3353 2713 3367 2727
rect 3293 2673 3307 2687
rect 3313 2673 3327 2687
rect 3233 2593 3247 2607
rect 3193 2553 3207 2567
rect 3273 2553 3287 2567
rect 3173 2493 3187 2507
rect 3213 2513 3227 2527
rect 3253 2513 3267 2527
rect 3273 2513 3287 2527
rect 3213 2493 3227 2507
rect 3193 2473 3207 2487
rect 3193 2413 3207 2427
rect 3193 2353 3207 2367
rect 3173 2333 3187 2347
rect 3193 2333 3207 2347
rect 3293 2453 3307 2467
rect 3253 2393 3267 2407
rect 3233 2353 3247 2367
rect 3193 2253 3207 2267
rect 3213 2253 3227 2267
rect 3113 2233 3127 2247
rect 3153 2233 3167 2247
rect 3193 2233 3207 2247
rect 3133 2173 3147 2187
rect 3173 2093 3187 2107
rect 3213 2073 3227 2087
rect 3193 2033 3207 2047
rect 3173 1933 3187 1947
rect 3153 1873 3167 1887
rect 3093 1813 3107 1827
rect 3113 1813 3127 1827
rect 3093 1773 3107 1787
rect 3073 1733 3087 1747
rect 3033 1613 3047 1627
rect 3053 1613 3067 1627
rect 2973 1573 2987 1587
rect 2973 1533 2987 1547
rect 3013 1513 3027 1527
rect 3033 1373 3047 1387
rect 2993 1353 3007 1367
rect 2973 1293 2987 1307
rect 3113 1753 3127 1767
rect 3173 1713 3187 1727
rect 3473 3493 3487 3507
rect 3513 3493 3527 3507
rect 3453 3473 3467 3487
rect 3493 3473 3507 3487
rect 3493 3433 3507 3447
rect 3453 3413 3467 3427
rect 3553 3373 3567 3387
rect 3613 4153 3627 4167
rect 3653 4153 3667 4167
rect 3813 4633 3827 4647
rect 3773 4613 3787 4627
rect 3813 4553 3827 4567
rect 3793 4473 3807 4487
rect 3753 4453 3767 4467
rect 3813 4453 3827 4467
rect 3773 4213 3787 4227
rect 3853 4673 3867 4687
rect 3893 4633 3907 4647
rect 3893 4613 3907 4627
rect 4033 5173 4047 5187
rect 3993 5153 4007 5167
rect 4013 5113 4027 5127
rect 3993 5073 4007 5087
rect 4013 4973 4027 4987
rect 4053 5153 4067 5167
rect 4093 5053 4107 5067
rect 4053 4953 4067 4967
rect 4033 4913 4047 4927
rect 4073 4913 4087 4927
rect 3973 4853 3987 4867
rect 3953 4793 3967 4807
rect 3953 4693 3967 4707
rect 3933 4593 3947 4607
rect 3933 4553 3947 4567
rect 3893 4493 3907 4507
rect 3853 4453 3867 4467
rect 3873 4433 3887 4447
rect 3913 4253 3927 4267
rect 4013 4693 4027 4707
rect 3993 4653 4007 4667
rect 3973 4233 3987 4247
rect 3913 4213 3927 4227
rect 3733 4173 3747 4187
rect 3633 4073 3647 4087
rect 3713 4073 3727 4087
rect 3733 4073 3747 4087
rect 3713 4053 3727 4067
rect 3793 4193 3807 4207
rect 3833 4193 3847 4207
rect 3933 4193 3947 4207
rect 3973 4173 3987 4187
rect 4073 4633 4087 4647
rect 4033 4593 4047 4607
rect 4013 4493 4027 4507
rect 4253 5393 4267 5407
rect 4353 5413 4367 5427
rect 4373 5393 4387 5407
rect 4413 5393 4427 5407
rect 4213 5353 4227 5367
rect 4273 5333 4287 5347
rect 4253 5173 4267 5187
rect 4213 5153 4227 5167
rect 4193 5133 4207 5147
rect 4173 5113 4187 5127
rect 4133 5013 4147 5027
rect 4133 4973 4147 4987
rect 4253 5133 4267 5147
rect 4233 5033 4247 5047
rect 4233 5013 4247 5027
rect 4113 4913 4127 4927
rect 4193 4933 4207 4947
rect 4173 4913 4187 4927
rect 4213 4913 4227 4927
rect 4153 4753 4167 4767
rect 4173 4693 4187 4707
rect 4173 4673 4187 4687
rect 4133 4633 4147 4647
rect 4173 4633 4187 4647
rect 4413 5213 4427 5227
rect 4293 5153 4307 5167
rect 4333 5153 4347 5167
rect 4353 5133 4367 5147
rect 4373 5133 4387 5147
rect 4313 5113 4327 5127
rect 4273 4953 4287 4967
rect 4293 4953 4307 4967
rect 4393 5073 4407 5087
rect 4373 4973 4387 4987
rect 4273 4893 4287 4907
rect 4273 4873 4287 4887
rect 4273 4713 4287 4727
rect 4353 4913 4367 4927
rect 4373 4913 4387 4927
rect 4333 4813 4347 4827
rect 4293 4673 4307 4687
rect 4333 4673 4347 4687
rect 4253 4613 4267 4627
rect 4233 4593 4247 4607
rect 4233 4573 4247 4587
rect 4113 4533 4127 4547
rect 4053 4513 4067 4527
rect 4093 4513 4107 4527
rect 4113 4493 4127 4507
rect 4033 4433 4047 4447
rect 4153 4413 4167 4427
rect 4033 4233 4047 4247
rect 3993 4153 4007 4167
rect 3873 4073 3887 4087
rect 3793 4053 3807 4067
rect 3773 4033 3787 4047
rect 3753 3993 3767 4007
rect 3673 3953 3687 3967
rect 3713 3933 3727 3947
rect 3633 3793 3647 3807
rect 3713 3733 3727 3747
rect 3633 3693 3647 3707
rect 3613 3673 3627 3687
rect 3633 3613 3647 3627
rect 3613 3573 3627 3587
rect 3693 3693 3707 3707
rect 3673 3633 3687 3647
rect 3673 3613 3687 3627
rect 3653 3553 3667 3567
rect 3693 3533 3707 3547
rect 3653 3493 3667 3507
rect 3593 3393 3607 3407
rect 3573 3313 3587 3327
rect 3453 3273 3467 3287
rect 3433 3173 3447 3187
rect 3433 3113 3447 3127
rect 3473 3253 3487 3267
rect 3473 3133 3487 3147
rect 3453 2993 3467 3007
rect 3433 2953 3447 2967
rect 3533 3233 3547 3247
rect 3533 3213 3547 3227
rect 3513 3153 3527 3167
rect 3553 3193 3567 3207
rect 3493 3033 3507 3047
rect 3673 3453 3687 3467
rect 3613 3273 3627 3287
rect 3693 3413 3707 3427
rect 3693 3393 3707 3407
rect 3673 3253 3687 3267
rect 3593 3233 3607 3247
rect 3633 3233 3647 3247
rect 3653 3213 3667 3227
rect 3693 3213 3707 3227
rect 3693 3193 3707 3207
rect 3613 3153 3627 3167
rect 3573 3133 3587 3147
rect 3613 3133 3627 3147
rect 3553 3033 3567 3047
rect 3513 2993 3527 3007
rect 3533 2993 3547 3007
rect 3473 2793 3487 2807
rect 3513 2793 3527 2807
rect 3413 2773 3427 2787
rect 3433 2773 3447 2787
rect 3433 2733 3447 2747
rect 3413 2713 3427 2727
rect 3393 2673 3407 2687
rect 3333 2653 3347 2667
rect 3373 2653 3387 2667
rect 3373 2553 3387 2567
rect 3453 2693 3467 2707
rect 3353 2513 3367 2527
rect 3393 2513 3407 2527
rect 3433 2513 3447 2527
rect 3353 2493 3367 2507
rect 3333 2473 3347 2487
rect 3333 2353 3347 2367
rect 3273 2293 3287 2307
rect 3313 2293 3327 2307
rect 3253 2273 3267 2287
rect 3293 2273 3307 2287
rect 3273 2253 3287 2267
rect 3313 2213 3327 2227
rect 3433 2453 3447 2467
rect 3393 2433 3407 2447
rect 3413 2433 3427 2447
rect 3373 2353 3387 2367
rect 3373 2293 3387 2307
rect 3393 2293 3407 2307
rect 3253 2173 3267 2187
rect 3333 2173 3347 2187
rect 3353 2173 3367 2187
rect 3293 2113 3307 2127
rect 3313 2113 3327 2127
rect 3273 2093 3287 2107
rect 3253 2073 3267 2087
rect 3233 2053 3247 2067
rect 3273 2053 3287 2067
rect 3253 1973 3267 1987
rect 3213 1793 3227 1807
rect 3193 1673 3207 1687
rect 3353 2093 3367 2107
rect 3313 2033 3327 2047
rect 3333 2033 3347 2047
rect 3313 1813 3327 1827
rect 3293 1773 3307 1787
rect 3293 1733 3307 1747
rect 3253 1713 3267 1727
rect 3513 2733 3527 2747
rect 3493 2713 3507 2727
rect 3473 2673 3487 2687
rect 3473 2653 3487 2667
rect 3473 2553 3487 2567
rect 3473 2473 3487 2487
rect 3453 2353 3467 2367
rect 3413 2273 3427 2287
rect 3473 2313 3487 2327
rect 3393 2213 3407 2227
rect 3393 2173 3407 2187
rect 3413 2173 3427 2187
rect 3433 2153 3447 2167
rect 3373 1833 3387 1847
rect 3373 1813 3387 1827
rect 3413 1813 3427 1827
rect 3353 1773 3367 1787
rect 3313 1673 3327 1687
rect 3113 1593 3127 1607
rect 3113 1573 3127 1587
rect 3113 1533 3127 1547
rect 3213 1653 3227 1667
rect 3233 1653 3247 1667
rect 3133 1513 3147 1527
rect 3233 1633 3247 1647
rect 3233 1573 3247 1587
rect 3393 1793 3407 1807
rect 3393 1753 3407 1767
rect 3413 1693 3427 1707
rect 3693 3113 3707 3127
rect 3653 3053 3667 3067
rect 3633 3033 3647 3047
rect 3673 2993 3687 3007
rect 3733 3713 3747 3727
rect 3733 3653 3747 3667
rect 3833 3973 3847 3987
rect 3893 4033 3907 4047
rect 3853 3933 3867 3947
rect 3773 3913 3787 3927
rect 3813 3833 3827 3847
rect 3773 3733 3787 3747
rect 3833 3753 3847 3767
rect 3793 3653 3807 3667
rect 3833 3653 3847 3667
rect 3773 3573 3787 3587
rect 3713 2833 3727 2847
rect 3753 3513 3767 3527
rect 3773 3473 3787 3487
rect 3833 3493 3847 3507
rect 3793 3453 3807 3467
rect 3833 3393 3847 3407
rect 3833 3233 3847 3247
rect 3833 3213 3847 3227
rect 3773 3153 3787 3167
rect 3793 3153 3807 3167
rect 3753 3053 3767 3067
rect 3773 3013 3787 3027
rect 3653 2793 3667 2807
rect 3733 2793 3747 2807
rect 3593 2733 3607 2747
rect 3613 2733 3627 2747
rect 3573 2713 3587 2727
rect 3593 2693 3607 2707
rect 3553 2673 3567 2687
rect 3533 2653 3547 2667
rect 3573 2653 3587 2667
rect 3513 2493 3527 2507
rect 3493 2253 3507 2267
rect 3493 2233 3507 2247
rect 3473 2113 3487 2127
rect 3453 2073 3467 2087
rect 3453 1973 3467 1987
rect 3433 1553 3447 1567
rect 3253 1473 3267 1487
rect 3273 1473 3287 1487
rect 3113 1393 3127 1407
rect 3053 1353 3067 1367
rect 3193 1353 3207 1367
rect 3013 1313 3027 1327
rect 3153 1313 3167 1327
rect 3033 1293 3047 1307
rect 3033 1273 3047 1287
rect 2953 1173 2967 1187
rect 2773 1093 2787 1107
rect 2893 1113 2907 1127
rect 2873 1033 2887 1047
rect 2953 1133 2967 1147
rect 2933 1113 2947 1127
rect 2993 1173 3007 1187
rect 2973 1073 2987 1087
rect 2913 973 2927 987
rect 2973 933 2987 947
rect 2933 873 2947 887
rect 2773 833 2787 847
rect 2673 813 2687 827
rect 2733 813 2747 827
rect 2853 853 2867 867
rect 2893 853 2907 867
rect 2693 773 2707 787
rect 2813 773 2827 787
rect 2653 753 2667 767
rect 2733 653 2747 667
rect 2613 613 2627 627
rect 2593 533 2607 547
rect 2733 613 2747 627
rect 2693 533 2707 547
rect 2633 513 2647 527
rect 2593 433 2607 447
rect 2533 413 2547 427
rect 2453 333 2467 347
rect 2313 313 2327 327
rect 2353 313 2367 327
rect 2433 313 2447 327
rect 2373 293 2387 307
rect 2253 173 2267 187
rect 1933 113 1947 127
rect 1973 113 1987 127
rect 2073 113 2087 127
rect 2133 113 2147 127
rect 193 93 207 107
rect 793 93 807 107
rect 1853 93 1867 107
rect 2093 93 2107 107
rect 2333 153 2347 167
rect 2453 153 2467 167
rect 2553 373 2567 387
rect 2533 353 2547 367
rect 2653 453 2667 467
rect 2633 393 2647 407
rect 2713 393 2727 407
rect 2573 313 2587 327
rect 2673 333 2687 347
rect 2693 333 2707 347
rect 2633 293 2647 307
rect 2873 653 2887 667
rect 2833 613 2847 627
rect 2793 573 2807 587
rect 2773 513 2787 527
rect 2793 513 2807 527
rect 2733 353 2747 367
rect 3013 833 3027 847
rect 3053 1133 3067 1147
rect 3133 1293 3147 1307
rect 3073 1113 3087 1127
rect 3113 1113 3127 1127
rect 3093 1073 3107 1087
rect 3193 1233 3207 1247
rect 3173 1213 3187 1227
rect 3153 1153 3167 1167
rect 3153 1073 3167 1087
rect 3133 1053 3147 1067
rect 3113 873 3127 887
rect 3053 833 3067 847
rect 2953 793 2967 807
rect 2993 793 3007 807
rect 2913 453 2927 467
rect 2833 413 2847 427
rect 2753 333 2767 347
rect 2513 193 2527 207
rect 2713 193 2727 207
rect 2653 173 2667 187
rect 2613 153 2627 167
rect 2873 373 2887 387
rect 2873 333 2887 347
rect 2933 333 2947 347
rect 2833 313 2847 327
rect 2893 313 2907 327
rect 2913 313 2927 327
rect 2913 153 2927 167
rect 2633 133 2647 147
rect 2673 133 2687 147
rect 2713 133 2727 147
rect 2833 133 2847 147
rect 2393 113 2407 127
rect 2473 113 2487 127
rect 2933 113 2947 127
rect 2773 93 2787 107
rect 2893 93 2907 107
rect 2273 33 2287 47
rect 2673 33 2687 47
rect 2633 13 2647 27
rect 3033 633 3047 647
rect 2993 613 3007 627
rect 2973 593 2987 607
rect 3013 593 3027 607
rect 2973 533 2987 547
rect 3013 353 3027 367
rect 2993 313 3007 327
rect 3133 833 3147 847
rect 3173 833 3187 847
rect 3113 793 3127 807
rect 3153 793 3167 807
rect 3093 653 3107 667
rect 3133 633 3147 647
rect 3153 633 3167 647
rect 3073 613 3087 627
rect 3113 613 3127 627
rect 3093 573 3107 587
rect 3053 393 3067 407
rect 3213 1173 3227 1187
rect 3293 1393 3307 1407
rect 3433 1493 3447 1507
rect 3413 1293 3427 1307
rect 3273 1273 3287 1287
rect 3313 1273 3327 1287
rect 3373 1233 3387 1247
rect 3413 1213 3427 1227
rect 3373 1153 3387 1167
rect 3253 1133 3267 1147
rect 3393 1133 3407 1147
rect 3233 1093 3247 1107
rect 3193 653 3207 667
rect 3313 1113 3327 1127
rect 3273 1053 3287 1067
rect 3253 913 3267 927
rect 3293 853 3307 867
rect 3273 773 3287 787
rect 3333 1033 3347 1047
rect 3633 2673 3647 2687
rect 3693 2773 3707 2787
rect 3713 2753 3727 2767
rect 3753 2753 3767 2767
rect 3673 2733 3687 2747
rect 3733 2733 3747 2747
rect 3673 2713 3687 2727
rect 3653 2553 3667 2567
rect 3613 2513 3627 2527
rect 3573 2473 3587 2487
rect 3573 2293 3587 2307
rect 3533 2253 3547 2267
rect 3573 2253 3587 2267
rect 3513 2193 3527 2207
rect 3593 2173 3607 2187
rect 3533 2093 3547 2107
rect 3573 2093 3587 2107
rect 3513 2053 3527 2067
rect 3553 2053 3567 2067
rect 3693 2673 3707 2687
rect 3673 2493 3687 2507
rect 3653 2473 3667 2487
rect 3673 2393 3687 2407
rect 3633 2373 3647 2387
rect 3653 2373 3667 2387
rect 3633 2253 3647 2267
rect 3773 2733 3787 2747
rect 3713 2573 3727 2587
rect 3753 2573 3767 2587
rect 3833 3053 3847 3067
rect 3813 3033 3827 3047
rect 3833 3013 3847 3027
rect 3813 2933 3827 2947
rect 3833 2893 3847 2907
rect 3933 3993 3947 4007
rect 3973 3993 3987 4007
rect 4013 3993 4027 4007
rect 3893 3813 3907 3827
rect 3913 3773 3927 3787
rect 3893 3633 3907 3647
rect 3893 3613 3907 3627
rect 3873 3593 3887 3607
rect 3873 3513 3887 3527
rect 3913 3513 3927 3527
rect 3913 3373 3927 3387
rect 3893 3233 3907 3247
rect 3873 3193 3887 3207
rect 3913 3193 3927 3207
rect 3913 3173 3927 3187
rect 3873 3073 3887 3087
rect 3873 3033 3887 3047
rect 3893 3033 3907 3047
rect 3893 2993 3907 3007
rect 3873 2973 3887 2987
rect 3853 2813 3867 2827
rect 3873 2813 3887 2827
rect 3813 2773 3827 2787
rect 3793 2693 3807 2707
rect 3833 2633 3847 2647
rect 3833 2613 3847 2627
rect 3813 2573 3827 2587
rect 3793 2533 3807 2547
rect 3733 2513 3747 2527
rect 3753 2513 3767 2527
rect 3793 2513 3807 2527
rect 3713 2433 3727 2447
rect 3693 2373 3707 2387
rect 3773 2473 3787 2487
rect 3753 2353 3767 2367
rect 3733 2273 3747 2287
rect 3673 2253 3687 2267
rect 3693 2253 3707 2267
rect 3653 2233 3667 2247
rect 3653 2213 3667 2227
rect 3633 2073 3647 2087
rect 3553 2033 3567 2047
rect 3613 2033 3627 2047
rect 3593 2013 3607 2027
rect 3493 1913 3507 1927
rect 3533 1913 3547 1927
rect 3493 1853 3507 1867
rect 3493 1793 3507 1807
rect 3573 1813 3587 1827
rect 3473 1733 3487 1747
rect 3473 1693 3487 1707
rect 3473 1553 3487 1567
rect 3473 1533 3487 1547
rect 3453 1453 3467 1467
rect 3453 1373 3467 1387
rect 3453 1293 3467 1307
rect 3453 1273 3467 1287
rect 3433 1193 3447 1207
rect 3433 1133 3447 1147
rect 3433 1013 3447 1027
rect 3413 833 3427 847
rect 3393 813 3407 827
rect 3333 793 3347 807
rect 3413 793 3427 807
rect 3433 773 3447 787
rect 3373 653 3387 667
rect 3413 653 3427 667
rect 3173 613 3187 627
rect 3153 533 3167 547
rect 3173 453 3187 467
rect 3133 413 3147 427
rect 3253 613 3267 627
rect 3233 593 3247 607
rect 3293 613 3307 627
rect 3253 553 3267 567
rect 3213 393 3227 407
rect 3333 613 3347 627
rect 3313 413 3327 427
rect 3153 353 3167 367
rect 3173 353 3187 367
rect 3253 353 3267 367
rect 3153 313 3167 327
rect 3273 313 3287 327
rect 3353 593 3367 607
rect 3353 553 3367 567
rect 3413 393 3427 407
rect 3553 1673 3567 1687
rect 3553 1613 3567 1627
rect 3533 1593 3547 1607
rect 3513 1533 3527 1547
rect 3533 1533 3547 1547
rect 3513 1513 3527 1527
rect 3493 1373 3507 1387
rect 3493 1213 3507 1227
rect 3473 1193 3487 1207
rect 3493 1173 3507 1187
rect 3533 1473 3547 1487
rect 3533 1433 3547 1447
rect 3533 1293 3547 1307
rect 3673 2093 3687 2107
rect 3653 2013 3667 2027
rect 3713 2053 3727 2067
rect 3673 1993 3687 2007
rect 3713 1973 3727 1987
rect 3633 1933 3647 1947
rect 3613 1893 3627 1907
rect 3613 1833 3627 1847
rect 3613 1773 3627 1787
rect 3693 1893 3707 1907
rect 3633 1753 3647 1767
rect 3653 1753 3667 1767
rect 3653 1733 3667 1747
rect 3633 1713 3647 1727
rect 3593 1613 3607 1627
rect 3713 1773 3727 1787
rect 3693 1713 3707 1727
rect 3673 1673 3687 1687
rect 3673 1613 3687 1627
rect 3593 1593 3607 1607
rect 3653 1573 3667 1587
rect 3613 1553 3627 1567
rect 3593 1533 3607 1547
rect 3573 1253 3587 1267
rect 3733 1653 3747 1667
rect 3813 2493 3827 2507
rect 3813 2413 3827 2427
rect 3793 2293 3807 2307
rect 3773 2233 3787 2247
rect 3793 2193 3807 2207
rect 3853 2573 3867 2587
rect 3853 2533 3867 2547
rect 3853 2513 3867 2527
rect 3853 2333 3867 2347
rect 3833 2293 3847 2307
rect 3833 2233 3847 2247
rect 3773 2173 3787 2187
rect 3813 2173 3827 2187
rect 3953 3973 3967 3987
rect 3993 3973 4007 3987
rect 4093 4233 4107 4247
rect 4053 4213 4067 4227
rect 4133 4213 4147 4227
rect 4053 4173 4067 4187
rect 3993 3953 4007 3967
rect 4033 3953 4047 3967
rect 4013 3713 4027 3727
rect 4313 4533 4327 4547
rect 4253 4473 4267 4487
rect 4233 4293 4247 4307
rect 4173 4253 4187 4267
rect 4193 4253 4207 4267
rect 4193 4193 4207 4207
rect 4193 4173 4207 4187
rect 4233 4173 4247 4187
rect 4153 4093 4167 4107
rect 4093 4053 4107 4067
rect 4133 4053 4147 4067
rect 4173 4053 4187 4067
rect 4073 3993 4087 4007
rect 4133 4033 4147 4047
rect 4113 3973 4127 3987
rect 4293 4453 4307 4467
rect 4273 4433 4287 4447
rect 4353 4453 4367 4467
rect 4273 4393 4287 4407
rect 4313 4393 4327 4407
rect 4333 4393 4347 4407
rect 4273 4373 4287 4387
rect 4253 4033 4267 4047
rect 4233 3973 4247 3987
rect 4193 3933 4207 3947
rect 4213 3933 4227 3947
rect 4253 3833 4267 3847
rect 4133 3713 4147 3727
rect 4073 3693 4087 3707
rect 3993 3633 4007 3647
rect 3973 3613 3987 3627
rect 3993 3513 4007 3527
rect 3973 3473 3987 3487
rect 3993 3373 4007 3387
rect 3953 3253 3967 3267
rect 3953 3233 3967 3247
rect 4133 3653 4147 3667
rect 4033 3613 4047 3627
rect 4153 3593 4167 3607
rect 4213 3693 4227 3707
rect 4193 3573 4207 3587
rect 4193 3553 4207 3567
rect 4053 3533 4067 3547
rect 4153 3533 4167 3547
rect 4033 3493 4047 3507
rect 4113 3493 4127 3507
rect 4173 3493 4187 3507
rect 4013 3353 4027 3367
rect 4013 3253 4027 3267
rect 3993 3153 4007 3167
rect 3933 3133 3947 3147
rect 3973 3133 3987 3147
rect 3933 3033 3947 3047
rect 3953 2973 3967 2987
rect 3993 3053 4007 3067
rect 3993 3033 4007 3047
rect 4033 3153 4047 3167
rect 4173 3473 4187 3487
rect 4073 3453 4087 3467
rect 4153 3333 4167 3347
rect 4133 3313 4147 3327
rect 4093 3233 4107 3247
rect 4073 3173 4087 3187
rect 4073 3113 4087 3127
rect 4053 3053 4067 3067
rect 4093 3053 4107 3067
rect 4033 3033 4047 3047
rect 4013 2893 4027 2907
rect 4013 2873 4027 2887
rect 3933 2793 3947 2807
rect 3973 2793 3987 2807
rect 3993 2793 4007 2807
rect 3913 2693 3927 2707
rect 3913 2573 3927 2587
rect 3893 2553 3907 2567
rect 3993 2773 4007 2787
rect 4013 2773 4027 2787
rect 3973 2753 3987 2767
rect 3993 2673 4007 2687
rect 3973 2653 3987 2667
rect 3953 2633 3967 2647
rect 3913 2533 3927 2547
rect 3893 2273 3907 2287
rect 3793 2073 3807 2087
rect 3833 2073 3847 2087
rect 3833 2053 3847 2067
rect 3813 2033 3827 2047
rect 3773 2013 3787 2027
rect 3793 1873 3807 1887
rect 3773 1773 3787 1787
rect 3773 1733 3787 1747
rect 3753 1633 3767 1647
rect 3753 1613 3767 1627
rect 3713 1593 3727 1607
rect 3693 1573 3707 1587
rect 3733 1573 3747 1587
rect 3773 1573 3787 1587
rect 3673 1553 3687 1567
rect 3733 1533 3747 1547
rect 3853 1833 3867 1847
rect 3833 1773 3847 1787
rect 3813 1753 3827 1767
rect 3833 1593 3847 1607
rect 3933 2493 3947 2507
rect 3953 2333 3967 2347
rect 4113 2973 4127 2987
rect 4093 2753 4107 2767
rect 4073 2713 4087 2727
rect 4113 2713 4127 2727
rect 4413 4933 4427 4947
rect 4493 5453 4507 5467
rect 4573 5593 4587 5607
rect 4813 5593 4827 5607
rect 4853 5593 4867 5607
rect 4573 5513 4587 5527
rect 4553 5493 4567 5507
rect 4713 5493 4727 5507
rect 4593 5433 4607 5447
rect 4753 5453 4767 5467
rect 4473 5413 4487 5427
rect 4513 5413 4527 5427
rect 4633 5413 4647 5427
rect 4513 5393 4527 5407
rect 4553 5393 4567 5407
rect 4733 5393 4747 5407
rect 4473 5353 4487 5367
rect 4473 5153 4487 5167
rect 4533 5133 4547 5147
rect 4453 5113 4467 5127
rect 4453 4973 4467 4987
rect 4493 4953 4507 4967
rect 4433 4873 4447 4887
rect 4673 5253 4687 5267
rect 4573 5193 4587 5207
rect 4593 5133 4607 5147
rect 4633 5153 4647 5167
rect 4653 5133 4667 5147
rect 4613 5113 4627 5127
rect 4613 5033 4627 5047
rect 4653 5033 4667 5047
rect 4593 4973 4607 4987
rect 4633 4953 4647 4967
rect 4693 5153 4707 5167
rect 4733 5153 4747 5167
rect 4793 5353 4807 5367
rect 4713 5113 4727 5127
rect 4753 5113 4767 5127
rect 4713 5033 4727 5047
rect 4553 4913 4567 4927
rect 4613 4913 4627 4927
rect 4613 4833 4627 4847
rect 4493 4813 4507 4827
rect 4593 4813 4607 4827
rect 4413 4713 4427 4727
rect 4493 4713 4507 4727
rect 4413 4693 4427 4707
rect 4433 4673 4447 4687
rect 4473 4673 4487 4687
rect 4453 4633 4467 4647
rect 4473 4533 4487 4547
rect 4473 4513 4487 4527
rect 4393 4473 4407 4487
rect 4413 4473 4427 4487
rect 4393 4453 4407 4467
rect 4433 4433 4447 4447
rect 4373 4413 4387 4427
rect 4533 4673 4547 4687
rect 4533 4593 4547 4607
rect 4573 4653 4587 4667
rect 4593 4633 4607 4647
rect 4553 4573 4567 4587
rect 4493 4433 4507 4447
rect 4513 4433 4527 4447
rect 4333 4193 4347 4207
rect 4313 4173 4327 4187
rect 4473 4193 4487 4207
rect 4393 4173 4407 4187
rect 4433 4173 4447 4187
rect 4373 4153 4387 4167
rect 4413 4153 4427 4167
rect 4693 4733 4707 4747
rect 4693 4673 4707 4687
rect 4673 4633 4687 4647
rect 4613 4353 4627 4367
rect 4653 4353 4667 4367
rect 4593 4333 4607 4347
rect 4553 4293 4567 4307
rect 4613 4293 4627 4307
rect 4553 4213 4567 4227
rect 4593 4213 4607 4227
rect 4493 4133 4507 4147
rect 4293 4113 4307 4127
rect 4333 4113 4347 4127
rect 4393 4113 4407 4127
rect 4293 4093 4307 4107
rect 4373 4033 4387 4047
rect 4333 3993 4347 4007
rect 4353 3973 4367 3987
rect 4393 3973 4407 3987
rect 4433 3973 4447 3987
rect 4413 3893 4427 3907
rect 4333 3873 4347 3887
rect 4373 3873 4387 3887
rect 4293 3573 4307 3587
rect 4213 3533 4227 3547
rect 4213 3313 4227 3327
rect 4273 3553 4287 3567
rect 4253 3533 4267 3547
rect 4373 3713 4387 3727
rect 4433 3733 4447 3747
rect 4513 3993 4527 4007
rect 4533 3993 4547 4007
rect 4473 3913 4487 3927
rect 4613 4193 4627 4207
rect 4573 4113 4587 4127
rect 4693 4393 4707 4407
rect 4733 4953 4747 4967
rect 4833 5333 4847 5347
rect 4873 5333 4887 5347
rect 4833 5133 4847 5147
rect 4873 5133 4887 5147
rect 4833 5093 4847 5107
rect 4853 5073 4867 5087
rect 5153 5753 5167 5767
rect 5133 5673 5147 5687
rect 4933 5593 4947 5607
rect 4913 5513 4927 5527
rect 4993 5613 5007 5627
rect 5053 5613 5067 5627
rect 5133 5613 5147 5627
rect 4933 5093 4947 5107
rect 4913 5053 4927 5067
rect 4893 5033 4907 5047
rect 4893 4993 4907 5007
rect 4773 4933 4787 4947
rect 4733 4633 4747 4647
rect 4813 4613 4827 4627
rect 4773 4433 4787 4447
rect 4793 4413 4807 4427
rect 4733 4313 4747 4327
rect 4673 4173 4687 4187
rect 4633 4153 4647 4167
rect 4653 4153 4667 4167
rect 4593 3993 4607 4007
rect 4653 3993 4667 4007
rect 4533 3833 4547 3847
rect 4493 3753 4507 3767
rect 4393 3693 4407 3707
rect 4433 3693 4447 3707
rect 4453 3693 4467 3707
rect 4513 3713 4527 3727
rect 4373 3673 4387 3687
rect 4413 3673 4427 3687
rect 4473 3673 4487 3687
rect 4553 3673 4567 3687
rect 4673 3953 4687 3967
rect 4753 4173 4767 4187
rect 4713 4133 4727 4147
rect 4713 4013 4727 4027
rect 4713 3913 4727 3927
rect 4753 4013 4767 4027
rect 4833 4573 4847 4587
rect 4873 4633 4887 4647
rect 4913 4953 4927 4967
rect 4953 4973 4967 4987
rect 5093 5593 5107 5607
rect 5033 5513 5047 5527
rect 5093 5473 5107 5487
rect 5133 5473 5147 5487
rect 5133 5433 5147 5447
rect 5173 5673 5187 5687
rect 5233 5773 5247 5787
rect 5393 5773 5407 5787
rect 5193 5633 5207 5647
rect 5213 5613 5227 5627
rect 5173 5433 5187 5447
rect 5113 5353 5127 5367
rect 5073 5173 5087 5187
rect 5073 5113 5087 5127
rect 5053 5073 5067 5087
rect 5013 4993 5027 5007
rect 5013 4953 5027 4967
rect 5053 4953 5067 4967
rect 4973 4913 4987 4927
rect 5053 4873 5067 4887
rect 5153 5393 5167 5407
rect 5133 5093 5147 5107
rect 5133 4973 5147 4987
rect 5093 4953 5107 4967
rect 5173 5333 5187 5347
rect 5153 4953 5167 4967
rect 5153 4933 5167 4947
rect 5133 4913 5147 4927
rect 5073 4793 5087 4807
rect 4953 4713 4967 4727
rect 5053 4713 5067 4727
rect 5033 4673 5047 4687
rect 5073 4673 5087 4687
rect 4953 4653 4967 4667
rect 5013 4653 5027 4667
rect 4933 4613 4947 4627
rect 4893 4593 4907 4607
rect 4853 4493 4867 4507
rect 4873 4473 4887 4487
rect 4933 4473 4947 4487
rect 4813 4133 4827 4147
rect 4753 3953 4767 3967
rect 4773 3953 4787 3967
rect 4813 3953 4827 3967
rect 4733 3893 4747 3907
rect 4813 3853 4827 3867
rect 4593 3793 4607 3807
rect 4693 3813 4707 3827
rect 4673 3793 4687 3807
rect 4633 3713 4647 3727
rect 4653 3693 4667 3707
rect 4753 3773 4767 3787
rect 4793 3713 4807 3727
rect 4733 3693 4747 3707
rect 4353 3573 4367 3587
rect 4313 3513 4327 3527
rect 4273 3493 4287 3507
rect 4313 3493 4327 3507
rect 4233 3253 4247 3267
rect 4293 3253 4307 3267
rect 4193 3233 4207 3247
rect 4233 3233 4247 3247
rect 4173 3113 4187 3127
rect 4213 3193 4227 3207
rect 4573 3533 4587 3547
rect 4393 3493 4407 3507
rect 4433 3493 4447 3507
rect 4473 3493 4487 3507
rect 4493 3493 4507 3507
rect 4533 3493 4547 3507
rect 4373 3453 4387 3467
rect 4353 3413 4367 3427
rect 4453 3473 4467 3487
rect 4373 3233 4387 3247
rect 4413 3233 4427 3247
rect 4253 3173 4267 3187
rect 4333 3173 4347 3187
rect 4273 3133 4287 3147
rect 4253 3113 4267 3127
rect 4193 3093 4207 3107
rect 4213 3073 4227 3087
rect 4153 3033 4167 3047
rect 4213 3033 4227 3047
rect 4193 2993 4207 3007
rect 4233 2973 4247 2987
rect 4253 2813 4267 2827
rect 4153 2773 4167 2787
rect 4173 2773 4187 2787
rect 4213 2773 4227 2787
rect 4253 2773 4267 2787
rect 4193 2753 4207 2767
rect 4233 2753 4247 2767
rect 4253 2733 4267 2747
rect 4233 2713 4247 2727
rect 4053 2693 4067 2707
rect 4093 2693 4107 2707
rect 4133 2693 4147 2707
rect 4073 2533 4087 2547
rect 4033 2513 4047 2527
rect 4013 2473 4027 2487
rect 4253 2533 4267 2547
rect 4093 2393 4107 2407
rect 3993 2353 4007 2367
rect 3953 2153 3967 2167
rect 3973 2073 3987 2087
rect 4253 2333 4267 2347
rect 4373 3173 4387 3187
rect 4333 3093 4347 3107
rect 4353 3093 4367 3107
rect 4293 3053 4307 3067
rect 4293 2793 4307 2807
rect 4353 3053 4367 3067
rect 4413 3173 4427 3187
rect 4413 3153 4427 3167
rect 4393 3053 4407 3067
rect 4453 3233 4467 3247
rect 4513 3473 4527 3487
rect 4513 3453 4527 3467
rect 4453 3113 4467 3127
rect 4433 3093 4447 3107
rect 4433 3033 4447 3047
rect 4473 3033 4487 3047
rect 4353 2993 4367 3007
rect 4373 2993 4387 3007
rect 4313 2433 4327 2447
rect 4413 2933 4427 2947
rect 4413 2753 4427 2767
rect 4393 2713 4407 2727
rect 4013 2293 4027 2307
rect 4173 2253 4187 2267
rect 4153 2233 4167 2247
rect 4033 2153 4047 2167
rect 4013 2073 4027 2087
rect 3933 2033 3947 2047
rect 3913 1993 3927 2007
rect 3933 1993 3947 2007
rect 3993 2053 4007 2067
rect 4013 2053 4027 2067
rect 4053 2113 4067 2127
rect 4073 2093 4087 2107
rect 4053 2033 4067 2047
rect 4033 1873 4047 1887
rect 4053 1873 4067 1887
rect 4013 1833 4027 1847
rect 3953 1813 3967 1827
rect 3953 1793 3967 1807
rect 3993 1793 4007 1807
rect 3933 1773 3947 1787
rect 3953 1733 3967 1747
rect 3893 1693 3907 1707
rect 3913 1653 3927 1667
rect 3873 1593 3887 1607
rect 3893 1573 3907 1587
rect 3853 1513 3867 1527
rect 3793 1413 3807 1427
rect 3833 1413 3847 1427
rect 3653 1393 3667 1407
rect 3693 1393 3707 1407
rect 3733 1373 3747 1387
rect 3773 1373 3787 1387
rect 3693 1313 3707 1327
rect 3673 1273 3687 1287
rect 3753 1293 3767 1307
rect 3733 1273 3747 1287
rect 3713 1253 3727 1267
rect 3793 1253 3807 1267
rect 3633 1193 3647 1207
rect 3593 1173 3607 1187
rect 3553 1153 3567 1167
rect 3533 1133 3547 1147
rect 3513 993 3527 1007
rect 3493 973 3507 987
rect 3473 853 3487 867
rect 3473 833 3487 847
rect 3453 353 3467 367
rect 3333 313 3347 327
rect 3433 293 3447 307
rect 3313 193 3327 207
rect 3033 173 3047 187
rect 3193 173 3207 187
rect 3053 133 3067 147
rect 3173 133 3187 147
rect 2993 113 3007 127
rect 3073 113 3087 127
rect 3373 193 3387 207
rect 3413 153 3427 167
rect 3213 133 3227 147
rect 3293 133 3307 147
rect 3333 133 3347 147
rect 3393 133 3407 147
rect 3433 133 3447 147
rect 3153 93 3167 107
rect 2953 13 2967 27
rect 3593 1113 3607 1127
rect 3813 1213 3827 1227
rect 3713 1193 3727 1207
rect 3773 1193 3787 1207
rect 3673 1173 3687 1187
rect 3573 1093 3587 1107
rect 3613 1093 3627 1107
rect 3653 1093 3667 1107
rect 3593 1073 3607 1087
rect 3533 913 3547 927
rect 3513 813 3527 827
rect 3533 793 3547 807
rect 3553 793 3567 807
rect 3553 673 3567 687
rect 3653 1033 3667 1047
rect 3653 913 3667 927
rect 3693 1113 3707 1127
rect 3733 1113 3747 1127
rect 3793 1173 3807 1187
rect 3993 1773 4007 1787
rect 3973 1693 3987 1707
rect 3993 1653 4007 1667
rect 3973 1613 3987 1627
rect 3953 1413 3967 1427
rect 3913 1353 3927 1367
rect 3893 1213 3907 1227
rect 3853 1173 3867 1187
rect 3853 1133 3867 1147
rect 3693 1073 3707 1087
rect 3793 1073 3807 1087
rect 3753 1033 3767 1047
rect 3693 973 3707 987
rect 3673 833 3687 847
rect 3793 933 3807 947
rect 3893 1113 3907 1127
rect 3833 1073 3847 1087
rect 3873 1073 3887 1087
rect 3713 853 3727 867
rect 3673 793 3687 807
rect 3513 633 3527 647
rect 3553 633 3567 647
rect 3493 613 3507 627
rect 3533 613 3547 627
rect 3493 433 3507 447
rect 3633 653 3647 667
rect 3593 633 3607 647
rect 3613 633 3627 647
rect 3673 633 3687 647
rect 3653 593 3667 607
rect 3493 393 3507 407
rect 3573 393 3587 407
rect 3593 393 3607 407
rect 3533 373 3547 387
rect 3693 613 3707 627
rect 3693 453 3707 467
rect 3673 373 3687 387
rect 3633 353 3647 367
rect 3813 893 3827 907
rect 3733 833 3747 847
rect 3793 833 3807 847
rect 3753 793 3767 807
rect 3793 793 3807 807
rect 3793 713 3807 727
rect 3853 933 3867 947
rect 3873 893 3887 907
rect 3913 1093 3927 1107
rect 3993 1593 4007 1607
rect 4013 1593 4027 1607
rect 4093 2073 4107 2087
rect 4133 2073 4147 2087
rect 4273 2273 4287 2287
rect 4253 2093 4267 2107
rect 4113 2033 4127 2047
rect 4093 1933 4107 1947
rect 4153 1913 4167 1927
rect 4133 1893 4147 1907
rect 4113 1833 4127 1847
rect 4133 1813 4147 1827
rect 4113 1793 4127 1807
rect 4213 2073 4227 2087
rect 4193 2053 4207 2067
rect 4173 1873 4187 1887
rect 4173 1833 4187 1847
rect 4153 1773 4167 1787
rect 4093 1693 4107 1707
rect 4073 1673 4087 1687
rect 4073 1633 4087 1647
rect 4013 1473 4027 1487
rect 4073 1353 4087 1367
rect 4133 1593 4147 1607
rect 4153 1553 4167 1567
rect 4113 1513 4127 1527
rect 4253 2053 4267 2067
rect 4273 2013 4287 2027
rect 4413 2433 4427 2447
rect 4413 2393 4427 2407
rect 4373 2313 4387 2327
rect 4353 2273 4367 2287
rect 4393 2253 4407 2267
rect 4373 2213 4387 2227
rect 4293 1973 4307 1987
rect 4293 1953 4307 1967
rect 4373 2073 4387 2087
rect 4453 2833 4467 2847
rect 4633 3673 4647 3687
rect 4753 3653 4767 3667
rect 4673 3593 4687 3607
rect 4733 3593 4747 3607
rect 4653 3553 4667 3567
rect 4613 3513 4627 3527
rect 4613 3453 4627 3467
rect 4593 3373 4607 3387
rect 4553 3273 4567 3287
rect 4573 3273 4587 3287
rect 4593 3213 4607 3227
rect 4673 3533 4687 3547
rect 4693 3533 4707 3547
rect 4573 3193 4587 3207
rect 4653 3193 4667 3207
rect 4553 3173 4567 3187
rect 4713 3273 4727 3287
rect 4773 3593 4787 3607
rect 4893 4433 4907 4447
rect 4933 4433 4947 4447
rect 4933 4393 4947 4407
rect 4913 4293 4927 4307
rect 4853 4153 4867 4167
rect 4873 4153 4887 4167
rect 4933 4093 4947 4107
rect 4913 4013 4927 4027
rect 4873 3973 4887 3987
rect 4893 3973 4907 3987
rect 4933 3953 4947 3967
rect 4913 3893 4927 3907
rect 4853 3873 4867 3887
rect 4853 3813 4867 3827
rect 4833 3453 4847 3467
rect 4813 3433 4827 3447
rect 4833 3413 4847 3427
rect 4813 3273 4827 3287
rect 4773 3213 4787 3227
rect 4793 3213 4807 3227
rect 4793 3193 4807 3207
rect 4673 3173 4687 3187
rect 4713 3093 4727 3107
rect 4713 3053 4727 3067
rect 4613 3033 4627 3047
rect 4693 3033 4707 3047
rect 4753 3033 4767 3047
rect 4773 3033 4787 3047
rect 4533 3013 4547 3027
rect 4633 3013 4647 3027
rect 4533 2713 4547 2727
rect 4553 2673 4567 2687
rect 4513 2653 4527 2667
rect 4613 2993 4627 3007
rect 4613 2813 4627 2827
rect 4593 2773 4607 2787
rect 4593 2733 4607 2747
rect 4573 2613 4587 2627
rect 4453 2493 4467 2507
rect 4453 2473 4467 2487
rect 4473 2433 4487 2447
rect 4513 2453 4527 2467
rect 4433 2313 4447 2327
rect 4473 2293 4487 2307
rect 4813 2993 4827 3007
rect 4793 2953 4807 2967
rect 4733 2933 4747 2947
rect 4693 2733 4707 2747
rect 4773 2733 4787 2747
rect 4633 2593 4647 2607
rect 4813 2673 4827 2687
rect 4833 2453 4847 2467
rect 4693 2393 4707 2407
rect 4613 2373 4627 2387
rect 4673 2353 4687 2367
rect 4553 2313 4567 2327
rect 4633 2313 4647 2327
rect 4593 2273 4607 2287
rect 4613 2253 4627 2267
rect 4593 2233 4607 2247
rect 4533 2193 4547 2207
rect 4513 2133 4527 2147
rect 4453 2093 4467 2107
rect 4513 2093 4527 2107
rect 4313 1913 4327 1927
rect 4213 1893 4227 1907
rect 4213 1853 4227 1867
rect 4273 1833 4287 1847
rect 4233 1793 4247 1807
rect 4253 1773 4267 1787
rect 4393 2053 4407 2067
rect 4433 2053 4447 2067
rect 4413 1913 4427 1927
rect 4353 1833 4367 1847
rect 4333 1753 4347 1767
rect 4333 1733 4347 1747
rect 4233 1673 4247 1687
rect 4333 1693 4347 1707
rect 4473 2073 4487 2087
rect 4573 2193 4587 2207
rect 4553 2073 4567 2087
rect 4493 2053 4507 2067
rect 4533 2053 4547 2067
rect 4453 1833 4467 1847
rect 4493 1833 4507 1847
rect 4553 1833 4567 1847
rect 4173 1373 4187 1387
rect 4133 1353 4147 1367
rect 4053 1313 4067 1327
rect 4093 1313 4107 1327
rect 4013 1273 4027 1287
rect 4013 1133 4027 1147
rect 3973 1113 3987 1127
rect 3973 1093 3987 1107
rect 3913 1013 3927 1027
rect 3833 833 3847 847
rect 3813 653 3827 667
rect 3773 633 3787 647
rect 3793 613 3807 627
rect 3733 593 3747 607
rect 3813 513 3827 527
rect 3733 393 3747 407
rect 3793 393 3807 407
rect 3713 333 3727 347
rect 3553 193 3567 207
rect 3553 173 3567 187
rect 3533 133 3547 147
rect 3673 293 3687 307
rect 3733 173 3747 187
rect 3893 853 3907 867
rect 3853 753 3867 767
rect 3913 833 3927 847
rect 3893 813 3907 827
rect 3993 893 4007 907
rect 4093 1133 4107 1147
rect 4113 1113 4127 1127
rect 4053 1053 4067 1067
rect 4153 1313 4167 1327
rect 4193 1313 4207 1327
rect 4173 1273 4187 1287
rect 4213 1233 4227 1247
rect 4213 1193 4227 1207
rect 4153 1113 4167 1127
rect 4173 1113 4187 1127
rect 4033 853 4047 867
rect 4013 833 4027 847
rect 3893 713 3907 727
rect 3873 693 3887 707
rect 3933 653 3947 667
rect 3913 633 3927 647
rect 3893 613 3907 627
rect 4093 873 4107 887
rect 4133 873 4147 887
rect 3993 793 4007 807
rect 4053 793 4067 807
rect 4073 773 4087 787
rect 4033 693 4047 707
rect 4073 633 4087 647
rect 3993 613 4007 627
rect 3913 533 3927 547
rect 3953 533 3967 547
rect 3853 413 3867 427
rect 3893 413 3907 427
rect 3833 393 3847 407
rect 3853 373 3867 387
rect 3833 333 3847 347
rect 3873 333 3887 347
rect 4053 613 4067 627
rect 4013 513 4027 527
rect 4113 853 4127 867
rect 4153 853 4167 867
rect 4213 913 4227 927
rect 4173 833 4187 847
rect 4133 793 4147 807
rect 4113 433 4127 447
rect 4193 813 4207 827
rect 4293 1653 4307 1667
rect 4253 1593 4267 1607
rect 4353 1653 4367 1667
rect 4333 1593 4347 1607
rect 4273 1573 4287 1587
rect 4273 1473 4287 1487
rect 4313 1473 4327 1487
rect 4353 1393 4367 1407
rect 4313 1313 4327 1327
rect 4293 1293 4307 1307
rect 4273 1273 4287 1287
rect 4333 1273 4347 1287
rect 4453 1793 4467 1807
rect 4433 1773 4447 1787
rect 4473 1773 4487 1787
rect 4453 1693 4467 1707
rect 4453 1613 4467 1627
rect 4473 1613 4487 1627
rect 4493 1593 4507 1607
rect 4433 1573 4447 1587
rect 4473 1473 4487 1487
rect 4493 1333 4507 1347
rect 4553 1773 4567 1787
rect 4533 1733 4547 1747
rect 4553 1713 4567 1727
rect 4553 1693 4567 1707
rect 4533 1613 4547 1627
rect 4633 2153 4647 2167
rect 4633 2053 4647 2067
rect 4613 2033 4627 2047
rect 4613 2013 4627 2027
rect 4593 1793 4607 1807
rect 4653 1993 4667 2007
rect 4733 2293 4747 2307
rect 4713 2253 4727 2267
rect 4713 2173 4727 2187
rect 4693 2093 4707 2107
rect 4673 1833 4687 1847
rect 4793 2393 4807 2407
rect 4773 2093 4787 2107
rect 4753 2053 4767 2067
rect 4733 2033 4747 2047
rect 4873 3673 4887 3687
rect 4893 3573 4907 3587
rect 4913 3493 4927 3507
rect 4893 3473 4907 3487
rect 4933 3353 4947 3367
rect 5053 4633 5067 4647
rect 5013 4613 5027 4627
rect 4973 4473 4987 4487
rect 5073 4593 5087 4607
rect 5113 4693 5127 4707
rect 5113 4653 5127 4667
rect 5313 5653 5327 5667
rect 5293 5613 5307 5627
rect 5313 5593 5327 5607
rect 5233 5553 5247 5567
rect 5253 5513 5267 5527
rect 5233 5473 5247 5487
rect 5293 5433 5307 5447
rect 5273 5413 5287 5427
rect 5233 5393 5247 5407
rect 5233 5373 5247 5387
rect 5213 5313 5227 5327
rect 5213 5153 5227 5167
rect 5293 5193 5307 5207
rect 5193 5113 5207 5127
rect 5193 5093 5207 5107
rect 5233 5073 5247 5087
rect 5213 4853 5227 4867
rect 5173 4833 5187 4847
rect 5233 4833 5247 4847
rect 5213 4733 5227 4747
rect 5193 4713 5207 4727
rect 5153 4693 5167 4707
rect 5173 4673 5187 4687
rect 5193 4633 5207 4647
rect 5133 4533 5147 4547
rect 5093 4513 5107 4527
rect 5153 4513 5167 4527
rect 5013 4433 5027 4447
rect 4993 4413 5007 4427
rect 4993 4193 5007 4207
rect 4993 4133 5007 4147
rect 4973 3993 4987 4007
rect 4973 3493 4987 3507
rect 5053 4413 5067 4427
rect 5053 4153 5067 4167
rect 5013 3973 5027 3987
rect 5013 3753 5027 3767
rect 5053 3733 5067 3747
rect 5033 3713 5047 3727
rect 5133 4453 5147 4467
rect 5133 4393 5147 4407
rect 5173 4493 5187 4507
rect 5213 4513 5227 4527
rect 5213 4473 5227 4487
rect 5293 4993 5307 5007
rect 5273 4733 5287 4747
rect 5373 5613 5387 5627
rect 5353 5593 5367 5607
rect 5353 5193 5367 5207
rect 5353 5153 5367 5167
rect 5333 5093 5347 5107
rect 5333 5053 5347 5067
rect 5253 4713 5267 4727
rect 5273 4713 5287 4727
rect 5313 4693 5327 4707
rect 5333 4693 5347 4707
rect 5313 4653 5327 4667
rect 5373 4773 5387 4787
rect 5373 4653 5387 4667
rect 5333 4633 5347 4647
rect 5353 4633 5367 4647
rect 5453 5693 5467 5707
rect 5593 5773 5607 5787
rect 5553 5753 5567 5767
rect 5633 5673 5647 5687
rect 5573 5653 5587 5667
rect 5633 5653 5647 5667
rect 5513 5613 5527 5627
rect 5433 5593 5447 5607
rect 5513 5593 5527 5607
rect 5413 5573 5427 5587
rect 5433 5473 5447 5487
rect 5473 5433 5487 5447
rect 5493 5433 5507 5447
rect 5453 5353 5467 5367
rect 5453 5153 5467 5167
rect 5473 5133 5487 5147
rect 5453 5113 5467 5127
rect 5473 5113 5487 5127
rect 5453 5053 5467 5067
rect 5453 4973 5467 4987
rect 5433 4913 5447 4927
rect 5433 4893 5447 4907
rect 5453 4773 5467 4787
rect 5413 4693 5427 4707
rect 5453 4693 5467 4707
rect 5433 4673 5447 4687
rect 5433 4653 5447 4667
rect 5313 4593 5327 4607
rect 5393 4593 5407 4607
rect 5153 4213 5167 4227
rect 5093 4193 5107 4207
rect 5193 4413 5207 4427
rect 5193 4393 5207 4407
rect 5193 4193 5207 4207
rect 5173 4153 5187 4167
rect 5113 4113 5127 4127
rect 5113 4093 5127 4107
rect 5153 4013 5167 4027
rect 5293 4553 5307 4567
rect 5293 4533 5307 4547
rect 5293 4513 5307 4527
rect 5293 4233 5307 4247
rect 5273 4213 5287 4227
rect 5253 4193 5267 4207
rect 5293 4193 5307 4207
rect 5353 4513 5367 4527
rect 5333 4493 5347 4507
rect 5213 4133 5227 4147
rect 5233 4093 5247 4107
rect 5273 4073 5287 4087
rect 5233 4053 5247 4067
rect 5293 4053 5307 4067
rect 5313 4053 5327 4067
rect 5193 4033 5207 4047
rect 5113 3973 5127 3987
rect 5133 3953 5147 3967
rect 5093 3933 5107 3947
rect 5073 3673 5087 3687
rect 5033 3553 5047 3567
rect 5073 3513 5087 3527
rect 5013 3493 5027 3507
rect 4993 3473 5007 3487
rect 5053 3453 5067 3467
rect 4973 3353 4987 3367
rect 4893 3273 4907 3287
rect 4953 3273 4967 3287
rect 4933 3253 4947 3267
rect 4913 3233 4927 3247
rect 5053 3233 5067 3247
rect 4873 3213 4887 3227
rect 4933 3213 4947 3227
rect 4953 3213 4967 3227
rect 4973 3213 4987 3227
rect 4893 3013 4907 3027
rect 4873 2993 4887 3007
rect 4913 2973 4927 2987
rect 4913 2713 4927 2727
rect 4853 2353 4867 2367
rect 4853 2333 4867 2347
rect 4813 2273 4827 2287
rect 4833 2233 4847 2247
rect 4813 2093 4827 2107
rect 4713 2013 4727 2027
rect 4713 1873 4727 1887
rect 4713 1853 4727 1867
rect 4633 1773 4647 1787
rect 4613 1693 4627 1707
rect 4613 1613 4627 1627
rect 4573 1593 4587 1607
rect 4653 1593 4667 1607
rect 4553 1573 4567 1587
rect 4533 1373 4547 1387
rect 4633 1573 4647 1587
rect 4593 1533 4607 1547
rect 4753 2013 4767 2027
rect 4813 2013 4827 2027
rect 4733 1813 4747 1827
rect 4693 1753 4707 1767
rect 4653 1333 4667 1347
rect 4673 1333 4687 1347
rect 4553 1313 4567 1327
rect 4593 1313 4607 1327
rect 4633 1313 4647 1327
rect 4453 1293 4467 1307
rect 4433 1253 4447 1267
rect 4473 1253 4487 1267
rect 4433 1213 4447 1227
rect 4413 1193 4427 1207
rect 4253 1173 4267 1187
rect 4373 1173 4387 1187
rect 4233 893 4247 907
rect 4353 1153 4367 1167
rect 4393 1153 4407 1167
rect 4353 1133 4367 1147
rect 4313 1113 4327 1127
rect 4333 1093 4347 1107
rect 4453 1133 4467 1147
rect 4453 1093 4467 1107
rect 4513 1293 4527 1307
rect 4573 1293 4587 1307
rect 4573 1273 4587 1287
rect 4493 1153 4507 1167
rect 4533 1153 4547 1167
rect 4493 1113 4507 1127
rect 4513 1093 4527 1107
rect 4413 1073 4427 1087
rect 4793 1873 4807 1887
rect 4793 1793 4807 1807
rect 4753 1753 4767 1767
rect 4813 1773 4827 1787
rect 4773 1733 4787 1747
rect 4773 1673 4787 1687
rect 4813 1693 4827 1707
rect 4793 1633 4807 1647
rect 4793 1613 4807 1627
rect 4753 1593 4767 1607
rect 4773 1593 4787 1607
rect 4733 1553 4747 1567
rect 4773 1513 4787 1527
rect 4733 1493 4747 1507
rect 4753 1413 4767 1427
rect 4713 1333 4727 1347
rect 4733 1313 4747 1327
rect 4893 2313 4907 2327
rect 4893 2293 4907 2307
rect 4873 2253 4887 2267
rect 5073 3213 5087 3227
rect 5133 3913 5147 3927
rect 5133 3793 5147 3807
rect 5153 3753 5167 3767
rect 5153 3693 5167 3707
rect 5113 3673 5127 3687
rect 5213 3873 5227 3887
rect 5173 3573 5187 3587
rect 5133 3513 5147 3527
rect 5153 3513 5167 3527
rect 5173 3493 5187 3507
rect 5153 3473 5167 3487
rect 5113 3453 5127 3467
rect 5133 3453 5147 3467
rect 4993 3033 5007 3047
rect 5033 3033 5047 3047
rect 5013 2993 5027 3007
rect 4973 2973 4987 2987
rect 4953 2773 4967 2787
rect 4973 2753 4987 2767
rect 5013 2753 5027 2767
rect 5053 2753 5067 2767
rect 4953 2733 4967 2747
rect 4993 2733 5007 2747
rect 4933 2293 4947 2307
rect 4913 2273 4927 2287
rect 4993 2713 5007 2727
rect 5053 2673 5067 2687
rect 4973 2433 4987 2447
rect 5193 3453 5207 3467
rect 5153 3253 5167 3267
rect 5153 3233 5167 3247
rect 5113 3053 5127 3067
rect 5173 3053 5187 3067
rect 5133 3033 5147 3047
rect 5193 3013 5207 3027
rect 5113 2993 5127 3007
rect 5173 2973 5187 2987
rect 5133 2773 5147 2787
rect 5173 2773 5187 2787
rect 5153 2753 5167 2767
rect 5173 2733 5187 2747
rect 5133 2433 5147 2447
rect 5073 2333 5087 2347
rect 5053 2273 5067 2287
rect 5093 2273 5107 2287
rect 5133 2273 5147 2287
rect 4973 2253 4987 2267
rect 4933 2233 4947 2247
rect 4893 2173 4907 2187
rect 4953 2133 4967 2147
rect 4873 2073 4887 2087
rect 4913 2073 4927 2087
rect 4853 2033 4867 2047
rect 4853 1833 4867 1847
rect 4833 1653 4847 1667
rect 4893 2053 4907 2067
rect 4933 2053 4947 2067
rect 5033 2193 5047 2207
rect 5033 2173 5047 2187
rect 4993 2153 5007 2167
rect 4893 1853 4907 1867
rect 4933 1813 4947 1827
rect 4913 1793 4927 1807
rect 4913 1733 4927 1747
rect 4853 1613 4867 1627
rect 4873 1613 4887 1627
rect 4893 1593 4907 1607
rect 4833 1553 4847 1567
rect 4853 1553 4867 1567
rect 4813 1533 4827 1547
rect 4933 1613 4947 1627
rect 4873 1513 4887 1527
rect 4813 1393 4827 1407
rect 4853 1393 4867 1407
rect 4853 1373 4867 1387
rect 4893 1313 4907 1327
rect 4693 1273 4707 1287
rect 4793 1273 4807 1287
rect 4793 1253 4807 1267
rect 4653 1173 4667 1187
rect 4693 1173 4707 1187
rect 4613 1133 4627 1147
rect 4653 1093 4667 1107
rect 4673 1093 4687 1107
rect 4593 873 4607 887
rect 4713 1153 4727 1167
rect 4713 1133 4727 1147
rect 4733 1133 4747 1147
rect 4773 1113 4787 1127
rect 4713 1093 4727 1107
rect 4893 1273 4907 1287
rect 4873 1193 4887 1207
rect 4813 1113 4827 1127
rect 4693 1073 4707 1087
rect 4753 1073 4767 1087
rect 4773 1073 4787 1087
rect 4813 1073 4827 1087
rect 4853 1073 4867 1087
rect 4613 853 4627 867
rect 4313 833 4327 847
rect 4393 833 4407 847
rect 4433 833 4447 847
rect 4513 833 4527 847
rect 4253 813 4267 827
rect 4293 793 4307 807
rect 4333 753 4347 767
rect 4353 673 4367 687
rect 4173 653 4187 667
rect 4213 653 4227 667
rect 4373 653 4387 667
rect 4213 633 4227 647
rect 4193 613 4207 627
rect 4233 613 4247 627
rect 4333 613 4347 627
rect 4213 593 4227 607
rect 4213 553 4227 567
rect 4193 433 4207 447
rect 3933 373 3947 387
rect 3913 353 3927 367
rect 3953 353 3967 367
rect 4013 353 4027 367
rect 3993 333 4007 347
rect 4013 253 4027 267
rect 3673 113 3687 127
rect 3633 93 3647 107
rect 3853 153 3867 167
rect 4053 193 4067 207
rect 4013 133 4027 147
rect 3993 113 4007 127
rect 4153 393 4167 407
rect 4173 393 4187 407
rect 4093 373 4107 387
rect 4133 373 4147 387
rect 4113 353 4127 367
rect 4193 353 4207 367
rect 4213 333 4227 347
rect 4173 313 4187 327
rect 4273 353 4287 367
rect 4253 333 4267 347
rect 4233 293 4247 307
rect 4413 793 4427 807
rect 4573 833 4587 847
rect 4533 813 4547 827
rect 4553 793 4567 807
rect 4513 733 4527 747
rect 4433 693 4447 707
rect 4593 673 4607 687
rect 4473 653 4487 667
rect 4793 873 4807 887
rect 4873 873 4887 887
rect 4653 853 4667 867
rect 4773 853 4787 867
rect 4693 833 4707 847
rect 4733 833 4747 847
rect 4673 733 4687 747
rect 4733 793 4747 807
rect 4773 793 4787 807
rect 4773 753 4787 767
rect 4713 673 4727 687
rect 4653 653 4667 667
rect 4633 633 4647 647
rect 4813 793 4827 807
rect 4853 773 4867 787
rect 4853 693 4867 707
rect 4833 673 4847 687
rect 4793 653 4807 667
rect 4713 633 4727 647
rect 4733 633 4747 647
rect 4773 633 4787 647
rect 4393 613 4407 627
rect 4453 613 4467 627
rect 4573 613 4587 627
rect 4613 613 4627 627
rect 4653 613 4667 627
rect 4913 1133 4927 1147
rect 4913 1073 4927 1087
rect 4893 853 4907 867
rect 4893 833 4907 847
rect 4973 1833 4987 1847
rect 5053 2133 5067 2147
rect 5013 2113 5027 2127
rect 5013 2073 5027 2087
rect 5113 2253 5127 2267
rect 5133 2233 5147 2247
rect 5073 2113 5087 2127
rect 5093 2113 5107 2127
rect 5113 2113 5127 2127
rect 5073 2033 5087 2047
rect 5013 2013 5027 2027
rect 5073 1913 5087 1927
rect 5033 1833 5047 1847
rect 4993 1813 5007 1827
rect 4973 1793 4987 1807
rect 5013 1773 5027 1787
rect 5053 1773 5067 1787
rect 4993 1753 5007 1767
rect 5053 1753 5067 1767
rect 5093 1753 5107 1767
rect 5013 1673 5027 1687
rect 5013 1613 5027 1627
rect 5033 1533 5047 1547
rect 4993 1513 5007 1527
rect 5033 1453 5047 1467
rect 5013 1293 5027 1307
rect 5013 1273 5027 1287
rect 4993 1233 5007 1247
rect 4973 1133 4987 1147
rect 4993 1133 5007 1147
rect 4953 1073 4967 1087
rect 5013 1053 5027 1067
rect 5013 953 5027 967
rect 4933 873 4947 887
rect 4933 833 4947 847
rect 4973 833 4987 847
rect 4953 813 4967 827
rect 5073 1653 5087 1667
rect 5153 2113 5167 2127
rect 5253 4033 5267 4047
rect 5293 3993 5307 4007
rect 5393 4473 5407 4487
rect 5353 4433 5367 4447
rect 5373 4413 5387 4427
rect 5413 4413 5427 4427
rect 5393 4193 5407 4207
rect 5373 4153 5387 4167
rect 5393 4153 5407 4167
rect 5373 4133 5387 4147
rect 5353 4113 5367 4127
rect 5333 3993 5347 4007
rect 5253 3793 5267 3807
rect 5233 3733 5247 3747
rect 5233 3713 5247 3727
rect 5293 3713 5307 3727
rect 5453 4633 5467 4647
rect 5433 4153 5447 4167
rect 5513 5113 5527 5127
rect 5493 5093 5507 5107
rect 5573 5613 5587 5627
rect 5673 5633 5687 5647
rect 5653 5573 5667 5587
rect 5673 5533 5687 5547
rect 5613 5413 5627 5427
rect 5633 5393 5647 5407
rect 5573 5353 5587 5367
rect 5593 5353 5607 5367
rect 5633 5353 5647 5367
rect 5593 5313 5607 5327
rect 5573 5193 5587 5207
rect 5633 5173 5647 5187
rect 5513 4933 5527 4947
rect 5573 4953 5587 4967
rect 5573 4933 5587 4947
rect 5613 4933 5627 4947
rect 5493 4873 5507 4887
rect 5633 4913 5647 4927
rect 5573 4733 5587 4747
rect 5613 4793 5627 4807
rect 5613 4733 5627 4747
rect 5673 5393 5687 5407
rect 5713 5633 5727 5647
rect 5793 5693 5807 5707
rect 5733 5533 5747 5547
rect 5733 5433 5747 5447
rect 5673 5193 5687 5207
rect 5753 5373 5767 5387
rect 5713 5193 5727 5207
rect 5733 5193 5747 5207
rect 5713 5153 5727 5167
rect 5693 5133 5707 5147
rect 5713 5133 5727 5147
rect 5753 5133 5767 5147
rect 5673 4913 5687 4927
rect 5553 4673 5567 4687
rect 5573 4653 5587 4667
rect 5593 4653 5607 4667
rect 5513 4613 5527 4627
rect 5493 4513 5507 4527
rect 5493 4493 5507 4507
rect 5473 4433 5487 4447
rect 5593 4513 5607 4527
rect 5573 4413 5587 4427
rect 5533 4393 5547 4407
rect 5553 4293 5567 4307
rect 5493 4193 5507 4207
rect 5473 4173 5487 4187
rect 5473 4113 5487 4127
rect 5453 4073 5467 4087
rect 5413 4033 5427 4047
rect 5413 4013 5427 4027
rect 5413 3973 5427 3987
rect 5393 3873 5407 3887
rect 5433 3813 5447 3827
rect 5353 3613 5367 3627
rect 5233 3573 5247 3587
rect 5313 3553 5327 3567
rect 5293 3513 5307 3527
rect 5333 3533 5347 3547
rect 5373 3533 5387 3547
rect 5253 3273 5267 3287
rect 5293 3253 5307 3267
rect 5273 3193 5287 3207
rect 5233 3133 5247 3147
rect 5253 3033 5267 3047
rect 5373 3473 5387 3487
rect 5373 3233 5387 3247
rect 5353 3053 5367 3067
rect 5213 2693 5227 2707
rect 5193 2673 5207 2687
rect 5233 2533 5247 2547
rect 5193 2473 5207 2487
rect 5313 2753 5327 2767
rect 5313 2733 5327 2747
rect 5353 2733 5367 2747
rect 5273 2353 5287 2367
rect 5353 2693 5367 2707
rect 5313 2333 5327 2347
rect 5233 2293 5247 2307
rect 5273 2293 5287 2307
rect 5213 2253 5227 2267
rect 5213 2193 5227 2207
rect 5153 2093 5167 2107
rect 5173 2093 5187 2107
rect 5193 2093 5207 2107
rect 5153 2053 5167 2067
rect 5173 2053 5187 2067
rect 5133 1793 5147 1807
rect 5133 1773 5147 1787
rect 5073 1553 5087 1567
rect 5073 1453 5087 1467
rect 5113 1633 5127 1647
rect 5113 1513 5127 1527
rect 5093 1413 5107 1427
rect 5193 2033 5207 2047
rect 5173 1793 5187 1807
rect 5173 1713 5187 1727
rect 5193 1673 5207 1687
rect 5193 1653 5207 1667
rect 5233 2113 5247 2127
rect 5273 2093 5287 2107
rect 5253 2073 5267 2087
rect 5313 2053 5327 2067
rect 5233 2013 5247 2027
rect 5253 1913 5267 1927
rect 5293 1893 5307 1907
rect 5253 1853 5267 1867
rect 5233 1733 5247 1747
rect 5233 1713 5247 1727
rect 5173 1553 5187 1567
rect 5193 1533 5207 1547
rect 5133 1373 5147 1387
rect 5133 1353 5147 1367
rect 5093 1333 5107 1347
rect 5113 1313 5127 1327
rect 5133 1173 5147 1187
rect 5053 953 5067 967
rect 5033 893 5047 907
rect 5133 893 5147 907
rect 5073 833 5087 847
rect 5033 813 5047 827
rect 5073 793 5087 807
rect 5113 793 5127 807
rect 4913 773 4927 787
rect 5113 773 5127 787
rect 4993 673 5007 687
rect 4873 653 4887 667
rect 4913 653 4927 667
rect 4953 653 4967 667
rect 5093 653 5107 667
rect 4853 633 4867 647
rect 4893 633 4907 647
rect 4753 613 4767 627
rect 4793 613 4807 627
rect 4833 613 4847 627
rect 4873 613 4887 627
rect 4813 593 4827 607
rect 4793 493 4807 507
rect 4493 453 4507 467
rect 4533 453 4547 467
rect 4513 393 4527 407
rect 4413 373 4427 387
rect 4373 353 4387 367
rect 4313 313 4327 327
rect 4173 273 4187 287
rect 4133 193 4147 207
rect 4073 153 4087 167
rect 4093 153 4107 167
rect 4113 153 4127 167
rect 4093 113 4107 127
rect 4413 293 4427 307
rect 4333 193 4347 207
rect 4293 153 4307 167
rect 4513 373 4527 387
rect 4493 353 4507 367
rect 4533 353 4547 367
rect 4573 353 4587 367
rect 4633 353 4647 367
rect 4673 353 4687 367
rect 4733 353 4747 367
rect 4593 333 4607 347
rect 4613 313 4627 327
rect 4753 313 4767 327
rect 4573 273 4587 287
rect 4453 253 4467 267
rect 4633 233 4647 247
rect 4593 213 4607 227
rect 4453 133 4467 147
rect 4393 113 4407 127
rect 4553 133 4567 147
rect 4613 133 4627 147
rect 4513 113 4527 127
rect 4573 113 4587 127
rect 4693 213 4707 227
rect 4753 173 4767 187
rect 4713 153 4727 167
rect 4813 373 4827 387
rect 5173 1433 5187 1447
rect 5153 673 5167 687
rect 5133 653 5147 667
rect 5153 653 5167 667
rect 5133 633 5147 647
rect 5093 473 5107 487
rect 5153 433 5167 447
rect 5133 413 5147 427
rect 5073 393 5087 407
rect 5013 373 5027 387
rect 4953 353 4967 367
rect 4813 313 4827 327
rect 4893 333 4907 347
rect 4973 313 4987 327
rect 4853 233 4867 247
rect 4953 213 4967 227
rect 4873 153 4887 167
rect 4833 133 4847 147
rect 5033 333 5047 347
rect 4993 193 5007 207
rect 5213 1513 5227 1527
rect 5373 2533 5387 2547
rect 5373 2313 5387 2327
rect 5353 2193 5367 2207
rect 5433 3713 5447 3727
rect 5453 3613 5467 3627
rect 5433 3433 5447 3447
rect 5433 3373 5447 3387
rect 5493 4073 5507 4087
rect 5573 4173 5587 4187
rect 5533 4153 5547 4167
rect 5513 4053 5527 4067
rect 5513 4033 5527 4047
rect 5513 3993 5527 4007
rect 5493 3973 5507 3987
rect 5493 3733 5507 3747
rect 5513 3693 5527 3707
rect 5553 3993 5567 4007
rect 5553 3653 5567 3667
rect 5613 4293 5627 4307
rect 5613 3773 5627 3787
rect 5613 3733 5627 3747
rect 5533 3513 5547 3527
rect 5573 3513 5587 3527
rect 5593 3513 5607 3527
rect 5513 3493 5527 3507
rect 5553 3493 5567 3507
rect 5493 3473 5507 3487
rect 5473 3373 5487 3387
rect 5533 3473 5547 3487
rect 5593 3453 5607 3467
rect 5573 3433 5587 3447
rect 5513 3273 5527 3287
rect 5553 3273 5567 3287
rect 5493 3233 5507 3247
rect 5473 3213 5487 3227
rect 5533 3053 5547 3067
rect 5513 3033 5527 3047
rect 5453 2913 5467 2927
rect 5493 2913 5507 2927
rect 5433 2833 5447 2847
rect 5433 2673 5447 2687
rect 5493 2833 5507 2847
rect 5473 2733 5487 2747
rect 5533 2733 5547 2747
rect 5453 2533 5467 2547
rect 5413 2413 5427 2427
rect 5413 2373 5427 2387
rect 5453 2293 5467 2307
rect 5393 2253 5407 2267
rect 5393 2233 5407 2247
rect 5373 2093 5387 2107
rect 5353 2073 5367 2087
rect 5453 2253 5467 2267
rect 5433 2113 5447 2127
rect 5433 2093 5447 2107
rect 5333 1853 5347 1867
rect 5353 1853 5367 1867
rect 5333 1833 5347 1847
rect 5293 1793 5307 1807
rect 5273 1773 5287 1787
rect 5313 1753 5327 1767
rect 5413 2013 5427 2027
rect 5393 1853 5407 1867
rect 5433 1833 5447 1847
rect 5373 1773 5387 1787
rect 5413 1773 5427 1787
rect 5353 1753 5367 1767
rect 5413 1753 5427 1767
rect 5373 1713 5387 1727
rect 5393 1713 5407 1727
rect 5273 1673 5287 1687
rect 5333 1673 5347 1687
rect 5253 1653 5267 1667
rect 5293 1653 5307 1667
rect 5273 1593 5287 1607
rect 5373 1633 5387 1647
rect 5333 1593 5347 1607
rect 5253 1533 5267 1547
rect 5233 1433 5247 1447
rect 5233 1413 5247 1427
rect 5213 1373 5227 1387
rect 5253 1353 5267 1367
rect 5313 1573 5327 1587
rect 5353 1573 5367 1587
rect 5333 1553 5347 1567
rect 5313 1513 5327 1527
rect 5273 1333 5287 1347
rect 5253 1313 5267 1327
rect 5213 1273 5227 1287
rect 5393 1533 5407 1547
rect 5433 1733 5447 1747
rect 5533 2693 5547 2707
rect 5493 2533 5507 2547
rect 5493 2373 5507 2387
rect 5573 2913 5587 2927
rect 5753 5093 5767 5107
rect 5753 4973 5767 4987
rect 5733 4913 5747 4927
rect 5713 4893 5727 4907
rect 5773 4893 5787 4907
rect 5773 4793 5787 4807
rect 5673 4713 5687 4727
rect 5693 4713 5707 4727
rect 5753 4713 5767 4727
rect 5693 4653 5707 4667
rect 5733 4653 5747 4667
rect 5773 4653 5787 4667
rect 5713 4613 5727 4627
rect 5673 4473 5687 4487
rect 5673 4433 5687 4447
rect 5673 4213 5687 4227
rect 5673 4193 5687 4207
rect 5653 4173 5667 4187
rect 5653 4153 5667 4167
rect 5733 4413 5747 4427
rect 5773 4173 5787 4187
rect 5713 4133 5727 4147
rect 5773 4133 5787 4147
rect 5693 4033 5707 4047
rect 5653 3933 5667 3947
rect 5733 3993 5747 4007
rect 5753 3973 5767 3987
rect 5713 3953 5727 3967
rect 5733 3953 5747 3967
rect 5673 3913 5687 3927
rect 5713 3913 5727 3927
rect 5693 3773 5707 3787
rect 5673 3653 5687 3667
rect 5633 3533 5647 3547
rect 5633 3513 5647 3527
rect 5653 3493 5667 3507
rect 5753 3933 5767 3947
rect 5713 3753 5727 3767
rect 5733 3753 5747 3767
rect 5753 3733 5767 3747
rect 5733 3713 5747 3727
rect 5713 3693 5727 3707
rect 5733 3493 5747 3507
rect 5713 3453 5727 3467
rect 5653 3433 5667 3447
rect 5613 3253 5627 3267
rect 5693 3253 5707 3267
rect 5633 3213 5647 3227
rect 5673 3033 5687 3047
rect 5613 3013 5627 3027
rect 5633 2753 5647 2767
rect 5733 2913 5747 2927
rect 5613 2713 5627 2727
rect 5673 2733 5687 2747
rect 5653 2693 5667 2707
rect 5613 2673 5627 2687
rect 5593 2533 5607 2547
rect 5553 2313 5567 2327
rect 5513 2293 5527 2307
rect 5553 2273 5567 2287
rect 5573 2273 5587 2287
rect 5513 2233 5527 2247
rect 5533 2153 5547 2167
rect 5533 2133 5547 2147
rect 5473 2033 5487 2047
rect 5473 2013 5487 2027
rect 5453 1713 5467 1727
rect 5433 1693 5447 1707
rect 5513 2053 5527 2067
rect 5513 2033 5527 2047
rect 5493 1873 5507 1887
rect 5493 1793 5507 1807
rect 5473 1653 5487 1667
rect 5473 1593 5487 1607
rect 5433 1553 5447 1567
rect 5453 1553 5467 1567
rect 5493 1553 5507 1567
rect 5453 1533 5467 1547
rect 5413 1493 5427 1507
rect 5433 1473 5447 1487
rect 5333 1453 5347 1467
rect 5313 1333 5327 1347
rect 5393 1333 5407 1347
rect 5293 1253 5307 1267
rect 5353 1313 5367 1327
rect 5413 1253 5427 1267
rect 5333 1153 5347 1167
rect 5373 1153 5387 1167
rect 5233 1133 5247 1147
rect 5293 1133 5307 1147
rect 5313 1133 5327 1147
rect 5273 1113 5287 1127
rect 5233 873 5247 887
rect 5213 673 5227 687
rect 5213 513 5227 527
rect 5153 373 5167 387
rect 5173 373 5187 387
rect 5133 353 5147 367
rect 5173 353 5187 367
rect 5153 333 5167 347
rect 5193 333 5207 347
rect 5133 313 5147 327
rect 5193 233 5207 247
rect 5093 193 5107 207
rect 5033 173 5047 187
rect 5073 173 5087 187
rect 4973 153 4987 167
rect 5013 153 5027 167
rect 5113 153 5127 167
rect 4993 133 5007 147
rect 5033 133 5047 147
rect 5253 813 5267 827
rect 5253 793 5267 807
rect 5273 793 5287 807
rect 5253 733 5267 747
rect 5413 1133 5427 1147
rect 5373 1113 5387 1127
rect 5313 873 5327 887
rect 5313 833 5327 847
rect 5313 813 5327 827
rect 5293 773 5307 787
rect 5273 673 5287 687
rect 5273 633 5287 647
rect 5393 1093 5407 1107
rect 5413 893 5427 907
rect 5373 833 5387 847
rect 5413 813 5427 827
rect 5333 793 5347 807
rect 5393 793 5407 807
rect 5433 733 5447 747
rect 5333 713 5347 727
rect 5253 613 5267 627
rect 5353 693 5367 707
rect 5373 693 5387 707
rect 5433 693 5447 707
rect 5293 593 5307 607
rect 5333 593 5347 607
rect 5413 633 5427 647
rect 5393 613 5407 627
rect 5533 1793 5547 1807
rect 5633 2333 5647 2347
rect 5653 2253 5667 2267
rect 5633 2233 5647 2247
rect 5713 2533 5727 2547
rect 5713 2293 5727 2307
rect 5693 2273 5707 2287
rect 5733 2273 5747 2287
rect 5633 2053 5647 2067
rect 5533 1773 5547 1787
rect 5533 1593 5547 1607
rect 5513 1473 5527 1487
rect 5593 1753 5607 1767
rect 5573 1733 5587 1747
rect 5573 1633 5587 1647
rect 5713 2233 5727 2247
rect 5673 2193 5687 2207
rect 5733 2193 5747 2207
rect 5733 2173 5747 2187
rect 5753 2133 5767 2147
rect 5673 2093 5687 2107
rect 5733 2093 5747 2107
rect 5733 2073 5747 2087
rect 5713 2053 5727 2067
rect 5673 2033 5687 2047
rect 5693 2033 5707 2047
rect 5653 1793 5667 1807
rect 5633 1613 5647 1627
rect 5653 1593 5667 1607
rect 5573 1573 5587 1587
rect 5613 1573 5627 1587
rect 5553 1553 5567 1567
rect 5593 1553 5607 1567
rect 5613 1533 5627 1547
rect 5573 1393 5587 1407
rect 5533 1373 5547 1387
rect 5553 1353 5567 1367
rect 5493 1333 5507 1347
rect 5493 1313 5507 1327
rect 5473 1173 5487 1187
rect 5473 1133 5487 1147
rect 5493 1133 5507 1147
rect 5533 1133 5547 1147
rect 5513 1113 5527 1127
rect 5593 1333 5607 1347
rect 5593 1193 5607 1207
rect 5593 1173 5607 1187
rect 5573 1073 5587 1087
rect 5493 913 5507 927
rect 5533 913 5547 927
rect 5533 873 5547 887
rect 5493 833 5507 847
rect 5573 833 5587 847
rect 5733 2033 5747 2047
rect 5773 2033 5787 2047
rect 5713 2013 5727 2027
rect 5693 1973 5707 1987
rect 5673 1533 5687 1547
rect 5653 1393 5667 1407
rect 5653 1373 5667 1387
rect 5633 1333 5647 1347
rect 5713 1613 5727 1627
rect 5693 1353 5707 1367
rect 5633 1273 5647 1287
rect 5633 1193 5647 1207
rect 5613 1113 5627 1127
rect 5673 1173 5687 1187
rect 5673 1153 5687 1167
rect 5713 1133 5727 1147
rect 5673 1093 5687 1107
rect 5693 1093 5707 1107
rect 5713 1093 5727 1107
rect 5653 1073 5667 1087
rect 5613 893 5627 907
rect 5693 873 5707 887
rect 5613 853 5627 867
rect 5653 853 5667 867
rect 5473 813 5487 827
rect 5493 773 5507 787
rect 5473 733 5487 747
rect 5453 653 5467 667
rect 5473 613 5487 627
rect 5493 533 5507 547
rect 5393 513 5407 527
rect 5253 453 5267 467
rect 5353 453 5367 467
rect 5233 353 5247 367
rect 5213 193 5227 207
rect 5353 413 5367 427
rect 5293 393 5307 407
rect 5333 353 5347 367
rect 5373 393 5387 407
rect 5373 333 5387 347
rect 5353 233 5367 247
rect 5313 213 5327 227
rect 5333 193 5347 207
rect 5233 153 5247 167
rect 5293 153 5307 167
rect 5553 813 5567 827
rect 5593 813 5607 827
rect 5593 693 5607 707
rect 5553 673 5567 687
rect 5533 633 5547 647
rect 5593 633 5607 647
rect 5573 613 5587 627
rect 5513 493 5527 507
rect 5413 473 5427 487
rect 5593 473 5607 487
rect 5513 393 5527 407
rect 5553 393 5567 407
rect 5433 373 5447 387
rect 5413 313 5427 327
rect 5233 133 5247 147
rect 5353 133 5367 147
rect 5473 353 5487 367
rect 5693 833 5707 847
rect 5673 813 5687 827
rect 5653 733 5667 747
rect 5633 653 5647 667
rect 5613 433 5627 447
rect 5673 713 5687 727
rect 5693 633 5707 647
rect 5653 593 5667 607
rect 5753 1633 5767 1647
rect 5813 5673 5827 5687
rect 5813 3933 5827 3947
rect 5813 3813 5827 3827
rect 5813 2133 5827 2147
rect 5793 1593 5807 1607
rect 5793 1573 5807 1587
rect 5773 1513 5787 1527
rect 5773 1493 5787 1507
rect 5753 1353 5767 1367
rect 5753 1153 5767 1167
rect 5753 1093 5767 1107
rect 5773 1093 5787 1107
rect 5753 873 5767 887
rect 5633 393 5647 407
rect 5613 373 5627 387
rect 5633 353 5647 367
rect 5613 333 5627 347
rect 5493 313 5507 327
rect 5453 173 5467 187
rect 5613 173 5627 187
rect 5673 533 5687 547
rect 5673 173 5687 187
rect 5493 133 5507 147
rect 5593 133 5607 147
rect 5653 133 5667 147
rect 5733 593 5747 607
rect 5713 393 5727 407
rect 5753 393 5767 407
rect 5733 353 5747 367
rect 5793 353 5807 367
rect 5733 173 5747 187
rect 5253 113 5267 127
rect 5373 113 5387 127
rect 5433 113 5447 127
rect 5673 113 5687 127
rect 4533 93 4547 107
rect 4633 93 4647 107
<< metal3 >>
rect 5087 5776 5233 5784
rect 5407 5776 5593 5784
rect 5167 5756 5553 5764
rect 5467 5696 5793 5704
rect 4847 5676 4973 5684
rect 5147 5676 5173 5684
rect 5187 5676 5633 5684
rect 5827 5676 5864 5684
rect 467 5656 513 5664
rect 847 5656 1333 5664
rect 1507 5656 1633 5664
rect 1947 5656 2073 5664
rect 2087 5656 2113 5664
rect 2387 5656 2453 5664
rect 2627 5656 2713 5664
rect 2767 5656 2793 5664
rect 2807 5656 2873 5664
rect 2887 5656 3253 5664
rect 3267 5656 3433 5664
rect 3447 5656 3493 5664
rect 3547 5656 4093 5664
rect 4456 5656 4584 5664
rect 4456 5647 4464 5656
rect 127 5636 213 5644
rect 227 5636 244 5644
rect 147 5616 193 5624
rect 236 5624 244 5636
rect 407 5636 533 5644
rect 707 5636 733 5644
rect 907 5636 933 5644
rect 1527 5636 1673 5644
rect 1687 5636 1753 5644
rect 2047 5636 2133 5644
rect 2147 5636 2173 5644
rect 2347 5636 2413 5644
rect 2487 5636 2593 5644
rect 2647 5636 2693 5644
rect 2987 5636 3073 5644
rect 3527 5636 3653 5644
rect 3867 5636 3953 5644
rect 4507 5636 4553 5644
rect 4576 5644 4584 5656
rect 4727 5656 4733 5664
rect 4747 5656 4873 5664
rect 4907 5656 5313 5664
rect 5587 5656 5633 5664
rect 5647 5656 5864 5664
rect 4576 5636 5193 5644
rect 5687 5636 5713 5644
rect 5856 5636 5864 5656
rect 236 5616 373 5624
rect 1216 5624 1224 5633
rect 787 5616 1224 5624
rect 1267 5616 1373 5624
rect 1387 5616 1393 5624
rect 1567 5616 1733 5624
rect 1887 5616 2213 5624
rect 3116 5624 3124 5633
rect 3116 5616 3233 5624
rect 3307 5616 3373 5624
rect 3387 5616 3493 5624
rect 4287 5616 4473 5624
rect 5007 5616 5053 5624
rect 5147 5616 5213 5624
rect 5307 5616 5373 5624
rect 5527 5616 5573 5624
rect 427 5596 493 5604
rect 547 5596 913 5604
rect 1007 5596 1073 5604
rect 1287 5596 1413 5604
rect 1547 5596 1693 5604
rect 1707 5596 1773 5604
rect 1787 5596 1833 5604
rect 1867 5596 1913 5604
rect 2127 5596 2153 5604
rect 2207 5596 2733 5604
rect 3147 5596 3393 5604
rect 3687 5596 3933 5604
rect 4007 5596 4073 5604
rect 4247 5596 4573 5604
rect 4827 5596 4853 5604
rect 4947 5596 5093 5604
rect 5327 5596 5353 5604
rect 5447 5596 5513 5604
rect 727 5576 893 5584
rect 907 5576 1093 5584
rect 1127 5576 1353 5584
rect 1927 5576 2313 5584
rect 3627 5576 3773 5584
rect 3787 5576 4133 5584
rect 5427 5576 5653 5584
rect 667 5556 793 5564
rect 807 5556 813 5564
rect 1827 5556 2273 5564
rect 2287 5556 2313 5564
rect 2787 5556 2813 5564
rect 2827 5556 3973 5564
rect 4527 5556 5233 5564
rect 267 5536 653 5544
rect 667 5536 1053 5544
rect 1067 5536 1393 5544
rect 2387 5536 2773 5544
rect 2787 5536 2873 5544
rect 3007 5536 3713 5544
rect 3747 5536 3973 5544
rect 5687 5536 5733 5544
rect 3407 5516 3793 5524
rect 3967 5516 4533 5524
rect 4587 5516 4913 5524
rect 4927 5516 5033 5524
rect 5047 5516 5253 5524
rect 1387 5496 3753 5504
rect 3787 5496 3853 5504
rect 3867 5496 3953 5504
rect 3987 5496 4553 5504
rect 4567 5496 4713 5504
rect 107 5476 393 5484
rect 547 5476 573 5484
rect 587 5476 693 5484
rect 1627 5476 1633 5484
rect 1647 5476 1693 5484
rect 1987 5476 2553 5484
rect 2567 5476 2933 5484
rect 3547 5476 3913 5484
rect 4447 5476 5093 5484
rect 5107 5476 5133 5484
rect 5247 5476 5433 5484
rect 87 5456 133 5464
rect 147 5456 573 5464
rect 587 5456 773 5464
rect 1147 5456 1173 5464
rect 1747 5456 1853 5464
rect 1867 5456 2053 5464
rect 2107 5456 2233 5464
rect 2247 5456 2413 5464
rect 2507 5456 2513 5464
rect 2527 5456 2853 5464
rect 2927 5456 3013 5464
rect 3027 5456 3253 5464
rect 3567 5456 3833 5464
rect 3847 5456 4313 5464
rect 4387 5456 4493 5464
rect 4507 5456 4753 5464
rect 287 5436 524 5444
rect 96 5407 104 5433
rect 127 5416 193 5424
rect 447 5416 493 5424
rect 516 5407 524 5436
rect 627 5436 833 5444
rect 967 5436 1293 5444
rect 1367 5436 1413 5444
rect 1516 5436 1553 5444
rect 607 5416 673 5424
rect 747 5416 813 5424
rect 867 5416 913 5424
rect 927 5416 933 5424
rect 987 5416 1073 5424
rect 1167 5416 1253 5424
rect 367 5396 413 5404
rect 536 5396 553 5404
rect 67 5376 73 5384
rect 536 5384 544 5396
rect 567 5396 673 5404
rect 1187 5396 1233 5404
rect 87 5376 544 5384
rect 1167 5376 1253 5384
rect 1516 5384 1524 5436
rect 1607 5436 1633 5444
rect 1656 5427 1664 5453
rect 1687 5436 1953 5444
rect 2487 5436 2553 5444
rect 2607 5436 2673 5444
rect 3107 5436 3273 5444
rect 3287 5436 3373 5444
rect 3447 5436 3533 5444
rect 3607 5436 3733 5444
rect 3827 5436 3864 5444
rect 3856 5427 3864 5436
rect 3907 5436 4093 5444
rect 4167 5436 4593 5444
rect 5147 5436 5173 5444
rect 5307 5436 5473 5444
rect 5507 5436 5733 5444
rect 1787 5416 1813 5424
rect 2047 5416 2073 5424
rect 2647 5416 2684 5424
rect 1536 5404 1544 5413
rect 1536 5396 1793 5404
rect 1987 5396 2053 5404
rect 2107 5396 2613 5404
rect 2676 5404 2684 5416
rect 2867 5416 2893 5424
rect 3147 5416 3173 5424
rect 3347 5416 3413 5424
rect 3587 5416 3693 5424
rect 3727 5416 3733 5424
rect 3807 5416 3833 5424
rect 4127 5416 4233 5424
rect 4367 5416 4473 5424
rect 4527 5416 4633 5424
rect 5287 5416 5613 5424
rect 2676 5396 2753 5404
rect 3047 5396 3113 5404
rect 3296 5404 3304 5413
rect 3296 5396 3433 5404
rect 3447 5396 3673 5404
rect 3736 5404 3744 5413
rect 3736 5396 3873 5404
rect 3907 5396 4153 5404
rect 4267 5396 4373 5404
rect 4427 5396 4513 5404
rect 4567 5396 4733 5404
rect 5167 5396 5233 5404
rect 5647 5396 5673 5404
rect 1516 5376 1533 5384
rect 2027 5376 2093 5384
rect 2656 5384 2664 5393
rect 2567 5376 2664 5384
rect 3167 5376 3333 5384
rect 3716 5384 3724 5393
rect 3716 5376 3773 5384
rect 4007 5376 4133 5384
rect 5247 5376 5753 5384
rect 427 5356 453 5364
rect 507 5356 713 5364
rect 4067 5356 4073 5364
rect 4087 5356 4213 5364
rect 4227 5356 4473 5364
rect 4807 5356 5113 5364
rect 5127 5356 5453 5364
rect 5587 5356 5593 5364
rect 5607 5356 5633 5364
rect 407 5336 473 5344
rect 4287 5336 4833 5344
rect 4887 5336 5173 5344
rect 67 5316 93 5324
rect 5227 5316 5593 5324
rect 2187 5296 2333 5304
rect 1567 5276 1593 5284
rect 3507 5256 3973 5264
rect 3987 5256 4673 5264
rect 187 5236 233 5244
rect 167 5216 233 5224
rect 247 5216 613 5224
rect 2027 5216 2193 5224
rect 3567 5216 4413 5224
rect 547 5196 993 5204
rect 2007 5196 2033 5204
rect 2107 5196 2213 5204
rect 2227 5196 2393 5204
rect 2407 5196 2553 5204
rect 3647 5196 3973 5204
rect 3996 5196 4573 5204
rect 96 5176 153 5184
rect 96 5167 104 5176
rect 207 5176 273 5184
rect 327 5176 453 5184
rect 507 5176 613 5184
rect 807 5176 1013 5184
rect 896 5167 904 5176
rect 1067 5176 1293 5184
rect 1707 5176 1893 5184
rect 1927 5176 2053 5184
rect 2067 5176 2313 5184
rect 2367 5176 2473 5184
rect 2827 5176 3553 5184
rect 3707 5176 3773 5184
rect 3996 5184 4004 5196
rect 5307 5196 5353 5204
rect 5587 5196 5673 5204
rect 5696 5196 5713 5204
rect 3927 5176 4004 5184
rect 4056 5176 4253 5184
rect 127 5156 193 5164
rect 367 5156 433 5164
rect 487 5156 573 5164
rect 767 5156 873 5164
rect 1087 5156 1153 5164
rect 1367 5156 1413 5164
rect 1467 5156 1513 5164
rect 1667 5156 1753 5164
rect 1807 5156 1833 5164
rect 2147 5156 2193 5164
rect 2287 5156 2333 5164
rect 2347 5156 2513 5164
rect 2747 5156 2893 5164
rect 3807 5156 3893 5164
rect 4036 5164 4044 5173
rect 4056 5167 4064 5176
rect 5087 5176 5633 5184
rect 4007 5156 4044 5164
rect 4227 5156 4293 5164
rect 4307 5156 4333 5164
rect 4487 5156 4633 5164
rect 4647 5156 4693 5164
rect 4856 5156 5213 5164
rect 427 5136 513 5144
rect 747 5136 813 5144
rect 867 5136 913 5144
rect 1347 5136 1433 5144
rect 1547 5136 1673 5144
rect 1727 5136 1753 5144
rect 1767 5136 1933 5144
rect 1947 5136 2073 5144
rect 2427 5136 2453 5144
rect 2567 5136 2873 5144
rect 2896 5144 2904 5153
rect 2896 5136 2993 5144
rect 3047 5136 3113 5144
rect 3127 5136 3653 5144
rect 3296 5127 3304 5136
rect 4016 5136 4193 5144
rect 4016 5127 4024 5136
rect 4267 5136 4353 5144
rect 4387 5136 4533 5144
rect 4547 5136 4593 5144
rect 4736 5144 4744 5153
rect 4667 5136 4744 5144
rect 4856 5144 4864 5156
rect 5236 5156 5353 5164
rect 4847 5136 4864 5144
rect 5236 5144 5244 5156
rect 5367 5156 5453 5164
rect 5696 5147 5704 5196
rect 5747 5196 5764 5204
rect 5756 5164 5764 5196
rect 5727 5156 5764 5164
rect 4887 5136 5244 5144
rect 5456 5136 5473 5144
rect 5456 5127 5464 5136
rect 5727 5136 5753 5144
rect 147 5116 213 5124
rect 547 5116 593 5124
rect 787 5116 853 5124
rect 907 5116 1133 5124
rect 1147 5116 1313 5124
rect 1327 5116 1353 5124
rect 1707 5116 1773 5124
rect 1787 5116 1873 5124
rect 2387 5116 2493 5124
rect 2507 5116 2553 5124
rect 2627 5116 2673 5124
rect 2687 5116 2713 5124
rect 2927 5116 3133 5124
rect 3387 5116 3513 5124
rect 3527 5116 3553 5124
rect 4187 5116 4313 5124
rect 4327 5116 4453 5124
rect 4627 5116 4713 5124
rect 4727 5116 4753 5124
rect 5087 5116 5193 5124
rect 5487 5116 5513 5124
rect 507 5096 733 5104
rect 767 5096 1033 5104
rect 1047 5096 1133 5104
rect 1147 5096 1273 5104
rect 2127 5096 2153 5104
rect 2167 5096 3033 5104
rect 3727 5096 3913 5104
rect 3927 5096 4833 5104
rect 4947 5096 5133 5104
rect 5207 5096 5333 5104
rect 5507 5096 5753 5104
rect 1127 5076 1153 5084
rect 4007 5076 4393 5084
rect 4407 5076 4853 5084
rect 5067 5076 5233 5084
rect 2367 5056 2653 5064
rect 2667 5056 3933 5064
rect 4107 5056 4913 5064
rect 5347 5056 5453 5064
rect 1787 5036 1913 5044
rect 1927 5036 2093 5044
rect 2107 5036 2433 5044
rect 2847 5036 3833 5044
rect 4247 5036 4613 5044
rect 4627 5036 4653 5044
rect 4727 5036 4893 5044
rect 47 5016 373 5024
rect 1427 5016 2433 5024
rect 2707 5016 2993 5024
rect 3007 5016 3273 5024
rect 4147 5016 4233 5024
rect 3067 4996 3113 5004
rect 3127 4996 3153 5004
rect 3167 4996 3393 5004
rect 3427 4996 3513 5004
rect 3527 4996 3773 5004
rect 3847 4996 4893 5004
rect 5027 4996 5293 5004
rect 87 4976 373 4984
rect 387 4976 413 4984
rect 967 4976 993 4984
rect 1007 4976 1233 4984
rect 1307 4976 1333 4984
rect 1587 4976 1713 4984
rect 1727 4976 1833 4984
rect 2147 4976 2373 4984
rect 2767 4976 2773 4984
rect 2787 4976 2853 4984
rect 3247 4976 3313 4984
rect 3447 4976 3493 4984
rect 3507 4976 3533 4984
rect 3867 4976 3953 4984
rect 3967 4976 4013 4984
rect 4027 4976 4133 4984
rect 4387 4976 4453 4984
rect 4467 4976 4593 4984
rect 4967 4976 5133 4984
rect 5467 4976 5753 4984
rect 176 4956 213 4964
rect 176 4924 184 4956
rect 587 4956 633 4964
rect 707 4956 773 4964
rect 827 4956 893 4964
rect 936 4956 1084 4964
rect 207 4936 233 4944
rect 307 4936 333 4944
rect 396 4927 404 4953
rect 936 4947 944 4956
rect 567 4936 653 4944
rect 807 4936 933 4944
rect 1007 4936 1053 4944
rect 1076 4944 1084 4956
rect 1127 4956 1173 4964
rect 1887 4956 1913 4964
rect 2427 4956 2453 4964
rect 2987 4956 3133 4964
rect 1076 4936 1213 4944
rect 1227 4936 1313 4944
rect 1407 4936 1433 4944
rect 1747 4936 1773 4944
rect 1807 4936 1853 4944
rect 1907 4936 1973 4944
rect 2127 4936 2193 4944
rect 2267 4936 2393 4944
rect 2527 4936 2633 4944
rect 2887 4936 2953 4944
rect 3176 4927 3184 4973
rect 3327 4956 3373 4964
rect 4067 4956 4273 4964
rect 4287 4956 4293 4964
rect 4507 4956 4633 4964
rect 4647 4956 4733 4964
rect 4927 4956 5013 4964
rect 5067 4956 5093 4964
rect 5107 4956 5153 4964
rect 5587 4956 5744 4964
rect 3387 4936 3413 4944
rect 3447 4936 3813 4944
rect 3827 4936 4193 4944
rect 4207 4936 4384 4944
rect 4376 4927 4384 4936
rect 4427 4936 4773 4944
rect 5167 4936 5513 4944
rect 5587 4936 5613 4944
rect 5736 4927 5744 4956
rect 176 4916 213 4924
rect 267 4916 313 4924
rect 327 4916 353 4924
rect 687 4916 773 4924
rect 1467 4916 1493 4924
rect 1507 4916 1533 4924
rect 1647 4916 1813 4924
rect 1927 4916 1953 4924
rect 2167 4916 2493 4924
rect 2547 4916 2593 4924
rect 2767 4916 2873 4924
rect 3527 4916 3573 4924
rect 3756 4916 3833 4924
rect 227 4896 293 4904
rect 607 4896 633 4904
rect 1427 4896 1553 4904
rect 1687 4896 1853 4904
rect 2536 4896 3433 4904
rect 2536 4887 2544 4896
rect 3587 4896 3613 4904
rect 3756 4904 3764 4916
rect 3847 4916 4033 4924
rect 4087 4916 4113 4924
rect 4187 4916 4204 4924
rect 3627 4896 3764 4904
rect 4196 4904 4204 4916
rect 4227 4916 4353 4924
rect 4567 4916 4613 4924
rect 4987 4916 5133 4924
rect 5147 4916 5433 4924
rect 5647 4916 5673 4924
rect 4196 4896 4273 4904
rect 5447 4896 5713 4904
rect 5727 4896 5773 4904
rect 127 4876 293 4884
rect 307 4876 493 4884
rect 1107 4876 1473 4884
rect 3187 4876 3293 4884
rect 3307 4876 3713 4884
rect 4287 4876 4433 4884
rect 5067 4876 5493 4884
rect 2607 4856 3313 4864
rect 3567 4856 3673 4864
rect 3987 4856 5213 4864
rect 147 4836 193 4844
rect 207 4836 553 4844
rect 3147 4836 4613 4844
rect 5187 4836 5233 4844
rect 3707 4816 3873 4824
rect 4347 4816 4493 4824
rect 4507 4816 4593 4824
rect 1827 4796 3433 4804
rect 3807 4796 3953 4804
rect 5087 4796 5613 4804
rect 5627 4796 5773 4804
rect 47 4776 113 4784
rect 187 4776 313 4784
rect 1307 4776 2113 4784
rect 3407 4776 3913 4784
rect 5387 4776 5453 4784
rect 107 4756 153 4764
rect 167 4756 413 4764
rect 427 4756 453 4764
rect 3467 4756 3473 4764
rect 3487 4756 4153 4764
rect 1367 4736 2133 4744
rect 2427 4736 2653 4744
rect 3207 4736 3653 4744
rect 3667 4736 4693 4744
rect 5227 4736 5273 4744
rect 5587 4736 5613 4744
rect 167 4716 193 4724
rect 387 4716 1013 4724
rect 1447 4716 1873 4724
rect 2247 4716 2533 4724
rect 3147 4716 3233 4724
rect 3427 4716 3593 4724
rect 3827 4716 4273 4724
rect 4427 4716 4493 4724
rect 4967 4716 5053 4724
rect 5067 4716 5193 4724
rect 5267 4716 5273 4724
rect 5287 4716 5673 4724
rect 5707 4716 5753 4724
rect 127 4696 264 4704
rect 47 4676 233 4684
rect 256 4664 264 4696
rect 407 4696 504 4704
rect 496 4687 504 4696
rect 527 4696 613 4704
rect 1567 4696 1593 4704
rect 1647 4696 1713 4704
rect 2507 4696 2573 4704
rect 2707 4696 2753 4704
rect 2807 4696 2953 4704
rect 2967 4696 3033 4704
rect 3167 4696 3193 4704
rect 3487 4696 3664 4704
rect 3656 4687 3664 4696
rect 3767 4696 3833 4704
rect 3967 4696 4013 4704
rect 4187 4696 4413 4704
rect 5127 4696 5153 4704
rect 5347 4696 5413 4704
rect 287 4676 373 4684
rect 667 4676 793 4684
rect 807 4676 1013 4684
rect 1167 4676 1213 4684
rect 1267 4676 1353 4684
rect 1367 4676 1493 4684
rect 1547 4676 1573 4684
rect 1787 4676 1993 4684
rect 2087 4676 2353 4684
rect 2407 4676 2433 4684
rect 2527 4676 2813 4684
rect 3087 4676 3253 4684
rect 3347 4676 3413 4684
rect 3507 4676 3633 4684
rect 3767 4676 3853 4684
rect 3867 4676 4173 4684
rect 4307 4676 4333 4684
rect 4347 4676 4433 4684
rect 4487 4676 4533 4684
rect 4707 4676 5033 4684
rect 5087 4676 5173 4684
rect 5316 4684 5324 4693
rect 5316 4676 5433 4684
rect 5456 4684 5464 4693
rect 5456 4676 5553 4684
rect 256 4656 273 4664
rect 467 4656 533 4664
rect 887 4656 1233 4664
rect 1627 4656 1713 4664
rect 1807 4656 1953 4664
rect 2107 4656 2193 4664
rect 2207 4656 2253 4664
rect 2267 4656 2273 4664
rect 2407 4656 2573 4664
rect 2587 4656 2633 4664
rect 2647 4656 2733 4664
rect 2787 4656 2964 4664
rect 127 4636 193 4644
rect 247 4636 313 4644
rect 367 4636 453 4644
rect 1067 4636 1133 4644
rect 1147 4636 1213 4644
rect 1267 4636 1373 4644
rect 1527 4636 1593 4644
rect 1727 4636 2033 4644
rect 2187 4636 2773 4644
rect 2956 4644 2964 4656
rect 3107 4656 3173 4664
rect 3547 4656 3613 4664
rect 4007 4656 4573 4664
rect 4967 4656 5013 4664
rect 5127 4656 5313 4664
rect 5387 4656 5433 4664
rect 5587 4656 5593 4664
rect 5607 4656 5693 4664
rect 5747 4656 5773 4664
rect 2956 4636 3173 4644
rect 3267 4636 3453 4644
rect 3507 4636 3633 4644
rect 3747 4636 3813 4644
rect 3907 4636 4073 4644
rect 4147 4636 4173 4644
rect 4467 4636 4593 4644
rect 4607 4636 4673 4644
rect 4687 4636 4733 4644
rect 4887 4636 5053 4644
rect 5207 4636 5333 4644
rect 5367 4636 5453 4644
rect 267 4616 353 4624
rect 1327 4616 1473 4624
rect 1607 4616 2244 4624
rect 527 4596 833 4604
rect 847 4596 893 4604
rect 907 4596 1673 4604
rect 2236 4604 2244 4616
rect 2327 4616 2673 4624
rect 2927 4616 3353 4624
rect 3787 4616 3893 4624
rect 4096 4616 4253 4624
rect 2236 4596 2513 4604
rect 2687 4596 3293 4604
rect 3307 4596 3653 4604
rect 3727 4596 3933 4604
rect 4096 4604 4104 4616
rect 4827 4616 4933 4624
rect 5027 4616 5513 4624
rect 5527 4616 5713 4624
rect 4047 4596 4104 4604
rect 4247 4596 4533 4604
rect 4907 4596 5073 4604
rect 5327 4596 5393 4604
rect 147 4576 493 4584
rect 1387 4576 1433 4584
rect 1847 4576 2093 4584
rect 2467 4576 2673 4584
rect 2687 4576 2893 4584
rect 2907 4576 3013 4584
rect 4247 4576 4553 4584
rect 4567 4576 4833 4584
rect 247 4556 413 4564
rect 427 4556 693 4564
rect 1007 4556 1933 4564
rect 2287 4556 2593 4564
rect 2767 4556 2833 4564
rect 2847 4556 3213 4564
rect 3827 4556 3933 4564
rect 3947 4556 5293 4564
rect 507 4536 573 4544
rect 647 4536 653 4544
rect 667 4536 853 4544
rect 867 4536 933 4544
rect 1287 4536 1393 4544
rect 1407 4536 1433 4544
rect 1447 4536 1753 4544
rect 1827 4536 2173 4544
rect 3227 4536 3253 4544
rect 4127 4536 4313 4544
rect 4327 4536 4473 4544
rect 5147 4536 5293 4544
rect 587 4516 713 4524
rect 907 4516 1533 4524
rect 1667 4516 1973 4524
rect 2027 4516 2493 4524
rect 2507 4516 2573 4524
rect 2887 4516 2913 4524
rect 3127 4516 3453 4524
rect 3467 4516 3473 4524
rect 3667 4516 4053 4524
rect 4067 4516 4093 4524
rect 4487 4516 5093 4524
rect 5167 4516 5213 4524
rect 5307 4516 5353 4524
rect 5507 4516 5593 4524
rect 107 4496 153 4504
rect 267 4496 353 4504
rect 687 4496 773 4504
rect 787 4496 813 4504
rect 827 4496 893 4504
rect 1187 4496 1273 4504
rect 1296 4496 1313 4504
rect 56 4424 64 4493
rect 116 4476 293 4484
rect 116 4467 124 4476
rect 307 4476 393 4484
rect 607 4476 673 4484
rect 727 4476 824 4484
rect 287 4456 333 4464
rect 387 4456 413 4464
rect 567 4456 693 4464
rect 707 4456 793 4464
rect 816 4464 824 4476
rect 947 4476 1013 4484
rect 1296 4484 1304 4496
rect 1807 4496 2213 4504
rect 2487 4496 2613 4504
rect 2727 4496 2853 4504
rect 3027 4496 3133 4504
rect 3147 4496 3213 4504
rect 3227 4496 3313 4504
rect 3527 4496 3893 4504
rect 4027 4496 4113 4504
rect 4867 4496 5173 4504
rect 5187 4496 5333 4504
rect 1187 4476 1304 4484
rect 1467 4476 1493 4484
rect 1567 4476 1913 4484
rect 1927 4476 2013 4484
rect 2047 4476 2173 4484
rect 2227 4476 2764 4484
rect 2756 4467 2764 4476
rect 2887 4476 2993 4484
rect 3387 4476 3533 4484
rect 3547 4476 3584 4484
rect 816 4456 913 4464
rect 927 4456 993 4464
rect 1047 4456 1153 4464
rect 1207 4456 1333 4464
rect 1347 4456 1413 4464
rect 1447 4456 1713 4464
rect 1847 4456 1933 4464
rect 2067 4456 2153 4464
rect 2367 4456 2413 4464
rect 2447 4456 2473 4464
rect 2527 4456 2733 4464
rect 2947 4456 2973 4464
rect 3356 4464 3364 4473
rect 3356 4456 3553 4464
rect 3576 4464 3584 4476
rect 3607 4476 3633 4484
rect 3707 4476 3793 4484
rect 4267 4476 4393 4484
rect 4427 4476 4524 4484
rect 3576 4456 3753 4464
rect 76 4444 84 4453
rect 3656 4447 3664 4456
rect 3827 4456 3853 4464
rect 4307 4456 4353 4464
rect 4367 4456 4393 4464
rect 4516 4447 4524 4476
rect 4887 4476 4933 4484
rect 4947 4476 4973 4484
rect 5227 4476 5393 4484
rect 5496 4464 5504 4493
rect 5147 4456 5504 4464
rect 5676 4447 5684 4473
rect 76 4436 173 4444
rect 187 4436 213 4444
rect 347 4436 393 4444
rect 467 4436 533 4444
rect 1087 4436 1293 4444
rect 1307 4436 1353 4444
rect 1796 4436 1813 4444
rect 56 4416 73 4424
rect 256 4424 264 4433
rect 1796 4427 1804 4436
rect 2607 4436 2713 4444
rect 3007 4436 3333 4444
rect 3347 4436 3593 4444
rect 3707 4436 3873 4444
rect 4047 4436 4273 4444
rect 4447 4436 4493 4444
rect 4787 4436 4893 4444
rect 4947 4436 5013 4444
rect 5367 4436 5473 4444
rect 256 4416 333 4424
rect 1107 4416 1153 4424
rect 1527 4416 1553 4424
rect 1567 4416 1593 4424
rect 2076 4424 2084 4433
rect 2067 4416 2084 4424
rect 2347 4416 3633 4424
rect 4167 4416 4373 4424
rect 4807 4416 4993 4424
rect 5067 4416 5193 4424
rect 5387 4416 5413 4424
rect 5587 4416 5733 4424
rect 1707 4396 2333 4404
rect 2667 4396 3333 4404
rect 3527 4396 3613 4404
rect 4287 4396 4313 4404
rect 4327 4396 4333 4404
rect 4707 4396 4933 4404
rect 4947 4396 5133 4404
rect 5207 4396 5533 4404
rect 1827 4376 1853 4384
rect 2647 4376 3153 4384
rect 3647 4376 4273 4384
rect 1367 4356 2333 4364
rect 2747 4356 3033 4364
rect 4627 4356 4653 4364
rect 1487 4336 2373 4344
rect 2467 4336 2933 4344
rect 2947 4336 2993 4344
rect 3047 4336 4593 4344
rect 2227 4316 2413 4324
rect 2427 4316 4733 4324
rect 907 4296 2433 4304
rect 2707 4296 4233 4304
rect 4567 4296 4613 4304
rect 4627 4296 4913 4304
rect 5567 4296 5613 4304
rect 1687 4276 1853 4284
rect 2167 4276 2193 4284
rect 2967 4276 3313 4284
rect 387 4256 433 4264
rect 1267 4256 1293 4264
rect 1327 4256 1733 4264
rect 1847 4256 1893 4264
rect 1947 4256 2093 4264
rect 2127 4256 2353 4264
rect 2467 4256 2513 4264
rect 2727 4256 3593 4264
rect 3927 4256 4173 4264
rect 4187 4256 4193 4264
rect 1187 4236 1373 4244
rect 1527 4236 2053 4244
rect 2187 4236 2233 4244
rect 2276 4236 2493 4244
rect 816 4216 1033 4224
rect 816 4207 824 4216
rect 1047 4216 1213 4224
rect 1267 4216 1293 4224
rect 1487 4216 1653 4224
rect 1767 4216 1793 4224
rect 2047 4216 2073 4224
rect 2276 4224 2284 4236
rect 2836 4236 2893 4244
rect 2836 4227 2844 4236
rect 3027 4236 3573 4244
rect 3987 4236 4033 4244
rect 4047 4236 4093 4244
rect 5307 4236 5524 4244
rect 2147 4216 2284 4224
rect 2407 4216 2713 4224
rect 147 4196 213 4204
rect 227 4196 273 4204
rect 467 4196 593 4204
rect 767 4196 813 4204
rect 867 4196 913 4204
rect 1147 4196 1233 4204
rect 47 4176 113 4184
rect 156 4176 173 4184
rect 156 4164 164 4176
rect 267 4176 333 4184
rect 736 4184 744 4193
rect 736 4176 833 4184
rect 1076 4184 1084 4193
rect 1356 4187 1364 4213
rect 2636 4207 2644 4216
rect 2727 4216 2773 4224
rect 2887 4216 2953 4224
rect 3687 4216 3773 4224
rect 3816 4216 3913 4224
rect 1387 4196 1433 4204
rect 1547 4196 1613 4204
rect 1787 4196 1933 4204
rect 1947 4196 1973 4204
rect 2027 4196 2124 4204
rect 2116 4187 2124 4196
rect 2167 4196 2193 4204
rect 2216 4196 2593 4204
rect 1076 4176 1273 4184
rect 1607 4176 1673 4184
rect 1747 4176 1873 4184
rect 2067 4176 2093 4184
rect 2216 4184 2224 4196
rect 2727 4196 2913 4204
rect 3247 4196 3264 4204
rect 2127 4176 2224 4184
rect 2247 4176 2273 4184
rect 2367 4176 2433 4184
rect 2607 4176 3033 4184
rect 147 4156 164 4164
rect 187 4156 233 4164
rect 247 4156 573 4164
rect 827 4156 913 4164
rect 927 4156 933 4164
rect 947 4156 1053 4164
rect 1207 4156 1613 4164
rect 1727 4156 1813 4164
rect 1907 4156 1993 4164
rect 2007 4156 2133 4164
rect 2307 4156 2333 4164
rect 2487 4156 2873 4164
rect 2907 4156 3113 4164
rect 3127 4156 3233 4164
rect 3256 4164 3264 4196
rect 3296 4196 3373 4204
rect 3296 4184 3304 4196
rect 3427 4196 3453 4204
rect 3507 4196 3533 4204
rect 3816 4204 3824 4216
rect 4067 4216 4133 4224
rect 4567 4216 4593 4224
rect 5167 4216 5184 4224
rect 3807 4196 3824 4204
rect 3847 4196 3933 4204
rect 4207 4196 4333 4204
rect 4347 4196 4444 4204
rect 4436 4187 4444 4196
rect 4487 4196 4613 4204
rect 5007 4196 5093 4204
rect 3287 4176 3304 4184
rect 3316 4176 3353 4184
rect 3316 4164 3324 4176
rect 3607 4176 3633 4184
rect 3647 4176 3733 4184
rect 3987 4176 4053 4184
rect 4207 4176 4233 4184
rect 4327 4176 4393 4184
rect 4687 4176 4753 4184
rect 5176 4184 5184 4216
rect 5287 4216 5304 4224
rect 5296 4207 5304 4216
rect 5207 4196 5253 4204
rect 5407 4196 5493 4204
rect 5516 4204 5524 4236
rect 5687 4216 5704 4224
rect 5516 4196 5673 4204
rect 5176 4176 5464 4184
rect 3256 4156 3324 4164
rect 3347 4156 3373 4164
rect 3487 4156 3513 4164
rect 3527 4156 3553 4164
rect 3627 4156 3653 4164
rect 3667 4156 3993 4164
rect 4387 4156 4413 4164
rect 4647 4156 4653 4164
rect 4667 4156 4853 4164
rect 4887 4156 5053 4164
rect 5187 4156 5373 4164
rect 5407 4156 5433 4164
rect 5456 4164 5464 4176
rect 5487 4176 5573 4184
rect 5696 4184 5704 4216
rect 5667 4176 5704 4184
rect 5456 4156 5533 4164
rect 5776 4164 5784 4173
rect 5667 4156 5784 4164
rect 227 4136 253 4144
rect 587 4136 1693 4144
rect 1716 4136 2413 4144
rect 67 4116 113 4124
rect 247 4116 413 4124
rect 427 4116 553 4124
rect 567 4116 653 4124
rect 1107 4116 1253 4124
rect 1567 4116 1613 4124
rect 1716 4124 1724 4136
rect 2427 4136 2553 4144
rect 2687 4136 2713 4144
rect 2867 4136 4493 4144
rect 4507 4136 4713 4144
rect 4827 4136 4993 4144
rect 5227 4136 5373 4144
rect 5727 4136 5773 4144
rect 1647 4116 1724 4124
rect 2407 4116 2513 4124
rect 2527 4116 2693 4124
rect 2767 4116 2953 4124
rect 3087 4116 3133 4124
rect 3167 4116 3213 4124
rect 3247 4116 3493 4124
rect 4307 4116 4333 4124
rect 4407 4116 4573 4124
rect 4587 4116 5113 4124
rect 5367 4116 5473 4124
rect 67 4096 93 4104
rect 107 4096 433 4104
rect 447 4096 453 4104
rect 647 4096 733 4104
rect 747 4096 1973 4104
rect 2067 4096 2253 4104
rect 2327 4096 2413 4104
rect 2847 4096 3053 4104
rect 3067 4096 3193 4104
rect 3287 4096 3393 4104
rect 3447 4096 3493 4104
rect 4167 4096 4293 4104
rect 4947 4096 5113 4104
rect 5127 4096 5233 4104
rect 167 4076 293 4084
rect 1247 4076 2833 4084
rect 2856 4076 3313 4084
rect 367 4056 413 4064
rect 427 4056 593 4064
rect 607 4056 1993 4064
rect 2856 4064 2864 4076
rect 3347 4076 3393 4084
rect 3647 4076 3713 4084
rect 3747 4076 3873 4084
rect 3887 4076 5273 4084
rect 5467 4076 5493 4084
rect 2047 4056 2864 4064
rect 2987 4056 3153 4064
rect 3227 4056 3333 4064
rect 3347 4056 3553 4064
rect 3727 4056 3793 4064
rect 3807 4056 4093 4064
rect 4147 4056 4173 4064
rect 5247 4056 5293 4064
rect 5327 4056 5513 4064
rect 167 4036 193 4044
rect 307 4036 553 4044
rect 567 4036 613 4044
rect 887 4036 953 4044
rect 967 4036 1493 4044
rect 1547 4036 1553 4044
rect 1567 4036 1813 4044
rect 2167 4036 2813 4044
rect 2887 4036 3133 4044
rect 3307 4036 3353 4044
rect 3587 4036 3773 4044
rect 3907 4036 4133 4044
rect 4147 4036 4253 4044
rect 4387 4036 5193 4044
rect 5267 4036 5413 4044
rect 5527 4036 5693 4044
rect 107 4016 173 4024
rect 987 4016 1093 4024
rect 1287 4016 1333 4024
rect 1347 4016 1633 4024
rect 1667 4016 1753 4024
rect 1767 4016 1833 4024
rect 2187 4016 2273 4024
rect 2287 4016 2493 4024
rect 2887 4016 2993 4024
rect 3047 4016 3093 4024
rect 3187 4016 3284 4024
rect 76 3984 84 4013
rect 167 3996 213 4004
rect 607 3996 713 4004
rect 867 3996 913 4004
rect 1407 3996 1453 4004
rect 1467 3996 1613 4004
rect 1887 3996 2293 4004
rect 2307 3996 2333 4004
rect 2387 3996 2433 4004
rect 2647 3996 2673 4004
rect 2827 3996 3253 4004
rect 76 3976 93 3984
rect 207 3976 253 3984
rect 267 3976 333 3984
rect 487 3976 553 3984
rect 747 3976 833 3984
rect 856 3976 1344 3984
rect 147 3956 173 3964
rect 856 3964 864 3976
rect 727 3956 864 3964
rect 987 3956 1073 3964
rect 1227 3956 1313 3964
rect 1336 3964 1344 3976
rect 1647 3976 1693 3984
rect 1867 3976 1893 3984
rect 1987 3976 2073 3984
rect 2207 3976 2233 3984
rect 1336 3956 2133 3964
rect 1167 3936 1313 3944
rect 1387 3936 1553 3944
rect 1987 3936 2013 3944
rect 2156 3944 2164 3973
rect 2416 3964 2424 3973
rect 2327 3956 2424 3964
rect 2476 3964 2484 3993
rect 3276 3987 3284 4016
rect 3327 4016 4713 4024
rect 4767 4016 4913 4024
rect 5167 4016 5413 4024
rect 3447 3996 3753 4004
rect 3947 3996 3973 4004
rect 4027 3996 4073 4004
rect 4087 3996 4333 4004
rect 4547 3996 4593 4004
rect 4667 3996 4973 4004
rect 5307 3996 5333 4004
rect 5347 3996 5513 4004
rect 5567 3996 5733 4004
rect 2507 3976 2613 3984
rect 2627 3976 2753 3984
rect 2787 3976 2913 3984
rect 2967 3976 2993 3984
rect 3327 3976 3413 3984
rect 3536 3976 3833 3984
rect 3536 3967 3544 3976
rect 3847 3976 3953 3984
rect 4007 3976 4113 3984
rect 4127 3976 4233 3984
rect 4247 3976 4353 3984
rect 4407 3976 4433 3984
rect 4516 3984 4524 3993
rect 4516 3976 4873 3984
rect 4816 3967 4824 3976
rect 4907 3976 5013 3984
rect 5036 3976 5113 3984
rect 2476 3956 2493 3964
rect 2527 3956 2553 3964
rect 2607 3956 2633 3964
rect 2767 3956 2793 3964
rect 2987 3956 3033 3964
rect 3267 3956 3484 3964
rect 2696 3944 2704 3953
rect 2156 3936 2873 3944
rect 2936 3944 2944 3953
rect 2936 3936 2953 3944
rect 3067 3936 3453 3944
rect 3476 3944 3484 3956
rect 3587 3956 3673 3964
rect 4007 3956 4033 3964
rect 4687 3956 4753 3964
rect 4767 3956 4773 3964
rect 5036 3964 5044 3976
rect 5427 3976 5493 3984
rect 4947 3956 5044 3964
rect 5147 3956 5713 3964
rect 5756 3964 5764 3973
rect 5747 3956 5764 3964
rect 3476 3936 3713 3944
rect 3867 3936 4193 3944
rect 4207 3936 4213 3944
rect 5107 3936 5653 3944
rect 5767 3936 5813 3944
rect 2467 3916 2613 3924
rect 2627 3916 2673 3924
rect 3007 3916 3493 3924
rect 3787 3916 4473 3924
rect 4727 3916 5133 3924
rect 5687 3916 5713 3924
rect 1307 3896 2993 3904
rect 3027 3896 4413 3904
rect 4747 3896 4913 3904
rect 2407 3876 2453 3884
rect 2487 3876 2513 3884
rect 2547 3876 2613 3884
rect 2667 3876 2953 3884
rect 2967 3876 3224 3884
rect 1107 3856 1253 3864
rect 1687 3856 2753 3864
rect 3216 3864 3224 3876
rect 3247 3876 4333 3884
rect 4387 3876 4853 3884
rect 5227 3876 5393 3884
rect 3216 3856 4813 3864
rect 1307 3836 3113 3844
rect 3147 3836 3233 3844
rect 3267 3836 3373 3844
rect 3827 3836 4253 3844
rect 4267 3836 4533 3844
rect 1087 3816 1173 3824
rect 2387 3816 2733 3824
rect 3307 3816 3333 3824
rect 3527 3816 3893 3824
rect 4707 3816 4853 3824
rect 5447 3816 5813 3824
rect 1047 3796 1213 3804
rect 2067 3796 2073 3804
rect 2087 3796 2393 3804
rect 2487 3796 2653 3804
rect 2827 3796 2953 3804
rect 3127 3796 3353 3804
rect 3647 3796 4593 3804
rect 4687 3796 5133 3804
rect 5147 3796 5253 3804
rect 67 3776 113 3784
rect 2707 3776 3913 3784
rect 3927 3776 4753 3784
rect 5627 3776 5693 3784
rect 127 3756 244 3764
rect 236 3747 244 3756
rect 967 3756 1013 3764
rect 1127 3756 1173 3764
rect 1256 3756 1333 3764
rect 1256 3747 1264 3756
rect 1407 3756 1533 3764
rect 1827 3756 1873 3764
rect 1907 3756 1993 3764
rect 2007 3756 2133 3764
rect 2347 3756 2573 3764
rect 2847 3756 3293 3764
rect 3387 3756 3553 3764
rect 3847 3756 4493 3764
rect 5027 3756 5153 3764
rect 5167 3756 5713 3764
rect 5747 3756 5784 3764
rect 87 3736 184 3744
rect 176 3724 184 3736
rect 207 3736 224 3744
rect 216 3724 224 3736
rect 247 3736 313 3744
rect 667 3736 733 3744
rect 747 3736 993 3744
rect 1167 3736 1193 3744
rect 1347 3736 1433 3744
rect 1687 3736 1873 3744
rect 1887 3736 2033 3744
rect 2067 3736 2173 3744
rect 2327 3736 2424 3744
rect 176 3716 204 3724
rect 216 3716 293 3724
rect 87 3696 133 3704
rect 196 3704 204 3716
rect 427 3716 493 3724
rect 607 3716 813 3724
rect 1116 3724 1124 3733
rect 867 3716 924 3724
rect 1116 3716 1233 3724
rect 196 3696 213 3704
rect 267 3696 333 3704
rect 447 3696 453 3704
rect 467 3696 533 3704
rect 567 3696 713 3704
rect 816 3704 824 3713
rect 747 3696 824 3704
rect 847 3696 893 3704
rect 916 3704 924 3716
rect 1427 3716 1453 3724
rect 1467 3716 1493 3724
rect 916 3696 1013 3704
rect 1376 3704 1384 3713
rect 1147 3696 1384 3704
rect 1396 3704 1404 3713
rect 1516 3707 1524 3733
rect 2416 3727 2424 3736
rect 2576 3736 2693 3744
rect 1587 3716 1733 3724
rect 1907 3716 1993 3724
rect 2107 3716 2273 3724
rect 2467 3716 2553 3724
rect 1396 3696 1433 3704
rect 1567 3696 1753 3704
rect 1967 3696 2093 3704
rect 2127 3696 2293 3704
rect 2576 3704 2584 3736
rect 2807 3736 3033 3744
rect 3247 3736 3313 3744
rect 3367 3736 3413 3744
rect 3467 3736 3573 3744
rect 3727 3736 3773 3744
rect 5067 3736 5233 3744
rect 5247 3736 5493 3744
rect 5627 3736 5753 3744
rect 2687 3716 2704 3724
rect 2487 3696 2584 3704
rect 2696 3704 2704 3716
rect 2727 3716 2833 3724
rect 3076 3724 3084 3733
rect 2927 3716 3213 3724
rect 3347 3716 3433 3724
rect 3747 3716 4013 3724
rect 4027 3716 4133 3724
rect 4436 3724 4444 3733
rect 4416 3716 4444 3724
rect 2696 3696 2713 3704
rect 2947 3696 2993 3704
rect 3047 3696 3113 3704
rect 3647 3696 3693 3704
rect 4087 3696 4213 3704
rect 4376 3687 4384 3713
rect 4416 3704 4424 3716
rect 4527 3716 4633 3724
rect 4807 3716 5033 3724
rect 5247 3716 5293 3724
rect 5307 3716 5364 3724
rect 4407 3696 4424 3704
rect 4447 3696 4453 3704
rect 4467 3696 4653 3704
rect 4747 3696 5153 3704
rect 5356 3704 5364 3716
rect 5447 3716 5544 3724
rect 5356 3696 5513 3704
rect 5536 3704 5544 3716
rect 5776 3724 5784 3756
rect 5747 3716 5784 3724
rect 5536 3696 5713 3704
rect 627 3676 773 3684
rect 1027 3676 1093 3684
rect 1276 3676 1484 3684
rect 1276 3664 1284 3676
rect 587 3656 1284 3664
rect 1296 3656 1393 3664
rect 1296 3644 1304 3656
rect 1476 3664 1484 3676
rect 1507 3676 1653 3684
rect 1987 3676 2033 3684
rect 2047 3676 2593 3684
rect 2707 3676 2793 3684
rect 2807 3676 2833 3684
rect 2987 3676 3133 3684
rect 3307 3676 3333 3684
rect 3567 3676 3613 3684
rect 4427 3676 4473 3684
rect 4567 3676 4633 3684
rect 4887 3676 5073 3684
rect 5087 3676 5113 3684
rect 1476 3656 1933 3664
rect 1947 3656 1993 3664
rect 2267 3656 2513 3664
rect 2527 3656 2633 3664
rect 2647 3656 2933 3664
rect 3087 3656 3733 3664
rect 3807 3656 3833 3664
rect 4147 3656 4753 3664
rect 5567 3656 5673 3664
rect 727 3636 1304 3644
rect 1327 3636 1373 3644
rect 1567 3636 1593 3644
rect 1907 3636 2433 3644
rect 2527 3636 2733 3644
rect 3267 3636 3273 3644
rect 3287 3636 3673 3644
rect 3907 3636 3993 3644
rect 1207 3616 1213 3624
rect 1227 3616 1273 3624
rect 1607 3616 2213 3624
rect 2607 3616 2733 3624
rect 2747 3616 3633 3624
rect 3687 3616 3893 3624
rect 3987 3616 4033 3624
rect 5367 3616 5453 3624
rect 107 3596 213 3604
rect 1387 3596 3073 3604
rect 3107 3596 3873 3604
rect 4167 3596 4673 3604
rect 4747 3596 4773 3604
rect 107 3576 273 3584
rect 307 3576 413 3584
rect 687 3576 893 3584
rect 907 3576 973 3584
rect 1767 3576 2253 3584
rect 2407 3576 2433 3584
rect 2907 3576 3173 3584
rect 3327 3576 3393 3584
rect 3547 3576 3613 3584
rect 3627 3576 3773 3584
rect 4207 3576 4293 3584
rect 4367 3576 4893 3584
rect 5187 3576 5233 3584
rect 147 3556 373 3564
rect 507 3556 1113 3564
rect 1727 3556 1993 3564
rect 2287 3556 3553 3564
rect 3667 3556 4193 3564
rect 4287 3556 4653 3564
rect 5047 3556 5313 3564
rect 116 3536 213 3544
rect 116 3507 124 3536
rect 387 3536 613 3544
rect 967 3536 1053 3544
rect 1667 3536 1713 3544
rect 1927 3536 1953 3544
rect 2187 3536 2333 3544
rect 2347 3536 2393 3544
rect 3007 3536 3033 3544
rect 3067 3536 3393 3544
rect 3427 3536 3493 3544
rect 3707 3536 4053 3544
rect 4167 3536 4213 3544
rect 4267 3536 4573 3544
rect 4687 3536 4693 3544
rect 4707 3536 5333 3544
rect 5387 3536 5633 3544
rect 147 3516 204 3524
rect 196 3507 204 3516
rect 267 3516 293 3524
rect 487 3516 593 3524
rect 927 3516 1093 3524
rect 1107 3516 1153 3524
rect 1347 3516 1413 3524
rect 1536 3516 1673 3524
rect 1536 3507 1544 3516
rect 1847 3516 2013 3524
rect 2067 3516 2153 3524
rect 2167 3516 2293 3524
rect 247 3496 273 3504
rect 407 3496 453 3504
rect 947 3496 993 3504
rect 1287 3496 1333 3504
rect 1587 3496 1613 3504
rect 1787 3496 1853 3504
rect 1887 3496 1913 3504
rect 2027 3496 2093 3504
rect 2147 3496 2173 3504
rect 76 3484 84 3493
rect -24 3476 553 3484
rect 1036 3484 1044 3493
rect 927 3476 1044 3484
rect 1187 3476 1253 3484
rect 1367 3476 1393 3484
rect 1456 3484 1464 3493
rect 1456 3476 1613 3484
rect 1667 3476 1693 3484
rect 1707 3476 1813 3484
rect 1987 3476 2213 3484
rect 2236 3484 2244 3516
rect 2367 3516 2533 3524
rect 2587 3516 2813 3524
rect 2887 3516 3053 3524
rect 3516 3524 3524 3533
rect 3207 3516 3524 3524
rect 3656 3516 3753 3524
rect 3656 3507 3664 3516
rect 3776 3516 3873 3524
rect 2267 3496 2333 3504
rect 2387 3496 2453 3504
rect 2476 3496 2673 3504
rect 2476 3484 2484 3496
rect 2696 3496 2733 3504
rect 2696 3487 2704 3496
rect 2807 3496 2873 3504
rect 3067 3496 3173 3504
rect 3227 3496 3253 3504
rect 3316 3496 3353 3504
rect 2236 3476 2484 3484
rect 2567 3476 2653 3484
rect 2727 3476 2833 3484
rect 2867 3476 3193 3484
rect 3316 3484 3324 3496
rect 3367 3496 3473 3504
rect 3527 3496 3653 3504
rect 3776 3487 3784 3516
rect 4007 3516 4313 3524
rect 4327 3516 4613 3524
rect 5087 3516 5133 3524
rect 5147 3516 5153 3524
rect 5307 3516 5533 3524
rect 5587 3516 5593 3524
rect 5607 3516 5633 3524
rect 3916 3504 3924 3513
rect 3847 3496 4033 3504
rect 4127 3496 4173 3504
rect 4187 3496 4273 3504
rect 4327 3496 4393 3504
rect 4447 3496 4473 3504
rect 4507 3496 4533 3504
rect 4927 3496 4973 3504
rect 5027 3496 5173 3504
rect 5527 3496 5553 3504
rect 5667 3496 5733 3504
rect 3247 3476 3324 3484
rect 3347 3476 3364 3484
rect 147 3456 173 3464
rect 807 3456 893 3464
rect 1107 3456 1293 3464
rect 1436 3464 1444 3473
rect 3356 3467 3364 3476
rect 3387 3476 3453 3484
rect 3507 3476 3764 3484
rect 1427 3456 1444 3464
rect 1647 3456 1753 3464
rect 1947 3456 2353 3464
rect 3027 3456 3053 3464
rect 3127 3456 3204 3464
rect 107 3436 113 3444
rect 567 3436 593 3444
rect 827 3436 873 3444
rect 887 3436 953 3444
rect 1307 3436 1373 3444
rect 2047 3436 2273 3444
rect 3196 3444 3204 3456
rect 3267 3456 3333 3464
rect 3427 3456 3673 3464
rect 3756 3464 3764 3476
rect 3987 3476 4173 3484
rect 4467 3476 4513 3484
rect 4527 3476 4893 3484
rect 4907 3476 4993 3484
rect 5167 3476 5373 3484
rect 5507 3476 5533 3484
rect 3756 3456 3793 3464
rect 4087 3456 4373 3464
rect 4527 3456 4613 3464
rect 4847 3456 5053 3464
rect 5127 3456 5133 3464
rect 5147 3456 5193 3464
rect 5607 3456 5713 3464
rect 2287 3436 3184 3444
rect 3196 3436 3413 3444
rect 2567 3416 2913 3424
rect 3176 3424 3184 3436
rect 3436 3436 3493 3444
rect 3436 3424 3444 3436
rect 4827 3436 5433 3444
rect 5587 3436 5653 3444
rect 3176 3416 3444 3424
rect 3467 3416 3693 3424
rect 4367 3416 4833 3424
rect 1487 3396 2113 3404
rect 3107 3396 3153 3404
rect 3236 3396 3313 3404
rect 2007 3376 2853 3384
rect 3236 3384 3244 3396
rect 3327 3396 3593 3404
rect 3707 3396 3833 3404
rect 2927 3376 3244 3384
rect 3567 3376 3913 3384
rect 4007 3376 4593 3384
rect 5447 3376 5473 3384
rect 1047 3356 2553 3364
rect 2667 3356 3353 3364
rect 3427 3356 4013 3364
rect 4947 3356 4973 3364
rect 2767 3336 2793 3344
rect 2807 3336 3113 3344
rect 3147 3336 3193 3344
rect 3247 3336 3293 3344
rect 3307 3336 4153 3344
rect 1087 3316 1233 3324
rect 2627 3316 2753 3324
rect 3047 3316 3153 3324
rect 3327 3316 3573 3324
rect 4147 3316 4213 3324
rect 367 3296 413 3304
rect 667 3296 673 3304
rect 687 3296 833 3304
rect 847 3296 1353 3304
rect 1787 3296 1933 3304
rect 2087 3296 2313 3304
rect 2327 3296 2413 3304
rect 2687 3296 2873 3304
rect 2927 3296 3324 3304
rect 267 3276 313 3284
rect 327 3276 393 3284
rect 1187 3276 1253 3284
rect 1267 3276 1493 3284
rect 1567 3276 1733 3284
rect 1656 3267 1664 3276
rect 1827 3276 2013 3284
rect 2207 3276 2253 3284
rect 2587 3276 2653 3284
rect 2787 3276 3073 3284
rect 3087 3276 3293 3284
rect 3316 3284 3324 3296
rect 3316 3276 3453 3284
rect 3467 3276 3613 3284
rect 4567 3276 4573 3284
rect 4587 3276 4713 3284
rect 4727 3276 4813 3284
rect 4827 3276 4893 3284
rect 4907 3276 4953 3284
rect 4967 3276 5253 3284
rect 5527 3276 5553 3284
rect 87 3256 273 3264
rect 327 3256 553 3264
rect 707 3256 873 3264
rect 887 3256 913 3264
rect 927 3256 953 3264
rect 1007 3256 1093 3264
rect 1227 3256 1473 3264
rect 1587 3256 1613 3264
rect 1927 3256 2133 3264
rect 2207 3256 2233 3264
rect 2487 3256 2713 3264
rect 2816 3256 2933 3264
rect 2816 3247 2824 3256
rect 2976 3256 3153 3264
rect 107 3236 173 3244
rect 227 3236 313 3244
rect 427 3236 513 3244
rect 1127 3236 1213 3244
rect 1267 3236 1373 3244
rect 1447 3236 1593 3244
rect 1647 3236 1713 3244
rect 1807 3236 2084 3244
rect 147 3216 173 3224
rect 247 3216 273 3224
rect 407 3216 453 3224
rect 727 3216 753 3224
rect 767 3216 913 3224
rect 1236 3224 1244 3233
rect 1187 3216 1244 3224
rect 1527 3216 1673 3224
rect 2076 3224 2084 3236
rect 2107 3236 2173 3244
rect 2767 3236 2793 3244
rect 2847 3236 2913 3244
rect 2076 3216 2193 3224
rect 2247 3216 2293 3224
rect 2407 3216 2573 3224
rect 2596 3224 2604 3233
rect 2596 3216 2693 3224
rect 107 3196 253 3204
rect 887 3196 973 3204
rect 1507 3196 1553 3204
rect 1807 3196 1893 3204
rect 1907 3196 1933 3204
rect 2227 3196 2373 3204
rect 2667 3196 2733 3204
rect 2976 3204 2984 3256
rect 3167 3256 3233 3264
rect 3407 3256 3473 3264
rect 3687 3256 3953 3264
rect 4027 3256 4233 3264
rect 4307 3256 4484 3264
rect 3387 3236 3533 3244
rect 3547 3236 3593 3244
rect 3847 3236 3893 3244
rect 3967 3236 4093 3244
rect 4207 3236 4233 3244
rect 4427 3236 4453 3244
rect 4476 3244 4484 3256
rect 4947 3256 5153 3264
rect 5307 3256 5613 3264
rect 5627 3256 5693 3264
rect 4476 3236 4913 3244
rect 5067 3236 5153 3244
rect 5387 3236 5493 3244
rect 3027 3216 3053 3224
rect 3347 3216 3533 3224
rect 2867 3196 2984 3204
rect 3047 3196 3353 3204
rect 3367 3196 3553 3204
rect 3636 3204 3644 3233
rect 3667 3216 3693 3224
rect 4376 3224 4384 3233
rect 3847 3216 4384 3224
rect 4607 3216 4773 3224
rect 4807 3216 4824 3224
rect 3636 3196 3693 3204
rect 3887 3196 3913 3204
rect 4227 3196 4573 3204
rect 4667 3196 4793 3204
rect 4816 3204 4824 3216
rect 4887 3216 4933 3224
rect 4967 3216 4973 3224
rect 4987 3216 5073 3224
rect 5087 3216 5473 3224
rect 5487 3216 5633 3224
rect 4816 3196 5273 3204
rect 87 3176 113 3184
rect 647 3176 973 3184
rect 1147 3176 1233 3184
rect 1247 3176 1793 3184
rect 2567 3176 2653 3184
rect 2927 3176 3093 3184
rect 3447 3176 3913 3184
rect 4087 3176 4253 3184
rect 4347 3176 4373 3184
rect 4427 3176 4553 3184
rect 4567 3176 4673 3184
rect 867 3156 933 3164
rect 947 3156 993 3164
rect 1007 3156 1213 3164
rect 1767 3156 1893 3164
rect 2327 3156 2613 3164
rect 2627 3156 3093 3164
rect 3147 3156 3193 3164
rect 3207 3156 3353 3164
rect 3527 3156 3613 3164
rect 3627 3156 3773 3164
rect 3807 3156 3993 3164
rect 4047 3156 4413 3164
rect 27 3136 1033 3144
rect 1187 3136 1233 3144
rect 1347 3136 1613 3144
rect 1847 3136 2033 3144
rect 2347 3136 2593 3144
rect 2607 3136 2853 3144
rect 3287 3136 3473 3144
rect 3587 3136 3613 3144
rect 3947 3136 3973 3144
rect 4287 3136 5233 3144
rect 587 3116 1124 3124
rect 867 3096 1073 3104
rect 1116 3104 1124 3116
rect 1147 3116 1293 3124
rect 1407 3116 1533 3124
rect 2187 3116 2253 3124
rect 2367 3116 2433 3124
rect 2527 3116 2573 3124
rect 2707 3116 2753 3124
rect 3047 3116 3213 3124
rect 3347 3116 3433 3124
rect 3707 3116 4073 3124
rect 4187 3116 4253 3124
rect 4267 3116 4453 3124
rect 1116 3096 1593 3104
rect 2147 3096 2513 3104
rect 2647 3096 4193 3104
rect 4207 3096 4333 3104
rect 4367 3096 4433 3104
rect 4447 3096 4713 3104
rect 407 3076 664 3084
rect 367 3056 573 3064
rect 587 3056 633 3064
rect 167 3036 253 3044
rect 307 3036 473 3044
rect 547 3036 613 3044
rect 656 3027 664 3076
rect 1027 3076 1153 3084
rect 1507 3076 1733 3084
rect 1747 3076 1933 3084
rect 2047 3076 2113 3084
rect 2127 3076 2633 3084
rect 2687 3076 2773 3084
rect 2787 3076 2873 3084
rect 2887 3076 2933 3084
rect 3167 3076 3273 3084
rect 3287 3076 3393 3084
rect 3887 3076 4213 3084
rect 687 3056 1173 3064
rect 1287 3056 1313 3064
rect 1527 3056 1573 3064
rect 1587 3056 1673 3064
rect 1987 3056 2073 3064
rect 2087 3056 2353 3064
rect 2487 3056 2553 3064
rect 2587 3056 2953 3064
rect 716 3036 773 3044
rect -24 3016 13 3024
rect 327 3016 513 3024
rect 567 3016 653 3024
rect 127 2996 213 3004
rect 267 2996 413 3004
rect 716 3004 724 3036
rect 827 3036 944 3044
rect 936 3027 944 3036
rect 967 3036 1293 3044
rect 1336 3036 1633 3044
rect 1336 3027 1344 3036
rect 1847 3036 1924 3044
rect 1916 3027 1924 3036
rect 2027 3036 2233 3044
rect 2416 3044 2424 3053
rect 2416 3036 2653 3044
rect 747 3016 753 3024
rect 767 3016 793 3024
rect 987 3016 1033 3024
rect 1547 3016 1653 3024
rect 1727 3016 1773 3024
rect 1827 3016 1873 3024
rect 2127 3016 2253 3024
rect 667 2996 724 3004
rect 836 3004 844 3013
rect 807 2996 844 3004
rect 1096 2987 1104 3013
rect 1167 2996 1413 3004
rect 1427 2996 1473 3004
rect 1707 2996 1733 3004
rect 2276 3004 2284 3033
rect 2416 3027 2424 3036
rect 2367 3016 2393 3024
rect 2456 3016 2533 3024
rect 2456 3004 2464 3016
rect 2696 3007 2704 3056
rect 2987 3056 3164 3064
rect 2787 3036 2844 3044
rect 2736 3024 2744 3033
rect 2836 3024 2844 3036
rect 2867 3036 2973 3044
rect 3087 3036 3133 3044
rect 3156 3044 3164 3056
rect 3267 3056 3653 3064
rect 3767 3056 3833 3064
rect 3847 3056 3993 3064
rect 4107 3056 4293 3064
rect 4367 3056 4393 3064
rect 4727 3056 5113 3064
rect 5187 3056 5264 3064
rect 3156 3036 3373 3044
rect 3507 3036 3544 3044
rect 2736 3016 2784 3024
rect 2836 3016 2873 3024
rect 2167 2996 2464 3004
rect 2487 2996 2673 3004
rect 2776 3004 2784 3016
rect 3536 3024 3544 3036
rect 3567 3036 3633 3044
rect 3827 3036 3873 3044
rect 3907 3036 3933 3044
rect 4007 3036 4033 3044
rect 3407 3016 3524 3024
rect 3536 3016 3773 3024
rect 3516 3007 3524 3016
rect 4056 3024 4064 3053
rect 5256 3047 5264 3056
rect 5367 3056 5533 3064
rect 4227 3036 4433 3044
rect 4447 3036 4473 3044
rect 4707 3036 4753 3044
rect 4787 3036 4993 3044
rect 5047 3036 5133 3044
rect 5527 3036 5673 3044
rect 3847 3016 4064 3024
rect 4156 3024 4164 3033
rect 4156 3016 4533 3024
rect 4616 3007 4624 3033
rect 4647 3016 4893 3024
rect 5207 3016 5613 3024
rect 2776 2996 3073 3004
rect 3087 2996 3233 3004
rect 3407 2996 3453 3004
rect 3547 2996 3673 3004
rect 3687 2996 3893 3004
rect 4207 2996 4353 3004
rect 4367 2996 4373 3004
rect 4827 2996 4873 3004
rect 5027 2996 5113 3004
rect 87 2976 113 2984
rect 227 2976 373 2984
rect 767 2976 1073 2984
rect 1567 2976 1693 2984
rect 1707 2976 1973 2984
rect 2727 2976 3113 2984
rect 3887 2976 3953 2984
rect 3967 2976 4113 2984
rect 4127 2976 4233 2984
rect 4927 2976 4973 2984
rect 4987 2976 5173 2984
rect 667 2956 1113 2964
rect 1127 2956 1273 2964
rect 1507 2956 1653 2964
rect 2207 2956 2713 2964
rect 2907 2956 3433 2964
rect 3676 2956 4793 2964
rect 607 2936 713 2944
rect 727 2936 1153 2944
rect 1987 2936 3293 2944
rect 3676 2944 3684 2956
rect 3387 2936 3684 2944
rect 3716 2936 3813 2944
rect 1047 2916 1393 2924
rect 2247 2916 2433 2924
rect 2447 2916 2593 2924
rect 2987 2916 3133 2924
rect 3716 2924 3724 2936
rect 4427 2936 4733 2944
rect 3176 2916 3724 2924
rect 487 2896 2133 2904
rect 3176 2904 3184 2916
rect 5467 2916 5493 2924
rect 5587 2916 5733 2924
rect 2207 2896 3184 2904
rect 3847 2896 4013 2904
rect 1627 2876 2853 2884
rect 2867 2876 2893 2884
rect 3147 2876 4013 2884
rect 1927 2856 2033 2864
rect 2787 2856 2873 2864
rect 1167 2836 2953 2844
rect 2967 2836 3273 2844
rect 3307 2836 3713 2844
rect 3727 2836 4453 2844
rect 5447 2836 5493 2844
rect 507 2816 853 2824
rect 1307 2816 2053 2824
rect 2127 2816 2173 2824
rect 2587 2816 3033 2824
rect 3127 2816 3853 2824
rect 3867 2816 3873 2824
rect 4267 2816 4613 2824
rect 87 2796 253 2804
rect 787 2796 813 2804
rect 827 2796 893 2804
rect 1947 2796 1993 2804
rect 2187 2796 2313 2804
rect 2447 2796 2753 2804
rect 2847 2796 2913 2804
rect 3187 2796 3253 2804
rect 3487 2796 3513 2804
rect 3667 2796 3733 2804
rect 3947 2796 3973 2804
rect 4007 2796 4293 2804
rect 76 2776 113 2784
rect 76 2744 84 2776
rect 316 2776 373 2784
rect 316 2764 324 2776
rect 627 2776 713 2784
rect 727 2776 793 2784
rect 807 2776 893 2784
rect 947 2776 1073 2784
rect 1327 2776 2013 2784
rect 2227 2776 2373 2784
rect 2387 2776 2453 2784
rect 2647 2776 2673 2784
rect 2767 2776 2993 2784
rect 3007 2776 3033 2784
rect 3087 2776 3113 2784
rect 3167 2776 3213 2784
rect 3236 2776 3313 2784
rect 107 2756 324 2764
rect 347 2756 413 2764
rect 467 2756 533 2764
rect 607 2756 653 2764
rect 847 2756 933 2764
rect 1287 2756 1333 2764
rect 1347 2756 1373 2764
rect 1427 2756 1473 2764
rect 1487 2756 1513 2764
rect 1636 2756 1813 2764
rect 1636 2747 1644 2756
rect 1827 2756 1953 2764
rect 2196 2764 2204 2773
rect 2196 2756 2224 2764
rect 2216 2747 2224 2756
rect 2367 2756 2413 2764
rect 2427 2756 2653 2764
rect 2816 2756 2833 2764
rect 76 2736 93 2744
rect 127 2736 153 2744
rect 227 2736 493 2744
rect 567 2736 573 2744
rect 587 2736 673 2744
rect 747 2736 773 2744
rect 1007 2736 1313 2744
rect 1407 2736 1493 2744
rect 1567 2736 1633 2744
rect 1656 2736 1773 2744
rect 207 2716 393 2724
rect 487 2716 753 2724
rect 907 2716 953 2724
rect 1656 2724 1664 2736
rect 1967 2736 1993 2744
rect 2167 2736 2193 2744
rect 2467 2736 2693 2744
rect 1347 2716 1664 2724
rect 1687 2716 1833 2724
rect 2307 2716 2653 2724
rect 2816 2707 2824 2756
rect 3236 2764 3244 2776
rect 3387 2776 3413 2784
rect 3447 2776 3693 2784
rect 3827 2776 3993 2784
rect 4027 2776 4153 2784
rect 4167 2776 4173 2784
rect 4227 2776 4253 2784
rect 4967 2776 5133 2784
rect 5187 2776 5864 2784
rect 3036 2756 3244 2764
rect 3036 2747 3044 2756
rect 3727 2756 3753 2764
rect 3987 2756 4093 2764
rect 4107 2756 4193 2764
rect 4247 2756 4413 2764
rect 2847 2736 2913 2744
rect 3107 2736 3133 2744
rect 3247 2736 3313 2744
rect 3336 2744 3344 2753
rect 4596 2747 4604 2773
rect 4987 2756 5013 2764
rect 5067 2756 5153 2764
rect 5176 2756 5313 2764
rect 5176 2747 5184 2756
rect 3336 2736 3433 2744
rect 3527 2736 3593 2744
rect 3627 2736 3673 2744
rect 3687 2736 3733 2744
rect 3787 2736 4253 2744
rect 4707 2736 4773 2744
rect 4967 2736 4993 2744
rect 5327 2736 5353 2744
rect 5487 2736 5533 2744
rect 5636 2744 5644 2753
rect 5636 2736 5673 2744
rect 2887 2716 2913 2724
rect 2927 2716 2993 2724
rect 3267 2716 3344 2724
rect 447 2696 633 2704
rect 647 2696 733 2704
rect 747 2696 933 2704
rect 1307 2696 1653 2704
rect 1767 2696 1793 2704
rect 2267 2696 2313 2704
rect 2327 2696 2473 2704
rect 2507 2696 2733 2704
rect 3336 2704 3344 2716
rect 3367 2716 3413 2724
rect 3427 2716 3493 2724
rect 3507 2716 3573 2724
rect 3687 2716 4073 2724
rect 4127 2716 4233 2724
rect 4407 2716 4533 2724
rect 4547 2716 4913 2724
rect 5007 2716 5613 2724
rect 3336 2696 3453 2704
rect 3607 2696 3793 2704
rect 3927 2696 4053 2704
rect 4107 2696 4133 2704
rect 5227 2696 5353 2704
rect 5547 2696 5653 2704
rect 547 2676 673 2684
rect 727 2676 873 2684
rect 1207 2676 2933 2684
rect 3067 2676 3293 2684
rect 3327 2676 3393 2684
rect 3487 2676 3553 2684
rect 3567 2676 3633 2684
rect 3707 2676 3993 2684
rect 4567 2676 4813 2684
rect 4827 2676 5053 2684
rect 5067 2676 5193 2684
rect 5207 2676 5433 2684
rect 5447 2676 5613 2684
rect 187 2656 273 2664
rect 287 2656 353 2664
rect 367 2656 633 2664
rect 1247 2656 1353 2664
rect 1367 2656 1593 2664
rect 1607 2656 1684 2664
rect 1587 2636 1653 2644
rect 1676 2644 1684 2656
rect 1787 2656 1913 2664
rect 2107 2656 3173 2664
rect 3347 2656 3373 2664
rect 3487 2656 3533 2664
rect 3587 2656 3884 2664
rect 1676 2636 3833 2644
rect 3876 2644 3884 2656
rect 3987 2656 4513 2664
rect 3876 2636 3953 2644
rect 1587 2616 1913 2624
rect 1927 2616 2513 2624
rect 2527 2616 3833 2624
rect 3847 2616 4573 2624
rect 167 2596 373 2604
rect 807 2596 993 2604
rect 1187 2596 1644 2604
rect 247 2576 473 2584
rect 487 2576 533 2584
rect 667 2576 753 2584
rect 767 2576 873 2584
rect 1107 2576 1173 2584
rect 1636 2584 1644 2596
rect 1667 2596 1693 2604
rect 1867 2596 1933 2604
rect 2207 2596 2313 2604
rect 2327 2596 2413 2604
rect 2587 2596 2613 2604
rect 2647 2596 2973 2604
rect 3007 2596 3193 2604
rect 3247 2596 4633 2604
rect 1636 2576 1973 2584
rect 2067 2576 2273 2584
rect 2367 2576 2553 2584
rect 2727 2576 2744 2584
rect 316 2556 393 2564
rect 187 2536 293 2544
rect 316 2544 324 2556
rect 656 2556 673 2564
rect 307 2536 324 2544
rect 347 2536 373 2544
rect 387 2536 433 2544
rect 656 2544 664 2556
rect 827 2556 973 2564
rect 996 2556 1093 2564
rect 567 2536 664 2544
rect 747 2536 773 2544
rect 887 2536 913 2544
rect 996 2544 1004 2556
rect 1427 2556 1693 2564
rect 1827 2556 1873 2564
rect 2147 2556 2233 2564
rect 2387 2556 2433 2564
rect 2627 2556 2673 2564
rect 2696 2556 2713 2564
rect 947 2536 1004 2544
rect 1127 2536 1193 2544
rect 1247 2536 1413 2544
rect 1547 2536 1613 2544
rect 1767 2536 1793 2544
rect 127 2516 173 2524
rect 287 2516 353 2524
rect 367 2516 413 2524
rect 987 2516 1033 2524
rect 1287 2516 1353 2524
rect 1527 2516 1553 2524
rect 1647 2516 1993 2524
rect 2016 2524 2024 2553
rect 2047 2536 2093 2544
rect 2127 2536 2144 2544
rect 2016 2516 2113 2524
rect 2136 2524 2144 2536
rect 2167 2536 2333 2544
rect 2507 2536 2593 2544
rect 2696 2544 2704 2556
rect 2736 2544 2744 2576
rect 2787 2576 3713 2584
rect 3767 2576 3813 2584
rect 3867 2576 3913 2584
rect 2847 2556 2884 2564
rect 2876 2547 2884 2556
rect 3107 2556 3153 2564
rect 3207 2556 3273 2564
rect 3387 2556 3473 2564
rect 3667 2556 3744 2564
rect 2616 2536 2704 2544
rect 2716 2536 2744 2544
rect 2136 2516 2164 2524
rect 2156 2507 2164 2516
rect 2187 2516 2293 2524
rect 2367 2516 2393 2524
rect 2447 2516 2473 2524
rect 2616 2524 2624 2536
rect 2716 2527 2724 2536
rect 2827 2536 2853 2544
rect 2947 2536 2973 2544
rect 3047 2536 3264 2544
rect 3256 2527 3264 2536
rect 3736 2527 3744 2556
rect 3807 2536 3853 2544
rect 3896 2544 3904 2553
rect 3896 2536 3913 2544
rect 4087 2536 4253 2544
rect 4267 2536 5233 2544
rect 5387 2536 5453 2544
rect 5467 2536 5493 2544
rect 5607 2536 5713 2544
rect 2507 2516 2624 2524
rect 3167 2516 3213 2524
rect 3287 2516 3353 2524
rect 3447 2516 3613 2524
rect 3627 2516 3704 2524
rect 1227 2496 1333 2504
rect 1347 2496 1473 2504
rect 1547 2496 1573 2504
rect 1727 2496 1793 2504
rect 2447 2496 2453 2504
rect 2467 2496 2753 2504
rect 3187 2496 3213 2504
rect 3236 2496 3353 2504
rect 1567 2476 1733 2484
rect 1747 2476 1764 2484
rect 1807 2476 1833 2484
rect 1856 2476 1893 2484
rect 1507 2456 1693 2464
rect 1856 2464 1864 2476
rect 1907 2476 2253 2484
rect 2347 2476 2493 2484
rect 2607 2476 2693 2484
rect 3236 2484 3244 2496
rect 3396 2504 3404 2513
rect 3396 2496 3513 2504
rect 3527 2496 3673 2504
rect 3696 2504 3704 2516
rect 3767 2516 3793 2524
rect 3867 2516 4033 2524
rect 3696 2496 3813 2504
rect 3947 2496 4453 2504
rect 3207 2476 3244 2484
rect 3347 2476 3473 2484
rect 3587 2476 3653 2484
rect 3787 2476 4013 2484
rect 4467 2476 5193 2484
rect 1747 2456 1864 2464
rect 1887 2456 2213 2464
rect 2247 2456 3073 2464
rect 3307 2456 3433 2464
rect 4527 2456 4833 2464
rect 167 2436 253 2444
rect 767 2436 893 2444
rect 1207 2436 1873 2444
rect 2076 2436 2773 2444
rect 2076 2424 2084 2436
rect 3176 2436 3393 2444
rect 1007 2416 2084 2424
rect 2107 2416 2553 2424
rect 3176 2424 3184 2436
rect 3427 2436 3713 2444
rect 4327 2436 4413 2444
rect 4427 2436 4473 2444
rect 4987 2436 5133 2444
rect 3027 2416 3184 2424
rect 3207 2416 3744 2424
rect 1107 2396 2833 2404
rect 3267 2396 3673 2404
rect 3736 2404 3744 2416
rect 3827 2416 5413 2424
rect 3736 2396 4093 2404
rect 4107 2396 4413 2404
rect 4427 2396 4693 2404
rect 4707 2396 4793 2404
rect 1467 2376 1973 2384
rect 2187 2376 2373 2384
rect 3107 2376 3633 2384
rect 3667 2376 3693 2384
rect 4627 2376 5413 2384
rect 5427 2376 5493 2384
rect 1647 2356 1684 2364
rect 1407 2336 1653 2344
rect 1676 2344 1684 2356
rect 1767 2356 2133 2364
rect 2527 2356 3193 2364
rect 3247 2356 3333 2364
rect 3387 2356 3453 2364
rect 3767 2356 3993 2364
rect 4687 2356 4853 2364
rect 4867 2356 5273 2364
rect 1676 2336 1713 2344
rect 1727 2336 1833 2344
rect 2127 2336 3173 2344
rect 3207 2336 3853 2344
rect 3967 2336 4253 2344
rect 4867 2336 5073 2344
rect 5327 2336 5633 2344
rect 307 2316 353 2324
rect 1607 2316 2053 2324
rect 2167 2316 2193 2324
rect 2987 2316 3044 2324
rect -24 2284 -16 2304
rect 87 2296 224 2304
rect 216 2287 224 2296
rect 247 2296 313 2304
rect 687 2296 893 2304
rect 907 2296 1013 2304
rect 1127 2296 1253 2304
rect 1347 2296 1413 2304
rect 1447 2296 1473 2304
rect 1727 2296 1864 2304
rect 1856 2287 1864 2296
rect 1887 2296 1913 2304
rect 1927 2296 2013 2304
rect 2147 2296 2653 2304
rect 2807 2296 3013 2304
rect 3036 2304 3044 2316
rect 3067 2316 3473 2324
rect 4387 2316 4433 2324
rect 4447 2316 4553 2324
rect 4647 2316 4893 2324
rect 5387 2316 5553 2324
rect 3036 2296 3273 2304
rect 3327 2296 3373 2304
rect 3407 2296 3573 2304
rect 3716 2296 3793 2304
rect -24 2276 93 2284
rect 236 2276 333 2284
rect -24 2256 73 2264
rect 236 2264 244 2276
rect 427 2276 453 2284
rect 827 2276 853 2284
rect 1287 2276 1453 2284
rect 1527 2276 1553 2284
rect 1567 2276 1713 2284
rect 1887 2276 2073 2284
rect 2467 2276 2533 2284
rect 2787 2276 2804 2284
rect 167 2256 244 2264
rect 267 2256 293 2264
rect 307 2256 313 2264
rect 636 2264 644 2273
rect 447 2256 644 2264
rect 967 2256 1153 2264
rect 1507 2256 1693 2264
rect 1736 2247 1744 2273
rect 1807 2256 1893 2264
rect 1927 2256 2033 2264
rect 2047 2256 2113 2264
rect 2647 2256 2773 2264
rect 2796 2264 2804 2276
rect 2847 2276 3033 2284
rect 3267 2276 3293 2284
rect 3307 2276 3413 2284
rect 3716 2284 3724 2296
rect 3847 2296 4013 2304
rect 4487 2296 4733 2304
rect 4907 2296 4933 2304
rect 5247 2296 5273 2304
rect 5467 2296 5513 2304
rect 5527 2296 5713 2304
rect 3676 2276 3724 2284
rect 3676 2267 3684 2276
rect 3747 2276 3893 2284
rect 4287 2276 4353 2284
rect 4827 2276 4913 2284
rect 4927 2276 5053 2284
rect 5107 2276 5133 2284
rect 5567 2276 5573 2284
rect 5587 2276 5664 2284
rect 2796 2256 2893 2264
rect 3047 2256 3193 2264
rect 3227 2256 3273 2264
rect 3507 2256 3533 2264
rect 3587 2256 3633 2264
rect 3707 2256 4164 2264
rect 4156 2247 4164 2256
rect 4187 2256 4393 2264
rect 4596 2247 4604 2273
rect 5656 2267 5664 2276
rect 5707 2276 5733 2284
rect 4627 2256 4713 2264
rect 4887 2256 4973 2264
rect 5127 2256 5213 2264
rect 5407 2256 5453 2264
rect 387 2236 473 2244
rect 507 2236 533 2244
rect 547 2236 653 2244
rect 1047 2236 1073 2244
rect 1307 2236 1433 2244
rect 1447 2236 1573 2244
rect 1767 2236 2173 2244
rect 2276 2236 2333 2244
rect 467 2216 513 2224
rect 587 2216 633 2224
rect 1067 2216 1093 2224
rect 1187 2216 1293 2224
rect 1427 2216 1513 2224
rect 1627 2216 1753 2224
rect 1796 2216 1813 2224
rect 347 2196 593 2204
rect 627 2196 773 2204
rect 1796 2204 1804 2216
rect 2276 2224 2284 2236
rect 2727 2236 2913 2244
rect 2927 2236 3113 2244
rect 3167 2236 3193 2244
rect 3507 2236 3653 2244
rect 3787 2236 3833 2244
rect 4847 2236 4933 2244
rect 5147 2236 5393 2244
rect 5527 2236 5633 2244
rect 5647 2236 5713 2244
rect 2107 2216 2284 2224
rect 2347 2216 2593 2224
rect 2727 2216 2853 2224
rect 2947 2216 3313 2224
rect 3327 2216 3393 2224
rect 3667 2216 4373 2224
rect 1727 2196 1804 2204
rect 1827 2196 1993 2204
rect 2787 2196 3513 2204
rect 3527 2196 3793 2204
rect 4547 2196 4573 2204
rect 4587 2196 5033 2204
rect 5227 2196 5353 2204
rect 5687 2196 5733 2204
rect 427 2176 473 2184
rect 1847 2176 1893 2184
rect 2287 2176 2513 2184
rect 2567 2176 3133 2184
rect 3267 2176 3333 2184
rect 3367 2176 3393 2184
rect 3427 2176 3593 2184
rect 3787 2176 3813 2184
rect 4727 2176 4893 2184
rect 5047 2176 5733 2184
rect 127 2156 1873 2164
rect 2167 2156 2233 2164
rect 2247 2156 2433 2164
rect 2447 2156 3433 2164
rect 3447 2156 3953 2164
rect 4047 2156 4633 2164
rect 5007 2156 5533 2164
rect 587 2136 913 2144
rect 1487 2136 1593 2144
rect 2436 2136 3033 2144
rect 87 2116 793 2124
rect 927 2116 1353 2124
rect 1587 2116 1773 2124
rect 1867 2116 1933 2124
rect 2436 2124 2444 2136
rect 3456 2136 4513 2144
rect 1987 2116 2444 2124
rect 2627 2116 2893 2124
rect 2967 2116 3293 2124
rect 3456 2124 3464 2136
rect 4967 2136 5053 2144
rect 5547 2136 5753 2144
rect 5767 2136 5813 2144
rect 3327 2116 3464 2124
rect 3487 2116 4053 2124
rect 5027 2116 5073 2124
rect 5107 2116 5113 2124
rect 5127 2116 5153 2124
rect 5247 2116 5433 2124
rect 5696 2116 5764 2124
rect 207 2096 273 2104
rect 307 2096 373 2104
rect 807 2096 893 2104
rect 1287 2096 1393 2104
rect 1527 2096 1693 2104
rect 1707 2096 1773 2104
rect 1787 2096 1893 2104
rect 2427 2096 2753 2104
rect 2867 2096 2913 2104
rect 3187 2096 3273 2104
rect 3287 2096 3344 2104
rect 427 2076 613 2084
rect 687 2076 753 2084
rect 847 2076 1113 2084
rect 1147 2076 1213 2084
rect 1267 2076 1393 2084
rect 1407 2076 1473 2084
rect 1496 2076 1653 2084
rect 1496 2067 1504 2076
rect 1687 2076 1933 2084
rect 2007 2076 2093 2084
rect 2207 2076 2884 2084
rect 2876 2067 2884 2076
rect 3227 2076 3253 2084
rect 3336 2084 3344 2096
rect 3367 2096 3533 2104
rect 3587 2096 3673 2104
rect 4087 2096 4253 2104
rect 4467 2096 4513 2104
rect 4707 2096 4773 2104
rect 4827 2096 5153 2104
rect 5207 2096 5273 2104
rect 5387 2096 5433 2104
rect 5636 2096 5673 2104
rect 3336 2076 3453 2084
rect 3467 2076 3524 2084
rect 3516 2067 3524 2076
rect 3647 2076 3793 2084
rect 3807 2076 3833 2084
rect 3987 2076 4013 2084
rect 4107 2076 4133 2084
rect 4147 2076 4213 2084
rect 4387 2076 4473 2084
rect 4496 2076 4553 2084
rect 4496 2067 4504 2076
rect 4887 2076 4913 2084
rect 4936 2076 5013 2084
rect 4936 2067 4944 2076
rect 5176 2084 5184 2093
rect 5156 2076 5184 2084
rect 5156 2067 5164 2076
rect 5267 2076 5353 2084
rect 5636 2067 5644 2096
rect 407 2056 473 2064
rect 827 2056 913 2064
rect 1007 2056 1073 2064
rect 1087 2056 1193 2064
rect 1247 2056 1273 2064
rect 1287 2056 1373 2064
rect 1547 2056 1633 2064
rect 1687 2056 1873 2064
rect 1927 2056 2053 2064
rect 2087 2056 2113 2064
rect 2487 2056 2613 2064
rect 2927 2056 3033 2064
rect 3247 2056 3273 2064
rect 3567 2056 3713 2064
rect 3847 2056 3993 2064
rect 4007 2056 4013 2064
rect 4207 2056 4253 2064
rect 4407 2056 4433 2064
rect 4547 2056 4633 2064
rect 4767 2056 4893 2064
rect 5187 2056 5313 2064
rect 5527 2056 5544 2064
rect 207 2036 233 2044
rect 256 2024 264 2053
rect 296 2044 304 2053
rect 296 2036 513 2044
rect 787 2036 853 2044
rect 907 2036 1053 2044
rect 1667 2036 1693 2044
rect 1767 2036 2073 2044
rect 2307 2036 3184 2044
rect 256 2016 293 2024
rect 307 2016 353 2024
rect 427 2016 713 2024
rect 827 2016 933 2024
rect 1096 2024 1104 2033
rect 967 2016 1613 2024
rect 1687 2016 1833 2024
rect 1856 2016 2353 2024
rect 1856 2004 1864 2016
rect 2847 2016 3053 2024
rect 3176 2024 3184 2036
rect 3207 2036 3313 2044
rect 3347 2036 3553 2044
rect 3627 2036 3813 2044
rect 3827 2036 3933 2044
rect 4067 2036 4113 2044
rect 4627 2036 4733 2044
rect 4747 2036 4853 2044
rect 5087 2036 5193 2044
rect 5487 2036 5513 2044
rect 5536 2044 5544 2056
rect 5696 2047 5704 2116
rect 5716 2096 5733 2104
rect 5716 2067 5724 2096
rect 5756 2084 5764 2116
rect 5747 2076 5764 2084
rect 5536 2036 5673 2044
rect 5747 2036 5773 2044
rect 3176 2016 3593 2024
rect 3607 2016 3653 2024
rect 3787 2016 4273 2024
rect 4627 2016 4713 2024
rect 4767 2016 4813 2024
rect 5027 2016 5233 2024
rect 5427 2016 5473 2024
rect 5487 2016 5713 2024
rect 127 1996 1864 2004
rect 2307 1996 2373 2004
rect 2967 1996 3033 2004
rect 3067 1996 3673 2004
rect 3687 1996 3913 2004
rect 3947 1996 4653 2004
rect 1487 1976 1713 1984
rect 2027 1976 3253 1984
rect 3467 1976 3713 1984
rect 4307 1976 5693 1984
rect 287 1956 333 1964
rect 1847 1956 2253 1964
rect 2627 1956 2773 1964
rect 2787 1956 3073 1964
rect 3087 1956 4293 1964
rect 387 1936 653 1944
rect 1407 1936 1573 1944
rect 1767 1936 1973 1944
rect 2067 1936 2333 1944
rect 2607 1936 2713 1944
rect 3027 1936 3173 1944
rect 3647 1936 4093 1944
rect 4107 1936 4244 1944
rect 1927 1916 3493 1924
rect 3547 1916 4153 1924
rect 4236 1924 4244 1936
rect 4236 1916 4313 1924
rect 4327 1916 4413 1924
rect 5087 1916 5253 1924
rect 2427 1896 2553 1904
rect 2707 1896 3613 1904
rect 3707 1896 4133 1904
rect 4227 1896 5293 1904
rect 407 1876 513 1884
rect 1027 1876 1933 1884
rect 1987 1876 2793 1884
rect 2827 1876 3153 1884
rect 3807 1876 4033 1884
rect 4067 1876 4173 1884
rect 4187 1876 4713 1884
rect 4807 1876 5493 1884
rect 227 1856 713 1864
rect 1707 1856 1853 1864
rect 2827 1856 2993 1864
rect 3507 1856 4213 1864
rect 4727 1856 4893 1864
rect 4907 1856 5253 1864
rect 5267 1856 5333 1864
rect 5367 1856 5393 1864
rect 207 1836 333 1844
rect 347 1836 493 1844
rect 727 1836 1133 1844
rect 1247 1836 2113 1844
rect 2227 1836 2613 1844
rect 2767 1836 3373 1844
rect 3387 1836 3613 1844
rect 3867 1836 4013 1844
rect 4127 1836 4173 1844
rect 4187 1836 4273 1844
rect 4367 1836 4453 1844
rect 4507 1836 4553 1844
rect 4687 1836 4853 1844
rect 4987 1836 5033 1844
rect 5347 1836 5433 1844
rect 127 1816 213 1824
rect 247 1816 264 1824
rect 107 1796 193 1804
rect 236 1784 244 1793
rect 147 1776 244 1784
rect 127 1756 213 1764
rect 256 1744 264 1816
rect 376 1804 384 1813
rect 356 1796 384 1804
rect 356 1787 364 1796
rect 416 1784 424 1813
rect 387 1776 424 1784
rect 516 1784 524 1833
rect 547 1816 953 1824
rect 1867 1816 1953 1824
rect 1967 1816 2153 1824
rect 2207 1816 2253 1824
rect 2787 1816 2833 1824
rect 2887 1816 3033 1824
rect 3056 1816 3093 1824
rect 567 1796 593 1804
rect 607 1796 833 1804
rect 947 1796 1033 1804
rect 1107 1796 1173 1804
rect 1187 1796 1233 1804
rect 1287 1796 1333 1804
rect 1647 1796 1753 1804
rect 2247 1796 2273 1804
rect 2587 1796 2653 1804
rect 2807 1796 2853 1804
rect 3056 1804 3064 1816
rect 3127 1816 3313 1824
rect 3387 1816 3413 1824
rect 3587 1816 3953 1824
rect 4147 1816 4733 1824
rect 4947 1816 4993 1824
rect 2987 1796 3064 1804
rect 3407 1796 3493 1804
rect 4007 1796 4113 1804
rect 4247 1796 4453 1804
rect 4467 1796 4593 1804
rect 4807 1796 4824 1804
rect 516 1776 553 1784
rect 707 1776 804 1784
rect 427 1756 684 1764
rect 227 1736 264 1744
rect 427 1736 473 1744
rect 676 1744 684 1756
rect 727 1756 773 1764
rect 796 1764 804 1776
rect 827 1776 973 1784
rect 1127 1776 1253 1784
rect 1267 1776 1393 1784
rect 1507 1776 1533 1784
rect 1547 1776 1553 1784
rect 1627 1776 1733 1784
rect 2187 1776 2633 1784
rect 2647 1776 2893 1784
rect 2967 1776 3093 1784
rect 3216 1784 3224 1793
rect 3107 1776 3224 1784
rect 3307 1776 3353 1784
rect 3627 1776 3713 1784
rect 3727 1776 3773 1784
rect 3847 1776 3933 1784
rect 3956 1784 3964 1793
rect 4816 1787 4824 1796
rect 4927 1796 4973 1804
rect 5016 1796 5133 1804
rect 5016 1787 5024 1796
rect 5187 1796 5284 1804
rect 5276 1787 5284 1796
rect 5307 1796 5384 1804
rect 5376 1787 5384 1796
rect 5507 1796 5533 1804
rect 5667 1796 5864 1804
rect 3956 1776 3993 1784
rect 4167 1776 4253 1784
rect 4447 1776 4473 1784
rect 4567 1776 4633 1784
rect 5067 1776 5133 1784
rect 5427 1776 5533 1784
rect 796 1756 993 1764
rect 1047 1756 1133 1764
rect 1147 1756 1193 1764
rect 1447 1756 1513 1764
rect 1527 1756 1773 1764
rect 1787 1756 1833 1764
rect 2467 1756 2553 1764
rect 2707 1756 2753 1764
rect 2827 1756 2993 1764
rect 3047 1756 3113 1764
rect 3407 1756 3633 1764
rect 3667 1756 3813 1764
rect 3827 1756 4333 1764
rect 4707 1756 4753 1764
rect 5007 1756 5053 1764
rect 5067 1756 5093 1764
rect 5327 1756 5353 1764
rect 5367 1756 5413 1764
rect 5427 1756 5593 1764
rect 527 1736 664 1744
rect 676 1736 853 1744
rect 267 1716 353 1724
rect 527 1716 553 1724
rect 656 1724 664 1736
rect 967 1736 1053 1744
rect 1367 1736 1413 1744
rect 1507 1736 1813 1744
rect 1947 1736 2573 1744
rect 2727 1736 2913 1744
rect 3087 1736 3293 1744
rect 3487 1736 3653 1744
rect 3787 1736 3953 1744
rect 4347 1736 4533 1744
rect 4547 1736 4773 1744
rect 4787 1736 4913 1744
rect 4927 1736 5233 1744
rect 5247 1736 5433 1744
rect 5447 1736 5573 1744
rect 656 1716 1313 1724
rect 1387 1716 1873 1724
rect 2607 1716 2813 1724
rect 2927 1716 3173 1724
rect 3267 1716 3633 1724
rect 3647 1716 3693 1724
rect 4336 1716 4553 1724
rect 4336 1707 4344 1716
rect 5187 1716 5233 1724
rect 5247 1716 5373 1724
rect 5407 1716 5453 1724
rect 147 1696 733 1704
rect 1867 1696 2233 1704
rect 2407 1696 2473 1704
rect 3427 1696 3473 1704
rect 3487 1696 3893 1704
rect 3987 1696 4093 1704
rect 4467 1696 4553 1704
rect 4627 1696 4813 1704
rect 5256 1696 5433 1704
rect 207 1676 293 1684
rect 1147 1676 1313 1684
rect 1447 1676 1593 1684
rect 1807 1676 1913 1684
rect 1936 1676 1993 1684
rect 947 1656 1093 1664
rect 1936 1664 1944 1676
rect 2527 1676 3193 1684
rect 3276 1676 3313 1684
rect 1107 1656 1944 1664
rect 2907 1656 3213 1664
rect 3247 1656 3264 1664
rect 87 1636 573 1644
rect 587 1636 613 1644
rect 1307 1636 2253 1644
rect 2507 1636 2853 1644
rect 3007 1636 3233 1644
rect 327 1616 373 1624
rect 567 1616 693 1624
rect 747 1616 753 1624
rect 767 1616 893 1624
rect 987 1616 1293 1624
rect 1347 1616 1453 1624
rect 1587 1616 1633 1624
rect 1747 1616 1833 1624
rect 2047 1616 2333 1624
rect 2547 1616 2713 1624
rect 2807 1616 3033 1624
rect 3047 1616 3053 1624
rect 287 1596 384 1604
rect 376 1587 384 1596
rect 887 1596 1033 1604
rect 1167 1596 1373 1604
rect 1607 1596 1633 1604
rect 2307 1596 2413 1604
rect 2607 1596 2724 1604
rect 47 1576 113 1584
rect 287 1576 353 1584
rect 507 1576 533 1584
rect 787 1576 853 1584
rect 927 1576 973 1584
rect 1047 1576 1173 1584
rect 1567 1576 1653 1584
rect 2136 1584 2144 1593
rect 2047 1576 2144 1584
rect 2267 1576 2313 1584
rect 2367 1576 2453 1584
rect -24 1556 13 1564
rect 147 1556 213 1564
rect 256 1564 264 1573
rect 2716 1567 2724 1596
rect 3096 1596 3113 1604
rect 2747 1576 2973 1584
rect 256 1556 393 1564
rect 607 1556 633 1564
rect 1207 1556 1253 1564
rect 1267 1556 1313 1564
rect 1487 1556 1773 1564
rect 3096 1564 3104 1596
rect 3127 1576 3233 1584
rect 3096 1556 3124 1564
rect 96 1544 104 1553
rect 3116 1547 3124 1556
rect 96 1536 113 1544
rect 207 1536 233 1544
rect 367 1536 753 1544
rect 2447 1536 2753 1544
rect 2767 1536 2793 1544
rect 2927 1536 2973 1544
rect 87 1516 373 1524
rect 967 1516 1253 1524
rect 2667 1516 2853 1524
rect 3027 1516 3133 1524
rect 27 1496 1393 1504
rect 3256 1487 3264 1656
rect 3276 1487 3284 1676
rect 3567 1676 3673 1684
rect 4087 1676 4233 1684
rect 4787 1676 5013 1684
rect 5256 1684 5264 1696
rect 5207 1676 5264 1684
rect 5287 1676 5333 1684
rect 3747 1656 3913 1664
rect 4007 1656 4293 1664
rect 4367 1656 4833 1664
rect 5087 1656 5193 1664
rect 5207 1656 5253 1664
rect 5307 1656 5473 1664
rect 3767 1636 4073 1644
rect 4096 1636 4793 1644
rect 3567 1616 3593 1624
rect 3687 1616 3753 1624
rect 4096 1624 4104 1636
rect 5127 1636 5373 1644
rect 5587 1636 5753 1644
rect 3987 1616 4104 1624
rect 4467 1616 4473 1624
rect 4547 1616 4613 1624
rect 4807 1616 4853 1624
rect 4887 1616 4933 1624
rect 5027 1616 5364 1624
rect 3547 1596 3593 1604
rect 3676 1596 3713 1604
rect 3676 1584 3684 1596
rect 3847 1596 3873 1604
rect 4007 1596 4013 1604
rect 4027 1596 4124 1604
rect 3667 1576 3684 1584
rect 3707 1576 3733 1584
rect 3787 1576 3893 1584
rect 3447 1556 3473 1564
rect 3627 1556 3673 1564
rect 4116 1564 4124 1596
rect 4147 1596 4253 1604
rect 4347 1596 4493 1604
rect 4507 1596 4573 1604
rect 4667 1596 4753 1604
rect 4856 1596 4893 1604
rect 4287 1576 4433 1584
rect 4447 1576 4553 1584
rect 4567 1576 4633 1584
rect 4776 1584 4784 1593
rect 4647 1576 4784 1584
rect 4856 1567 4864 1596
rect 5287 1596 5333 1604
rect 5356 1587 5364 1616
rect 5647 1616 5713 1624
rect 5487 1596 5533 1604
rect 5667 1596 5793 1604
rect 5327 1576 5344 1584
rect 5336 1567 5344 1576
rect 5456 1576 5573 1584
rect 5456 1567 5464 1576
rect 5627 1576 5793 1584
rect 4116 1556 4153 1564
rect 4747 1556 4833 1564
rect 5087 1556 5173 1564
rect 5347 1556 5433 1564
rect 5507 1556 5553 1564
rect 5567 1556 5593 1564
rect 3487 1536 3513 1544
rect 3547 1536 3593 1544
rect 3747 1536 4593 1544
rect 4607 1536 4813 1544
rect 4827 1536 5033 1544
rect 5207 1536 5253 1544
rect 5407 1536 5453 1544
rect 5627 1536 5673 1544
rect 3527 1516 3853 1524
rect 3867 1516 4113 1524
rect 4787 1516 4873 1524
rect 4887 1516 4993 1524
rect 5127 1516 5213 1524
rect 5327 1516 5773 1524
rect 3447 1496 4733 1504
rect 5427 1496 5773 1504
rect 307 1476 393 1484
rect 2047 1476 2113 1484
rect 3547 1476 4013 1484
rect 4027 1476 4273 1484
rect 4287 1476 4313 1484
rect 4327 1476 4473 1484
rect 5447 1476 5513 1484
rect 327 1456 353 1464
rect 2547 1456 3453 1464
rect 3467 1456 5033 1464
rect 5047 1456 5073 1464
rect 5087 1456 5333 1464
rect 2307 1436 3533 1444
rect 5187 1436 5233 1444
rect 127 1416 313 1424
rect 1387 1416 2593 1424
rect 2607 1416 2733 1424
rect 2747 1416 2933 1424
rect 3807 1416 3833 1424
rect 3967 1416 4753 1424
rect 5107 1416 5233 1424
rect 2567 1396 2613 1404
rect 2847 1396 2873 1404
rect 3127 1396 3293 1404
rect 3667 1396 3693 1404
rect 3707 1396 4353 1404
rect 4827 1396 4853 1404
rect 5587 1396 5653 1404
rect 1707 1376 1753 1384
rect 1767 1376 1793 1384
rect 1807 1376 2073 1384
rect 2147 1376 2233 1384
rect 2927 1376 3033 1384
rect 3467 1376 3493 1384
rect 3747 1376 3773 1384
rect 3787 1376 4173 1384
rect 4547 1376 4853 1384
rect 5147 1376 5213 1384
rect 5547 1376 5653 1384
rect 827 1356 913 1364
rect 927 1356 1013 1364
rect 1716 1356 1733 1364
rect 1716 1347 1724 1356
rect 1747 1356 1984 1364
rect 1976 1347 1984 1356
rect 2647 1356 2853 1364
rect 2867 1356 2913 1364
rect 3007 1356 3053 1364
rect 3207 1356 3913 1364
rect 4087 1356 4133 1364
rect 5147 1356 5253 1364
rect 5267 1356 5553 1364
rect 5707 1356 5753 1364
rect 207 1336 473 1344
rect 516 1336 533 1344
rect 107 1316 193 1324
rect 247 1316 273 1324
rect 407 1316 493 1324
rect 516 1307 524 1336
rect 887 1336 953 1344
rect 967 1336 1193 1344
rect 1467 1336 1673 1344
rect 1887 1336 1933 1344
rect 2027 1336 2193 1344
rect 2247 1336 2293 1344
rect 2387 1336 4493 1344
rect 4507 1336 4653 1344
rect 4667 1336 4673 1344
rect 4727 1336 5093 1344
rect 5107 1336 5273 1344
rect 5287 1336 5313 1344
rect 5407 1336 5493 1344
rect 5607 1336 5633 1344
rect 547 1316 573 1324
rect 587 1316 673 1324
rect 1067 1316 1133 1324
rect 1187 1316 1213 1324
rect 1567 1316 1693 1324
rect 1707 1316 1953 1324
rect 2067 1316 2253 1324
rect 2407 1316 2673 1324
rect 2747 1316 2873 1324
rect 2887 1316 3013 1324
rect 3027 1316 3153 1324
rect 3707 1316 3764 1324
rect 267 1296 433 1304
rect 567 1296 633 1304
rect 647 1296 793 1304
rect 1167 1296 1293 1304
rect 2227 1296 2353 1304
rect 2567 1296 2613 1304
rect 2716 1287 2724 1313
rect 3756 1307 3764 1316
rect 4107 1316 4153 1324
rect 4567 1316 4593 1324
rect 4647 1316 4733 1324
rect 4907 1316 5113 1324
rect 5267 1316 5353 1324
rect 5376 1316 5493 1324
rect 2787 1296 2813 1304
rect 2847 1296 2893 1304
rect 2987 1296 3033 1304
rect 3147 1296 3413 1304
rect 3467 1296 3533 1304
rect 4056 1304 4064 1313
rect 4196 1304 4204 1313
rect 4056 1296 4293 1304
rect 4316 1304 4324 1313
rect 4316 1296 4453 1304
rect 4527 1296 4573 1304
rect 5376 1304 5384 1316
rect 5027 1296 5384 1304
rect 387 1276 553 1284
rect 1267 1276 1313 1284
rect 2007 1276 2093 1284
rect 2107 1276 2313 1284
rect 2347 1276 2453 1284
rect 2467 1276 2533 1284
rect 2787 1276 2853 1284
rect 3047 1276 3273 1284
rect 3327 1276 3453 1284
rect 3687 1276 3733 1284
rect 4027 1276 4173 1284
rect 4287 1276 4333 1284
rect 4587 1276 4693 1284
rect 4807 1276 4893 1284
rect 4907 1276 5013 1284
rect 5227 1276 5633 1284
rect 187 1256 233 1264
rect 327 1256 373 1264
rect 467 1256 513 1264
rect 547 1256 653 1264
rect 2107 1256 2273 1264
rect 2367 1256 3573 1264
rect 3727 1256 3793 1264
rect 4447 1256 4473 1264
rect 4487 1256 4793 1264
rect 5307 1256 5413 1264
rect 127 1236 273 1244
rect 287 1236 473 1244
rect 1807 1236 2373 1244
rect 3207 1236 3373 1244
rect 4227 1236 4993 1244
rect 147 1216 213 1224
rect 227 1216 533 1224
rect 2527 1216 2733 1224
rect 2807 1216 3173 1224
rect 3427 1216 3493 1224
rect 3827 1216 3893 1224
rect 3907 1216 4433 1224
rect 2327 1196 2693 1204
rect 2767 1196 3433 1204
rect 3487 1196 3633 1204
rect 3647 1196 3713 1204
rect 3787 1196 4213 1204
rect 4427 1196 4873 1204
rect 5607 1196 5633 1204
rect 107 1176 433 1184
rect 1567 1176 1613 1184
rect 1627 1176 2013 1184
rect 2087 1176 2493 1184
rect 2727 1176 2813 1184
rect 2827 1176 2953 1184
rect 2967 1176 2993 1184
rect 3007 1176 3213 1184
rect 3507 1176 3593 1184
rect 3607 1176 3673 1184
rect 3807 1176 3853 1184
rect 4267 1176 4373 1184
rect 4667 1176 4693 1184
rect 5147 1176 5473 1184
rect 5607 1176 5673 1184
rect 227 1156 293 1164
rect 667 1156 773 1164
rect 787 1156 933 1164
rect 1147 1156 1433 1164
rect 1527 1156 1633 1164
rect 3167 1156 3373 1164
rect 3567 1156 4353 1164
rect 4407 1156 4493 1164
rect 4507 1156 4533 1164
rect 4547 1156 4713 1164
rect 5347 1156 5373 1164
rect 5687 1156 5753 1164
rect 47 1136 173 1144
rect 447 1136 613 1144
rect 687 1136 893 1144
rect 947 1136 993 1144
rect 1207 1136 1273 1144
rect 1287 1136 1333 1144
rect 1387 1136 1533 1144
rect 1847 1136 2213 1144
rect 2227 1136 2253 1144
rect 2447 1136 2553 1144
rect 2967 1136 3053 1144
rect 3236 1136 3253 1144
rect 176 1116 353 1124
rect 87 1096 153 1104
rect 176 1104 184 1116
rect 407 1116 613 1124
rect 847 1116 1053 1124
rect 1227 1116 2033 1124
rect 2187 1116 2313 1124
rect 2387 1116 2453 1124
rect 2607 1116 2753 1124
rect 2907 1116 2933 1124
rect 3087 1116 3113 1124
rect 3236 1107 3244 1136
rect 3407 1136 3433 1144
rect 3547 1136 3853 1144
rect 4027 1136 4093 1144
rect 4367 1136 4453 1144
rect 4627 1136 4664 1144
rect 3327 1116 3593 1124
rect 3707 1116 3733 1124
rect 3907 1116 3973 1124
rect 4127 1116 4153 1124
rect 4187 1116 4313 1124
rect 4336 1116 4493 1124
rect 4336 1107 4344 1116
rect 4656 1107 4664 1136
rect 4727 1136 4733 1144
rect 4747 1136 4913 1144
rect 4927 1136 4973 1144
rect 5007 1136 5233 1144
rect 5307 1136 5313 1144
rect 5327 1136 5413 1144
rect 5427 1136 5473 1144
rect 5507 1136 5533 1144
rect 5727 1136 5784 1144
rect 4787 1116 4813 1124
rect 5287 1116 5373 1124
rect 5396 1116 5513 1124
rect 5396 1107 5404 1116
rect 5627 1116 5744 1124
rect 167 1096 184 1104
rect 207 1096 273 1104
rect 296 1096 373 1104
rect 296 1084 304 1096
rect 387 1096 493 1104
rect 787 1096 873 1104
rect 1127 1096 1293 1104
rect 1307 1096 1373 1104
rect 1547 1096 1913 1104
rect 2067 1096 2113 1104
rect 2287 1096 2333 1104
rect 2367 1096 2393 1104
rect 2487 1096 2533 1104
rect 2647 1096 2673 1104
rect 2747 1096 2773 1104
rect 3627 1096 3653 1104
rect 3927 1096 3973 1104
rect 4467 1096 4513 1104
rect 4687 1096 4713 1104
rect 5687 1096 5693 1104
rect 5707 1096 5713 1104
rect 5736 1104 5744 1116
rect 5776 1107 5784 1136
rect 5736 1096 5753 1104
rect 87 1076 304 1084
rect 327 1076 453 1084
rect 547 1076 593 1084
rect 647 1076 673 1084
rect 707 1076 893 1084
rect 1036 1084 1044 1093
rect 1036 1076 1253 1084
rect 1267 1076 1413 1084
rect 1467 1076 1753 1084
rect 1887 1076 1933 1084
rect 2016 1084 2024 1093
rect 1967 1076 2153 1084
rect 2207 1076 2613 1084
rect 2627 1076 2973 1084
rect 3107 1076 3153 1084
rect 3576 1084 3584 1093
rect 3576 1076 3593 1084
rect 3607 1076 3693 1084
rect 3807 1076 3833 1084
rect 3887 1076 4413 1084
rect 4707 1076 4753 1084
rect 4787 1076 4813 1084
rect 4867 1076 4913 1084
rect 4927 1076 4953 1084
rect 5587 1076 5653 1084
rect 1267 1056 1493 1064
rect 1867 1056 1893 1064
rect 2087 1056 3133 1064
rect 3287 1056 4053 1064
rect 4067 1056 5013 1064
rect 1307 1036 1353 1044
rect 2427 1036 2513 1044
rect 2887 1036 3333 1044
rect 3667 1036 3753 1044
rect 367 1016 393 1024
rect 427 1016 633 1024
rect 647 1016 673 1024
rect 3447 1016 3913 1024
rect 1827 996 3513 1004
rect 2927 976 3493 984
rect 3507 976 3693 984
rect 487 956 513 964
rect 3516 956 5013 964
rect 3516 944 3524 956
rect 5027 956 5053 964
rect 2987 936 3524 944
rect 3807 936 3853 944
rect 2247 916 2293 924
rect 3267 916 3533 924
rect 3667 916 4213 924
rect 5507 916 5533 924
rect 587 896 613 904
rect 627 896 733 904
rect 2147 896 2213 904
rect 2307 896 2553 904
rect 3827 896 3873 904
rect 3896 896 3993 904
rect 147 876 173 884
rect 887 876 1213 884
rect 1347 876 1364 884
rect 96 856 233 864
rect 96 847 104 856
rect 447 856 553 864
rect 687 856 713 864
rect 727 856 793 864
rect 916 856 1133 864
rect 916 847 924 856
rect 1356 864 1364 876
rect 1447 876 1853 884
rect 2016 876 2273 884
rect 1356 856 1373 864
rect 1427 856 1453 864
rect 1487 856 1553 864
rect 1647 856 1713 864
rect 2016 864 2024 876
rect 2947 876 3113 884
rect 3896 884 3904 896
rect 4007 896 4233 904
rect 5047 896 5133 904
rect 5427 896 5613 904
rect 3127 876 3904 884
rect 4107 876 4133 884
rect 4607 876 4793 884
rect 4887 876 4933 884
rect 5247 876 5313 884
rect 5547 876 5684 884
rect 1907 856 2024 864
rect 2047 856 2053 864
rect 2067 856 2133 864
rect 2527 856 2633 864
rect 2867 856 2893 864
rect 3307 856 3473 864
rect 3727 856 3893 864
rect 4047 856 4113 864
rect 4127 856 4153 864
rect 4627 856 4653 864
rect 4667 856 4773 864
rect 4907 856 5613 864
rect 5627 856 5653 864
rect 5676 864 5684 876
rect 5707 876 5753 884
rect 5676 856 5724 864
rect 147 836 193 844
rect 387 836 513 844
rect 567 836 853 844
rect 967 836 1013 844
rect 1087 836 1133 844
rect 1367 836 1573 844
rect 1787 836 1833 844
rect 1847 836 1913 844
rect 1927 836 1973 844
rect 2587 836 2773 844
rect 3027 836 3053 844
rect 3147 836 3173 844
rect 3427 836 3473 844
rect 3687 836 3733 844
rect 3807 836 3833 844
rect 3927 836 4013 844
rect 4187 836 4313 844
rect 4407 836 4433 844
rect 4527 836 4573 844
rect 4707 836 4733 844
rect 4756 836 4893 844
rect 267 816 313 824
rect 507 816 613 824
rect 827 816 893 824
rect 1196 824 1204 833
rect 1027 816 1204 824
rect 1227 816 1293 824
rect 1747 816 1813 824
rect 1887 816 2013 824
rect 2027 816 2073 824
rect 2167 816 2433 824
rect 2687 816 2733 824
rect 3407 816 3444 824
rect 127 796 213 804
rect 247 796 273 804
rect 347 796 373 804
rect 407 796 533 804
rect 547 796 933 804
rect 1107 796 1233 804
rect 1467 796 1613 804
rect 1787 796 2113 804
rect 2127 796 2313 804
rect 2967 796 2993 804
rect 3127 796 3153 804
rect 3347 796 3413 804
rect 3436 804 3444 816
rect 3527 816 3893 824
rect 4207 816 4253 824
rect 4756 824 4764 836
rect 4907 836 4933 844
rect 4987 836 5073 844
rect 4547 816 4764 824
rect 4967 816 5033 824
rect 3436 796 3533 804
rect 3567 796 3673 804
rect 3687 796 3753 804
rect 3807 796 3993 804
rect 4007 796 4053 804
rect 4147 796 4293 804
rect 4307 796 4413 804
rect 4567 796 4733 804
rect 4787 796 4813 804
rect 5056 804 5064 836
rect 5327 836 5373 844
rect 5396 836 5493 844
rect 5267 816 5313 824
rect 5396 807 5404 836
rect 5587 836 5693 844
rect 5427 816 5473 824
rect 5567 816 5593 824
rect 5716 824 5724 856
rect 5687 816 5724 824
rect 4827 796 5073 804
rect 5127 796 5253 804
rect 5287 796 5333 804
rect 667 776 733 784
rect 747 776 953 784
rect 1767 776 1993 784
rect 2707 776 2813 784
rect 2827 776 3273 784
rect 3447 776 4073 784
rect 4867 776 4913 784
rect 4927 776 5113 784
rect 5307 776 5493 784
rect 687 756 773 764
rect 787 756 1033 764
rect 1987 756 2093 764
rect 2447 756 2653 764
rect 3867 756 4333 764
rect 4347 756 4773 764
rect 1347 736 1953 744
rect 2007 736 4513 744
rect 4527 736 4673 744
rect 5267 736 5433 744
rect 5447 736 5473 744
rect 5487 736 5653 744
rect 147 716 353 724
rect 3807 716 3893 724
rect 5347 716 5673 724
rect 1467 696 1813 704
rect 1867 696 2373 704
rect 3887 696 4033 704
rect 4047 696 4433 704
rect 4867 696 5353 704
rect 5367 696 5373 704
rect 5447 696 5593 704
rect 947 676 1113 684
rect 1127 676 1213 684
rect 1227 676 1533 684
rect 1827 676 2173 684
rect 3567 676 4353 684
rect 4367 676 4593 684
rect 4727 676 4833 684
rect 4847 676 4993 684
rect 5167 676 5213 684
rect 5287 676 5553 684
rect 167 656 273 664
rect 467 656 653 664
rect 987 656 993 664
rect 1007 656 1184 664
rect 127 636 533 644
rect 296 627 304 636
rect 1107 636 1153 644
rect 1176 644 1184 656
rect 1407 656 1513 664
rect 1667 656 1933 664
rect 2007 656 2093 664
rect 2127 656 2253 664
rect 2747 656 2844 664
rect 1176 636 1353 644
rect 1236 627 1244 636
rect 1527 636 1673 644
rect 1727 636 1733 644
rect 1747 636 1993 644
rect 2087 636 2233 644
rect 2247 636 2273 644
rect 2836 627 2844 656
rect 2887 656 3093 664
rect 3107 656 3193 664
rect 3207 656 3373 664
rect 3427 656 3633 664
rect 3827 656 3933 664
rect 4187 656 4213 664
rect 4387 656 4473 664
rect 4667 656 4793 664
rect 4887 656 4913 664
rect 4927 656 4953 664
rect 5107 656 5133 664
rect 5167 656 5453 664
rect 5467 656 5633 664
rect 3047 636 3133 644
rect 3167 636 3513 644
rect 3567 636 3593 644
rect 3687 636 3773 644
rect 4087 636 4204 644
rect 67 616 93 624
rect 107 616 253 624
rect 327 616 393 624
rect 607 616 673 624
rect 696 616 793 624
rect 47 596 73 604
rect 516 604 524 613
rect 427 596 633 604
rect 696 604 704 616
rect 987 616 1013 624
rect 1147 616 1193 624
rect 1427 616 1533 624
rect 1607 616 1653 624
rect 1707 616 1773 624
rect 1867 616 1913 624
rect 1967 616 1993 624
rect 2356 616 2473 624
rect 2356 607 2364 616
rect 2627 616 2733 624
rect 2747 616 2824 624
rect 647 596 704 604
rect 867 596 1073 604
rect 1207 596 1553 604
rect 1727 596 1833 604
rect 1847 596 2053 604
rect 2816 604 2824 616
rect 3007 616 3073 624
rect 3127 616 3173 624
rect 3307 616 3333 624
rect 3347 616 3493 624
rect 3616 624 3624 633
rect 3547 616 3664 624
rect 2816 596 2973 604
rect 3027 596 3233 604
rect 3256 604 3264 613
rect 3256 596 3353 604
rect 87 576 153 584
rect 687 576 773 584
rect 787 576 1313 584
rect 1427 576 1793 584
rect 2187 576 2793 584
rect 2807 576 3093 584
rect 3496 584 3504 613
rect 3656 607 3664 616
rect 3707 616 3793 624
rect 3807 616 3893 624
rect 3916 604 3924 633
rect 4196 627 4204 636
rect 4647 636 4713 644
rect 4787 636 4853 644
rect 5147 636 5273 644
rect 5296 636 5413 644
rect 4007 616 4053 624
rect 4216 607 4224 633
rect 4247 616 4333 624
rect 4407 616 4453 624
rect 4627 616 4653 624
rect 4736 624 4744 633
rect 4676 616 4744 624
rect 3747 596 3924 604
rect 4576 604 4584 613
rect 4676 604 4684 616
rect 4767 616 4793 624
rect 4847 616 4873 624
rect 4236 596 4684 604
rect 4236 584 4244 596
rect 4896 604 4904 633
rect 5296 624 5304 636
rect 5427 636 5533 644
rect 5607 636 5693 644
rect 5267 616 5304 624
rect 5407 616 5473 624
rect 5487 616 5573 624
rect 4827 596 4904 604
rect 5307 596 5333 604
rect 5667 596 5733 604
rect 3496 576 4244 584
rect 1247 556 1373 564
rect 1387 556 1473 564
rect 1847 556 2493 564
rect 3267 556 3353 564
rect 3367 556 4213 564
rect 167 536 453 544
rect 467 536 513 544
rect 1127 536 1153 544
rect 2347 536 2593 544
rect 2607 536 2693 544
rect 2707 536 2973 544
rect 2987 536 3153 544
rect 3927 536 3953 544
rect 5507 536 5673 544
rect 2647 516 2773 524
rect 2787 516 2793 524
rect 3827 516 4013 524
rect 5227 516 5393 524
rect 2087 496 2293 504
rect 4807 496 5513 504
rect 5107 476 5413 484
rect 5427 476 5593 484
rect 2667 456 2913 464
rect 3187 456 3693 464
rect 4507 456 4533 464
rect 5267 456 5353 464
rect 2607 436 3493 444
rect 4127 436 4193 444
rect 5167 436 5613 444
rect 307 416 553 424
rect 1027 416 1633 424
rect 2267 416 2533 424
rect 2847 416 3133 424
rect 3147 416 3313 424
rect 3867 416 3893 424
rect 5147 416 5353 424
rect 747 396 813 404
rect 1487 396 1913 404
rect 2367 396 2633 404
rect 2727 396 3053 404
rect 3227 396 3413 404
rect 3507 396 3573 404
rect 3607 396 3733 404
rect 3807 396 3833 404
rect 4136 396 4153 404
rect 4136 387 4144 396
rect 4187 396 4513 404
rect 5087 396 5293 404
rect 5387 396 5513 404
rect 5527 396 5553 404
rect 5567 396 5633 404
rect 5727 396 5753 404
rect 216 376 413 384
rect 216 367 224 376
rect 556 376 793 384
rect 107 356 213 364
rect 267 356 293 364
rect 467 356 533 364
rect 556 364 564 376
rect 967 376 1033 384
rect 1047 376 1073 384
rect 1116 376 1353 384
rect 547 356 564 364
rect 1007 356 1093 364
rect 1116 364 1124 376
rect 1407 376 1513 384
rect 1527 376 1593 384
rect 1667 376 1693 384
rect 1787 376 1853 384
rect 1867 376 1993 384
rect 2007 376 2553 384
rect 2567 376 2873 384
rect 2887 376 3533 384
rect 3547 376 3673 384
rect 3867 376 3933 384
rect 3947 376 4093 384
rect 4147 376 4413 384
rect 4527 376 4813 384
rect 5027 376 5144 384
rect 5136 367 5144 376
rect 5187 376 5433 384
rect 5627 376 5644 384
rect 1107 356 1124 364
rect 1387 356 1453 364
rect 1627 356 1713 364
rect 2047 356 2133 364
rect 2227 356 2293 364
rect 2307 356 2413 364
rect 2547 356 2733 364
rect 3027 356 3153 364
rect 3187 356 3253 364
rect 3467 356 3633 364
rect 3927 356 3953 364
rect 4027 356 4113 364
rect 4207 356 4244 364
rect 127 336 313 344
rect 327 336 373 344
rect 416 344 424 353
rect 416 336 653 344
rect 976 344 984 353
rect 947 336 984 344
rect 1267 336 1333 344
rect 1687 336 1733 344
rect 1827 336 1913 344
rect 1927 336 2273 344
rect 2467 336 2673 344
rect 2707 336 2753 344
rect 2887 336 2933 344
rect 3727 336 3833 344
rect 3887 336 3993 344
rect 4007 336 4213 344
rect 4236 344 4244 356
rect 4387 356 4484 364
rect 4236 336 4253 344
rect 267 316 293 324
rect 307 316 433 324
rect 1547 316 1613 324
rect 2327 316 2353 324
rect 2447 316 2573 324
rect 2847 316 2893 324
rect 2927 316 2993 324
rect 3167 316 3273 324
rect 3287 316 3333 324
rect 4276 324 4284 353
rect 4476 344 4484 356
rect 4507 356 4533 364
rect 4587 356 4633 364
rect 4687 356 4733 364
rect 4896 356 4953 364
rect 4896 347 4904 356
rect 5156 364 5164 373
rect 5636 367 5644 376
rect 5156 356 5173 364
rect 5247 356 5333 364
rect 5747 356 5793 364
rect 4476 336 4593 344
rect 5047 336 5153 344
rect 5207 336 5373 344
rect 5476 344 5484 353
rect 5476 336 5613 344
rect 4187 316 4284 324
rect 4327 316 4613 324
rect 4767 316 4813 324
rect 4987 316 5133 324
rect 5427 316 5493 324
rect 347 296 393 304
rect 987 296 1053 304
rect 1067 296 1633 304
rect 2387 296 2633 304
rect 3447 296 3673 304
rect 3687 296 4233 304
rect 4247 296 4413 304
rect 827 276 1073 284
rect 1087 276 1193 284
rect 4187 276 4573 284
rect 287 256 373 264
rect 387 256 593 264
rect 4027 256 4453 264
rect 487 236 573 244
rect 4647 236 4853 244
rect 5207 236 5353 244
rect 527 216 833 224
rect 847 216 913 224
rect 927 216 1013 224
rect 4607 216 4693 224
rect 4707 216 4953 224
rect 4967 216 5313 224
rect 427 196 553 204
rect 567 196 673 204
rect 867 196 1133 204
rect 1607 196 2173 204
rect 2527 196 2713 204
rect 3327 196 3373 204
rect 3387 196 3553 204
rect 4067 196 4133 204
rect 4147 196 4333 204
rect 4347 196 4993 204
rect 5016 196 5093 204
rect 167 176 213 184
rect 227 176 533 184
rect 587 176 633 184
rect 647 176 873 184
rect 907 176 1173 184
rect 1247 176 1313 184
rect 1347 176 1433 184
rect 1747 176 1893 184
rect 2187 176 2253 184
rect 2667 176 3033 184
rect 3207 176 3553 184
rect 3567 176 3733 184
rect 5016 184 5024 196
rect 5227 196 5333 204
rect 4767 176 5024 184
rect 5047 176 5073 184
rect 5087 176 5453 184
rect 5627 176 5673 184
rect 5687 176 5733 184
rect 107 156 173 164
rect 656 156 953 164
rect 656 147 664 156
rect 1287 156 1293 164
rect 1307 156 1413 164
rect 1707 156 1793 164
rect 1807 156 1913 164
rect 2127 156 2153 164
rect 2167 156 2333 164
rect 2347 156 2453 164
rect 2476 156 2613 164
rect 96 136 113 144
rect 96 124 104 136
rect 147 136 193 144
rect 407 136 473 144
rect 567 136 653 144
rect 707 136 833 144
rect 887 136 1193 144
rect 1207 136 1233 144
rect 1587 136 1673 144
rect 1727 136 1753 144
rect 2476 144 2484 156
rect 2636 156 2913 164
rect 2636 147 2644 156
rect 2936 156 3413 164
rect 1967 136 2484 144
rect 2687 136 2713 144
rect 2936 144 2944 156
rect 3867 156 4073 164
rect 4107 156 4113 164
rect 4127 156 4293 164
rect 4307 156 4713 164
rect 4887 156 4973 164
rect 5027 156 5113 164
rect 5127 156 5233 164
rect 5247 156 5293 164
rect 2847 136 2944 144
rect 2936 127 2944 136
rect 3067 136 3173 144
rect 3227 136 3293 144
rect 3347 136 3393 144
rect 3447 136 3533 144
rect 3676 136 4013 144
rect 3676 127 3684 136
rect 4467 136 4553 144
rect 4567 136 4604 144
rect 87 116 104 124
rect 127 116 153 124
rect 187 116 233 124
rect 847 116 893 124
rect 907 116 933 124
rect 967 116 1033 124
rect 1047 116 1493 124
rect 1987 116 2073 124
rect 2147 116 2393 124
rect 2407 116 2473 124
rect 3007 116 3073 124
rect 4007 116 4093 124
rect 4407 116 4513 124
rect 4596 124 4604 136
rect 4627 136 4833 144
rect 5007 136 5033 144
rect 5056 136 5233 144
rect 5056 124 5064 136
rect 5367 136 5493 144
rect 5607 136 5653 144
rect 4596 116 5064 124
rect 5267 116 5373 124
rect 5447 116 5673 124
rect 207 96 793 104
rect 1936 104 1944 113
rect 1867 96 2093 104
rect 2787 96 2893 104
rect 2907 96 3153 104
rect 3647 96 4533 104
rect 4576 104 4584 113
rect 4576 96 4633 104
rect 2287 36 2673 44
rect 2647 16 2953 24
use INVX2  _920_
timestamp 0
transform -1 0 3730 0 -1 2170
box -6 -8 66 248
use AND2X2  _921_
timestamp 0
transform 1 0 4110 0 -1 4570
box -6 -8 106 248
use NAND2X1  _922_
timestamp 0
transform -1 0 3970 0 1 4090
box -6 -8 86 248
use INVX1  _923_
timestamp 0
transform -1 0 3970 0 -1 5050
box -6 -8 66 248
use INVX2  _924_
timestamp 0
transform 1 0 4290 0 1 2650
box -6 -8 66 248
use NOR2X1  _925_
timestamp 0
transform -1 0 3710 0 1 3610
box -6 -8 86 248
use NAND2X1  _926_
timestamp 0
transform 1 0 2370 0 1 4570
box -6 -8 86 248
use OR2X2  _927_
timestamp 0
transform -1 0 1290 0 1 5530
box -6 -8 106 248
use NAND3X1  _928_
timestamp 0
transform 1 0 2250 0 -1 4090
box -6 -8 106 248
use NAND3X1  _929_
timestamp 0
transform 1 0 2110 0 1 4090
box -6 -8 106 248
use NOR2X1  _930_
timestamp 0
transform -1 0 2330 0 1 4090
box -6 -8 86 248
use INVX1  _931_
timestamp 0
transform -1 0 1070 0 -1 4570
box -6 -8 66 248
use NAND3X1  _932_
timestamp 0
transform -1 0 1850 0 -1 4570
box -6 -8 106 248
use INVX2  _933_
timestamp 0
transform 1 0 3950 0 -1 2170
box -6 -8 66 248
use NAND2X1  _934_
timestamp 0
transform -1 0 2610 0 -1 4090
box -6 -8 86 248
use OAI21X1  _935_
timestamp 0
transform -1 0 2490 0 -1 4090
box -6 -8 106 248
use INVX1  _936_
timestamp 0
transform 1 0 1470 0 1 4570
box -6 -8 66 248
use OAI21X1  _937_
timestamp 0
transform -1 0 1290 0 1 4570
box -6 -8 106 248
use NAND3X1  _938_
timestamp 0
transform -1 0 2210 0 1 4570
box -6 -8 106 248
use INVX1  _939_
timestamp 0
transform 1 0 1130 0 1 5050
box -6 -8 66 248
use NAND3X1  _940_
timestamp 0
transform -1 0 2650 0 1 4090
box -6 -8 106 248
use NAND3X1  _941_
timestamp 0
transform -1 0 1930 0 1 4090
box -6 -8 106 248
use NOR2X1  _942_
timestamp 0
transform -1 0 1650 0 1 4090
box -6 -8 86 248
use INVX1  _943_
timestamp 0
transform -1 0 1150 0 1 4570
box -6 -8 66 248
use INVX1  _944_
timestamp 0
transform 1 0 2450 0 1 1210
box -6 -8 66 248
use NAND2X1  _945_
timestamp 0
transform 1 0 2530 0 1 3610
box -6 -8 86 248
use OAI21X1  _946_
timestamp 0
transform -1 0 2490 0 1 4090
box -6 -8 106 248
use NAND3X1  _947_
timestamp 0
transform -1 0 1090 0 1 5050
box -6 -8 106 248
use INVX1  _948_
timestamp 0
transform -1 0 1350 0 -1 5050
box -6 -8 66 248
use OAI21X1  _949_
timestamp 0
transform -1 0 970 0 -1 5050
box -6 -8 106 248
use NAND3X1  _950_
timestamp 0
transform 1 0 850 0 1 5050
box -6 -8 106 248
use INVX1  _951_
timestamp 0
transform -1 0 4050 0 1 3610
box -6 -8 66 248
use NAND2X1  _952_
timestamp 0
transform 1 0 2490 0 1 4570
box -6 -8 86 248
use OAI21X1  _953_
timestamp 0
transform -1 0 1490 0 1 5050
box -6 -8 106 248
use NAND2X1  _954_
timestamp 0
transform -1 0 850 0 1 5530
box -6 -8 86 248
use AOI21X1  _955_
timestamp 0
transform -1 0 810 0 1 5050
box -6 -8 106 248
use OAI21X1  _956_
timestamp 0
transform 1 0 790 0 -1 5530
box -6 -8 106 248
use OAI21X1  _957_
timestamp 0
transform -1 0 830 0 -1 5050
box -6 -8 106 248
use NAND3X1  _958_
timestamp 0
transform 1 0 1970 0 1 4090
box -6 -8 106 248
use NAND3X1  _959_
timestamp 0
transform -1 0 2210 0 -1 4090
box -6 -8 106 248
use OR2X2  _960_
timestamp 0
transform -1 0 750 0 1 4090
box -6 -8 106 248
use INVX1  _961_
timestamp 0
transform -1 0 5170 0 -1 4090
box -6 -8 66 248
use NAND2X1  _962_
timestamp 0
transform 1 0 2650 0 -1 4090
box -6 -8 86 248
use OAI21X1  _963_
timestamp 0
transform -1 0 2050 0 -1 4090
box -6 -8 106 248
use NAND3X1  _964_
timestamp 0
transform -1 0 1790 0 1 4090
box -6 -8 106 248
use INVX1  _965_
timestamp 0
transform -1 0 110 0 -1 4090
box -6 -8 66 248
use NAND3X1  _966_
timestamp 0
transform -1 0 470 0 1 4090
box -6 -8 106 248
use NOR2X1  _967_
timestamp 0
transform -1 0 650 0 -1 4090
box -6 -8 86 248
use INVX1  _968_
timestamp 0
transform -1 0 370 0 -1 4090
box -6 -8 66 248
use OAI21X1  _969_
timestamp 0
transform -1 0 310 0 1 4090
box -6 -8 106 248
use NAND3X1  _970_
timestamp 0
transform -1 0 290 0 -1 4570
box -6 -8 106 248
use AOI21X1  _971_
timestamp 0
transform -1 0 1110 0 -1 5050
box -6 -8 106 248
use OAI21X1  _972_
timestamp 0
transform -1 0 170 0 1 4090
box -6 -8 106 248
use NAND3X1  _973_
timestamp 0
transform -1 0 610 0 1 4090
box -6 -8 106 248
use NAND3X1  _974_
timestamp 0
transform -1 0 290 0 1 4570
box -6 -8 106 248
use NAND2X1  _975_
timestamp 0
transform 1 0 4170 0 1 2650
box -6 -8 86 248
use INVX2  _976_
timestamp 0
transform -1 0 3990 0 1 2650
box -6 -8 66 248
use NAND2X1  _977_
timestamp 0
transform -1 0 1710 0 -1 4570
box -6 -8 86 248
use INVX1  _978_
timestamp 0
transform 1 0 890 0 1 4570
box -6 -8 66 248
use NAND3X1  _979_
timestamp 0
transform -1 0 2270 0 -1 4570
box -6 -8 106 248
use NAND3X1  _980_
timestamp 0
transform -1 0 2110 0 -1 4570
box -6 -8 106 248
use NOR2X1  _981_
timestamp 0
transform -1 0 1970 0 -1 4570
box -6 -8 86 248
use OAI21X1  _982_
timestamp 0
transform 1 0 1490 0 -1 4570
box -6 -8 106 248
use INVX1  _983_
timestamp 0
transform 1 0 770 0 -1 4570
box -6 -8 66 248
use OAI21X1  _984_
timestamp 0
transform -1 0 730 0 -1 4570
box -6 -8 106 248
use INVX1  _985_
timestamp 0
transform 1 0 990 0 1 4570
box -6 -8 66 248
use NAND3X1  _986_
timestamp 0
transform -1 0 850 0 1 4570
box -6 -8 106 248
use NAND2X1  _987_
timestamp 0
transform -1 0 690 0 -1 5050
box -6 -8 86 248
use NAND3X1  _988_
timestamp 0
transform -1 0 290 0 -1 5050
box -6 -8 106 248
use AOI21X1  _989_
timestamp 0
transform 1 0 330 0 1 4570
box -6 -8 106 248
use AOI21X1  _990_
timestamp 0
transform 1 0 330 0 -1 4570
box -6 -8 106 248
use NAND3X1  _991_
timestamp 0
transform -1 0 690 0 1 4570
box -6 -8 106 248
use OAI21X1  _992_
timestamp 0
transform -1 0 590 0 -1 4570
box -6 -8 106 248
use NAND2X1  _993_
timestamp 0
transform 1 0 470 0 1 4570
box -6 -8 86 248
use OAI21X1  _994_
timestamp 0
transform -1 0 150 0 -1 5050
box -6 -8 106 248
use NAND3X1  _995_
timestamp 0
transform -1 0 150 0 1 5050
box -6 -8 106 248
use AOI21X1  _996_
timestamp 0
transform 1 0 190 0 1 5050
box -6 -8 106 248
use OAI21X1  _997_
timestamp 0
transform -1 0 150 0 -1 5530
box -6 -8 106 248
use OAI21X1  _998_
timestamp 0
transform -1 0 150 0 -1 4570
box -6 -8 106 248
use AOI21X1  _999_
timestamp 0
transform 1 0 430 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1000_
timestamp 0
transform -1 0 1930 0 1 730
box -6 -8 106 248
use NAND3X1  _1001_
timestamp 0
transform -1 0 2230 0 -1 1210
box -6 -8 106 248
use NOR2X1  _1002_
timestamp 0
transform 1 0 1290 0 -1 250
box -6 -8 86 248
use AND2X2  _1003_
timestamp 0
transform 1 0 1410 0 -1 250
box -6 -8 106 248
use NAND3X1  _1004_
timestamp 0
transform -1 0 1790 0 1 730
box -6 -8 106 248
use INVX1  _1005_
timestamp 0
transform 1 0 910 0 -1 250
box -6 -8 66 248
use OAI21X1  _1006_
timestamp 0
transform 1 0 630 0 -1 250
box -6 -8 106 248
use OR2X2  _1007_
timestamp 0
transform -1 0 1290 0 1 250
box -6 -8 106 248
use OAI21X1  _1008_
timestamp 0
transform -1 0 2090 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1009_
timestamp 0
transform -1 0 870 0 1 250
box -6 -8 106 248
use NAND3X1  _1010_
timestamp 0
transform -1 0 590 0 1 250
box -6 -8 106 248
use OAI21X1  _1011_
timestamp 0
transform 1 0 170 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1012_
timestamp 0
transform -1 0 870 0 -1 250
box -6 -8 106 248
use OAI21X1  _1013_
timestamp 0
transform -1 0 590 0 -1 250
box -6 -8 106 248
use NAND3X1  _1014_
timestamp 0
transform -1 0 150 0 -1 250
box -6 -8 106 248
use NAND3X1  _1015_
timestamp 0
transform -1 0 1830 0 -1 1210
box -6 -8 106 248
use INVX1  _1016_
timestamp 0
transform -1 0 1450 0 -1 1210
box -6 -8 66 248
use NAND3X1  _1017_
timestamp 0
transform -1 0 2270 0 1 1210
box -6 -8 106 248
use NAND3X1  _1018_
timestamp 0
transform -1 0 2330 0 -1 2170
box -6 -8 106 248
use NOR2X1  _1019_
timestamp 0
transform -1 0 1570 0 -1 1210
box -6 -8 86 248
use OAI21X1  _1020_
timestamp 0
transform -1 0 1510 0 1 1690
box -6 -8 106 248
use INVX1  _1021_
timestamp 0
transform -1 0 1210 0 -1 1210
box -6 -8 66 248
use OAI21X1  _1022_
timestamp 0
transform -1 0 1110 0 -1 1210
box -6 -8 106 248
use INVX1  _1023_
timestamp 0
transform 1 0 1450 0 1 730
box -6 -8 66 248
use INVX1  _1024_
timestamp 0
transform 1 0 1630 0 -1 1210
box -6 -8 66 248
use NAND2X1  _1025_
timestamp 0
transform 1 0 1550 0 1 730
box -6 -8 86 248
use NAND3X1  _1026_
timestamp 0
transform -1 0 1410 0 1 730
box -6 -8 106 248
use NAND2X1  _1027_
timestamp 0
transform 1 0 770 0 -1 730
box -6 -8 86 248
use NAND3X1  _1028_
timestamp 0
transform -1 0 450 0 -1 730
box -6 -8 106 248
use AOI21X1  _1029_
timestamp 0
transform 1 0 190 0 -1 250
box -6 -8 106 248
use AOI21X1  _1030_
timestamp 0
transform -1 0 450 0 -1 250
box -6 -8 106 248
use AND2X2  _1031_
timestamp 0
transform -1 0 730 0 1 250
box -6 -8 106 248
use OAI21X1  _1032_
timestamp 0
transform -1 0 290 0 1 250
box -6 -8 106 248
use AOI21X1  _1033_
timestamp 0
transform 1 0 190 0 1 730
box -6 -8 106 248
use AOI21X1  _1034_
timestamp 0
transform -1 0 150 0 1 4570
box -6 -8 106 248
use OAI21X1  _1035_
timestamp 0
transform -1 0 590 0 -1 730
box -6 -8 106 248
use NAND3X1  _1036_
timestamp 0
transform -1 0 150 0 1 250
box -6 -8 106 248
use AOI21X1  _1037_
timestamp 0
transform -1 0 310 0 -1 730
box -6 -8 106 248
use NAND2X1  _1038_
timestamp 0
transform -1 0 3070 0 1 2170
box -6 -8 86 248
use AOI21X1  _1039_
timestamp 0
transform 1 0 870 0 -1 4570
box -6 -8 106 248
use OR2X2  _1040_
timestamp 0
transform -1 0 1090 0 1 2170
box -6 -8 106 248
use INVX1  _1041_
timestamp 0
transform 1 0 5330 0 1 5050
box -6 -8 66 248
use NOR2X1  _1042_
timestamp 0
transform 1 0 4830 0 1 5050
box -6 -8 86 248
use INVX4  _1043_
timestamp 0
transform -1 0 2170 0 1 1690
box -6 -8 86 248
use OAI21X1  _1044_
timestamp 0
transform -1 0 1150 0 -1 2650
box -6 -8 106 248
use NAND2X1  _1045_
timestamp 0
transform -1 0 950 0 1 2170
box -6 -8 86 248
use INVX1  _1046_
timestamp 0
transform -1 0 110 0 -1 1210
box -6 -8 66 248
use OAI21X1  _1047_
timestamp 0
transform 1 0 290 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1048_
timestamp 0
transform -1 0 150 0 -1 730
box -6 -8 106 248
use NAND3X1  _1049_
timestamp 0
transform -1 0 150 0 1 730
box -6 -8 106 248
use NAND3X1  _1050_
timestamp 0
transform 1 0 70 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1051_
timestamp 0
transform 1 0 310 0 1 2170
box -6 -8 86 248
use NAND2X1  _1052_
timestamp 0
transform -1 0 130 0 1 2650
box -6 -8 86 248
use INVX1  _1053_
timestamp 0
transform 1 0 150 0 -1 2650
box -6 -8 66 248
use INVX1  _1054_
timestamp 0
transform -1 0 550 0 -1 2170
box -6 -8 66 248
use AOI21X1  _1055_
timestamp 0
transform 1 0 150 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1056_
timestamp 0
transform -1 0 450 0 1 250
box -6 -8 106 248
use AOI21X1  _1057_
timestamp 0
transform 1 0 1150 0 -1 250
box -6 -8 106 248
use NAND3X1  _1058_
timestamp 0
transform -1 0 2370 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1059_
timestamp 0
transform -1 0 2650 0 -1 1210
box -6 -8 106 248
use NOR2X1  _1060_
timestamp 0
transform -1 0 2130 0 -1 730
box -6 -8 86 248
use AND2X2  _1061_
timestamp 0
transform 1 0 2250 0 1 730
box -6 -8 106 248
use NAND3X1  _1062_
timestamp 0
transform 1 0 1970 0 1 730
box -6 -8 106 248
use INVX1  _1063_
timestamp 0
transform -1 0 1550 0 1 250
box -6 -8 66 248
use OAI21X1  _1064_
timestamp 0
transform -1 0 1730 0 -1 730
box -6 -8 106 248
use OR2X2  _1065_
timestamp 0
transform -1 0 2270 0 -1 730
box -6 -8 106 248
use NAND2X1  _1066_
timestamp 0
transform 1 0 2690 0 1 1690
box -6 -8 86 248
use OAI21X1  _1067_
timestamp 0
transform -1 0 2510 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1068_
timestamp 0
transform -1 0 1870 0 -1 730
box -6 -8 106 248
use NAND3X1  _1069_
timestamp 0
transform 1 0 1490 0 -1 730
box -6 -8 106 248
use OAI21X1  _1070_
timestamp 0
transform 1 0 1010 0 -1 250
box -6 -8 106 248
use NAND3X1  _1071_
timestamp 0
transform -1 0 1430 0 1 250
box -6 -8 106 248
use OAI21X1  _1072_
timestamp 0
transform -1 0 1690 0 1 250
box -6 -8 106 248
use NAND3X1  _1073_
timestamp 0
transform 1 0 1050 0 1 250
box -6 -8 106 248
use NAND3X1  _1074_
timestamp 0
transform -1 0 2410 0 1 1210
box -6 -8 106 248
use INVX1  _1075_
timestamp 0
transform -1 0 2110 0 1 1210
box -6 -8 66 248
use NAND3X1  _1076_
timestamp 0
transform 1 0 3790 0 -1 2170
box -6 -8 106 248
use INVX1  _1077_
timestamp 0
transform 1 0 3890 0 1 3610
box -6 -8 66 248
use NAND3X1  _1078_
timestamp 0
transform 1 0 2250 0 1 3610
box -6 -8 106 248
use OAI21X1  _1079_
timestamp 0
transform -1 0 2490 0 1 3610
box -6 -8 106 248
use OAI21X1  _1080_
timestamp 0
transform -1 0 1790 0 1 1690
box -6 -8 106 248
use NAND2X1  _1081_
timestamp 0
transform 1 0 1790 0 1 1210
box -6 -8 86 248
use INVX1  _1082_
timestamp 0
transform -1 0 1590 0 -1 1690
box -6 -8 66 248
use NAND2X1  _1083_
timestamp 0
transform -1 0 1590 0 1 1210
box -6 -8 86 248
use NAND3X1  _1084_
timestamp 0
transform -1 0 2010 0 1 1210
box -6 -8 106 248
use NAND2X1  _1085_
timestamp 0
transform -1 0 1950 0 -1 1210
box -6 -8 86 248
use NAND3X1  _1086_
timestamp 0
transform -1 0 1150 0 -1 730
box -6 -8 106 248
use AOI21X1  _1087_
timestamp 0
transform -1 0 1010 0 1 250
box -6 -8 106 248
use AOI21X1  _1088_
timestamp 0
transform -1 0 1430 0 -1 730
box -6 -8 106 248
use NAND3X1  _1089_
timestamp 0
transform -1 0 1750 0 1 1210
box -6 -8 106 248
use NAND2X1  _1090_
timestamp 0
transform -1 0 2390 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1091_
timestamp 0
transform 1 0 1550 0 1 1690
box -6 -8 106 248
use NAND2X1  _1092_
timestamp 0
transform -1 0 1470 0 1 1210
box -6 -8 86 248
use OAI21X1  _1093_
timestamp 0
transform -1 0 990 0 1 730
box -6 -8 106 248
use AOI21X1  _1094_
timestamp 0
transform -1 0 570 0 1 730
box -6 -8 106 248
use AOI21X1  _1095_
timestamp 0
transform 1 0 630 0 -1 730
box -6 -8 106 248
use OAI21X1  _1096_
timestamp 0
transform -1 0 1010 0 -1 730
box -6 -8 106 248
use NAND3X1  _1097_
timestamp 0
transform -1 0 1130 0 1 730
box -6 -8 106 248
use AOI21X1  _1098_
timestamp 0
transform 1 0 750 0 1 730
box -6 -8 106 248
use NAND2X1  _1099_
timestamp 0
transform -1 0 2030 0 1 1690
box -6 -8 86 248
use INVX1  _1100_
timestamp 0
transform -1 0 1090 0 1 1210
box -6 -8 66 248
use AOI21X1  _1101_
timestamp 0
transform 1 0 1250 0 -1 1210
box -6 -8 106 248
use INVX1  _1102_
timestamp 0
transform -1 0 970 0 1 1690
box -6 -8 66 248
use OAI21X1  _1103_
timestamp 0
transform -1 0 1270 0 1 1690
box -6 -8 106 248
use NAND2X1  _1104_
timestamp 0
transform -1 0 1910 0 1 1690
box -6 -8 86 248
use INVX1  _1105_
timestamp 0
transform -1 0 1370 0 1 1690
box -6 -8 66 248
use NAND2X1  _1106_
timestamp 0
transform 1 0 1270 0 1 1210
box -6 -8 86 248
use NAND3X1  _1107_
timestamp 0
transform 1 0 1130 0 1 1210
box -6 -8 106 248
use NAND2X1  _1108_
timestamp 0
transform -1 0 1210 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1109_
timestamp 0
transform -1 0 1130 0 1 1690
box -6 -8 106 248
use NAND3X1  _1110_
timestamp 0
transform -1 0 1090 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1111_
timestamp 0
transform 1 0 910 0 1 1210
box -6 -8 86 248
use OAI21X1  _1112_
timestamp 0
transform 1 0 710 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1113_
timestamp 0
transform -1 0 710 0 1 730
box -6 -8 106 248
use NAND3X1  _1114_
timestamp 0
transform -1 0 430 0 1 730
box -6 -8 106 248
use AND2X2  _1115_
timestamp 0
transform -1 0 870 0 1 1210
box -6 -8 106 248
use NAND3X1  _1116_
timestamp 0
transform -1 0 430 0 1 1210
box -6 -8 106 248
use NAND3X1  _1117_
timestamp 0
transform -1 0 310 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1118_
timestamp 0
transform 1 0 430 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1119_
timestamp 0
transform -1 0 670 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1120_
timestamp 0
transform -1 0 710 0 1 1210
box -6 -8 106 248
use NAND3X1  _1121_
timestamp 0
transform -1 0 150 0 1 1210
box -6 -8 106 248
use NAND3X1  _1122_
timestamp 0
transform -1 0 310 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1123_
timestamp 0
transform 1 0 190 0 1 1210
box -6 -8 106 248
use AOI21X1  _1124_
timestamp 0
transform 1 0 350 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1125_
timestamp 0
transform 1 0 430 0 1 2170
box -6 -8 106 248
use NAND3X1  _1126_
timestamp 0
transform 1 0 390 0 -1 2650
box -6 -8 106 248
use AOI21X1  _1127_
timestamp 0
transform -1 0 350 0 -1 2650
box -6 -8 106 248
use NOR2X1  _1128_
timestamp 0
transform 1 0 1370 0 -1 5530
box -6 -8 86 248
use INVX1  _1129_
timestamp 0
transform -1 0 1450 0 -1 4570
box -6 -8 66 248
use AOI21X1  _1130_
timestamp 0
transform -1 0 1350 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1131_
timestamp 0
transform -1 0 1250 0 -1 5050
box -6 -8 106 248
use NAND3X1  _1132_
timestamp 0
transform -1 0 1330 0 1 5050
box -6 -8 106 248
use AOI21X1  _1133_
timestamp 0
transform -1 0 1170 0 -1 5530
box -6 -8 106 248
use AND2X2  _1134_
timestamp 0
transform -1 0 1430 0 1 5530
box -6 -8 106 248
use NOR2X1  _1135_
timestamp 0
transform 1 0 1050 0 1 5530
box -6 -8 86 248
use NAND3X1  _1136_
timestamp 0
transform 1 0 1210 0 -1 5530
box -6 -8 106 248
use AOI21X1  _1137_
timestamp 0
transform -1 0 990 0 1 5530
box -6 -8 106 248
use OAI21X1  _1138_
timestamp 0
transform 1 0 470 0 -1 5050
box -6 -8 106 248
use NAND3X1  _1139_
timestamp 0
transform 1 0 330 0 -1 5050
box -6 -8 106 248
use NAND3X1  _1140_
timestamp 0
transform 1 0 490 0 1 5530
box -6 -8 106 248
use NAND3X1  _1141_
timestamp 0
transform 1 0 650 0 -1 5530
box -6 -8 106 248
use NAND3X1  _1142_
timestamp 0
transform 1 0 930 0 -1 5530
box -6 -8 106 248
use NAND3X1  _1143_
timestamp 0
transform -1 0 1210 0 -1 4570
box -6 -8 106 248
use NAND3X1  _1144_
timestamp 0
transform 1 0 2770 0 -1 4090
box -6 -8 106 248
use INVX1  _1145_
timestamp 0
transform -1 0 3350 0 1 3610
box -6 -8 66 248
use NAND3X1  _1146_
timestamp 0
transform 1 0 2910 0 -1 4090
box -6 -8 106 248
use INVX1  _1147_
timestamp 0
transform -1 0 3110 0 -1 4090
box -6 -8 66 248
use NAND2X1  _1148_
timestamp 0
transform -1 0 3250 0 1 3610
box -6 -8 86 248
use NAND2X1  _1149_
timestamp 0
transform -1 0 3170 0 1 3130
box -6 -8 86 248
use OAI21X1  _1150_
timestamp 0
transform 1 0 2650 0 1 3610
box -6 -8 106 248
use INVX1  _1151_
timestamp 0
transform -1 0 2850 0 1 3610
box -6 -8 66 248
use OAI21X1  _1152_
timestamp 0
transform -1 0 2990 0 1 3610
box -6 -8 106 248
use OAI21X1  _1153_
timestamp 0
transform 1 0 1330 0 1 4570
box -6 -8 106 248
use NAND3X1  _1154_
timestamp 0
transform -1 0 1290 0 1 4090
box -6 -8 106 248
use NAND2X1  _1155_
timestamp 0
transform -1 0 1530 0 1 4090
box -6 -8 86 248
use AOI21X1  _1156_
timestamp 0
transform -1 0 1130 0 1 4090
box -6 -8 106 248
use OAI21X1  _1157_
timestamp 0
transform -1 0 890 0 1 4090
box -6 -8 106 248
use OAI21X1  _1158_
timestamp 0
transform -1 0 730 0 1 5530
box -6 -8 106 248
use NAND3X1  _1159_
timestamp 0
transform -1 0 530 0 1 5050
box -6 -8 106 248
use INVX1  _1160_
timestamp 0
transform 1 0 330 0 1 5050
box -6 -8 66 248
use AOI21X1  _1161_
timestamp 0
transform -1 0 450 0 1 5530
box -6 -8 106 248
use OAI21X1  _1162_
timestamp 0
transform -1 0 150 0 1 5530
box -6 -8 106 248
use NAND3X1  _1163_
timestamp 0
transform -1 0 450 0 -1 5530
box -6 -8 106 248
use INVX1  _1164_
timestamp 0
transform -1 0 110 0 1 3130
box -6 -8 66 248
use INVX1  _1165_
timestamp 0
transform -1 0 110 0 -1 2650
box -6 -8 66 248
use NAND3X1  _1166_
timestamp 0
transform -1 0 270 0 1 2170
box -6 -8 106 248
use AND2X2  _1167_
timestamp 0
transform -1 0 170 0 -1 3130
box -6 -8 106 248
use INVX1  _1168_
timestamp 0
transform 1 0 950 0 -1 4090
box -6 -8 66 248
use INVX1  _1169_
timestamp 0
transform 1 0 930 0 1 4090
box -6 -8 66 248
use NAND3X1  _1170_
timestamp 0
transform 1 0 1050 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1171_
timestamp 0
transform 1 0 3030 0 1 3610
box -6 -8 86 248
use OR2X2  _1172_
timestamp 0
transform 1 0 3330 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1173_
timestamp 0
transform 1 0 3610 0 -1 2650
box -6 -8 86 248
use NAND2X1  _1174_
timestamp 0
transform -1 0 3310 0 1 3130
box -6 -8 86 248
use NOR2X1  _1175_
timestamp 0
transform 1 0 3550 0 1 2650
box -6 -8 86 248
use INVX1  _1176_
timestamp 0
transform 1 0 4390 0 1 2650
box -6 -8 66 248
use OAI21X1  _1177_
timestamp 0
transform -1 0 4130 0 1 2650
box -6 -8 106 248
use NAND3X1  _1178_
timestamp 0
transform -1 0 3430 0 -1 2650
box -6 -8 106 248
use INVX1  _1179_
timestamp 0
transform -1 0 3010 0 -1 2650
box -6 -8 66 248
use INVX1  _1180_
timestamp 0
transform -1 0 770 0 -1 4090
box -6 -8 66 248
use OAI21X1  _1181_
timestamp 0
transform 1 0 810 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1182_
timestamp 0
transform -1 0 1210 0 -1 3610
box -6 -8 106 248
use AOI21X1  _1183_
timestamp 0
transform 1 0 570 0 1 5050
box -6 -8 106 248
use NOR3X1  _1184_
timestamp 0
transform -1 0 490 0 1 3610
box -6 -8 186 248
use OAI21X1  _1185_
timestamp 0
transform 1 0 190 0 1 5530
box -6 -8 106 248
use NAND3X1  _1186_
timestamp 0
transform -1 0 590 0 -1 5530
box -6 -8 106 248
use NAND3X1  _1187_
timestamp 0
transform -1 0 310 0 -1 5530
box -6 -8 106 248
use NAND3X1  _1188_
timestamp 0
transform -1 0 270 0 1 3610
box -6 -8 106 248
use INVX1  _1189_
timestamp 0
transform -1 0 350 0 1 3130
box -6 -8 66 248
use OAI21X1  _1190_
timestamp 0
transform -1 0 250 0 1 3130
box -6 -8 106 248
use OAI21X1  _1191_
timestamp 0
transform 1 0 170 0 1 2650
box -6 -8 106 248
use AOI21X1  _1192_
timestamp 0
transform 1 0 350 0 -1 2170
box -6 -8 106 248
use NOR2X1  _1193_
timestamp 0
transform 1 0 1270 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1194_
timestamp 0
transform -1 0 950 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1195_
timestamp 0
transform -1 0 570 0 1 1210
box -6 -8 106 248
use INVX1  _1196_
timestamp 0
transform 1 0 5110 0 1 3610
box -6 -8 66 248
use NOR2X1  _1197_
timestamp 0
transform 1 0 4610 0 1 3610
box -6 -8 86 248
use NAND2X1  _1198_
timestamp 0
transform 1 0 3810 0 1 2650
box -6 -8 86 248
use INVX1  _1199_
timestamp 0
transform 1 0 1590 0 -1 2650
box -6 -8 66 248
use NAND2X1  _1200_
timestamp 0
transform -1 0 1990 0 1 2650
box -6 -8 86 248
use AOI22X1  _1201_
timestamp 0
transform 1 0 1630 0 -1 1690
box -6 -8 126 248
use OR2X2  _1202_
timestamp 0
transform -1 0 1590 0 1 2650
box -6 -8 106 248
use OAI21X1  _1203_
timestamp 0
transform -1 0 1930 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1204_
timestamp 0
transform -1 0 1550 0 -1 2650
box -6 -8 106 248
use NOR2X1  _1205_
timestamp 0
transform 1 0 1630 0 1 2650
box -6 -8 86 248
use AND2X2  _1206_
timestamp 0
transform -1 0 1850 0 1 2650
box -6 -8 106 248
use OAI21X1  _1207_
timestamp 0
transform -1 0 1310 0 1 2650
box -6 -8 106 248
use NAND2X1  _1208_
timestamp 0
transform -1 0 1270 0 -1 2650
box -6 -8 86 248
use AOI21X1  _1209_
timestamp 0
transform 1 0 1190 0 -1 730
box -6 -8 106 248
use NAND3X1  _1210_
timestamp 0
transform 1 0 2950 0 1 3130
box -6 -8 106 248
use NAND3X1  _1211_
timestamp 0
transform 1 0 4170 0 -1 3130
box -6 -8 106 248
use NOR2X1  _1212_
timestamp 0
transform 1 0 4050 0 -1 3130
box -6 -8 86 248
use AND2X2  _1213_
timestamp 0
transform -1 0 4010 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1214_
timestamp 0
transform -1 0 3710 0 -1 3130
box -6 -8 106 248
use INVX1  _1215_
timestamp 0
transform 1 0 3350 0 1 3130
box -6 -8 66 248
use OR2X2  _1216_
timestamp 0
transform -1 0 3850 0 -1 3130
box -6 -8 106 248
use INVX1  _1217_
timestamp 0
transform 1 0 3870 0 1 3130
box -6 -8 66 248
use OAI21X1  _1218_
timestamp 0
transform -1 0 3830 0 1 3130
box -6 -8 106 248
use NAND3X1  _1219_
timestamp 0
transform -1 0 3550 0 1 3130
box -6 -8 106 248
use NAND2X1  _1220_
timestamp 0
transform 1 0 3070 0 -1 3130
box -6 -8 86 248
use AOI21X1  _1221_
timestamp 0
transform 1 0 1910 0 -1 730
box -6 -8 106 248
use NAND3X1  _1222_
timestamp 0
transform 1 0 2810 0 1 3130
box -6 -8 106 248
use NAND3X1  _1223_
timestamp 0
transform -1 0 3110 0 1 2650
box -6 -8 106 248
use NOR2X1  _1224_
timestamp 0
transform 1 0 2930 0 -1 3130
box -6 -8 86 248
use AND2X2  _1225_
timestamp 0
transform -1 0 2810 0 1 2650
box -6 -8 106 248
use NOR2X1  _1226_
timestamp 0
transform 1 0 2450 0 1 2650
box -6 -8 86 248
use NAND2X1  _1227_
timestamp 0
transform 1 0 2390 0 -1 2650
box -6 -8 86 248
use OAI21X1  _1228_
timestamp 0
transform 1 0 2110 0 1 730
box -6 -8 106 248
use OAI21X1  _1229_
timestamp 0
transform 1 0 2670 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1230_
timestamp 0
transform -1 0 2210 0 -1 2650
box -6 -8 106 248
use AND2X2  _1231_
timestamp 0
transform -1 0 3290 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1232_
timestamp 0
transform -1 0 2390 0 1 2650
box -6 -8 86 248
use OAI21X1  _1233_
timestamp 0
transform -1 0 2630 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1234_
timestamp 0
transform -1 0 2670 0 1 2650
box -6 -8 106 248
use NAND3X1  _1235_
timestamp 0
transform -1 0 2050 0 1 2170
box -6 -8 106 248
use OAI21X1  _1236_
timestamp 0
transform 1 0 1170 0 1 730
box -6 -8 106 248
use AOI22X1  _1237_
timestamp 0
transform -1 0 2750 0 -1 3130
box -6 -8 126 248
use AOI21X1  _1238_
timestamp 0
transform -1 0 2350 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1239_
timestamp 0
transform -1 0 1630 0 1 2170
box -6 -8 106 248
use NAND3X1  _1240_
timestamp 0
transform -1 0 1330 0 1 2170
box -6 -8 106 248
use AND2X2  _1241_
timestamp 0
transform 1 0 1310 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1242_
timestamp 0
transform -1 0 1910 0 1 2170
box -6 -8 106 248
use OAI21X1  _1243_
timestamp 0
transform 1 0 1730 0 -1 2170
box -6 -8 106 248
use NAND3X1  _1244_
timestamp 0
transform -1 0 1690 0 -1 2170
box -6 -8 106 248
use NAND3X1  _1245_
timestamp 0
transform -1 0 570 0 1 1690
box -6 -8 106 248
use AOI21X1  _1246_
timestamp 0
transform 1 0 870 0 -1 1210
box -6 -8 106 248
use AOI21X1  _1247_
timestamp 0
transform -1 0 1550 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1248_
timestamp 0
transform -1 0 1470 0 1 2170
box -6 -8 106 248
use OAI21X1  _1249_
timestamp 0
transform -1 0 1270 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1250_
timestamp 0
transform 1 0 190 0 1 1690
box -6 -8 106 248
use INVX1  _1251_
timestamp 0
transform 1 0 750 0 -1 1690
box -6 -8 66 248
use NAND3X1  _1252_
timestamp 0
transform -1 0 1130 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1253_
timestamp 0
transform -1 0 1410 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1254_
timestamp 0
transform -1 0 830 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1255_
timestamp 0
transform -1 0 690 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1256_
timestamp 0
transform -1 0 670 0 1 2170
box -6 -8 106 248
use NAND3X1  _1257_
timestamp 0
transform 1 0 870 0 -1 2170
box -6 -8 106 248
use NAND3X1  _1258_
timestamp 0
transform -1 0 150 0 1 1690
box -6 -8 106 248
use NAND3X1  _1259_
timestamp 0
transform -1 0 830 0 1 2170
box -6 -8 106 248
use AND2X2  _1260_
timestamp 0
transform 1 0 670 0 1 2650
box -6 -8 106 248
use NAND2X1  _1261_
timestamp 0
transform 1 0 810 0 1 2650
box -6 -8 86 248
use INVX1  _1262_
timestamp 0
transform 1 0 530 0 -1 2650
box -6 -8 66 248
use INVX1  _1263_
timestamp 0
transform -1 0 370 0 1 2650
box -6 -8 66 248
use NAND2X1  _1264_
timestamp 0
transform 1 0 370 0 -1 3130
box -6 -8 86 248
use NAND3X1  _1265_
timestamp 0
transform 1 0 230 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1266_
timestamp 0
transform -1 0 590 0 -1 3130
box -6 -8 106 248
use AOI21X1  _1267_
timestamp 0
transform 1 0 410 0 1 2650
box -6 -8 106 248
use NAND2X1  _1268_
timestamp 0
transform -1 0 630 0 1 2650
box -6 -8 86 248
use NAND2X1  _1269_
timestamp 0
transform -1 0 1130 0 -1 3130
box -6 -8 86 248
use NAND2X1  _1270_
timestamp 0
transform 1 0 1070 0 1 2650
box -6 -8 86 248
use NOR2X1  _1271_
timestamp 0
transform -1 0 3270 0 -1 1210
box -6 -8 86 248
use INVX1  _1272_
timestamp 0
transform 1 0 2710 0 -1 1210
box -6 -8 66 248
use INVX2  _1273_
timestamp 0
transform 1 0 1130 0 1 2170
box -6 -8 66 248
use OAI21X1  _1274_
timestamp 0
transform -1 0 2950 0 1 1210
box -6 -8 106 248
use NAND3X1  _1275_
timestamp 0
transform -1 0 2910 0 1 1690
box -6 -8 106 248
use OAI21X1  _1276_
timestamp 0
transform -1 0 2910 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1277_
timestamp 0
transform 1 0 2430 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1278_
timestamp 0
transform 1 0 2290 0 -1 1690
box -6 -8 106 248
use AND2X2  _1279_
timestamp 0
transform -1 0 3510 0 1 2650
box -6 -8 106 248
use OAI21X1  _1280_
timestamp 0
transform -1 0 3370 0 1 2650
box -6 -8 106 248
use MUX2X1  _1281_
timestamp 0
transform 1 0 3210 0 1 1690
box -6 -8 126 248
use AOI21X1  _1282_
timestamp 0
transform -1 0 3350 0 1 2170
box -6 -8 106 248
use NAND2X1  _1283_
timestamp 0
transform 1 0 3150 0 1 2650
box -6 -8 86 248
use NAND2X1  _1284_
timestamp 0
transform 1 0 630 0 -1 1690
box -6 -8 86 248
use NOR2X1  _1285_
timestamp 0
transform -1 0 710 0 1 1690
box -6 -8 86 248
use AOI21X1  _1286_
timestamp 0
transform 1 0 750 0 1 1690
box -6 -8 106 248
use OAI21X1  _1287_
timestamp 0
transform 1 0 1350 0 1 2650
box -6 -8 106 248
use INVX1  _1288_
timestamp 0
transform -1 0 1410 0 1 3130
box -6 -8 66 248
use NOR3X1  _1289_
timestamp 0
transform -1 0 2190 0 -1 2170
box -6 -8 186 248
use AOI21X1  _1290_
timestamp 0
transform 1 0 1870 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1291_
timestamp 0
transform 1 0 3770 0 1 3610
box -6 -8 86 248
use INVX1  _1292_
timestamp 0
transform 1 0 3530 0 1 3610
box -6 -8 66 248
use INVX1  _1293_
timestamp 0
transform 1 0 2690 0 1 4090
box -6 -8 66 248
use OAI21X1  _1294_
timestamp 0
transform -1 0 3570 0 -1 3130
box -6 -8 106 248
use NAND3X1  _1295_
timestamp 0
transform 1 0 3170 0 -1 3610
box -6 -8 106 248
use INVX1  _1296_
timestamp 0
transform 1 0 4150 0 -1 3610
box -6 -8 66 248
use AOI21X1  _1297_
timestamp 0
transform 1 0 3590 0 1 3130
box -6 -8 106 248
use OAI21X1  _1298_
timestamp 0
transform -1 0 4110 0 -1 3610
box -6 -8 106 248
use NAND3X1  _1299_
timestamp 0
transform -1 0 3410 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1300_
timestamp 0
transform -1 0 3130 0 -1 3610
box -6 -8 86 248
use NOR2X1  _1301_
timestamp 0
transform 1 0 3870 0 -1 3610
box -6 -8 86 248
use AND2X2  _1302_
timestamp 0
transform -1 0 3830 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1303_
timestamp 0
transform -1 0 3690 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1304_
timestamp 0
transform 1 0 2650 0 -1 3610
box -6 -8 86 248
use NAND3X1  _1305_
timestamp 0
transform -1 0 4490 0 1 4570
box -6 -8 106 248
use INVX1  _1306_
timestamp 0
transform 1 0 4130 0 1 4570
box -6 -8 66 248
use NAND3X1  _1307_
timestamp 0
transform -1 0 3870 0 -1 5050
box -6 -8 106 248
use NAND3X1  _1308_
timestamp 0
transform 1 0 3610 0 1 4090
box -6 -8 106 248
use OR2X2  _1309_
timestamp 0
transform 1 0 3510 0 -1 5050
box -6 -8 106 248
use INVX1  _1310_
timestamp 0
transform -1 0 3790 0 1 5530
box -6 -8 66 248
use OAI21X1  _1311_
timestamp 0
transform -1 0 3590 0 1 5050
box -6 -8 106 248
use AOI21X1  _1312_
timestamp 0
transform -1 0 3530 0 1 4570
box -6 -8 106 248
use NAND3X1  _1313_
timestamp 0
transform 1 0 3750 0 1 4090
box -6 -8 106 248
use AND2X2  _1314_
timestamp 0
transform -1 0 4330 0 1 4570
box -6 -8 106 248
use NAND3X1  _1315_
timestamp 0
transform 1 0 3990 0 1 4570
box -6 -8 106 248
use AOI21X1  _1316_
timestamp 0
transform -1 0 3810 0 1 4570
box -6 -8 106 248
use NAND3X1  _1317_
timestamp 0
transform 1 0 2730 0 1 4570
box -6 -8 106 248
use OAI22X1  _1318_
timestamp 0
transform 1 0 3010 0 1 4570
box -6 -8 126 248
use NAND3X1  _1319_
timestamp 0
transform 1 0 3850 0 1 4570
box -6 -8 106 248
use NAND3X1  _1320_
timestamp 0
transform -1 0 3670 0 1 4570
box -6 -8 106 248
use NOR2X1  _1321_
timestamp 0
transform -1 0 2950 0 1 4570
box -6 -8 86 248
use NAND3X1  _1322_
timestamp 0
transform -1 0 3390 0 1 4570
box -6 -8 106 248
use NAND2X1  _1323_
timestamp 0
transform 1 0 2410 0 1 3130
box -6 -8 86 248
use AOI21X1  _1324_
timestamp 0
transform -1 0 2450 0 -1 3130
box -6 -8 106 248
use OR2X2  _1325_
timestamp 0
transform -1 0 2890 0 -1 3130
box -6 -8 106 248
use INVX2  _1326_
timestamp 0
transform 1 0 4870 0 1 3610
box -6 -8 66 248
use OAI21X1  _1327_
timestamp 0
transform -1 0 2870 0 -1 3610
box -6 -8 106 248
use AOI21X1  _1328_
timestamp 0
transform -1 0 2770 0 1 3130
box -6 -8 106 248
use OAI21X1  _1329_
timestamp 0
transform -1 0 2630 0 1 3130
box -6 -8 106 248
use AOI21X1  _1330_
timestamp 0
transform -1 0 2470 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1331_
timestamp 0
transform 1 0 2230 0 -1 3610
box -6 -8 106 248
use AND2X2  _1332_
timestamp 0
transform -1 0 2610 0 -1 3610
box -6 -8 106 248
use AND2X2  _1333_
timestamp 0
transform -1 0 2270 0 1 2650
box -6 -8 106 248
use AND2X2  _1334_
timestamp 0
transform -1 0 2370 0 1 3130
box -6 -8 106 248
use OAI21X1  _1335_
timestamp 0
transform -1 0 2290 0 -1 3130
box -6 -8 106 248
use AOI21X1  _1336_
timestamp 0
transform -1 0 2590 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1337_
timestamp 0
transform -1 0 1970 0 1 3130
box -6 -8 86 248
use NAND3X1  _1338_
timestamp 0
transform -1 0 1890 0 -1 3610
box -6 -8 106 248
use NAND3X1  _1339_
timestamp 0
transform -1 0 1550 0 1 3130
box -6 -8 106 248
use AOI21X1  _1340_
timestamp 0
transform -1 0 1770 0 1 2170
box -6 -8 106 248
use OAI21X1  _1341_
timestamp 0
transform 1 0 1690 0 -1 2650
box -6 -8 106 248
use AOI21X1  _1342_
timestamp 0
transform -1 0 1830 0 1 3130
box -6 -8 106 248
use NAND2X1  _1343_
timestamp 0
transform 1 0 2150 0 1 3130
box -6 -8 86 248
use OAI21X1  _1344_
timestamp 0
transform -1 0 2150 0 -1 3130
box -6 -8 106 248
use AOI21X1  _1345_
timestamp 0
transform -1 0 2110 0 1 3130
box -6 -8 106 248
use OAI21X1  _1346_
timestamp 0
transform -1 0 1850 0 -1 3130
box -6 -8 106 248
use AOI21X1  _1347_
timestamp 0
transform 1 0 1210 0 1 3130
box -6 -8 106 248
use NAND3X1  _1348_
timestamp 0
transform -1 0 1690 0 1 3130
box -6 -8 106 248
use OAI21X1  _1349_
timestamp 0
transform 1 0 1890 0 -1 3130
box -6 -8 106 248
use AOI21X1  _1350_
timestamp 0
transform -1 0 1710 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1351_
timestamp 0
transform 1 0 1310 0 -1 3130
box -6 -8 106 248
use AOI21X1  _1352_
timestamp 0
transform -1 0 590 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1353_
timestamp 0
transform -1 0 430 0 1 1690
box -6 -8 106 248
use NAND3X1  _1354_
timestamp 0
transform -1 0 1550 0 -1 3130
box -6 -8 106 248
use NAND3X1  _1355_
timestamp 0
transform -1 0 1170 0 1 3130
box -6 -8 106 248
use NAND3X1  _1356_
timestamp 0
transform -1 0 1030 0 1 3130
box -6 -8 106 248
use NAND2X1  _1357_
timestamp 0
transform -1 0 890 0 1 3130
box -6 -8 86 248
use AOI21X1  _1358_
timestamp 0
transform 1 0 930 0 1 2650
box -6 -8 106 248
use OAI21X1  _1359_
timestamp 0
transform 1 0 770 0 -1 3130
box -6 -8 106 248
use AND2X2  _1360_
timestamp 0
transform 1 0 650 0 1 3130
box -6 -8 106 248
use OAI21X1  _1361_
timestamp 0
transform 1 0 910 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1362_
timestamp 0
transform 1 0 2030 0 1 2650
box -6 -8 106 248
use NAND2X1  _1363_
timestamp 0
transform -1 0 810 0 -1 3610
box -6 -8 86 248
use NAND2X1  _1364_
timestamp 0
transform -1 0 930 0 -1 3610
box -6 -8 86 248
use NAND2X1  _1365_
timestamp 0
transform -1 0 750 0 1 3610
box -6 -8 86 248
use OAI21X1  _1366_
timestamp 0
transform -1 0 630 0 1 3610
box -6 -8 106 248
use OAI21X1  _1367_
timestamp 0
transform -1 0 3550 0 -1 3610
box -6 -8 106 248
use INVX1  _1368_
timestamp 0
transform -1 0 1590 0 1 5050
box -6 -8 66 248
use AOI21X1  _1369_
timestamp 0
transform 1 0 1930 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1370_
timestamp 0
transform -1 0 2810 0 -1 5050
box -6 -8 86 248
use INVX1  _1371_
timestamp 0
transform 1 0 2850 0 -1 5050
box -6 -8 66 248
use NOR2X1  _1372_
timestamp 0
transform -1 0 3430 0 1 5050
box -6 -8 86 248
use INVX1  _1373_
timestamp 0
transform 1 0 4670 0 1 4570
box -6 -8 66 248
use NOR2X1  _1374_
timestamp 0
transform -1 0 3730 0 -1 5050
box -6 -8 86 248
use NAND2X1  _1375_
timestamp 0
transform 1 0 3630 0 1 5050
box -6 -8 86 248
use INVX1  _1376_
timestamp 0
transform -1 0 3310 0 1 5050
box -6 -8 66 248
use OAI21X1  _1377_
timestamp 0
transform -1 0 3330 0 -1 5050
box -6 -8 106 248
use AOI21X1  _1378_
timestamp 0
transform -1 0 3470 0 -1 5050
box -6 -8 106 248
use OAI21X1  _1379_
timestamp 0
transform -1 0 3190 0 -1 5050
box -6 -8 106 248
use NAND3X1  _1380_
timestamp 0
transform 1 0 2950 0 -1 5050
box -6 -8 106 248
use NOR2X1  _1381_
timestamp 0
transform 1 0 3110 0 1 5050
box -6 -8 86 248
use AND2X2  _1382_
timestamp 0
transform -1 0 3070 0 1 5050
box -6 -8 106 248
use OAI21X1  _1383_
timestamp 0
transform -1 0 2930 0 1 5050
box -6 -8 106 248
use NAND2X1  _1384_
timestamp 0
transform 1 0 2170 0 1 5050
box -6 -8 86 248
use NAND3X1  _1385_
timestamp 0
transform 1 0 4010 0 -1 5050
box -6 -8 106 248
use INVX1  _1386_
timestamp 0
transform 1 0 4450 0 1 5050
box -6 -8 66 248
use NAND3X1  _1387_
timestamp 0
transform 1 0 4150 0 -1 5050
box -6 -8 106 248
use NAND3X1  _1388_
timestamp 0
transform 1 0 4530 0 1 4570
box -6 -8 106 248
use OR2X2  _1389_
timestamp 0
transform 1 0 4450 0 -1 5050
box -6 -8 106 248
use INVX1  _1390_
timestamp 0
transform 1 0 5090 0 -1 5530
box -6 -8 66 248
use OAI21X1  _1391_
timestamp 0
transform -1 0 4810 0 -1 5050
box -6 -8 106 248
use NAND3X1  _1392_
timestamp 0
transform -1 0 4650 0 1 5050
box -6 -8 106 248
use NOR2X1  _1393_
timestamp 0
transform 1 0 4590 0 -1 5050
box -6 -8 86 248
use AND2X2  _1394_
timestamp 0
transform -1 0 4390 0 -1 5050
box -6 -8 106 248
use OAI21X1  _1395_
timestamp 0
transform -1 0 4250 0 1 5050
box -6 -8 106 248
use NAND2X1  _1396_
timestamp 0
transform -1 0 3970 0 1 5050
box -6 -8 86 248
use AOI21X1  _1397_
timestamp 0
transform -1 0 2530 0 1 5050
box -6 -8 106 248
use NAND3X1  _1398_
timestamp 0
transform -1 0 2390 0 1 5050
box -6 -8 106 248
use INVX1  _1399_
timestamp 0
transform 1 0 1910 0 1 5530
box -6 -8 66 248
use OAI21X1  _1400_
timestamp 0
transform -1 0 2110 0 1 5530
box -6 -8 106 248
use AND2X2  _1401_
timestamp 0
transform -1 0 2390 0 -1 5530
box -6 -8 106 248
use INVX1  _1402_
timestamp 0
transform -1 0 2250 0 -1 5530
box -6 -8 66 248
use NAND3X1  _1403_
timestamp 0
transform -1 0 1870 0 1 5530
box -6 -8 106 248
use NAND3X1  _1404_
timestamp 0
transform -1 0 1870 0 -1 5530
box -6 -8 106 248
use OAI21X1  _1405_
timestamp 0
transform -1 0 2170 0 -1 3610
box -6 -8 106 248
use AOI22X1  _1406_
timestamp 0
transform -1 0 2130 0 1 5050
box -6 -8 126 248
use INVX1  _1407_
timestamp 0
transform -1 0 2670 0 -1 5050
box -6 -8 66 248
use NAND3X1  _1408_
timestamp 0
transform -1 0 2570 0 -1 5050
box -6 -8 106 248
use INVX1  _1409_
timestamp 0
transform -1 0 2290 0 -1 5050
box -6 -8 66 248
use OAI21X1  _1410_
timestamp 0
transform -1 0 2430 0 -1 5050
box -6 -8 106 248
use AOI21X1  _1411_
timestamp 0
transform -1 0 2170 0 -1 5050
box -6 -8 106 248
use OAI21X1  _1412_
timestamp 0
transform -1 0 1730 0 1 5050
box -6 -8 106 248
use NAND3X1  _1413_
timestamp 0
transform -1 0 1590 0 -1 5530
box -6 -8 106 248
use NAND3X1  _1414_
timestamp 0
transform -1 0 1570 0 1 5530
box -6 -8 106 248
use OAI21X1  _1415_
timestamp 0
transform -1 0 1770 0 -1 5050
box -6 -8 106 248
use NAND3X1  _1416_
timestamp 0
transform -1 0 1630 0 -1 5050
box -6 -8 106 248
use NAND2X1  _1417_
timestamp 0
transform -1 0 1470 0 -1 5050
box -6 -8 86 248
use NAND3X1  _1418_
timestamp 0
transform -1 0 1470 0 -1 3610
box -6 -8 106 248
use AOI21X1  _1419_
timestamp 0
transform -1 0 1750 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1420_
timestamp 0
transform 1 0 1510 0 -1 3610
box -6 -8 106 248
use NAND3X1  _1421_
timestamp 0
transform 1 0 1570 0 1 4570
box -6 -8 106 248
use NAND2X1  _1422_
timestamp 0
transform 1 0 1370 0 -1 4090
box -6 -8 86 248
use INVX1  _1423_
timestamp 0
transform 1 0 1650 0 1 3610
box -6 -8 66 248
use NAND2X1  _1424_
timestamp 0
transform 1 0 1870 0 1 3610
box -6 -8 86 248
use OR2X2  _1425_
timestamp 0
transform 1 0 1990 0 1 3610
box -6 -8 106 248
use NAND2X1  _1426_
timestamp 0
transform 1 0 2130 0 1 3610
box -6 -8 86 248
use AND2X2  _1427_
timestamp 0
transform 1 0 3470 0 -1 2650
box -6 -8 106 248
use NOR2X1  _1428_
timestamp 0
transform 1 0 3390 0 1 2170
box -6 -8 86 248
use OAI21X1  _1429_
timestamp 0
transform 1 0 3530 0 1 2170
box -6 -8 106 248
use NOR2X1  _1430_
timestamp 0
transform 1 0 3090 0 1 1690
box -6 -8 86 248
use OAI21X1  _1431_
timestamp 0
transform -1 0 3090 0 1 1210
box -6 -8 106 248
use OAI21X1  _1432_
timestamp 0
transform -1 0 3050 0 1 1690
box -6 -8 106 248
use NAND2X1  _1433_
timestamp 0
transform -1 0 3070 0 -1 2170
box -6 -8 86 248
use OAI21X1  _1434_
timestamp 0
transform 1 0 2850 0 -1 2170
box -6 -8 106 248
use NOR3X1  _1435_
timestamp 0
transform -1 0 1970 0 1 5050
box -6 -8 186 248
use AOI21X1  _1436_
timestamp 0
transform 1 0 1810 0 -1 5050
box -6 -8 106 248
use OAI21X1  _1437_
timestamp 0
transform -1 0 2770 0 1 5050
box -6 -8 106 248
use INVX1  _1438_
timestamp 0
transform -1 0 2630 0 1 5050
box -6 -8 66 248
use AOI21X1  _1439_
timestamp 0
transform 1 0 2290 0 1 5530
box -6 -8 106 248
use NAND2X1  _1440_
timestamp 0
transform -1 0 3830 0 1 5050
box -6 -8 86 248
use INVX1  _1441_
timestamp 0
transform 1 0 4610 0 -1 5530
box -6 -8 66 248
use OAI21X1  _1442_
timestamp 0
transform 1 0 4310 0 1 5050
box -6 -8 106 248
use NAND3X1  _1443_
timestamp 0
transform 1 0 4010 0 1 5050
box -6 -8 106 248
use AOI21X1  _1444_
timestamp 0
transform 1 0 4690 0 1 5050
box -6 -8 106 248
use OAI21X1  _1445_
timestamp 0
transform 1 0 4710 0 -1 5530
box -6 -8 106 248
use NAND3X1  _1446_
timestamp 0
transform -1 0 4410 0 -1 5530
box -6 -8 106 248
use INVX1  _1447_
timestamp 0
transform 1 0 3830 0 1 5530
box -6 -8 66 248
use AOI21X1  _1448_
timestamp 0
transform 1 0 4470 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1449_
timestamp 0
transform -1 0 4330 0 -1 4570
box -6 -8 86 248
use NAND2X1  _1450_
timestamp 0
transform -1 0 4230 0 1 4090
box -6 -8 86 248
use OR2X2  _1451_
timestamp 0
transform 1 0 4410 0 1 4090
box -6 -8 106 248
use OAI21X1  _1452_
timestamp 0
transform -1 0 4470 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1453_
timestamp 0
transform 1 0 4510 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1454_
timestamp 0
transform 1 0 3930 0 1 5530
box -6 -8 106 248
use INVX1  _1455_
timestamp 0
transform -1 0 3690 0 1 5530
box -6 -8 66 248
use INVX1  _1456_
timestamp 0
transform 1 0 4070 0 1 5530
box -6 -8 66 248
use NAND3X1  _1457_
timestamp 0
transform -1 0 3570 0 1 5530
box -6 -8 106 248
use NAND3X1  _1458_
timestamp 0
transform -1 0 2830 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1459_
timestamp 0
transform 1 0 2830 0 1 5530
box -6 -8 86 248
use OAI21X1  _1460_
timestamp 0
transform 1 0 2430 0 -1 5530
box -6 -8 106 248
use NAND3X1  _1461_
timestamp 0
transform -1 0 2690 0 -1 5530
box -6 -8 106 248
use OAI21X1  _1462_
timestamp 0
transform 1 0 2150 0 1 5530
box -6 -8 106 248
use NAND3X1  _1463_
timestamp 0
transform -1 0 2790 0 1 5530
box -6 -8 106 248
use NAND2X1  _1464_
timestamp 0
transform -1 0 2510 0 1 5530
box -6 -8 86 248
use NAND3X1  _1465_
timestamp 0
transform -1 0 2650 0 1 5530
box -6 -8 106 248
use NAND2X1  _1466_
timestamp 0
transform 1 0 2050 0 -1 5530
box -6 -8 86 248
use NAND2X1  _1467_
timestamp 0
transform 1 0 1950 0 -1 5050
box -6 -8 86 248
use AOI21X1  _1468_
timestamp 0
transform -1 0 1730 0 1 5530
box -6 -8 106 248
use OAI21X1  _1469_
timestamp 0
transform 1 0 1630 0 -1 5530
box -6 -8 106 248
use NAND3X1  _1470_
timestamp 0
transform -1 0 2010 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1471_
timestamp 0
transform -1 0 1930 0 1 4570
box -6 -8 86 248
use NAND3X1  _1472_
timestamp 0
transform 1 0 1810 0 -1 4090
box -6 -8 106 248
use INVX1  _1473_
timestamp 0
transform -1 0 1550 0 -1 4090
box -6 -8 66 248
use NOR2X1  _1474_
timestamp 0
transform -1 0 1270 0 -1 3130
box -6 -8 86 248
use NAND2X1  _1475_
timestamp 0
transform 1 0 1110 0 1 3610
box -6 -8 86 248
use AOI21X1  _1476_
timestamp 0
transform 1 0 1370 0 1 3610
box -6 -8 106 248
use INVX1  _1477_
timestamp 0
transform -1 0 1770 0 -1 4090
box -6 -8 66 248
use OAI21X1  _1478_
timestamp 0
transform 1 0 1510 0 1 3610
box -6 -8 106 248
use NAND2X1  _1479_
timestamp 0
transform -1 0 1830 0 1 3610
box -6 -8 86 248
use NAND2X1  _1480_
timestamp 0
transform 1 0 1250 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1481_
timestamp 0
transform 1 0 2870 0 1 2650
box -6 -8 106 248
use AOI21X1  _1482_
timestamp 0
transform -1 0 2910 0 -1 2650
box -6 -8 106 248
use INVX1  _1483_
timestamp 0
transform 1 0 2390 0 1 730
box -6 -8 66 248
use OAI21X1  _1484_
timestamp 0
transform -1 0 3230 0 1 1210
box -6 -8 106 248
use AOI21X1  _1485_
timestamp 0
transform 1 0 2710 0 1 1210
box -6 -8 106 248
use OAI21X1  _1486_
timestamp 0
transform 1 0 2850 0 1 2170
box -6 -8 106 248
use OAI21X1  _1487_
timestamp 0
transform 1 0 2710 0 1 2170
box -6 -8 106 248
use OAI21X1  _1488_
timestamp 0
transform 1 0 2870 0 -1 5530
box -6 -8 106 248
use INVX1  _1489_
timestamp 0
transform 1 0 3010 0 -1 5530
box -6 -8 66 248
use NAND2X1  _1490_
timestamp 0
transform -1 0 4270 0 -1 5530
box -6 -8 86 248
use OAI21X1  _1491_
timestamp 0
transform -1 0 4150 0 -1 5530
box -6 -8 106 248
use INVX1  _1492_
timestamp 0
transform -1 0 3010 0 1 5530
box -6 -8 66 248
use NAND2X1  _1493_
timestamp 0
transform 1 0 4490 0 1 3610
box -6 -8 86 248
use NAND2X1  _1494_
timestamp 0
transform -1 0 4110 0 1 4090
box -6 -8 86 248
use OAI21X1  _1495_
timestamp 0
transform -1 0 4370 0 1 4090
box -6 -8 106 248
use OAI21X1  _1496_
timestamp 0
transform -1 0 4650 0 1 4090
box -6 -8 106 248
use OR2X2  _1497_
timestamp 0
transform 1 0 4610 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1498_
timestamp 0
transform 1 0 4470 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1499_
timestamp 0
transform -1 0 4830 0 -1 4090
box -6 -8 86 248
use OAI21X1  _1500_
timestamp 0
transform 1 0 4710 0 1 4090
box -6 -8 106 248
use INVX1  _1501_
timestamp 0
transform 1 0 4750 0 -1 4570
box -6 -8 66 248
use NAND2X1  _1502_
timestamp 0
transform 1 0 4850 0 -1 4570
box -6 -8 86 248
use INVX1  _1503_
timestamp 0
transform 1 0 5010 0 -1 4090
box -6 -8 66 248
use NAND3X1  _1504_
timestamp 0
transform 1 0 4870 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1505_
timestamp 0
transform -1 0 4710 0 -1 4570
box -6 -8 86 248
use NOR2X1  _1506_
timestamp 0
transform -1 0 3430 0 1 5530
box -6 -8 86 248
use AND2X2  _1507_
timestamp 0
transform -1 0 3310 0 1 5530
box -6 -8 106 248
use OAI21X1  _1508_
timestamp 0
transform -1 0 3150 0 1 5530
box -6 -8 106 248
use OR2X2  _1509_
timestamp 0
transform 1 0 3510 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1510_
timestamp 0
transform 1 0 3930 0 -1 5530
box -6 -8 86 248
use NAND3X1  _1511_
timestamp 0
transform -1 0 3750 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1512_
timestamp 0
transform 1 0 3390 0 -1 5530
box -6 -8 86 248
use NAND2X1  _1513_
timestamp 0
transform 1 0 3110 0 -1 5530
box -6 -8 86 248
use NAND3X1  _1514_
timestamp 0
transform 1 0 3250 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1515_
timestamp 0
transform -1 0 3250 0 1 4570
box -6 -8 86 248
use INVX1  _1516_
timestamp 0
transform -1 0 2770 0 -1 4570
box -6 -8 66 248
use NAND2X1  _1517_
timestamp 0
transform -1 0 1410 0 1 4090
box -6 -8 86 248
use OAI21X1  _1518_
timestamp 0
transform 1 0 1970 0 1 4570
box -6 -8 106 248
use OAI21X1  _1519_
timestamp 0
transform -1 0 1810 0 1 4570
box -6 -8 106 248
use AOI22X1  _1520_
timestamp 0
transform -1 0 1070 0 1 3610
box -6 -8 126 248
use OAI21X1  _1521_
timestamp 0
transform 1 0 790 0 1 3610
box -6 -8 106 248
use NAND3X1  _1522_
timestamp 0
transform -1 0 2530 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1523_
timestamp 0
transform 1 0 970 0 -1 3610
box -6 -8 106 248
use NOR2X1  _1524_
timestamp 0
transform -1 0 1670 0 -1 4090
box -6 -8 86 248
use AOI22X1  _1525_
timestamp 0
transform 1 0 1190 0 -1 4090
box -6 -8 126 248
use NAND3X1  _1526_
timestamp 0
transform 1 0 1230 0 1 3610
box -6 -8 106 248
use NAND3X1  _1527_
timestamp 0
transform 1 0 2810 0 1 4090
box -6 -8 106 248
use NAND2X1  _1528_
timestamp 0
transform 1 0 2950 0 1 4090
box -6 -8 86 248
use INVX1  _1529_
timestamp 0
transform 1 0 330 0 -1 3610
box -6 -8 66 248
use OAI21X1  _1530_
timestamp 0
transform 1 0 430 0 -1 3610
box -6 -8 106 248
use NAND3X1  _1531_
timestamp 0
transform 1 0 570 0 -1 3610
box -6 -8 106 248
use NOR2X1  _1532_
timestamp 0
transform 1 0 2810 0 -1 1210
box -6 -8 86 248
use OAI21X1  _1533_
timestamp 0
transform -1 0 2670 0 1 1210
box -6 -8 106 248
use OAI21X1  _1534_
timestamp 0
transform -1 0 2650 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1535_
timestamp 0
transform -1 0 2770 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1536_
timestamp 0
transform -1 0 3050 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1537_
timestamp 0
transform -1 0 130 0 1 3610
box -6 -8 86 248
use OAI21X1  _1538_
timestamp 0
transform -1 0 150 0 -1 3610
box -6 -8 106 248
use AOI21X1  _1539_
timestamp 0
transform 1 0 190 0 -1 3610
box -6 -8 106 248
use NOR2X1  _1540_
timestamp 0
transform 1 0 3250 0 -1 2170
box -6 -8 86 248
use AND2X2  _1541_
timestamp 0
transform -1 0 3470 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1542_
timestamp 0
transform 1 0 3050 0 -1 2650
box -6 -8 106 248
use AOI21X1  _1543_
timestamp 0
transform -1 0 3890 0 -1 5530
box -6 -8 106 248
use INVX1  _1544_
timestamp 0
transform 1 0 4970 0 1 4090
box -6 -8 66 248
use NOR2X1  _1545_
timestamp 0
transform 1 0 4850 0 1 4090
box -6 -8 86 248
use AOI21X1  _1546_
timestamp 0
transform 1 0 5090 0 1 4090
box -6 -8 106 248
use NAND2X1  _1547_
timestamp 0
transform 1 0 4210 0 -1 4090
box -6 -8 86 248
use OAI22X1  _1548_
timestamp 0
transform -1 0 4450 0 1 3610
box -6 -8 126 248
use OAI21X1  _1549_
timestamp 0
transform 1 0 4330 0 -1 4090
box -6 -8 106 248
use OR2X2  _1550_
timestamp 0
transform 1 0 5490 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1551_
timestamp 0
transform 1 0 4970 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1552_
timestamp 0
transform 1 0 5530 0 1 4570
box -6 -8 86 248
use NAND2X1  _1553_
timestamp 0
transform 1 0 5410 0 1 4570
box -6 -8 86 248
use INVX1  _1554_
timestamp 0
transform 1 0 5650 0 1 5530
box -6 -8 66 248
use NAND3X1  _1555_
timestamp 0
transform -1 0 5750 0 1 4570
box -6 -8 106 248
use NAND2X1  _1556_
timestamp 0
transform 1 0 5270 0 1 4570
box -6 -8 86 248
use NAND2X1  _1557_
timestamp 0
transform 1 0 3870 0 -1 4570
box -6 -8 86 248
use OR2X2  _1558_
timestamp 0
transform -1 0 3830 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1559_
timestamp 0
transform 1 0 3610 0 -1 4570
box -6 -8 86 248
use NAND3X1  _1560_
timestamp 0
transform -1 0 3030 0 -1 4570
box -6 -8 106 248
use INVX1  _1561_
timestamp 0
transform 1 0 3210 0 -1 4570
box -6 -8 66 248
use AOI21X1  _1562_
timestamp 0
transform 1 0 3210 0 1 4090
box -6 -8 106 248
use AND2X2  _1563_
timestamp 0
transform -1 0 3550 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1564_
timestamp 0
transform 1 0 3350 0 1 4090
box -6 -8 106 248
use NAND3X1  _1565_
timestamp 0
transform 1 0 3390 0 1 3610
box -6 -8 106 248
use NAND2X1  _1566_
timestamp 0
transform 1 0 3210 0 -1 2650
box -6 -8 86 248
use NAND2X1  _1567_
timestamp 0
transform 1 0 390 0 1 3130
box -6 -8 86 248
use AOI21X1  _1568_
timestamp 0
transform 1 0 510 0 1 3130
box -6 -8 106 248
use OAI21X1  _1569_
timestamp 0
transform 1 0 630 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1570_
timestamp 0
transform 1 0 3110 0 -1 2170
box -6 -8 86 248
use OAI21X1  _1571_
timestamp 0
transform 1 0 1970 0 -1 2650
box -6 -8 106 248
use NAND2X1  _1572_
timestamp 0
transform 1 0 3130 0 1 2170
box -6 -8 86 248
use NAND3X1  _1573_
timestamp 0
transform -1 0 3170 0 -1 4570
box -6 -8 106 248
use AOI21X1  _1574_
timestamp 0
transform 1 0 3070 0 1 4090
box -6 -8 106 248
use OAI21X1  _1575_
timestamp 0
transform 1 0 3310 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1576_
timestamp 0
transform 1 0 5230 0 1 4090
box -6 -8 106 248
use AOI21X1  _1577_
timestamp 0
transform -1 0 4170 0 -1 4090
box -6 -8 106 248
use OR2X2  _1578_
timestamp 0
transform -1 0 3750 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1579_
timestamp 0
transform 1 0 3810 0 -1 4090
box -6 -8 86 248
use NAND2X1  _1580_
timestamp 0
transform 1 0 3530 0 -1 4090
box -6 -8 86 248
use INVX1  _1581_
timestamp 0
transform -1 0 3350 0 -1 4090
box -6 -8 66 248
use OAI21X1  _1582_
timestamp 0
transform -1 0 3490 0 -1 4090
box -6 -8 106 248
use NOR2X1  _1583_
timestamp 0
transform -1 0 2890 0 -1 4570
box -6 -8 86 248
use NAND3X1  _1584_
timestamp 0
transform 1 0 2570 0 -1 4570
box -6 -8 106 248
use INVX1  _1585_
timestamp 0
transform 1 0 3510 0 1 4090
box -6 -8 66 248
use NAND3X1  _1586_
timestamp 0
transform -1 0 3250 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1587_
timestamp 0
transform 1 0 3670 0 1 2650
box -6 -8 106 248
use NAND2X1  _1588_
timestamp 0
transform 1 0 3670 0 1 2170
box -6 -8 86 248
use OAI21X1  _1589_
timestamp 0
transform -1 0 4030 0 -1 4090
box -6 -8 106 248
use NOR2X1  _1590_
timestamp 0
transform 1 0 3890 0 -1 2650
box -6 -8 86 248
use NOR2X1  _1591_
timestamp 0
transform 1 0 630 0 -1 2650
box -6 -8 86 248
use AOI21X1  _1592_
timestamp 0
transform 1 0 910 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1593_
timestamp 0
transform 1 0 750 0 -1 2650
box -6 -8 106 248
use AOI21X1  _1594_
timestamp 0
transform 1 0 3510 0 -1 2170
box -6 -8 106 248
use AOI22X1  _1595_
timestamp 0
transform 1 0 3730 0 -1 2650
box -6 -8 126 248
use INVX4  _1596_
timestamp 0
transform 1 0 5650 0 1 1690
box -6 -8 86 248
use INVX1  _1597_
timestamp 0
transform -1 0 5790 0 -1 1210
box -6 -8 66 248
use NAND2X1  _1598_
timestamp 0
transform -1 0 5710 0 1 3130
box -6 -8 86 248
use OAI21X1  _1599_
timestamp 0
transform 1 0 5610 0 1 2650
box -6 -8 106 248
use INVX1  _1600_
timestamp 0
transform -1 0 5650 0 -1 2170
box -6 -8 66 248
use NAND2X1  _1601_
timestamp 0
transform 1 0 5530 0 1 5530
box -6 -8 86 248
use OAI21X1  _1602_
timestamp 0
transform 1 0 5630 0 -1 3610
box -6 -8 106 248
use INVX1  _1603_
timestamp 0
transform 1 0 4930 0 1 2170
box -6 -8 66 248
use NAND2X1  _1604_
timestamp 0
transform 1 0 5130 0 1 2650
box -6 -8 86 248
use OAI21X1  _1605_
timestamp 0
transform 1 0 4990 0 1 2650
box -6 -8 106 248
use INVX1  _1606_
timestamp 0
transform -1 0 5190 0 1 3130
box -6 -8 66 248
use NAND2X1  _1607_
timestamp 0
transform -1 0 4950 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1608_
timestamp 0
transform -1 0 5090 0 1 3130
box -6 -8 106 248
use INVX1  _1609_
timestamp 0
transform 1 0 5350 0 1 3130
box -6 -8 66 248
use NAND2X1  _1610_
timestamp 0
transform -1 0 5590 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1611_
timestamp 0
transform 1 0 5470 0 1 3130
box -6 -8 106 248
use INVX1  _1612_
timestamp 0
transform -1 0 5630 0 -1 250
box -6 -8 66 248
use NAND2X1  _1613_
timestamp 0
transform -1 0 5650 0 1 5050
box -6 -8 86 248
use OAI21X1  _1614_
timestamp 0
transform -1 0 5730 0 -1 4570
box -6 -8 106 248
use INVX1  _1615_
timestamp 0
transform 1 0 5370 0 1 4090
box -6 -8 66 248
use NAND2X1  _1616_
timestamp 0
transform 1 0 5590 0 -1 5050
box -6 -8 86 248
use OAI21X1  _1617_
timestamp 0
transform 1 0 5470 0 1 4090
box -6 -8 106 248
use NAND2X1  _1618_
timestamp 0
transform 1 0 5590 0 -1 5530
box -6 -8 86 248
use OAI21X1  _1619_
timestamp 0
transform 1 0 5190 0 1 5050
box -6 -8 106 248
use NAND2X1  _1620_
timestamp 0
transform -1 0 5310 0 1 3130
box -6 -8 86 248
use OAI21X1  _1621_
timestamp 0
transform 1 0 4730 0 1 3130
box -6 -8 106 248
use NAND2X1  _1622_
timestamp 0
transform -1 0 4950 0 1 3130
box -6 -8 86 248
use OAI21X1  _1623_
timestamp 0
transform 1 0 4210 0 1 3130
box -6 -8 106 248
use NAND2X1  _1624_
timestamp 0
transform -1 0 4930 0 -1 3130
box -6 -8 86 248
use OAI21X1  _1625_
timestamp 0
transform 1 0 4570 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1626_
timestamp 0
transform 1 0 4510 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1627_
timestamp 0
transform 1 0 4250 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1628_
timestamp 0
transform 1 0 5150 0 1 4570
box -6 -8 86 248
use OAI21X1  _1629_
timestamp 0
transform 1 0 5010 0 1 4570
box -6 -8 106 248
use NAND2X1  _1630_
timestamp 0
transform 1 0 5170 0 1 5530
box -6 -8 86 248
use OAI21X1  _1631_
timestamp 0
transform -1 0 4530 0 1 5530
box -6 -8 106 248
use NAND2X1  _1632_
timestamp 0
transform 1 0 5710 0 -1 5530
box -6 -8 86 248
use OAI21X1  _1633_
timestamp 0
transform 1 0 5430 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1634_
timestamp 0
transform -1 0 5550 0 -1 5050
box -6 -8 86 248
use OAI21X1  _1635_
timestamp 0
transform 1 0 5090 0 -1 5050
box -6 -8 106 248
use NAND2X1  _1636_
timestamp 0
transform -1 0 5770 0 1 3610
box -6 -8 86 248
use OAI21X1  _1637_
timestamp 0
transform 1 0 5690 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1638_
timestamp 0
transform 1 0 5150 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1639_
timestamp 0
transform -1 0 5090 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1640_
timestamp 0
transform 1 0 4970 0 -1 3130
box -6 -8 86 248
use OAI21X1  _1641_
timestamp 0
transform 1 0 4710 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1642_
timestamp 0
transform -1 0 4470 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1643_
timestamp 0
transform 1 0 4350 0 1 3130
box -6 -8 106 248
use NAND2X1  _1644_
timestamp 0
transform -1 0 5070 0 1 3610
box -6 -8 86 248
use OAI21X1  _1645_
timestamp 0
transform 1 0 4730 0 1 3610
box -6 -8 106 248
use INVX1  _1646_
timestamp 0
transform -1 0 4870 0 1 5530
box -6 -8 66 248
use NAND2X1  _1647_
timestamp 0
transform -1 0 5130 0 1 5530
box -6 -8 86 248
use OAI21X1  _1648_
timestamp 0
transform -1 0 5010 0 1 5530
box -6 -8 106 248
use NAND2X1  _1649_
timestamp 0
transform 1 0 5690 0 1 5050
box -6 -8 86 248
use OAI21X1  _1650_
timestamp 0
transform 1 0 5430 0 1 5050
box -6 -8 106 248
use NAND2X1  _1651_
timestamp 0
transform 1 0 5730 0 -1 5050
box -6 -8 86 248
use OAI21X1  _1652_
timestamp 0
transform 1 0 5350 0 -1 4570
box -6 -8 106 248
use DFFPOSX1  _1653_
timestamp 0
transform -1 0 5570 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _1654_
timestamp 0
transform -1 0 5650 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _1655_
timestamp 0
transform 1 0 4930 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _1656_
timestamp 0
transform 1 0 5050 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _1657_
timestamp 0
transform -1 0 5770 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _1658_
timestamp 0
transform 1 0 5570 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _1659_
timestamp 0
transform -1 0 5410 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _1660_
timestamp 0
transform -1 0 5150 0 1 5050
box -6 -8 246 248
use DFFSR  _1661_
timestamp 0
transform -1 0 2230 0 -1 1690
box -6 -8 486 248
use DFFSR  _1662_
timestamp 0
transform -1 0 2530 0 1 2170
box -6 -8 486 248
use DFFSR  _1663_
timestamp 0
transform -1 0 2810 0 -1 2170
box -6 -8 486 248
use DFFSR  _1664_
timestamp 0
transform -1 0 2650 0 1 1690
box -6 -8 486 248
use DFFSR  _1665_
timestamp 0
transform 1 0 3050 0 -1 1690
box -6 -8 486 248
use DFFSR  _1666_
timestamp 0
transform 1 0 4450 0 -1 2650
box -6 -8 486 248
use DFFSR  _1667_
timestamp 0
transform -1 0 4350 0 1 2170
box -6 -8 486 248
use DFFSR  _1668_
timestamp 0
transform -1 0 4450 0 -1 2650
box -6 -8 486 248
use DFFPOSX1  _1669_
timestamp 0
transform -1 0 4690 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _1670_
timestamp 0
transform -1 0 4170 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _1671_
timestamp 0
transform -1 0 4690 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _1672_
timestamp 0
transform -1 0 4290 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _1673_
timestamp 0
transform -1 0 4970 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _1674_
timestamp 0
transform -1 0 4370 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _1675_
timestamp 0
transform -1 0 5390 0 -1 5530
box -6 -8 246 248
use DFFPOSX1  _1676_
timestamp 0
transform -1 0 5050 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _1677_
timestamp 0
transform -1 0 5650 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _1678_
timestamp 0
transform 1 0 5230 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1679_
timestamp 0
transform 1 0 4690 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _1680_
timestamp 0
transform 1 0 4270 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _1681_
timestamp 0
transform -1 0 4830 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1682_
timestamp 0
transform -1 0 5050 0 -1 5530
box -6 -8 246 248
use DFFPOSX1  _1683_
timestamp 0
transform -1 0 5430 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _1684_
timestamp 0
transform -1 0 5310 0 -1 4570
box -6 -8 246 248
use INVX1  _1685_
timestamp 0
transform 1 0 5090 0 -1 1210
box -6 -8 66 248
use INVX4  _1686_
timestamp 0
transform 1 0 5250 0 1 2650
box -6 -8 86 248
use OAI21X1  _1687_
timestamp 0
transform 1 0 5470 0 1 1210
box -6 -8 106 248
use NOR2X1  _1688_
timestamp 0
transform 1 0 5470 0 -1 1210
box -6 -8 86 248
use INVX1  _1689_
timestamp 0
transform -1 0 5410 0 1 730
box -6 -8 66 248
use INVX2  _1690_
timestamp 0
transform 1 0 5710 0 -1 2650
box -6 -8 66 248
use NAND2X1  _1691_
timestamp 0
transform 1 0 5370 0 -1 2170
box -6 -8 86 248
use INVX2  _1692_
timestamp 0
transform 1 0 5310 0 1 2170
box -6 -8 66 248
use NAND2X1  _1693_
timestamp 0
transform -1 0 4950 0 1 1690
box -6 -8 86 248
use NAND2X1  _1694_
timestamp 0
transform 1 0 5410 0 1 2170
box -6 -8 86 248
use AOI22X1  _1695_
timestamp 0
transform -1 0 5110 0 1 1690
box -6 -8 126 248
use INVX2  _1696_
timestamp 0
transform -1 0 5790 0 -1 1690
box -6 -8 66 248
use INVX1  _1697_
timestamp 0
transform 1 0 5530 0 1 2170
box -6 -8 66 248
use INVX1  _1698_
timestamp 0
transform 1 0 5490 0 -1 2170
box -6 -8 66 248
use OAI21X1  _1699_
timestamp 0
transform -1 0 5610 0 1 1690
box -6 -8 106 248
use NAND2X1  _1700_
timestamp 0
transform 1 0 5450 0 -1 1690
box -6 -8 86 248
use NAND2X1  _1701_
timestamp 0
transform 1 0 5670 0 -1 250
box -6 -8 86 248
use OAI21X1  _1702_
timestamp 0
transform 1 0 5630 0 1 1210
box -6 -8 106 248
use OAI21X1  _1703_
timestamp 0
transform -1 0 5010 0 1 730
box -6 -8 106 248
use AOI21X1  _1704_
timestamp 0
transform 1 0 5050 0 1 730
box -6 -8 106 248
use NOR2X1  _1705_
timestamp 0
transform 1 0 4970 0 1 1210
box -6 -8 86 248
use OAI21X1  _1706_
timestamp 0
transform 1 0 5370 0 -1 730
box -6 -8 106 248
use OAI21X1  _1707_
timestamp 0
transform -1 0 5610 0 -1 730
box -6 -8 106 248
use OR2X2  _1708_
timestamp 0
transform -1 0 5290 0 1 730
box -6 -8 106 248
use OAI21X1  _1709_
timestamp 0
transform -1 0 5430 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1710_
timestamp 0
transform -1 0 5270 0 -1 1210
box -6 -8 86 248
use INVX1  _1711_
timestamp 0
transform 1 0 4990 0 -1 1210
box -6 -8 66 248
use NOR2X1  _1712_
timestamp 0
transform 1 0 5650 0 -1 730
box -6 -8 86 248
use OAI21X1  _1713_
timestamp 0
transform -1 0 5330 0 -1 730
box -6 -8 106 248
use NAND2X1  _1714_
timestamp 0
transform -1 0 5290 0 1 1210
box -6 -8 86 248
use NAND3X1  _1715_
timestamp 0
transform 1 0 5150 0 -1 1690
box -6 -8 106 248
use AOI22X1  _1716_
timestamp 0
transform 1 0 5290 0 -1 1690
box -6 -8 126 248
use INVX1  _1717_
timestamp 0
transform -1 0 5210 0 1 1690
box -6 -8 66 248
use NOR2X1  _1718_
timestamp 0
transform -1 0 5330 0 1 1690
box -6 -8 86 248
use OAI21X1  _1719_
timestamp 0
transform 1 0 5370 0 1 1690
box -6 -8 106 248
use OAI21X1  _1720_
timestamp 0
transform -1 0 5430 0 1 1210
box -6 -8 106 248
use OAI21X1  _1721_
timestamp 0
transform 1 0 5570 0 1 250
box -6 -8 106 248
use AOI21X1  _1722_
timestamp 0
transform -1 0 5530 0 1 250
box -6 -8 106 248
use INVX1  _1723_
timestamp 0
transform 1 0 5470 0 -1 250
box -6 -8 66 248
use OAI21X1  _1724_
timestamp 0
transform 1 0 5290 0 1 5530
box -6 -8 106 248
use MUX2X1  _1725_
timestamp 0
transform 1 0 5310 0 -1 250
box -6 -8 126 248
use NAND2X1  _1726_
timestamp 0
transform -1 0 5270 0 -1 250
box -6 -8 86 248
use INVX1  _1727_
timestamp 0
transform 1 0 5430 0 1 5530
box -6 -8 66 248
use OAI21X1  _1728_
timestamp 0
transform 1 0 5630 0 1 730
box -6 -8 106 248
use MUX2X1  _1729_
timestamp 0
transform 1 0 5630 0 1 2170
box -6 -8 126 248
use OAI21X1  _1730_
timestamp 0
transform 1 0 5690 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1731_
timestamp 0
transform 1 0 5710 0 1 250
box -6 -8 86 248
use NAND3X1  _1732_
timestamp 0
transform 1 0 5570 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1733_
timestamp 0
transform -1 0 5690 0 -1 1210
box -6 -8 106 248
use AOI22X1  _1734_
timestamp 0
transform -1 0 5570 0 1 730
box -6 -8 126 248
use OAI21X1  _1735_
timestamp 0
transform 1 0 5270 0 1 250
box -6 -8 106 248
use OAI21X1  _1736_
timestamp 0
transform -1 0 5030 0 -1 250
box -6 -8 106 248
use NAND2X1  _1737_
timestamp 0
transform 1 0 4810 0 -1 250
box -6 -8 86 248
use NAND2X1  _1738_
timestamp 0
transform 1 0 4390 0 -1 250
box -6 -8 86 248
use INVX1  _1739_
timestamp 0
transform -1 0 3450 0 1 250
box -6 -8 66 248
use NOR2X1  _1740_
timestamp 0
transform 1 0 5070 0 -1 250
box -6 -8 86 248
use OAI21X1  _1741_
timestamp 0
transform -1 0 4770 0 -1 250
box -6 -8 106 248
use NAND2X1  _1742_
timestamp 0
transform 1 0 4730 0 -1 2170
box -6 -8 86 248
use INVX1  _1743_
timestamp 0
transform 1 0 5150 0 -1 2170
box -6 -8 66 248
use NOR2X1  _1744_
timestamp 0
transform 1 0 5250 0 -1 2170
box -6 -8 86 248
use NAND2X1  _1745_
timestamp 0
transform 1 0 5190 0 1 2170
box -6 -8 86 248
use AOI22X1  _1746_
timestamp 0
transform 1 0 5030 0 1 2170
box -6 -8 126 248
use OAI21X1  _1747_
timestamp 0
transform -1 0 5110 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1748_
timestamp 0
transform -1 0 4970 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1749_
timestamp 0
transform -1 0 4610 0 1 730
box -6 -8 106 248
use AOI21X1  _1750_
timestamp 0
transform 1 0 4650 0 1 730
box -6 -8 106 248
use INVX1  _1751_
timestamp 0
transform 1 0 4990 0 -1 730
box -6 -8 66 248
use OAI21X1  _1752_
timestamp 0
transform -1 0 5210 0 1 250
box -6 -8 106 248
use MUX2X1  _1753_
timestamp 0
transform 1 0 4950 0 1 250
box -6 -8 126 248
use NAND2X1  _1754_
timestamp 0
transform -1 0 4050 0 -1 250
box -6 -8 86 248
use OAI21X1  _1755_
timestamp 0
transform 1 0 4850 0 -1 730
box -6 -8 106 248
use OAI21X1  _1756_
timestamp 0
transform -1 0 4910 0 1 250
box -6 -8 106 248
use NAND3X1  _1757_
timestamp 0
transform -1 0 4610 0 -1 250
box -6 -8 106 248
use NAND2X1  _1758_
timestamp 0
transform -1 0 3690 0 -1 250
box -6 -8 86 248
use INVX1  _1759_
timestamp 0
transform -1 0 3330 0 1 1210
box -6 -8 66 248
use INVX1  _1760_
timestamp 0
transform -1 0 4770 0 1 250
box -6 -8 66 248
use AND2X2  _1761_
timestamp 0
transform 1 0 4110 0 -1 250
box -6 -8 106 248
use NAND2X1  _1762_
timestamp 0
transform 1 0 4610 0 -1 2170
box -6 -8 86 248
use AND2X2  _1763_
timestamp 0
transform 1 0 4390 0 1 2170
box -6 -8 106 248
use NAND2X1  _1764_
timestamp 0
transform 1 0 4690 0 1 2170
box -6 -8 86 248
use AOI22X1  _1765_
timestamp 0
transform 1 0 4530 0 1 2170
box -6 -8 126 248
use OAI21X1  _1766_
timestamp 0
transform -1 0 4430 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1767_
timestamp 0
transform 1 0 4470 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1768_
timestamp 0
transform -1 0 4550 0 -1 1210
box -6 -8 106 248
use AOI21X1  _1769_
timestamp 0
transform -1 0 4390 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1770_
timestamp 0
transform -1 0 4350 0 1 730
box -6 -8 106 248
use OAI21X1  _1771_
timestamp 0
transform -1 0 4210 0 1 730
box -6 -8 106 248
use INVX1  _1772_
timestamp 0
transform -1 0 4410 0 1 250
box -6 -8 66 248
use OAI21X1  _1773_
timestamp 0
transform -1 0 4670 0 1 250
box -6 -8 106 248
use NAND3X1  _1774_
timestamp 0
transform -1 0 4170 0 1 250
box -6 -8 106 248
use NAND2X1  _1775_
timestamp 0
transform 1 0 3930 0 1 250
box -6 -8 86 248
use INVX1  _1776_
timestamp 0
transform -1 0 3950 0 1 1210
box -6 -8 66 248
use INVX1  _1777_
timestamp 0
transform -1 0 3170 0 1 730
box -6 -8 66 248
use AOI21X1  _1778_
timestamp 0
transform 1 0 3650 0 1 250
box -6 -8 106 248
use NAND3X1  _1779_
timestamp 0
transform -1 0 3890 0 1 250
box -6 -8 106 248
use NAND2X1  _1780_
timestamp 0
transform -1 0 4530 0 1 250
box -6 -8 86 248
use INVX1  _1781_
timestamp 0
transform 1 0 4410 0 1 730
box -6 -8 66 248
use AOI21X1  _1782_
timestamp 0
transform -1 0 4510 0 -1 730
box -6 -8 106 248
use NAND2X1  _1783_
timestamp 0
transform -1 0 4150 0 1 1690
box -6 -8 86 248
use AND2X2  _1784_
timestamp 0
transform -1 0 4070 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1785_
timestamp 0
transform 1 0 4110 0 -1 1690
box -6 -8 86 248
use AOI22X1  _1786_
timestamp 0
transform -1 0 4350 0 -1 1690
box -6 -8 126 248
use OAI21X1  _1787_
timestamp 0
transform -1 0 3890 0 1 1690
box -6 -8 106 248
use OAI21X1  _1788_
timestamp 0
transform 1 0 3930 0 1 1690
box -6 -8 106 248
use OAI21X1  _1789_
timestamp 0
transform -1 0 4510 0 1 1210
box -6 -8 106 248
use AOI21X1  _1790_
timestamp 0
transform -1 0 4370 0 1 1210
box -6 -8 106 248
use OAI21X1  _1791_
timestamp 0
transform -1 0 4230 0 1 1210
box -6 -8 106 248
use OAI21X1  _1792_
timestamp 0
transform -1 0 4090 0 1 1210
box -6 -8 106 248
use AOI21X1  _1793_
timestamp 0
transform 1 0 4010 0 -1 730
box -6 -8 106 248
use NOR2X1  _1794_
timestamp 0
transform -1 0 4350 0 -1 250
box -6 -8 86 248
use OAI21X1  _1795_
timestamp 0
transform -1 0 4310 0 1 250
box -6 -8 106 248
use NAND2X1  _1796_
timestamp 0
transform 1 0 3990 0 1 730
box -6 -8 86 248
use OAI21X1  _1797_
timestamp 0
transform -1 0 3950 0 1 730
box -6 -8 106 248
use INVX1  _1798_
timestamp 0
transform -1 0 3810 0 1 730
box -6 -8 66 248
use NOR2X1  _1799_
timestamp 0
transform -1 0 3570 0 1 730
box -6 -8 86 248
use NOR2X1  _1800_
timestamp 0
transform -1 0 3450 0 1 730
box -6 -8 86 248
use INVX1  _1801_
timestamp 0
transform 1 0 4190 0 -1 1210
box -6 -8 66 248
use NAND2X1  _1802_
timestamp 0
transform 1 0 4710 0 1 1210
box -6 -8 86 248
use AND2X2  _1803_
timestamp 0
transform -1 0 4710 0 1 1690
box -6 -8 106 248
use NAND2X1  _1804_
timestamp 0
transform -1 0 4430 0 1 1690
box -6 -8 86 248
use AOI22X1  _1805_
timestamp 0
transform -1 0 4510 0 -1 1690
box -6 -8 126 248
use OAI21X1  _1806_
timestamp 0
transform 1 0 4470 0 1 1690
box -6 -8 106 248
use OAI21X1  _1807_
timestamp 0
transform 1 0 4570 0 1 1210
box -6 -8 106 248
use OAI21X1  _1808_
timestamp 0
transform 1 0 4730 0 -1 1210
box -6 -8 106 248
use AOI21X1  _1809_
timestamp 0
transform -1 0 4690 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1810_
timestamp 0
transform -1 0 4790 0 -1 730
box -6 -8 106 248
use OAI21X1  _1811_
timestamp 0
transform -1 0 4650 0 -1 730
box -6 -8 106 248
use INVX1  _1812_
timestamp 0
transform -1 0 4370 0 -1 730
box -6 -8 66 248
use OAI21X1  _1813_
timestamp 0
transform 1 0 4170 0 -1 730
box -6 -8 106 248
use AOI21X1  _1814_
timestamp 0
transform -1 0 3710 0 1 730
box -6 -8 106 248
use NAND2X1  _1815_
timestamp 0
transform 1 0 3610 0 -1 730
box -6 -8 86 248
use NAND2X1  _1816_
timestamp 0
transform 1 0 3350 0 -1 730
box -6 -8 86 248
use INVX1  _1817_
timestamp 0
transform 1 0 3370 0 1 1210
box -6 -8 66 248
use OAI21X1  _1818_
timestamp 0
transform -1 0 3570 0 -1 730
box -6 -8 106 248
use INVX1  _1819_
timestamp 0
transform -1 0 3430 0 1 1690
box -6 -8 66 248
use AND2X2  _1820_
timestamp 0
transform -1 0 4170 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1821_
timestamp 0
transform -1 0 4290 0 -1 2170
box -6 -8 86 248
use AOI22X1  _1822_
timestamp 0
transform -1 0 4310 0 1 1690
box -6 -8 126 248
use OAI21X1  _1823_
timestamp 0
transform -1 0 3730 0 1 1690
box -6 -8 106 248
use OAI22X1  _1824_
timestamp 0
transform 1 0 3470 0 1 1690
box -6 -8 126 248
use OAI21X1  _1825_
timestamp 0
transform 1 0 3750 0 1 1210
box -6 -8 106 248
use AOI21X1  _1826_
timestamp 0
transform -1 0 3710 0 1 1210
box -6 -8 106 248
use OAI21X1  _1827_
timestamp 0
transform -1 0 3790 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1828_
timestamp 0
transform -1 0 3650 0 -1 1210
box -6 -8 106 248
use INVX1  _1829_
timestamp 0
transform -1 0 2830 0 1 250
box -6 -8 66 248
use NAND2X1  _1830_
timestamp 0
transform -1 0 2650 0 -1 730
box -6 -8 86 248
use NAND3X1  _1831_
timestamp 0
transform -1 0 3310 0 -1 730
box -6 -8 106 248
use NAND2X1  _1832_
timestamp 0
transform -1 0 3030 0 -1 730
box -6 -8 86 248
use INVX1  _1833_
timestamp 0
transform 1 0 3010 0 1 730
box -6 -8 66 248
use INVX1  _1834_
timestamp 0
transform -1 0 2450 0 1 250
box -6 -8 66 248
use AOI21X1  _1835_
timestamp 0
transform -1 0 3190 0 1 250
box -6 -8 106 248
use NAND2X1  _1836_
timestamp 0
transform 1 0 5090 0 1 1210
box -6 -8 86 248
use AND2X2  _1837_
timestamp 0
transform -1 0 5090 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1838_
timestamp 0
transform 1 0 4730 0 -1 1690
box -6 -8 86 248
use AOI22X1  _1839_
timestamp 0
transform 1 0 4570 0 -1 1690
box -6 -8 126 248
use OAI21X1  _1840_
timestamp 0
transform 1 0 4850 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1841_
timestamp 0
transform 1 0 4830 0 1 1210
box -6 -8 106 248
use OAI21X1  _1842_
timestamp 0
transform 1 0 3710 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1843_
timestamp 0
transform -1 0 3670 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1844_
timestamp 0
transform 1 0 3870 0 -1 730
box -6 -8 106 248
use OAI21X1  _1845_
timestamp 0
transform -1 0 3830 0 -1 730
box -6 -8 106 248
use INVX1  _1846_
timestamp 0
transform 1 0 2010 0 1 250
box -6 -8 66 248
use OAI21X1  _1847_
timestamp 0
transform -1 0 2210 0 1 250
box -6 -8 106 248
use NAND3X1  _1848_
timestamp 0
transform -1 0 2590 0 1 250
box -6 -8 106 248
use AND2X2  _1849_
timestamp 0
transform 1 0 2450 0 -1 250
box -6 -8 106 248
use NOR2X1  _1850_
timestamp 0
transform 1 0 4070 0 -1 1210
box -6 -8 86 248
use NAND2X1  _1851_
timestamp 0
transform 1 0 3950 0 -1 1210
box -6 -8 86 248
use NOR2X1  _1852_
timestamp 0
transform -1 0 3410 0 -1 1210
box -6 -8 86 248
use NOR2X1  _1853_
timestamp 0
transform -1 0 2770 0 -1 730
box -6 -8 86 248
use OAI21X1  _1854_
timestamp 0
transform 1 0 2810 0 -1 730
box -6 -8 106 248
use NOR2X1  _1855_
timestamp 0
transform 1 0 2930 0 -1 1210
box -6 -8 86 248
use AND2X2  _1856_
timestamp 0
transform 1 0 3050 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1857_
timestamp 0
transform -1 0 2410 0 -1 250
box -6 -8 86 248
use NAND2X1  _1858_
timestamp 0
transform -1 0 2950 0 1 730
box -6 -8 86 248
use OAI21X1  _1859_
timestamp 0
transform 1 0 3510 0 1 250
box -6 -8 106 248
use INVX1  _1860_
timestamp 0
transform -1 0 3330 0 -1 250
box -6 -8 66 248
use NOR2X1  _1861_
timestamp 0
transform -1 0 2950 0 1 250
box -6 -8 86 248
use NAND2X1  _1862_
timestamp 0
transform -1 0 3090 0 -1 250
box -6 -8 86 248
use NOR2X1  _1863_
timestamp 0
transform -1 0 4830 0 1 1690
box -6 -8 86 248
use NAND3X1  _1864_
timestamp 0
transform -1 0 3230 0 -1 250
box -6 -8 106 248
use INVX1  _1865_
timestamp 0
transform 1 0 2990 0 1 250
box -6 -8 66 248
use AOI21X1  _1866_
timestamp 0
transform 1 0 3250 0 1 250
box -6 -8 106 248
use INVX1  _1867_
timestamp 0
transform -1 0 3570 0 -1 250
box -6 -8 66 248
use OAI21X1  _1868_
timestamp 0
transform 1 0 3370 0 -1 250
box -6 -8 106 248
use AND2X2  _1869_
timestamp 0
transform -1 0 2830 0 -1 250
box -6 -8 106 248
use OAI21X1  _1870_
timestamp 0
transform 1 0 2630 0 1 250
box -6 -8 106 248
use AOI21X1  _1871_
timestamp 0
transform 1 0 3070 0 -1 730
box -6 -8 106 248
use NAND2X1  _1872_
timestamp 0
transform 1 0 2890 0 -1 250
box -6 -8 86 248
use AOI21X1  _1873_
timestamp 0
transform -1 0 2690 0 -1 250
box -6 -8 106 248
use AOI21X1  _1874_
timestamp 0
transform -1 0 2350 0 1 250
box -6 -8 106 248
use NOR2X1  _1875_
timestamp 0
transform 1 0 1870 0 1 250
box -6 -8 86 248
use AND2X2  _1876_
timestamp 0
transform -1 0 1830 0 1 250
box -6 -8 106 248
use INVX1  _1877_
timestamp 0
transform -1 0 3510 0 -1 1210
box -6 -8 66 248
use NAND2X1  _1878_
timestamp 0
transform 1 0 3830 0 -1 1210
box -6 -8 86 248
use NAND2X1  _1879_
timestamp 0
transform -1 0 3310 0 1 730
box -6 -8 86 248
use NAND2X1  _1880_
timestamp 0
transform 1 0 2750 0 1 730
box -6 -8 86 248
use OR2X2  _1881_
timestamp 0
transform -1 0 2710 0 1 730
box -6 -8 106 248
use NAND2X1  _1882_
timestamp 0
transform -1 0 2570 0 1 730
box -6 -8 86 248
use INVX1  _1883_
timestamp 0
transform -1 0 1610 0 -1 250
box -6 -8 66 248
use OAI21X1  _1884_
timestamp 0
transform -1 0 1750 0 -1 250
box -6 -8 106 248
use NAND3X1  _1885_
timestamp 0
transform -1 0 2170 0 -1 250
box -6 -8 106 248
use NAND3X1  _1886_
timestamp 0
transform 1 0 1910 0 -1 250
box -6 -8 106 248
use NAND2X1  _1887_
timestamp 0
transform -1 0 1870 0 -1 250
box -6 -8 86 248
use NAND2X1  _1888_
timestamp 0
transform 1 0 2450 0 -1 730
box -6 -8 86 248
use AND2X2  _1889_
timestamp 0
transform 1 0 2310 0 -1 730
box -6 -8 106 248
use BUFX2  _1890_
timestamp 0
transform -1 0 1470 0 -1 1690
box -6 -8 86 248
use BUFX2  _1891_
timestamp 0
transform -1 0 130 0 1 2170
box -6 -8 86 248
use BUFX2  _1892_
timestamp 0
transform -1 0 150 0 -1 2170
box -6 -8 86 248
use BUFX2  _1893_
timestamp 0
transform 1 0 2210 0 -1 250
box -6 -8 86 248
use BUFX2  _1894_
timestamp 0
transform -1 0 3550 0 1 1210
box -6 -8 86 248
use BUFX2  _1895_
timestamp 0
transform -1 0 3810 0 -1 250
box -6 -8 86 248
use BUFX2  _1896_
timestamp 0
transform -1 0 3930 0 -1 1690
box -6 -8 86 248
use BUFX2  _1897_
timestamp 0
transform 1 0 3850 0 -1 250
box -6 -8 86 248
use BUFX2  BUFX2_insert5
timestamp 0
transform 1 0 3790 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert6
timestamp 0
transform -1 0 2330 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert7
timestamp 0
transform -1 0 4070 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert8
timestamp 0
transform -1 0 3010 0 -1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert9
timestamp 0
transform -1 0 2650 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert10
timestamp 0
transform -1 0 2690 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert11
timestamp 0
transform 1 0 4870 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert12
timestamp 0
transform -1 0 4890 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert13
timestamp 0
transform -1 0 4870 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert14
timestamp 0
transform 1 0 5110 0 -1 730
box -6 -8 86 248
use CLKBUF1  CLKBUF1_insert0
timestamp 0
transform -1 0 5410 0 -1 2650
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert1
timestamp 0
transform 1 0 5470 0 -1 2650
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert2
timestamp 0
transform -1 0 5410 0 1 3610
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert3
timestamp 0
transform -1 0 4770 0 1 5530
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert4
timestamp 0
transform -1 0 5530 0 -1 3130
box -6 -8 206 248
use FILL  FILL85650x39750
timestamp 0
transform 1 0 5710 0 1 2650
box -6 -8 26 248
use FILL  FILL85650x46950
timestamp 0
transform 1 0 5710 0 1 3130
box -6 -8 26 248
use FILL  FILL85650x82950
timestamp 0
transform 1 0 5710 0 1 5530
box -6 -8 26 248
use FILL  FILL85950x7350
timestamp 0
transform -1 0 5750 0 -1 730
box -6 -8 26 248
use FILL  FILL85950x10950
timestamp 0
transform 1 0 5730 0 1 730
box -6 -8 26 248
use FILL  FILL85950x18150
timestamp 0
transform 1 0 5730 0 1 1210
box -6 -8 26 248
use FILL  FILL85950x25350
timestamp 0
transform 1 0 5730 0 1 1690
box -6 -8 26 248
use FILL  FILL85950x39750
timestamp 0
transform 1 0 5730 0 1 2650
box -6 -8 26 248
use FILL  FILL85950x46950
timestamp 0
transform 1 0 5730 0 1 3130
box -6 -8 26 248
use FILL  FILL85950x50550
timestamp 0
transform -1 0 5750 0 -1 3610
box -6 -8 26 248
use FILL  FILL85950x64950
timestamp 0
transform -1 0 5750 0 -1 4570
box -6 -8 26 248
use FILL  FILL85950x82950
timestamp 0
transform 1 0 5730 0 1 5530
box -6 -8 26 248
use FILL  FILL86250x150
timestamp 0
transform -1 0 5770 0 -1 250
box -6 -8 26 248
use FILL  FILL86250x7350
timestamp 0
transform -1 0 5770 0 -1 730
box -6 -8 26 248
use FILL  FILL86250x10950
timestamp 0
transform 1 0 5750 0 1 730
box -6 -8 26 248
use FILL  FILL86250x18150
timestamp 0
transform 1 0 5750 0 1 1210
box -6 -8 26 248
use FILL  FILL86250x25350
timestamp 0
transform 1 0 5750 0 1 1690
box -6 -8 26 248
use FILL  FILL86250x32550
timestamp 0
transform 1 0 5750 0 1 2170
box -6 -8 26 248
use FILL  FILL86250x39750
timestamp 0
transform 1 0 5750 0 1 2650
box -6 -8 26 248
use FILL  FILL86250x46950
timestamp 0
transform 1 0 5750 0 1 3130
box -6 -8 26 248
use FILL  FILL86250x50550
timestamp 0
transform -1 0 5770 0 -1 3610
box -6 -8 26 248
use FILL  FILL86250x64950
timestamp 0
transform -1 0 5770 0 -1 4570
box -6 -8 26 248
use FILL  FILL86250x68550
timestamp 0
transform 1 0 5750 0 1 4570
box -6 -8 26 248
use FILL  FILL86250x82950
timestamp 0
transform 1 0 5750 0 1 5530
box -6 -8 26 248
use FILL  FILL86550x150
timestamp 0
transform -1 0 5790 0 -1 250
box -6 -8 26 248
use FILL  FILL86550x7350
timestamp 0
transform -1 0 5790 0 -1 730
box -6 -8 26 248
use FILL  FILL86550x10950
timestamp 0
transform 1 0 5770 0 1 730
box -6 -8 26 248
use FILL  FILL86550x18150
timestamp 0
transform 1 0 5770 0 1 1210
box -6 -8 26 248
use FILL  FILL86550x25350
timestamp 0
transform 1 0 5770 0 1 1690
box -6 -8 26 248
use FILL  FILL86550x32550
timestamp 0
transform 1 0 5770 0 1 2170
box -6 -8 26 248
use FILL  FILL86550x36150
timestamp 0
transform -1 0 5790 0 -1 2650
box -6 -8 26 248
use FILL  FILL86550x39750
timestamp 0
transform 1 0 5770 0 1 2650
box -6 -8 26 248
use FILL  FILL86550x43350
timestamp 0
transform -1 0 5790 0 -1 3130
box -6 -8 26 248
use FILL  FILL86550x46950
timestamp 0
transform 1 0 5770 0 1 3130
box -6 -8 26 248
use FILL  FILL86550x50550
timestamp 0
transform -1 0 5790 0 -1 3610
box -6 -8 26 248
use FILL  FILL86550x54150
timestamp 0
transform 1 0 5770 0 1 3610
box -6 -8 26 248
use FILL  FILL86550x64950
timestamp 0
transform -1 0 5790 0 -1 4570
box -6 -8 26 248
use FILL  FILL86550x68550
timestamp 0
transform 1 0 5770 0 1 4570
box -6 -8 26 248
use FILL  FILL86550x75750
timestamp 0
transform 1 0 5770 0 1 5050
box -6 -8 26 248
use FILL  FILL86550x82950
timestamp 0
transform 1 0 5770 0 1 5530
box -6 -8 26 248
use FILL  FILL86850x150
timestamp 0
transform -1 0 5810 0 -1 250
box -6 -8 26 248
use FILL  FILL86850x3750
timestamp 0
transform 1 0 5790 0 1 250
box -6 -8 26 248
use FILL  FILL86850x7350
timestamp 0
transform -1 0 5810 0 -1 730
box -6 -8 26 248
use FILL  FILL86850x10950
timestamp 0
transform 1 0 5790 0 1 730
box -6 -8 26 248
use FILL  FILL86850x14550
timestamp 0
transform -1 0 5810 0 -1 1210
box -6 -8 26 248
use FILL  FILL86850x18150
timestamp 0
transform 1 0 5790 0 1 1210
box -6 -8 26 248
use FILL  FILL86850x21750
timestamp 0
transform -1 0 5810 0 -1 1690
box -6 -8 26 248
use FILL  FILL86850x25350
timestamp 0
transform 1 0 5790 0 1 1690
box -6 -8 26 248
use FILL  FILL86850x28950
timestamp 0
transform -1 0 5810 0 -1 2170
box -6 -8 26 248
use FILL  FILL86850x32550
timestamp 0
transform 1 0 5790 0 1 2170
box -6 -8 26 248
use FILL  FILL86850x36150
timestamp 0
transform -1 0 5810 0 -1 2650
box -6 -8 26 248
use FILL  FILL86850x39750
timestamp 0
transform 1 0 5790 0 1 2650
box -6 -8 26 248
use FILL  FILL86850x43350
timestamp 0
transform -1 0 5810 0 -1 3130
box -6 -8 26 248
use FILL  FILL86850x46950
timestamp 0
transform 1 0 5790 0 1 3130
box -6 -8 26 248
use FILL  FILL86850x50550
timestamp 0
transform -1 0 5810 0 -1 3610
box -6 -8 26 248
use FILL  FILL86850x54150
timestamp 0
transform 1 0 5790 0 1 3610
box -6 -8 26 248
use FILL  FILL86850x57750
timestamp 0
transform -1 0 5810 0 -1 4090
box -6 -8 26 248
use FILL  FILL86850x64950
timestamp 0
transform -1 0 5810 0 -1 4570
box -6 -8 26 248
use FILL  FILL86850x68550
timestamp 0
transform 1 0 5790 0 1 4570
box -6 -8 26 248
use FILL  FILL86850x75750
timestamp 0
transform 1 0 5790 0 1 5050
box -6 -8 26 248
use FILL  FILL86850x79350
timestamp 0
transform -1 0 5810 0 -1 5530
box -6 -8 26 248
use FILL  FILL86850x82950
timestamp 0
transform 1 0 5790 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__920_
timestamp 0
transform -1 0 3630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__921_
timestamp 0
transform 1 0 4070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__922_
timestamp 0
transform -1 0 3870 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__923_
timestamp 0
transform -1 0 3890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__924_
timestamp 0
transform 1 0 4250 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__925_
timestamp 0
transform -1 0 3610 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__926_
timestamp 0
transform 1 0 2330 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__927_
timestamp 0
transform -1 0 1150 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__928_
timestamp 0
transform 1 0 2210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__929_
timestamp 0
transform 1 0 2070 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__930_
timestamp 0
transform -1 0 2230 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__931_
timestamp 0
transform -1 0 990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__932_
timestamp 0
transform -1 0 1730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__933_
timestamp 0
transform 1 0 3890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__934_
timestamp 0
transform -1 0 2510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__935_
timestamp 0
transform -1 0 2370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__936_
timestamp 0
transform 1 0 1430 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__937_
timestamp 0
transform -1 0 1170 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__938_
timestamp 0
transform -1 0 2090 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__939_
timestamp 0
transform 1 0 1090 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__940_
timestamp 0
transform -1 0 2510 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__941_
timestamp 0
transform -1 0 1810 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__942_
timestamp 0
transform -1 0 1550 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__943_
timestamp 0
transform -1 0 1070 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__944_
timestamp 0
transform 1 0 2410 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__945_
timestamp 0
transform 1 0 2490 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__946_
timestamp 0
transform -1 0 2350 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__947_
timestamp 0
transform -1 0 970 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__948_
timestamp 0
transform -1 0 1270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__949_
timestamp 0
transform -1 0 850 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__950_
timestamp 0
transform 1 0 810 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__951_
timestamp 0
transform -1 0 3970 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__952_
timestamp 0
transform 1 0 2450 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__953_
timestamp 0
transform -1 0 1350 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__954_
timestamp 0
transform -1 0 750 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__955_
timestamp 0
transform -1 0 690 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__956_
timestamp 0
transform 1 0 750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__957_
timestamp 0
transform -1 0 710 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__958_
timestamp 0
transform 1 0 1930 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__959_
timestamp 0
transform -1 0 2070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__960_
timestamp 0
transform -1 0 630 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__961_
timestamp 0
transform -1 0 5090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__962_
timestamp 0
transform 1 0 2610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__963_
timestamp 0
transform -1 0 1930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__964_
timestamp 0
transform -1 0 1670 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__965_
timestamp 0
transform -1 0 30 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__966_
timestamp 0
transform -1 0 330 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__967_
timestamp 0
transform -1 0 550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__968_
timestamp 0
transform -1 0 290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__969_
timestamp 0
transform -1 0 190 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__970_
timestamp 0
transform -1 0 170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__971_
timestamp 0
transform -1 0 990 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__972_
timestamp 0
transform -1 0 30 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__973_
timestamp 0
transform -1 0 490 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__974_
timestamp 0
transform -1 0 170 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__975_
timestamp 0
transform 1 0 4130 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__976_
timestamp 0
transform -1 0 3910 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__977_
timestamp 0
transform -1 0 1610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__978_
timestamp 0
transform 1 0 850 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__979_
timestamp 0
transform -1 0 2130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__980_
timestamp 0
transform -1 0 1990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__981_
timestamp 0
transform -1 0 1870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__982_
timestamp 0
transform 1 0 1450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__983_
timestamp 0
transform 1 0 730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__984_
timestamp 0
transform -1 0 610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__985_
timestamp 0
transform 1 0 950 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__986_
timestamp 0
transform -1 0 710 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__987_
timestamp 0
transform -1 0 590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__988_
timestamp 0
transform -1 0 170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__989_
timestamp 0
transform 1 0 290 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__990_
timestamp 0
transform 1 0 290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__991_
timestamp 0
transform -1 0 570 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__992_
timestamp 0
transform -1 0 450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__993_
timestamp 0
transform 1 0 430 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__994_
timestamp 0
transform -1 0 30 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__995_
timestamp 0
transform -1 0 30 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__996_
timestamp 0
transform 1 0 150 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__997_
timestamp 0
transform -1 0 30 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__998_
timestamp 0
transform -1 0 30 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__999_
timestamp 0
transform 1 0 370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1000_
timestamp 0
transform -1 0 1810 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1001_
timestamp 0
transform -1 0 2110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1002_
timestamp 0
transform 1 0 1250 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1003_
timestamp 0
transform 1 0 1370 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1004_
timestamp 0
transform -1 0 1650 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1005_
timestamp 0
transform 1 0 870 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1006_
timestamp 0
transform 1 0 590 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1007_
timestamp 0
transform -1 0 1170 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1008_
timestamp 0
transform -1 0 1970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1009_
timestamp 0
transform -1 0 750 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1010_
timestamp 0
transform -1 0 470 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1011_
timestamp 0
transform 1 0 110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1012_
timestamp 0
transform -1 0 750 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1013_
timestamp 0
transform -1 0 470 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1014_
timestamp 0
transform -1 0 30 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1015_
timestamp 0
transform -1 0 1710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1016_
timestamp 0
transform -1 0 1370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1017_
timestamp 0
transform -1 0 2130 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1018_
timestamp 0
transform -1 0 2210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1019_
timestamp 0
transform -1 0 1470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1020_
timestamp 0
transform -1 0 1390 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1021_
timestamp 0
transform -1 0 1130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1022_
timestamp 0
transform -1 0 990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1023_
timestamp 0
transform 1 0 1410 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1024_
timestamp 0
transform 1 0 1570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1025_
timestamp 0
transform 1 0 1510 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1026_
timestamp 0
transform -1 0 1290 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1027_
timestamp 0
transform 1 0 730 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1028_
timestamp 0
transform -1 0 330 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1029_
timestamp 0
transform 1 0 150 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1030_
timestamp 0
transform -1 0 310 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1031_
timestamp 0
transform -1 0 610 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1032_
timestamp 0
transform -1 0 170 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1033_
timestamp 0
transform 1 0 150 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1034_
timestamp 0
transform -1 0 30 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1035_
timestamp 0
transform -1 0 470 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1036_
timestamp 0
transform -1 0 30 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1037_
timestamp 0
transform -1 0 170 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1038_
timestamp 0
transform -1 0 2970 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1039_
timestamp 0
transform 1 0 830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1040_
timestamp 0
transform -1 0 970 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1041_
timestamp 0
transform 1 0 5290 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1042_
timestamp 0
transform 1 0 4790 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1043_
timestamp 0
transform -1 0 2050 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1044_
timestamp 0
transform -1 0 1030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1045_
timestamp 0
transform -1 0 850 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1046_
timestamp 0
transform -1 0 30 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1047_
timestamp 0
transform 1 0 250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1048_
timestamp 0
transform -1 0 30 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1049_
timestamp 0
transform -1 0 30 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1050_
timestamp 0
transform 1 0 10 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1051_
timestamp 0
transform 1 0 270 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1052_
timestamp 0
transform -1 0 30 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1053_
timestamp 0
transform 1 0 110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1054_
timestamp 0
transform -1 0 470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1055_
timestamp 0
transform 1 0 110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1056_
timestamp 0
transform -1 0 310 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1057_
timestamp 0
transform 1 0 1110 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1058_
timestamp 0
transform -1 0 2250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1059_
timestamp 0
transform -1 0 2530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1060_
timestamp 0
transform -1 0 2030 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1061_
timestamp 0
transform 1 0 2210 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1062_
timestamp 0
transform 1 0 1930 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1063_
timestamp 0
transform -1 0 1450 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1064_
timestamp 0
transform -1 0 1610 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1065_
timestamp 0
transform -1 0 2150 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1066_
timestamp 0
transform 1 0 2650 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1067_
timestamp 0
transform -1 0 2390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1068_
timestamp 0
transform -1 0 1750 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1069_
timestamp 0
transform 1 0 1430 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1070_
timestamp 0
transform 1 0 970 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1071_
timestamp 0
transform -1 0 1310 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1072_
timestamp 0
transform -1 0 1570 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1073_
timestamp 0
transform 1 0 1010 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1074_
timestamp 0
transform -1 0 2290 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1075_
timestamp 0
transform -1 0 2030 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1076_
timestamp 0
transform 1 0 3730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1077_
timestamp 0
transform 1 0 3850 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1078_
timestamp 0
transform 1 0 2210 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1079_
timestamp 0
transform -1 0 2370 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1080_
timestamp 0
transform -1 0 1670 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1081_
timestamp 0
transform 1 0 1750 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1082_
timestamp 0
transform -1 0 1490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1083_
timestamp 0
transform -1 0 1490 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1084_
timestamp 0
transform -1 0 1890 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1085_
timestamp 0
transform -1 0 1850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1086_
timestamp 0
transform -1 0 1030 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1087_
timestamp 0
transform -1 0 890 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1088_
timestamp 0
transform -1 0 1310 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1089_
timestamp 0
transform -1 0 1610 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1090_
timestamp 0
transform -1 0 2290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1091_
timestamp 0
transform 1 0 1510 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1092_
timestamp 0
transform -1 0 1370 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1093_
timestamp 0
transform -1 0 870 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1094_
timestamp 0
transform -1 0 450 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1095_
timestamp 0
transform 1 0 590 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1096_
timestamp 0
transform -1 0 870 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1097_
timestamp 0
transform -1 0 1010 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1098_
timestamp 0
transform 1 0 710 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1099_
timestamp 0
transform -1 0 1930 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1100_
timestamp 0
transform -1 0 1010 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1101_
timestamp 0
transform 1 0 1210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1102_
timestamp 0
transform -1 0 870 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1103_
timestamp 0
transform -1 0 1150 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1104_
timestamp 0
transform -1 0 1810 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1105_
timestamp 0
transform -1 0 1290 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1106_
timestamp 0
transform 1 0 1230 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1107_
timestamp 0
transform 1 0 1090 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1108_
timestamp 0
transform -1 0 1110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1109_
timestamp 0
transform -1 0 990 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1110_
timestamp 0
transform -1 0 970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1111_
timestamp 0
transform 1 0 870 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1112_
timestamp 0
transform 1 0 670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1113_
timestamp 0
transform -1 0 590 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1114_
timestamp 0
transform -1 0 310 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1115_
timestamp 0
transform -1 0 730 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1116_
timestamp 0
transform -1 0 310 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1117_
timestamp 0
transform -1 0 190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1118_
timestamp 0
transform 1 0 390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1119_
timestamp 0
transform -1 0 550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1120_
timestamp 0
transform -1 0 590 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1121_
timestamp 0
transform -1 0 30 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1122_
timestamp 0
transform -1 0 170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1123_
timestamp 0
transform 1 0 150 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1124_
timestamp 0
transform 1 0 310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1125_
timestamp 0
transform 1 0 390 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1126_
timestamp 0
transform 1 0 350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1127_
timestamp 0
transform -1 0 230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1128_
timestamp 0
transform 1 0 1310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1129_
timestamp 0
transform -1 0 1370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1130_
timestamp 0
transform -1 0 1230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1131_
timestamp 0
transform -1 0 1130 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1132_
timestamp 0
transform -1 0 1210 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1133_
timestamp 0
transform -1 0 1050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1134_
timestamp 0
transform -1 0 1310 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1135_
timestamp 0
transform 1 0 990 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1136_
timestamp 0
transform 1 0 1170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1137_
timestamp 0
transform -1 0 870 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1138_
timestamp 0
transform 1 0 430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1139_
timestamp 0
transform 1 0 290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1140_
timestamp 0
transform 1 0 450 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1141_
timestamp 0
transform 1 0 590 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1142_
timestamp 0
transform 1 0 890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1143_
timestamp 0
transform -1 0 1090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1144_
timestamp 0
transform 1 0 2730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1145_
timestamp 0
transform -1 0 3270 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1146_
timestamp 0
transform 1 0 2870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1147_
timestamp 0
transform -1 0 3030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1148_
timestamp 0
transform -1 0 3130 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1149_
timestamp 0
transform -1 0 3070 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1150_
timestamp 0
transform 1 0 2610 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1151_
timestamp 0
transform -1 0 2770 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1152_
timestamp 0
transform -1 0 2870 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1153_
timestamp 0
transform 1 0 1290 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1154_
timestamp 0
transform -1 0 1150 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1155_
timestamp 0
transform -1 0 1430 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1156_
timestamp 0
transform -1 0 1010 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1157_
timestamp 0
transform -1 0 770 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1158_
timestamp 0
transform -1 0 610 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1159_
timestamp 0
transform -1 0 410 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1160_
timestamp 0
transform 1 0 290 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1161_
timestamp 0
transform -1 0 310 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1162_
timestamp 0
transform -1 0 30 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1163_
timestamp 0
transform -1 0 330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1164_
timestamp 0
transform -1 0 30 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1165_
timestamp 0
transform -1 0 30 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1166_
timestamp 0
transform -1 0 150 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1167_
timestamp 0
transform -1 0 30 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1168_
timestamp 0
transform 1 0 910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1169_
timestamp 0
transform 1 0 890 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1170_
timestamp 0
transform 1 0 1010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1171_
timestamp 0
transform 1 0 2990 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1172_
timestamp 0
transform 1 0 3290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1173_
timestamp 0
transform 1 0 3570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1174_
timestamp 0
transform -1 0 3190 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1175_
timestamp 0
transform 1 0 3510 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1176_
timestamp 0
transform 1 0 4350 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1177_
timestamp 0
transform -1 0 4010 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1178_
timestamp 0
transform -1 0 3310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1179_
timestamp 0
transform -1 0 2930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1180_
timestamp 0
transform -1 0 670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1181_
timestamp 0
transform 1 0 770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1182_
timestamp 0
transform -1 0 1090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1183_
timestamp 0
transform 1 0 530 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1184_
timestamp 0
transform -1 0 290 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1185_
timestamp 0
transform 1 0 150 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1186_
timestamp 0
transform -1 0 470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1187_
timestamp 0
transform -1 0 170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1188_
timestamp 0
transform -1 0 150 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1189_
timestamp 0
transform -1 0 270 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1190_
timestamp 0
transform -1 0 130 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1191_
timestamp 0
transform 1 0 130 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1192_
timestamp 0
transform 1 0 310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1193_
timestamp 0
transform 1 0 1210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1194_
timestamp 0
transform -1 0 830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1195_
timestamp 0
transform -1 0 450 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1196_
timestamp 0
transform 1 0 5070 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1197_
timestamp 0
transform 1 0 4570 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1198_
timestamp 0
transform 1 0 3770 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1199_
timestamp 0
transform 1 0 1550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1200_
timestamp 0
transform -1 0 1870 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1201_
timestamp 0
transform 1 0 1590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1202_
timestamp 0
transform -1 0 1470 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1203_
timestamp 0
transform -1 0 1810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1204_
timestamp 0
transform -1 0 1430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1205_
timestamp 0
transform 1 0 1590 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1206_
timestamp 0
transform -1 0 1730 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1207_
timestamp 0
transform -1 0 1170 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1208_
timestamp 0
transform -1 0 1170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1209_
timestamp 0
transform 1 0 1150 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1210_
timestamp 0
transform 1 0 2910 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1211_
timestamp 0
transform 1 0 4130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1212_
timestamp 0
transform 1 0 4010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1213_
timestamp 0
transform -1 0 3870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1214_
timestamp 0
transform -1 0 3590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1215_
timestamp 0
transform 1 0 3310 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1216_
timestamp 0
transform -1 0 3730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1217_
timestamp 0
transform 1 0 3830 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1218_
timestamp 0
transform -1 0 3710 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1219_
timestamp 0
transform -1 0 3430 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1220_
timestamp 0
transform 1 0 3010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1221_
timestamp 0
transform 1 0 1870 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1222_
timestamp 0
transform 1 0 2770 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1223_
timestamp 0
transform -1 0 2990 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1224_
timestamp 0
transform 1 0 2890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1225_
timestamp 0
transform -1 0 2690 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1226_
timestamp 0
transform 1 0 2390 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1227_
timestamp 0
transform 1 0 2350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1228_
timestamp 0
transform 1 0 2070 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1229_
timestamp 0
transform 1 0 2630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1230_
timestamp 0
transform -1 0 2090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1231_
timestamp 0
transform -1 0 3170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1232_
timestamp 0
transform -1 0 2290 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1233_
timestamp 0
transform -1 0 2490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1234_
timestamp 0
transform -1 0 2550 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1235_
timestamp 0
transform -1 0 1930 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1236_
timestamp 0
transform 1 0 1130 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1237_
timestamp 0
transform -1 0 2610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1238_
timestamp 0
transform -1 0 2230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1239_
timestamp 0
transform -1 0 1490 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1240_
timestamp 0
transform -1 0 1210 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1241_
timestamp 0
transform 1 0 1270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1242_
timestamp 0
transform -1 0 1790 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1243_
timestamp 0
transform 1 0 1690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1244_
timestamp 0
transform -1 0 1570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1245_
timestamp 0
transform -1 0 450 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1246_
timestamp 0
transform 1 0 810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1247_
timestamp 0
transform -1 0 1430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1248_
timestamp 0
transform -1 0 1350 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1249_
timestamp 0
transform -1 0 1150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1250_
timestamp 0
transform 1 0 150 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1251_
timestamp 0
transform 1 0 710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1252_
timestamp 0
transform -1 0 990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1253_
timestamp 0
transform -1 0 1290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1254_
timestamp 0
transform -1 0 710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1255_
timestamp 0
transform -1 0 570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1256_
timestamp 0
transform -1 0 550 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1257_
timestamp 0
transform 1 0 830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1258_
timestamp 0
transform -1 0 30 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1259_
timestamp 0
transform -1 0 690 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1260_
timestamp 0
transform 1 0 630 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1261_
timestamp 0
transform 1 0 770 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1262_
timestamp 0
transform 1 0 490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1263_
timestamp 0
transform -1 0 290 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1264_
timestamp 0
transform 1 0 330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1265_
timestamp 0
transform 1 0 170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1266_
timestamp 0
transform -1 0 470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1267_
timestamp 0
transform 1 0 370 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1268_
timestamp 0
transform -1 0 530 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1269_
timestamp 0
transform -1 0 1030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1270_
timestamp 0
transform 1 0 1030 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1271_
timestamp 0
transform -1 0 3170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1272_
timestamp 0
transform 1 0 2650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1273_
timestamp 0
transform 1 0 1090 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1274_
timestamp 0
transform -1 0 2830 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1275_
timestamp 0
transform -1 0 2790 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1276_
timestamp 0
transform -1 0 2790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1277_
timestamp 0
transform 1 0 2390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1278_
timestamp 0
transform 1 0 2230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1279_
timestamp 0
transform -1 0 3390 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1280_
timestamp 0
transform -1 0 3250 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1281_
timestamp 0
transform 1 0 3170 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1282_
timestamp 0
transform -1 0 3230 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1283_
timestamp 0
transform 1 0 3110 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1284_
timestamp 0
transform 1 0 590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1285_
timestamp 0
transform -1 0 590 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1286_
timestamp 0
transform 1 0 710 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1287_
timestamp 0
transform 1 0 1310 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1288_
timestamp 0
transform -1 0 1330 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1289_
timestamp 0
transform -1 0 1990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1290_
timestamp 0
transform 1 0 1830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1291_
timestamp 0
transform 1 0 3710 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1292_
timestamp 0
transform 1 0 3490 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1293_
timestamp 0
transform 1 0 2650 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1294_
timestamp 0
transform -1 0 3450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1295_
timestamp 0
transform 1 0 3130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1296_
timestamp 0
transform 1 0 4110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1297_
timestamp 0
transform 1 0 3550 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1298_
timestamp 0
transform -1 0 3970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1299_
timestamp 0
transform -1 0 3290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1300_
timestamp 0
transform -1 0 3030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1301_
timestamp 0
transform 1 0 3830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1302_
timestamp 0
transform -1 0 3710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1303_
timestamp 0
transform -1 0 3570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1304_
timestamp 0
transform 1 0 2610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1305_
timestamp 0
transform -1 0 4350 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1306_
timestamp 0
transform 1 0 4090 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1307_
timestamp 0
transform -1 0 3750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1308_
timestamp 0
transform 1 0 3570 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1309_
timestamp 0
transform 1 0 3470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1310_
timestamp 0
transform -1 0 3710 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1311_
timestamp 0
transform -1 0 3450 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1312_
timestamp 0
transform -1 0 3410 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1313_
timestamp 0
transform 1 0 3710 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1314_
timestamp 0
transform -1 0 4210 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1315_
timestamp 0
transform 1 0 3950 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1316_
timestamp 0
transform -1 0 3690 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1317_
timestamp 0
transform 1 0 2690 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1318_
timestamp 0
transform 1 0 2950 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1319_
timestamp 0
transform 1 0 3810 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1320_
timestamp 0
transform -1 0 3550 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1321_
timestamp 0
transform -1 0 2850 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1322_
timestamp 0
transform -1 0 3270 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1323_
timestamp 0
transform 1 0 2370 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1324_
timestamp 0
transform -1 0 2310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1325_
timestamp 0
transform -1 0 2770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1326_
timestamp 0
transform 1 0 4830 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1327_
timestamp 0
transform -1 0 2750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1328_
timestamp 0
transform -1 0 2650 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1329_
timestamp 0
transform -1 0 2510 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1330_
timestamp 0
transform -1 0 2350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1331_
timestamp 0
transform 1 0 2170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1332_
timestamp 0
transform -1 0 2490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1333_
timestamp 0
transform -1 0 2150 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1334_
timestamp 0
transform -1 0 2250 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1335_
timestamp 0
transform -1 0 2170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1336_
timestamp 0
transform -1 0 2470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1337_
timestamp 0
transform -1 0 1850 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1338_
timestamp 0
transform -1 0 1770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1339_
timestamp 0
transform -1 0 1430 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1340_
timestamp 0
transform -1 0 1650 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1341_
timestamp 0
transform 1 0 1650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1342_
timestamp 0
transform -1 0 1710 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1343_
timestamp 0
transform 1 0 2110 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1344_
timestamp 0
transform -1 0 2010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1345_
timestamp 0
transform -1 0 1990 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1346_
timestamp 0
transform -1 0 1730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1347_
timestamp 0
transform 1 0 1170 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1348_
timestamp 0
transform -1 0 1570 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1349_
timestamp 0
transform 1 0 1850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1350_
timestamp 0
transform -1 0 1570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1351_
timestamp 0
transform 1 0 1270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1352_
timestamp 0
transform -1 0 470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1353_
timestamp 0
transform -1 0 310 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1354_
timestamp 0
transform -1 0 1430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1355_
timestamp 0
transform -1 0 1050 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1356_
timestamp 0
transform -1 0 910 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1357_
timestamp 0
transform -1 0 770 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1358_
timestamp 0
transform 1 0 890 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1359_
timestamp 0
transform 1 0 730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1360_
timestamp 0
transform 1 0 610 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1361_
timestamp 0
transform 1 0 870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1362_
timestamp 0
transform 1 0 1990 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1363_
timestamp 0
transform -1 0 690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1364_
timestamp 0
transform -1 0 830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1365_
timestamp 0
transform -1 0 650 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1366_
timestamp 0
transform -1 0 510 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1367_
timestamp 0
transform -1 0 3430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1368_
timestamp 0
transform -1 0 1510 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1369_
timestamp 0
transform 1 0 1890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1370_
timestamp 0
transform -1 0 2690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1371_
timestamp 0
transform 1 0 2810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1372_
timestamp 0
transform -1 0 3330 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1373_
timestamp 0
transform 1 0 4630 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1374_
timestamp 0
transform -1 0 3630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1375_
timestamp 0
transform 1 0 3590 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1376_
timestamp 0
transform -1 0 3210 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1377_
timestamp 0
transform -1 0 3210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1378_
timestamp 0
transform -1 0 3350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1379_
timestamp 0
transform -1 0 3070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1380_
timestamp 0
transform 1 0 2910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1381_
timestamp 0
transform 1 0 3070 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1382_
timestamp 0
transform -1 0 2950 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1383_
timestamp 0
transform -1 0 2790 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1384_
timestamp 0
transform 1 0 2130 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1385_
timestamp 0
transform 1 0 3970 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1386_
timestamp 0
transform 1 0 4410 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1387_
timestamp 0
transform 1 0 4110 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1388_
timestamp 0
transform 1 0 4490 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1389_
timestamp 0
transform 1 0 4390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1390_
timestamp 0
transform 1 0 5050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1391_
timestamp 0
transform -1 0 4690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1392_
timestamp 0
transform -1 0 4530 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1393_
timestamp 0
transform 1 0 4550 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1394_
timestamp 0
transform -1 0 4270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1395_
timestamp 0
transform -1 0 4130 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1396_
timestamp 0
transform -1 0 3850 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1397_
timestamp 0
transform -1 0 2410 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1398_
timestamp 0
transform -1 0 2270 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1399_
timestamp 0
transform 1 0 1870 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1400_
timestamp 0
transform -1 0 1990 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1401_
timestamp 0
transform -1 0 2270 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1402_
timestamp 0
transform -1 0 2150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1403_
timestamp 0
transform -1 0 1750 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1404_
timestamp 0
transform -1 0 1750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1405_
timestamp 0
transform -1 0 2050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1406_
timestamp 0
transform -1 0 1990 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1407_
timestamp 0
transform -1 0 2590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1408_
timestamp 0
transform -1 0 2450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1409_
timestamp 0
transform -1 0 2190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1410_
timestamp 0
transform -1 0 2310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1411_
timestamp 0
transform -1 0 2050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1412_
timestamp 0
transform -1 0 1610 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1413_
timestamp 0
transform -1 0 1470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1414_
timestamp 0
transform -1 0 1450 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1415_
timestamp 0
transform -1 0 1650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1416_
timestamp 0
transform -1 0 1490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1417_
timestamp 0
transform -1 0 1370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1418_
timestamp 0
transform -1 0 1350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1419_
timestamp 0
transform -1 0 1630 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1420_
timestamp 0
transform 1 0 1470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1421_
timestamp 0
transform 1 0 1530 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1422_
timestamp 0
transform 1 0 1310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1423_
timestamp 0
transform 1 0 1610 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1424_
timestamp 0
transform 1 0 1830 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1425_
timestamp 0
transform 1 0 1950 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1426_
timestamp 0
transform 1 0 2090 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1427_
timestamp 0
transform 1 0 3430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1428_
timestamp 0
transform 1 0 3350 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1429_
timestamp 0
transform 1 0 3470 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1430_
timestamp 0
transform 1 0 3050 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1431_
timestamp 0
transform -1 0 2970 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1432_
timestamp 0
transform -1 0 2930 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1433_
timestamp 0
transform -1 0 2970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1434_
timestamp 0
transform 1 0 2810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1435_
timestamp 0
transform -1 0 1750 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1436_
timestamp 0
transform 1 0 1770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1437_
timestamp 0
transform -1 0 2650 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1438_
timestamp 0
transform -1 0 2550 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1439_
timestamp 0
transform 1 0 2250 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1440_
timestamp 0
transform -1 0 3730 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1441_
timestamp 0
transform 1 0 4570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1442_
timestamp 0
transform 1 0 4250 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1443_
timestamp 0
transform 1 0 3970 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1444_
timestamp 0
transform 1 0 4650 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1445_
timestamp 0
transform 1 0 4670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1446_
timestamp 0
transform -1 0 4290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1447_
timestamp 0
transform 1 0 3790 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1448_
timestamp 0
transform 1 0 4410 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1449_
timestamp 0
transform -1 0 4230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1450_
timestamp 0
transform -1 0 4130 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1451_
timestamp 0
transform 1 0 4370 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1452_
timestamp 0
transform -1 0 4350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1453_
timestamp 0
transform 1 0 4470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1454_
timestamp 0
transform 1 0 3890 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1455_
timestamp 0
transform -1 0 3590 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1456_
timestamp 0
transform 1 0 4030 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1457_
timestamp 0
transform -1 0 3450 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1458_
timestamp 0
transform -1 0 2710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1459_
timestamp 0
transform 1 0 2790 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1460_
timestamp 0
transform 1 0 2390 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1461_
timestamp 0
transform -1 0 2550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1462_
timestamp 0
transform 1 0 2110 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1463_
timestamp 0
transform -1 0 2670 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1464_
timestamp 0
transform -1 0 2410 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1465_
timestamp 0
transform -1 0 2530 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1466_
timestamp 0
transform 1 0 2010 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1467_
timestamp 0
transform 1 0 1910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1468_
timestamp 0
transform -1 0 1590 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1469_
timestamp 0
transform 1 0 1590 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1470_
timestamp 0
transform -1 0 1890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1471_
timestamp 0
transform -1 0 1830 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1472_
timestamp 0
transform 1 0 1770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1473_
timestamp 0
transform -1 0 1470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1474_
timestamp 0
transform -1 0 1150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1475_
timestamp 0
transform 1 0 1070 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1476_
timestamp 0
transform 1 0 1330 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1477_
timestamp 0
transform -1 0 1690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1478_
timestamp 0
transform 1 0 1470 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1479_
timestamp 0
transform -1 0 1730 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1480_
timestamp 0
transform 1 0 1210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1481_
timestamp 0
transform 1 0 2810 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1482_
timestamp 0
transform -1 0 2790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1483_
timestamp 0
transform 1 0 2350 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1484_
timestamp 0
transform -1 0 3110 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1485_
timestamp 0
transform 1 0 2670 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1486_
timestamp 0
transform 1 0 2810 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1487_
timestamp 0
transform 1 0 2650 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1488_
timestamp 0
transform 1 0 2830 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1489_
timestamp 0
transform 1 0 2970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1490_
timestamp 0
transform -1 0 4170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1491_
timestamp 0
transform -1 0 4030 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1492_
timestamp 0
transform -1 0 2930 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1493_
timestamp 0
transform 1 0 4450 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1494_
timestamp 0
transform -1 0 3990 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1495_
timestamp 0
transform -1 0 4250 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1496_
timestamp 0
transform -1 0 4530 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1497_
timestamp 0
transform 1 0 4570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1498_
timestamp 0
transform 1 0 4430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1499_
timestamp 0
transform -1 0 4730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1500_
timestamp 0
transform 1 0 4650 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1501_
timestamp 0
transform 1 0 4710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1502_
timestamp 0
transform 1 0 4810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1503_
timestamp 0
transform 1 0 4970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1504_
timestamp 0
transform 1 0 4830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1505_
timestamp 0
transform -1 0 4610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1506_
timestamp 0
transform -1 0 3330 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1507_
timestamp 0
transform -1 0 3170 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1508_
timestamp 0
transform -1 0 3030 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1509_
timestamp 0
transform 1 0 3470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1510_
timestamp 0
transform 1 0 3890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1511_
timestamp 0
transform -1 0 3630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1512_
timestamp 0
transform 1 0 3350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1513_
timestamp 0
transform 1 0 3070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1514_
timestamp 0
transform 1 0 3190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1515_
timestamp 0
transform -1 0 3150 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1516_
timestamp 0
transform -1 0 2690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1517_
timestamp 0
transform -1 0 1310 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1518_
timestamp 0
transform 1 0 1930 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1519_
timestamp 0
transform -1 0 1690 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1520_
timestamp 0
transform -1 0 910 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1521_
timestamp 0
transform 1 0 750 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1522_
timestamp 0
transform -1 0 2410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1523_
timestamp 0
transform 1 0 930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1524_
timestamp 0
transform -1 0 1570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1525_
timestamp 0
transform 1 0 1150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1526_
timestamp 0
transform 1 0 1190 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1527_
timestamp 0
transform 1 0 2750 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1528_
timestamp 0
transform 1 0 2910 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1529_
timestamp 0
transform 1 0 290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1530_
timestamp 0
transform 1 0 390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1531_
timestamp 0
transform 1 0 530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1532_
timestamp 0
transform 1 0 2770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1533_
timestamp 0
transform -1 0 2530 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1534_
timestamp 0
transform -1 0 2530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1535_
timestamp 0
transform -1 0 2670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1536_
timestamp 0
transform -1 0 2930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1537_
timestamp 0
transform -1 0 30 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1538_
timestamp 0
transform -1 0 30 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1539_
timestamp 0
transform 1 0 150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1540_
timestamp 0
transform 1 0 3190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1541_
timestamp 0
transform -1 0 3350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1542_
timestamp 0
transform 1 0 3010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1543_
timestamp 0
transform -1 0 3770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1544_
timestamp 0
transform 1 0 4930 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1545_
timestamp 0
transform 1 0 4810 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1546_
timestamp 0
transform 1 0 5030 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1547_
timestamp 0
transform 1 0 4170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1548_
timestamp 0
transform -1 0 4310 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1549_
timestamp 0
transform 1 0 4290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1550_
timestamp 0
transform 1 0 5450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1551_
timestamp 0
transform 1 0 4930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1552_
timestamp 0
transform 1 0 5490 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1553_
timestamp 0
transform 1 0 5350 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1554_
timestamp 0
transform 1 0 5610 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1555_
timestamp 0
transform -1 0 5630 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1556_
timestamp 0
transform 1 0 5230 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1557_
timestamp 0
transform 1 0 3830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1558_
timestamp 0
transform -1 0 3710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1559_
timestamp 0
transform 1 0 3550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1560_
timestamp 0
transform -1 0 2910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1561_
timestamp 0
transform 1 0 3170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1562_
timestamp 0
transform 1 0 3170 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1563_
timestamp 0
transform -1 0 3430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1564_
timestamp 0
transform 1 0 3310 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1565_
timestamp 0
transform 1 0 3350 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1566_
timestamp 0
transform 1 0 3150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1567_
timestamp 0
transform 1 0 350 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1568_
timestamp 0
transform 1 0 470 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1569_
timestamp 0
transform 1 0 590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1570_
timestamp 0
transform 1 0 3070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1571_
timestamp 0
transform 1 0 1930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1572_
timestamp 0
transform 1 0 3070 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1573_
timestamp 0
transform -1 0 3050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1574_
timestamp 0
transform 1 0 3030 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1575_
timestamp 0
transform 1 0 3270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1576_
timestamp 0
transform 1 0 5190 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1577_
timestamp 0
transform -1 0 4050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1578_
timestamp 0
transform -1 0 3630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1579_
timestamp 0
transform 1 0 3750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1580_
timestamp 0
transform 1 0 3490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1581_
timestamp 0
transform -1 0 3270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1582_
timestamp 0
transform -1 0 3370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1583_
timestamp 0
transform -1 0 2790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1584_
timestamp 0
transform 1 0 2530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1585_
timestamp 0
transform 1 0 3450 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1586_
timestamp 0
transform -1 0 3130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1587_
timestamp 0
transform 1 0 3630 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1588_
timestamp 0
transform 1 0 3630 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1589_
timestamp 0
transform -1 0 3910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1590_
timestamp 0
transform 1 0 3850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1591_
timestamp 0
transform 1 0 590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1592_
timestamp 0
transform 1 0 850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1593_
timestamp 0
transform 1 0 710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1594_
timestamp 0
transform 1 0 3470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1595_
timestamp 0
transform 1 0 3690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1596_
timestamp 0
transform 1 0 5610 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1597_
timestamp 0
transform -1 0 5710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1598_
timestamp 0
transform -1 0 5590 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1599_
timestamp 0
transform 1 0 5570 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1600_
timestamp 0
transform -1 0 5570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1601_
timestamp 0
transform 1 0 5490 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1602_
timestamp 0
transform 1 0 5590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1603_
timestamp 0
transform 1 0 4890 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1604_
timestamp 0
transform 1 0 5090 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1605_
timestamp 0
transform 1 0 4930 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1606_
timestamp 0
transform -1 0 5110 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1607_
timestamp 0
transform -1 0 4850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1608_
timestamp 0
transform -1 0 4970 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1609_
timestamp 0
transform 1 0 5310 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1610_
timestamp 0
transform -1 0 5490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1611_
timestamp 0
transform 1 0 5410 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1612_
timestamp 0
transform -1 0 5550 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1613_
timestamp 0
transform -1 0 5550 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1614_
timestamp 0
transform -1 0 5610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1615_
timestamp 0
transform 1 0 5330 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1616_
timestamp 0
transform 1 0 5550 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1617_
timestamp 0
transform 1 0 5430 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1618_
timestamp 0
transform 1 0 5530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1619_
timestamp 0
transform 1 0 5150 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1620_
timestamp 0
transform -1 0 5210 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1621_
timestamp 0
transform 1 0 4690 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1622_
timestamp 0
transform -1 0 4850 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1623_
timestamp 0
transform 1 0 4170 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1624_
timestamp 0
transform -1 0 4830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1625_
timestamp 0
transform 1 0 4510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1626_
timestamp 0
transform 1 0 4470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1627_
timestamp 0
transform 1 0 4210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1628_
timestamp 0
transform 1 0 5110 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1629_
timestamp 0
transform 1 0 4970 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1630_
timestamp 0
transform 1 0 5130 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1631_
timestamp 0
transform -1 0 4390 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1632_
timestamp 0
transform 1 0 5670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1633_
timestamp 0
transform 1 0 5390 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1634_
timestamp 0
transform -1 0 5450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1635_
timestamp 0
transform 1 0 5050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1636_
timestamp 0
transform -1 0 5670 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1637_
timestamp 0
transform 1 0 5650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1638_
timestamp 0
transform 1 0 5090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1639_
timestamp 0
transform -1 0 4970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1640_
timestamp 0
transform 1 0 4930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1641_
timestamp 0
transform 1 0 4670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1642_
timestamp 0
transform -1 0 4370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1643_
timestamp 0
transform 1 0 4310 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1644_
timestamp 0
transform -1 0 4950 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1645_
timestamp 0
transform 1 0 4690 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1646_
timestamp 0
transform -1 0 4790 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1647_
timestamp 0
transform -1 0 5030 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1648_
timestamp 0
transform -1 0 4890 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1649_
timestamp 0
transform 1 0 5650 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1650_
timestamp 0
transform 1 0 5390 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1651_
timestamp 0
transform 1 0 5670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1652_
timestamp 0
transform 1 0 5310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1685_
timestamp 0
transform 1 0 5050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1686_
timestamp 0
transform 1 0 5210 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1687_
timestamp 0
transform 1 0 5430 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1688_
timestamp 0
transform 1 0 5430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1689_
timestamp 0
transform -1 0 5310 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1690_
timestamp 0
transform 1 0 5670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1691_
timestamp 0
transform 1 0 5330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1692_
timestamp 0
transform 1 0 5270 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1693_
timestamp 0
transform -1 0 4850 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1694_
timestamp 0
transform 1 0 5370 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1695_
timestamp 0
transform -1 0 4970 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1696_
timestamp 0
transform -1 0 5690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1697_
timestamp 0
transform 1 0 5490 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1698_
timestamp 0
transform 1 0 5450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1699_
timestamp 0
transform -1 0 5490 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1700_
timestamp 0
transform 1 0 5410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1701_
timestamp 0
transform 1 0 5630 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1702_
timestamp 0
transform 1 0 5570 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1703_
timestamp 0
transform -1 0 4890 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1704_
timestamp 0
transform 1 0 5010 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1705_
timestamp 0
transform 1 0 4930 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1706_
timestamp 0
transform 1 0 5330 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1707_
timestamp 0
transform -1 0 5490 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1708_
timestamp 0
transform -1 0 5170 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1709_
timestamp 0
transform -1 0 5290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1710_
timestamp 0
transform -1 0 5170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1711_
timestamp 0
transform 1 0 4950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1712_
timestamp 0
transform 1 0 5610 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1713_
timestamp 0
transform -1 0 5210 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1714_
timestamp 0
transform -1 0 5190 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1715_
timestamp 0
transform 1 0 5090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1716_
timestamp 0
transform 1 0 5250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1717_
timestamp 0
transform -1 0 5130 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1718_
timestamp 0
transform -1 0 5230 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1719_
timestamp 0
transform 1 0 5330 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1720_
timestamp 0
transform -1 0 5310 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1721_
timestamp 0
transform 1 0 5530 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1722_
timestamp 0
transform -1 0 5390 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1723_
timestamp 0
transform 1 0 5430 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1724_
timestamp 0
transform 1 0 5250 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1725_
timestamp 0
transform 1 0 5270 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1726_
timestamp 0
transform -1 0 5170 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1727_
timestamp 0
transform 1 0 5390 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1728_
timestamp 0
transform 1 0 5570 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1729_
timestamp 0
transform 1 0 5590 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1730_
timestamp 0
transform 1 0 5650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1731_
timestamp 0
transform 1 0 5670 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1732_
timestamp 0
transform 1 0 5530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1733_
timestamp 0
transform -1 0 5570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1734_
timestamp 0
transform -1 0 5430 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1735_
timestamp 0
transform 1 0 5210 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1736_
timestamp 0
transform -1 0 4910 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1737_
timestamp 0
transform 1 0 4770 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1738_
timestamp 0
transform 1 0 4350 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1739_
timestamp 0
transform -1 0 3370 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1740_
timestamp 0
transform 1 0 5030 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1741_
timestamp 0
transform -1 0 4630 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1742_
timestamp 0
transform 1 0 4690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1743_
timestamp 0
transform 1 0 5110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1744_
timestamp 0
transform 1 0 5210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1745_
timestamp 0
transform 1 0 5150 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1746_
timestamp 0
transform 1 0 4990 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1747_
timestamp 0
transform -1 0 4990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1748_
timestamp 0
transform -1 0 4830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1749_
timestamp 0
transform -1 0 4490 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1750_
timestamp 0
transform 1 0 4610 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1751_
timestamp 0
transform 1 0 4950 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1752_
timestamp 0
transform -1 0 5090 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1753_
timestamp 0
transform 1 0 4910 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1754_
timestamp 0
transform -1 0 3950 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1755_
timestamp 0
transform 1 0 4790 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1756_
timestamp 0
transform -1 0 4790 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1757_
timestamp 0
transform -1 0 4490 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1758_
timestamp 0
transform -1 0 3590 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1759_
timestamp 0
transform -1 0 3250 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1760_
timestamp 0
transform -1 0 4690 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1761_
timestamp 0
transform 1 0 4050 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1762_
timestamp 0
transform 1 0 4570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1763_
timestamp 0
transform 1 0 4350 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1764_
timestamp 0
transform 1 0 4650 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1765_
timestamp 0
transform 1 0 4490 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1766_
timestamp 0
transform -1 0 4310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1767_
timestamp 0
transform 1 0 4430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1768_
timestamp 0
transform -1 0 4410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1769_
timestamp 0
transform -1 0 4270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1770_
timestamp 0
transform -1 0 4230 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1771_
timestamp 0
transform -1 0 4090 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1772_
timestamp 0
transform -1 0 4330 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1773_
timestamp 0
transform -1 0 4550 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1774_
timestamp 0
transform -1 0 4030 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1775_
timestamp 0
transform 1 0 3890 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1776_
timestamp 0
transform -1 0 3870 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1777_
timestamp 0
transform -1 0 3090 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1778_
timestamp 0
transform 1 0 3610 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1779_
timestamp 0
transform -1 0 3770 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1780_
timestamp 0
transform -1 0 4430 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1781_
timestamp 0
transform 1 0 4350 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1782_
timestamp 0
transform -1 0 4390 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1783_
timestamp 0
transform -1 0 4050 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1784_
timestamp 0
transform -1 0 3950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1785_
timestamp 0
transform 1 0 4070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1786_
timestamp 0
transform -1 0 4210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1787_
timestamp 0
transform -1 0 3750 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1788_
timestamp 0
transform 1 0 3890 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1789_
timestamp 0
transform -1 0 4390 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1790_
timestamp 0
transform -1 0 4250 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1791_
timestamp 0
transform -1 0 4110 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1792_
timestamp 0
transform -1 0 3970 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1793_
timestamp 0
transform 1 0 3970 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1794_
timestamp 0
transform -1 0 4230 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1795_
timestamp 0
transform -1 0 4190 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1796_
timestamp 0
transform 1 0 3950 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1797_
timestamp 0
transform -1 0 3830 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1798_
timestamp 0
transform -1 0 3730 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1799_
timestamp 0
transform -1 0 3470 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1800_
timestamp 0
transform -1 0 3330 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1801_
timestamp 0
transform 1 0 4150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1802_
timestamp 0
transform 1 0 4670 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1803_
timestamp 0
transform -1 0 4590 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1804_
timestamp 0
transform -1 0 4330 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1805_
timestamp 0
transform -1 0 4370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1806_
timestamp 0
transform 1 0 4430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1807_
timestamp 0
transform 1 0 4510 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1808_
timestamp 0
transform 1 0 4690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1809_
timestamp 0
transform -1 0 4570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1810_
timestamp 0
transform -1 0 4670 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1811_
timestamp 0
transform -1 0 4530 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1812_
timestamp 0
transform -1 0 4290 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1813_
timestamp 0
transform 1 0 4110 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1814_
timestamp 0
transform -1 0 3590 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1815_
timestamp 0
transform 1 0 3570 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1816_
timestamp 0
transform 1 0 3310 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1817_
timestamp 0
transform 1 0 3330 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1818_
timestamp 0
transform -1 0 3450 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1819_
timestamp 0
transform -1 0 3350 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1820_
timestamp 0
transform -1 0 4030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1821_
timestamp 0
transform -1 0 4190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1822_
timestamp 0
transform -1 0 4170 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1823_
timestamp 0
transform -1 0 3610 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1824_
timestamp 0
transform 1 0 3430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1825_
timestamp 0
transform 1 0 3710 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1826_
timestamp 0
transform -1 0 3570 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1827_
timestamp 0
transform -1 0 3670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1828_
timestamp 0
transform -1 0 3530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1829_
timestamp 0
transform -1 0 2750 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1830_
timestamp 0
transform -1 0 2550 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1831_
timestamp 0
transform -1 0 3190 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1832_
timestamp 0
transform -1 0 2930 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1833_
timestamp 0
transform 1 0 2950 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1834_
timestamp 0
transform -1 0 2370 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1835_
timestamp 0
transform -1 0 3070 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1836_
timestamp 0
transform 1 0 5050 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1837_
timestamp 0
transform -1 0 4970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1838_
timestamp 0
transform 1 0 4690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1839_
timestamp 0
transform 1 0 4510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1840_
timestamp 0
transform 1 0 4810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1841_
timestamp 0
transform 1 0 4790 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1842_
timestamp 0
transform 1 0 3670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1843_
timestamp 0
transform -1 0 3550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1844_
timestamp 0
transform 1 0 3830 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1845_
timestamp 0
transform -1 0 3710 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1846_
timestamp 0
transform 1 0 1950 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1847_
timestamp 0
transform -1 0 2090 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1848_
timestamp 0
transform -1 0 2470 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1849_
timestamp 0
transform 1 0 2410 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1850_
timestamp 0
transform 1 0 4030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1851_
timestamp 0
transform 1 0 3910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1852_
timestamp 0
transform -1 0 3290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1853_
timestamp 0
transform -1 0 2670 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1854_
timestamp 0
transform 1 0 2770 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1855_
timestamp 0
transform 1 0 2890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1856_
timestamp 0
transform 1 0 3010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1857_
timestamp 0
transform -1 0 2310 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1858_
timestamp 0
transform -1 0 2850 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1859_
timestamp 0
transform 1 0 3450 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1860_
timestamp 0
transform -1 0 3250 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1861_
timestamp 0
transform -1 0 2850 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1862_
timestamp 0
transform -1 0 2990 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1863_
timestamp 0
transform -1 0 4730 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1864_
timestamp 0
transform -1 0 3110 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1865_
timestamp 0
transform 1 0 2950 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1866_
timestamp 0
transform 1 0 3190 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1867_
timestamp 0
transform -1 0 3490 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1868_
timestamp 0
transform 1 0 3330 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1869_
timestamp 0
transform -1 0 2710 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1870_
timestamp 0
transform 1 0 2590 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1871_
timestamp 0
transform 1 0 3030 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1872_
timestamp 0
transform 1 0 2830 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1873_
timestamp 0
transform -1 0 2570 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1874_
timestamp 0
transform -1 0 2230 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1875_
timestamp 0
transform 1 0 1830 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1876_
timestamp 0
transform -1 0 1710 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1877_
timestamp 0
transform -1 0 3430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1878_
timestamp 0
transform 1 0 3790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1879_
timestamp 0
transform -1 0 3190 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1880_
timestamp 0
transform 1 0 2710 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1881_
timestamp 0
transform -1 0 2590 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1882_
timestamp 0
transform -1 0 2470 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1883_
timestamp 0
transform -1 0 1530 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1884_
timestamp 0
transform -1 0 1630 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1885_
timestamp 0
transform -1 0 2030 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1886_
timestamp 0
transform 1 0 1870 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1887_
timestamp 0
transform -1 0 1770 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1888_
timestamp 0
transform 1 0 2410 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1889_
timestamp 0
transform 1 0 2270 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1890_
timestamp 0
transform -1 0 1370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1891_
timestamp 0
transform -1 0 30 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1892_
timestamp 0
transform -1 0 30 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1893_
timestamp 0
transform 1 0 2170 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1894_
timestamp 0
transform -1 0 3450 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1895_
timestamp 0
transform -1 0 3710 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1896_
timestamp 0
transform -1 0 3830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1897_
timestamp 0
transform 1 0 3810 0 -1 250
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert5
timestamp 0
transform 1 0 3750 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert6
timestamp 0
transform -1 0 2230 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert7
timestamp 0
transform -1 0 3970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert8
timestamp 0
transform -1 0 2890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert9
timestamp 0
transform -1 0 2550 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert10
timestamp 0
transform -1 0 2590 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert11
timestamp 0
transform 1 0 4830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert12
timestamp 0
transform -1 0 4790 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert13
timestamp 0
transform -1 0 4770 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert14
timestamp 0
transform 1 0 5050 0 -1 730
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert0
timestamp 0
transform -1 0 5190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert1
timestamp 0
transform 1 0 5410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert2
timestamp 0
transform -1 0 5190 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert3
timestamp 0
transform -1 0 4550 0 1 5530
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert4
timestamp 0
transform -1 0 5310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__920_
timestamp 0
transform -1 0 3650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__921_
timestamp 0
transform 1 0 4090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__922_
timestamp 0
transform -1 0 3890 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__923_
timestamp 0
transform -1 0 3910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__924_
timestamp 0
transform 1 0 4270 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__925_
timestamp 0
transform -1 0 3630 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__926_
timestamp 0
transform 1 0 2350 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__927_
timestamp 0
transform -1 0 1170 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__928_
timestamp 0
transform 1 0 2230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__929_
timestamp 0
transform 1 0 2090 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__930_
timestamp 0
transform -1 0 2250 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__931_
timestamp 0
transform -1 0 1010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__932_
timestamp 0
transform -1 0 1750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__933_
timestamp 0
transform 1 0 3910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__934_
timestamp 0
transform -1 0 2530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__935_
timestamp 0
transform -1 0 2390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__936_
timestamp 0
transform 1 0 1450 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__937_
timestamp 0
transform -1 0 1190 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__938_
timestamp 0
transform -1 0 2110 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__939_
timestamp 0
transform 1 0 1110 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__940_
timestamp 0
transform -1 0 2530 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__941_
timestamp 0
transform -1 0 1830 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__942_
timestamp 0
transform -1 0 1570 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__943_
timestamp 0
transform -1 0 1090 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__944_
timestamp 0
transform 1 0 2430 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__945_
timestamp 0
transform 1 0 2510 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__946_
timestamp 0
transform -1 0 2370 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__947_
timestamp 0
transform -1 0 990 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__948_
timestamp 0
transform -1 0 1290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__949_
timestamp 0
transform -1 0 870 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__950_
timestamp 0
transform 1 0 830 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__951_
timestamp 0
transform -1 0 3990 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__952_
timestamp 0
transform 1 0 2470 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__953_
timestamp 0
transform -1 0 1370 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__954_
timestamp 0
transform -1 0 770 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__955_
timestamp 0
transform -1 0 710 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__956_
timestamp 0
transform 1 0 770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__957_
timestamp 0
transform -1 0 730 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__958_
timestamp 0
transform 1 0 1950 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__959_
timestamp 0
transform -1 0 2090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__960_
timestamp 0
transform -1 0 650 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__961_
timestamp 0
transform -1 0 5110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__962_
timestamp 0
transform 1 0 2630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__963_
timestamp 0
transform -1 0 1950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__964_
timestamp 0
transform -1 0 1690 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__965_
timestamp 0
transform -1 0 50 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__966_
timestamp 0
transform -1 0 350 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__967_
timestamp 0
transform -1 0 570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__968_
timestamp 0
transform -1 0 310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__969_
timestamp 0
transform -1 0 210 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__970_
timestamp 0
transform -1 0 190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__971_
timestamp 0
transform -1 0 1010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__972_
timestamp 0
transform -1 0 50 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__973_
timestamp 0
transform -1 0 510 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__974_
timestamp 0
transform -1 0 190 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__975_
timestamp 0
transform 1 0 4150 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__976_
timestamp 0
transform -1 0 3930 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__977_
timestamp 0
transform -1 0 1630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__978_
timestamp 0
transform 1 0 870 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__979_
timestamp 0
transform -1 0 2150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__980_
timestamp 0
transform -1 0 2010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__981_
timestamp 0
transform -1 0 1890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__982_
timestamp 0
transform 1 0 1470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__983_
timestamp 0
transform 1 0 750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__984_
timestamp 0
transform -1 0 630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__985_
timestamp 0
transform 1 0 970 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__986_
timestamp 0
transform -1 0 730 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__987_
timestamp 0
transform -1 0 610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__988_
timestamp 0
transform -1 0 190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__989_
timestamp 0
transform 1 0 310 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__990_
timestamp 0
transform 1 0 310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__991_
timestamp 0
transform -1 0 590 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__992_
timestamp 0
transform -1 0 470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__993_
timestamp 0
transform 1 0 450 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__994_
timestamp 0
transform -1 0 50 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__995_
timestamp 0
transform -1 0 50 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__996_
timestamp 0
transform 1 0 170 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__997_
timestamp 0
transform -1 0 50 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__998_
timestamp 0
transform -1 0 50 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__999_
timestamp 0
transform 1 0 390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1000_
timestamp 0
transform -1 0 1830 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1001_
timestamp 0
transform -1 0 2130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1002_
timestamp 0
transform 1 0 1270 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1003_
timestamp 0
transform 1 0 1390 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1004_
timestamp 0
transform -1 0 1670 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1005_
timestamp 0
transform 1 0 890 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1006_
timestamp 0
transform 1 0 610 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1007_
timestamp 0
transform -1 0 1190 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1008_
timestamp 0
transform -1 0 1990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1009_
timestamp 0
transform -1 0 770 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1010_
timestamp 0
transform -1 0 490 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1011_
timestamp 0
transform 1 0 130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1012_
timestamp 0
transform -1 0 770 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1013_
timestamp 0
transform -1 0 490 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1014_
timestamp 0
transform -1 0 50 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1015_
timestamp 0
transform -1 0 1730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1016_
timestamp 0
transform -1 0 1390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1017_
timestamp 0
transform -1 0 2150 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1018_
timestamp 0
transform -1 0 2230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1019_
timestamp 0
transform -1 0 1490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1020_
timestamp 0
transform -1 0 1410 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1021_
timestamp 0
transform -1 0 1150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1022_
timestamp 0
transform -1 0 1010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1023_
timestamp 0
transform 1 0 1430 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1024_
timestamp 0
transform 1 0 1590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1025_
timestamp 0
transform 1 0 1530 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1026_
timestamp 0
transform -1 0 1310 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1027_
timestamp 0
transform 1 0 750 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1028_
timestamp 0
transform -1 0 350 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1029_
timestamp 0
transform 1 0 170 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1030_
timestamp 0
transform -1 0 330 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1031_
timestamp 0
transform -1 0 630 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1032_
timestamp 0
transform -1 0 190 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1033_
timestamp 0
transform 1 0 170 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1034_
timestamp 0
transform -1 0 50 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1035_
timestamp 0
transform -1 0 490 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1036_
timestamp 0
transform -1 0 50 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1037_
timestamp 0
transform -1 0 190 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1038_
timestamp 0
transform -1 0 2990 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1039_
timestamp 0
transform 1 0 850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1040_
timestamp 0
transform -1 0 990 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1041_
timestamp 0
transform 1 0 5310 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1042_
timestamp 0
transform 1 0 4810 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1043_
timestamp 0
transform -1 0 2070 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1044_
timestamp 0
transform -1 0 1050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1045_
timestamp 0
transform -1 0 870 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1046_
timestamp 0
transform -1 0 50 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1047_
timestamp 0
transform 1 0 270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1048_
timestamp 0
transform -1 0 50 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1049_
timestamp 0
transform -1 0 50 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1050_
timestamp 0
transform 1 0 30 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1051_
timestamp 0
transform 1 0 290 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1052_
timestamp 0
transform -1 0 50 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1053_
timestamp 0
transform 1 0 130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1054_
timestamp 0
transform -1 0 490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1055_
timestamp 0
transform 1 0 130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1056_
timestamp 0
transform -1 0 330 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1057_
timestamp 0
transform 1 0 1130 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1058_
timestamp 0
transform -1 0 2270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1059_
timestamp 0
transform -1 0 2550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1060_
timestamp 0
transform -1 0 2050 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1061_
timestamp 0
transform 1 0 2230 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1062_
timestamp 0
transform 1 0 1950 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1063_
timestamp 0
transform -1 0 1470 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1064_
timestamp 0
transform -1 0 1630 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1065_
timestamp 0
transform -1 0 2170 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1066_
timestamp 0
transform 1 0 2670 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1067_
timestamp 0
transform -1 0 2410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1068_
timestamp 0
transform -1 0 1770 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1069_
timestamp 0
transform 1 0 1450 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1070_
timestamp 0
transform 1 0 990 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1071_
timestamp 0
transform -1 0 1330 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1072_
timestamp 0
transform -1 0 1590 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1073_
timestamp 0
transform 1 0 1030 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1074_
timestamp 0
transform -1 0 2310 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1075_
timestamp 0
transform -1 0 2050 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1076_
timestamp 0
transform 1 0 3750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1077_
timestamp 0
transform 1 0 3870 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1078_
timestamp 0
transform 1 0 2230 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1079_
timestamp 0
transform -1 0 2390 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1080_
timestamp 0
transform -1 0 1690 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1081_
timestamp 0
transform 1 0 1770 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1082_
timestamp 0
transform -1 0 1510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1083_
timestamp 0
transform -1 0 1510 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1084_
timestamp 0
transform -1 0 1910 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1085_
timestamp 0
transform -1 0 1870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1086_
timestamp 0
transform -1 0 1050 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1087_
timestamp 0
transform -1 0 910 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1088_
timestamp 0
transform -1 0 1330 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1089_
timestamp 0
transform -1 0 1630 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1090_
timestamp 0
transform -1 0 2310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1091_
timestamp 0
transform 1 0 1530 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1092_
timestamp 0
transform -1 0 1390 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1093_
timestamp 0
transform -1 0 890 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1094_
timestamp 0
transform -1 0 470 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1095_
timestamp 0
transform 1 0 610 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1096_
timestamp 0
transform -1 0 890 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1097_
timestamp 0
transform -1 0 1030 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1098_
timestamp 0
transform 1 0 730 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1099_
timestamp 0
transform -1 0 1950 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1100_
timestamp 0
transform -1 0 1030 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1101_
timestamp 0
transform 1 0 1230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1102_
timestamp 0
transform -1 0 890 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1103_
timestamp 0
transform -1 0 1170 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1104_
timestamp 0
transform -1 0 1830 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1105_
timestamp 0
transform -1 0 1310 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1106_
timestamp 0
transform 1 0 1250 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1107_
timestamp 0
transform 1 0 1110 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1108_
timestamp 0
transform -1 0 1130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1109_
timestamp 0
transform -1 0 1010 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1110_
timestamp 0
transform -1 0 990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1111_
timestamp 0
transform 1 0 890 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1112_
timestamp 0
transform 1 0 690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1113_
timestamp 0
transform -1 0 610 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1114_
timestamp 0
transform -1 0 330 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1115_
timestamp 0
transform -1 0 750 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1116_
timestamp 0
transform -1 0 330 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1117_
timestamp 0
transform -1 0 210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1118_
timestamp 0
transform 1 0 410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1119_
timestamp 0
transform -1 0 570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1120_
timestamp 0
transform -1 0 610 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1121_
timestamp 0
transform -1 0 50 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1122_
timestamp 0
transform -1 0 190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1123_
timestamp 0
transform 1 0 170 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1124_
timestamp 0
transform 1 0 330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1125_
timestamp 0
transform 1 0 410 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1126_
timestamp 0
transform 1 0 370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1127_
timestamp 0
transform -1 0 250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1128_
timestamp 0
transform 1 0 1330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1129_
timestamp 0
transform -1 0 1390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1130_
timestamp 0
transform -1 0 1250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1131_
timestamp 0
transform -1 0 1150 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1132_
timestamp 0
transform -1 0 1230 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1133_
timestamp 0
transform -1 0 1070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1134_
timestamp 0
transform -1 0 1330 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1135_
timestamp 0
transform 1 0 1010 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1136_
timestamp 0
transform 1 0 1190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1137_
timestamp 0
transform -1 0 890 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1138_
timestamp 0
transform 1 0 450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1139_
timestamp 0
transform 1 0 310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1140_
timestamp 0
transform 1 0 470 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1141_
timestamp 0
transform 1 0 610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1142_
timestamp 0
transform 1 0 910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1143_
timestamp 0
transform -1 0 1110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1144_
timestamp 0
transform 1 0 2750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1145_
timestamp 0
transform -1 0 3290 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1146_
timestamp 0
transform 1 0 2890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1147_
timestamp 0
transform -1 0 3050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1148_
timestamp 0
transform -1 0 3150 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1149_
timestamp 0
transform -1 0 3090 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1150_
timestamp 0
transform 1 0 2630 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1151_
timestamp 0
transform -1 0 2790 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1152_
timestamp 0
transform -1 0 2890 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1153_
timestamp 0
transform 1 0 1310 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1154_
timestamp 0
transform -1 0 1170 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1155_
timestamp 0
transform -1 0 1450 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1156_
timestamp 0
transform -1 0 1030 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1157_
timestamp 0
transform -1 0 790 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1158_
timestamp 0
transform -1 0 630 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1159_
timestamp 0
transform -1 0 430 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1160_
timestamp 0
transform 1 0 310 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1161_
timestamp 0
transform -1 0 330 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1162_
timestamp 0
transform -1 0 50 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1163_
timestamp 0
transform -1 0 350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1164_
timestamp 0
transform -1 0 50 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1165_
timestamp 0
transform -1 0 50 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1166_
timestamp 0
transform -1 0 170 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1167_
timestamp 0
transform -1 0 50 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1168_
timestamp 0
transform 1 0 930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1169_
timestamp 0
transform 1 0 910 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1170_
timestamp 0
transform 1 0 1030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1171_
timestamp 0
transform 1 0 3010 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1172_
timestamp 0
transform 1 0 3310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1173_
timestamp 0
transform 1 0 3590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1174_
timestamp 0
transform -1 0 3210 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1175_
timestamp 0
transform 1 0 3530 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1176_
timestamp 0
transform 1 0 4370 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1177_
timestamp 0
transform -1 0 4030 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1178_
timestamp 0
transform -1 0 3330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1179_
timestamp 0
transform -1 0 2950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1180_
timestamp 0
transform -1 0 690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1181_
timestamp 0
transform 1 0 790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1182_
timestamp 0
transform -1 0 1110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1183_
timestamp 0
transform 1 0 550 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1184_
timestamp 0
transform -1 0 310 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1185_
timestamp 0
transform 1 0 170 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1186_
timestamp 0
transform -1 0 490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1187_
timestamp 0
transform -1 0 190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1188_
timestamp 0
transform -1 0 170 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1189_
timestamp 0
transform -1 0 290 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1190_
timestamp 0
transform -1 0 150 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1191_
timestamp 0
transform 1 0 150 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1192_
timestamp 0
transform 1 0 330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1193_
timestamp 0
transform 1 0 1230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1194_
timestamp 0
transform -1 0 850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1195_
timestamp 0
transform -1 0 470 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1196_
timestamp 0
transform 1 0 5090 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1197_
timestamp 0
transform 1 0 4590 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1198_
timestamp 0
transform 1 0 3790 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1199_
timestamp 0
transform 1 0 1570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1200_
timestamp 0
transform -1 0 1890 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1201_
timestamp 0
transform 1 0 1610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1202_
timestamp 0
transform -1 0 1490 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1203_
timestamp 0
transform -1 0 1830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1204_
timestamp 0
transform -1 0 1450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1205_
timestamp 0
transform 1 0 1610 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1206_
timestamp 0
transform -1 0 1750 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1207_
timestamp 0
transform -1 0 1190 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1208_
timestamp 0
transform -1 0 1190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1209_
timestamp 0
transform 1 0 1170 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1210_
timestamp 0
transform 1 0 2930 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1211_
timestamp 0
transform 1 0 4150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1212_
timestamp 0
transform 1 0 4030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1213_
timestamp 0
transform -1 0 3890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1214_
timestamp 0
transform -1 0 3610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1215_
timestamp 0
transform 1 0 3330 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1216_
timestamp 0
transform -1 0 3750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1217_
timestamp 0
transform 1 0 3850 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1218_
timestamp 0
transform -1 0 3730 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1219_
timestamp 0
transform -1 0 3450 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1220_
timestamp 0
transform 1 0 3030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1221_
timestamp 0
transform 1 0 1890 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1222_
timestamp 0
transform 1 0 2790 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1223_
timestamp 0
transform -1 0 3010 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1224_
timestamp 0
transform 1 0 2910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1225_
timestamp 0
transform -1 0 2710 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1226_
timestamp 0
transform 1 0 2410 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1227_
timestamp 0
transform 1 0 2370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1228_
timestamp 0
transform 1 0 2090 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1229_
timestamp 0
transform 1 0 2650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1230_
timestamp 0
transform -1 0 2110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1231_
timestamp 0
transform -1 0 3190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1232_
timestamp 0
transform -1 0 2310 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1233_
timestamp 0
transform -1 0 2510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1234_
timestamp 0
transform -1 0 2570 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1235_
timestamp 0
transform -1 0 1950 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1236_
timestamp 0
transform 1 0 1150 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1237_
timestamp 0
transform -1 0 2630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1238_
timestamp 0
transform -1 0 2250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1239_
timestamp 0
transform -1 0 1510 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1240_
timestamp 0
transform -1 0 1230 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1241_
timestamp 0
transform 1 0 1290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1242_
timestamp 0
transform -1 0 1810 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1243_
timestamp 0
transform 1 0 1710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1244_
timestamp 0
transform -1 0 1590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1245_
timestamp 0
transform -1 0 470 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1246_
timestamp 0
transform 1 0 830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1247_
timestamp 0
transform -1 0 1450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1248_
timestamp 0
transform -1 0 1370 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1249_
timestamp 0
transform -1 0 1170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1250_
timestamp 0
transform 1 0 170 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1251_
timestamp 0
transform 1 0 730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1252_
timestamp 0
transform -1 0 1010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1253_
timestamp 0
transform -1 0 1310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1254_
timestamp 0
transform -1 0 730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1255_
timestamp 0
transform -1 0 590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1256_
timestamp 0
transform -1 0 570 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1257_
timestamp 0
transform 1 0 850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1258_
timestamp 0
transform -1 0 50 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1259_
timestamp 0
transform -1 0 710 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1260_
timestamp 0
transform 1 0 650 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1261_
timestamp 0
transform 1 0 790 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1262_
timestamp 0
transform 1 0 510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1263_
timestamp 0
transform -1 0 310 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1264_
timestamp 0
transform 1 0 350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1265_
timestamp 0
transform 1 0 190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1266_
timestamp 0
transform -1 0 490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1267_
timestamp 0
transform 1 0 390 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1268_
timestamp 0
transform -1 0 550 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1269_
timestamp 0
transform -1 0 1050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1270_
timestamp 0
transform 1 0 1050 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1271_
timestamp 0
transform -1 0 3190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1272_
timestamp 0
transform 1 0 2670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1273_
timestamp 0
transform 1 0 1110 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1274_
timestamp 0
transform -1 0 2850 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1275_
timestamp 0
transform -1 0 2810 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1276_
timestamp 0
transform -1 0 2810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1277_
timestamp 0
transform 1 0 2410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1278_
timestamp 0
transform 1 0 2250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1279_
timestamp 0
transform -1 0 3410 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1280_
timestamp 0
transform -1 0 3270 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1281_
timestamp 0
transform 1 0 3190 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1282_
timestamp 0
transform -1 0 3250 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1283_
timestamp 0
transform 1 0 3130 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1284_
timestamp 0
transform 1 0 610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1285_
timestamp 0
transform -1 0 610 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1286_
timestamp 0
transform 1 0 730 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1287_
timestamp 0
transform 1 0 1330 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1288_
timestamp 0
transform -1 0 1350 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1289_
timestamp 0
transform -1 0 2010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1290_
timestamp 0
transform 1 0 1850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1291_
timestamp 0
transform 1 0 3730 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1292_
timestamp 0
transform 1 0 3510 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1293_
timestamp 0
transform 1 0 2670 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1294_
timestamp 0
transform -1 0 3470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1295_
timestamp 0
transform 1 0 3150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1296_
timestamp 0
transform 1 0 4130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1297_
timestamp 0
transform 1 0 3570 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1298_
timestamp 0
transform -1 0 3990 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1299_
timestamp 0
transform -1 0 3310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1300_
timestamp 0
transform -1 0 3050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1301_
timestamp 0
transform 1 0 3850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1302_
timestamp 0
transform -1 0 3730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1303_
timestamp 0
transform -1 0 3590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1304_
timestamp 0
transform 1 0 2630 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1305_
timestamp 0
transform -1 0 4370 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1306_
timestamp 0
transform 1 0 4110 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1307_
timestamp 0
transform -1 0 3770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1308_
timestamp 0
transform 1 0 3590 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1309_
timestamp 0
transform 1 0 3490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1310_
timestamp 0
transform -1 0 3730 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1311_
timestamp 0
transform -1 0 3470 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1312_
timestamp 0
transform -1 0 3430 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1313_
timestamp 0
transform 1 0 3730 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1314_
timestamp 0
transform -1 0 4230 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1315_
timestamp 0
transform 1 0 3970 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1316_
timestamp 0
transform -1 0 3710 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1317_
timestamp 0
transform 1 0 2710 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1318_
timestamp 0
transform 1 0 2970 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1319_
timestamp 0
transform 1 0 3830 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1320_
timestamp 0
transform -1 0 3570 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1321_
timestamp 0
transform -1 0 2870 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1322_
timestamp 0
transform -1 0 3290 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1323_
timestamp 0
transform 1 0 2390 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1324_
timestamp 0
transform -1 0 2330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1325_
timestamp 0
transform -1 0 2790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1326_
timestamp 0
transform 1 0 4850 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1327_
timestamp 0
transform -1 0 2770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1328_
timestamp 0
transform -1 0 2670 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1329_
timestamp 0
transform -1 0 2530 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1330_
timestamp 0
transform -1 0 2370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1331_
timestamp 0
transform 1 0 2190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1332_
timestamp 0
transform -1 0 2510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1333_
timestamp 0
transform -1 0 2170 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1334_
timestamp 0
transform -1 0 2270 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1335_
timestamp 0
transform -1 0 2190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1336_
timestamp 0
transform -1 0 2490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1337_
timestamp 0
transform -1 0 1870 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1338_
timestamp 0
transform -1 0 1790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1339_
timestamp 0
transform -1 0 1450 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1340_
timestamp 0
transform -1 0 1670 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1341_
timestamp 0
transform 1 0 1670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1342_
timestamp 0
transform -1 0 1730 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1343_
timestamp 0
transform 1 0 2130 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1344_
timestamp 0
transform -1 0 2030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1345_
timestamp 0
transform -1 0 2010 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1346_
timestamp 0
transform -1 0 1750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1347_
timestamp 0
transform 1 0 1190 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1348_
timestamp 0
transform -1 0 1590 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1349_
timestamp 0
transform 1 0 1870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1350_
timestamp 0
transform -1 0 1590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1351_
timestamp 0
transform 1 0 1290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1352_
timestamp 0
transform -1 0 490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1353_
timestamp 0
transform -1 0 330 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1354_
timestamp 0
transform -1 0 1450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1355_
timestamp 0
transform -1 0 1070 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1356_
timestamp 0
transform -1 0 930 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1357_
timestamp 0
transform -1 0 790 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1358_
timestamp 0
transform 1 0 910 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1359_
timestamp 0
transform 1 0 750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1360_
timestamp 0
transform 1 0 630 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1361_
timestamp 0
transform 1 0 890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1362_
timestamp 0
transform 1 0 2010 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1363_
timestamp 0
transform -1 0 710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1364_
timestamp 0
transform -1 0 850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1365_
timestamp 0
transform -1 0 670 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1366_
timestamp 0
transform -1 0 530 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1367_
timestamp 0
transform -1 0 3450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1368_
timestamp 0
transform -1 0 1530 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1369_
timestamp 0
transform 1 0 1910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1370_
timestamp 0
transform -1 0 2710 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1371_
timestamp 0
transform 1 0 2830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1372_
timestamp 0
transform -1 0 3350 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1373_
timestamp 0
transform 1 0 4650 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1374_
timestamp 0
transform -1 0 3650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1375_
timestamp 0
transform 1 0 3610 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1376_
timestamp 0
transform -1 0 3230 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1377_
timestamp 0
transform -1 0 3230 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1378_
timestamp 0
transform -1 0 3370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1379_
timestamp 0
transform -1 0 3090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1380_
timestamp 0
transform 1 0 2930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1381_
timestamp 0
transform 1 0 3090 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1382_
timestamp 0
transform -1 0 2970 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1383_
timestamp 0
transform -1 0 2810 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1384_
timestamp 0
transform 1 0 2150 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1385_
timestamp 0
transform 1 0 3990 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1386_
timestamp 0
transform 1 0 4430 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1387_
timestamp 0
transform 1 0 4130 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1388_
timestamp 0
transform 1 0 4510 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1389_
timestamp 0
transform 1 0 4410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1390_
timestamp 0
transform 1 0 5070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1391_
timestamp 0
transform -1 0 4710 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1392_
timestamp 0
transform -1 0 4550 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1393_
timestamp 0
transform 1 0 4570 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1394_
timestamp 0
transform -1 0 4290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1395_
timestamp 0
transform -1 0 4150 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1396_
timestamp 0
transform -1 0 3870 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1397_
timestamp 0
transform -1 0 2430 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1398_
timestamp 0
transform -1 0 2290 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1399_
timestamp 0
transform 1 0 1890 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1400_
timestamp 0
transform -1 0 2010 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1401_
timestamp 0
transform -1 0 2290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1402_
timestamp 0
transform -1 0 2170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1403_
timestamp 0
transform -1 0 1770 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1404_
timestamp 0
transform -1 0 1770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1405_
timestamp 0
transform -1 0 2070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1406_
timestamp 0
transform -1 0 2010 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1407_
timestamp 0
transform -1 0 2610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1408_
timestamp 0
transform -1 0 2470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1409_
timestamp 0
transform -1 0 2210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1410_
timestamp 0
transform -1 0 2330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1411_
timestamp 0
transform -1 0 2070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1412_
timestamp 0
transform -1 0 1630 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1413_
timestamp 0
transform -1 0 1490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1414_
timestamp 0
transform -1 0 1470 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1415_
timestamp 0
transform -1 0 1670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1416_
timestamp 0
transform -1 0 1510 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1417_
timestamp 0
transform -1 0 1390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1418_
timestamp 0
transform -1 0 1370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1419_
timestamp 0
transform -1 0 1650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1420_
timestamp 0
transform 1 0 1490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1421_
timestamp 0
transform 1 0 1550 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1422_
timestamp 0
transform 1 0 1330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1423_
timestamp 0
transform 1 0 1630 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1424_
timestamp 0
transform 1 0 1850 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1425_
timestamp 0
transform 1 0 1970 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1426_
timestamp 0
transform 1 0 2110 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1427_
timestamp 0
transform 1 0 3450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1428_
timestamp 0
transform 1 0 3370 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1429_
timestamp 0
transform 1 0 3490 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1430_
timestamp 0
transform 1 0 3070 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1431_
timestamp 0
transform -1 0 2990 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1432_
timestamp 0
transform -1 0 2950 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1433_
timestamp 0
transform -1 0 2990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1434_
timestamp 0
transform 1 0 2830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1435_
timestamp 0
transform -1 0 1770 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1436_
timestamp 0
transform 1 0 1790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1437_
timestamp 0
transform -1 0 2670 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1438_
timestamp 0
transform -1 0 2570 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1439_
timestamp 0
transform 1 0 2270 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1440_
timestamp 0
transform -1 0 3750 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1441_
timestamp 0
transform 1 0 4590 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1442_
timestamp 0
transform 1 0 4270 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1443_
timestamp 0
transform 1 0 3990 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1444_
timestamp 0
transform 1 0 4670 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1445_
timestamp 0
transform 1 0 4690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1446_
timestamp 0
transform -1 0 4310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1447_
timestamp 0
transform 1 0 3810 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1448_
timestamp 0
transform 1 0 4430 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1449_
timestamp 0
transform -1 0 4250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1450_
timestamp 0
transform -1 0 4150 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1451_
timestamp 0
transform 1 0 4390 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1452_
timestamp 0
transform -1 0 4370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1453_
timestamp 0
transform 1 0 4490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1454_
timestamp 0
transform 1 0 3910 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1455_
timestamp 0
transform -1 0 3610 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1456_
timestamp 0
transform 1 0 4050 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1457_
timestamp 0
transform -1 0 3470 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1458_
timestamp 0
transform -1 0 2730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1459_
timestamp 0
transform 1 0 2810 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1460_
timestamp 0
transform 1 0 2410 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1461_
timestamp 0
transform -1 0 2570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1462_
timestamp 0
transform 1 0 2130 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1463_
timestamp 0
transform -1 0 2690 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1464_
timestamp 0
transform -1 0 2430 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1465_
timestamp 0
transform -1 0 2550 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1466_
timestamp 0
transform 1 0 2030 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1467_
timestamp 0
transform 1 0 1930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1468_
timestamp 0
transform -1 0 1610 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1469_
timestamp 0
transform 1 0 1610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1470_
timestamp 0
transform -1 0 1910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1471_
timestamp 0
transform -1 0 1850 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1472_
timestamp 0
transform 1 0 1790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1473_
timestamp 0
transform -1 0 1490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1474_
timestamp 0
transform -1 0 1170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1475_
timestamp 0
transform 1 0 1090 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1476_
timestamp 0
transform 1 0 1350 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1477_
timestamp 0
transform -1 0 1710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1478_
timestamp 0
transform 1 0 1490 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1479_
timestamp 0
transform -1 0 1750 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1480_
timestamp 0
transform 1 0 1230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1481_
timestamp 0
transform 1 0 2830 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1482_
timestamp 0
transform -1 0 2810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1483_
timestamp 0
transform 1 0 2370 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1484_
timestamp 0
transform -1 0 3130 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1485_
timestamp 0
transform 1 0 2690 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1486_
timestamp 0
transform 1 0 2830 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1487_
timestamp 0
transform 1 0 2670 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1488_
timestamp 0
transform 1 0 2850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1489_
timestamp 0
transform 1 0 2990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1490_
timestamp 0
transform -1 0 4190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1491_
timestamp 0
transform -1 0 4050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1492_
timestamp 0
transform -1 0 2950 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1493_
timestamp 0
transform 1 0 4470 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1494_
timestamp 0
transform -1 0 4010 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1495_
timestamp 0
transform -1 0 4270 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1496_
timestamp 0
transform -1 0 4550 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1497_
timestamp 0
transform 1 0 4590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1498_
timestamp 0
transform 1 0 4450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1499_
timestamp 0
transform -1 0 4750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1500_
timestamp 0
transform 1 0 4670 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1501_
timestamp 0
transform 1 0 4730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1502_
timestamp 0
transform 1 0 4830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1503_
timestamp 0
transform 1 0 4990 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1504_
timestamp 0
transform 1 0 4850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1505_
timestamp 0
transform -1 0 4630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1506_
timestamp 0
transform -1 0 3350 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1507_
timestamp 0
transform -1 0 3190 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1508_
timestamp 0
transform -1 0 3050 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1509_
timestamp 0
transform 1 0 3490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1510_
timestamp 0
transform 1 0 3910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1511_
timestamp 0
transform -1 0 3650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1512_
timestamp 0
transform 1 0 3370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1513_
timestamp 0
transform 1 0 3090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1514_
timestamp 0
transform 1 0 3210 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1515_
timestamp 0
transform -1 0 3170 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1516_
timestamp 0
transform -1 0 2710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1517_
timestamp 0
transform -1 0 1330 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1518_
timestamp 0
transform 1 0 1950 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1519_
timestamp 0
transform -1 0 1710 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1520_
timestamp 0
transform -1 0 930 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1521_
timestamp 0
transform 1 0 770 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1522_
timestamp 0
transform -1 0 2430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1523_
timestamp 0
transform 1 0 950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1524_
timestamp 0
transform -1 0 1590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1525_
timestamp 0
transform 1 0 1170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1526_
timestamp 0
transform 1 0 1210 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1527_
timestamp 0
transform 1 0 2770 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1528_
timestamp 0
transform 1 0 2930 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1529_
timestamp 0
transform 1 0 310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1530_
timestamp 0
transform 1 0 410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1531_
timestamp 0
transform 1 0 550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1532_
timestamp 0
transform 1 0 2790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1533_
timestamp 0
transform -1 0 2550 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1534_
timestamp 0
transform -1 0 2550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1535_
timestamp 0
transform -1 0 2690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1536_
timestamp 0
transform -1 0 2950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1537_
timestamp 0
transform -1 0 50 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1538_
timestamp 0
transform -1 0 50 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1539_
timestamp 0
transform 1 0 170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1540_
timestamp 0
transform 1 0 3210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1541_
timestamp 0
transform -1 0 3370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1542_
timestamp 0
transform 1 0 3030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1543_
timestamp 0
transform -1 0 3790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1544_
timestamp 0
transform 1 0 4950 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1545_
timestamp 0
transform 1 0 4830 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1546_
timestamp 0
transform 1 0 5050 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1547_
timestamp 0
transform 1 0 4190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1548_
timestamp 0
transform -1 0 4330 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1549_
timestamp 0
transform 1 0 4310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1550_
timestamp 0
transform 1 0 5470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1551_
timestamp 0
transform 1 0 4950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1552_
timestamp 0
transform 1 0 5510 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1553_
timestamp 0
transform 1 0 5370 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1554_
timestamp 0
transform 1 0 5630 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1555_
timestamp 0
transform -1 0 5650 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1556_
timestamp 0
transform 1 0 5250 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1557_
timestamp 0
transform 1 0 3850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1558_
timestamp 0
transform -1 0 3730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1559_
timestamp 0
transform 1 0 3570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1560_
timestamp 0
transform -1 0 2930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1561_
timestamp 0
transform 1 0 3190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1562_
timestamp 0
transform 1 0 3190 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1563_
timestamp 0
transform -1 0 3450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1564_
timestamp 0
transform 1 0 3330 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1565_
timestamp 0
transform 1 0 3370 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1566_
timestamp 0
transform 1 0 3170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1567_
timestamp 0
transform 1 0 370 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1568_
timestamp 0
transform 1 0 490 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1569_
timestamp 0
transform 1 0 610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1570_
timestamp 0
transform 1 0 3090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1571_
timestamp 0
transform 1 0 1950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1572_
timestamp 0
transform 1 0 3090 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1573_
timestamp 0
transform -1 0 3070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1574_
timestamp 0
transform 1 0 3050 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1575_
timestamp 0
transform 1 0 3290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1576_
timestamp 0
transform 1 0 5210 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1577_
timestamp 0
transform -1 0 4070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1578_
timestamp 0
transform -1 0 3650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1579_
timestamp 0
transform 1 0 3770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1580_
timestamp 0
transform 1 0 3510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1581_
timestamp 0
transform -1 0 3290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1582_
timestamp 0
transform -1 0 3390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1583_
timestamp 0
transform -1 0 2810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1584_
timestamp 0
transform 1 0 2550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1585_
timestamp 0
transform 1 0 3470 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1586_
timestamp 0
transform -1 0 3150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1587_
timestamp 0
transform 1 0 3650 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1588_
timestamp 0
transform 1 0 3650 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1589_
timestamp 0
transform -1 0 3930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1590_
timestamp 0
transform 1 0 3870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1591_
timestamp 0
transform 1 0 610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1592_
timestamp 0
transform 1 0 870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1593_
timestamp 0
transform 1 0 730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1594_
timestamp 0
transform 1 0 3490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1595_
timestamp 0
transform 1 0 3710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1596_
timestamp 0
transform 1 0 5630 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1597_
timestamp 0
transform -1 0 5730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1598_
timestamp 0
transform -1 0 5610 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1599_
timestamp 0
transform 1 0 5590 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1600_
timestamp 0
transform -1 0 5590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1601_
timestamp 0
transform 1 0 5510 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1602_
timestamp 0
transform 1 0 5610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1603_
timestamp 0
transform 1 0 4910 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1604_
timestamp 0
transform 1 0 5110 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1605_
timestamp 0
transform 1 0 4950 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1606_
timestamp 0
transform -1 0 5130 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1607_
timestamp 0
transform -1 0 4870 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1608_
timestamp 0
transform -1 0 4990 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1609_
timestamp 0
transform 1 0 5330 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1610_
timestamp 0
transform -1 0 5510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1611_
timestamp 0
transform 1 0 5430 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1612_
timestamp 0
transform -1 0 5570 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1613_
timestamp 0
transform -1 0 5570 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1614_
timestamp 0
transform -1 0 5630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1615_
timestamp 0
transform 1 0 5350 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1616_
timestamp 0
transform 1 0 5570 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1617_
timestamp 0
transform 1 0 5450 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1618_
timestamp 0
transform 1 0 5550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1619_
timestamp 0
transform 1 0 5170 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1620_
timestamp 0
transform -1 0 5230 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1621_
timestamp 0
transform 1 0 4710 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1622_
timestamp 0
transform -1 0 4870 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1623_
timestamp 0
transform 1 0 4190 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1624_
timestamp 0
transform -1 0 4850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1625_
timestamp 0
transform 1 0 4530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1626_
timestamp 0
transform 1 0 4490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1627_
timestamp 0
transform 1 0 4230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1628_
timestamp 0
transform 1 0 5130 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1629_
timestamp 0
transform 1 0 4990 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1630_
timestamp 0
transform 1 0 5150 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1631_
timestamp 0
transform -1 0 4410 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1632_
timestamp 0
transform 1 0 5690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1633_
timestamp 0
transform 1 0 5410 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1634_
timestamp 0
transform -1 0 5470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1635_
timestamp 0
transform 1 0 5070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1636_
timestamp 0
transform -1 0 5690 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1637_
timestamp 0
transform 1 0 5670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1638_
timestamp 0
transform 1 0 5110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1639_
timestamp 0
transform -1 0 4990 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1640_
timestamp 0
transform 1 0 4950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1641_
timestamp 0
transform 1 0 4690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1642_
timestamp 0
transform -1 0 4390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1643_
timestamp 0
transform 1 0 4330 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1644_
timestamp 0
transform -1 0 4970 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1645_
timestamp 0
transform 1 0 4710 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1646_
timestamp 0
transform -1 0 4810 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1647_
timestamp 0
transform -1 0 5050 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1648_
timestamp 0
transform -1 0 4910 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1649_
timestamp 0
transform 1 0 5670 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1650_
timestamp 0
transform 1 0 5410 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1651_
timestamp 0
transform 1 0 5690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1652_
timestamp 0
transform 1 0 5330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1685_
timestamp 0
transform 1 0 5070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1686_
timestamp 0
transform 1 0 5230 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1687_
timestamp 0
transform 1 0 5450 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1688_
timestamp 0
transform 1 0 5450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1689_
timestamp 0
transform -1 0 5330 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1690_
timestamp 0
transform 1 0 5690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1691_
timestamp 0
transform 1 0 5350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1692_
timestamp 0
transform 1 0 5290 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1693_
timestamp 0
transform -1 0 4870 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1694_
timestamp 0
transform 1 0 5390 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1695_
timestamp 0
transform -1 0 4990 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1696_
timestamp 0
transform -1 0 5710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1697_
timestamp 0
transform 1 0 5510 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1698_
timestamp 0
transform 1 0 5470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1699_
timestamp 0
transform -1 0 5510 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1700_
timestamp 0
transform 1 0 5430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1701_
timestamp 0
transform 1 0 5650 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1702_
timestamp 0
transform 1 0 5590 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1703_
timestamp 0
transform -1 0 4910 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1704_
timestamp 0
transform 1 0 5030 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1705_
timestamp 0
transform 1 0 4950 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1706_
timestamp 0
transform 1 0 5350 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1707_
timestamp 0
transform -1 0 5510 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1708_
timestamp 0
transform -1 0 5190 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1709_
timestamp 0
transform -1 0 5310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1710_
timestamp 0
transform -1 0 5190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1711_
timestamp 0
transform 1 0 4970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1712_
timestamp 0
transform 1 0 5630 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1713_
timestamp 0
transform -1 0 5230 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1714_
timestamp 0
transform -1 0 5210 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1715_
timestamp 0
transform 1 0 5110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1716_
timestamp 0
transform 1 0 5270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1717_
timestamp 0
transform -1 0 5150 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1718_
timestamp 0
transform -1 0 5250 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1719_
timestamp 0
transform 1 0 5350 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1720_
timestamp 0
transform -1 0 5330 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1721_
timestamp 0
transform 1 0 5550 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1722_
timestamp 0
transform -1 0 5410 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1723_
timestamp 0
transform 1 0 5450 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1724_
timestamp 0
transform 1 0 5270 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1725_
timestamp 0
transform 1 0 5290 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1726_
timestamp 0
transform -1 0 5190 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1727_
timestamp 0
transform 1 0 5410 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1728_
timestamp 0
transform 1 0 5590 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1729_
timestamp 0
transform 1 0 5610 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1730_
timestamp 0
transform 1 0 5670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1731_
timestamp 0
transform 1 0 5690 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1732_
timestamp 0
transform 1 0 5550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1733_
timestamp 0
transform -1 0 5590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1734_
timestamp 0
transform -1 0 5450 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1735_
timestamp 0
transform 1 0 5230 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1736_
timestamp 0
transform -1 0 4930 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1737_
timestamp 0
transform 1 0 4790 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1738_
timestamp 0
transform 1 0 4370 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1739_
timestamp 0
transform -1 0 3390 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1740_
timestamp 0
transform 1 0 5050 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1741_
timestamp 0
transform -1 0 4650 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1742_
timestamp 0
transform 1 0 4710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1743_
timestamp 0
transform 1 0 5130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1744_
timestamp 0
transform 1 0 5230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1745_
timestamp 0
transform 1 0 5170 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1746_
timestamp 0
transform 1 0 5010 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1747_
timestamp 0
transform -1 0 5010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1748_
timestamp 0
transform -1 0 4850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1749_
timestamp 0
transform -1 0 4510 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1750_
timestamp 0
transform 1 0 4630 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1751_
timestamp 0
transform 1 0 4970 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1752_
timestamp 0
transform -1 0 5110 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1753_
timestamp 0
transform 1 0 4930 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1754_
timestamp 0
transform -1 0 3970 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1755_
timestamp 0
transform 1 0 4810 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1756_
timestamp 0
transform -1 0 4810 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1757_
timestamp 0
transform -1 0 4510 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1758_
timestamp 0
transform -1 0 3610 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1759_
timestamp 0
transform -1 0 3270 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1760_
timestamp 0
transform -1 0 4710 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1761_
timestamp 0
transform 1 0 4070 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1762_
timestamp 0
transform 1 0 4590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1763_
timestamp 0
transform 1 0 4370 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1764_
timestamp 0
transform 1 0 4670 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1765_
timestamp 0
transform 1 0 4510 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1766_
timestamp 0
transform -1 0 4330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1767_
timestamp 0
transform 1 0 4450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1768_
timestamp 0
transform -1 0 4430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1769_
timestamp 0
transform -1 0 4290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1770_
timestamp 0
transform -1 0 4250 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1771_
timestamp 0
transform -1 0 4110 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1772_
timestamp 0
transform -1 0 4350 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1773_
timestamp 0
transform -1 0 4570 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1774_
timestamp 0
transform -1 0 4050 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1775_
timestamp 0
transform 1 0 3910 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1776_
timestamp 0
transform -1 0 3890 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1777_
timestamp 0
transform -1 0 3110 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1778_
timestamp 0
transform 1 0 3630 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1779_
timestamp 0
transform -1 0 3790 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1780_
timestamp 0
transform -1 0 4450 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1781_
timestamp 0
transform 1 0 4370 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1782_
timestamp 0
transform -1 0 4410 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1783_
timestamp 0
transform -1 0 4070 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1784_
timestamp 0
transform -1 0 3970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1785_
timestamp 0
transform 1 0 4090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1786_
timestamp 0
transform -1 0 4230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1787_
timestamp 0
transform -1 0 3770 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1788_
timestamp 0
transform 1 0 3910 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1789_
timestamp 0
transform -1 0 4410 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1790_
timestamp 0
transform -1 0 4270 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1791_
timestamp 0
transform -1 0 4130 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1792_
timestamp 0
transform -1 0 3990 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1793_
timestamp 0
transform 1 0 3990 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1794_
timestamp 0
transform -1 0 4250 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1795_
timestamp 0
transform -1 0 4210 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1796_
timestamp 0
transform 1 0 3970 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1797_
timestamp 0
transform -1 0 3850 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1798_
timestamp 0
transform -1 0 3750 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1799_
timestamp 0
transform -1 0 3490 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1800_
timestamp 0
transform -1 0 3350 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1801_
timestamp 0
transform 1 0 4170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1802_
timestamp 0
transform 1 0 4690 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1803_
timestamp 0
transform -1 0 4610 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1804_
timestamp 0
transform -1 0 4350 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1805_
timestamp 0
transform -1 0 4390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1806_
timestamp 0
transform 1 0 4450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1807_
timestamp 0
transform 1 0 4530 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1808_
timestamp 0
transform 1 0 4710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1809_
timestamp 0
transform -1 0 4590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1810_
timestamp 0
transform -1 0 4690 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1811_
timestamp 0
transform -1 0 4550 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1812_
timestamp 0
transform -1 0 4310 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1813_
timestamp 0
transform 1 0 4130 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1814_
timestamp 0
transform -1 0 3610 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1815_
timestamp 0
transform 1 0 3590 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1816_
timestamp 0
transform 1 0 3330 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1817_
timestamp 0
transform 1 0 3350 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1818_
timestamp 0
transform -1 0 3470 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1819_
timestamp 0
transform -1 0 3370 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1820_
timestamp 0
transform -1 0 4050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1821_
timestamp 0
transform -1 0 4210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1822_
timestamp 0
transform -1 0 4190 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1823_
timestamp 0
transform -1 0 3630 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1824_
timestamp 0
transform 1 0 3450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1825_
timestamp 0
transform 1 0 3730 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1826_
timestamp 0
transform -1 0 3590 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1827_
timestamp 0
transform -1 0 3690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1828_
timestamp 0
transform -1 0 3550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1829_
timestamp 0
transform -1 0 2770 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1830_
timestamp 0
transform -1 0 2570 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1831_
timestamp 0
transform -1 0 3210 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1832_
timestamp 0
transform -1 0 2950 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1833_
timestamp 0
transform 1 0 2970 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1834_
timestamp 0
transform -1 0 2390 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1835_
timestamp 0
transform -1 0 3090 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1836_
timestamp 0
transform 1 0 5070 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1837_
timestamp 0
transform -1 0 4990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1838_
timestamp 0
transform 1 0 4710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1839_
timestamp 0
transform 1 0 4530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1840_
timestamp 0
transform 1 0 4830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1841_
timestamp 0
transform 1 0 4810 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1842_
timestamp 0
transform 1 0 3690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1843_
timestamp 0
transform -1 0 3570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1844_
timestamp 0
transform 1 0 3850 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1845_
timestamp 0
transform -1 0 3730 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1846_
timestamp 0
transform 1 0 1970 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1847_
timestamp 0
transform -1 0 2110 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1848_
timestamp 0
transform -1 0 2490 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1849_
timestamp 0
transform 1 0 2430 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1850_
timestamp 0
transform 1 0 4050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1851_
timestamp 0
transform 1 0 3930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1852_
timestamp 0
transform -1 0 3310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1853_
timestamp 0
transform -1 0 2690 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1854_
timestamp 0
transform 1 0 2790 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1855_
timestamp 0
transform 1 0 2910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1856_
timestamp 0
transform 1 0 3030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1857_
timestamp 0
transform -1 0 2330 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1858_
timestamp 0
transform -1 0 2870 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1859_
timestamp 0
transform 1 0 3470 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1860_
timestamp 0
transform -1 0 3270 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1861_
timestamp 0
transform -1 0 2870 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1862_
timestamp 0
transform -1 0 3010 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1863_
timestamp 0
transform -1 0 4750 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1864_
timestamp 0
transform -1 0 3130 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1865_
timestamp 0
transform 1 0 2970 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1866_
timestamp 0
transform 1 0 3210 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1867_
timestamp 0
transform -1 0 3510 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1868_
timestamp 0
transform 1 0 3350 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1869_
timestamp 0
transform -1 0 2730 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1870_
timestamp 0
transform 1 0 2610 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1871_
timestamp 0
transform 1 0 3050 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1872_
timestamp 0
transform 1 0 2850 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1873_
timestamp 0
transform -1 0 2590 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1874_
timestamp 0
transform -1 0 2250 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1875_
timestamp 0
transform 1 0 1850 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1876_
timestamp 0
transform -1 0 1730 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1877_
timestamp 0
transform -1 0 3450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1878_
timestamp 0
transform 1 0 3810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1879_
timestamp 0
transform -1 0 3210 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1880_
timestamp 0
transform 1 0 2730 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1881_
timestamp 0
transform -1 0 2610 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1882_
timestamp 0
transform -1 0 2490 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1883_
timestamp 0
transform -1 0 1550 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1884_
timestamp 0
transform -1 0 1650 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1885_
timestamp 0
transform -1 0 2050 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1886_
timestamp 0
transform 1 0 1890 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1887_
timestamp 0
transform -1 0 1790 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1888_
timestamp 0
transform 1 0 2430 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1889_
timestamp 0
transform 1 0 2290 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1890_
timestamp 0
transform -1 0 1390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1891_
timestamp 0
transform -1 0 50 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1892_
timestamp 0
transform -1 0 50 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1893_
timestamp 0
transform 1 0 2190 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1894_
timestamp 0
transform -1 0 3470 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1895_
timestamp 0
transform -1 0 3730 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1896_
timestamp 0
transform -1 0 3850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1897_
timestamp 0
transform 1 0 3830 0 -1 250
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert5
timestamp 0
transform 1 0 3770 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert6
timestamp 0
transform -1 0 2250 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert7
timestamp 0
transform -1 0 3990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert8
timestamp 0
transform -1 0 2910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert9
timestamp 0
transform -1 0 2570 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert10
timestamp 0
transform -1 0 2610 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert11
timestamp 0
transform 1 0 4850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert12
timestamp 0
transform -1 0 4810 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert13
timestamp 0
transform -1 0 4790 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert14
timestamp 0
transform 1 0 5070 0 -1 730
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert0
timestamp 0
transform -1 0 5210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert1
timestamp 0
transform 1 0 5430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert2
timestamp 0
transform -1 0 5210 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert3
timestamp 0
transform -1 0 4570 0 1 5530
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert4
timestamp 0
transform -1 0 5330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__920_
timestamp 0
transform -1 0 3670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__927_
timestamp 0
transform -1 0 1190 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__933_
timestamp 0
transform 1 0 3930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__940_
timestamp 0
transform -1 0 2550 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__946_
timestamp 0
transform -1 0 2390 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__953_
timestamp 0
transform -1 0 1390 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__959_
timestamp 0
transform -1 0 2110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__966_
timestamp 0
transform -1 0 370 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__972_
timestamp 0
transform -1 0 70 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__979_
timestamp 0
transform -1 0 2170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__986_
timestamp 0
transform -1 0 750 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__992_
timestamp 0
transform -1 0 490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__999_
timestamp 0
transform 1 0 410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1004_
timestamp 0
transform -1 0 1690 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1011_
timestamp 0
transform 1 0 150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1017_
timestamp 0
transform -1 0 2170 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1024_
timestamp 0
transform 1 0 1610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__1030_
timestamp 0
transform -1 0 350 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1037_
timestamp 0
transform -1 0 210 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1043_
timestamp 0
transform -1 0 2090 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__1050_
timestamp 0
transform 1 0 50 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1056_
timestamp 0
transform -1 0 350 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1063_
timestamp 0
transform -1 0 1490 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1069_
timestamp 0
transform 1 0 1470 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1076_
timestamp 0
transform 1 0 3770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1082_
timestamp 0
transform -1 0 1530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1089_
timestamp 0
transform -1 0 1650 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1096_
timestamp 0
transform -1 0 910 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1102_
timestamp 0
transform -1 0 910 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__1109_
timestamp 0
transform -1 0 1030 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__1115_
timestamp 0
transform -1 0 770 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1122_
timestamp 0
transform -1 0 210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1128_
timestamp 0
transform 1 0 1350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1135_
timestamp 0
transform 1 0 1030 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__1141_
timestamp 0
transform 1 0 630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1148_
timestamp 0
transform -1 0 3170 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1154_
timestamp 0
transform -1 0 1190 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1161_
timestamp 0
transform -1 0 350 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__1167_
timestamp 0
transform -1 0 70 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1174_
timestamp 0
transform -1 0 3230 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__1180_
timestamp 0
transform -1 0 710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1187_
timestamp 0
transform -1 0 210 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1193_
timestamp 0
transform 1 0 1250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1200_
timestamp 0
transform -1 0 1910 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__1207_
timestamp 0
transform -1 0 1210 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__1213_
timestamp 0
transform -1 0 3910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1220_
timestamp 0
transform 1 0 3050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1226_
timestamp 0
transform 1 0 2430 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__1233_
timestamp 0
transform -1 0 2530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__1239_
timestamp 0
transform -1 0 1530 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__1246_
timestamp 0
transform 1 0 850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__1252_
timestamp 0
transform -1 0 1030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1259_
timestamp 0
transform -1 0 730 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__1265_
timestamp 0
transform 1 0 210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1272_
timestamp 0
transform 1 0 2690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__1278_
timestamp 0
transform 1 0 2270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1285_
timestamp 0
transform -1 0 630 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__1291_
timestamp 0
transform 1 0 3750 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1298_
timestamp 0
transform -1 0 4010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1305_
timestamp 0
transform -1 0 4390 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1311_
timestamp 0
transform -1 0 3490 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1318_
timestamp 0
transform 1 0 2990 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1324_
timestamp 0
transform -1 0 2350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1331_
timestamp 0
transform 1 0 2210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1337_
timestamp 0
transform -1 0 1890 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__1344_
timestamp 0
transform -1 0 2050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1350_
timestamp 0
transform -1 0 1610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1357_
timestamp 0
transform -1 0 810 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__1363_
timestamp 0
transform -1 0 730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1370_
timestamp 0
transform -1 0 2730 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1376_
timestamp 0
transform -1 0 3250 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1383_
timestamp 0
transform -1 0 2830 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1389_
timestamp 0
transform 1 0 4430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1396_
timestamp 0
transform -1 0 3890 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1402_
timestamp 0
transform -1 0 2190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1409_
timestamp 0
transform -1 0 2230 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1416_
timestamp 0
transform -1 0 1530 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1422_
timestamp 0
transform 1 0 1350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1429_
timestamp 0
transform 1 0 3510 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__1435_
timestamp 0
transform -1 0 1790 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1442_
timestamp 0
transform 1 0 4290 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__1448_
timestamp 0
transform 1 0 4450 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1455_
timestamp 0
transform -1 0 3630 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__1461_
timestamp 0
transform -1 0 2590 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1468_
timestamp 0
transform -1 0 1630 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__1474_
timestamp 0
transform -1 0 1190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1481_
timestamp 0
transform 1 0 2850 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__1487_
timestamp 0
transform 1 0 2690 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__1494_
timestamp 0
transform -1 0 4030 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1500_
timestamp 0
transform 1 0 4690 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1507_
timestamp 0
transform -1 0 3210 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__1514_
timestamp 0
transform 1 0 3230 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1520_
timestamp 0
transform -1 0 950 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1527_
timestamp 0
transform 1 0 2790 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1533_
timestamp 0
transform -1 0 2570 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1540_
timestamp 0
transform 1 0 3230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1546_
timestamp 0
transform 1 0 5070 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1553_
timestamp 0
transform 1 0 5390 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__1559_
timestamp 0
transform 1 0 3590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__1566_
timestamp 0
transform 1 0 3190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__1572_
timestamp 0
transform 1 0 3110 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__1579_
timestamp 0
transform 1 0 3790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__1585_
timestamp 0
transform 1 0 3490 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__1592_
timestamp 0
transform 1 0 890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__1598_
timestamp 0
transform -1 0 5630 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__1605_
timestamp 0
transform 1 0 4970 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__1611_
timestamp 0
transform 1 0 5450 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__1618_
timestamp 0
transform 1 0 5570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__1625_
timestamp 0
transform 1 0 4550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__1631_
timestamp 0
transform -1 0 4430 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__1638_
timestamp 0
transform 1 0 5130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__1644_
timestamp 0
transform -1 0 4990 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__1651_
timestamp 0
transform 1 0 5710 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__1689_
timestamp 0
transform -1 0 5350 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1696_
timestamp 0
transform -1 0 5730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1702_
timestamp 0
transform 1 0 5610 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1709_
timestamp 0
transform -1 0 5330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__1715_
timestamp 0
transform 1 0 5130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1722_
timestamp 0
transform -1 0 5430 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1728_
timestamp 0
transform 1 0 5610 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1735_
timestamp 0
transform 1 0 5250 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1741_
timestamp 0
transform -1 0 4670 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1748_
timestamp 0
transform -1 0 4870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1755_
timestamp 0
transform 1 0 4830 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1761_
timestamp 0
transform 1 0 4090 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1768_
timestamp 0
transform -1 0 4450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__1774_
timestamp 0
transform -1 0 4070 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1781_
timestamp 0
transform 1 0 4390 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1787_
timestamp 0
transform -1 0 3790 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__1794_
timestamp 0
transform -1 0 4270 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1800_
timestamp 0
transform -1 0 3370 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1807_
timestamp 0
transform 1 0 4550 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1813_
timestamp 0
transform 1 0 4150 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__1820_
timestamp 0
transform -1 0 4070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__1826_
timestamp 0
transform -1 0 3610 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__1833_
timestamp 0
transform 1 0 2990 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1839_
timestamp 0
transform 1 0 4550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__1846_
timestamp 0
transform 1 0 1990 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1852_
timestamp 0
transform -1 0 3330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__1859_
timestamp 0
transform 1 0 3490 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1866_
timestamp 0
transform 1 0 3230 0 1 250
box -6 -8 26 248
use FILL  FILL_2__1872_
timestamp 0
transform 1 0 2870 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1879_
timestamp 0
transform -1 0 3230 0 1 730
box -6 -8 26 248
use FILL  FILL_2__1885_
timestamp 0
transform -1 0 2070 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__1892_
timestamp 0
transform -1 0 70 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert8
timestamp 0
transform -1 0 2930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert14
timestamp 0
transform 1 0 5090 0 -1 730
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert1
timestamp 0
transform 1 0 5450 0 -1 2650
box -6 -8 26 248
<< labels >>
flabel metal1 s 5822 2 5882 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 5737 5817 5743 5823 3 FreeSans 16 90 0 0 ABCmd_i[7]
port 2 nsew
flabel metal2 s 5697 5817 5703 5823 3 FreeSans 16 90 0 0 ABCmd_i[6]
port 3 nsew
flabel metal2 s 5637 5817 5643 5823 3 FreeSans 16 90 0 0 ABCmd_i[5]
port 4 nsew
flabel metal2 s 5597 5817 5603 5823 3 FreeSans 16 90 0 0 ABCmd_i[4]
port 5 nsew
flabel metal2 s 5557 5817 5563 5823 3 FreeSans 16 90 0 0 ABCmd_i[3]
port 6 nsew
flabel metal3 s 5856 2776 5864 2784 3 FreeSans 16 0 0 0 ABCmd_i[2]
port 7 nsew
flabel metal3 s 5856 5636 5864 5644 3 FreeSans 16 0 0 0 ABCmd_i[1]
port 8 nsew
flabel metal3 s 5856 5676 5864 5684 3 FreeSans 16 0 0 0 ABCmd_i[0]
port 9 nsew
flabel metal2 s 3897 -23 3903 -17 7 FreeSans 16 270 0 0 ACC_o[7]
port 10 nsew
flabel metal2 s 3857 -23 3863 -17 7 FreeSans 16 270 0 0 ACC_o[6]
port 11 nsew
flabel metal2 s 3757 -23 3763 -17 7 FreeSans 16 270 0 0 ACC_o[5]
port 12 nsew
flabel metal2 s 3497 -23 3503 -17 7 FreeSans 16 270 0 0 ACC_o[4]
port 13 nsew
flabel metal2 s 2677 -23 2683 -17 7 FreeSans 16 270 0 0 ACC_o[3]
port 14 nsew
flabel metal3 s -24 2296 -16 2304 7 FreeSans 16 0 0 0 ACC_o[2]
port 15 nsew
flabel metal3 s -24 2256 -16 2264 7 FreeSans 16 0 0 0 ACC_o[1]
port 16 nsew
flabel metal3 s -24 1556 -16 1564 7 FreeSans 16 0 0 0 ACC_o[0]
port 17 nsew
flabel metal2 s 2637 -23 2643 -17 7 FreeSans 16 270 0 0 Flag_i
port 18 nsew
flabel metal2 s 5197 5817 5203 5823 3 FreeSans 16 90 0 0 LoadA_i
port 19 nsew
flabel metal2 s 5237 5817 5243 5823 3 FreeSans 16 90 0 0 LoadB_i
port 20 nsew
flabel metal2 s 5517 5817 5523 5823 3 FreeSans 16 90 0 0 LoadCmd_i
port 21 nsew
flabel metal3 s -24 3016 -16 3024 7 FreeSans 16 0 0 0 MulH_i
port 22 nsew
flabel metal3 s -24 3476 -16 3484 7 FreeSans 16 0 0 0 MulL_i
port 23 nsew
flabel metal2 s 4717 5817 4723 5823 3 FreeSans 16 90 0 0 clk
port 24 nsew
flabel metal3 s 5856 1796 5864 1804 3 FreeSans 16 0 0 0 reset
port 25 nsew
<< properties >>
string FIXED_BBOX -40 -40 5860 5820
<< end >>
