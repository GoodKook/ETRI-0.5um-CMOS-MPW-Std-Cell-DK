magic
tech scmos
magscale 1 30
timestamp 1726646330
<< checkpaint >>
rect 18300 186927 44800 197000
rect 13915 181835 44800 186927
rect 46919 186419 142100 190000
rect 46919 181835 143266 186419
rect 6771 176042 185015 181835
rect 6771 175958 328570 176042
rect 205 167042 328570 175958
rect 205 160774 185015 167042
rect 6771 143081 185015 160774
rect 0 142100 185015 143081
rect 0 102896 190000 142100
rect -13866 102380 190000 102896
rect -25613 89180 190000 102380
rect -24170 89077 190000 89180
rect -17472 83925 190000 89077
rect 0 47900 190000 83925
rect 6771 46919 190000 47900
rect 6771 32547 185015 46919
rect 6771 31724 186496 32547
rect -4457 10781 186496 31724
rect -4457 8670 185015 10781
rect -4457 7765 35955 8670
rect 205 1458 35955 7765
rect -600 -600 630 630
rect 46919 0 142100 8670
rect 149430 7830 171960 8670
<< metal1 >>
rect 45700 132200 51200 135800
rect 139100 90300 143700 99700
rect 45700 53700 51200 57900
<< m2contact >>
rect 44200 132200 45700 135800
rect 143700 90300 145500 99700
rect 44200 53700 45700 57900
<< metal2 >>
rect 59800 140800 60200 145900
rect 73300 139800 73700 145900
rect 86800 141900 87200 145900
rect 100300 143000 100700 145900
rect 100300 142600 103500 143000
rect 81200 140400 98100 140800
rect 87800 139300 95600 139800
rect 95200 136400 95600 139300
rect 97700 136400 98100 140400
rect 100000 136400 100400 141500
rect 103100 136400 103500 142600
rect 109900 136400 110300 142600
rect 113800 141600 114200 145900
rect 110600 141200 114200 141600
rect 110600 136400 111000 141200
rect 127300 140500 127700 145900
rect 140800 143000 141200 145900
rect 114500 136400 114900 140100
rect 141700 130000 145900 130400
rect 44100 116300 49300 116700
rect 143100 116500 145900 116900
rect 44100 102800 49400 103200
rect 143200 103000 145900 103400
rect 44100 89300 47000 89700
rect 145500 90300 145900 99700
rect 48100 76200 48500 87300
rect 44100 75800 48500 76200
rect 142300 76000 145900 76400
rect 49400 62700 49800 70900
rect 44100 62300 49800 62700
rect 141200 62500 145900 62900
rect 44100 53700 44200 57900
rect 87800 51800 88100 53400
rect 76300 51400 88100 51800
rect 59800 44100 60200 51400
rect 89300 50700 89600 53400
rect 101300 50500 101600 53400
rect 73300 44100 73700 50300
rect 100300 50100 101600 50500
rect 86800 44100 87200 48800
rect 100300 44100 100700 50100
rect 101900 49200 102200 53400
rect 113600 48200 113900 53400
rect 114200 49400 114500 53400
rect 103000 47800 113900 48200
rect 115700 48200 116000 53400
rect 103000 44100 103400 47800
rect 116900 46100 117200 53400
rect 133400 49000 145900 49400
rect 116500 45700 117200 46100
rect 116500 44100 116900 45700
rect 130000 44100 130400 47800
<< m3contact >>
rect 59800 140400 61000 140800
rect 86800 141500 87800 141900
rect 99400 141500 100400 141900
rect 79800 140400 81200 140800
rect 73300 139300 74800 139800
rect 86400 139300 87800 139800
rect 109900 142600 111500 143000
rect 139900 142600 141200 143000
rect 114500 140100 115900 140500
rect 126300 140100 127700 140500
rect 141300 129000 141700 130400
rect 49300 115500 49700 116700
rect 142700 115600 143100 116900
rect 49400 102800 49800 103900
rect 142700 103000 143200 104500
rect 47000 89300 47400 90400
rect 48100 87300 48500 88400
rect 141900 76000 142300 77300
rect 49400 70900 49800 72300
rect 140800 62500 141200 63800
rect 59800 51400 60900 51800
rect 75200 51400 76300 51800
rect 73300 50300 74400 50700
rect 88500 50300 89600 50700
rect 86800 48800 87700 49200
rect 101300 48800 102200 49200
rect 114200 49000 115200 49400
rect 115700 47800 116700 48200
rect 132100 49000 133400 49400
rect 129100 47800 130400 48200
<< metal3 >>
rect 111500 142600 139900 143000
rect 87800 141500 99400 141900
rect 61000 140400 79800 140800
rect 115900 140100 126300 140500
rect 74800 139300 86400 139800
rect 49300 107200 49700 115500
rect 141300 115100 141700 129000
rect 138900 114700 141700 115100
rect 142700 114400 143100 115600
rect 138900 114000 143100 114400
rect 138900 110200 143200 110600
rect 49300 106900 51700 107200
rect 49400 106300 51700 106600
rect 49400 103900 49800 106300
rect 142700 104500 143200 110200
rect 47000 99100 51700 99400
rect 47000 90400 47400 99100
rect 48100 98500 51700 98800
rect 138800 98500 142300 98900
rect 48100 88400 48500 98500
rect 138800 94600 141200 95000
rect 49400 82900 51700 83200
rect 49400 72300 49800 82900
rect 140800 63800 141200 94600
rect 141900 77300 142300 98500
rect 60900 51400 75200 51800
rect 74400 50300 88500 50700
rect 87700 48800 101300 49200
rect 115200 49000 132100 49400
rect 116700 47800 129100 48200
use PIC  CIN_0 ~/ETRI050_DesignKit/pads_ETRI050
timestamp 1537935238
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_1
timestamp 1537935238
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_2
timestamp 1537935238
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_3
timestamp 1537935238
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_4
timestamp 1537935238
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_5
timestamp 1537935238
transform 1 0 129500 0 -1 171100
box -100 -9150 12100 25300
use PIC  CLK
timestamp 1537935238
transform 1 0 48500 0 -1 171100
box -100 -9150 12100 25300
use fir_pe_Core  fir_pe_Core_0
timestamp 1726639203
transform 1 0 51945 0 1 53660
box -945 -360 87345 82845
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/pads_ETRI050
timestamp 1725930584
transform 0 -1 171100 -1 0 75646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_1
timestamp 1725930584
transform 0 -1 171098 -1 0 62146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_2
timestamp 1725930584
transform 0 -1 171100 -1 0 102646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_3
timestamp 1725930584
transform 0 -1 171100 -1 0 89146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_4
timestamp 1725930584
transform 0 -1 171102 -1 0 129646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_5
timestamp 1725930584
transform 0 -1 171100 -1 0 116146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_6
timestamp 1725930584
transform 1 0 73845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_7
timestamp 1725930584
transform 1 0 60345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_8
timestamp 1725930584
transform 1 0 100845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_9
timestamp 1725930584
transform 1 0 87345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_10
timestamp 1725930584
transform 1 0 127845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_11
timestamp 1725930584
transform 1 0 114345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_12
timestamp 1725930584
transform 0 1 18899 -1 0 75655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_13
timestamp 1725930584
transform 0 1 18899 -1 0 62155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_14
timestamp 1725930584
transform 0 1 18900 -1 0 102655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_15
timestamp 1725930584
transform 0 1 18900 -1 0 89155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_16
timestamp 1725930584
transform 1 0 73845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_17
timestamp 1725930584
transform 0 1 18897 -1 0 116155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_18
timestamp 1725930584
transform 0 1 18900 -1 0 129655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_19
timestamp 1725930584
transform 1 0 60345 0 -1 171101
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_20
timestamp 1725930584
transform 1 0 100845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_21
timestamp 1725930584
transform 1 0 87344 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_22
timestamp 1725930584
transform 1 0 127845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_23
timestamp 1725930584
transform 1 0 114345 0 -1 171100
box -60 0 1860 25060
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1537935238
transform 1 0 43621 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1537935238
transform 1 0 141360 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1537935238
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1537935238
transform 1 0 43638 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1537935238
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1537935238
transform 0 1 18900 -1 0 146379
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1537935238
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1537935238
transform 0 -1 171100 -1 0 146346
box -35 0 5035 25060
use MY_LOGO  MY_LOGO_0
timestamp 1724157349
transform 1 0 147600 0 1 9285
box 180 225 21510 9045
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1537935238
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1537935238
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1537935238
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1537935238
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
use PIC  RDY_I
timestamp 1537935238
transform 0 1 18900 -1 0 74000
box -100 -9150 12100 25300
use PVDD  VDD_0 ~/ETRI050_DesignKit/pads_ETRI050
timestamp 1537935238
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use PVDD  VDD_1
timestamp 1537935238
transform 0 1 18900 -1 0 141500
box -100 -9150 12100 25300
use POB8  VLD_O ~/ETRI050_DesignKit/pads_ETRI050
timestamp 1537935238
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use PVSS  VSS_0 ~/ETRI050_DesignKit/pads_ETRI050
timestamp 1537935238
transform 0 -1 171100 1 0 89000
box -100 -9150 12100 25300
use PIC  XIN_0
timestamp 1537935238
transform 0 1 18900 -1 0 87500
box -100 -9150 12100 25300
use PIC  XIN_1
timestamp 1537935238
transform 0 1 18900 -1 0 101000
box -100 -9150 12100 25300
use PIC  XIN_2
timestamp 1537935238
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use PIC  XIN_3
timestamp 1537935238
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use POB8  XOUT_0
timestamp 1537935238
transform 0 -1 171100 1 0 75500
box -100 -9150 12100 25300
use POB8  XOUT_1
timestamp 1537935238
transform 0 -1 171100 1 0 102500
box -100 -9150 12100 25300
use POB8  XOUT_2
timestamp 1537935238
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
use POB8  XOUT_3
timestamp 1537935238
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
use PIC  YIN_0
timestamp 1537935238
transform 1 0 48500 0 1 18900
box -100 -9150 12100 25300
use PIC  YIN_1
timestamp 1537935238
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use PIC  YIN_2
timestamp 1537935238
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use PIC  YIN_3
timestamp 1537935238
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use POB8  YOUT_0
timestamp 1537935238
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use POB8  YOUT_1
timestamp 1537935238
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use POB8  YOUT_2
timestamp 1537935238
transform 1 0 129500 0 1 18900
box -100 -9150 12100 25300
use POB8  YOUT_3
timestamp 1537935238
transform 0 -1 171100 1 0 48500
box -100 -9150 12100 25300
<< end >>
