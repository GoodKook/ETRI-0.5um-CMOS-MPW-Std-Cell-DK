/* Verilog module written by vlog2Verilog (qflow) */
/* With bit-blasted vectors */
/* With power connections converted to binary 1, 0 */

module cpu(
    output [15:0] AB,
    input [7:0] DI,
    output [7:0] DO,
    input IRQ,
    input NMI,
    input RDY,
    output WE,
    input clk,
    input reset
);

wire C ;
wire D ;
wire I ;
wire N ;
wire V ;
wire Z ;
wire _1677_ ;
wire _1257_ ;
wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _397_ ;
wire _1295_ ;
wire _703_ ;
wire _1389_ ;
wire _19_ ;
wire _1601_ ;
wire _932_ ;
wire _512_ ;
wire _1198_ ;
wire _1410_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _1504_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _929_ ;
wire _509_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _1407_ ;
wire _738_ ;
wire _318_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _1674_ ;
wire _1254_ ;
wire _585_ ;
wire _165_ ;
wire [5:0] _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _1539_ ;
wire _1119_ ;
wire _1292_ ;
wire _1348_ ;
wire _679_ ;
wire _259_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _700_ ;
wire _1386_ ;
wire _297_ ;
wire _16_ ;
wire _1195_ ;
wire _54_ ;
wire _603_ ;
wire _1289_ ;
wire _1501_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire _1098_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire _926_ ;
wire _506_ ;
wire _1404_ ;
wire _735_ ;
wire _315_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire IRQ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _1307_ ;
wire _638_ ;
wire _218_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _1__bF$buf10 ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire WE ;
wire _1383_ ;
wire _294_ ;
wire _13_ ;
wire _1439_ ;
wire _1019_ ;
wire php ;
wire _1192_ ;
wire _1668_ ;
wire _1248_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _600_ ;
wire _1286_ ;
wire _197_ ;
wire _1095_ ;
wire _7_ ;
wire RDY ;
wire _923_ ;
wire _503_ ;
wire _1189_ ;
wire _1401_ ;
wire _732_ ;
wire _312_ ;
wire adc_sbc ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _1304_ ;
wire _635_ ;
wire _215_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _1627_ ;
wire _1207_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _1380_ ;
wire _291_ ;
wire _10_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire _887__bF$buf0 ;
wire _887__bF$buf1 ;
wire _887__bF$buf2 ;
wire _887__bF$buf3 ;
wire _887__bF$buf4 ;
wire _1283_ ;
wire _194_ ;
wire _1339_ ;
wire _1092_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire write_back ;
wire _1377_ ;
wire _288_ ;
wire _4_ ;
wire _920_ ;
wire _500_ ;
wire _1186_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _1089_ ;
wire _1301_ ;
wire _632_ ;
wire _212_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _1624_ ;
wire _1204_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _1527_ ;
wire _1107_ ;
wire _858_ ;
wire _438_ ;
wire _1280_ ;
wire _191_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _1374_ ;
wire _285_ ;
wire _1_ ;
wire index_y ;
wire _1183_ ;
wire _1659_ ;
wire _1239_ ;
wire _42_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _1277_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _1086_ ;
wire _914_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire clc ;
wire cld ;
wire cli ;
wire clk ;
wire clv ;
wire _817_ ;
wire _77_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _1618_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _1371_ ;
wire _282_ ;
wire _1427_ ;
wire _1007_ ;
wire _758_ ;
wire _338_ ;
wire _1180_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _1274_ ;
wire _185_ ;
wire _1083_ ;
wire _1559_ ;
wire _1139_ ;
wire _830__bF$buf0 ;
wire _830__bF$buf1 ;
wire _830__bF$buf2 ;
wire _830__bF$buf3 ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire _1597_ ;
wire _1177_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _908_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _1615_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _1518_ ;
wire _849_ ;
wire _429_ ;
wire _1271_ ;
wire _182_ ;
wire _1327_ ;
wire _658_ ;
wire _238_ ;
wire _1080_ ;
wire IRHOLD_valid_bF$buf0 ;
wire IRHOLD_valid_bF$buf1 ;
wire IRHOLD_valid_bF$buf2 ;
wire IRHOLD_valid_bF$buf3 ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _1594_ ;
wire _1174_ ;
wire HC ;
wire _33_ ;
wire _1459_ ;
wire _1039_ ;
wire _1268_ ;
wire _691__bF$buf0 ;
wire _691__bF$buf1 ;
wire _691__bF$buf2 ;
wire _691__bF$buf3 ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _620_ ;
wire _200_ ;
wire _905_ ;
wire _714_ ;
wire [7:0] ADD ;
wire _1612_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _1609_ ;
wire _1362_ ;
wire RDY_bF$buf0 ;
wire RDY_bF$buf1 ;
wire RDY_bF$buf2 ;
wire RDY_bF$buf3 ;
wire RDY_bF$buf4 ;
wire RDY_bF$buf5 ;
wire RDY_bF$buf6 ;
wire RDY_bF$buf7 ;
wire RDY_bF$buf8 ;
wire _693_ ;
wire _273_ ;
wire _1418_ ;
wire _749_ ;
wire _329_ ;
wire _1591_ ;
wire _1171_ ;
wire _1647_ ;
wire _1227_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _1456_ ;
wire _1036_ ;
wire res ;
wire _787_ ;
wire _367_ ;
wire rotate ;
wire [15:0] _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _1494_ ;
wire _1074_ ;
wire [3:0] alu_op ;
wire _1359_ ;
wire _902_ ;
wire _1588_ ;
wire _1168_ ;
wire _499_ ;
wire _711_ ;
wire _1397_ ;
wire _27_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire [1:0] dst_reg ;
wire \u_ALU8.BI7  ;
wire _805_ ;
wire [7:0] DIHOLD ;
wire _65_ ;
wire _614_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _1606_ ;
wire _937_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire [7:0] BI ;
wire _1453_ ;
wire _1033_ ;
wire _918__bF$buf0 ;
wire _918__bF$buf1 ;
wire _918__bF$buf2 ;
wire _918__bF$buf3 ;
wire _784_ ;
wire _364_ ;
wire _1509_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _1318_ ;
wire _649_ ;
wire _229_ ;
wire _1491_ ;
wire _1071_ ;
wire _1547_ ;
wire _1127_ ;
wire _878_ ;
wire _458_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _1394_ ;
wire _24_ ;
wire _1679_ ;
wire _1259_ ;
wire _802_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _399_ ;
wire _611_ ;
wire _1297_ ;
wire _840_ ;
wire _420_ ;
wire \u_ALU8.AI7  ;
wire _705_ ;
wire _1603_ ;
wire _934_ ;
wire _514_ ;
wire _1412_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _1506_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire _1544_ ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire \u_ALU8.BCD  ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _1409_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _1638_ ;
wire _1218_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _1391_ ;
wire _21_ ;
wire _1447_ ;
wire _1027_ ;
wire _778_ ;
wire _358_ ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _1485_ ;
wire _1065_ ;
wire _396_ ;
wire _1294_ ;
wire [7:0] \AXYS[1]  ;
wire _1579_ ;
wire _1159_ ;
wire _702_ ;
wire _1388_ ;
wire _299_ ;
wire _18_ ;
wire _1600_ ;
wire _931_ ;
wire _511_ ;
wire _1197_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _1503_ ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _928_ ;
wire _508_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _1406_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _1309_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _1538_ ;
wire _1118_ ;
wire _869_ ;
wire _449_ ;
wire _1291_ ;
wire _1347_ ;
wire _678_ ;
wire _258_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _1385_ ;
wire _296_ ;
wire _15_ ;
wire _1194_ ;
wire _1129__bF$buf0 ;
wire _1129__bF$buf1 ;
wire _1129__bF$buf2 ;
wire _1129__bF$buf3 ;
wire _1129__bF$buf4 ;
wire _853__bF$buf0 ;
wire _853__bF$buf1 ;
wire _853__bF$buf2 ;
wire _853__bF$buf3 ;
wire _853__bF$buf4 ;
wire _853__bF$buf5 ;
wire _853__bF$buf6 ;
wire _853__bF$buf7 ;
wire _53_ ;
wire _1479_ ;
wire _1059_ ;
wire store ;
wire _602_ ;
wire _1288_ ;
wire _199_ ;
wire _1500_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _1097_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _925_ ;
wire _505_ ;
wire IRHOLD_valid ;
wire _1403_ ;
wire _734_ ;
wire _314_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _1306_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _1629_ ;
wire _1209_ ;
wire _1382_ ;
wire _293_ ;
wire _12_ ;
wire _1438_ ;
wire _1018_ ;
wire _769_ ;
wire _349_ ;
wire _1191_ ;
wire _1667_ ;
wire _1247_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _1002__bF$buf0 ;
wire _1002__bF$buf1 ;
wire _1002__bF$buf2 ;
wire _1002__bF$buf3 ;
wire _1002__bF$buf4 ;
wire _50_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _1285_ ;
wire _196_ ;
wire _1094_ ;
wire _1379_ ;
wire _6_ ;
wire _922_ ;
wire _502_ ;
wire _1188_ ;
wire _1400_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _1303_ ;
wire _634_ ;
wire _214_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _1__bF$buf0 ;
wire _1__bF$buf1 ;
wire _1__bF$buf2 ;
wire _1__bF$buf3 ;
wire _1__bF$buf4 ;
wire _1__bF$buf5 ;
wire _1__bF$buf6 ;
wire _1__bF$buf7 ;
wire _1__bF$buf8 ;
wire _1__bF$buf9 ;
wire _919_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _1626_ ;
wire _1206_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire backwards ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _1529_ ;
wire _1109_ ;
wire _1282_ ;
wire _193_ ;
wire _1338_ ;
wire _669_ ;
wire _249_ ;
wire _1091_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _1376_ ;
wire _287_ ;
wire _3_ ;
wire _1185_ ;
wire _44_ ;
wire _1279_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _1088_ ;
wire _1300_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _916_ ;
wire _926__bF$buf0 ;
wire _926__bF$buf1 ;
wire _926__bF$buf2 ;
wire _926__bF$buf3 ;
wire _725_ ;
wire _305_ ;
wire [15:0] PC ;
wire _1623_ ;
wire _1203_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _1432_ ;
wire _1012_ ;
wire _882__bF$buf0 ;
wire _882__bF$buf1 ;
wire _882__bF$buf2 ;
wire _882__bF$buf3 ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _1373_ ;
wire _284_ ;
wire _0_ ;
wire _1429_ ;
wire _1009_ ;
wire _1182_ ;
wire _1658_ ;
wire _1238_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire adj_bcd ;
wire _41_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _1276_ ;
wire _187_ ;
wire _1085_ ;
wire _913_ ;
wire [7:0] \AXYS[3]  ;
wire _1599_ ;
wire _1179_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire compare ;
wire _816_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire load_only ;
wire clk_bF$buf10 ;
wire shift ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _1617_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _1370_ ;
wire _281_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire [1:0] src_reg ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _1273_ ;
wire _184_ ;
wire _1329_ ;
wire _1082_ ;
wire _1558_ ;
wire _1138_ ;
wire _889_ ;
wire _469_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _1596_ ;
wire _1176_ ;
wire _869__bF$buf0 ;
wire _869__bF$buf1 ;
wire _869__bF$buf2 ;
wire _869__bF$buf3 ;
wire _35_ ;
wire _813_ ;
wire _73_ ;
wire _1499_ ;
wire _1079_ ;
wire _622_ ;
wire _202_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _1614_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _1517_ ;
wire _848_ ;
wire _428_ ;
wire _1270_ ;
wire _181_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _1593_ ;
wire _1173_ ;
wire _1649_ ;
wire _1229_ ;
wire _32_ ;
wire _1458_ ;
wire _1038_ ;
wire [2:0] cond_code ;
wire _789_ ;
wire _369_ ;
wire _1687_ ;
wire _1267_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _904_ ;
wire _713_ ;
wire _1399_ ;
wire _29_ ;
wire _1611_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire [5:0] state ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire bit_ins ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _1608_ ;
wire _939_ ;
wire _519_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _1417_ ;
wire _748_ ;
wire _328_ ;
wire _1590_ ;
wire _1170_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire [7:0] DI ;
wire [7:0] DO ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _1493_ ;
wire _1073_ ;
wire _1549_ ;
wire _1129_ ;
wire _1358_ ;
wire _689_ ;
wire _269_ ;
wire _901_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _710_ ;
wire _1396_ ;
wire _26_ ;
wire _804_ ;
wire _64_ ;
wire _613_ ;
wire _1299_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _1605_ ;
wire _936_ ;
wire _516_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire [15:0] AB ;
wire [7:0] AI ;
wire AN ;
wire AV ;
wire AZ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _1508_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _1317_ ;
wire _648_ ;
wire _228_ ;
wire _1490_ ;
wire _1070_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _1393_ ;
wire _23_ ;
wire _1449_ ;
wire _1029_ ;
wire _1678_ ;
wire _1258_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _610_ ;
wire _1296_ ;
wire _886__bF$buf0 ;
wire _886__bF$buf1 ;
wire _886__bF$buf2 ;
wire _886__bF$buf3 ;
wire _704_ ;
wire _1602_ ;
wire _933_ ;
wire _513_ ;
wire _1199_ ;
wire _1411_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _1640_ ;
wire _1220_ ;
wire _1051__bF$buf0 ;
wire _1051__bF$buf1 ;
wire _1051__bF$buf2 ;
wire _1051__bF$buf3 ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _1505_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire NMI ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _1408_ ;
wire _739_ ;
wire _319_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _1637_ ;
wire _1217_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _1390_ ;
wire _20_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire _1293_ ;
wire _1349_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _701_ ;
wire _1387_ ;
wire _298_ ;
wire _17_ ;
wire _930_ ;
wire _510_ ;
wire plp ;
wire _1196_ ;
wire _55_ ;
wire _604_ ;
wire _1502_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _1099_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _927_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _1405_ ;
wire _736_ ;
wire _316_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _1308_ ;
wire _639_ ;
wire _219_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire _1537_ ;
wire _1117_ ;
wire _868_ ;
wire _448_ ;
wire _1290_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _1384_ ;
wire _295_ ;
wire _14_ ;
wire _1193_ ;
wire _1669_ ;
wire _1249_ ;
wire _52_ ;
wire _1478_ ;
wire _1058_ ;
wire _389_ ;
wire _601_ ;
wire _1287_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _1096_ ;
wire _8_ ;
wire _924_ ;
wire _504_ ;
wire _1402_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _1305_ ;
wire _636_ ;
wire _216_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _1628_ ;
wire _1208_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _1381_ ;
wire _292_ ;
wire _11_ ;
wire _1437_ ;
wire _1017_ ;
wire _768_ ;
wire _348_ ;
wire _1190_ ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire _1284_ ;
wire _195_ ;
wire _1093_ ;
wire [7:0] \AXYS[0]  ;
wire _1569_ ;
wire _1149_ ;
wire _1378_ ;
wire _289_ ;
wire _5_ ;
wire _921_ ;
wire _501_ ;
wire _1187_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _1302_ ;
wire _633_ ;
wire _213_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _918_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _1625_ ;
wire _1205_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _1528_ ;
wire _1108_ ;
wire shift_right ;
wire _859_ ;
wire _439_ ;
wire _1281_ ;
wire _192_ ;
wire _1337_ ;
wire _668_ ;
wire _248_ ;
wire _1090_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _1375_ ;
wire _286_ ;
wire _2_ ;
wire _1184_ ;
wire _43_ ;
wire _1469_ ;
wire _1049_ ;
wire [7:0] DIMUX ;
wire _1278_ ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _1087_ ;
wire [3:0] op ;
wire _630_ ;
wire _210_ ;
wire _915_ ;
wire _724_ ;
wire _304_ ;
wire _1622_ ;
wire _1202_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _1619_ ;
wire _1372_ ;
wire _283_ ;
wire _1428_ ;
wire _1008_ ;
wire _759_ ;
wire _339_ ;
wire _1181_ ;
wire _1657_ ;
wire _1237_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire sec ;
wire sed ;
wire sei ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire [7:0] IRHOLD ;
wire _1275_ ;
wire _186_ ;
wire alu_shift_right ;
wire _1084_ ;
wire _1369_ ;
wire _912_ ;
wire _1598_ ;
wire _1178_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _909_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _1616_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _374_ ;
wire _1519_ ;
wire _1272_ ;
wire _183_ ;
wire _1328_ ;
wire _659_ ;
wire _239_ ;
wire _1081_ ;
wire _1557_ ;
wire _1137_ ;
wire _888_ ;
wire _468_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _1595_ ;
wire _1175_ ;
wire _34_ ;
wire _1269_ ;
wire NMI_1 ;
wire _812_ ;
wire _72_ ;
wire _1649__bF$buf0 ;
wire _1649__bF$buf1 ;
wire _1649__bF$buf2 ;
wire _1498_ ;
wire _1649__bF$buf3 ;
wire _1078_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _906_ ;
wire _715_ ;
wire _1613_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _1219__bF$buf0 ;
wire _1219__bF$buf1 ;
wire _1219__bF$buf2 ;
wire _1219__bF$buf3 ;
wire adc_bcd ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _1419_ ;
wire _1592_ ;
wire _1172_ ;
wire _1648_ ;
wire _1228_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _1457_ ;
wire _1037_ ;
wire _788_ ;
wire _368_ ;
wire [7:0] _1686_ ;
wire _1266_ ;
wire _597_ ;
wire _177_ ;
wire _1495_ ;
wire _1075_ ;
wire _903_ ;
wire [7:0] \AXYS[2]  ;
wire _1589_ ;
wire _1169_ ;
wire _712_ ;
wire [7:0] ABH ;
wire [7:0] ABL ;
wire _1398_ ;
wire _28_ ;
wire _1610_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire NMI_edge ;
wire _806_ ;
wire _66_ ;
wire _615_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire load_reg ;
wire _709_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _1607_ ;
wire _938_ ;
wire _518_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire CI ;
wire CO ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _1319_ ;
wire _1492_ ;
wire _1072_ ;
wire inc ;
wire _1548_ ;
wire _1128_ ;
wire _879_ ;
wire _459_ ;
wire _1357_ ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire _1395_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _1489_ ;
wire _1069_ ;
wire _612_ ;
wire _1298_ ;
wire reset ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _1604_ ;
wire _935_ ;
wire _515_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _1507_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _1639_ ;
wire _1219_ ;
wire _1392_ ;
wire _22_ ;
wire _1448_ ;
wire _1028_ ;
wire _779_ ;
wire _359_ ;

BUFX2 BUFX2_insert97 (
    .A(_1219_),
    .Y(_1219__bF$buf0)
);

BUFX2 BUFX2_insert96 (
    .A(_1219_),
    .Y(_1219__bF$buf1)
);

BUFX2 BUFX2_insert95 (
    .A(_1219_),
    .Y(_1219__bF$buf2)
);

BUFX2 BUFX2_insert94 (
    .A(_1219_),
    .Y(_1219__bF$buf3)
);

BUFX2 BUFX2_insert93 (
    .A(_691_),
    .Y(_691__bF$buf0)
);

BUFX2 BUFX2_insert92 (
    .A(_691_),
    .Y(_691__bF$buf1)
);

BUFX2 BUFX2_insert91 (
    .A(_691_),
    .Y(_691__bF$buf2)
);

BUFX2 BUFX2_insert90 (
    .A(_691_),
    .Y(_691__bF$buf3)
);

BUFX2 BUFX2_insert89 (
    .A(_882_),
    .Y(_882__bF$buf0)
);

BUFX2 BUFX2_insert88 (
    .A(_882_),
    .Y(_882__bF$buf1)
);

BUFX2 BUFX2_insert87 (
    .A(_882_),
    .Y(_882__bF$buf2)
);

BUFX2 BUFX2_insert86 (
    .A(_882_),
    .Y(_882__bF$buf3)
);

BUFX2 BUFX2_insert85 (
    .A(_1002_),
    .Y(_1002__bF$buf0)
);

BUFX2 BUFX2_insert84 (
    .A(_1002_),
    .Y(_1002__bF$buf1)
);

BUFX2 BUFX2_insert83 (
    .A(_1002_),
    .Y(_1002__bF$buf2)
);

BUFX2 BUFX2_insert82 (
    .A(_1002_),
    .Y(_1002__bF$buf3)
);

BUFX2 BUFX2_insert81 (
    .A(_1002_),
    .Y(_1002__bF$buf4)
);

BUFX2 BUFX2_insert80 (
    .A(_853_),
    .Y(_853__bF$buf0)
);

BUFX2 BUFX2_insert79 (
    .A(_853_),
    .Y(_853__bF$buf1)
);

BUFX2 BUFX2_insert78 (
    .A(_853_),
    .Y(_853__bF$buf2)
);

BUFX2 BUFX2_insert77 (
    .A(_853_),
    .Y(_853__bF$buf3)
);

BUFX2 BUFX2_insert76 (
    .A(_853_),
    .Y(_853__bF$buf4)
);

BUFX2 BUFX2_insert75 (
    .A(_853_),
    .Y(_853__bF$buf5)
);

BUFX2 BUFX2_insert74 (
    .A(_853_),
    .Y(_853__bF$buf6)
);

BUFX2 BUFX2_insert73 (
    .A(_853_),
    .Y(_853__bF$buf7)
);

BUFX2 BUFX2_insert72 (
    .A(_918_),
    .Y(_918__bF$buf0)
);

BUFX2 BUFX2_insert71 (
    .A(_918_),
    .Y(_918__bF$buf1)
);

BUFX2 BUFX2_insert70 (
    .A(_918_),
    .Y(_918__bF$buf2)
);

BUFX2 BUFX2_insert69 (
    .A(_918_),
    .Y(_918__bF$buf3)
);

BUFX2 BUFX2_insert68 (
    .A(_830_),
    .Y(_830__bF$buf0)
);

BUFX2 BUFX2_insert67 (
    .A(_830_),
    .Y(_830__bF$buf1)
);

BUFX2 BUFX2_insert66 (
    .A(_830_),
    .Y(_830__bF$buf2)
);

BUFX2 BUFX2_insert65 (
    .A(_830_),
    .Y(_830__bF$buf3)
);

BUFX2 BUFX2_insert64 (
    .A(_1129_),
    .Y(_1129__bF$buf0)
);

BUFX2 BUFX2_insert63 (
    .A(_1129_),
    .Y(_1129__bF$buf1)
);

BUFX2 BUFX2_insert62 (
    .A(_1129_),
    .Y(_1129__bF$buf2)
);

BUFX2 BUFX2_insert61 (
    .A(_1129_),
    .Y(_1129__bF$buf3)
);

BUFX2 BUFX2_insert60 (
    .A(_1129_),
    .Y(_1129__bF$buf4)
);

BUFX2 BUFX2_insert59 (
    .A(_1649_),
    .Y(_1649__bF$buf0)
);

BUFX2 BUFX2_insert58 (
    .A(_1649_),
    .Y(_1649__bF$buf1)
);

BUFX2 BUFX2_insert57 (
    .A(_1649_),
    .Y(_1649__bF$buf2)
);

BUFX2 BUFX2_insert56 (
    .A(_1649_),
    .Y(_1649__bF$buf3)
);

BUFX2 BUFX2_insert55 (
    .A(_886_),
    .Y(_886__bF$buf0)
);

BUFX2 BUFX2_insert54 (
    .A(_886_),
    .Y(_886__bF$buf1)
);

BUFX2 BUFX2_insert53 (
    .A(_886_),
    .Y(_886__bF$buf2)
);

BUFX2 BUFX2_insert52 (
    .A(_886_),
    .Y(_886__bF$buf3)
);

BUFX2 BUFX2_insert51 (
    .A(IRHOLD_valid),
    .Y(IRHOLD_valid_bF$buf0)
);

BUFX2 BUFX2_insert50 (
    .A(IRHOLD_valid),
    .Y(IRHOLD_valid_bF$buf1)
);

BUFX2 BUFX2_insert49 (
    .A(IRHOLD_valid),
    .Y(IRHOLD_valid_bF$buf2)
);

BUFX2 BUFX2_insert48 (
    .A(IRHOLD_valid),
    .Y(IRHOLD_valid_bF$buf3)
);

BUFX2 BUFX2_insert47 (
    .A(_869_),
    .Y(_869__bF$buf0)
);

BUFX2 BUFX2_insert46 (
    .A(_869_),
    .Y(_869__bF$buf1)
);

BUFX2 BUFX2_insert45 (
    .A(_869_),
    .Y(_869__bF$buf2)
);

BUFX2 BUFX2_insert44 (
    .A(_869_),
    .Y(_869__bF$buf3)
);

BUFX2 BUFX2_insert43 (
    .A(_887_),
    .Y(_887__bF$buf0)
);

BUFX2 BUFX2_insert42 (
    .A(_887_),
    .Y(_887__bF$buf1)
);

BUFX2 BUFX2_insert41 (
    .A(_887_),
    .Y(_887__bF$buf2)
);

BUFX2 BUFX2_insert40 (
    .A(_887_),
    .Y(_887__bF$buf3)
);

BUFX2 BUFX2_insert39 (
    .A(_887_),
    .Y(_887__bF$buf4)
);

CLKBUF1 CLKBUF1_insert38 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert37 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert36 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert35 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert34 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert33 (
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert32 (
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert31 (
    .A(clk),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert30 (
    .A(clk),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert29 (
    .A(clk),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert28 (
    .A(clk),
    .Y(clk_bF$buf10)
);

BUFX2 BUFX2_insert27 (
    .A(_1_),
    .Y(_1__bF$buf0)
);

BUFX2 BUFX2_insert26 (
    .A(_1_),
    .Y(_1__bF$buf1)
);

BUFX2 BUFX2_insert25 (
    .A(_1_),
    .Y(_1__bF$buf2)
);

BUFX2 BUFX2_insert24 (
    .A(_1_),
    .Y(_1__bF$buf3)
);

BUFX2 BUFX2_insert23 (
    .A(_1_),
    .Y(_1__bF$buf4)
);

BUFX2 BUFX2_insert22 (
    .A(_1_),
    .Y(_1__bF$buf5)
);

BUFX2 BUFX2_insert21 (
    .A(_1_),
    .Y(_1__bF$buf6)
);

BUFX2 BUFX2_insert20 (
    .A(_1_),
    .Y(_1__bF$buf7)
);

BUFX2 BUFX2_insert19 (
    .A(_1_),
    .Y(_1__bF$buf8)
);

BUFX2 BUFX2_insert18 (
    .A(_1_),
    .Y(_1__bF$buf9)
);

BUFX2 BUFX2_insert17 (
    .A(_1_),
    .Y(_1__bF$buf10)
);

BUFX2 BUFX2_insert16 (
    .A(_1051_),
    .Y(_1051__bF$buf0)
);

BUFX2 BUFX2_insert15 (
    .A(_1051_),
    .Y(_1051__bF$buf1)
);

BUFX2 BUFX2_insert14 (
    .A(_1051_),
    .Y(_1051__bF$buf2)
);

BUFX2 BUFX2_insert13 (
    .A(_1051_),
    .Y(_1051__bF$buf3)
);

BUFX2 BUFX2_insert12 (
    .A(RDY),
    .Y(RDY_bF$buf0)
);

BUFX2 BUFX2_insert11 (
    .A(RDY),
    .Y(RDY_bF$buf1)
);

BUFX2 BUFX2_insert10 (
    .A(RDY),
    .Y(RDY_bF$buf2)
);

BUFX2 BUFX2_insert9 (
    .A(RDY),
    .Y(RDY_bF$buf3)
);

BUFX2 BUFX2_insert8 (
    .A(RDY),
    .Y(RDY_bF$buf4)
);

BUFX2 BUFX2_insert7 (
    .A(RDY),
    .Y(RDY_bF$buf5)
);

BUFX2 BUFX2_insert6 (
    .A(RDY),
    .Y(RDY_bF$buf6)
);

BUFX2 BUFX2_insert5 (
    .A(RDY),
    .Y(RDY_bF$buf7)
);

BUFX2 BUFX2_insert4 (
    .A(RDY),
    .Y(RDY_bF$buf8)
);

BUFX2 BUFX2_insert3 (
    .A(_926_),
    .Y(_926__bF$buf0)
);

BUFX2 BUFX2_insert2 (
    .A(_926_),
    .Y(_926__bF$buf1)
);

BUFX2 BUFX2_insert1 (
    .A(_926_),
    .Y(_926__bF$buf2)
);

BUFX2 BUFX2_insert0 (
    .A(_926_),
    .Y(_926__bF$buf3)
);

INVX1 _1688_ (
    .A(DIHOLD[0]),
    .Y(_849_)
);

NAND2X1 _1689_ (
    .A(DI[0]),
    .B(RDY_bF$buf8),
    .Y(_850_)
);

OAI21X1 _1690_ (
    .A(RDY_bF$buf7),
    .B(_849_),
    .C(_850_),
    .Y(DIMUX[0])
);

INVX1 _1691_ (
    .A(DIHOLD[1]),
    .Y(_851_)
);

NAND2X1 _1692_ (
    .A(RDY_bF$buf6),
    .B(DI[1]),
    .Y(_852_)
);

OAI21X1 _1693_ (
    .A(RDY_bF$buf5),
    .B(_851_),
    .C(_852_),
    .Y(DIMUX[1])
);

INVX8 _1694_ (
    .A(RDY_bF$buf4),
    .Y(_853_)
);

OR2X2 _1695_ (
    .A(RDY_bF$buf3),
    .B(DIHOLD[2]),
    .Y(_854_)
);

OAI21X1 _1696_ (
    .A(_853__bF$buf7),
    .B(DI[2]),
    .C(_854_),
    .Y(_855_)
);

INVX1 _1697_ (
    .A(_855_),
    .Y(DIMUX[2])
);

OR2X2 _1698_ (
    .A(RDY_bF$buf2),
    .B(DIHOLD[3]),
    .Y(_856_)
);

OAI21X1 _1699_ (
    .A(_853__bF$buf6),
    .B(DI[3]),
    .C(_856_),
    .Y(_857_)
);

INVX1 _1700_ (
    .A(_857_),
    .Y(DIMUX[3])
);

OR2X2 _1701_ (
    .A(RDY_bF$buf1),
    .B(DIHOLD[4]),
    .Y(_858_)
);

OAI21X1 _1702_ (
    .A(_853__bF$buf5),
    .B(DI[4]),
    .C(_858_),
    .Y(_859_)
);

INVX1 _1703_ (
    .A(_859_),
    .Y(DIMUX[4])
);

OR2X2 _1704_ (
    .A(RDY_bF$buf0),
    .B(DIHOLD[5]),
    .Y(_860_)
);

OAI21X1 _1705_ (
    .A(_853__bF$buf4),
    .B(DI[5]),
    .C(_860_),
    .Y(_861_)
);

INVX1 _1706_ (
    .A(_861_),
    .Y(DIMUX[5])
);

OR2X2 _1707_ (
    .A(RDY_bF$buf8),
    .B(DIHOLD[6]),
    .Y(_862_)
);

OAI21X1 _1708_ (
    .A(_853__bF$buf3),
    .B(DI[6]),
    .C(_862_),
    .Y(_863_)
);

INVX1 _1709_ (
    .A(_863_),
    .Y(DIMUX[6])
);

MUX2X1 _1710_ (
    .A(DI[7]),
    .B(DIHOLD[7]),
    .S(RDY_bF$buf7),
    .Y(_864_)
);

INVX1 _1711_ (
    .A(_864_),
    .Y(DIMUX[7])
);

INVX1 _1712_ (
    .A(CO),
    .Y(_865_)
);

INVX1 _1713_ (
    .A(state[3]),
    .Y(_866_)
);

NAND2X1 _1714_ (
    .A(state[2]),
    .B(_866_),
    .Y(_867_)
);

INVX1 _1715_ (
    .A(_867_),
    .Y(_868_)
);

NOR2X1 _1716_ (
    .A(state[5]),
    .B(state[4]),
    .Y(_869_)
);

INVX1 _1717_ (
    .A(state[1]),
    .Y(_870_)
);

NOR2X1 _1718_ (
    .A(state[0]),
    .B(_870_),
    .Y(_871_)
);

NAND3X1 _1719_ (
    .A(_869__bF$buf3),
    .B(_871_),
    .C(_868_),
    .Y(_872_)
);

INVX1 _1720_ (
    .A(state[2]),
    .Y(_873_)
);

NAND2X1 _1721_ (
    .A(_873_),
    .B(_866_),
    .Y(_874_)
);

NAND2X1 _1722_ (
    .A(state[1]),
    .B(state[0]),
    .Y(_875_)
);

NOR2X1 _1723_ (
    .A(_875_),
    .B(_874_),
    .Y(_876_)
);

NAND2X1 _1724_ (
    .A(_869__bF$buf2),
    .B(_876_),
    .Y(_877_)
);

INVX1 _1725_ (
    .A(_877_),
    .Y(_878_)
);

NOR2X1 _1726_ (
    .A(state[1]),
    .B(state[0]),
    .Y(_879_)
);

NAND2X1 _1727_ (
    .A(_879_),
    .B(_868_),
    .Y(_880_)
);

INVX2 _1728_ (
    .A(state[5]),
    .Y(_881_)
);

NAND2X1 _1729_ (
    .A(state[4]),
    .B(_881_),
    .Y(_882_)
);

NOR2X1 _1730_ (
    .A(_882__bF$buf3),
    .B(_880_),
    .Y(_883_)
);

NOR2X1 _1731_ (
    .A(_883_),
    .B(_878_),
    .Y(_884_)
);

AND2X2 _1732_ (
    .A(_884_),
    .B(_872_),
    .Y(_885_)
);

NOR2X1 _1733_ (
    .A(state[4]),
    .B(_881_),
    .Y(_886_)
);

INVX8 _1734_ (
    .A(_886__bF$buf3),
    .Y(_887_)
);

INVX1 _1735_ (
    .A(state[0]),
    .Y(_888_)
);

NAND2X1 _1736_ (
    .A(state[1]),
    .B(_888_),
    .Y(_889_)
);

NOR2X1 _1737_ (
    .A(_867_),
    .B(_889_),
    .Y(_890_)
);

INVX2 _1738_ (
    .A(_890_),
    .Y(_891_)
);

NAND2X1 _1739_ (
    .A(state[3]),
    .B(_873_),
    .Y(_892_)
);

NOR2X1 _1740_ (
    .A(_889_),
    .B(_892_),
    .Y(_893_)
);

NAND2X1 _1741_ (
    .A(_886__bF$buf2),
    .B(_893_),
    .Y(_894_)
);

OAI21X1 _1742_ (
    .A(_887__bF$buf4),
    .B(_891_),
    .C(_894_),
    .Y(_895_)
);

NAND2X1 _1743_ (
    .A(state[2]),
    .B(state[3]),
    .Y(_896_)
);

NOR2X1 _1744_ (
    .A(_875_),
    .B(_896_),
    .Y(_897_)
);

NAND2X1 _1745_ (
    .A(_869__bF$buf1),
    .B(_897_),
    .Y(_898_)
);

NAND2X1 _1746_ (
    .A(state[0]),
    .B(_870_),
    .Y(_899_)
);

NOR2X1 _1747_ (
    .A(_867_),
    .B(_899_),
    .Y(_900_)
);

INVX1 _1748_ (
    .A(_900_),
    .Y(_901_)
);

OAI21X1 _1749_ (
    .A(_887__bF$buf3),
    .B(_901_),
    .C(_898_),
    .Y(_902_)
);

NOR2X1 _1750_ (
    .A(_902_),
    .B(_895_),
    .Y(_903_)
);

OAI21X1 _1751_ (
    .A(_865_),
    .B(_885_),
    .C(_903_),
    .Y(_904_)
);

NOR2X1 _1752_ (
    .A(_875_),
    .B(_867_),
    .Y(_905_)
);

NOR2X1 _1753_ (
    .A(_875_),
    .B(_892_),
    .Y(_906_)
);

OAI21X1 _1754_ (
    .A(_905_),
    .B(_906_),
    .C(_886__bF$buf1),
    .Y(_907_)
);

INVX1 _1755_ (
    .A(rotate),
    .Y(_908_)
);

NAND2X1 _1756_ (
    .A(_870_),
    .B(_888_),
    .Y(_909_)
);

NOR2X1 _1757_ (
    .A(_867_),
    .B(_909_),
    .Y(_910_)
);

OAI21X1 _1758_ (
    .A(_876_),
    .B(_910_),
    .C(_886__bF$buf0),
    .Y(_911_)
);

INVX1 _1759_ (
    .A(shift),
    .Y(_912_)
);

AOI21X1 _1760_ (
    .A(_912_),
    .B(inc),
    .C(rotate),
    .Y(_913_)
);

AND2X2 _1761_ (
    .A(state[2]),
    .B(state[3]),
    .Y(_914_)
);

NOR2X1 _1762_ (
    .A(state[1]),
    .B(_888_),
    .Y(_915_)
);

NAND2X1 _1763_ (
    .A(_914_),
    .B(_915_),
    .Y(_916_)
);

INVX4 _1764_ (
    .A(state[4]),
    .Y(_917_)
);

NAND2X1 _1765_ (
    .A(_881_),
    .B(_917_),
    .Y(_918_)
);

NOR2X1 _1766_ (
    .A(_918__bF$buf3),
    .B(_916_),
    .Y(_919_)
);

INVX1 _1767_ (
    .A(compare),
    .Y(_920_)
);

NAND2X1 _1768_ (
    .A(C),
    .B(_912_),
    .Y(_921_)
);

OAI21X1 _1769_ (
    .A(load_only),
    .B(_921_),
    .C(_920_),
    .Y(_922_)
);

OAI21X1 _1770_ (
    .A(rotate),
    .B(_922_),
    .C(_919_),
    .Y(_923_)
);

OAI21X1 _1771_ (
    .A(_911_),
    .B(_913_),
    .C(_923_),
    .Y(_924_)
);

OAI21X1 _1772_ (
    .A(C),
    .B(_908_),
    .C(_924_),
    .Y(_925_)
);

NOR2X1 _1773_ (
    .A(state[5]),
    .B(_917_),
    .Y(_926_)
);

NOR2X1 _1774_ (
    .A(_889_),
    .B(_874_),
    .Y(_927_)
);

NOR2X1 _1775_ (
    .A(_896_),
    .B(_889_),
    .Y(_928_)
);

OAI21X1 _1776_ (
    .A(_928_),
    .B(_927_),
    .C(_926__bF$buf3),
    .Y(_929_)
);

NAND3X1 _1777_ (
    .A(_907_),
    .B(_929_),
    .C(_925_),
    .Y(_930_)
);

OR2X2 _1778_ (
    .A(_904_),
    .B(_930_),
    .Y(CI)
);

INVX2 _1779_ (
    .A(PC[0]),
    .Y(_931_)
);

INVX1 _1780_ (
    .A(DIMUX[0]),
    .Y(_932_)
);

NAND2X1 _1781_ (
    .A(_869__bF$buf0),
    .B(_900_),
    .Y(_933_)
);

NAND2X1 _1782_ (
    .A(_926__bF$buf2),
    .B(_928_),
    .Y(_934_)
);

NOR2X1 _1783_ (
    .A(_899_),
    .B(_874_),
    .Y(_935_)
);

INVX2 _1784_ (
    .A(_935_),
    .Y(_936_)
);

OAI21X1 _1785_ (
    .A(_918__bF$buf2),
    .B(_936_),
    .C(_934_),
    .Y(_937_)
);

NAND2X1 _1786_ (
    .A(_886__bF$buf3),
    .B(_900_),
    .Y(_938_)
);

OAI21X1 _1787_ (
    .A(_887__bF$buf2),
    .B(_936_),
    .C(_938_),
    .Y(_939_)
);

OR2X2 _1788_ (
    .A(_939_),
    .B(_937_),
    .Y(_940_)
);

INVX1 _1789_ (
    .A(_876_),
    .Y(_941_)
);

NOR2X1 _1790_ (
    .A(_887__bF$buf1),
    .B(_941_),
    .Y(_942_)
);

INVX1 _1791_ (
    .A(_933_),
    .Y(_943_)
);

NOR2X1 _1792_ (
    .A(_943_),
    .B(_942_),
    .Y(_944_)
);

NOR2X1 _1793_ (
    .A(state[2]),
    .B(_866_),
    .Y(_945_)
);

NAND2X1 _1794_ (
    .A(_915_),
    .B(_945_),
    .Y(_946_)
);

OAI21X1 _1795_ (
    .A(_918__bF$buf1),
    .B(_946_),
    .C(_944_),
    .Y(_947_)
);

NOR2X1 _1796_ (
    .A(_940_),
    .B(_947_),
    .Y(_948_)
);

NAND2X1 _1797_ (
    .A(_881_),
    .B(_893_),
    .Y(_949_)
);

INVX1 _1798_ (
    .A(_949_),
    .Y(_950_)
);

NOR2X1 _1799_ (
    .A(_887__bF$buf0),
    .B(_880_),
    .Y(_951_)
);

INVX1 _1800_ (
    .A(_951_),
    .Y(_952_)
);

AND2X2 _1801_ (
    .A(_914_),
    .B(_879_),
    .Y(_953_)
);

NAND2X1 _1802_ (
    .A(_926__bF$buf1),
    .B(_953_),
    .Y(_954_)
);

NOR2X1 _1803_ (
    .A(_892_),
    .B(_909_),
    .Y(_955_)
);

OAI21X1 _1804_ (
    .A(_953_),
    .B(_955_),
    .C(_869__bF$buf3),
    .Y(_956_)
);

NAND3X1 _1805_ (
    .A(_952_),
    .B(_954_),
    .C(_956_),
    .Y(_957_)
);

NOR2X1 _1806_ (
    .A(_950_),
    .B(_957_),
    .Y(_958_)
);

INVX1 _1807_ (
    .A(_898_),
    .Y(_959_)
);

INVX1 _1808_ (
    .A(_875_),
    .Y(_960_)
);

NAND2X1 _1809_ (
    .A(_960_),
    .B(_945_),
    .Y(_961_)
);

OAI21X1 _1810_ (
    .A(_882__bF$buf2),
    .B(_961_),
    .C(_907_),
    .Y(_962_)
);

OR2X2 _1811_ (
    .A(_962_),
    .B(_959_),
    .Y(_963_)
);

OAI21X1 _1812_ (
    .A(_893_),
    .B(_927_),
    .C(_886__bF$buf2),
    .Y(_964_)
);

OAI21X1 _1813_ (
    .A(state[4]),
    .B(_891_),
    .C(_964_),
    .Y(_965_)
);

NOR2X1 _1814_ (
    .A(_965_),
    .B(_963_),
    .Y(_966_)
);

NAND3X1 _1815_ (
    .A(_958_),
    .B(_966_),
    .C(_948_),
    .Y(_967_)
);

OAI22X1 _1816_ (
    .A(_931_),
    .B(_933_),
    .C(_932_),
    .D(_967_),
    .Y(BI[0])
);

INVX2 _1817_ (
    .A(PC[1]),
    .Y(_968_)
);

INVX2 _1818_ (
    .A(DIMUX[1]),
    .Y(_969_)
);

OAI22X1 _1819_ (
    .A(_968_),
    .B(_933_),
    .C(_969_),
    .D(_967_),
    .Y(BI[1])
);

INVX1 _1820_ (
    .A(PC[2]),
    .Y(_970_)
);

OAI22X1 _1821_ (
    .A(_970_),
    .B(_933_),
    .C(_855_),
    .D(_967_),
    .Y(BI[2])
);

INVX2 _1822_ (
    .A(PC[3]),
    .Y(_971_)
);

OAI22X1 _1823_ (
    .A(_971_),
    .B(_933_),
    .C(_857_),
    .D(_967_),
    .Y(BI[3])
);

INVX1 _1824_ (
    .A(PC[4]),
    .Y(_972_)
);

OAI22X1 _1825_ (
    .A(_972_),
    .B(_933_),
    .C(_859_),
    .D(_967_),
    .Y(BI[4])
);

INVX2 _1826_ (
    .A(PC[5]),
    .Y(_973_)
);

OAI22X1 _1827_ (
    .A(_973_),
    .B(_933_),
    .C(_861_),
    .D(_967_),
    .Y(BI[5])
);

INVX2 _1828_ (
    .A(PC[6]),
    .Y(_974_)
);

OAI22X1 _1829_ (
    .A(_974_),
    .B(_933_),
    .C(_863_),
    .D(_967_),
    .Y(BI[6])
);

INVX2 _1830_ (
    .A(PC[7]),
    .Y(_975_)
);

OAI22X1 _1831_ (
    .A(_975_),
    .B(_933_),
    .C(_864_),
    .D(_967_),
    .Y(BI[7])
);

OAI21X1 _1832_ (
    .A(_886__bF$buf1),
    .B(_926__bF$buf0),
    .C(_953_),
    .Y(_976_)
);

NAND2X1 _1833_ (
    .A(_926__bF$buf3),
    .B(_897_),
    .Y(_977_)
);

NAND2X1 _1834_ (
    .A(_869__bF$buf2),
    .B(_906_),
    .Y(_978_)
);

NAND3X1 _1835_ (
    .A(_976_),
    .B(_977_),
    .C(_978_),
    .Y(_979_)
);

INVX1 _1836_ (
    .A(_979_),
    .Y(_980_)
);

NAND2X1 _1837_ (
    .A(_926__bF$buf2),
    .B(_893_),
    .Y(_981_)
);

NAND3X1 _1838_ (
    .A(_934_),
    .B(_938_),
    .C(_981_),
    .Y(_982_)
);

INVX1 _1839_ (
    .A(_982_),
    .Y(_983_)
);

NAND2X1 _1840_ (
    .A(_917_),
    .B(_955_),
    .Y(_984_)
);

NAND2X1 _1841_ (
    .A(_984_),
    .B(_964_),
    .Y(_985_)
);

INVX1 _1842_ (
    .A(_985_),
    .Y(_986_)
);

NAND3X1 _1843_ (
    .A(_980_),
    .B(_983_),
    .C(_986_),
    .Y(_987_)
);

NAND2X1 _1844_ (
    .A(_879_),
    .B(_914_),
    .Y(_988_)
);

NAND2X1 _1845_ (
    .A(_914_),
    .B(_871_),
    .Y(_989_)
);

NAND2X1 _1846_ (
    .A(_926__bF$buf1),
    .B(_876_),
    .Y(_990_)
);

OAI21X1 _1847_ (
    .A(_918__bF$buf0),
    .B(_989_),
    .C(_990_),
    .Y(_991_)
);

NAND2X1 _1848_ (
    .A(_869__bF$buf1),
    .B(_927_),
    .Y(_992_)
);

NOR2X1 _1849_ (
    .A(_881_),
    .B(_917_),
    .Y(_993_)
);

INVX1 _1850_ (
    .A(_993_),
    .Y(_994_)
);

NOR2X1 _1851_ (
    .A(state[2]),
    .B(state[3]),
    .Y(_995_)
);

NAND2X1 _1852_ (
    .A(_995_),
    .B(_879_),
    .Y(_996_)
);

OAI21X1 _1853_ (
    .A(_994_),
    .B(_996_),
    .C(_992_),
    .Y(_997_)
);

NOR2X1 _1854_ (
    .A(_991_),
    .B(_997_),
    .Y(_998_)
);

OAI21X1 _1855_ (
    .A(_918__bF$buf3),
    .B(_988_),
    .C(_998_),
    .Y(_999_)
);

NOR2X1 _1856_ (
    .A(_987_),
    .B(_999_),
    .Y(_1000_)
);

INVX1 _1857_ (
    .A(dst_reg[1]),
    .Y(_1001_)
);

NAND3X1 _1858_ (
    .A(_879_),
    .B(_914_),
    .C(_869__bF$buf0),
    .Y(_1002_)
);

OAI21X1 _1859_ (
    .A(_1001_),
    .B(_1002__bF$buf4),
    .C(_998_),
    .Y(_1003_)
);

AOI21X1 _1860_ (
    .A(_1000_),
    .B(src_reg[1]),
    .C(_1003_),
    .Y(_1004_)
);

NOR3X1 _1861_ (
    .A(_979_),
    .B(_982_),
    .C(_985_),
    .Y(_1005_)
);

NAND3X1 _1862_ (
    .A(_1002__bF$buf3),
    .B(_998_),
    .C(_1005_),
    .Y(_1006_)
);

OAI21X1 _1863_ (
    .A(_991_),
    .B(_997_),
    .C(index_y),
    .Y(_1007_)
);

INVX2 _1864_ (
    .A(_1002__bF$buf2),
    .Y(_1008_)
);

NAND2X1 _1865_ (
    .A(dst_reg[0]),
    .B(_1008_),
    .Y(_1009_)
);

NAND3X1 _1866_ (
    .A(_1007_),
    .B(_1009_),
    .C(_1005_),
    .Y(_1010_)
);

MUX2X1 _1867_ (
    .A(_1010_),
    .B(src_reg[0]),
    .S(_1006_),
    .Y(_1011_)
);

NOR2X1 _1868_ (
    .A(_1004_),
    .B(_1011_),
    .Y(_1012_)
);

NAND2X1 _1869_ (
    .A(\AXYS[3] [0]),
    .B(_1012_),
    .Y(_1013_)
);

INVX1 _1870_ (
    .A(src_reg[1]),
    .Y(_1014_)
);

INVX1 _1871_ (
    .A(_1003_),
    .Y(_1015_)
);

OAI21X1 _1872_ (
    .A(_1014_),
    .B(_1006_),
    .C(_1015_),
    .Y(_1016_)
);

AND2X2 _1873_ (
    .A(_1005_),
    .B(_1009_),
    .Y(_1017_)
);

NAND3X1 _1874_ (
    .A(_1006_),
    .B(_1007_),
    .C(_1017_),
    .Y(_1018_)
);

OR2X2 _1875_ (
    .A(_1006_),
    .B(src_reg[0]),
    .Y(_1019_)
);

AOI21X1 _1876_ (
    .A(_1019_),
    .B(_1018_),
    .C(_1016_),
    .Y(_1020_)
);

NAND2X1 _1877_ (
    .A(\AXYS[0] [0]),
    .B(_1020_),
    .Y(_1021_)
);

NOR2X1 _1878_ (
    .A(_1016_),
    .B(_1011_),
    .Y(_1022_)
);

AOI21X1 _1879_ (
    .A(_1018_),
    .B(_1019_),
    .C(_1004_),
    .Y(_1023_)
);

AOI22X1 _1880_ (
    .A(\AXYS[2] [0]),
    .B(_1023_),
    .C(_1022_),
    .D(\AXYS[1] [0]),
    .Y(_1024_)
);

NAND3X1 _1881_ (
    .A(_1013_),
    .B(_1021_),
    .C(_1024_),
    .Y(_1025_)
);

INVX1 _1882_ (
    .A(_1025_),
    .Y(_1026_)
);

INVX1 _1883_ (
    .A(_991_),
    .Y(_1027_)
);

OAI21X1 _1884_ (
    .A(_887__bF$buf4),
    .B(_901_),
    .C(_1027_),
    .Y(_1028_)
);

INVX1 _1885_ (
    .A(_954_),
    .Y(_1029_)
);

NOR2X1 _1886_ (
    .A(_1029_),
    .B(_951_),
    .Y(_1030_)
);

INVX1 _1887_ (
    .A(_919_),
    .Y(_1031_)
);

NAND2X1 _1888_ (
    .A(_995_),
    .B(_871_),
    .Y(_1032_)
);

OAI22X1 _1889_ (
    .A(state[4]),
    .B(_1032_),
    .C(load_only),
    .D(_1031_),
    .Y(_1033_)
);

OAI21X1 _1890_ (
    .A(_886__bF$buf0),
    .B(_926__bF$buf0),
    .C(_893_),
    .Y(_1034_)
);

NAND2X1 _1891_ (
    .A(_879_),
    .B(_945_),
    .Y(_1035_)
);

NOR2X1 _1892_ (
    .A(_918__bF$buf2),
    .B(_1035_),
    .Y(_1036_)
);

INVX2 _1893_ (
    .A(_996_),
    .Y(_1037_)
);

NAND2X1 _1894_ (
    .A(_993_),
    .B(_1037_),
    .Y(_1038_)
);

INVX1 _1895_ (
    .A(_1038_),
    .Y(_1039_)
);

NOR2X1 _1896_ (
    .A(_1036_),
    .B(_1039_),
    .Y(_1040_)
);

NAND2X1 _1897_ (
    .A(_1034_),
    .B(_1040_),
    .Y(_1041_)
);

NOR2X1 _1898_ (
    .A(_1033_),
    .B(_1041_),
    .Y(_1042_)
);

INVX1 _1899_ (
    .A(_934_),
    .Y(_1043_)
);

NOR2X1 _1900_ (
    .A(_887__bF$buf3),
    .B(_936_),
    .Y(_1044_)
);

NOR2X1 _1901_ (
    .A(_1043_),
    .B(_1044_),
    .Y(_1045_)
);

NAND3X1 _1902_ (
    .A(_1030_),
    .B(_1045_),
    .C(_1042_),
    .Y(_1046_)
);

NOR2X1 _1903_ (
    .A(_1028_),
    .B(_1046_),
    .Y(_1047_)
);

NOR2X1 _1904_ (
    .A(_918__bF$buf1),
    .B(_946_),
    .Y(_1048_)
);

INVX1 _1905_ (
    .A(_1048_),
    .Y(_1049_)
);

INVX1 _1906_ (
    .A(_963_),
    .Y(_1050_)
);

NAND2X1 _1907_ (
    .A(_869__bF$buf3),
    .B(_893_),
    .Y(_1051_)
);

OAI21X1 _1908_ (
    .A(_887__bF$buf2),
    .B(_891_),
    .C(_1051__bF$buf3),
    .Y(_1052_)
);

INVX1 _1909_ (
    .A(_1052_),
    .Y(_1053_)
);

NAND3X1 _1910_ (
    .A(_1049_),
    .B(_1053_),
    .C(_1050_),
    .Y(_1054_)
);

INVX1 _1911_ (
    .A(ABH[0]),
    .Y(_1055_)
);

NOR2X1 _1912_ (
    .A(_1055_),
    .B(_872_),
    .Y(_1056_)
);

INVX1 _1913_ (
    .A(_1056_),
    .Y(_1057_)
);

OAI21X1 _1914_ (
    .A(_932_),
    .B(_944_),
    .C(_1057_),
    .Y(_1058_)
);

AOI21X1 _1915_ (
    .A(_1054_),
    .B(ADD[0]),
    .C(_1058_),
    .Y(_1059_)
);

OAI21X1 _1916_ (
    .A(_1047_),
    .B(_1026_),
    .C(_1059_),
    .Y(AI[0])
);

NAND2X1 _1917_ (
    .A(\AXYS[1] [1]),
    .B(_1022_),
    .Y(_1060_)
);

AOI22X1 _1918_ (
    .A(\AXYS[2] [1]),
    .B(_1023_),
    .C(_1012_),
    .D(\AXYS[3] [1]),
    .Y(_1061_)
);

NAND2X1 _1919_ (
    .A(\AXYS[0] [1]),
    .B(_1020_),
    .Y(_1062_)
);

NAND3X1 _1920_ (
    .A(_1060_),
    .B(_1062_),
    .C(_1061_),
    .Y(_1063_)
);

INVX1 _1921_ (
    .A(_1063_),
    .Y(_1064_)
);

INVX1 _1922_ (
    .A(ABH[1]),
    .Y(_1065_)
);

NOR2X1 _1923_ (
    .A(_1065_),
    .B(_872_),
    .Y(_1066_)
);

INVX1 _1924_ (
    .A(_1066_),
    .Y(_1067_)
);

OAI21X1 _1925_ (
    .A(_969_),
    .B(_944_),
    .C(_1067_),
    .Y(_1068_)
);

AOI21X1 _1926_ (
    .A(_1054_),
    .B(ADD[1]),
    .C(_1068_),
    .Y(_1069_)
);

OAI21X1 _1927_ (
    .A(_1047_),
    .B(_1064_),
    .C(_1069_),
    .Y(AI[1])
);

NAND2X1 _1928_ (
    .A(\AXYS[1] [2]),
    .B(_1022_),
    .Y(_1070_)
);

AOI22X1 _1929_ (
    .A(\AXYS[2] [2]),
    .B(_1023_),
    .C(_1012_),
    .D(\AXYS[3] [2]),
    .Y(_1071_)
);

NAND2X1 _1930_ (
    .A(\AXYS[0] [2]),
    .B(_1020_),
    .Y(_1072_)
);

NAND3X1 _1931_ (
    .A(_1070_),
    .B(_1072_),
    .C(_1071_),
    .Y(_1073_)
);

INVX1 _1932_ (
    .A(_1073_),
    .Y(_1074_)
);

NOR3X1 _1933_ (
    .A(_867_),
    .B(_918__bF$buf0),
    .C(_889_),
    .Y(_1075_)
);

NAND2X1 _1934_ (
    .A(ABH[2]),
    .B(_1075_),
    .Y(_1076_)
);

OAI21X1 _1935_ (
    .A(_855_),
    .B(_944_),
    .C(_1076_),
    .Y(_1077_)
);

AOI21X1 _1936_ (
    .A(_1054_),
    .B(ADD[2]),
    .C(_1077_),
    .Y(_1078_)
);

OAI21X1 _1937_ (
    .A(_1047_),
    .B(_1074_),
    .C(_1078_),
    .Y(AI[2])
);

NAND2X1 _1938_ (
    .A(\AXYS[1] [3]),
    .B(_1022_),
    .Y(_1079_)
);

AOI22X1 _1939_ (
    .A(\AXYS[2] [3]),
    .B(_1023_),
    .C(_1012_),
    .D(\AXYS[3] [3]),
    .Y(_1080_)
);

NAND2X1 _1940_ (
    .A(\AXYS[0] [3]),
    .B(_1020_),
    .Y(_1081_)
);

NAND3X1 _1941_ (
    .A(_1079_),
    .B(_1081_),
    .C(_1080_),
    .Y(_1082_)
);

INVX1 _1942_ (
    .A(_1082_),
    .Y(_1083_)
);

NAND2X1 _1943_ (
    .A(ABH[3]),
    .B(_1075_),
    .Y(_1084_)
);

OAI21X1 _1944_ (
    .A(_857_),
    .B(_944_),
    .C(_1084_),
    .Y(_1085_)
);

AOI21X1 _1945_ (
    .A(_1054_),
    .B(ADD[3]),
    .C(_1085_),
    .Y(_1086_)
);

OAI21X1 _1946_ (
    .A(_1047_),
    .B(_1083_),
    .C(_1086_),
    .Y(AI[3])
);

NAND2X1 _1947_ (
    .A(\AXYS[1] [4]),
    .B(_1022_),
    .Y(_1087_)
);

AOI22X1 _1948_ (
    .A(\AXYS[2] [4]),
    .B(_1023_),
    .C(_1012_),
    .D(\AXYS[3] [4]),
    .Y(_1088_)
);

NAND2X1 _1949_ (
    .A(\AXYS[0] [4]),
    .B(_1020_),
    .Y(_1089_)
);

NAND3X1 _1950_ (
    .A(_1087_),
    .B(_1089_),
    .C(_1088_),
    .Y(_1090_)
);

INVX1 _1951_ (
    .A(_1090_),
    .Y(_1091_)
);

NAND2X1 _1952_ (
    .A(ABH[4]),
    .B(_1075_),
    .Y(_1092_)
);

OAI21X1 _1953_ (
    .A(_859_),
    .B(_944_),
    .C(_1092_),
    .Y(_1093_)
);

AOI21X1 _1954_ (
    .A(_1054_),
    .B(ADD[4]),
    .C(_1093_),
    .Y(_1094_)
);

OAI21X1 _1955_ (
    .A(_1047_),
    .B(_1091_),
    .C(_1094_),
    .Y(AI[4])
);

NAND2X1 _1956_ (
    .A(\AXYS[1] [5]),
    .B(_1022_),
    .Y(_1095_)
);

AOI22X1 _1957_ (
    .A(\AXYS[2] [5]),
    .B(_1023_),
    .C(_1012_),
    .D(\AXYS[3] [5]),
    .Y(_1096_)
);

NAND2X1 _1958_ (
    .A(\AXYS[0] [5]),
    .B(_1020_),
    .Y(_1097_)
);

NAND3X1 _1959_ (
    .A(_1095_),
    .B(_1097_),
    .C(_1096_),
    .Y(_1098_)
);

INVX1 _1960_ (
    .A(_1098_),
    .Y(_1099_)
);

NAND2X1 _1961_ (
    .A(ABH[5]),
    .B(_1075_),
    .Y(_1100_)
);

OAI21X1 _1962_ (
    .A(_861_),
    .B(_944_),
    .C(_1100_),
    .Y(_1101_)
);

AOI21X1 _1963_ (
    .A(_1054_),
    .B(ADD[5]),
    .C(_1101_),
    .Y(_1102_)
);

OAI21X1 _1964_ (
    .A(_1047_),
    .B(_1099_),
    .C(_1102_),
    .Y(AI[5])
);

NAND2X1 _1965_ (
    .A(\AXYS[1] [6]),
    .B(_1022_),
    .Y(_1103_)
);

AOI22X1 _1966_ (
    .A(\AXYS[2] [6]),
    .B(_1023_),
    .C(_1012_),
    .D(\AXYS[3] [6]),
    .Y(_1104_)
);

NAND2X1 _1967_ (
    .A(\AXYS[0] [6]),
    .B(_1020_),
    .Y(_1105_)
);

NAND3X1 _1968_ (
    .A(_1103_),
    .B(_1105_),
    .C(_1104_),
    .Y(_1106_)
);

INVX1 _1969_ (
    .A(_1106_),
    .Y(_1107_)
);

INVX1 _1970_ (
    .A(ABH[6]),
    .Y(_1108_)
);

NOR2X1 _1971_ (
    .A(_1108_),
    .B(_872_),
    .Y(_1109_)
);

INVX1 _1972_ (
    .A(_1109_),
    .Y(_1110_)
);

OAI21X1 _1973_ (
    .A(_863_),
    .B(_944_),
    .C(_1110_),
    .Y(_1111_)
);

AOI21X1 _1974_ (
    .A(_1054_),
    .B(ADD[6]),
    .C(_1111_),
    .Y(_1112_)
);

OAI21X1 _1975_ (
    .A(_1047_),
    .B(_1107_),
    .C(_1112_),
    .Y(AI[6])
);

NAND2X1 _1976_ (
    .A(\AXYS[1] [7]),
    .B(_1022_),
    .Y(_1113_)
);

AOI22X1 _1977_ (
    .A(\AXYS[2] [7]),
    .B(_1023_),
    .C(_1012_),
    .D(\AXYS[3] [7]),
    .Y(_1114_)
);

NAND2X1 _1978_ (
    .A(\AXYS[0] [7]),
    .B(_1020_),
    .Y(_1115_)
);

NAND3X1 _1979_ (
    .A(_1113_),
    .B(_1115_),
    .C(_1114_),
    .Y(_1116_)
);

INVX1 _1980_ (
    .A(_1116_),
    .Y(_1117_)
);

INVX1 _1981_ (
    .A(ABH[7]),
    .Y(_1118_)
);

NOR2X1 _1982_ (
    .A(_1118_),
    .B(_872_),
    .Y(_1119_)
);

INVX1 _1983_ (
    .A(_1119_),
    .Y(_1120_)
);

OAI21X1 _1984_ (
    .A(_864_),
    .B(_944_),
    .C(_1120_),
    .Y(_1121_)
);

AOI21X1 _1985_ (
    .A(_1054_),
    .B(AN),
    .C(_1121_),
    .Y(_1122_)
);

OAI21X1 _1986_ (
    .A(_1047_),
    .B(_1117_),
    .C(_1122_),
    .Y(AI[7])
);

NAND2X1 _1987_ (
    .A(_926__bF$buf3),
    .B(_900_),
    .Y(_1123_)
);

INVX1 _1988_ (
    .A(_1123_),
    .Y(_1124_)
);

OR2X2 _1989_ (
    .A(CO),
    .B(store),
    .Y(_1125_)
);

AND2X2 _1990_ (
    .A(_883_),
    .B(RDY_bF$buf6),
    .Y(_1126_)
);

AOI22X1 _1991_ (
    .A(_853__bF$buf2),
    .B(_1124_),
    .C(_1126_),
    .D(_1125_),
    .Y(_1127_)
);

OR2X2 _1992_ (
    .A(_938_),
    .B(RDY_bF$buf5),
    .Y(_1128_)
);

NOR2X1 _1993_ (
    .A(_853__bF$buf1),
    .B(_1002__bF$buf1),
    .Y(_1129_)
);

INVX1 _1994_ (
    .A(IRHOLD[1]),
    .Y(_1130_)
);

INVX1 _1995_ (
    .A(IRQ),
    .Y(_1131_)
);

INVX1 _1996_ (
    .A(NMI_edge),
    .Y(_1132_)
);

OAI21X1 _1997_ (
    .A(I),
    .B(_1131_),
    .C(_1132_),
    .Y(_1133_)
);

AOI21X1 _1998_ (
    .A(IRHOLD_valid_bF$buf3),
    .B(_1130_),
    .C(_1133_),
    .Y(_1134_)
);

OAI21X1 _1999_ (
    .A(IRHOLD_valid_bF$buf2),
    .B(DIMUX[1]),
    .C(_1134_),
    .Y(_1135_)
);

INVX1 _2000_ (
    .A(IRHOLD[0]),
    .Y(_1136_)
);

AOI21X1 _2001_ (
    .A(_1136_),
    .B(IRHOLD_valid_bF$buf1),
    .C(_1133_),
    .Y(_1137_)
);

OAI21X1 _2002_ (
    .A(IRHOLD_valid_bF$buf0),
    .B(DIMUX[0]),
    .C(_1137_),
    .Y(_1138_)
);

NAND2X1 _2003_ (
    .A(_1135_),
    .B(_1138_),
    .Y(_1139_)
);

INVX1 _2004_ (
    .A(IRHOLD[3]),
    .Y(_1140_)
);

AOI21X1 _2005_ (
    .A(IRHOLD_valid_bF$buf3),
    .B(_1140_),
    .C(_1133_),
    .Y(_1141_)
);

OAI21X1 _2006_ (
    .A(IRHOLD_valid_bF$buf2),
    .B(DIMUX[3]),
    .C(_1141_),
    .Y(_1142_)
);

INVX1 _2007_ (
    .A(I),
    .Y(_1143_)
);

NAND2X1 _2008_ (
    .A(_1131_),
    .B(_1132_),
    .Y(_1144_)
);

OAI21X1 _2009_ (
    .A(_1143_),
    .B(NMI_edge),
    .C(_1144_),
    .Y(_1145_)
);

NAND2X1 _2010_ (
    .A(IRHOLD_valid_bF$buf1),
    .B(IRHOLD[2]),
    .Y(_1146_)
);

OAI21X1 _2011_ (
    .A(IRHOLD_valid_bF$buf0),
    .B(_855_),
    .C(_1146_),
    .Y(_1147_)
);

NAND2X1 _2012_ (
    .A(_1145_),
    .B(_1147_),
    .Y(_1148_)
);

NAND2X1 _2013_ (
    .A(_1142_),
    .B(_1148_),
    .Y(_1149_)
);

NOR2X1 _2014_ (
    .A(_1139_),
    .B(_1149_),
    .Y(_1150_)
);

NAND2X1 _2015_ (
    .A(IRHOLD_valid_bF$buf3),
    .B(IRHOLD[4]),
    .Y(_1151_)
);

OAI21X1 _2016_ (
    .A(IRHOLD_valid_bF$buf2),
    .B(_859_),
    .C(_1151_),
    .Y(_1152_)
);

NAND2X1 _2017_ (
    .A(IRHOLD_valid_bF$buf1),
    .B(IRHOLD[5]),
    .Y(_1153_)
);

OAI21X1 _2018_ (
    .A(IRHOLD_valid_bF$buf0),
    .B(_861_),
    .C(_1153_),
    .Y(_1154_)
);

OAI21X1 _2019_ (
    .A(_1152_),
    .B(_1154_),
    .C(_1145_),
    .Y(_1155_)
);

INVX1 _2020_ (
    .A(_1155_),
    .Y(_1156_)
);

NAND2X1 _2021_ (
    .A(IRHOLD_valid_bF$buf3),
    .B(IRHOLD[7]),
    .Y(_1157_)
);

OAI21X1 _2022_ (
    .A(IRHOLD_valid_bF$buf2),
    .B(_864_),
    .C(_1157_),
    .Y(_1158_)
);

NAND2X1 _2023_ (
    .A(_1145_),
    .B(_1158_),
    .Y(_1159_)
);

NAND2X1 _2024_ (
    .A(IRHOLD_valid_bF$buf1),
    .B(IRHOLD[6]),
    .Y(_1160_)
);

OAI21X1 _2025_ (
    .A(IRHOLD_valid_bF$buf0),
    .B(_863_),
    .C(_1160_),
    .Y(_1161_)
);

AND2X2 _2026_ (
    .A(_1161_),
    .B(_1145_),
    .Y(_1162_)
);

NAND2X1 _2027_ (
    .A(_1159_),
    .B(_1162_),
    .Y(_1163_)
);

NOR2X1 _2028_ (
    .A(_1156_),
    .B(_1163_),
    .Y(_1164_)
);

NAND3X1 _2029_ (
    .A(_1129__bF$buf4),
    .B(_1150_),
    .C(_1164_),
    .Y(_1165_)
);

NAND3X1 _2030_ (
    .A(_1127_),
    .B(_1128_),
    .C(_1165_),
    .Y(_1166_)
);

INVX1 _2031_ (
    .A(_1166_),
    .Y(_1167_)
);

NAND2X1 _2032_ (
    .A(_1145_),
    .B(_1152_),
    .Y(_1168_)
);

INVX1 _2033_ (
    .A(IRHOLD_valid_bF$buf3),
    .Y(_1169_)
);

OAI21X1 _2034_ (
    .A(_1169_),
    .B(IRHOLD[3]),
    .C(_1145_),
    .Y(_1170_)
);

AOI21X1 _2035_ (
    .A(_1169_),
    .B(_857_),
    .C(_1170_),
    .Y(_1171_)
);

NAND2X1 _2036_ (
    .A(_1148_),
    .B(_1171_),
    .Y(_1172_)
);

INVX1 _2037_ (
    .A(_1172_),
    .Y(_1173_)
);

INVX1 _2038_ (
    .A(_1135_),
    .Y(_1174_)
);

NOR2X1 _2039_ (
    .A(_1138_),
    .B(_1174_),
    .Y(_1175_)
);

NAND2X1 _2040_ (
    .A(_1175_),
    .B(_1173_),
    .Y(_1176_)
);

NAND2X1 _2041_ (
    .A(_1138_),
    .B(_1148_),
    .Y(_1177_)
);

INVX1 _2042_ (
    .A(_1159_),
    .Y(_1178_)
);

NAND2X1 _2043_ (
    .A(_1142_),
    .B(_1178_),
    .Y(_1179_)
);

OAI21X1 _2044_ (
    .A(_1177_),
    .B(_1179_),
    .C(_1176_),
    .Y(_1180_)
);

NAND3X1 _2045_ (
    .A(_1129__bF$buf3),
    .B(_1168_),
    .C(_1180_),
    .Y(_1181_)
);

NOR2X1 _2046_ (
    .A(_917_),
    .B(_936_),
    .Y(_1182_)
);

INVX1 _2047_ (
    .A(_1182_),
    .Y(_1183_)
);

NAND2X1 _2048_ (
    .A(_886__bF$buf3),
    .B(_897_),
    .Y(_1184_)
);

INVX1 _2049_ (
    .A(_1184_),
    .Y(_1185_)
);

NAND2X1 _2050_ (
    .A(_869__bF$buf2),
    .B(_910_),
    .Y(_1186_)
);

OAI21X1 _2051_ (
    .A(_918__bF$buf3),
    .B(_936_),
    .C(_1186_),
    .Y(_1187_)
);

NOR2X1 _2052_ (
    .A(_1185_),
    .B(_1187_),
    .Y(_1188_)
);

OAI21X1 _2053_ (
    .A(_881_),
    .B(_1183_),
    .C(_1188_),
    .Y(_1189_)
);

INVX1 _2054_ (
    .A(_1189_),
    .Y(_1190_)
);

NOR2X1 _2055_ (
    .A(_887__bF$buf1),
    .B(_989_),
    .Y(_1191_)
);

INVX1 _2056_ (
    .A(_1191_),
    .Y(_1192_)
);

NOR2X1 _2057_ (
    .A(_896_),
    .B(_899_),
    .Y(_1193_)
);

OAI21X1 _2058_ (
    .A(_886__bF$buf2),
    .B(_926__bF$buf2),
    .C(_1193_),
    .Y(_1194_)
);

OAI21X1 _2059_ (
    .A(_900_),
    .B(_935_),
    .C(_926__bF$buf1),
    .Y(_1195_)
);

NAND3X1 _2060_ (
    .A(_1194_),
    .B(_1195_),
    .C(_1192_),
    .Y(_1196_)
);

NAND3X1 _2061_ (
    .A(RDY_bF$buf4),
    .B(_1196_),
    .C(_1190_),
    .Y(_1197_)
);

NOR2X1 _2062_ (
    .A(write_back),
    .B(_853__bF$buf0),
    .Y(_1198_)
);

NAND2X1 _2063_ (
    .A(RDY_bF$buf3),
    .B(_883_),
    .Y(_1199_)
);

NOR2X1 _2064_ (
    .A(write_back),
    .B(_1125_),
    .Y(_1200_)
);

NAND3X1 _2065_ (
    .A(RDY_bF$buf2),
    .B(_1200_),
    .C(_878_),
    .Y(_1201_)
);

OAI21X1 _2066_ (
    .A(_1125_),
    .B(_1199_),
    .C(_1201_),
    .Y(_1202_)
);

OAI21X1 _2067_ (
    .A(_882__bF$buf1),
    .B(_916_),
    .C(_853__bF$buf7),
    .Y(_1203_)
);

OAI21X1 _2068_ (
    .A(_853__bF$buf6),
    .B(_1029_),
    .C(_1203_),
    .Y(_1204_)
);

OAI21X1 _2069_ (
    .A(_988_),
    .B(_887__bF$buf0),
    .C(RDY_bF$buf1),
    .Y(_1205_)
);

OAI21X1 _2070_ (
    .A(_887__bF$buf4),
    .B(_916_),
    .C(_853__bF$buf5),
    .Y(_1206_)
);

NAND2X1 _2071_ (
    .A(_1205_),
    .B(_1206_),
    .Y(_1207_)
);

NAND2X1 _2072_ (
    .A(_853__bF$buf4),
    .B(_919_),
    .Y(_1208_)
);

NAND3X1 _2073_ (
    .A(_1208_),
    .B(_1207_),
    .C(_1204_),
    .Y(_1209_)
);

OR2X2 _2074_ (
    .A(_1202_),
    .B(_1209_),
    .Y(_1210_)
);

AOI21X1 _2075_ (
    .A(_1189_),
    .B(_1198_),
    .C(_1210_),
    .Y(_1211_)
);

AND2X2 _2076_ (
    .A(_1211_),
    .B(_1197_),
    .Y(_1212_)
);

NAND3X1 _2077_ (
    .A(_1167_),
    .B(_1181_),
    .C(_1212_),
    .Y(_1213_)
);

INVX1 _2078_ (
    .A(_1139_),
    .Y(_1214_)
);

NAND2X1 _2079_ (
    .A(_1214_),
    .B(_1173_),
    .Y(_1215_)
);

NAND2X1 _2080_ (
    .A(_1159_),
    .B(_1155_),
    .Y(_1216_)
);

NOR2X1 _2081_ (
    .A(_1216_),
    .B(_1215_),
    .Y(_1217_)
);

AOI22X1 _2082_ (
    .A(_853__bF$buf3),
    .B(_1044_),
    .C(_1217_),
    .D(_1129__bF$buf2),
    .Y(_1218_)
);

INVX8 _2083_ (
    .A(_1129__bF$buf1),
    .Y(_1219_)
);

INVX2 _2084_ (
    .A(_1168_),
    .Y(_1220_)
);

NAND2X1 _2085_ (
    .A(_1220_),
    .B(_1150_),
    .Y(_1221_)
);

NOR2X1 _2086_ (
    .A(_1219__bF$buf3),
    .B(_1221_),
    .Y(_1222_)
);

AOI21X1 _2087_ (
    .A(_853__bF$buf2),
    .B(_943_),
    .C(_1222_),
    .Y(_1223_)
);

NOR2X1 _2088_ (
    .A(_882__bF$buf0),
    .B(_1035_),
    .Y(_1224_)
);

OAI21X1 _2089_ (
    .A(_882__bF$buf3),
    .B(_946_),
    .C(_853__bF$buf1),
    .Y(_1225_)
);

OAI21X1 _2090_ (
    .A(_853__bF$buf0),
    .B(_1224_),
    .C(_1225_),
    .Y(_1226_)
);

NAND2X1 _2091_ (
    .A(_886__bF$buf1),
    .B(_955_),
    .Y(_1227_)
);

NOR2X1 _2092_ (
    .A(_887__bF$buf3),
    .B(_946_),
    .Y(_1228_)
);

NAND2X1 _2093_ (
    .A(_853__bF$buf7),
    .B(_1228_),
    .Y(_1229_)
);

OAI21X1 _2094_ (
    .A(_853__bF$buf6),
    .B(_1227_),
    .C(_1229_),
    .Y(_1230_)
);

NAND2X1 _2095_ (
    .A(RDY_bF$buf0),
    .B(_1036_),
    .Y(_1231_)
);

OAI21X1 _2096_ (
    .A(RDY_bF$buf8),
    .B(_1049_),
    .C(_1231_),
    .Y(_1232_)
);

NOR2X1 _2097_ (
    .A(_1230_),
    .B(_1232_),
    .Y(_1233_)
);

AND2X2 _2098_ (
    .A(_1233_),
    .B(_1226_),
    .Y(_1234_)
);

NAND2X1 _2099_ (
    .A(_993_),
    .B(_935_),
    .Y(_1235_)
);

NAND2X1 _2100_ (
    .A(RDY_bF$buf7),
    .B(_1039_),
    .Y(_1236_)
);

OAI21X1 _2101_ (
    .A(RDY_bF$buf6),
    .B(_1235_),
    .C(_1236_),
    .Y(_1237_)
);

NAND2X1 _2102_ (
    .A(_926__bF$buf0),
    .B(_935_),
    .Y(_1238_)
);

NAND2X1 _2103_ (
    .A(_926__bF$buf3),
    .B(_1037_),
    .Y(_1239_)
);

INVX1 _2104_ (
    .A(_1239_),
    .Y(_1240_)
);

NAND2X1 _2105_ (
    .A(RDY_bF$buf5),
    .B(_1240_),
    .Y(_1241_)
);

OAI21X1 _2106_ (
    .A(RDY_bF$buf4),
    .B(_1238_),
    .C(_1241_),
    .Y(_1242_)
);

NOR2X1 _2107_ (
    .A(_1237_),
    .B(_1242_),
    .Y(_1243_)
);

NOR2X1 _2108_ (
    .A(_918__bF$buf2),
    .B(_936_),
    .Y(_1244_)
);

OAI21X1 _2109_ (
    .A(_918__bF$buf1),
    .B(_996_),
    .C(RDY_bF$buf3),
    .Y(_1245_)
);

OAI21X1 _2110_ (
    .A(RDY_bF$buf2),
    .B(_1244_),
    .C(_1245_),
    .Y(_1246_)
);

AND2X2 _2111_ (
    .A(_1243_),
    .B(_1246_),
    .Y(_1247_)
);

AND2X2 _2112_ (
    .A(_1247_),
    .B(_1234_),
    .Y(_1248_)
);

NAND3X1 _2113_ (
    .A(_1218_),
    .B(_1223_),
    .C(_1248_),
    .Y(_1249_)
);

INVX1 _2114_ (
    .A(write_back),
    .Y(_1250_)
);

OAI21X1 _2115_ (
    .A(_1250_),
    .B(_1190_),
    .C(RDY_bF$buf1),
    .Y(_1251_)
);

OAI21X1 _2116_ (
    .A(RDY_bF$buf0),
    .B(_942_),
    .C(_1251_),
    .Y(_1252_)
);

NOR2X1 _2117_ (
    .A(_1148_),
    .B(_1171_),
    .Y(_1253_)
);

NOR2X1 _2118_ (
    .A(_1219__bF$buf2),
    .B(_1220_),
    .Y(_1254_)
);

AOI22X1 _2119_ (
    .A(_853__bF$buf5),
    .B(_1185_),
    .C(_1254_),
    .D(_1253_),
    .Y(_1255_)
);

OAI21X1 _2120_ (
    .A(_918__bF$buf0),
    .B(_989_),
    .C(RDY_bF$buf8),
    .Y(_1256_)
);

OAI21X1 _2121_ (
    .A(RDY_bF$buf7),
    .B(_959_),
    .C(_1256_),
    .Y(_1257_)
);

NAND2X1 _2122_ (
    .A(_1257_),
    .B(_1255_),
    .Y(_1258_)
);

NAND2X1 _2123_ (
    .A(_960_),
    .B(_868_),
    .Y(_1259_)
);

NOR2X1 _2124_ (
    .A(_887__bF$buf2),
    .B(_1259_),
    .Y(_1260_)
);

OAI21X1 _2125_ (
    .A(_887__bF$buf1),
    .B(_891_),
    .C(RDY_bF$buf6),
    .Y(_1261_)
);

OAI21X1 _2126_ (
    .A(RDY_bF$buf5),
    .B(_1260_),
    .C(_1261_),
    .Y(_1262_)
);

OAI21X1 _2127_ (
    .A(_882__bF$buf2),
    .B(_891_),
    .C(RDY_bF$buf4),
    .Y(_1263_)
);

NOR3X1 _2128_ (
    .A(_875_),
    .B(_867_),
    .C(_882__bF$buf1),
    .Y(_1264_)
);

OAI21X1 _2129_ (
    .A(RDY_bF$buf3),
    .B(_1264_),
    .C(_1263_),
    .Y(_1265_)
);

NAND2X1 _2130_ (
    .A(_1265_),
    .B(_1262_),
    .Y(_1266_)
);

NAND2X1 _2131_ (
    .A(_869__bF$buf1),
    .B(_905_),
    .Y(_1267_)
);

XOR2X1 _2132_ (
    .A(CO),
    .B(backwards),
    .Y(_1268_)
);

NAND2X1 _2133_ (
    .A(RDY_bF$buf2),
    .B(_1268_),
    .Y(_1269_)
);

OAI22X1 _2134_ (
    .A(_872_),
    .B(_1269_),
    .C(RDY_bF$buf1),
    .D(_1267_),
    .Y(_1270_)
);

NOR3X1 _2135_ (
    .A(_1266_),
    .B(_1270_),
    .C(_1258_),
    .Y(_1271_)
);

OAI21X1 _2136_ (
    .A(_918__bF$buf3),
    .B(_1032_),
    .C(RDY_bF$buf0),
    .Y(_1272_)
);

OAI21X1 _2137_ (
    .A(RDY_bF$buf8),
    .B(_878_),
    .C(_1272_),
    .Y(_1273_)
);

INVX1 _2138_ (
    .A(_977_),
    .Y(_1274_)
);

OAI21X1 _2139_ (
    .A(_882__bF$buf0),
    .B(_989_),
    .C(RDY_bF$buf7),
    .Y(_1275_)
);

OAI21X1 _2140_ (
    .A(RDY_bF$buf6),
    .B(_1274_),
    .C(_1275_),
    .Y(_1276_)
);

INVX1 _2141_ (
    .A(_990_),
    .Y(_1277_)
);

OAI21X1 _2142_ (
    .A(_882__bF$buf3),
    .B(_1032_),
    .C(RDY_bF$buf5),
    .Y(_1278_)
);

OAI21X1 _2143_ (
    .A(RDY_bF$buf4),
    .B(_1277_),
    .C(_1278_),
    .Y(_1279_)
);

NAND3X1 _2144_ (
    .A(_1276_),
    .B(_1273_),
    .C(_1279_),
    .Y(_1280_)
);

INVX4 _2145_ (
    .A(_981_),
    .Y(_1281_)
);

OAI21X1 _2146_ (
    .A(_882__bF$buf2),
    .B(_961_),
    .C(_853__bF$buf4),
    .Y(_1282_)
);

OAI21X1 _2147_ (
    .A(_853__bF$buf3),
    .B(_1281_),
    .C(_1282_),
    .Y(_1283_)
);

INVX2 _2148_ (
    .A(_1051__bF$buf2),
    .Y(_1284_)
);

NAND2X1 _2149_ (
    .A(RDY_bF$buf3),
    .B(_1284_),
    .Y(_1285_)
);

OAI21X1 _2150_ (
    .A(RDY_bF$buf2),
    .B(_978_),
    .C(_1285_),
    .Y(_1286_)
);

NOR2X1 _2151_ (
    .A(_887__bF$buf0),
    .B(_961_),
    .Y(_1287_)
);

NAND2X1 _2152_ (
    .A(_853__bF$buf2),
    .B(_1287_),
    .Y(_1288_)
);

OAI21X1 _2153_ (
    .A(_853__bF$buf1),
    .B(_894_),
    .C(_1288_),
    .Y(_1289_)
);

NOR2X1 _2154_ (
    .A(_1289_),
    .B(_1286_),
    .Y(_1290_)
);

NAND2X1 _2155_ (
    .A(_1283_),
    .B(_1290_),
    .Y(_1291_)
);

NOR2X1 _2156_ (
    .A(_1280_),
    .B(_1291_),
    .Y(_1292_)
);

NAND3X1 _2157_ (
    .A(_1252_),
    .B(_1292_),
    .C(_1271_),
    .Y(_1293_)
);

NOR3X1 _2158_ (
    .A(_1293_),
    .B(_1249_),
    .C(_1213_),
    .Y(_1294_)
);

INVX1 _2159_ (
    .A(_1294_),
    .Y(_1483_[0])
);

INVX1 _2160_ (
    .A(_1150_),
    .Y(_1295_)
);

OAI21X1 _2161_ (
    .A(_1158_),
    .B(_1152_),
    .C(_1145_),
    .Y(_1296_)
);

NAND2X1 _2162_ (
    .A(_1145_),
    .B(_1154_),
    .Y(_1297_)
);

NOR2X1 _2163_ (
    .A(_1297_),
    .B(_1162_),
    .Y(_1298_)
);

NAND2X1 _2164_ (
    .A(_1296_),
    .B(_1298_),
    .Y(_1299_)
);

NOR2X1 _2165_ (
    .A(_1299_),
    .B(_1295_),
    .Y(_1300_)
);

AOI22X1 _2166_ (
    .A(_853__bF$buf0),
    .B(_1281_),
    .C(_1300_),
    .D(_1129__bF$buf0),
    .Y(_1301_)
);

INVX1 _2167_ (
    .A(_894_),
    .Y(_1302_)
);

NAND2X1 _2168_ (
    .A(_1145_),
    .B(_1161_),
    .Y(_1303_)
);

NOR2X1 _2169_ (
    .A(_1297_),
    .B(_1303_),
    .Y(_1304_)
);

NAND2X1 _2170_ (
    .A(_1296_),
    .B(_1304_),
    .Y(_1305_)
);

NOR2X1 _2171_ (
    .A(_1305_),
    .B(_1295_),
    .Y(_1306_)
);

AOI22X1 _2172_ (
    .A(_853__bF$buf7),
    .B(_1302_),
    .C(_1306_),
    .D(_1129__bF$buf4),
    .Y(_1307_)
);

NAND2X1 _2173_ (
    .A(_1307_),
    .B(_1301_),
    .Y(_1308_)
);

OAI21X1 _2174_ (
    .A(_882__bF$buf1),
    .B(_946_),
    .C(_978_),
    .Y(_1309_)
);

NAND3X1 _2175_ (
    .A(RDY_bF$buf1),
    .B(_1235_),
    .C(_1188_),
    .Y(_1310_)
);

NOR2X1 _2176_ (
    .A(_1196_),
    .B(_1310_),
    .Y(_1311_)
);

NAND2X1 _2177_ (
    .A(_1309_),
    .B(_1311_),
    .Y(_1312_)
);

NAND3X1 _2178_ (
    .A(_853__bF$buf6),
    .B(_926__bF$buf2),
    .C(_890_),
    .Y(_1313_)
);

AND2X2 _2179_ (
    .A(_1147_),
    .B(_1145_),
    .Y(_1314_)
);

NAND2X1 _2180_ (
    .A(_1171_),
    .B(_1314_),
    .Y(_1315_)
);

NOR2X1 _2181_ (
    .A(_1139_),
    .B(_1315_),
    .Y(_1316_)
);

NAND2X1 _2182_ (
    .A(_1164_),
    .B(_1316_),
    .Y(_1317_)
);

OR2X2 _2183_ (
    .A(_1317_),
    .B(_1219__bF$buf1),
    .Y(_1318_)
);

NAND3X1 _2184_ (
    .A(_1312_),
    .B(_1313_),
    .C(_1318_),
    .Y(_1319_)
);

INVX1 _2185_ (
    .A(_1296_),
    .Y(_1320_)
);

NOR2X1 _2186_ (
    .A(_1297_),
    .B(_1320_),
    .Y(_1321_)
);

INVX1 _2187_ (
    .A(_1321_),
    .Y(_1322_)
);

NOR2X1 _2188_ (
    .A(_1139_),
    .B(_1172_),
    .Y(_1323_)
);

NAND2X1 _2189_ (
    .A(_1129__bF$buf3),
    .B(_1323_),
    .Y(_1324_)
);

OAI22X1 _2190_ (
    .A(RDY_bF$buf0),
    .B(_934_),
    .C(_1324_),
    .D(_1322_),
    .Y(_1325_)
);

INVX1 _2191_ (
    .A(_1254_),
    .Y(_1326_)
);

NOR2X1 _2192_ (
    .A(state[4]),
    .B(_989_),
    .Y(_1327_)
);

MUX2X1 _2193_ (
    .A(_942_),
    .B(_1327_),
    .S(RDY_bF$buf8),
    .Y(_1328_)
);

INVX1 _2194_ (
    .A(_1149_),
    .Y(_1329_)
);

NAND2X1 _2195_ (
    .A(_1175_),
    .B(_1329_),
    .Y(_1330_)
);

OAI21X1 _2196_ (
    .A(_1330_),
    .B(_1326_),
    .C(_1328_),
    .Y(_1331_)
);

NOR2X1 _2197_ (
    .A(_1331_),
    .B(_1325_),
    .Y(_1332_)
);

NAND3X1 _2198_ (
    .A(_853__bF$buf5),
    .B(_886__bF$buf0),
    .C(_890_),
    .Y(_1333_)
);

OAI21X1 _2199_ (
    .A(_853__bF$buf4),
    .B(_938_),
    .C(_1333_),
    .Y(_1334_)
);

AND2X2 _2200_ (
    .A(cond_code[2]),
    .B(Z),
    .Y(_1335_)
);

INVX1 _2201_ (
    .A(V),
    .Y(_1336_)
);

NOR2X1 _2202_ (
    .A(cond_code[2]),
    .B(_1336_),
    .Y(_1337_)
);

OAI21X1 _2203_ (
    .A(_1335_),
    .B(_1337_),
    .C(cond_code[1]),
    .Y(_1338_)
);

MUX2X1 _2204_ (
    .A(C),
    .B(N),
    .S(cond_code[2]),
    .Y(_1339_)
);

OAI21X1 _2205_ (
    .A(cond_code[1]),
    .B(_1339_),
    .C(_1338_),
    .Y(_1340_)
);

XOR2X1 _2206_ (
    .A(_1340_),
    .B(cond_code[0]),
    .Y(_1341_)
);

NAND2X1 _2207_ (
    .A(RDY_bF$buf7),
    .B(_943_),
    .Y(_1342_)
);

OAI22X1 _2208_ (
    .A(RDY_bF$buf6),
    .B(_872_),
    .C(_1342_),
    .D(_1341_),
    .Y(_1343_)
);

NOR2X1 _2209_ (
    .A(_1334_),
    .B(_1343_),
    .Y(_1344_)
);

NAND2X1 _2210_ (
    .A(_1344_),
    .B(_1332_),
    .Y(_1345_)
);

NOR3X1 _2211_ (
    .A(_1319_),
    .B(_1308_),
    .C(_1345_),
    .Y(_1346_)
);

NOR2X1 _2212_ (
    .A(_882__bF$buf0),
    .B(_1032_),
    .Y(_1347_)
);

NOR2X1 _2213_ (
    .A(_1168_),
    .B(_1330_),
    .Y(_1348_)
);

AOI22X1 _2214_ (
    .A(_853__bF$buf3),
    .B(_1347_),
    .C(_1348_),
    .D(_1129__bF$buf2),
    .Y(_1349_)
);

INVX1 _2215_ (
    .A(_1175_),
    .Y(_1350_)
);

OAI21X1 _2216_ (
    .A(_1172_),
    .B(_1350_),
    .C(_1315_),
    .Y(_1351_)
);

NOR2X1 _2217_ (
    .A(_1219__bF$buf0),
    .B(_1168_),
    .Y(_1352_)
);

NOR2X1 _2218_ (
    .A(_887__bF$buf4),
    .B(_1032_),
    .Y(_1353_)
);

OAI21X1 _2219_ (
    .A(_887__bF$buf3),
    .B(_936_),
    .C(RDY_bF$buf5),
    .Y(_1354_)
);

OAI21X1 _2220_ (
    .A(RDY_bF$buf4),
    .B(_1353_),
    .C(_1354_),
    .Y(_1355_)
);

OAI21X1 _2221_ (
    .A(_918__bF$buf2),
    .B(_946_),
    .C(RDY_bF$buf3),
    .Y(_1356_)
);

OAI21X1 _2222_ (
    .A(RDY_bF$buf2),
    .B(_1284_),
    .C(_1356_),
    .Y(_1357_)
);

NAND3X1 _2223_ (
    .A(_869__bF$buf0),
    .B(_927_),
    .C(_1356_),
    .Y(_1358_)
);

NAND3X1 _2224_ (
    .A(_1358_),
    .B(_1357_),
    .C(_1355_),
    .Y(_1359_)
);

AOI21X1 _2225_ (
    .A(_1351_),
    .B(_1352_),
    .C(_1359_),
    .Y(_1360_)
);

AND2X2 _2226_ (
    .A(_1349_),
    .B(_1360_),
    .Y(_1361_)
);

NAND2X1 _2227_ (
    .A(_1361_),
    .B(_1346_),
    .Y(_1362_)
);

OR2X2 _2228_ (
    .A(_1362_),
    .B(_1293_),
    .Y(_1483_[1])
);

INVX1 _2229_ (
    .A(_1228_),
    .Y(_1363_)
);

OAI21X1 _2230_ (
    .A(_927_),
    .B(_1037_),
    .C(_886__bF$buf3),
    .Y(_1364_)
);

NAND2X1 _2231_ (
    .A(_881_),
    .B(_905_),
    .Y(_1365_)
);

OAI21X1 _2232_ (
    .A(_916_),
    .B(_918__bF$buf1),
    .C(_1365_),
    .Y(_1366_)
);

NOR2X1 _2233_ (
    .A(_951_),
    .B(_1366_),
    .Y(_1367_)
);

NAND3X1 _2234_ (
    .A(_1363_),
    .B(_1364_),
    .C(_1367_),
    .Y(_1368_)
);

NAND3X1 _2235_ (
    .A(RDY_bF$buf1),
    .B(_943_),
    .C(_1341_),
    .Y(_1369_)
);

OAI21X1 _2236_ (
    .A(_988_),
    .B(_887__bF$buf2),
    .C(_853__bF$buf2),
    .Y(_1370_)
);

NOR2X1 _2237_ (
    .A(_1268_),
    .B(_872_),
    .Y(_1371_)
);

NAND2X1 _2238_ (
    .A(_1370_),
    .B(_1371_),
    .Y(_1372_)
);

OAI21X1 _2239_ (
    .A(_882__bF$buf3),
    .B(_961_),
    .C(RDY_bF$buf0),
    .Y(_1373_)
);

OAI21X1 _2240_ (
    .A(RDY_bF$buf8),
    .B(_1029_),
    .C(_1373_),
    .Y(_1374_)
);

INVX1 _2241_ (
    .A(_1374_),
    .Y(_1375_)
);

OAI21X1 _2242_ (
    .A(_853__bF$buf1),
    .B(_1287_),
    .C(_1370_),
    .Y(_1376_)
);

OAI21X1 _2243_ (
    .A(RDY_bF$buf7),
    .B(_1002__bF$buf0),
    .C(_1376_),
    .Y(_1377_)
);

NOR2X1 _2244_ (
    .A(_1377_),
    .B(_1375_),
    .Y(_1378_)
);

NAND3X1 _2245_ (
    .A(_1369_),
    .B(_1372_),
    .C(_1378_),
    .Y(_1379_)
);

AOI21X1 _2246_ (
    .A(_1311_),
    .B(_1368_),
    .C(_1379_),
    .Y(_1380_)
);

NAND2X1 _2247_ (
    .A(_1220_),
    .B(_1351_),
    .Y(_1381_)
);

INVX1 _2248_ (
    .A(_1138_),
    .Y(_1382_)
);

NOR2X1 _2249_ (
    .A(_1135_),
    .B(_1382_),
    .Y(_1383_)
);

NAND2X1 _2250_ (
    .A(_1383_),
    .B(_1173_),
    .Y(_1384_)
);

OAI21X1 _2251_ (
    .A(_1296_),
    .B(_1215_),
    .C(_1384_),
    .Y(_1385_)
);

AOI21X1 _2252_ (
    .A(_1168_),
    .B(_1180_),
    .C(_1385_),
    .Y(_1386_)
);

NAND2X1 _2253_ (
    .A(_1381_),
    .B(_1386_),
    .Y(_1387_)
);

INVX1 _2254_ (
    .A(_1387_),
    .Y(_1388_)
);

OAI21X1 _2255_ (
    .A(_1150_),
    .B(_1323_),
    .C(_1321_),
    .Y(_1389_)
);

NOR2X1 _2256_ (
    .A(_1219__bF$buf3),
    .B(_1253_),
    .Y(_1390_)
);

NAND3X1 _2257_ (
    .A(_1221_),
    .B(_1390_),
    .C(_1389_),
    .Y(_1391_)
);

INVX1 _2258_ (
    .A(_1316_),
    .Y(_1392_)
);

OR2X2 _2259_ (
    .A(_1392_),
    .B(_1305_),
    .Y(_1393_)
);

NAND2X1 _2260_ (
    .A(_1159_),
    .B(_1303_),
    .Y(_1394_)
);

NOR2X1 _2261_ (
    .A(_1394_),
    .B(_1156_),
    .Y(_1395_)
);

NAND2X1 _2262_ (
    .A(_1150_),
    .B(_1395_),
    .Y(_1396_)
);

NAND3X1 _2263_ (
    .A(_1330_),
    .B(_1396_),
    .C(_1393_),
    .Y(_1397_)
);

NOR2X1 _2264_ (
    .A(_1391_),
    .B(_1397_),
    .Y(_1398_)
);

OAI21X1 _2265_ (
    .A(_1220_),
    .B(_1159_),
    .C(_1299_),
    .Y(_1399_)
);

INVX1 _2266_ (
    .A(_1383_),
    .Y(_1400_)
);

NAND2X1 _2267_ (
    .A(_1350_),
    .B(_1400_),
    .Y(_1401_)
);

NOR2X1 _2268_ (
    .A(_1220_),
    .B(_1315_),
    .Y(_1402_)
);

AOI22X1 _2269_ (
    .A(_1401_),
    .B(_1402_),
    .C(_1399_),
    .D(_1316_),
    .Y(_1403_)
);

AOI21X1 _2270_ (
    .A(_1150_),
    .B(_1164_),
    .C(_1217_),
    .Y(_1404_)
);

NAND3X1 _2271_ (
    .A(_1317_),
    .B(_1403_),
    .C(_1404_),
    .Y(_1405_)
);

INVX1 _2272_ (
    .A(_1405_),
    .Y(_1406_)
);

NAND3X1 _2273_ (
    .A(_1388_),
    .B(_1406_),
    .C(_1398_),
    .Y(_1407_)
);

AOI22X1 _2274_ (
    .A(_853__bF$buf0),
    .B(_951_),
    .C(_1385_),
    .D(_1129__bF$buf1),
    .Y(_1408_)
);

NOR2X1 _2275_ (
    .A(_853__bF$buf7),
    .B(_1200_),
    .Y(_1409_)
);

OAI21X1 _2276_ (
    .A(_882__bF$buf2),
    .B(_880_),
    .C(_853__bF$buf6),
    .Y(_1410_)
);

OAI21X1 _2277_ (
    .A(_853__bF$buf5),
    .B(_1277_),
    .C(_1410_),
    .Y(_1411_)
);

OAI21X1 _2278_ (
    .A(RDY_bF$buf6),
    .B(_1186_),
    .C(_1411_),
    .Y(_1412_)
);

AOI21X1 _2279_ (
    .A(_878_),
    .B(_1409_),
    .C(_1412_),
    .Y(_1413_)
);

AND2X2 _2280_ (
    .A(_1408_),
    .B(_1413_),
    .Y(_1414_)
);

NAND3X1 _2281_ (
    .A(_1380_),
    .B(_1414_),
    .C(_1407_),
    .Y(_1415_)
);

INVX1 _2282_ (
    .A(_1213_),
    .Y(_1416_)
);

NOR2X1 _2283_ (
    .A(_1319_),
    .B(_1345_),
    .Y(_1417_)
);

AND2X2 _2284_ (
    .A(_1223_),
    .B(_1276_),
    .Y(_1418_)
);

AND2X2 _2285_ (
    .A(_1418_),
    .B(_1271_),
    .Y(_1419_)
);

NAND3X1 _2286_ (
    .A(_1416_),
    .B(_1417_),
    .C(_1419_),
    .Y(_1420_)
);

OR2X2 _2287_ (
    .A(_1415_),
    .B(_1420_),
    .Y(_1483_[2])
);

AOI22X1 _2288_ (
    .A(_853__bF$buf4),
    .B(_1039_),
    .C(_1253_),
    .D(_1352_),
    .Y(_1421_)
);

MUX2X1 _2289_ (
    .A(_1240_),
    .B(_959_),
    .S(_853__bF$buf3),
    .Y(_1422_)
);

NAND2X1 _2290_ (
    .A(_1422_),
    .B(_1421_),
    .Y(_1423_)
);

NAND2X1 _2291_ (
    .A(_869__bF$buf3),
    .B(_1037_),
    .Y(_1424_)
);

OAI21X1 _2292_ (
    .A(_996_),
    .B(_887__bF$buf1),
    .C(_853__bF$buf2),
    .Y(_1425_)
);

OAI21X1 _2293_ (
    .A(_853__bF$buf1),
    .B(_1274_),
    .C(_1425_),
    .Y(_1426_)
);

OAI21X1 _2294_ (
    .A(RDY_bF$buf5),
    .B(_1424_),
    .C(_1426_),
    .Y(_1427_)
);

NOR2X1 _2295_ (
    .A(_1427_),
    .B(_1423_),
    .Y(_1428_)
);

NAND2X1 _2296_ (
    .A(_1428_),
    .B(_1361_),
    .Y(_1429_)
);

NOR2X1 _2297_ (
    .A(_1305_),
    .B(_1392_),
    .Y(_1430_)
);

AOI22X1 _2298_ (
    .A(_853__bF$buf0),
    .B(_1224_),
    .C(_1430_),
    .D(_1129__bF$buf0),
    .Y(_1431_)
);

OAI21X1 _2299_ (
    .A(_887__bF$buf0),
    .B(_1035_),
    .C(_853__bF$buf7),
    .Y(_1432_)
);

OAI21X1 _2300_ (
    .A(_853__bF$buf6),
    .B(_1260_),
    .C(_1432_),
    .Y(_1433_)
);

OR2X2 _2301_ (
    .A(_1403_),
    .B(_1219__bF$buf2),
    .Y(_1434_)
);

NAND3X1 _2302_ (
    .A(_1433_),
    .B(_1431_),
    .C(_1434_),
    .Y(_1435_)
);

NOR2X1 _2303_ (
    .A(_1429_),
    .B(_1435_),
    .Y(_1436_)
);

NAND3X1 _2304_ (
    .A(_1346_),
    .B(_1436_),
    .C(_1294_),
    .Y(_1437_)
);

NOR2X1 _2305_ (
    .A(_1219__bF$buf1),
    .B(_1217_),
    .Y(_1438_)
);

NAND3X1 _2306_ (
    .A(_1381_),
    .B(_1438_),
    .C(_1386_),
    .Y(_1439_)
);

NAND2X1 _2307_ (
    .A(_1396_),
    .B(_1317_),
    .Y(_1440_)
);

NOR2X1 _2308_ (
    .A(_1440_),
    .B(_1430_),
    .Y(_1441_)
);

OAI21X1 _2309_ (
    .A(_1314_),
    .B(_1175_),
    .C(_1142_),
    .Y(_1442_)
);

NAND2X1 _2310_ (
    .A(_1442_),
    .B(_1389_),
    .Y(_1443_)
);

INVX1 _2311_ (
    .A(_1164_),
    .Y(_1444_)
);

OAI21X1 _2312_ (
    .A(_1295_),
    .B(_1444_),
    .C(_1221_),
    .Y(_1445_)
);

NOR2X1 _2313_ (
    .A(_1443_),
    .B(_1445_),
    .Y(_1446_)
);

NAND3X1 _2314_ (
    .A(_1403_),
    .B(_1446_),
    .C(_1441_),
    .Y(_1447_)
);

OAI21X1 _2315_ (
    .A(_1439_),
    .B(_1447_),
    .C(_1380_),
    .Y(_1448_)
);

NAND2X1 _2316_ (
    .A(_1433_),
    .B(_1431_),
    .Y(_1449_)
);

INVX1 _2317_ (
    .A(_1449_),
    .Y(_1450_)
);

NAND3X1 _2318_ (
    .A(_1197_),
    .B(_1181_),
    .C(_1211_),
    .Y(_1451_)
);

OR2X2 _2319_ (
    .A(_1258_),
    .B(_1291_),
    .Y(_1452_)
);

NAND3X1 _2320_ (
    .A(_1276_),
    .B(_1357_),
    .C(_1234_),
    .Y(_1453_)
);

NOR3X1 _2321_ (
    .A(_1453_),
    .B(_1452_),
    .C(_1451_),
    .Y(_1454_)
);

INVX1 _2322_ (
    .A(_1332_),
    .Y(_1455_)
);

NOR2X1 _2323_ (
    .A(_1308_),
    .B(_1455_),
    .Y(_1456_)
);

NAND3X1 _2324_ (
    .A(_1450_),
    .B(_1454_),
    .C(_1456_),
    .Y(_1457_)
);

NOR2X1 _2325_ (
    .A(_1448_),
    .B(_1457_),
    .Y(_1458_)
);

OAI21X1 _2326_ (
    .A(_1415_),
    .B(_1437_),
    .C(_1458_),
    .Y(_1483_[3])
);

NAND2X1 _2327_ (
    .A(_1349_),
    .B(_1431_),
    .Y(_1459_)
);

NOR2X1 _2328_ (
    .A(_1319_),
    .B(_1459_),
    .Y(_1460_)
);

NAND3X1 _2329_ (
    .A(_1374_),
    .B(_1204_),
    .C(_1411_),
    .Y(_1461_)
);

AND2X2 _2330_ (
    .A(_1283_),
    .B(_1279_),
    .Y(_1462_)
);

NAND3X1 _2331_ (
    .A(_1265_),
    .B(_1127_),
    .C(_1462_),
    .Y(_1463_)
);

NAND3X1 _2332_ (
    .A(_1226_),
    .B(_1276_),
    .C(_1243_),
    .Y(_1464_)
);

OR2X2 _2333_ (
    .A(_1464_),
    .B(_1463_),
    .Y(_1465_)
);

NOR2X1 _2334_ (
    .A(_1461_),
    .B(_1465_),
    .Y(_1466_)
);

AND2X2 _2335_ (
    .A(_1466_),
    .B(_1301_),
    .Y(_1467_)
);

NOR2X1 _2336_ (
    .A(_1423_),
    .B(_1325_),
    .Y(_1468_)
);

NAND3X1 _2337_ (
    .A(_1460_),
    .B(_1468_),
    .C(_1467_),
    .Y(_1483_[4])
);

AND2X2 _2338_ (
    .A(_1165_),
    .B(_1128_),
    .Y(_1469_)
);

NAND3X1 _2339_ (
    .A(_1469_),
    .B(_1218_),
    .C(_1307_),
    .Y(_1470_)
);

INVX1 _2340_ (
    .A(_942_),
    .Y(_1471_)
);

OAI21X1 _2341_ (
    .A(_853__bF$buf5),
    .B(_1471_),
    .C(_1376_),
    .Y(_1472_)
);

OAI21X1 _2342_ (
    .A(RDY_bF$buf4),
    .B(_1192_),
    .C(_1426_),
    .Y(_1473_)
);

NOR2X1 _2343_ (
    .A(_1473_),
    .B(_1472_),
    .Y(_1474_)
);

NAND3X1 _2344_ (
    .A(_1421_),
    .B(_1255_),
    .C(_1474_),
    .Y(_1475_)
);

NAND2X1 _2345_ (
    .A(_1433_),
    .B(_1355_),
    .Y(_1476_)
);

NOR2X1 _2346_ (
    .A(_1334_),
    .B(_1476_),
    .Y(_1477_)
);

AOI21X1 _2347_ (
    .A(_1205_),
    .B(_1206_),
    .C(_1289_),
    .Y(_1478_)
);

AND2X2 _2348_ (
    .A(_1478_),
    .B(_1262_),
    .Y(_1479_)
);

NOR2X1 _2349_ (
    .A(_1230_),
    .B(_1237_),
    .Y(_1480_)
);

NAND3X1 _2350_ (
    .A(_1477_),
    .B(_1480_),
    .C(_1479_),
    .Y(_1481_)
);

NOR2X1 _2351_ (
    .A(_1475_),
    .B(_1481_),
    .Y(_1482_)
);

NAND3X1 _2352_ (
    .A(_1252_),
    .B(_1408_),
    .C(_1482_),
    .Y(_117_)
);

OR2X2 _2353_ (
    .A(_117_),
    .B(_1470_),
    .Y(_1483_[5])
);

INVX1 _2354_ (
    .A(op[0]),
    .Y(_118_)
);

OAI21X1 _2355_ (
    .A(_916_),
    .B(_918__bF$buf0),
    .C(_911_),
    .Y(_119_)
);

INVX2 _2356_ (
    .A(_119_),
    .Y(_120_)
);

INVX1 _2357_ (
    .A(_1244_),
    .Y(_121_)
);

NAND3X1 _2358_ (
    .A(_1002__bF$buf4),
    .B(_121_),
    .C(_120_),
    .Y(_122_)
);

OAI21X1 _2359_ (
    .A(_118_),
    .B(_120_),
    .C(_122_),
    .Y(alu_op[0])
);

INVX1 _2360_ (
    .A(op[1]),
    .Y(_123_)
);

OAI21X1 _2361_ (
    .A(_123_),
    .B(_120_),
    .C(_122_),
    .Y(alu_op[1])
);

INVX1 _2362_ (
    .A(op[2]),
    .Y(_124_)
);

NOR2X1 _2363_ (
    .A(_882__bF$buf1),
    .B(_961_),
    .Y(_125_)
);

INVX1 _2364_ (
    .A(_125_),
    .Y(_126_)
);

OAI21X1 _2365_ (
    .A(_918__bF$buf3),
    .B(_946_),
    .C(_126_),
    .Y(_127_)
);

INVX2 _2366_ (
    .A(_127_),
    .Y(_128_)
);

NOR2X1 _2367_ (
    .A(_1036_),
    .B(_1353_),
    .Y(_129_)
);

NAND3X1 _2368_ (
    .A(_949_),
    .B(_129_),
    .C(_128_),
    .Y(_130_)
);

AOI21X1 _2369_ (
    .A(backwards),
    .B(_1075_),
    .C(_130_),
    .Y(_131_)
);

OAI21X1 _2370_ (
    .A(_124_),
    .B(_120_),
    .C(_131_),
    .Y(alu_op[2])
);

INVX1 _2371_ (
    .A(op[3]),
    .Y(_132_)
);

NOR2X1 _2372_ (
    .A(_132_),
    .B(_120_),
    .Y(alu_op[3])
);

NOR2X1 _2373_ (
    .A(_1191_),
    .B(_130_),
    .Y(_133_)
);

OAI21X1 _2374_ (
    .A(_882__bF$buf0),
    .B(_901_),
    .C(_1188_),
    .Y(_134_)
);

OAI21X1 _2375_ (
    .A(_1182_),
    .B(_134_),
    .C(store),
    .Y(_135_)
);

NAND2X1 _2376_ (
    .A(_135_),
    .B(_133_),
    .Y(_1687_)
);

NAND2X1 _2377_ (
    .A(_133_),
    .B(_1025_),
    .Y(_136_)
);

OAI21X1 _2378_ (
    .A(_1036_),
    .B(_1281_),
    .C(PC[8]),
    .Y(_137_)
);

NAND2X1 _2379_ (
    .A(_886__bF$buf2),
    .B(_927_),
    .Y(_138_)
);

OAI21X1 _2380_ (
    .A(php),
    .B(_138_),
    .C(_1192_),
    .Y(_139_)
);

INVX1 _2381_ (
    .A(php),
    .Y(_140_)
);

OAI21X1 _2382_ (
    .A(_140_),
    .B(_138_),
    .C(_1051__bF$buf1),
    .Y(_141_)
);

NAND2X1 _2383_ (
    .A(C),
    .B(_141_),
    .Y(_142_)
);

OAI21X1 _2384_ (
    .A(_931_),
    .B(_128_),
    .C(_142_),
    .Y(_143_)
);

AOI21X1 _2385_ (
    .A(ADD[0]),
    .B(_139_),
    .C(_143_),
    .Y(_144_)
);

NAND3X1 _2386_ (
    .A(_137_),
    .B(_144_),
    .C(_136_),
    .Y(_1686_[0])
);

NAND2X1 _2387_ (
    .A(_133_),
    .B(_1063_),
    .Y(_145_)
);

OAI21X1 _2388_ (
    .A(_1036_),
    .B(_1281_),
    .C(PC[9]),
    .Y(_146_)
);

NAND2X1 _2389_ (
    .A(Z),
    .B(_141_),
    .Y(_147_)
);

OAI21X1 _2390_ (
    .A(_968_),
    .B(_128_),
    .C(_147_),
    .Y(_148_)
);

AOI21X1 _2391_ (
    .A(ADD[1]),
    .B(_139_),
    .C(_148_),
    .Y(_149_)
);

NAND3X1 _2392_ (
    .A(_146_),
    .B(_149_),
    .C(_145_),
    .Y(_1686_[1])
);

NAND2X1 _2393_ (
    .A(_133_),
    .B(_1073_),
    .Y(_150_)
);

OAI21X1 _2394_ (
    .A(_1036_),
    .B(_1281_),
    .C(PC[10]),
    .Y(_151_)
);

NAND2X1 _2395_ (
    .A(I),
    .B(_141_),
    .Y(_152_)
);

OAI21X1 _2396_ (
    .A(_970_),
    .B(_128_),
    .C(_152_),
    .Y(_153_)
);

AOI21X1 _2397_ (
    .A(ADD[2]),
    .B(_139_),
    .C(_153_),
    .Y(_154_)
);

NAND3X1 _2398_ (
    .A(_151_),
    .B(_154_),
    .C(_150_),
    .Y(_1686_[2])
);

NAND2X1 _2399_ (
    .A(_133_),
    .B(_1082_),
    .Y(_155_)
);

OAI21X1 _2400_ (
    .A(_1036_),
    .B(_1281_),
    .C(PC[11]),
    .Y(_156_)
);

NAND2X1 _2401_ (
    .A(D),
    .B(_141_),
    .Y(_157_)
);

OAI21X1 _2402_ (
    .A(_971_),
    .B(_128_),
    .C(_157_),
    .Y(_158_)
);

AOI21X1 _2403_ (
    .A(ADD[3]),
    .B(_139_),
    .C(_158_),
    .Y(_159_)
);

NAND3X1 _2404_ (
    .A(_156_),
    .B(_159_),
    .C(_155_),
    .Y(_1686_[3])
);

INVX1 _2405_ (
    .A(_133_),
    .Y(_160_)
);

OAI22X1 _2406_ (
    .A(_140_),
    .B(_138_),
    .C(_1051__bF$buf0),
    .D(_1144_),
    .Y(_161_)
);

AOI21X1 _2407_ (
    .A(_127_),
    .B(PC[4]),
    .C(_161_),
    .Y(_162_)
);

OAI21X1 _2408_ (
    .A(_918__bF$buf2),
    .B(_1035_),
    .C(_981_),
    .Y(_163_)
);

OAI21X1 _2409_ (
    .A(_887__bF$buf4),
    .B(_989_),
    .C(_138_),
    .Y(_164_)
);

AOI22X1 _2410_ (
    .A(_164_),
    .B(ADD[4]),
    .C(PC[12]),
    .D(_163_),
    .Y(_165_)
);

AND2X2 _2411_ (
    .A(_162_),
    .B(_165_),
    .Y(_166_)
);

OAI21X1 _2412_ (
    .A(_160_),
    .B(_1091_),
    .C(_166_),
    .Y(_1686_[4])
);

AOI22X1 _2413_ (
    .A(_164_),
    .B(ADD[5]),
    .C(PC[13]),
    .D(_163_),
    .Y(_167_)
);

OAI21X1 _2414_ (
    .A(_973_),
    .B(_128_),
    .C(_167_),
    .Y(_168_)
);

NOR2X1 _2415_ (
    .A(_141_),
    .B(_168_),
    .Y(_169_)
);

OAI21X1 _2416_ (
    .A(_160_),
    .B(_1099_),
    .C(_169_),
    .Y(_1686_[5])
);

NAND2X1 _2417_ (
    .A(_133_),
    .B(_1106_),
    .Y(_170_)
);

OAI21X1 _2418_ (
    .A(_1036_),
    .B(_1281_),
    .C(PC[14]),
    .Y(_171_)
);

NAND2X1 _2419_ (
    .A(V),
    .B(_141_),
    .Y(_172_)
);

OAI21X1 _2420_ (
    .A(_974_),
    .B(_128_),
    .C(_172_),
    .Y(_173_)
);

AOI21X1 _2421_ (
    .A(ADD[6]),
    .B(_139_),
    .C(_173_),
    .Y(_174_)
);

NAND3X1 _2422_ (
    .A(_171_),
    .B(_174_),
    .C(_170_),
    .Y(_1686_[6])
);

NAND2X1 _2423_ (
    .A(_133_),
    .B(_1116_),
    .Y(_175_)
);

OAI21X1 _2424_ (
    .A(_1036_),
    .B(_1281_),
    .C(PC[15]),
    .Y(_176_)
);

NAND2X1 _2425_ (
    .A(N),
    .B(_141_),
    .Y(_177_)
);

OAI21X1 _2426_ (
    .A(_975_),
    .B(_128_),
    .C(_177_),
    .Y(_178_)
);

AOI21X1 _2427_ (
    .A(AN),
    .B(_139_),
    .C(_178_),
    .Y(_179_)
);

NAND3X1 _2428_ (
    .A(_176_),
    .B(_179_),
    .C(_175_),
    .Y(_1686_[7])
);

INVX1 _2429_ (
    .A(_129_),
    .Y(_180_)
);

OAI21X1 _2430_ (
    .A(_887__bF$buf3),
    .B(_901_),
    .C(_1034_),
    .Y(_181_)
);

OR2X2 _2431_ (
    .A(_180_),
    .B(_181_),
    .Y(_182_)
);

NAND2X1 _2432_ (
    .A(_886__bF$buf1),
    .B(_953_),
    .Y(_183_)
);

NOR2X1 _2433_ (
    .A(_1274_),
    .B(_1048_),
    .Y(_184_)
);

NAND3X1 _2434_ (
    .A(_183_),
    .B(_1227_),
    .C(_184_),
    .Y(_185_)
);

OR2X2 _2435_ (
    .A(_962_),
    .B(_1052_),
    .Y(_186_)
);

NOR2X1 _2436_ (
    .A(_185_),
    .B(_186_),
    .Y(_187_)
);

NAND3X1 _2437_ (
    .A(_898_),
    .B(_990_),
    .C(_1235_),
    .Y(_188_)
);

NOR2X1 _2438_ (
    .A(_1240_),
    .B(_188_),
    .Y(_189_)
);

NAND2X1 _2439_ (
    .A(_189_),
    .B(_187_),
    .Y(_190_)
);

NAND2X1 _2440_ (
    .A(_926__bF$buf1),
    .B(_905_),
    .Y(_191_)
);

NAND3X1 _2441_ (
    .A(_191_),
    .B(_1238_),
    .C(_1363_),
    .Y(_192_)
);

NOR2X1 _2442_ (
    .A(_899_),
    .B(_892_),
    .Y(_193_)
);

NAND2X1 _2443_ (
    .A(_926__bF$buf0),
    .B(_193_),
    .Y(_194_)
);

NAND3X1 _2444_ (
    .A(_194_),
    .B(_121_),
    .C(_884_),
    .Y(_195_)
);

NOR2X1 _2445_ (
    .A(_192_),
    .B(_195_),
    .Y(_196_)
);

OAI21X1 _2446_ (
    .A(_918__bF$buf1),
    .B(_891_),
    .C(_196_),
    .Y(_197_)
);

NOR2X1 _2447_ (
    .A(_190_),
    .B(_197_),
    .Y(_198_)
);

OAI21X1 _2448_ (
    .A(_887__bF$buf2),
    .B(_989_),
    .C(_911_),
    .Y(_199_)
);

NAND3X1 _2449_ (
    .A(_1267_),
    .B(_1123_),
    .C(_1186_),
    .Y(_200_)
);

NOR2X1 _2450_ (
    .A(_200_),
    .B(_199_),
    .Y(_201_)
);

INVX2 _2451_ (
    .A(_201_),
    .Y(_202_)
);

INVX1 _2452_ (
    .A(_182_),
    .Y(_203_)
);

OAI21X1 _2453_ (
    .A(_882__bF$buf3),
    .B(_1032_),
    .C(_1184_),
    .Y(_204_)
);

INVX1 _2454_ (
    .A(_204_),
    .Y(_205_)
);

NAND2X1 _2455_ (
    .A(_205_),
    .B(_203_),
    .Y(_206_)
);

NOR2X1 _2456_ (
    .A(_202_),
    .B(_206_),
    .Y(_207_)
);

NAND2X1 _2457_ (
    .A(_198_),
    .B(_207_),
    .Y(_208_)
);

OAI21X1 _2458_ (
    .A(_190_),
    .B(_197_),
    .C(ADD[0]),
    .Y(_209_)
);

AOI22X1 _2459_ (
    .A(DIMUX[0]),
    .B(_204_),
    .C(_202_),
    .D(ABL[0]),
    .Y(_210_)
);

AND2X2 _2460_ (
    .A(_209_),
    .B(_210_),
    .Y(_211_)
);

OAI21X1 _2461_ (
    .A(_931_),
    .B(_208_),
    .C(_211_),
    .Y(_212_)
);

AOI21X1 _2462_ (
    .A(_1025_),
    .B(_182_),
    .C(_212_),
    .Y(_213_)
);

INVX1 _2463_ (
    .A(_213_),
    .Y(_1685_[0])
);

OAI21X1 _2464_ (
    .A(_190_),
    .B(_197_),
    .C(ADD[1]),
    .Y(_214_)
);

AOI22X1 _2465_ (
    .A(DIMUX[1]),
    .B(_204_),
    .C(_202_),
    .D(ABL[1]),
    .Y(_215_)
);

AND2X2 _2466_ (
    .A(_214_),
    .B(_215_),
    .Y(_216_)
);

OAI21X1 _2467_ (
    .A(_968_),
    .B(_208_),
    .C(_216_),
    .Y(_217_)
);

AOI21X1 _2468_ (
    .A(_1063_),
    .B(_182_),
    .C(_217_),
    .Y(_218_)
);

INVX1 _2469_ (
    .A(_218_),
    .Y(_1685_[1])
);

OAI21X1 _2470_ (
    .A(_190_),
    .B(_197_),
    .C(ADD[2]),
    .Y(_219_)
);

AOI22X1 _2471_ (
    .A(DIMUX[2]),
    .B(_204_),
    .C(_202_),
    .D(ABL[2]),
    .Y(_220_)
);

AND2X2 _2472_ (
    .A(_219_),
    .B(_220_),
    .Y(_221_)
);

OAI21X1 _2473_ (
    .A(_970_),
    .B(_208_),
    .C(_221_),
    .Y(_222_)
);

AOI21X1 _2474_ (
    .A(_1073_),
    .B(_182_),
    .C(_222_),
    .Y(_223_)
);

INVX1 _2475_ (
    .A(_223_),
    .Y(_1685_[2])
);

INVX1 _2476_ (
    .A(_190_),
    .Y(_224_)
);

OR2X2 _2477_ (
    .A(_195_),
    .B(_192_),
    .Y(_225_)
);

NOR2X1 _2478_ (
    .A(_1075_),
    .B(_225_),
    .Y(_226_)
);

NAND2X1 _2479_ (
    .A(_224_),
    .B(_226_),
    .Y(_227_)
);

INVX1 _2480_ (
    .A(ABL[3]),
    .Y(_228_)
);

OAI22X1 _2481_ (
    .A(_857_),
    .B(_205_),
    .C(_228_),
    .D(_201_),
    .Y(_229_)
);

AOI21X1 _2482_ (
    .A(_227_),
    .B(ADD[3]),
    .C(_229_),
    .Y(_230_)
);

OAI21X1 _2483_ (
    .A(_971_),
    .B(_208_),
    .C(_230_),
    .Y(_231_)
);

AOI21X1 _2484_ (
    .A(_1082_),
    .B(_182_),
    .C(_231_),
    .Y(_232_)
);

INVX1 _2485_ (
    .A(_232_),
    .Y(_1685_[3])
);

OAI21X1 _2486_ (
    .A(_190_),
    .B(_197_),
    .C(ADD[4]),
    .Y(_233_)
);

AOI22X1 _2487_ (
    .A(DIMUX[4]),
    .B(_204_),
    .C(_202_),
    .D(ABL[4]),
    .Y(_234_)
);

AND2X2 _2488_ (
    .A(_233_),
    .B(_234_),
    .Y(_235_)
);

OAI21X1 _2489_ (
    .A(_972_),
    .B(_208_),
    .C(_235_),
    .Y(_236_)
);

AOI21X1 _2490_ (
    .A(_1090_),
    .B(_182_),
    .C(_236_),
    .Y(_237_)
);

INVX1 _2491_ (
    .A(_237_),
    .Y(_1685_[4])
);

OAI21X1 _2492_ (
    .A(_190_),
    .B(_197_),
    .C(ADD[5]),
    .Y(_238_)
);

INVX1 _2493_ (
    .A(ABL[5]),
    .Y(_239_)
);

INVX2 _2494_ (
    .A(_200_),
    .Y(_240_)
);

OAI22X1 _2495_ (
    .A(_861_),
    .B(_205_),
    .C(_239_),
    .D(_240_),
    .Y(_241_)
);

AOI21X1 _2496_ (
    .A(ABL[5]),
    .B(_199_),
    .C(_241_),
    .Y(_242_)
);

AND2X2 _2497_ (
    .A(_238_),
    .B(_242_),
    .Y(_243_)
);

OAI21X1 _2498_ (
    .A(_973_),
    .B(_208_),
    .C(_243_),
    .Y(_244_)
);

AOI21X1 _2499_ (
    .A(_1098_),
    .B(_182_),
    .C(_244_),
    .Y(_245_)
);

INVX1 _2500_ (
    .A(_245_),
    .Y(_1685_[5])
);

INVX1 _2501_ (
    .A(ADD[6]),
    .Y(_246_)
);

AOI22X1 _2502_ (
    .A(DIMUX[6]),
    .B(_204_),
    .C(_202_),
    .D(ABL[6]),
    .Y(_247_)
);

OAI21X1 _2503_ (
    .A(_246_),
    .B(_226_),
    .C(_247_),
    .Y(_248_)
);

AOI21X1 _2504_ (
    .A(ADD[6]),
    .B(_190_),
    .C(_248_),
    .Y(_249_)
);

OAI21X1 _2505_ (
    .A(_974_),
    .B(_208_),
    .C(_249_),
    .Y(_250_)
);

AOI21X1 _2506_ (
    .A(_1106_),
    .B(_182_),
    .C(_250_),
    .Y(_251_)
);

INVX1 _2507_ (
    .A(_251_),
    .Y(_1685_[6])
);

NAND2X1 _2508_ (
    .A(AN),
    .B(_190_),
    .Y(_252_)
);

INVX1 _2509_ (
    .A(ABL[7]),
    .Y(_253_)
);

OAI22X1 _2510_ (
    .A(_864_),
    .B(_205_),
    .C(_253_),
    .D(_201_),
    .Y(_254_)
);

AOI21X1 _2511_ (
    .A(_197_),
    .B(AN),
    .C(_254_),
    .Y(_255_)
);

NAND2X1 _2512_ (
    .A(_252_),
    .B(_255_),
    .Y(_256_)
);

INVX1 _2513_ (
    .A(_256_),
    .Y(_257_)
);

OAI21X1 _2514_ (
    .A(_975_),
    .B(_208_),
    .C(_257_),
    .Y(_258_)
);

AOI21X1 _2515_ (
    .A(_1116_),
    .B(_182_),
    .C(_258_),
    .Y(_259_)
);

INVX1 _2516_ (
    .A(_259_),
    .Y(_1685_[7])
);

INVX1 _2517_ (
    .A(PC[8]),
    .Y(_260_)
);

NOR2X1 _2518_ (
    .A(_260_),
    .B(_208_),
    .Y(_261_)
);

AOI21X1 _2519_ (
    .A(ABH[0]),
    .B(_199_),
    .C(_182_),
    .Y(_262_)
);

INVX1 _2520_ (
    .A(ADD[0]),
    .Y(_263_)
);

OAI21X1 _2521_ (
    .A(_263_),
    .B(_240_),
    .C(_1057_),
    .Y(_264_)
);

AOI21X1 _2522_ (
    .A(_225_),
    .B(DIMUX[0]),
    .C(_264_),
    .Y(_265_)
);

NAND3X1 _2523_ (
    .A(_187_),
    .B(_262_),
    .C(_265_),
    .Y(_266_)
);

OR2X2 _2524_ (
    .A(_261_),
    .B(_266_),
    .Y(_1685_[8])
);

INVX1 _2525_ (
    .A(PC[9]),
    .Y(_267_)
);

INVX2 _2526_ (
    .A(_199_),
    .Y(_268_)
);

AOI21X1 _2527_ (
    .A(_200_),
    .B(ADD[1]),
    .C(_1066_),
    .Y(_269_)
);

OAI21X1 _2528_ (
    .A(_1065_),
    .B(_268_),
    .C(_269_),
    .Y(_270_)
);

AOI21X1 _2529_ (
    .A(_225_),
    .B(DIMUX[1]),
    .C(_270_),
    .Y(_271_)
);

OAI21X1 _2530_ (
    .A(_267_),
    .B(_208_),
    .C(_271_),
    .Y(_1685_[9])
);

INVX1 _2531_ (
    .A(PC[10]),
    .Y(_272_)
);

INVX1 _2532_ (
    .A(ABH[2]),
    .Y(_273_)
);

AOI22X1 _2533_ (
    .A(ABH[2]),
    .B(_1075_),
    .C(_200_),
    .D(ADD[2]),
    .Y(_274_)
);

OAI21X1 _2534_ (
    .A(_273_),
    .B(_268_),
    .C(_274_),
    .Y(_275_)
);

AOI21X1 _2535_ (
    .A(_225_),
    .B(DIMUX[2]),
    .C(_275_),
    .Y(_276_)
);

OAI21X1 _2536_ (
    .A(_272_),
    .B(_208_),
    .C(_276_),
    .Y(_1685_[10])
);

INVX1 _2537_ (
    .A(PC[11]),
    .Y(_277_)
);

NAND2X1 _2538_ (
    .A(ABH[3]),
    .B(_199_),
    .Y(_278_)
);

AOI22X1 _2539_ (
    .A(ABH[3]),
    .B(_1075_),
    .C(_200_),
    .D(ADD[3]),
    .Y(_279_)
);

AND2X2 _2540_ (
    .A(_279_),
    .B(_278_),
    .Y(_280_)
);

OAI21X1 _2541_ (
    .A(_857_),
    .B(_196_),
    .C(_280_),
    .Y(_281_)
);

INVX1 _2542_ (
    .A(_281_),
    .Y(_282_)
);

OAI21X1 _2543_ (
    .A(_277_),
    .B(_208_),
    .C(_282_),
    .Y(_1685_[11])
);

INVX1 _2544_ (
    .A(PC[12]),
    .Y(_283_)
);

INVX1 _2545_ (
    .A(ABH[4]),
    .Y(_284_)
);

INVX1 _2546_ (
    .A(ADD[4]),
    .Y(_285_)
);

OAI21X1 _2547_ (
    .A(_192_),
    .B(_195_),
    .C(DIMUX[4]),
    .Y(_286_)
);

OAI21X1 _2548_ (
    .A(_285_),
    .B(_240_),
    .C(_286_),
    .Y(_287_)
);

AOI21X1 _2549_ (
    .A(ABH[4]),
    .B(_1075_),
    .C(_287_),
    .Y(_288_)
);

OAI21X1 _2550_ (
    .A(_284_),
    .B(_268_),
    .C(_288_),
    .Y(_289_)
);

INVX1 _2551_ (
    .A(_289_),
    .Y(_290_)
);

OAI21X1 _2552_ (
    .A(_283_),
    .B(_208_),
    .C(_290_),
    .Y(_1685_[12])
);

INVX1 _2553_ (
    .A(PC[13]),
    .Y(_291_)
);

INVX1 _2554_ (
    .A(ABH[5]),
    .Y(_292_)
);

INVX1 _2555_ (
    .A(ADD[5]),
    .Y(_293_)
);

OAI21X1 _2556_ (
    .A(_192_),
    .B(_195_),
    .C(DIMUX[5]),
    .Y(_294_)
);

OAI21X1 _2557_ (
    .A(_293_),
    .B(_240_),
    .C(_294_),
    .Y(_295_)
);

AOI21X1 _2558_ (
    .A(ABH[5]),
    .B(_1075_),
    .C(_295_),
    .Y(_296_)
);

OAI21X1 _2559_ (
    .A(_292_),
    .B(_268_),
    .C(_296_),
    .Y(_297_)
);

INVX1 _2560_ (
    .A(_297_),
    .Y(_298_)
);

OAI21X1 _2561_ (
    .A(_291_),
    .B(_208_),
    .C(_298_),
    .Y(_1685_[13])
);

INVX1 _2562_ (
    .A(PC[14]),
    .Y(_299_)
);

AOI21X1 _2563_ (
    .A(_200_),
    .B(ADD[6]),
    .C(_1109_),
    .Y(_300_)
);

OAI21X1 _2564_ (
    .A(_1108_),
    .B(_268_),
    .C(_300_),
    .Y(_301_)
);

AOI21X1 _2565_ (
    .A(_225_),
    .B(DIMUX[6]),
    .C(_301_),
    .Y(_302_)
);

OAI21X1 _2566_ (
    .A(_299_),
    .B(_208_),
    .C(_302_),
    .Y(_1685_[14])
);

INVX1 _2567_ (
    .A(PC[15]),
    .Y(_303_)
);

INVX1 _2568_ (
    .A(AN),
    .Y(_304_)
);

OAI21X1 _2569_ (
    .A(_192_),
    .B(_195_),
    .C(DIMUX[7]),
    .Y(_305_)
);

OAI21X1 _2570_ (
    .A(_304_),
    .B(_240_),
    .C(_305_),
    .Y(_306_)
);

NOR2X1 _2571_ (
    .A(_1119_),
    .B(_306_),
    .Y(_307_)
);

OAI21X1 _2572_ (
    .A(_1118_),
    .B(_268_),
    .C(_307_),
    .Y(_308_)
);

INVX1 _2573_ (
    .A(_308_),
    .Y(_309_)
);

OAI21X1 _2574_ (
    .A(_303_),
    .B(_208_),
    .C(_309_),
    .Y(_1685_[15])
);

AND2X2 _2575_ (
    .A(adc_sbc),
    .B(D),
    .Y(_0_)
);

INVX1 _2576_ (
    .A(adc_bcd),
    .Y(_310_)
);

NOR2X1 _2577_ (
    .A(_310_),
    .B(_1031_),
    .Y(\u_ALU8.BCD )
);

INVX1 _2578_ (
    .A(shift_right),
    .Y(_311_)
);

NOR2X1 _2579_ (
    .A(_311_),
    .B(_120_),
    .Y(alu_shift_right)
);

INVX8 _2580_ (
    .A(reset),
    .Y(_1_)
);

OAI21X1 _2581_ (
    .A(_900_),
    .B(_1037_),
    .C(_869__bF$buf2),
    .Y(_312_)
);

OAI21X1 _2582_ (
    .A(_872_),
    .B(_1268_),
    .C(_312_),
    .Y(_313_)
);

AOI21X1 _2583_ (
    .A(_917_),
    .B(_1193_),
    .C(_313_),
    .Y(_314_)
);

OAI21X1 _2584_ (
    .A(_886__bF$buf0),
    .B(_926__bF$buf3),
    .C(_193_),
    .Y(_315_)
);

OAI21X1 _2585_ (
    .A(_1002__bF$buf3),
    .B(_1133_),
    .C(_315_),
    .Y(_316_)
);

NAND3X1 _2586_ (
    .A(_978_),
    .B(_1365_),
    .C(_992_),
    .Y(_317_)
);

NOR2X1 _2587_ (
    .A(_316_),
    .B(_317_),
    .Y(_318_)
);

NAND2X1 _2588_ (
    .A(_318_),
    .B(_314_),
    .Y(_319_)
);

OAI22X1 _2589_ (
    .A(_886__bF$buf3),
    .B(_926__bF$buf2),
    .C(_1193_),
    .D(_193_),
    .Y(_320_)
);

NAND3X1 _2590_ (
    .A(_872_),
    .B(_191_),
    .C(_320_),
    .Y(_321_)
);

NAND3X1 _2591_ (
    .A(_1002__bF$buf2),
    .B(_1267_),
    .C(_1051__bF$buf3),
    .Y(_322_)
);

NOR2X1 _2592_ (
    .A(_322_),
    .B(_321_),
    .Y(_323_)
);

INVX2 _2593_ (
    .A(_323_),
    .Y(_324_)
);

NOR3X1 _2594_ (
    .A(_875_),
    .B(_867_),
    .C(_918__bF$buf0),
    .Y(_325_)
);

AOI22X1 _2595_ (
    .A(PC[0]),
    .B(_325_),
    .C(_321_),
    .D(ADD[0]),
    .Y(_326_)
);

AND2X2 _2596_ (
    .A(_1133_),
    .B(ABL[0]),
    .Y(_327_)
);

NOR2X1 _2597_ (
    .A(_931_),
    .B(_1133_),
    .Y(_328_)
);

OAI21X1 _2598_ (
    .A(_328_),
    .B(_327_),
    .C(_1008_),
    .Y(_329_)
);

NAND3X1 _2599_ (
    .A(_326_),
    .B(_329_),
    .C(_324_),
    .Y(_330_)
);

NAND2X1 _2600_ (
    .A(_931_),
    .B(_323_),
    .Y(_331_)
);

AOI21X1 _2601_ (
    .A(_330_),
    .B(_331_),
    .C(_319_),
    .Y(_332_)
);

NAND3X1 _2602_ (
    .A(_869__bF$buf1),
    .B(_953_),
    .C(_1145_),
    .Y(_333_)
);

OAI21X1 _2603_ (
    .A(_918__bF$buf3),
    .B(_1259_),
    .C(_333_),
    .Y(_334_)
);

INVX1 _2604_ (
    .A(_334_),
    .Y(_335_)
);

OAI21X1 _2605_ (
    .A(_322_),
    .B(_321_),
    .C(_335_),
    .Y(_336_)
);

NAND2X1 _2606_ (
    .A(PC[0]),
    .B(_336_),
    .Y(_337_)
);

NOR2X1 _2607_ (
    .A(_1002__bF$buf1),
    .B(_1145_),
    .Y(_338_)
);

AOI22X1 _2608_ (
    .A(ABL[0]),
    .B(_338_),
    .C(_321_),
    .D(ADD[0]),
    .Y(_339_)
);

AOI22X1 _2609_ (
    .A(_314_),
    .B(_318_),
    .C(_337_),
    .D(_339_),
    .Y(_340_)
);

INVX1 _2610_ (
    .A(_340_),
    .Y(_341_)
);

NAND2X1 _2611_ (
    .A(RDY_bF$buf3),
    .B(_341_),
    .Y(_342_)
);

OAI22X1 _2612_ (
    .A(RDY_bF$buf2),
    .B(_931_),
    .C(_332_),
    .D(_342_),
    .Y(_2_)
);

INVX2 _2613_ (
    .A(_336_),
    .Y(_343_)
);

NAND2X1 _2614_ (
    .A(ABL[1]),
    .B(_338_),
    .Y(_344_)
);

OAI21X1 _2615_ (
    .A(res),
    .B(_1051__bF$buf2),
    .C(_344_),
    .Y(_345_)
);

AOI21X1 _2616_ (
    .A(ADD[1]),
    .B(_321_),
    .C(_345_),
    .Y(_346_)
);

OAI21X1 _2617_ (
    .A(_968_),
    .B(_343_),
    .C(_346_),
    .Y(_347_)
);

NOR2X1 _2618_ (
    .A(_347_),
    .B(_340_),
    .Y(_348_)
);

NAND2X1 _2619_ (
    .A(_347_),
    .B(_340_),
    .Y(_349_)
);

NAND2X1 _2620_ (
    .A(RDY_bF$buf1),
    .B(_349_),
    .Y(_350_)
);

OAI22X1 _2621_ (
    .A(RDY_bF$buf0),
    .B(_968_),
    .C(_348_),
    .D(_350_),
    .Y(_3_)
);

NAND2X1 _2622_ (
    .A(PC[2]),
    .B(_853__bF$buf4),
    .Y(_351_)
);

NOR2X1 _2623_ (
    .A(res),
    .B(_1132_),
    .Y(_352_)
);

NAND2X1 _2624_ (
    .A(ABL[2]),
    .B(_338_),
    .Y(_353_)
);

OAI21X1 _2625_ (
    .A(_1051__bF$buf1),
    .B(_352_),
    .C(_353_),
    .Y(_354_)
);

AOI21X1 _2626_ (
    .A(ADD[2]),
    .B(_321_),
    .C(_354_),
    .Y(_355_)
);

OAI21X1 _2627_ (
    .A(_970_),
    .B(_343_),
    .C(_355_),
    .Y(_356_)
);

XOR2X1 _2628_ (
    .A(_349_),
    .B(_356_),
    .Y(_357_)
);

OAI21X1 _2629_ (
    .A(_853__bF$buf3),
    .B(_357_),
    .C(_351_),
    .Y(_4_)
);

INVX1 _2630_ (
    .A(_349_),
    .Y(_358_)
);

INVX2 _2631_ (
    .A(_338_),
    .Y(_359_)
);

OAI21X1 _2632_ (
    .A(_228_),
    .B(_359_),
    .C(_1051__bF$buf0),
    .Y(_360_)
);

AOI21X1 _2633_ (
    .A(ADD[3]),
    .B(_321_),
    .C(_360_),
    .Y(_361_)
);

OAI21X1 _2634_ (
    .A(_971_),
    .B(_343_),
    .C(_361_),
    .Y(_362_)
);

AOI21X1 _2635_ (
    .A(_358_),
    .B(_356_),
    .C(_362_),
    .Y(_363_)
);

NAND2X1 _2636_ (
    .A(PC[2]),
    .B(_336_),
    .Y(_364_)
);

NAND2X1 _2637_ (
    .A(PC[3]),
    .B(_336_),
    .Y(_365_)
);

AOI22X1 _2638_ (
    .A(_364_),
    .B(_355_),
    .C(_365_),
    .D(_361_),
    .Y(_366_)
);

NAND3X1 _2639_ (
    .A(_347_),
    .B(_340_),
    .C(_366_),
    .Y(_367_)
);

NAND2X1 _2640_ (
    .A(RDY_bF$buf8),
    .B(_367_),
    .Y(_368_)
);

OAI22X1 _2641_ (
    .A(RDY_bF$buf7),
    .B(_971_),
    .C(_368_),
    .D(_363_),
    .Y(_5_)
);

NAND2X1 _2642_ (
    .A(PC[4]),
    .B(_853__bF$buf2),
    .Y(_369_)
);

INVX1 _2643_ (
    .A(ABL[4]),
    .Y(_370_)
);

OAI21X1 _2644_ (
    .A(_370_),
    .B(_359_),
    .C(_1051__bF$buf3),
    .Y(_371_)
);

AOI21X1 _2645_ (
    .A(ADD[4]),
    .B(_321_),
    .C(_371_),
    .Y(_372_)
);

OAI21X1 _2646_ (
    .A(_972_),
    .B(_343_),
    .C(_372_),
    .Y(_373_)
);

XOR2X1 _2647_ (
    .A(_367_),
    .B(_373_),
    .Y(_374_)
);

OAI21X1 _2648_ (
    .A(_853__bF$buf1),
    .B(_374_),
    .C(_369_),
    .Y(_6_)
);

INVX1 _2649_ (
    .A(_367_),
    .Y(_375_)
);

OAI21X1 _2650_ (
    .A(_239_),
    .B(_359_),
    .C(_1051__bF$buf2),
    .Y(_376_)
);

AOI21X1 _2651_ (
    .A(ADD[5]),
    .B(_321_),
    .C(_376_),
    .Y(_377_)
);

OAI21X1 _2652_ (
    .A(_973_),
    .B(_343_),
    .C(_377_),
    .Y(_378_)
);

AOI21X1 _2653_ (
    .A(_375_),
    .B(_373_),
    .C(_378_),
    .Y(_379_)
);

NAND2X1 _2654_ (
    .A(PC[4]),
    .B(_336_),
    .Y(_380_)
);

NAND2X1 _2655_ (
    .A(PC[5]),
    .B(_336_),
    .Y(_381_)
);

AOI22X1 _2656_ (
    .A(_380_),
    .B(_372_),
    .C(_381_),
    .D(_377_),
    .Y(_382_)
);

INVX1 _2657_ (
    .A(_382_),
    .Y(_383_)
);

OAI21X1 _2658_ (
    .A(_383_),
    .B(_367_),
    .C(RDY_bF$buf6),
    .Y(_384_)
);

OAI22X1 _2659_ (
    .A(RDY_bF$buf5),
    .B(_973_),
    .C(_384_),
    .D(_379_),
    .Y(_7_)
);

NOR2X1 _2660_ (
    .A(_383_),
    .B(_367_),
    .Y(_385_)
);

INVX1 _2661_ (
    .A(ABL[6]),
    .Y(_386_)
);

OAI21X1 _2662_ (
    .A(_386_),
    .B(_359_),
    .C(_1051__bF$buf1),
    .Y(_387_)
);

AOI21X1 _2663_ (
    .A(ADD[6]),
    .B(_321_),
    .C(_387_),
    .Y(_388_)
);

OAI21X1 _2664_ (
    .A(_974_),
    .B(_343_),
    .C(_388_),
    .Y(_389_)
);

NOR2X1 _2665_ (
    .A(_389_),
    .B(_385_),
    .Y(_390_)
);

NAND2X1 _2666_ (
    .A(_389_),
    .B(_385_),
    .Y(_391_)
);

NAND2X1 _2667_ (
    .A(RDY_bF$buf4),
    .B(_391_),
    .Y(_392_)
);

OAI22X1 _2668_ (
    .A(RDY_bF$buf3),
    .B(_974_),
    .C(_390_),
    .D(_392_),
    .Y(_8_)
);

OAI21X1 _2669_ (
    .A(_253_),
    .B(_359_),
    .C(_1051__bF$buf0),
    .Y(_393_)
);

AOI21X1 _2670_ (
    .A(AN),
    .B(_321_),
    .C(_393_),
    .Y(_394_)
);

OAI21X1 _2671_ (
    .A(_975_),
    .B(_343_),
    .C(_394_),
    .Y(_395_)
);

INVX1 _2672_ (
    .A(_395_),
    .Y(_396_)
);

NAND2X1 _2673_ (
    .A(_396_),
    .B(_391_),
    .Y(_397_)
);

NAND3X1 _2674_ (
    .A(_389_),
    .B(_395_),
    .C(_385_),
    .Y(_398_)
);

NAND3X1 _2675_ (
    .A(RDY_bF$buf2),
    .B(_398_),
    .C(_397_),
    .Y(_399_)
);

OAI21X1 _2676_ (
    .A(RDY_bF$buf1),
    .B(_975_),
    .C(_399_),
    .Y(_9_)
);

AOI21X1 _2677_ (
    .A(_320_),
    .B(_191_),
    .C(_932_),
    .Y(_400_)
);

OAI22X1 _2678_ (
    .A(_1055_),
    .B(_872_),
    .C(_260_),
    .D(_333_),
    .Y(_401_)
);

NAND3X1 _2679_ (
    .A(ADD[0]),
    .B(_869__bF$buf0),
    .C(_905_),
    .Y(_402_)
);

NAND3X1 _2680_ (
    .A(ABH[0]),
    .B(_1133_),
    .C(_1008_),
    .Y(_403_)
);

NAND3X1 _2681_ (
    .A(_1051__bF$buf3),
    .B(_402_),
    .C(_403_),
    .Y(_404_)
);

NOR3X1 _2682_ (
    .A(_401_),
    .B(_404_),
    .C(_400_),
    .Y(_405_)
);

OAI21X1 _2683_ (
    .A(_260_),
    .B(_324_),
    .C(_405_),
    .Y(_406_)
);

NAND2X1 _2684_ (
    .A(PC[6]),
    .B(_336_),
    .Y(_407_)
);

NAND2X1 _2685_ (
    .A(PC[7]),
    .B(_336_),
    .Y(_408_)
);

AOI22X1 _2686_ (
    .A(_407_),
    .B(_388_),
    .C(_408_),
    .D(_394_),
    .Y(_409_)
);

NAND2X1 _2687_ (
    .A(_382_),
    .B(_409_),
    .Y(_410_)
);

OR2X2 _2688_ (
    .A(_367_),
    .B(_410_),
    .Y(_411_)
);

NOR2X1 _2689_ (
    .A(_406_),
    .B(_411_),
    .Y(_412_)
);

AOI22X1 _2690_ (
    .A(_887__bF$buf1),
    .B(_882__bF$buf2),
    .C(_946_),
    .D(_916_),
    .Y(_413_)
);

NOR3X1 _2691_ (
    .A(_1075_),
    .B(_1264_),
    .C(_413_),
    .Y(_414_)
);

INVX1 _2692_ (
    .A(_322_),
    .Y(_415_)
);

NAND3X1 _2693_ (
    .A(PC[8]),
    .B(_415_),
    .C(_414_),
    .Y(_416_)
);

NOR2X1 _2694_ (
    .A(_410_),
    .B(_367_),
    .Y(_417_)
);

AOI21X1 _2695_ (
    .A(_405_),
    .B(_416_),
    .C(_417_),
    .Y(_418_)
);

OAI21X1 _2696_ (
    .A(_418_),
    .B(_412_),
    .C(RDY_bF$buf0),
    .Y(_419_)
);

OAI21X1 _2697_ (
    .A(RDY_bF$buf8),
    .B(_260_),
    .C(_419_),
    .Y(_10_)
);

INVX1 _2698_ (
    .A(_398_),
    .Y(_420_)
);

AOI21X1 _2699_ (
    .A(_320_),
    .B(_191_),
    .C(_969_),
    .Y(_421_)
);

OAI22X1 _2700_ (
    .A(_1065_),
    .B(_872_),
    .C(_267_),
    .D(_333_),
    .Y(_422_)
);

NAND3X1 _2701_ (
    .A(ADD[1]),
    .B(_869__bF$buf3),
    .C(_905_),
    .Y(_423_)
);

NAND3X1 _2702_ (
    .A(ABH[1]),
    .B(_1133_),
    .C(_1008_),
    .Y(_424_)
);

NAND3X1 _2703_ (
    .A(_1051__bF$buf2),
    .B(_423_),
    .C(_424_),
    .Y(_425_)
);

NOR3X1 _2704_ (
    .A(_422_),
    .B(_425_),
    .C(_421_),
    .Y(_426_)
);

OAI21X1 _2705_ (
    .A(_267_),
    .B(_324_),
    .C(_426_),
    .Y(_427_)
);

AOI21X1 _2706_ (
    .A(_420_),
    .B(_406_),
    .C(_427_),
    .Y(_428_)
);

NAND3X1 _2707_ (
    .A(PC[9]),
    .B(_415_),
    .C(_414_),
    .Y(_429_)
);

AOI22X1 _2708_ (
    .A(_405_),
    .B(_416_),
    .C(_426_),
    .D(_429_),
    .Y(_430_)
);

INVX1 _2709_ (
    .A(_430_),
    .Y(_431_)
);

OAI21X1 _2710_ (
    .A(_431_),
    .B(_398_),
    .C(RDY_bF$buf7),
    .Y(_432_)
);

OAI22X1 _2711_ (
    .A(RDY_bF$buf6),
    .B(_267_),
    .C(_432_),
    .D(_428_),
    .Y(_11_)
);

NAND2X1 _2712_ (
    .A(PC[10]),
    .B(_853__bF$buf0),
    .Y(_433_)
);

OAI21X1 _2713_ (
    .A(_1264_),
    .B(_413_),
    .C(DIMUX[2]),
    .Y(_434_)
);

NOR3X1 _2714_ (
    .A(_273_),
    .B(_1002__bF$buf0),
    .C(_1145_),
    .Y(_435_)
);

OAI21X1 _2715_ (
    .A(_272_),
    .B(_333_),
    .C(_1076_),
    .Y(_436_)
);

INVX1 _2716_ (
    .A(ADD[2]),
    .Y(_437_)
);

OAI21X1 _2717_ (
    .A(_437_),
    .B(_1267_),
    .C(_1051__bF$buf1),
    .Y(_438_)
);

NOR3X1 _2718_ (
    .A(_435_),
    .B(_438_),
    .C(_436_),
    .Y(_439_)
);

NAND3X1 _2719_ (
    .A(PC[10]),
    .B(_415_),
    .C(_414_),
    .Y(_440_)
);

NAND3X1 _2720_ (
    .A(_434_),
    .B(_440_),
    .C(_439_),
    .Y(_441_)
);

NAND2X1 _2721_ (
    .A(_430_),
    .B(_417_),
    .Y(_442_)
);

XOR2X1 _2722_ (
    .A(_442_),
    .B(_441_),
    .Y(_443_)
);

OAI21X1 _2723_ (
    .A(_853__bF$buf7),
    .B(_443_),
    .C(_433_),
    .Y(_12_)
);

NOR2X1 _2724_ (
    .A(_431_),
    .B(_398_),
    .Y(_444_)
);

AOI22X1 _2725_ (
    .A(_1008_),
    .B(_1145_),
    .C(_414_),
    .D(_415_),
    .Y(_445_)
);

OAI21X1 _2726_ (
    .A(_882__bF$buf1),
    .B(_1259_),
    .C(_320_),
    .Y(_446_)
);

AOI22X1 _2727_ (
    .A(ADD[3]),
    .B(_325_),
    .C(_338_),
    .D(ABH[3]),
    .Y(_447_)
);

NAND3X1 _2728_ (
    .A(_1051__bF$buf0),
    .B(_1084_),
    .C(_447_),
    .Y(_448_)
);

AOI21X1 _2729_ (
    .A(DIMUX[3]),
    .B(_446_),
    .C(_448_),
    .Y(_449_)
);

OAI21X1 _2730_ (
    .A(_277_),
    .B(_445_),
    .C(_449_),
    .Y(_450_)
);

AOI21X1 _2731_ (
    .A(_444_),
    .B(_441_),
    .C(_450_),
    .Y(_451_)
);

NAND3X1 _2732_ (
    .A(_441_),
    .B(_450_),
    .C(_430_),
    .Y(_452_)
);

OAI21X1 _2733_ (
    .A(_452_),
    .B(_398_),
    .C(RDY_bF$buf5),
    .Y(_453_)
);

OAI22X1 _2734_ (
    .A(RDY_bF$buf4),
    .B(_277_),
    .C(_453_),
    .D(_451_),
    .Y(_13_)
);

OAI21X1 _2735_ (
    .A(_283_),
    .B(_333_),
    .C(_1092_),
    .Y(_454_)
);

AOI21X1 _2736_ (
    .A(ADD[4]),
    .B(_325_),
    .C(_1284_),
    .Y(_455_)
);

OAI21X1 _2737_ (
    .A(_284_),
    .B(_359_),
    .C(_455_),
    .Y(_456_)
);

OR2X2 _2738_ (
    .A(_456_),
    .B(_454_),
    .Y(_457_)
);

AOI21X1 _2739_ (
    .A(DIMUX[4]),
    .B(_446_),
    .C(_457_),
    .Y(_458_)
);

OAI21X1 _2740_ (
    .A(_283_),
    .B(_324_),
    .C(_458_),
    .Y(_459_)
);

NOR3X1 _2741_ (
    .A(_452_),
    .B(_410_),
    .C(_367_),
    .Y(_460_)
);

XOR2X1 _2742_ (
    .A(_460_),
    .B(_459_),
    .Y(_461_)
);

NAND2X1 _2743_ (
    .A(RDY_bF$buf3),
    .B(_461_),
    .Y(_462_)
);

OAI21X1 _2744_ (
    .A(RDY_bF$buf2),
    .B(_283_),
    .C(_462_),
    .Y(_14_)
);

NAND2X1 _2745_ (
    .A(PC[13]),
    .B(_853__bF$buf6),
    .Y(_463_)
);

OAI21X1 _2746_ (
    .A(_291_),
    .B(_333_),
    .C(_1100_),
    .Y(_464_)
);

AOI21X1 _2747_ (
    .A(ADD[5]),
    .B(_325_),
    .C(_1284_),
    .Y(_465_)
);

OAI21X1 _2748_ (
    .A(_292_),
    .B(_359_),
    .C(_465_),
    .Y(_466_)
);

OR2X2 _2749_ (
    .A(_466_),
    .B(_464_),
    .Y(_467_)
);

AOI21X1 _2750_ (
    .A(DIMUX[5]),
    .B(_446_),
    .C(_467_),
    .Y(_468_)
);

OAI21X1 _2751_ (
    .A(_291_),
    .B(_324_),
    .C(_468_),
    .Y(_469_)
);

NAND2X1 _2752_ (
    .A(_459_),
    .B(_460_),
    .Y(_470_)
);

XOR2X1 _2753_ (
    .A(_470_),
    .B(_469_),
    .Y(_471_)
);

OAI21X1 _2754_ (
    .A(_853__bF$buf5),
    .B(_471_),
    .C(_463_),
    .Y(_15_)
);

NAND2X1 _2755_ (
    .A(PC[12]),
    .B(_323_),
    .Y(_472_)
);

NAND2X1 _2756_ (
    .A(PC[13]),
    .B(_323_),
    .Y(_473_)
);

AOI22X1 _2757_ (
    .A(_458_),
    .B(_472_),
    .C(_468_),
    .D(_473_),
    .Y(_474_)
);

NOR2X1 _2758_ (
    .A(_299_),
    .B(_445_),
    .Y(_475_)
);

OAI21X1 _2759_ (
    .A(_1264_),
    .B(_413_),
    .C(DIMUX[6]),
    .Y(_476_)
);

NOR2X1 _2760_ (
    .A(_1284_),
    .B(_1109_),
    .Y(_477_)
);

AOI22X1 _2761_ (
    .A(ADD[6]),
    .B(_325_),
    .C(_338_),
    .D(ABH[6]),
    .Y(_478_)
);

NAND3X1 _2762_ (
    .A(_476_),
    .B(_478_),
    .C(_477_),
    .Y(_479_)
);

NOR2X1 _2763_ (
    .A(_479_),
    .B(_475_),
    .Y(_480_)
);

NAND3X1 _2764_ (
    .A(_474_),
    .B(_480_),
    .C(_460_),
    .Y(_481_)
);

NAND2X1 _2765_ (
    .A(_474_),
    .B(_460_),
    .Y(_482_)
);

OAI21X1 _2766_ (
    .A(_475_),
    .B(_479_),
    .C(_482_),
    .Y(_483_)
);

NAND3X1 _2767_ (
    .A(RDY_bF$buf1),
    .B(_481_),
    .C(_483_),
    .Y(_484_)
);

NAND2X1 _2768_ (
    .A(_853__bF$buf4),
    .B(_299_),
    .Y(_485_)
);

AND2X2 _2769_ (
    .A(_484_),
    .B(_485_),
    .Y(_16_)
);

AOI22X1 _2770_ (
    .A(AN),
    .B(_325_),
    .C(_338_),
    .D(ABH[7]),
    .Y(_486_)
);

NAND3X1 _2771_ (
    .A(_1051__bF$buf3),
    .B(_486_),
    .C(_1120_),
    .Y(_487_)
);

AOI21X1 _2772_ (
    .A(DIMUX[7]),
    .B(_446_),
    .C(_487_),
    .Y(_488_)
);

OAI21X1 _2773_ (
    .A(_303_),
    .B(_445_),
    .C(_488_),
    .Y(_489_)
);

INVX1 _2774_ (
    .A(_480_),
    .Y(_490_)
);

NAND3X1 _2775_ (
    .A(_474_),
    .B(_490_),
    .C(_460_),
    .Y(_491_)
);

XOR2X1 _2776_ (
    .A(_491_),
    .B(_489_),
    .Y(_492_)
);

NAND2X1 _2777_ (
    .A(PC[15]),
    .B(_853__bF$buf3),
    .Y(_493_)
);

OAI21X1 _2778_ (
    .A(_853__bF$buf2),
    .B(_492_),
    .C(_493_),
    .Y(_17_)
);

INVX1 _2779_ (
    .A(NMI_1),
    .Y(_494_)
);

NAND2X1 _2780_ (
    .A(NMI),
    .B(_494_),
    .Y(_495_)
);

OAI21X1 _2781_ (
    .A(_918__bF$buf2),
    .B(_961_),
    .C(NMI_edge),
    .Y(_496_)
);

OAI21X1 _2782_ (
    .A(NMI_edge),
    .B(_495_),
    .C(_496_),
    .Y(_18_)
);

INVX1 _2783_ (
    .A(cond_code[0]),
    .Y(_497_)
);

INVX2 _2784_ (
    .A(_1297_),
    .Y(_498_)
);

NAND2X1 _2785_ (
    .A(RDY_bF$buf0),
    .B(_498_),
    .Y(_499_)
);

OAI21X1 _2786_ (
    .A(RDY_bF$buf8),
    .B(_497_),
    .C(_499_),
    .Y(_19_)
);

NAND2X1 _2787_ (
    .A(cond_code[1]),
    .B(_853__bF$buf1),
    .Y(_500_)
);

OAI21X1 _2788_ (
    .A(_853__bF$buf0),
    .B(_1303_),
    .C(_500_),
    .Y(_20_)
);

NAND2X1 _2789_ (
    .A(cond_code[2]),
    .B(_853__bF$buf7),
    .Y(_501_)
);

OAI21X1 _2790_ (
    .A(_853__bF$buf6),
    .B(_1159_),
    .C(_501_),
    .Y(_21_)
);

INVX1 _2791_ (
    .A(plp),
    .Y(_502_)
);

OAI22X1 _2792_ (
    .A(_502_),
    .B(_1129__bF$buf4),
    .C(_1299_),
    .D(_1324_),
    .Y(_22_)
);

INVX1 _2793_ (
    .A(_1324_),
    .Y(_503_)
);

NAND2X1 _2794_ (
    .A(_1395_),
    .B(_503_),
    .Y(_504_)
);

OAI21X1 _2795_ (
    .A(_140_),
    .B(_1129__bF$buf3),
    .C(_504_),
    .Y(_23_)
);

OAI21X1 _2796_ (
    .A(_853__bF$buf5),
    .B(_1002__bF$buf4),
    .C(clc),
    .Y(_505_)
);

NAND2X1 _2797_ (
    .A(_1297_),
    .B(_1352_),
    .Y(_506_)
);

OR2X2 _2798_ (
    .A(_1215_),
    .B(_1394_),
    .Y(_507_)
);

OAI21X1 _2799_ (
    .A(_506_),
    .B(_507_),
    .C(_505_),
    .Y(_24_)
);

INVX1 _2800_ (
    .A(sec),
    .Y(_508_)
);

NOR2X1 _2801_ (
    .A(_1002__bF$buf3),
    .B(_499_),
    .Y(_509_)
);

NAND2X1 _2802_ (
    .A(_1220_),
    .B(_509_),
    .Y(_510_)
);

OAI22X1 _2803_ (
    .A(_508_),
    .B(_1129__bF$buf2),
    .C(_510_),
    .D(_507_),
    .Y(_25_)
);

OAI21X1 _2804_ (
    .A(_853__bF$buf4),
    .B(_1002__bF$buf2),
    .C(cld),
    .Y(_511_)
);

NOR2X1 _2805_ (
    .A(_1159_),
    .B(_1303_),
    .Y(_512_)
);

NAND2X1 _2806_ (
    .A(_512_),
    .B(_1323_),
    .Y(_513_)
);

OAI21X1 _2807_ (
    .A(_506_),
    .B(_513_),
    .C(_511_),
    .Y(_26_)
);

INVX1 _2808_ (
    .A(sed),
    .Y(_514_)
);

OAI22X1 _2809_ (
    .A(_514_),
    .B(_1129__bF$buf1),
    .C(_513_),
    .D(_510_),
    .Y(_27_)
);

INVX1 _2810_ (
    .A(cli),
    .Y(_515_)
);

INVX1 _2811_ (
    .A(_1163_),
    .Y(_516_)
);

NAND2X1 _2812_ (
    .A(_516_),
    .B(_1323_),
    .Y(_517_)
);

OAI22X1 _2813_ (
    .A(_515_),
    .B(_1129__bF$buf0),
    .C(_506_),
    .D(_517_),
    .Y(_28_)
);

OAI21X1 _2814_ (
    .A(_853__bF$buf3),
    .B(_1002__bF$buf1),
    .C(sei),
    .Y(_518_)
);

OAI21X1 _2815_ (
    .A(_517_),
    .B(_510_),
    .C(_518_),
    .Y(_29_)
);

OAI21X1 _2816_ (
    .A(_853__bF$buf2),
    .B(_1002__bF$buf0),
    .C(clv),
    .Y(_519_)
);

NOR2X1 _2817_ (
    .A(_1159_),
    .B(_1162_),
    .Y(_520_)
);

NAND2X1 _2818_ (
    .A(_498_),
    .B(_520_),
    .Y(_521_)
);

NOR2X1 _2819_ (
    .A(_1168_),
    .B(_521_),
    .Y(_522_)
);

INVX1 _2820_ (
    .A(_522_),
    .Y(_523_)
);

OAI21X1 _2821_ (
    .A(_1324_),
    .B(_523_),
    .C(_519_),
    .Y(_30_)
);

INVX1 _2822_ (
    .A(bit_ins),
    .Y(_524_)
);

NAND3X1 _2823_ (
    .A(_1314_),
    .B(_1296_),
    .C(_1298_),
    .Y(_525_)
);

NOR2X1 _2824_ (
    .A(_1139_),
    .B(_525_),
    .Y(_526_)
);

NOR2X1 _2825_ (
    .A(_1219__bF$buf0),
    .B(_526_),
    .Y(_527_)
);

AOI21X1 _2826_ (
    .A(_524_),
    .B(_1219__bF$buf3),
    .C(_527_),
    .Y(_31_)
);

NOR2X1 _2827_ (
    .A(_1178_),
    .B(_1304_),
    .Y(_528_)
);

AND2X2 _2828_ (
    .A(_528_),
    .B(_1175_),
    .Y(_529_)
);

INVX1 _2829_ (
    .A(_529_),
    .Y(_530_)
);

NOR2X1 _2830_ (
    .A(_1178_),
    .B(_1400_),
    .Y(_531_)
);

NOR2X1 _2831_ (
    .A(_531_),
    .B(_526_),
    .Y(_532_)
);

OAI21X1 _2832_ (
    .A(_1297_),
    .B(_530_),
    .C(_532_),
    .Y(_533_)
);

INVX1 _2833_ (
    .A(_533_),
    .Y(_534_)
);

INVX1 _2834_ (
    .A(_531_),
    .Y(_535_)
);

NOR2X1 _2835_ (
    .A(_529_),
    .B(_526_),
    .Y(_536_)
);

AOI21X1 _2836_ (
    .A(_536_),
    .B(_535_),
    .C(_1219__bF$buf2),
    .Y(_537_)
);

AOI22X1 _2837_ (
    .A(_118_),
    .B(_1219__bF$buf1),
    .C(_534_),
    .D(_537_),
    .Y(_32_)
);

NAND2X1 _2838_ (
    .A(_1297_),
    .B(_1162_),
    .Y(_538_)
);

NOR2X1 _2839_ (
    .A(_538_),
    .B(_1350_),
    .Y(_539_)
);

OAI21X1 _2840_ (
    .A(_1383_),
    .B(_539_),
    .C(_1159_),
    .Y(_540_)
);

AOI22X1 _2841_ (
    .A(_123_),
    .B(_1219__bF$buf0),
    .C(_537_),
    .D(_540_),
    .Y(_33_)
);

NAND2X1 _2842_ (
    .A(_1314_),
    .B(_1383_),
    .Y(_541_)
);

OAI21X1 _2843_ (
    .A(_498_),
    .B(_541_),
    .C(_1350_),
    .Y(_542_)
);

NAND2X1 _2844_ (
    .A(_512_),
    .B(_542_),
    .Y(_543_)
);

NAND2X1 _2845_ (
    .A(_1155_),
    .B(_512_),
    .Y(_544_)
);

OAI21X1 _2846_ (
    .A(_1384_),
    .B(_544_),
    .C(_543_),
    .Y(_545_)
);

NAND2X1 _2847_ (
    .A(_1297_),
    .B(_1178_),
    .Y(_546_)
);

NAND2X1 _2848_ (
    .A(_1168_),
    .B(_1323_),
    .Y(_547_)
);

NOR2X1 _2849_ (
    .A(_546_),
    .B(_547_),
    .Y(_548_)
);

INVX1 _2850_ (
    .A(_548_),
    .Y(_549_)
);

INVX1 _2851_ (
    .A(_512_),
    .Y(_550_)
);

NOR2X1 _2852_ (
    .A(_1220_),
    .B(_550_),
    .Y(_551_)
);

NAND2X1 _2853_ (
    .A(_1316_),
    .B(_551_),
    .Y(_552_)
);

NAND3X1 _2854_ (
    .A(_1142_),
    .B(_1168_),
    .C(_1214_),
    .Y(_553_)
);

OAI21X1 _2855_ (
    .A(_550_),
    .B(_553_),
    .C(_552_),
    .Y(_554_)
);

INVX1 _2856_ (
    .A(_554_),
    .Y(_555_)
);

OAI21X1 _2857_ (
    .A(_1162_),
    .B(_549_),
    .C(_555_),
    .Y(_556_)
);

NOR2X1 _2858_ (
    .A(_545_),
    .B(_556_),
    .Y(_557_)
);

AOI21X1 _2859_ (
    .A(_516_),
    .B(_1383_),
    .C(_1219__bF$buf3),
    .Y(_558_)
);

AND2X2 _2860_ (
    .A(_536_),
    .B(_558_),
    .Y(_559_)
);

AOI22X1 _2861_ (
    .A(_124_),
    .B(_1219__bF$buf2),
    .C(_557_),
    .D(_559_),
    .Y(_34_)
);

INVX1 _2862_ (
    .A(_537_),
    .Y(_560_)
);

OAI21X1 _2863_ (
    .A(_132_),
    .B(_1129__bF$buf4),
    .C(_560_),
    .Y(_35_)
);

OAI21X1 _2864_ (
    .A(_1171_),
    .B(_1314_),
    .C(_509_),
    .Y(_561_)
);

OAI22X1 _2865_ (
    .A(_908_),
    .B(_1129__bF$buf3),
    .C(_561_),
    .D(_535_),
    .Y(_36_)
);

AOI21X1 _2866_ (
    .A(_311_),
    .B(_1219__bF$buf1),
    .C(_558_),
    .Y(_37_)
);

AND2X2 _2867_ (
    .A(_539_),
    .B(_1178_),
    .Y(_562_)
);

OAI21X1 _2868_ (
    .A(_562_),
    .B(_554_),
    .C(_1129__bF$buf2),
    .Y(_563_)
);

OAI21X1 _2869_ (
    .A(_920_),
    .B(_1129__bF$buf1),
    .C(_563_),
    .Y(_38_)
);

NAND2X1 _2870_ (
    .A(_1129__bF$buf0),
    .B(_531_),
    .Y(_564_)
);

OAI22X1 _2871_ (
    .A(_912_),
    .B(_1129__bF$buf4),
    .C(_1329_),
    .D(_564_),
    .Y(_39_)
);

OAI21X1 _2872_ (
    .A(_1008_),
    .B(_1036_),
    .C(RDY_bF$buf7),
    .Y(_565_)
);

INVX1 _2873_ (
    .A(_565_),
    .Y(_566_)
);

NAND2X1 _2874_ (
    .A(D),
    .B(_1159_),
    .Y(_567_)
);

NAND3X1 _2875_ (
    .A(_1304_),
    .B(_566_),
    .C(_1175_),
    .Y(_568_)
);

OAI22X1 _2876_ (
    .A(_310_),
    .B(_566_),
    .C(_567_),
    .D(_568_),
    .Y(_40_)
);

INVX1 _2877_ (
    .A(adc_sbc),
    .Y(_569_)
);

OAI21X1 _2878_ (
    .A(_569_),
    .B(_566_),
    .C(_568_),
    .Y(_41_)
);

OAI21X1 _2879_ (
    .A(_853__bF$buf1),
    .B(_1002__bF$buf4),
    .C(inc),
    .Y(_570_)
);

NOR2X1 _2880_ (
    .A(_550_),
    .B(_541_),
    .Y(_571_)
);

AOI22X1 _2881_ (
    .A(_1323_),
    .B(_551_),
    .C(_571_),
    .D(_498_),
    .Y(_572_)
);

OAI21X1 _2882_ (
    .A(_1219__bF$buf0),
    .B(_572_),
    .C(_570_),
    .Y(_42_)
);

OAI21X1 _2883_ (
    .A(_853__bF$buf0),
    .B(_1002__bF$buf3),
    .C(load_only),
    .Y(_573_)
);

OAI21X1 _2884_ (
    .A(_1219__bF$buf3),
    .B(_521_),
    .C(_573_),
    .Y(_43_)
);

OR2X2 _2885_ (
    .A(_541_),
    .B(_1219__bF$buf2),
    .Y(_574_)
);

OAI22X1 _2886_ (
    .A(_1250_),
    .B(_1129__bF$buf3),
    .C(_520_),
    .D(_574_),
    .Y(_44_)
);

NAND2X1 _2887_ (
    .A(_1129__bF$buf2),
    .B(_1178_),
    .Y(_575_)
);

OAI21X1 _2888_ (
    .A(_853__bF$buf7),
    .B(_1002__bF$buf2),
    .C(store),
    .Y(_576_)
);

OAI21X1 _2889_ (
    .A(_1154_),
    .B(_1161_),
    .C(_1145_),
    .Y(_577_)
);

NOR2X1 _2890_ (
    .A(_1148_),
    .B(_1382_),
    .Y(_578_)
);

OAI21X1 _2891_ (
    .A(_1175_),
    .B(_578_),
    .C(_577_),
    .Y(_579_)
);

OAI21X1 _2892_ (
    .A(_575_),
    .B(_579_),
    .C(_576_),
    .Y(_45_)
);

INVX1 _2893_ (
    .A(index_y),
    .Y(_580_)
);

NAND2X1 _2894_ (
    .A(_1220_),
    .B(_520_),
    .Y(_581_)
);

NOR2X1 _2895_ (
    .A(_541_),
    .B(_581_),
    .Y(_582_)
);

OAI21X1 _2896_ (
    .A(_1168_),
    .B(_1330_),
    .C(_1176_),
    .Y(_583_)
);

OAI21X1 _2897_ (
    .A(_583_),
    .B(_582_),
    .C(_1129__bF$buf1),
    .Y(_584_)
);

OAI21X1 _2898_ (
    .A(_580_),
    .B(_1129__bF$buf0),
    .C(_584_),
    .Y(_46_)
);

NAND2X1 _2899_ (
    .A(_1303_),
    .B(_1314_),
    .Y(_585_)
);

OAI21X1 _2900_ (
    .A(_546_),
    .B(_585_),
    .C(_544_),
    .Y(_586_)
);

OR2X2 _2901_ (
    .A(_581_),
    .B(_498_),
    .Y(_587_)
);

OAI21X1 _2902_ (
    .A(_1215_),
    .B(_587_),
    .C(_549_),
    .Y(_588_)
);

AOI21X1 _2903_ (
    .A(_1214_),
    .B(_586_),
    .C(_588_),
    .Y(_589_)
);

OAI21X1 _2904_ (
    .A(_1384_),
    .B(_523_),
    .C(_589_),
    .Y(_590_)
);

INVX1 _2905_ (
    .A(_590_),
    .Y(_591_)
);

OAI21X1 _2906_ (
    .A(_853__bF$buf6),
    .B(_1002__bF$buf1),
    .C(src_reg[0]),
    .Y(_592_)
);

OAI21X1 _2907_ (
    .A(_1219__bF$buf1),
    .B(_591_),
    .C(_592_),
    .Y(_47_)
);

OAI21X1 _2908_ (
    .A(_544_),
    .B(_1384_),
    .C(_1129__bF$buf4),
    .Y(_593_)
);

NAND3X1 _2909_ (
    .A(_1214_),
    .B(_498_),
    .C(_551_),
    .Y(_594_)
);

NAND3X1 _2910_ (
    .A(_1149_),
    .B(_1297_),
    .C(_520_),
    .Y(_595_)
);

OAI21X1 _2911_ (
    .A(_1400_),
    .B(_595_),
    .C(_594_),
    .Y(_596_)
);

NOR2X1 _2912_ (
    .A(_593_),
    .B(_596_),
    .Y(_597_)
);

AOI22X1 _2913_ (
    .A(_1014_),
    .B(_1219__bF$buf0),
    .C(_589_),
    .D(_597_),
    .Y(_48_)
);

INVX1 _2914_ (
    .A(dst_reg[0]),
    .Y(_598_)
);

OAI21X1 _2915_ (
    .A(_1314_),
    .B(_1168_),
    .C(_1214_),
    .Y(_599_)
);

OAI21X1 _2916_ (
    .A(_521_),
    .B(_599_),
    .C(_549_),
    .Y(_600_)
);

OAI21X1 _2917_ (
    .A(_1384_),
    .B(_587_),
    .C(_1438_),
    .Y(_601_)
);

NOR2X1 _2918_ (
    .A(_600_),
    .B(_601_),
    .Y(_602_)
);

AOI21X1 _2919_ (
    .A(_598_),
    .B(_1219__bF$buf3),
    .C(_602_),
    .Y(_49_)
);

INVX1 _2920_ (
    .A(_521_),
    .Y(_603_)
);

AOI21X1 _2921_ (
    .A(_1383_),
    .B(_603_),
    .C(_593_),
    .Y(_604_)
);

OAI21X1 _2922_ (
    .A(_1172_),
    .B(_594_),
    .C(_604_),
    .Y(_605_)
);

NOR2X1 _2923_ (
    .A(_600_),
    .B(_605_),
    .Y(_606_)
);

AOI21X1 _2924_ (
    .A(_1001_),
    .B(_1219__bF$buf2),
    .C(_606_),
    .Y(_50_)
);

INVX1 _2925_ (
    .A(load_reg),
    .Y(_607_)
);

OAI21X1 _2926_ (
    .A(_1384_),
    .B(_523_),
    .C(_547_),
    .Y(_608_)
);

NAND2X1 _2927_ (
    .A(_578_),
    .B(_522_),
    .Y(_609_)
);

OAI21X1 _2928_ (
    .A(_1320_),
    .B(_1384_),
    .C(_609_),
    .Y(_610_)
);

NOR2X1 _2929_ (
    .A(_610_),
    .B(_608_),
    .Y(_611_)
);

NOR2X1 _2930_ (
    .A(_1382_),
    .B(_498_),
    .Y(_612_)
);

NAND3X1 _2931_ (
    .A(_1173_),
    .B(_520_),
    .C(_612_),
    .Y(_613_)
);

NAND3X1 _2932_ (
    .A(_1138_),
    .B(_1168_),
    .C(_603_),
    .Y(_614_)
);

OAI21X1 _2933_ (
    .A(_498_),
    .B(_1159_),
    .C(_1175_),
    .Y(_615_)
);

NAND3X1 _2934_ (
    .A(_613_),
    .B(_615_),
    .C(_614_),
    .Y(_616_)
);

NOR2X1 _2935_ (
    .A(_593_),
    .B(_616_),
    .Y(_617_)
);

AOI22X1 _2936_ (
    .A(_607_),
    .B(_1219__bF$buf1),
    .C(_611_),
    .D(_617_),
    .Y(_51_)
);

AND2X2 _2937_ (
    .A(_1002__bF$buf0),
    .B(res),
    .Y(_52_)
);

OAI21X1 _2938_ (
    .A(_1043_),
    .B(_1044_),
    .C(RDY_bF$buf6),
    .Y(_618_)
);

NOR2X1 _2939_ (
    .A(reset),
    .B(_618_),
    .Y(_619_)
);

INVX2 _2940_ (
    .A(_619_),
    .Y(_620_)
);

OAI21X1 _2941_ (
    .A(reset),
    .B(_618_),
    .C(IRHOLD[0]),
    .Y(_621_)
);

OAI21X1 _2942_ (
    .A(_932_),
    .B(_620_),
    .C(_621_),
    .Y(_53_)
);

OAI21X1 _2943_ (
    .A(reset),
    .B(_618_),
    .C(IRHOLD[1]),
    .Y(_622_)
);

OAI21X1 _2944_ (
    .A(_969_),
    .B(_620_),
    .C(_622_),
    .Y(_54_)
);

OAI21X1 _2945_ (
    .A(reset),
    .B(_618_),
    .C(IRHOLD[2]),
    .Y(_623_)
);

OAI21X1 _2946_ (
    .A(_855_),
    .B(_620_),
    .C(_623_),
    .Y(_55_)
);

OAI21X1 _2947_ (
    .A(reset),
    .B(_618_),
    .C(IRHOLD[3]),
    .Y(_624_)
);

OAI21X1 _2948_ (
    .A(_857_),
    .B(_620_),
    .C(_624_),
    .Y(_56_)
);

OAI21X1 _2949_ (
    .A(reset),
    .B(_618_),
    .C(IRHOLD[4]),
    .Y(_625_)
);

OAI21X1 _2950_ (
    .A(_859_),
    .B(_620_),
    .C(_625_),
    .Y(_57_)
);

OAI21X1 _2951_ (
    .A(reset),
    .B(_618_),
    .C(IRHOLD[5]),
    .Y(_626_)
);

OAI21X1 _2952_ (
    .A(_861_),
    .B(_620_),
    .C(_626_),
    .Y(_58_)
);

OAI21X1 _2953_ (
    .A(reset),
    .B(_618_),
    .C(IRHOLD[6]),
    .Y(_627_)
);

OAI21X1 _2954_ (
    .A(_863_),
    .B(_620_),
    .C(_627_),
    .Y(_59_)
);

OAI21X1 _2955_ (
    .A(reset),
    .B(_618_),
    .C(IRHOLD[7]),
    .Y(_628_)
);

OAI21X1 _2956_ (
    .A(_864_),
    .B(_620_),
    .C(_628_),
    .Y(_60_)
);

OAI21X1 _2957_ (
    .A(_1169_),
    .B(_1129__bF$buf3),
    .C(_618_),
    .Y(_61_)
);

OAI21X1 _2958_ (
    .A(_887__bF$buf0),
    .B(_1259_),
    .C(_1002__bF$buf4),
    .Y(_629_)
);

INVX1 _2959_ (
    .A(_629_),
    .Y(_630_)
);

OAI21X1 _2960_ (
    .A(_524_),
    .B(_1031_),
    .C(_630_),
    .Y(_631_)
);

NOR2X1 _2961_ (
    .A(plp),
    .B(_1002__bF$buf3),
    .Y(_632_)
);

INVX1 _2962_ (
    .A(_632_),
    .Y(_633_)
);

NOR2X1 _2963_ (
    .A(clv),
    .B(_633_),
    .Y(_634_)
);

INVX1 _2964_ (
    .A(_634_),
    .Y(_635_)
);

OAI21X1 _2965_ (
    .A(adc_sbc),
    .B(_635_),
    .C(_631_),
    .Y(_636_)
);

OAI21X1 _2966_ (
    .A(_918__bF$buf1),
    .B(_988_),
    .C(DIMUX[6]),
    .Y(_637_)
);

NAND2X1 _2967_ (
    .A(plp),
    .B(ADD[6]),
    .Y(_638_)
);

OAI21X1 _2968_ (
    .A(_1002__bF$buf2),
    .B(_638_),
    .C(_637_),
    .Y(_639_)
);

AOI21X1 _2969_ (
    .A(_634_),
    .B(AV),
    .C(_639_),
    .Y(_640_)
);

NAND2X1 _2970_ (
    .A(V),
    .B(_636_),
    .Y(_641_)
);

OAI21X1 _2971_ (
    .A(_636_),
    .B(_640_),
    .C(_641_),
    .Y(_62_)
);

NOR2X1 _2972_ (
    .A(plp),
    .B(cld),
    .Y(_642_)
);

NAND2X1 _2973_ (
    .A(_514_),
    .B(_642_),
    .Y(_643_)
);

OAI21X1 _2974_ (
    .A(_1002__bF$buf1),
    .B(_643_),
    .C(_629_),
    .Y(_644_)
);

NAND2X1 _2975_ (
    .A(D),
    .B(_644_),
    .Y(_645_)
);

NAND2X1 _2976_ (
    .A(plp),
    .B(ADD[3]),
    .Y(_646_)
);

OAI21X1 _2977_ (
    .A(plp),
    .B(cld),
    .C(_646_),
    .Y(_647_)
);

MUX2X1 _2978_ (
    .A(DIMUX[3]),
    .B(_647_),
    .S(_1260_),
    .Y(_648_)
);

OAI21X1 _2979_ (
    .A(_644_),
    .B(_648_),
    .C(_645_),
    .Y(_63_)
);

NAND2X1 _2980_ (
    .A(_515_),
    .B(_951_),
    .Y(_649_)
);

AOI21X1 _2981_ (
    .A(_630_),
    .B(_978_),
    .C(_632_),
    .Y(_650_)
);

OAI22X1 _2982_ (
    .A(sei),
    .B(_649_),
    .C(_951_),
    .D(_650_),
    .Y(_651_)
);

INVX1 _2983_ (
    .A(_1260_),
    .Y(_652_)
);

OAI21X1 _2984_ (
    .A(_437_),
    .B(_951_),
    .C(_649_),
    .Y(_653_)
);

OAI21X1 _2985_ (
    .A(_855_),
    .B(_652_),
    .C(_978_),
    .Y(_654_)
);

AOI21X1 _2986_ (
    .A(_653_),
    .B(_652_),
    .C(_654_),
    .Y(_655_)
);

NAND2X1 _2987_ (
    .A(I),
    .B(_651_),
    .Y(_656_)
);

OAI21X1 _2988_ (
    .A(_651_),
    .B(_655_),
    .C(_656_),
    .Y(_64_)
);

NOR2X1 _2989_ (
    .A(compare),
    .B(_633_),
    .Y(_657_)
);

OAI21X1 _2990_ (
    .A(_607_),
    .B(_1022_),
    .C(_657_),
    .Y(_658_)
);

OAI21X1 _2991_ (
    .A(_1191_),
    .B(_631_),
    .C(_658_),
    .Y(_659_)
);

OAI21X1 _2992_ (
    .A(_502_),
    .B(AN),
    .C(_1008_),
    .Y(_660_)
);

OAI21X1 _2993_ (
    .A(_864_),
    .B(_1008_),
    .C(_660_),
    .Y(_661_)
);

INVX1 _2994_ (
    .A(AN),
    .Y(_662_)
);

OAI21X1 _2995_ (
    .A(_632_),
    .B(_1191_),
    .C(_662_),
    .Y(_663_)
);

OAI21X1 _2996_ (
    .A(_1191_),
    .B(_661_),
    .C(_663_),
    .Y(_664_)
);

NAND2X1 _2997_ (
    .A(N),
    .B(_659_),
    .Y(_665_)
);

OAI21X1 _2998_ (
    .A(_659_),
    .B(_664_),
    .C(_665_),
    .Y(_65_)
);

OAI22X1 _2999_ (
    .A(_1191_),
    .B(_629_),
    .C(bit_ins),
    .D(_658_),
    .Y(_666_)
);

MUX2X1 _3000_ (
    .A(ADD[1]),
    .B(AZ),
    .S(plp),
    .Y(_667_)
);

NAND2X1 _3001_ (
    .A(DIMUX[1]),
    .B(_1260_),
    .Y(_668_)
);

OAI21X1 _3002_ (
    .A(_1260_),
    .B(_667_),
    .C(_668_),
    .Y(_669_)
);

MUX2X1 _3003_ (
    .A(_669_),
    .B(AZ),
    .S(_1192_),
    .Y(_670_)
);

NAND2X1 _3004_ (
    .A(Z),
    .B(_666_),
    .Y(_671_)
);

OAI21X1 _3005_ (
    .A(_666_),
    .B(_670_),
    .C(_671_),
    .Y(_66_)
);

NOR2X1 _3006_ (
    .A(write_back),
    .B(_1002__bF$buf0),
    .Y(_672_)
);

NAND3X1 _3007_ (
    .A(_569_),
    .B(_912_),
    .C(_920_),
    .Y(_673_)
);

NOR2X1 _3008_ (
    .A(plp),
    .B(clc),
    .Y(_674_)
);

NAND2X1 _3009_ (
    .A(_508_),
    .B(_674_),
    .Y(_675_)
);

OAI21X1 _3010_ (
    .A(_673_),
    .B(_675_),
    .C(_672_),
    .Y(_676_)
);

AOI21X1 _3011_ (
    .A(shift),
    .B(_1191_),
    .C(_1260_),
    .Y(_677_)
);

AND2X2 _3012_ (
    .A(_677_),
    .B(_676_),
    .Y(_678_)
);

AOI21X1 _3013_ (
    .A(plp),
    .B(ADD[0]),
    .C(_674_),
    .Y(_679_)
);

NAND2X1 _3014_ (
    .A(CO),
    .B(_673_),
    .Y(_680_)
);

OAI21X1 _3015_ (
    .A(_673_),
    .B(_679_),
    .C(_680_),
    .Y(_681_)
);

NAND2X1 _3016_ (
    .A(_932_),
    .B(_1260_),
    .Y(_682_)
);

OAI21X1 _3017_ (
    .A(_1260_),
    .B(_681_),
    .C(_682_),
    .Y(_683_)
);

NAND2X1 _3018_ (
    .A(C),
    .B(_678_),
    .Y(_684_)
);

OAI21X1 _3019_ (
    .A(_678_),
    .B(_683_),
    .C(_684_),
    .Y(_67_)
);

INVX1 _3020_ (
    .A(backwards),
    .Y(_685_)
);

NAND2X1 _3021_ (
    .A(RDY_bF$buf5),
    .B(DI[7]),
    .Y(_686_)
);

OAI21X1 _3022_ (
    .A(RDY_bF$buf4),
    .B(_685_),
    .C(_686_),
    .Y(_68_)
);

NOR2X1 _3023_ (
    .A(_607_),
    .B(_633_),
    .Y(_687_)
);

OAI21X1 _3024_ (
    .A(_887__bF$buf4),
    .B(_1035_),
    .C(_981_),
    .Y(_688_)
);

NOR2X1 _3025_ (
    .A(_979_),
    .B(_688_),
    .Y(_689_)
);

INVX1 _3026_ (
    .A(_689_),
    .Y(_690_)
);

OAI21X1 _3027_ (
    .A(_687_),
    .B(_690_),
    .C(RDY_bF$buf3),
    .Y(_691_)
);

INVX1 _3028_ (
    .A(_691__bF$buf3),
    .Y(_692_)
);

NAND2X1 _3029_ (
    .A(_692_),
    .B(_1020_),
    .Y(_693_)
);

OAI21X1 _3030_ (
    .A(_917_),
    .B(_949_),
    .C(_263_),
    .Y(_694_)
);

OAI21X1 _3031_ (
    .A(DIMUX[0]),
    .B(_981_),
    .C(_694_),
    .Y(_695_)
);

NAND2X1 _3032_ (
    .A(\AXYS[0] [0]),
    .B(_693_),
    .Y(_696_)
);

OAI21X1 _3033_ (
    .A(_693_),
    .B(_695_),
    .C(_696_),
    .Y(_69_)
);

NAND3X1 _3034_ (
    .A(adj_bcd),
    .B(adc_bcd),
    .C(HC),
    .Y(_697_)
);

NAND2X1 _3035_ (
    .A(adj_bcd),
    .B(_310_),
    .Y(_698_)
);

OAI21X1 _3036_ (
    .A(HC),
    .B(_698_),
    .C(_697_),
    .Y(_699_)
);

INVX1 _3037_ (
    .A(_697_),
    .Y(_700_)
);

NOR2X1 _3038_ (
    .A(HC),
    .B(_698_),
    .Y(_701_)
);

OAI21X1 _3039_ (
    .A(_700_),
    .B(_701_),
    .C(ADD[1]),
    .Y(_702_)
);

INVX1 _3040_ (
    .A(_702_),
    .Y(_703_)
);

NOR2X1 _3041_ (
    .A(_1281_),
    .B(_703_),
    .Y(_704_)
);

OAI21X1 _3042_ (
    .A(ADD[1]),
    .B(_699_),
    .C(_704_),
    .Y(_705_)
);

OAI21X1 _3043_ (
    .A(_969_),
    .B(_981_),
    .C(_705_),
    .Y(_706_)
);

INVX1 _3044_ (
    .A(_706_),
    .Y(_707_)
);

NAND2X1 _3045_ (
    .A(\AXYS[0] [1]),
    .B(_693_),
    .Y(_708_)
);

OAI21X1 _3046_ (
    .A(_693_),
    .B(_707_),
    .C(_708_),
    .Y(_70_)
);

XNOR2X1 _3047_ (
    .A(_697_),
    .B(ADD[2]),
    .Y(_709_)
);

INVX1 _3048_ (
    .A(_709_),
    .Y(_710_)
);

NAND2X1 _3049_ (
    .A(_710_),
    .B(_702_),
    .Y(_711_)
);

NOR2X1 _3050_ (
    .A(_710_),
    .B(_702_),
    .Y(_712_)
);

NOR2X1 _3051_ (
    .A(_1281_),
    .B(_712_),
    .Y(_713_)
);

AOI22X1 _3052_ (
    .A(DIMUX[2]),
    .B(_1281_),
    .C(_713_),
    .D(_711_),
    .Y(_714_)
);

NAND2X1 _3053_ (
    .A(\AXYS[0] [2]),
    .B(_693_),
    .Y(_715_)
);

OAI21X1 _3054_ (
    .A(_693_),
    .B(_714_),
    .C(_715_),
    .Y(_71_)
);

INVX1 _3055_ (
    .A(_712_),
    .Y(_716_)
);

OAI21X1 _3056_ (
    .A(_437_),
    .B(_697_),
    .C(_716_),
    .Y(_717_)
);

XNOR2X1 _3057_ (
    .A(_701_),
    .B(ADD[3]),
    .Y(_718_)
);

AND2X2 _3058_ (
    .A(_717_),
    .B(_718_),
    .Y(_719_)
);

OAI21X1 _3059_ (
    .A(_718_),
    .B(_717_),
    .C(_981_),
    .Y(_720_)
);

OAI22X1 _3060_ (
    .A(DIMUX[3]),
    .B(_981_),
    .C(_720_),
    .D(_719_),
    .Y(_721_)
);

NAND2X1 _3061_ (
    .A(\AXYS[0] [3]),
    .B(_693_),
    .Y(_722_)
);

OAI21X1 _3062_ (
    .A(_693_),
    .B(_721_),
    .C(_722_),
    .Y(_72_)
);

OAI21X1 _3063_ (
    .A(_917_),
    .B(_949_),
    .C(_285_),
    .Y(_723_)
);

OAI21X1 _3064_ (
    .A(DIMUX[4]),
    .B(_981_),
    .C(_723_),
    .Y(_724_)
);

NAND2X1 _3065_ (
    .A(\AXYS[0] [4]),
    .B(_693_),
    .Y(_725_)
);

OAI21X1 _3066_ (
    .A(_693_),
    .B(_724_),
    .C(_725_),
    .Y(_73_)
);

NAND3X1 _3067_ (
    .A(adj_bcd),
    .B(adc_bcd),
    .C(CO),
    .Y(_726_)
);

OAI21X1 _3068_ (
    .A(CO),
    .B(_698_),
    .C(_726_),
    .Y(_727_)
);

INVX1 _3069_ (
    .A(_727_),
    .Y(_728_)
);

NAND2X1 _3070_ (
    .A(_293_),
    .B(_728_),
    .Y(_729_)
);

NOR2X1 _3071_ (
    .A(_293_),
    .B(_728_),
    .Y(_730_)
);

NOR2X1 _3072_ (
    .A(_1281_),
    .B(_730_),
    .Y(_731_)
);

AOI22X1 _3073_ (
    .A(DIMUX[5]),
    .B(_1281_),
    .C(_731_),
    .D(_729_),
    .Y(_732_)
);

NAND2X1 _3074_ (
    .A(\AXYS[0] [5]),
    .B(_693_),
    .Y(_733_)
);

OAI21X1 _3075_ (
    .A(_693_),
    .B(_732_),
    .C(_733_),
    .Y(_74_)
);

XNOR2X1 _3076_ (
    .A(_726_),
    .B(ADD[6]),
    .Y(_734_)
);

AOI21X1 _3077_ (
    .A(_730_),
    .B(_734_),
    .C(_1281_),
    .Y(_735_)
);

OAI21X1 _3078_ (
    .A(_730_),
    .B(_734_),
    .C(_735_),
    .Y(_736_)
);

OAI21X1 _3079_ (
    .A(_863_),
    .B(_981_),
    .C(_736_),
    .Y(_737_)
);

INVX1 _3080_ (
    .A(_737_),
    .Y(_738_)
);

NAND2X1 _3081_ (
    .A(\AXYS[0] [6]),
    .B(_693_),
    .Y(_739_)
);

OAI21X1 _3082_ (
    .A(_693_),
    .B(_738_),
    .C(_739_),
    .Y(_75_)
);

NAND2X1 _3083_ (
    .A(_734_),
    .B(_730_),
    .Y(_740_)
);

OAI21X1 _3084_ (
    .A(_246_),
    .B(_726_),
    .C(_740_),
    .Y(_741_)
);

NOR2X1 _3085_ (
    .A(CO),
    .B(_698_),
    .Y(_742_)
);

XOR2X1 _3086_ (
    .A(_742_),
    .B(AN),
    .Y(_743_)
);

XOR2X1 _3087_ (
    .A(_741_),
    .B(_743_),
    .Y(_744_)
);

MUX2X1 _3088_ (
    .A(_744_),
    .B(DIMUX[7]),
    .S(_981_),
    .Y(_745_)
);

NAND2X1 _3089_ (
    .A(\AXYS[0] [7]),
    .B(_693_),
    .Y(_746_)
);

OAI21X1 _3090_ (
    .A(_693_),
    .B(_745_),
    .C(_746_),
    .Y(_76_)
);

NAND2X1 _3091_ (
    .A(_692_),
    .B(_1022_),
    .Y(_747_)
);

INVX2 _3092_ (
    .A(_1022_),
    .Y(_748_)
);

OAI21X1 _3093_ (
    .A(_691__bF$buf2),
    .B(_748_),
    .C(\AXYS[1] [0]),
    .Y(_749_)
);

OAI21X1 _3094_ (
    .A(_695_),
    .B(_747_),
    .C(_749_),
    .Y(_77_)
);

OAI21X1 _3095_ (
    .A(_691__bF$buf1),
    .B(_748_),
    .C(\AXYS[1] [1]),
    .Y(_750_)
);

OAI21X1 _3096_ (
    .A(_707_),
    .B(_747_),
    .C(_750_),
    .Y(_78_)
);

OAI21X1 _3097_ (
    .A(_691__bF$buf0),
    .B(_748_),
    .C(\AXYS[1] [2]),
    .Y(_751_)
);

OAI21X1 _3098_ (
    .A(_714_),
    .B(_747_),
    .C(_751_),
    .Y(_79_)
);

OAI21X1 _3099_ (
    .A(_691__bF$buf3),
    .B(_748_),
    .C(\AXYS[1] [3]),
    .Y(_752_)
);

OAI21X1 _3100_ (
    .A(_721_),
    .B(_747_),
    .C(_752_),
    .Y(_80_)
);

OAI21X1 _3101_ (
    .A(_691__bF$buf2),
    .B(_748_),
    .C(\AXYS[1] [4]),
    .Y(_753_)
);

OAI21X1 _3102_ (
    .A(_724_),
    .B(_747_),
    .C(_753_),
    .Y(_81_)
);

OAI21X1 _3103_ (
    .A(_691__bF$buf1),
    .B(_748_),
    .C(\AXYS[1] [5]),
    .Y(_754_)
);

OAI21X1 _3104_ (
    .A(_732_),
    .B(_747_),
    .C(_754_),
    .Y(_82_)
);

OAI21X1 _3105_ (
    .A(_691__bF$buf0),
    .B(_748_),
    .C(\AXYS[1] [6]),
    .Y(_755_)
);

OAI21X1 _3106_ (
    .A(_738_),
    .B(_747_),
    .C(_755_),
    .Y(_83_)
);

OAI21X1 _3107_ (
    .A(_691__bF$buf3),
    .B(_748_),
    .C(\AXYS[1] [7]),
    .Y(_756_)
);

OAI21X1 _3108_ (
    .A(_745_),
    .B(_747_),
    .C(_756_),
    .Y(_84_)
);

NAND2X1 _3109_ (
    .A(_692_),
    .B(_1023_),
    .Y(_757_)
);

INVX2 _3110_ (
    .A(_1023_),
    .Y(_758_)
);

OAI21X1 _3111_ (
    .A(_691__bF$buf2),
    .B(_758_),
    .C(\AXYS[2] [0]),
    .Y(_759_)
);

OAI21X1 _3112_ (
    .A(_695_),
    .B(_757_),
    .C(_759_),
    .Y(_85_)
);

OAI21X1 _3113_ (
    .A(_691__bF$buf1),
    .B(_758_),
    .C(\AXYS[2] [1]),
    .Y(_760_)
);

OAI21X1 _3114_ (
    .A(_707_),
    .B(_757_),
    .C(_760_),
    .Y(_86_)
);

OAI21X1 _3115_ (
    .A(_691__bF$buf0),
    .B(_758_),
    .C(\AXYS[2] [2]),
    .Y(_761_)
);

OAI21X1 _3116_ (
    .A(_714_),
    .B(_757_),
    .C(_761_),
    .Y(_87_)
);

OAI21X1 _3117_ (
    .A(_691__bF$buf3),
    .B(_758_),
    .C(\AXYS[2] [3]),
    .Y(_762_)
);

OAI21X1 _3118_ (
    .A(_721_),
    .B(_757_),
    .C(_762_),
    .Y(_88_)
);

OAI21X1 _3119_ (
    .A(_691__bF$buf2),
    .B(_758_),
    .C(\AXYS[2] [4]),
    .Y(_763_)
);

OAI21X1 _3120_ (
    .A(_724_),
    .B(_757_),
    .C(_763_),
    .Y(_89_)
);

OAI21X1 _3121_ (
    .A(_691__bF$buf1),
    .B(_758_),
    .C(\AXYS[2] [5]),
    .Y(_764_)
);

OAI21X1 _3122_ (
    .A(_732_),
    .B(_757_),
    .C(_764_),
    .Y(_90_)
);

OAI21X1 _3123_ (
    .A(_691__bF$buf0),
    .B(_758_),
    .C(\AXYS[2] [6]),
    .Y(_765_)
);

OAI21X1 _3124_ (
    .A(_738_),
    .B(_757_),
    .C(_765_),
    .Y(_91_)
);

OAI21X1 _3125_ (
    .A(_691__bF$buf3),
    .B(_758_),
    .C(\AXYS[2] [7]),
    .Y(_766_)
);

OAI21X1 _3126_ (
    .A(_745_),
    .B(_757_),
    .C(_766_),
    .Y(_92_)
);

NAND2X1 _3127_ (
    .A(_692_),
    .B(_1012_),
    .Y(_767_)
);

NAND2X1 _3128_ (
    .A(\AXYS[3] [0]),
    .B(_767_),
    .Y(_768_)
);

OAI21X1 _3129_ (
    .A(_695_),
    .B(_767_),
    .C(_768_),
    .Y(_93_)
);

NAND2X1 _3130_ (
    .A(\AXYS[3] [1]),
    .B(_767_),
    .Y(_769_)
);

OAI21X1 _3131_ (
    .A(_707_),
    .B(_767_),
    .C(_769_),
    .Y(_94_)
);

NAND2X1 _3132_ (
    .A(\AXYS[3] [2]),
    .B(_767_),
    .Y(_770_)
);

OAI21X1 _3133_ (
    .A(_714_),
    .B(_767_),
    .C(_770_),
    .Y(_95_)
);

NAND2X1 _3134_ (
    .A(\AXYS[3] [3]),
    .B(_767_),
    .Y(_771_)
);

OAI21X1 _3135_ (
    .A(_721_),
    .B(_767_),
    .C(_771_),
    .Y(_96_)
);

NAND2X1 _3136_ (
    .A(\AXYS[3] [4]),
    .B(_767_),
    .Y(_772_)
);

OAI21X1 _3137_ (
    .A(_724_),
    .B(_767_),
    .C(_772_),
    .Y(_97_)
);

NAND2X1 _3138_ (
    .A(\AXYS[3] [5]),
    .B(_767_),
    .Y(_773_)
);

OAI21X1 _3139_ (
    .A(_732_),
    .B(_767_),
    .C(_773_),
    .Y(_98_)
);

NAND2X1 _3140_ (
    .A(\AXYS[3] [6]),
    .B(_767_),
    .Y(_774_)
);

OAI21X1 _3141_ (
    .A(_738_),
    .B(_767_),
    .C(_774_),
    .Y(_99_)
);

NAND2X1 _3142_ (
    .A(\AXYS[3] [7]),
    .B(_767_),
    .Y(_775_)
);

OAI21X1 _3143_ (
    .A(_745_),
    .B(_767_),
    .C(_775_),
    .Y(_100_)
);

AOI21X1 _3144_ (
    .A(_910_),
    .B(_869__bF$buf2),
    .C(_1224_),
    .Y(_776_)
);

OAI21X1 _3145_ (
    .A(state[4]),
    .B(_1035_),
    .C(_776_),
    .Y(_777_)
);

NOR2X1 _3146_ (
    .A(_1037_),
    .B(_777_),
    .Y(_778_)
);

OAI21X1 _3147_ (
    .A(_882__bF$buf0),
    .B(_880_),
    .C(_1002__bF$buf4),
    .Y(_779_)
);

NOR2X1 _3148_ (
    .A(_779_),
    .B(_951_),
    .Y(_780_)
);

OAI21X1 _3149_ (
    .A(_881_),
    .B(_917_),
    .C(_927_),
    .Y(_781_)
);

NAND3X1 _3150_ (
    .A(_781_),
    .B(_780_),
    .C(_778_),
    .Y(_782_)
);

OAI21X1 _3151_ (
    .A(_890_),
    .B(_1327_),
    .C(_994_),
    .Y(_783_)
);

OAI21X1 _3152_ (
    .A(_881_),
    .B(_917_),
    .C(_893_),
    .Y(_784_)
);

NAND3X1 _3153_ (
    .A(_976_),
    .B(_784_),
    .C(_783_),
    .Y(_785_)
);

NOR2X1 _3154_ (
    .A(_785_),
    .B(_782_),
    .Y(_786_)
);

INVX1 _3155_ (
    .A(_786_),
    .Y(_787_)
);

OAI21X1 _3156_ (
    .A(_917_),
    .B(_936_),
    .C(_1184_),
    .Y(_788_)
);

AOI21X1 _3157_ (
    .A(_869__bF$buf1),
    .B(_906_),
    .C(_1044_),
    .Y(_789_)
);

NAND3X1 _3158_ (
    .A(_1049_),
    .B(_990_),
    .C(_789_),
    .Y(_790_)
);

NOR2X1 _3159_ (
    .A(_788_),
    .B(_790_),
    .Y(_791_)
);

OAI21X1 _3160_ (
    .A(_886__bF$buf2),
    .B(_926__bF$buf1),
    .C(_900_),
    .Y(_792_)
);

OAI21X1 _3161_ (
    .A(state[4]),
    .B(_941_),
    .C(_792_),
    .Y(_793_)
);

INVX1 _3162_ (
    .A(_793_),
    .Y(_794_)
);

NOR2X1 _3163_ (
    .A(_943_),
    .B(_937_),
    .Y(_795_)
);

AND2X2 _3164_ (
    .A(_795_),
    .B(_794_),
    .Y(_796_)
);

NAND2X1 _3165_ (
    .A(_917_),
    .B(_1193_),
    .Y(_797_)
);

AOI22X1 _3166_ (
    .A(_1193_),
    .B(_926__bF$buf0),
    .C(_881_),
    .D(_905_),
    .Y(_798_)
);

NAND3X1 _3167_ (
    .A(_797_),
    .B(_315_),
    .C(_798_),
    .Y(_799_)
);

NOR2X1 _3168_ (
    .A(_799_),
    .B(_963_),
    .Y(_800_)
);

NAND3X1 _3169_ (
    .A(_796_),
    .B(_800_),
    .C(_791_),
    .Y(_801_)
);

NOR2X1 _3170_ (
    .A(_801_),
    .B(_787_),
    .Y(_802_)
);

NOR2X1 _3171_ (
    .A(_1185_),
    .B(_1277_),
    .Y(_803_)
);

AND2X2 _3172_ (
    .A(_803_),
    .B(_798_),
    .Y(_804_)
);

OAI21X1 _3173_ (
    .A(state[4]),
    .B(_916_),
    .C(_794_),
    .Y(_805_)
);

NOR2X1 _3174_ (
    .A(_963_),
    .B(_805_),
    .Y(_806_)
);

AND2X2 _3175_ (
    .A(_806_),
    .B(_804_),
    .Y(_807_)
);

NAND3X1 _3176_ (
    .A(_977_),
    .B(_978_),
    .C(_807_),
    .Y(_808_)
);

NOR2X1 _3177_ (
    .A(_1347_),
    .B(_1284_),
    .Y(_809_)
);

AND2X2 _3178_ (
    .A(_809_),
    .B(_992_),
    .Y(_810_)
);

NAND3X1 _3179_ (
    .A(_780_),
    .B(_810_),
    .C(_778_),
    .Y(_811_)
);

INVX1 _3180_ (
    .A(_779_),
    .Y(_812_)
);

NAND2X1 _3181_ (
    .A(_776_),
    .B(_812_),
    .Y(_813_)
);

OAI21X1 _3182_ (
    .A(state[5]),
    .B(_996_),
    .C(_952_),
    .Y(_814_)
);

OAI21X1 _3183_ (
    .A(state[4]),
    .B(_1032_),
    .C(_1227_),
    .Y(_815_)
);

NOR2X1 _3184_ (
    .A(_815_),
    .B(_814_),
    .Y(_816_)
);

NAND3X1 _3185_ (
    .A(_1040_),
    .B(_809_),
    .C(_816_),
    .Y(_817_)
);

OAI21X1 _3186_ (
    .A(_813_),
    .B(_817_),
    .C(_811_),
    .Y(_818_)
);

INVX1 _3187_ (
    .A(_976_),
    .Y(_819_)
);

INVX1 _3188_ (
    .A(_1034_),
    .Y(_820_)
);

OAI21X1 _3189_ (
    .A(_946_),
    .B(_993_),
    .C(_933_),
    .Y(_821_)
);

OR2X2 _3190_ (
    .A(_821_),
    .B(_935_),
    .Y(_822_)
);

NOR2X1 _3191_ (
    .A(_820_),
    .B(_822_),
    .Y(_823_)
);

NAND3X1 _3192_ (
    .A(_934_),
    .B(_783_),
    .C(_823_),
    .Y(_824_)
);

NOR2X1 _3193_ (
    .A(_819_),
    .B(_824_),
    .Y(_825_)
);

OAI21X1 _3194_ (
    .A(_937_),
    .B(_821_),
    .C(_822_),
    .Y(_826_)
);

AND2X2 _3195_ (
    .A(_826_),
    .B(_1183_),
    .Y(_827_)
);

AOI22X1 _3196_ (
    .A(_786_),
    .B(_827_),
    .C(_825_),
    .D(_818_),
    .Y(_828_)
);

OAI21X1 _3197_ (
    .A(_808_),
    .B(_828_),
    .C(RDY_bF$buf2),
    .Y(_829_)
);

NOR2X1 _3198_ (
    .A(_802_),
    .B(_829_),
    .Y(_830_)
);

INVX2 _3199_ (
    .A(_830__bF$buf3),
    .Y(_831_)
);

OAI21X1 _3200_ (
    .A(_802_),
    .B(_829_),
    .C(ABL[0]),
    .Y(_832_)
);

OAI21X1 _3201_ (
    .A(_831_),
    .B(_213_),
    .C(_832_),
    .Y(_101_)
);

OAI21X1 _3202_ (
    .A(_802_),
    .B(_829_),
    .C(ABL[1]),
    .Y(_833_)
);

OAI21X1 _3203_ (
    .A(_831_),
    .B(_218_),
    .C(_833_),
    .Y(_102_)
);

OAI21X1 _3204_ (
    .A(_802_),
    .B(_829_),
    .C(ABL[2]),
    .Y(_834_)
);

OAI21X1 _3205_ (
    .A(_831_),
    .B(_223_),
    .C(_834_),
    .Y(_103_)
);

OAI21X1 _3206_ (
    .A(_802_),
    .B(_829_),
    .C(ABL[3]),
    .Y(_835_)
);

OAI21X1 _3207_ (
    .A(_831_),
    .B(_232_),
    .C(_835_),
    .Y(_104_)
);

OAI21X1 _3208_ (
    .A(_802_),
    .B(_829_),
    .C(ABL[4]),
    .Y(_836_)
);

OAI21X1 _3209_ (
    .A(_831_),
    .B(_237_),
    .C(_836_),
    .Y(_105_)
);

OAI21X1 _3210_ (
    .A(_802_),
    .B(_829_),
    .C(ABL[5]),
    .Y(_837_)
);

OAI21X1 _3211_ (
    .A(_831_),
    .B(_245_),
    .C(_837_),
    .Y(_106_)
);

OAI21X1 _3212_ (
    .A(_802_),
    .B(_829_),
    .C(ABL[6]),
    .Y(_838_)
);

OAI21X1 _3213_ (
    .A(_831_),
    .B(_251_),
    .C(_838_),
    .Y(_107_)
);

OAI21X1 _3214_ (
    .A(_802_),
    .B(_829_),
    .C(ABL[7]),
    .Y(_839_)
);

OAI21X1 _3215_ (
    .A(_831_),
    .B(_259_),
    .C(_839_),
    .Y(_108_)
);

OAI21X1 _3216_ (
    .A(_261_),
    .B(_266_),
    .C(_830__bF$buf2),
    .Y(_840_)
);

OAI21X1 _3217_ (
    .A(_1055_),
    .B(_830__bF$buf1),
    .C(_840_),
    .Y(_109_)
);

NAND2X1 _3218_ (
    .A(_1685_[9]),
    .B(_830__bF$buf0),
    .Y(_841_)
);

OAI21X1 _3219_ (
    .A(_1065_),
    .B(_830__bF$buf3),
    .C(_841_),
    .Y(_110_)
);

NAND2X1 _3220_ (
    .A(_1685_[10]),
    .B(_830__bF$buf2),
    .Y(_842_)
);

OAI21X1 _3221_ (
    .A(_273_),
    .B(_830__bF$buf1),
    .C(_842_),
    .Y(_111_)
);

INVX1 _3222_ (
    .A(ABH[3]),
    .Y(_843_)
);

NAND2X1 _3223_ (
    .A(_1685_[11]),
    .B(_830__bF$buf0),
    .Y(_844_)
);

OAI21X1 _3224_ (
    .A(_843_),
    .B(_830__bF$buf3),
    .C(_844_),
    .Y(_112_)
);

NAND2X1 _3225_ (
    .A(_1685_[12]),
    .B(_830__bF$buf2),
    .Y(_845_)
);

OAI21X1 _3226_ (
    .A(_284_),
    .B(_830__bF$buf1),
    .C(_845_),
    .Y(_113_)
);

NAND2X1 _3227_ (
    .A(_1685_[13]),
    .B(_830__bF$buf0),
    .Y(_846_)
);

OAI21X1 _3228_ (
    .A(_292_),
    .B(_830__bF$buf3),
    .C(_846_),
    .Y(_114_)
);

NAND2X1 _3229_ (
    .A(_1685_[14]),
    .B(_830__bF$buf2),
    .Y(_847_)
);

OAI21X1 _3230_ (
    .A(_1108_),
    .B(_830__bF$buf1),
    .C(_847_),
    .Y(_115_)
);

NAND2X1 _3231_ (
    .A(_1685_[15]),
    .B(_830__bF$buf0),
    .Y(_848_)
);

OAI21X1 _3232_ (
    .A(_1118_),
    .B(_830__bF$buf3),
    .C(_848_),
    .Y(_116_)
);

DFFSR _3233_ (
    .CLK(clk_bF$buf10),
    .D(_1483_[0]),
    .Q(state[0]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3234_ (
    .CLK(clk_bF$buf9),
    .D(_1483_[1]),
    .Q(state[1]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3235_ (
    .CLK(clk_bF$buf8),
    .D(_1483_[2]),
    .Q(state[2]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3236_ (
    .CLK(clk_bF$buf7),
    .D(_1483_[3]),
    .Q(state[3]),
    .R(vdd),
    .S(_1__bF$buf7)
);

DFFSR _3237_ (
    .CLK(clk_bF$buf6),
    .D(_1483_[4]),
    .Q(state[4]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3238_ (
    .CLK(clk_bF$buf5),
    .D(_1483_[5]),
    .Q(state[5]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3239_ (
    .CLK(clk_bF$buf4),
    .D(_2_),
    .Q(PC[0]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3240_ (
    .CLK(clk_bF$buf3),
    .D(_3_),
    .Q(PC[1]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3241_ (
    .CLK(clk_bF$buf2),
    .D(_4_),
    .Q(PC[2]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3242_ (
    .CLK(clk_bF$buf1),
    .D(_5_),
    .Q(PC[3]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3243_ (
    .CLK(clk_bF$buf0),
    .D(_6_),
    .Q(PC[4]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3244_ (
    .CLK(clk_bF$buf10),
    .D(_7_),
    .Q(PC[5]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3245_ (
    .CLK(clk_bF$buf9),
    .D(_8_),
    .Q(PC[6]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3246_ (
    .CLK(clk_bF$buf8),
    .D(_9_),
    .Q(PC[7]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3247_ (
    .CLK(clk_bF$buf7),
    .D(_10_),
    .Q(PC[8]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3248_ (
    .CLK(clk_bF$buf6),
    .D(_11_),
    .Q(PC[9]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3249_ (
    .CLK(clk_bF$buf5),
    .D(_12_),
    .Q(PC[10]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3250_ (
    .CLK(clk_bF$buf4),
    .D(_13_),
    .Q(PC[11]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3251_ (
    .CLK(clk_bF$buf3),
    .D(_14_),
    .Q(PC[12]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3252_ (
    .CLK(clk_bF$buf2),
    .D(_15_),
    .Q(PC[13]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3253_ (
    .CLK(clk_bF$buf1),
    .D(_16_),
    .Q(PC[14]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3254_ (
    .CLK(clk_bF$buf0),
    .D(_17_),
    .Q(PC[15]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3255_ (
    .CLK(clk_bF$buf10),
    .D(NMI),
    .Q(NMI_1),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3256_ (
    .CLK(clk_bF$buf9),
    .D(_18_),
    .Q(NMI_edge),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3257_ (
    .CLK(clk_bF$buf8),
    .D(_19_),
    .Q(cond_code[0]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3258_ (
    .CLK(clk_bF$buf7),
    .D(_20_),
    .Q(cond_code[1]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3259_ (
    .CLK(clk_bF$buf6),
    .D(_21_),
    .Q(cond_code[2]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3260_ (
    .CLK(clk_bF$buf5),
    .D(_22_),
    .Q(plp),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3261_ (
    .CLK(clk_bF$buf4),
    .D(_23_),
    .Q(php),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3262_ (
    .CLK(clk_bF$buf3),
    .D(_24_),
    .Q(clc),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3263_ (
    .CLK(clk_bF$buf2),
    .D(_25_),
    .Q(sec),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3264_ (
    .CLK(clk_bF$buf1),
    .D(_26_),
    .Q(cld),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3265_ (
    .CLK(clk_bF$buf0),
    .D(_27_),
    .Q(sed),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3266_ (
    .CLK(clk_bF$buf10),
    .D(_28_),
    .Q(cli),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3267_ (
    .CLK(clk_bF$buf9),
    .D(_29_),
    .Q(sei),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3268_ (
    .CLK(clk_bF$buf8),
    .D(_30_),
    .Q(clv),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3269_ (
    .CLK(clk_bF$buf7),
    .D(_31_),
    .Q(bit_ins),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3270_ (
    .CLK(clk_bF$buf6),
    .D(_32_),
    .Q(op[0]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3271_ (
    .CLK(clk_bF$buf5),
    .D(_33_),
    .Q(op[1]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3272_ (
    .CLK(clk_bF$buf4),
    .D(_34_),
    .Q(op[2]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3273_ (
    .CLK(clk_bF$buf3),
    .D(_35_),
    .Q(op[3]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3274_ (
    .CLK(clk_bF$buf2),
    .D(_36_),
    .Q(rotate),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3275_ (
    .CLK(clk_bF$buf1),
    .D(_37_),
    .Q(shift_right),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3276_ (
    .CLK(clk_bF$buf0),
    .D(_38_),
    .Q(compare),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3277_ (
    .CLK(clk_bF$buf10),
    .D(_39_),
    .Q(shift),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3278_ (
    .CLK(clk_bF$buf9),
    .D(_40_),
    .Q(adc_bcd),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3279_ (
    .CLK(clk_bF$buf8),
    .D(_41_),
    .Q(adc_sbc),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3280_ (
    .CLK(clk_bF$buf7),
    .D(_42_),
    .Q(inc),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3281_ (
    .CLK(clk_bF$buf6),
    .D(_43_),
    .Q(load_only),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3282_ (
    .CLK(clk_bF$buf5),
    .D(_44_),
    .Q(write_back),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3283_ (
    .CLK(clk_bF$buf4),
    .D(_45_),
    .Q(store),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3284_ (
    .CLK(clk_bF$buf3),
    .D(_46_),
    .Q(index_y),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3285_ (
    .CLK(clk_bF$buf2),
    .D(_47_),
    .Q(src_reg[0]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3286_ (
    .CLK(clk_bF$buf1),
    .D(_48_),
    .Q(src_reg[1]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3287_ (
    .CLK(clk_bF$buf0),
    .D(_49_),
    .Q(dst_reg[0]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3288_ (
    .CLK(clk_bF$buf10),
    .D(_50_),
    .Q(dst_reg[1]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3289_ (
    .CLK(clk_bF$buf9),
    .D(_51_),
    .Q(load_reg),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3290_ (
    .CLK(clk_bF$buf8),
    .D(DIMUX[0]),
    .Q(DIHOLD[0]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3291_ (
    .CLK(clk_bF$buf7),
    .D(DIMUX[1]),
    .Q(DIHOLD[1]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3292_ (
    .CLK(clk_bF$buf6),
    .D(DIMUX[2]),
    .Q(DIHOLD[2]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3293_ (
    .CLK(clk_bF$buf5),
    .D(DIMUX[3]),
    .Q(DIHOLD[3]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3294_ (
    .CLK(clk_bF$buf4),
    .D(DIMUX[4]),
    .Q(DIHOLD[4]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3295_ (
    .CLK(clk_bF$buf3),
    .D(DIMUX[5]),
    .Q(DIHOLD[5]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3296_ (
    .CLK(clk_bF$buf2),
    .D(DIMUX[6]),
    .Q(DIHOLD[6]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3297_ (
    .CLK(clk_bF$buf1),
    .D(DIMUX[7]),
    .Q(DIHOLD[7]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3298_ (
    .CLK(clk_bF$buf0),
    .D(_52_),
    .Q(res),
    .R(vdd),
    .S(_1__bF$buf0)
);

DFFPOSX1 _3299_ (
    .CLK(clk_bF$buf10),
    .D(_53_),
    .Q(IRHOLD[0])
);

DFFPOSX1 _3300_ (
    .CLK(clk_bF$buf9),
    .D(_54_),
    .Q(IRHOLD[1])
);

DFFPOSX1 _3301_ (
    .CLK(clk_bF$buf8),
    .D(_55_),
    .Q(IRHOLD[2])
);

DFFPOSX1 _3302_ (
    .CLK(clk_bF$buf7),
    .D(_56_),
    .Q(IRHOLD[3])
);

DFFPOSX1 _3303_ (
    .CLK(clk_bF$buf6),
    .D(_57_),
    .Q(IRHOLD[4])
);

DFFPOSX1 _3304_ (
    .CLK(clk_bF$buf5),
    .D(_58_),
    .Q(IRHOLD[5])
);

DFFPOSX1 _3305_ (
    .CLK(clk_bF$buf4),
    .D(_59_),
    .Q(IRHOLD[6])
);

DFFPOSX1 _3306_ (
    .CLK(clk_bF$buf3),
    .D(_60_),
    .Q(IRHOLD[7])
);

DFFSR _3307_ (
    .CLK(clk_bF$buf2),
    .D(_61_),
    .Q(IRHOLD_valid),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3308_ (
    .CLK(clk_bF$buf1),
    .D(_62_),
    .Q(V),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3309_ (
    .CLK(clk_bF$buf0),
    .D(_63_),
    .Q(D),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3310_ (
    .CLK(clk_bF$buf10),
    .D(_64_),
    .Q(I),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3311_ (
    .CLK(clk_bF$buf9),
    .D(_65_),
    .Q(N),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3312_ (
    .CLK(clk_bF$buf8),
    .D(_66_),
    .Q(Z),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3313_ (
    .CLK(clk_bF$buf7),
    .D(_67_),
    .Q(C),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3314_ (
    .CLK(clk_bF$buf6),
    .D(_68_),
    .Q(backwards),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3315_ (
    .CLK(clk_bF$buf5),
    .D(_69_),
    .Q(\AXYS[0] [0]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3316_ (
    .CLK(clk_bF$buf4),
    .D(_70_),
    .Q(\AXYS[0] [1]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3317_ (
    .CLK(clk_bF$buf3),
    .D(_71_),
    .Q(\AXYS[0] [2]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3318_ (
    .CLK(clk_bF$buf2),
    .D(_72_),
    .Q(\AXYS[0] [3]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3319_ (
    .CLK(clk_bF$buf1),
    .D(_73_),
    .Q(\AXYS[0] [4]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3320_ (
    .CLK(clk_bF$buf0),
    .D(_74_),
    .Q(\AXYS[0] [5]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3321_ (
    .CLK(clk_bF$buf10),
    .D(_75_),
    .Q(\AXYS[0] [6]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3322_ (
    .CLK(clk_bF$buf9),
    .D(_76_),
    .Q(\AXYS[0] [7]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3323_ (
    .CLK(clk_bF$buf8),
    .D(_77_),
    .Q(\AXYS[1] [0]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3324_ (
    .CLK(clk_bF$buf7),
    .D(_78_),
    .Q(\AXYS[1] [1]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3325_ (
    .CLK(clk_bF$buf6),
    .D(_79_),
    .Q(\AXYS[1] [2]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3326_ (
    .CLK(clk_bF$buf5),
    .D(_80_),
    .Q(\AXYS[1] [3]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3327_ (
    .CLK(clk_bF$buf4),
    .D(_81_),
    .Q(\AXYS[1] [4]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3328_ (
    .CLK(clk_bF$buf3),
    .D(_82_),
    .Q(\AXYS[1] [5]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3329_ (
    .CLK(clk_bF$buf2),
    .D(_83_),
    .Q(\AXYS[1] [6]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3330_ (
    .CLK(clk_bF$buf1),
    .D(_84_),
    .Q(\AXYS[1] [7]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3331_ (
    .CLK(clk_bF$buf0),
    .D(_85_),
    .Q(\AXYS[2] [0]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3332_ (
    .CLK(clk_bF$buf10),
    .D(_86_),
    .Q(\AXYS[2] [1]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3333_ (
    .CLK(clk_bF$buf9),
    .D(_87_),
    .Q(\AXYS[2] [2]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3334_ (
    .CLK(clk_bF$buf8),
    .D(_88_),
    .Q(\AXYS[2] [3]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3335_ (
    .CLK(clk_bF$buf7),
    .D(_89_),
    .Q(\AXYS[2] [4]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3336_ (
    .CLK(clk_bF$buf6),
    .D(_90_),
    .Q(\AXYS[2] [5]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3337_ (
    .CLK(clk_bF$buf5),
    .D(_91_),
    .Q(\AXYS[2] [6]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3338_ (
    .CLK(clk_bF$buf4),
    .D(_92_),
    .Q(\AXYS[2] [7]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3339_ (
    .CLK(clk_bF$buf3),
    .D(_0_),
    .Q(adj_bcd),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3340_ (
    .CLK(clk_bF$buf2),
    .D(_93_),
    .Q(\AXYS[3] [0]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3341_ (
    .CLK(clk_bF$buf1),
    .D(_94_),
    .Q(\AXYS[3] [1]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3342_ (
    .CLK(clk_bF$buf0),
    .D(_95_),
    .Q(\AXYS[3] [2]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3343_ (
    .CLK(clk_bF$buf10),
    .D(_96_),
    .Q(\AXYS[3] [3]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3344_ (
    .CLK(clk_bF$buf9),
    .D(_97_),
    .Q(\AXYS[3] [4]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3345_ (
    .CLK(clk_bF$buf8),
    .D(_98_),
    .Q(\AXYS[3] [5]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3346_ (
    .CLK(clk_bF$buf7),
    .D(_99_),
    .Q(\AXYS[3] [6]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3347_ (
    .CLK(clk_bF$buf6),
    .D(_100_),
    .Q(\AXYS[3] [7]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3348_ (
    .CLK(clk_bF$buf5),
    .D(_101_),
    .Q(ABL[0]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3349_ (
    .CLK(clk_bF$buf4),
    .D(_102_),
    .Q(ABL[1]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3350_ (
    .CLK(clk_bF$buf3),
    .D(_103_),
    .Q(ABL[2]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3351_ (
    .CLK(clk_bF$buf2),
    .D(_104_),
    .Q(ABL[3]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3352_ (
    .CLK(clk_bF$buf1),
    .D(_105_),
    .Q(ABL[4]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3353_ (
    .CLK(clk_bF$buf0),
    .D(_106_),
    .Q(ABL[5]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3354_ (
    .CLK(clk_bF$buf10),
    .D(_107_),
    .Q(ABL[6]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3355_ (
    .CLK(clk_bF$buf9),
    .D(_108_),
    .Q(ABL[7]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3356_ (
    .CLK(clk_bF$buf8),
    .D(_109_),
    .Q(ABH[0]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3357_ (
    .CLK(clk_bF$buf7),
    .D(_110_),
    .Q(ABH[1]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3358_ (
    .CLK(clk_bF$buf6),
    .D(_111_),
    .Q(ABH[2]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3359_ (
    .CLK(clk_bF$buf5),
    .D(_112_),
    .Q(ABH[3]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3360_ (
    .CLK(clk_bF$buf4),
    .D(_113_),
    .Q(ABH[4]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3361_ (
    .CLK(clk_bF$buf3),
    .D(_114_),
    .Q(ABH[5]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3362_ (
    .CLK(clk_bF$buf2),
    .D(_115_),
    .Q(ABH[6]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3363_ (
    .CLK(clk_bF$buf1),
    .D(_116_),
    .Q(ABH[7]),
    .R(_1__bF$buf9),
    .S(vdd)
);

OR2X2 _3364_ (
    .A(ADD[0]),
    .B(ADD[3]),
    .Y(_1642_)
);

NOR2X1 _3365_ (
    .A(ADD[5]),
    .B(ADD[4]),
    .Y(_1643_)
);

NOR2X1 _3366_ (
    .A(AN),
    .B(ADD[6]),
    .Y(_1644_)
);

NOR2X1 _3367_ (
    .A(ADD[1]),
    .B(ADD[2]),
    .Y(_1645_)
);

NAND3X1 _3368_ (
    .A(_1643_),
    .B(_1644_),
    .C(_1645_),
    .Y(_1646_)
);

NOR2X1 _3369_ (
    .A(_1642_),
    .B(_1646_),
    .Y(AZ)
);

XOR2X1 _3370_ (
    .A(\u_ALU8.AI7 ),
    .B(CO),
    .Y(_1647_)
);

XNOR2X1 _3371_ (
    .A(AN),
    .B(\u_ALU8.BI7 ),
    .Y(_1648_)
);

XNOR2X1 _3372_ (
    .A(_1647_),
    .B(_1648_),
    .Y(AV)
);

INVX4 _3373_ (
    .A(reset),
    .Y(_1484_)
);

INVX4 _3374_ (
    .A(RDY_bF$buf1),
    .Y(_1649_)
);

NAND2X1 _3375_ (
    .A(alu_shift_right),
    .B(CI),
    .Y(_1650_)
);

INVX2 _3376_ (
    .A(alu_op[1]),
    .Y(_1651_)
);

NAND2X1 _3377_ (
    .A(alu_op[0]),
    .B(_1651_),
    .Y(_1652_)
);

INVX2 _3378_ (
    .A(alu_op[0]),
    .Y(_1653_)
);

AND2X2 _3379_ (
    .A(_1653_),
    .B(BI[7]),
    .Y(_1654_)
);

NAND2X1 _3380_ (
    .A(AI[7]),
    .B(_1654_),
    .Y(_1655_)
);

AOI22X1 _3381_ (
    .A(_1651_),
    .B(BI[7]),
    .C(_1655_),
    .D(_1652_),
    .Y(_1656_)
);

INVX2 _3382_ (
    .A(alu_shift_right),
    .Y(_1657_)
);

OAI21X1 _3383_ (
    .A(AI[7]),
    .B(_1654_),
    .C(_1657_),
    .Y(_1658_)
);

OAI21X1 _3384_ (
    .A(_1658_),
    .B(_1656_),
    .C(_1650_),
    .Y(_1659_)
);

INVX4 _3385_ (
    .A(alu_op[3]),
    .Y(_1660_)
);

OAI21X1 _3386_ (
    .A(alu_op[2]),
    .B(BI[7]),
    .C(_1660_),
    .Y(_1661_)
);

AOI21X1 _3387_ (
    .A(alu_op[2]),
    .B(BI[7]),
    .C(_1661_),
    .Y(_1662_)
);

NOR2X1 _3388_ (
    .A(alu_op[2]),
    .B(_1660_),
    .Y(_1663_)
);

AOI21X1 _3389_ (
    .A(_1659_),
    .B(_1663_),
    .C(_1662_),
    .Y(_1664_)
);

NAND2X1 _3390_ (
    .A(\u_ALU8.BI7 ),
    .B(_1649__bF$buf3),
    .Y(_1665_)
);

OAI21X1 _3391_ (
    .A(_1649__bF$buf2),
    .B(_1664_),
    .C(_1665_),
    .Y(_1485_)
);

INVX1 _3392_ (
    .A(CO),
    .Y(_1666_)
);

OAI21X1 _3393_ (
    .A(_1662_),
    .B(_1663_),
    .C(_1659_),
    .Y(_1667_)
);

NAND2X1 _3394_ (
    .A(alu_shift_right),
    .B(AI[7]),
    .Y(_1668_)
);

AND2X2 _3395_ (
    .A(_1653_),
    .B(BI[6]),
    .Y(_1669_)
);

NAND2X1 _3396_ (
    .A(AI[6]),
    .B(_1669_),
    .Y(_1670_)
);

AOI22X1 _3397_ (
    .A(_1651_),
    .B(BI[6]),
    .C(_1670_),
    .D(_1652_),
    .Y(_1671_)
);

OAI21X1 _3398_ (
    .A(AI[6]),
    .B(_1669_),
    .C(_1657_),
    .Y(_1672_)
);

OAI21X1 _3399_ (
    .A(_1672_),
    .B(_1671_),
    .C(_1668_),
    .Y(_1673_)
);

NAND2X1 _3400_ (
    .A(alu_op[2]),
    .B(_1660_),
    .Y(_1674_)
);

INVX2 _3401_ (
    .A(alu_op[2]),
    .Y(_1675_)
);

OAI21X1 _3402_ (
    .A(alu_op[3]),
    .B(BI[6]),
    .C(_1675_),
    .Y(_1676_)
);

OAI21X1 _3403_ (
    .A(BI[6]),
    .B(_1674_),
    .C(_1676_),
    .Y(_1677_)
);

NAND2X1 _3404_ (
    .A(alu_shift_right),
    .B(AI[6]),
    .Y(_1678_)
);

AND2X2 _3405_ (
    .A(_1653_),
    .B(BI[5]),
    .Y(_1679_)
);

NAND2X1 _3406_ (
    .A(AI[5]),
    .B(_1679_),
    .Y(_1680_)
);

AOI22X1 _3407_ (
    .A(_1651_),
    .B(BI[5]),
    .C(_1680_),
    .D(_1652_),
    .Y(_1681_)
);

OAI21X1 _3408_ (
    .A(AI[5]),
    .B(_1679_),
    .C(_1657_),
    .Y(_1682_)
);

OAI21X1 _3409_ (
    .A(_1682_),
    .B(_1681_),
    .C(_1678_),
    .Y(_1683_)
);

OAI21X1 _3410_ (
    .A(alu_op[3]),
    .B(BI[5]),
    .C(_1675_),
    .Y(_1684_)
);

OAI21X1 _3411_ (
    .A(BI[5]),
    .B(_1674_),
    .C(_1684_),
    .Y(_1497_)
);

NAND2X1 _3412_ (
    .A(_1497_),
    .B(_1683_),
    .Y(_1498_)
);

NAND2X1 _3413_ (
    .A(alu_shift_right),
    .B(AI[5]),
    .Y(_1499_)
);

AND2X2 _3414_ (
    .A(_1653_),
    .B(BI[4]),
    .Y(_1500_)
);

NAND2X1 _3415_ (
    .A(AI[4]),
    .B(_1500_),
    .Y(_1501_)
);

AOI22X1 _3416_ (
    .A(_1651_),
    .B(BI[4]),
    .C(_1501_),
    .D(_1652_),
    .Y(_1502_)
);

OAI21X1 _3417_ (
    .A(AI[4]),
    .B(_1500_),
    .C(_1657_),
    .Y(_1503_)
);

OAI21X1 _3418_ (
    .A(_1503_),
    .B(_1502_),
    .C(_1499_),
    .Y(_1504_)
);

OAI21X1 _3419_ (
    .A(alu_op[3]),
    .B(BI[4]),
    .C(_1675_),
    .Y(_1505_)
);

OAI21X1 _3420_ (
    .A(BI[4]),
    .B(_1674_),
    .C(_1505_),
    .Y(_1506_)
);

NAND2X1 _3421_ (
    .A(alu_shift_right),
    .B(AI[4]),
    .Y(_1507_)
);

AND2X2 _3422_ (
    .A(_1653_),
    .B(BI[3]),
    .Y(_1508_)
);

NAND2X1 _3423_ (
    .A(AI[3]),
    .B(_1508_),
    .Y(_1509_)
);

AOI22X1 _3424_ (
    .A(_1651_),
    .B(BI[3]),
    .C(_1509_),
    .D(_1652_),
    .Y(_1510_)
);

OAI21X1 _3425_ (
    .A(AI[3]),
    .B(_1508_),
    .C(_1657_),
    .Y(_1511_)
);

OAI21X1 _3426_ (
    .A(_1511_),
    .B(_1510_),
    .C(_1507_),
    .Y(_1512_)
);

OAI21X1 _3427_ (
    .A(alu_op[3]),
    .B(BI[3]),
    .C(_1675_),
    .Y(_1513_)
);

OAI21X1 _3428_ (
    .A(BI[3]),
    .B(_1674_),
    .C(_1513_),
    .Y(_1514_)
);

NAND2X1 _3429_ (
    .A(_1514_),
    .B(_1512_),
    .Y(_1515_)
);

INVX1 _3430_ (
    .A(_1663_),
    .Y(_1516_)
);

AND2X2 _3431_ (
    .A(_1514_),
    .B(_1516_),
    .Y(_1517_)
);

OAI21X1 _3432_ (
    .A(_1512_),
    .B(_1517_),
    .C(_1515_),
    .Y(_1518_)
);

INVX1 _3433_ (
    .A(_1518_),
    .Y(_1519_)
);

NAND2X1 _3434_ (
    .A(AI[3]),
    .B(alu_shift_right),
    .Y(_1520_)
);

NAND3X1 _3435_ (
    .A(BI[2]),
    .B(AI[2]),
    .C(_1653_),
    .Y(_1521_)
);

AOI22X1 _3436_ (
    .A(BI[2]),
    .B(_1651_),
    .C(_1521_),
    .D(_1652_),
    .Y(_1522_)
);

INVX1 _3437_ (
    .A(BI[2]),
    .Y(_1523_)
);

INVX1 _3438_ (
    .A(AI[2]),
    .Y(_1524_)
);

OAI21X1 _3439_ (
    .A(alu_op[0]),
    .B(_1523_),
    .C(_1524_),
    .Y(_1525_)
);

NAND2X1 _3440_ (
    .A(_1657_),
    .B(_1525_),
    .Y(_1526_)
);

OAI21X1 _3441_ (
    .A(_1526_),
    .B(_1522_),
    .C(_1520_),
    .Y(_1527_)
);

NOR2X1 _3442_ (
    .A(BI[2]),
    .B(alu_op[3]),
    .Y(_1528_)
);

XOR2X1 _3443_ (
    .A(_1528_),
    .B(_1675_),
    .Y(_1529_)
);

NAND3X1 _3444_ (
    .A(BI[1]),
    .B(AI[1]),
    .C(_1653_),
    .Y(_1530_)
);

AOI22X1 _3445_ (
    .A(_1651_),
    .B(BI[1]),
    .C(_1530_),
    .D(_1652_),
    .Y(_1531_)
);

INVX1 _3446_ (
    .A(BI[1]),
    .Y(_1532_)
);

NOR2X1 _3447_ (
    .A(alu_op[0]),
    .B(_1532_),
    .Y(_1533_)
);

OAI21X1 _3448_ (
    .A(AI[1]),
    .B(_1533_),
    .C(_1657_),
    .Y(_1534_)
);

OAI22X1 _3449_ (
    .A(_1524_),
    .B(_1657_),
    .C(_1531_),
    .D(_1534_),
    .Y(_1535_)
);

OAI21X1 _3450_ (
    .A(alu_op[2]),
    .B(BI[1]),
    .C(_1660_),
    .Y(_1536_)
);

AOI21X1 _3451_ (
    .A(alu_op[2]),
    .B(BI[1]),
    .C(_1536_),
    .Y(_1537_)
);

OAI21X1 _3452_ (
    .A(_1663_),
    .B(_1537_),
    .C(_1535_),
    .Y(_1538_)
);

NAND2X1 _3453_ (
    .A(BI[0]),
    .B(_1653_),
    .Y(_1539_)
);

NAND2X1 _3454_ (
    .A(alu_op[1]),
    .B(AI[0]),
    .Y(_1540_)
);

AOI22X1 _3455_ (
    .A(BI[0]),
    .B(_1540_),
    .C(_1652_),
    .D(_1539_),
    .Y(_1541_)
);

INVX1 _3456_ (
    .A(BI[0]),
    .Y(_1542_)
);

INVX1 _3457_ (
    .A(AI[0]),
    .Y(_1543_)
);

OAI21X1 _3458_ (
    .A(alu_op[0]),
    .B(_1542_),
    .C(_1543_),
    .Y(_1544_)
);

NAND2X1 _3459_ (
    .A(_1657_),
    .B(_1544_),
    .Y(_1545_)
);

NAND2X1 _3460_ (
    .A(alu_shift_right),
    .B(AI[1]),
    .Y(_1546_)
);

OAI21X1 _3461_ (
    .A(_1541_),
    .B(_1545_),
    .C(_1546_),
    .Y(_1547_)
);

OAI21X1 _3462_ (
    .A(alu_op[2]),
    .B(BI[0]),
    .C(_1660_),
    .Y(_1548_)
);

INVX1 _3463_ (
    .A(_1548_),
    .Y(_1549_)
);

OAI21X1 _3464_ (
    .A(_1675_),
    .B(_1542_),
    .C(_1549_),
    .Y(_1550_)
);

OAI21X1 _3465_ (
    .A(_1660_),
    .B(alu_op[2]),
    .C(_1550_),
    .Y(_1551_)
);

OAI21X1 _3466_ (
    .A(_1660_),
    .B(_1675_),
    .C(CI),
    .Y(_1552_)
);

NOR2X1 _3467_ (
    .A(alu_shift_right),
    .B(_1552_),
    .Y(_1553_)
);

MUX2X1 _3468_ (
    .A(alu_op[1]),
    .B(_1542_),
    .S(alu_op[0]),
    .Y(_1554_)
);

NAND2X1 _3469_ (
    .A(BI[0]),
    .B(_1540_),
    .Y(_1555_)
);

NAND2X1 _3470_ (
    .A(_1555_),
    .B(_1554_),
    .Y(_1556_)
);

AOI21X1 _3471_ (
    .A(_1539_),
    .B(_1543_),
    .C(alu_shift_right),
    .Y(_1557_)
);

NAND2X1 _3472_ (
    .A(_1557_),
    .B(_1556_),
    .Y(_1558_)
);

NAND3X1 _3473_ (
    .A(_1546_),
    .B(_1550_),
    .C(_1558_),
    .Y(_1559_)
);

AOI22X1 _3474_ (
    .A(_1547_),
    .B(_1551_),
    .C(_1559_),
    .D(_1553_),
    .Y(_1560_)
);

NOR2X1 _3475_ (
    .A(_1537_),
    .B(_1535_),
    .Y(_1561_)
);

OAI21X1 _3476_ (
    .A(_1561_),
    .B(_1560_),
    .C(_1538_),
    .Y(_1562_)
);

NAND2X1 _3477_ (
    .A(_1529_),
    .B(_1527_),
    .Y(_1563_)
);

NAND2X1 _3478_ (
    .A(_1660_),
    .B(_1529_),
    .Y(_1564_)
);

INVX1 _3479_ (
    .A(_1564_),
    .Y(_1565_)
);

OAI21X1 _3480_ (
    .A(_1527_),
    .B(_1565_),
    .C(_1563_),
    .Y(_1566_)
);

INVX1 _3481_ (
    .A(_1566_),
    .Y(_1567_)
);

AOI22X1 _3482_ (
    .A(_1527_),
    .B(_1529_),
    .C(_1562_),
    .D(_1567_),
    .Y(_1568_)
);

XOR2X1 _3483_ (
    .A(_1568_),
    .B(_1519_),
    .Y(_1569_)
);

AOI21X1 _3484_ (
    .A(alu_op[2]),
    .B(BI[0]),
    .C(_1548_),
    .Y(_1570_)
);

OAI21X1 _3485_ (
    .A(_1663_),
    .B(_1570_),
    .C(_1547_),
    .Y(_1571_)
);

INVX1 _3486_ (
    .A(_1553_),
    .Y(_1572_)
);

NOR2X1 _3487_ (
    .A(_1570_),
    .B(_1547_),
    .Y(_1573_)
);

OAI21X1 _3488_ (
    .A(_1572_),
    .B(_1573_),
    .C(_1571_),
    .Y(_1574_)
);

INVX1 _3489_ (
    .A(_1537_),
    .Y(_1575_)
);

OAI21X1 _3490_ (
    .A(_1660_),
    .B(alu_op[2]),
    .C(_1575_),
    .Y(_1576_)
);

MUX2X1 _3491_ (
    .A(_1576_),
    .B(_1575_),
    .S(_1535_),
    .Y(_1577_)
);

NAND2X1 _3492_ (
    .A(_1577_),
    .B(_1574_),
    .Y(_1578_)
);

OAI21X1 _3493_ (
    .A(_1535_),
    .B(_1537_),
    .C(_1538_),
    .Y(_1579_)
);

NAND2X1 _3494_ (
    .A(_1560_),
    .B(_1579_),
    .Y(_1580_)
);

NAND2X1 _3495_ (
    .A(_1580_),
    .B(_1578_),
    .Y(_1581_)
);

NAND2X1 _3496_ (
    .A(_1566_),
    .B(_1562_),
    .Y(_1582_)
);

NAND3X1 _3497_ (
    .A(_1538_),
    .B(_1567_),
    .C(_1578_),
    .Y(_1583_)
);

NAND3X1 _3498_ (
    .A(_1582_),
    .B(_1581_),
    .C(_1583_),
    .Y(_1584_)
);

NAND2X1 _3499_ (
    .A(\u_ALU8.BCD ),
    .B(_1584_),
    .Y(_1585_)
);

OAI21X1 _3500_ (
    .A(_1518_),
    .B(_1568_),
    .C(_1515_),
    .Y(_1586_)
);

INVX1 _3501_ (
    .A(_1586_),
    .Y(_1587_)
);

OAI21X1 _3502_ (
    .A(_1585_),
    .B(_1569_),
    .C(_1587_),
    .Y(_1588_)
);

NAND2X1 _3503_ (
    .A(_1506_),
    .B(_1504_),
    .Y(_1589_)
);

OAI21X1 _3504_ (
    .A(_1660_),
    .B(alu_op[2]),
    .C(_1506_),
    .Y(_1590_)
);

INVX1 _3505_ (
    .A(_1590_),
    .Y(_1591_)
);

OAI21X1 _3506_ (
    .A(_1504_),
    .B(_1591_),
    .C(_1589_),
    .Y(_1592_)
);

INVX1 _3507_ (
    .A(_1592_),
    .Y(_1593_)
);

AOI22X1 _3508_ (
    .A(_1504_),
    .B(_1506_),
    .C(_1588_),
    .D(_1593_),
    .Y(_1594_)
);

OAI21X1 _3509_ (
    .A(_1660_),
    .B(alu_op[2]),
    .C(_1497_),
    .Y(_1595_)
);

INVX1 _3510_ (
    .A(_1595_),
    .Y(_1596_)
);

OAI21X1 _3511_ (
    .A(_1683_),
    .B(_1596_),
    .C(_1498_),
    .Y(_1597_)
);

OAI21X1 _3512_ (
    .A(_1597_),
    .B(_1594_),
    .C(_1498_),
    .Y(_1598_)
);

NAND2X1 _3513_ (
    .A(_1677_),
    .B(_1673_),
    .Y(_1599_)
);

OAI21X1 _3514_ (
    .A(_1660_),
    .B(alu_op[2]),
    .C(_1677_),
    .Y(_1600_)
);

INVX1 _3515_ (
    .A(_1600_),
    .Y(_1601_)
);

OAI21X1 _3516_ (
    .A(_1673_),
    .B(_1601_),
    .C(_1599_),
    .Y(_1602_)
);

INVX1 _3517_ (
    .A(_1602_),
    .Y(_1603_)
);

AOI22X1 _3518_ (
    .A(_1673_),
    .B(_1677_),
    .C(_1598_),
    .D(_1603_),
    .Y(_1604_)
);

OAI21X1 _3519_ (
    .A(_1659_),
    .B(_1662_),
    .C(_1667_),
    .Y(_1605_)
);

OAI21X1 _3520_ (
    .A(_1605_),
    .B(_1604_),
    .C(_1667_),
    .Y(_1606_)
);

NAND2X1 _3521_ (
    .A(alu_shift_right),
    .B(AI[0]),
    .Y(_1607_)
);

XOR2X1 _3522_ (
    .A(_1606_),
    .B(_1607_),
    .Y(_1608_)
);

XOR2X1 _3523_ (
    .A(_1604_),
    .B(_1605_),
    .Y(_1609_)
);

INVX1 _3524_ (
    .A(\u_ALU8.BCD ),
    .Y(_1610_)
);

XOR2X1 _3525_ (
    .A(_1568_),
    .B(_1518_),
    .Y(_1611_)
);

XOR2X1 _3526_ (
    .A(_1562_),
    .B(_1566_),
    .Y(_1612_)
);

AOI21X1 _3527_ (
    .A(_1612_),
    .B(_1581_),
    .C(_1610_),
    .Y(_1613_)
);

AOI21X1 _3528_ (
    .A(_1613_),
    .B(_1611_),
    .C(_1586_),
    .Y(_1614_)
);

OAI21X1 _3529_ (
    .A(_1592_),
    .B(_1614_),
    .C(_1589_),
    .Y(_1615_)
);

INVX1 _3530_ (
    .A(_1597_),
    .Y(_1616_)
);

NAND2X1 _3531_ (
    .A(_1616_),
    .B(_1615_),
    .Y(_1617_)
);

NAND2X1 _3532_ (
    .A(_1597_),
    .B(_1594_),
    .Y(_1618_)
);

NAND2X1 _3533_ (
    .A(_1618_),
    .B(_1617_),
    .Y(_1619_)
);

NAND2X1 _3534_ (
    .A(_1603_),
    .B(_1598_),
    .Y(_1620_)
);

NAND3X1 _3535_ (
    .A(_1498_),
    .B(_1602_),
    .C(_1617_),
    .Y(_1621_)
);

NAND2X1 _3536_ (
    .A(_1621_),
    .B(_1620_),
    .Y(_1622_)
);

AOI21X1 _3537_ (
    .A(_1622_),
    .B(_1619_),
    .C(_1610_),
    .Y(_1623_)
);

AOI21X1 _3538_ (
    .A(_1609_),
    .B(_1623_),
    .C(_1649__bF$buf1),
    .Y(_1624_)
);

AOI22X1 _3539_ (
    .A(_1666_),
    .B(_1649__bF$buf0),
    .C(_1624_),
    .D(_1608_),
    .Y(_1486_)
);

NAND2X1 _3540_ (
    .A(HC),
    .B(_1649__bF$buf3),
    .Y(_1625_)
);

OAI21X1 _3541_ (
    .A(_1649__bF$buf2),
    .B(_1614_),
    .C(_1625_),
    .Y(_1487_)
);

NAND2X1 _3542_ (
    .A(ADD[0]),
    .B(_1649__bF$buf1),
    .Y(_1626_)
);

AOI21X1 _3543_ (
    .A(_1571_),
    .B(_1559_),
    .C(_1553_),
    .Y(_1627_)
);

OAI21X1 _3544_ (
    .A(_1547_),
    .B(_1570_),
    .C(_1571_),
    .Y(_1628_)
);

OAI21X1 _3545_ (
    .A(_1572_),
    .B(_1628_),
    .C(RDY_bF$buf0),
    .Y(_1629_)
);

OAI21X1 _3546_ (
    .A(_1627_),
    .B(_1629_),
    .C(_1626_),
    .Y(_1488_)
);

NAND2X1 _3547_ (
    .A(ADD[1]),
    .B(_1649__bF$buf0),
    .Y(_1630_)
);

OAI21X1 _3548_ (
    .A(_1649__bF$buf3),
    .B(_1581_),
    .C(_1630_),
    .Y(_1489_)
);

NAND2X1 _3549_ (
    .A(ADD[2]),
    .B(_1649__bF$buf2),
    .Y(_1631_)
);

OAI21X1 _3550_ (
    .A(_1649__bF$buf1),
    .B(_1612_),
    .C(_1631_),
    .Y(_1490_)
);

NAND2X1 _3551_ (
    .A(ADD[3]),
    .B(_1649__bF$buf0),
    .Y(_1632_)
);

OAI21X1 _3552_ (
    .A(_1649__bF$buf3),
    .B(_1569_),
    .C(_1632_),
    .Y(_1491_)
);

NAND2X1 _3553_ (
    .A(ADD[4]),
    .B(_1649__bF$buf2),
    .Y(_1633_)
);

NOR2X1 _3554_ (
    .A(_1593_),
    .B(_1588_),
    .Y(_1634_)
);

OAI21X1 _3555_ (
    .A(_1592_),
    .B(_1614_),
    .C(RDY_bF$buf8),
    .Y(_1635_)
);

OAI21X1 _3556_ (
    .A(_1634_),
    .B(_1635_),
    .C(_1633_),
    .Y(_1492_)
);

NAND2X1 _3557_ (
    .A(ADD[5]),
    .B(_1649__bF$buf1),
    .Y(_1636_)
);

OAI21X1 _3558_ (
    .A(_1649__bF$buf0),
    .B(_1619_),
    .C(_1636_),
    .Y(_1493_)
);

NAND2X1 _3559_ (
    .A(ADD[6]),
    .B(_1649__bF$buf3),
    .Y(_1637_)
);

OAI21X1 _3560_ (
    .A(_1649__bF$buf2),
    .B(_1622_),
    .C(_1637_),
    .Y(_1494_)
);

INVX1 _3561_ (
    .A(AN),
    .Y(_1638_)
);

NAND2X1 _3562_ (
    .A(RDY_bF$buf7),
    .B(_1609_),
    .Y(_1639_)
);

OAI21X1 _3563_ (
    .A(_1638_),
    .B(RDY_bF$buf6),
    .C(_1639_),
    .Y(_1495_)
);

INVX1 _3564_ (
    .A(\u_ALU8.AI7 ),
    .Y(_1640_)
);

NAND2X1 _3565_ (
    .A(AI[7]),
    .B(RDY_bF$buf5),
    .Y(_1641_)
);

OAI21X1 _3566_ (
    .A(RDY_bF$buf4),
    .B(_1640_),
    .C(_1641_),
    .Y(_1496_)
);

DFFSR _3567_ (
    .CLK(clk_bF$buf0),
    .D(_1485_),
    .Q(\u_ALU8.BI7 ),
    .R(_1484_),
    .S(vdd)
);

DFFSR _3568_ (
    .CLK(clk_bF$buf10),
    .D(_1486_),
    .Q(CO),
    .R(_1484_),
    .S(vdd)
);

DFFSR _3569_ (
    .CLK(clk_bF$buf9),
    .D(_1487_),
    .Q(HC),
    .R(_1484_),
    .S(vdd)
);

DFFSR _3570_ (
    .CLK(clk_bF$buf8),
    .D(_1488_),
    .Q(ADD[0]),
    .R(_1484_),
    .S(vdd)
);

DFFSR _3571_ (
    .CLK(clk_bF$buf7),
    .D(_1489_),
    .Q(ADD[1]),
    .R(_1484_),
    .S(vdd)
);

DFFSR _3572_ (
    .CLK(clk_bF$buf6),
    .D(_1490_),
    .Q(ADD[2]),
    .R(_1484_),
    .S(vdd)
);

DFFSR _3573_ (
    .CLK(clk_bF$buf5),
    .D(_1491_),
    .Q(ADD[3]),
    .R(_1484_),
    .S(vdd)
);

DFFSR _3574_ (
    .CLK(clk_bF$buf4),
    .D(_1492_),
    .Q(ADD[4]),
    .R(_1484_),
    .S(vdd)
);

DFFSR _3575_ (
    .CLK(clk_bF$buf3),
    .D(_1493_),
    .Q(ADD[5]),
    .R(_1484_),
    .S(vdd)
);

DFFSR _3576_ (
    .CLK(clk_bF$buf2),
    .D(_1494_),
    .Q(ADD[6]),
    .R(_1484_),
    .S(vdd)
);

DFFSR _3577_ (
    .CLK(clk_bF$buf1),
    .D(_1495_),
    .Q(AN),
    .R(_1484_),
    .S(vdd)
);

DFFSR _3578_ (
    .CLK(clk_bF$buf0),
    .D(_1496_),
    .Q(\u_ALU8.AI7 ),
    .R(_1484_),
    .S(vdd)
);

BUFX2 _3579_ (
    .A(_1685_[0]),
    .Y(AB[0])
);

BUFX2 _3580_ (
    .A(_1685_[1]),
    .Y(AB[1])
);

BUFX2 _3581_ (
    .A(_1685_[10]),
    .Y(AB[10])
);

BUFX2 _3582_ (
    .A(_1685_[11]),
    .Y(AB[11])
);

BUFX2 _3583_ (
    .A(_1685_[12]),
    .Y(AB[12])
);

BUFX2 _3584_ (
    .A(_1685_[13]),
    .Y(AB[13])
);

BUFX2 _3585_ (
    .A(_1685_[14]),
    .Y(AB[14])
);

BUFX2 _3586_ (
    .A(_1685_[15]),
    .Y(AB[15])
);

BUFX2 _3587_ (
    .A(_1685_[2]),
    .Y(AB[2])
);

BUFX2 _3588_ (
    .A(_1685_[3]),
    .Y(AB[3])
);

BUFX2 _3589_ (
    .A(_1685_[4]),
    .Y(AB[4])
);

BUFX2 _3590_ (
    .A(_1685_[5]),
    .Y(AB[5])
);

BUFX2 _3591_ (
    .A(_1685_[6]),
    .Y(AB[6])
);

BUFX2 _3592_ (
    .A(_1685_[7]),
    .Y(AB[7])
);

BUFX2 _3593_ (
    .A(_1685_[8]),
    .Y(AB[8])
);

BUFX2 _3594_ (
    .A(_1685_[9]),
    .Y(AB[9])
);

BUFX2 _3595_ (
    .A(_1686_[0]),
    .Y(DO[0])
);

BUFX2 _3596_ (
    .A(_1686_[1]),
    .Y(DO[1])
);

BUFX2 _3597_ (
    .A(_1686_[2]),
    .Y(DO[2])
);

BUFX2 _3598_ (
    .A(_1686_[3]),
    .Y(DO[3])
);

BUFX2 _3599_ (
    .A(_1686_[4]),
    .Y(DO[4])
);

BUFX2 _3600_ (
    .A(_1686_[5]),
    .Y(DO[5])
);

BUFX2 _3601_ (
    .A(_1686_[6]),
    .Y(DO[6])
);

BUFX2 _3602_ (
    .A(_1686_[7]),
    .Y(DO[7])
);

BUFX2 _3603_ (
    .A(_1687_),
    .Y(WE)
);

endmodule
