magic
tech scmos
magscale 1 2
timestamp 1739518439
<< error_s >>
rect 4 11284 11356 11296
rect 4 11044 11356 11056
rect 4 10804 11356 10816
rect 4 10564 11356 10576
rect 4 10324 11356 10336
rect 4 10084 11356 10096
rect 4 9844 11356 9856
rect 4 9604 11356 9616
rect 4 9364 11356 9376
rect 4 9124 11356 9136
rect 4 8884 11356 8896
rect 4 8644 11356 8656
rect 4 8404 11356 8416
rect 4 8164 11356 8176
rect 4 7924 11356 7936
rect 4 7684 11356 7696
rect 4 7444 11356 7456
rect 4 7204 11356 7216
rect 4 6964 11356 6976
rect 4 6724 11356 6736
rect 4 6484 11356 6496
rect 4 6244 11356 6256
rect 4 6004 11356 6016
rect 4 5764 11356 5776
rect 4 5524 11356 5536
rect 4 5284 11356 5296
rect 4 5044 11356 5056
rect 4 4804 11356 4816
rect 4 4564 11356 4576
rect 4 4324 11356 4336
rect 4 4084 11356 4096
rect 4 3844 11356 3856
rect 4 3604 11356 3616
rect 4 3364 11356 3376
rect 4 3124 11356 3136
rect 4 2884 11356 2896
rect 4 2644 11356 2656
rect 4 2404 11356 2416
rect 4 2164 11356 2176
rect 4 1924 11356 1936
rect 4 1684 11356 1696
rect 4 1444 11356 1456
rect 4 1204 11356 1216
rect 4 964 11356 976
rect 4 724 11356 736
rect 4 484 11356 496
rect 4 244 11356 256
rect 4 4 11356 16
<< metal1 >>
rect -62 11058 -2 11298
rect 11330 11282 11422 11298
rect 1347 11217 1433 11223
rect 8947 11197 9133 11203
rect -62 11042 30 11058
rect -62 10578 -2 11042
rect 11362 10818 11422 11282
rect 11330 10802 11422 10818
rect 10967 10777 11073 10783
rect 4567 10717 4613 10723
rect 8767 10677 8833 10683
rect -62 10562 30 10578
rect -62 10098 -2 10562
rect 6257 10543 6263 10563
rect 6207 10537 6263 10543
rect 10947 10457 11013 10463
rect 6247 10417 6273 10423
rect 11362 10338 11422 10802
rect 11330 10322 11422 10338
rect -62 10082 30 10098
rect -62 9618 -2 10082
rect 737 10063 743 10083
rect 737 10057 773 10063
rect 8467 9977 8513 9983
rect 2627 9877 2753 9883
rect 11362 9858 11422 10322
rect 11330 9842 11422 9858
rect -62 9602 30 9618
rect -62 9138 -2 9602
rect 397 9583 403 9603
rect 307 9577 403 9583
rect 4027 9497 4073 9503
rect 2987 9437 3073 9443
rect 5347 9437 5493 9443
rect 5827 9437 5893 9443
rect 10587 9437 10633 9443
rect 11362 9378 11422 9842
rect 11330 9362 11422 9378
rect 3767 9297 3853 9303
rect 6787 9297 6833 9303
rect -62 9122 30 9138
rect -62 8658 -2 9122
rect 5687 9097 5713 9103
rect 8827 9057 8853 9063
rect 2127 9017 2213 9023
rect 4507 8937 4533 8943
rect 11362 8898 11422 9362
rect 11330 8882 11422 8898
rect 5567 8797 5653 8803
rect 2147 8757 2213 8763
rect -62 8642 30 8658
rect -62 8178 -2 8642
rect 177 8623 183 8643
rect 87 8617 183 8623
rect 6247 8577 6293 8583
rect 5947 8497 6033 8503
rect 6547 8497 6613 8503
rect 9367 8477 9413 8483
rect 11362 8418 11422 8882
rect 11330 8402 11422 8418
rect 6927 8377 7013 8383
rect 3607 8317 3673 8323
rect -62 8162 30 8178
rect -62 7698 -2 8162
rect 6107 8097 6193 8103
rect 6227 8077 6273 8083
rect 5907 8057 5953 8063
rect 5387 7997 5413 8003
rect 5427 7997 5433 8003
rect 6127 7997 6293 8003
rect 4727 7977 4813 7983
rect 5207 7957 5273 7963
rect 11362 7938 11422 8402
rect 11330 7922 11422 7938
rect 6507 7877 6553 7883
rect 7207 7877 7313 7883
rect 2447 7857 2533 7863
rect 4087 7857 4173 7863
rect 7967 7857 8073 7863
rect 4787 7777 4913 7783
rect 5927 7757 6013 7763
rect 87 7717 93 7723
rect 107 7717 163 7723
rect -62 7682 30 7698
rect 157 7697 163 7717
rect -62 7218 -2 7682
rect 7397 7617 7413 7623
rect 5727 7577 5773 7583
rect 747 7537 893 7543
rect 7397 7543 7403 7617
rect 7397 7537 7413 7543
rect 7527 7517 7593 7523
rect 11362 7458 11422 7922
rect 11330 7442 11422 7458
rect 5527 7417 5573 7423
rect 3747 7377 3893 7383
rect 1817 7357 1833 7363
rect 1817 7283 1823 7357
rect 7727 7337 7873 7343
rect 7987 7317 8033 7323
rect 2167 7297 2313 7303
rect 1817 7277 1833 7283
rect -62 7202 30 7218
rect -62 6738 -2 7202
rect 4827 7137 4953 7143
rect 5827 7037 5953 7043
rect 5327 6997 5433 7003
rect 11362 6978 11422 7442
rect 11330 6962 11422 6978
rect 8567 6917 8593 6923
rect 4127 6877 4293 6883
rect 8007 6877 8053 6883
rect 1867 6857 1893 6863
rect 4707 6837 4813 6843
rect 3427 6817 3533 6823
rect 787 6797 813 6803
rect 567 6757 633 6763
rect 647 6757 663 6763
rect -62 6722 30 6738
rect 657 6737 663 6757
rect -62 6258 -2 6722
rect 6767 6617 6793 6623
rect 11362 6498 11422 6962
rect 11330 6482 11422 6498
rect 287 6423 293 6441
rect 287 6417 433 6423
rect 8347 6337 8393 6343
rect -62 6242 30 6258
rect -62 5778 -2 6242
rect 4057 6223 4063 6243
rect 3987 6217 4063 6223
rect 6967 6177 7133 6183
rect 1287 6157 1393 6163
rect 8087 6137 8153 6143
rect 1007 6097 1093 6103
rect 11362 6018 11422 6482
rect 11330 6002 11422 6018
rect 5347 5977 5373 5983
rect 11187 5897 11213 5903
rect 1927 5797 2083 5803
rect -62 5762 30 5778
rect 2077 5777 2083 5797
rect -62 5298 -2 5762
rect 6127 5657 6193 5663
rect 1647 5637 1713 5643
rect 3047 5617 3073 5623
rect 6487 5597 6633 5603
rect 10047 5597 10113 5603
rect 11362 5538 11422 6002
rect 11330 5522 11422 5538
rect 3007 5497 3113 5503
rect 9867 5437 9993 5443
rect 6147 5417 6253 5423
rect 2747 5397 2773 5403
rect 8907 5397 8973 5403
rect 2327 5317 2383 5323
rect -62 5282 30 5298
rect 2377 5297 2383 5317
rect -62 4818 -2 5282
rect 157 5263 163 5283
rect 87 5257 163 5263
rect 8267 5257 8333 5263
rect 7787 5197 7813 5203
rect 9687 5137 9773 5143
rect 6867 5097 6893 5103
rect 11362 5058 11422 5522
rect 11330 5042 11422 5058
rect 8447 4957 8553 4963
rect -62 4802 30 4818
rect -62 4338 -2 4802
rect 11107 4637 11193 4643
rect 11362 4578 11422 5042
rect 11330 4562 11422 4578
rect 9257 4497 9413 4503
rect 7787 4477 7833 4483
rect 9257 4483 9263 4497
rect 9227 4477 9263 4483
rect 4187 4437 4393 4443
rect 4747 4437 4773 4443
rect 9627 4417 9673 4423
rect -62 4322 30 4338
rect -62 3858 -2 4322
rect 6137 4303 6143 4323
rect 6137 4297 6213 4303
rect 3787 4177 3953 4183
rect 5547 4157 5573 4163
rect 9327 4157 9353 4163
rect 11362 4098 11422 4562
rect 11330 4082 11422 4098
rect 6767 4057 6813 4063
rect 11127 4017 11173 4023
rect 7647 3957 7753 3963
rect 10487 3937 10513 3943
rect 5847 3897 5873 3903
rect -62 3842 30 3858
rect -62 3378 -2 3842
rect 1737 3823 1743 3843
rect 1737 3817 1833 3823
rect 9127 3737 9193 3743
rect 6687 3717 6773 3723
rect 8567 3677 8713 3683
rect 9287 3657 9313 3663
rect 9027 3637 9113 3643
rect 11362 3618 11422 4082
rect 11330 3602 11422 3618
rect 10147 3537 10253 3543
rect -62 3362 30 3378
rect -62 2898 -2 3362
rect 687 3257 813 3263
rect 6327 3257 6353 3263
rect 6287 3217 6373 3223
rect 10167 3217 10233 3223
rect 10307 3197 10353 3203
rect 11362 3138 11422 3602
rect 11330 3122 11422 3138
rect 7827 3077 7893 3083
rect 6407 3057 6433 3063
rect 8067 3057 8133 3063
rect 10627 3057 10793 3063
rect 3107 3017 3193 3023
rect 9987 2997 10093 3003
rect 10067 2977 10093 2983
rect 10507 2957 10553 2963
rect -62 2882 30 2898
rect -62 2418 -2 2882
rect 8601 2717 8673 2723
rect 11362 2658 11422 3122
rect 11330 2642 11422 2658
rect 11107 2597 11133 2603
rect 3127 2577 3273 2583
rect 6367 2577 6413 2583
rect 6667 2577 6693 2583
rect 2087 2517 2153 2523
rect 10647 2517 10753 2523
rect 9947 2477 9993 2483
rect 1767 2437 1783 2443
rect -62 2402 30 2418
rect 1777 2417 1783 2437
rect -62 1938 -2 2402
rect 9147 2217 9253 2223
rect 11362 2178 11422 2642
rect 11330 2162 11422 2178
rect 2747 2097 2793 2103
rect 6907 2097 6953 2103
rect 8207 2097 8353 2103
rect 9687 2097 9713 2103
rect 10727 2097 10773 2103
rect 11067 2097 11133 2103
rect 9787 2017 9853 2023
rect -62 1922 30 1938
rect -62 1458 -2 1922
rect 8737 1783 8743 1793
rect 8737 1777 8873 1783
rect 11362 1698 11422 2162
rect 11330 1682 11422 1698
rect -62 1442 30 1458
rect -62 978 -2 1442
rect 2967 1357 3053 1363
rect 11362 1218 11422 1682
rect 11330 1202 11422 1218
rect 2347 1157 2413 1163
rect 5787 1137 5873 1143
rect 5927 1137 6093 1143
rect 6307 1137 6333 1143
rect 6547 1137 6593 1143
rect 7687 1137 7873 1143
rect 8287 1137 8453 1143
rect 9507 1117 9613 1123
rect -62 962 30 978
rect -62 498 -2 962
rect 8397 807 8403 853
rect 8607 817 8633 823
rect 6361 797 6453 803
rect 10207 797 10253 803
rect 11362 738 11422 1202
rect 11330 722 11422 738
rect 8707 657 8853 663
rect 9547 577 9593 583
rect -62 482 30 498
rect -62 18 -2 482
rect 8367 317 8513 323
rect 11362 258 11422 722
rect 11330 242 11422 258
rect 5827 157 6013 163
rect 10587 117 10633 123
rect -62 2 30 18
rect 11362 2 11422 242
<< m2contact >>
rect 1333 11213 1347 11227
rect 1433 11213 1447 11227
rect 8933 11193 8947 11207
rect 9133 11193 9147 11207
rect 533 11033 547 11047
rect 1553 11033 1567 11047
rect 2193 11033 2207 11047
rect 2813 11033 2827 11047
rect 3193 11033 3207 11047
rect 4713 11033 4727 11047
rect 6213 11033 6227 11047
rect 7573 11033 7587 11047
rect 10953 10773 10967 10787
rect 11073 10773 11087 10787
rect 4553 10713 4567 10727
rect 4613 10713 4627 10727
rect 8753 10673 8767 10687
rect 8833 10673 8847 10687
rect 4733 10553 4747 10567
rect 5233 10553 5247 10567
rect 6193 10533 6207 10547
rect 7033 10553 7047 10567
rect 7873 10553 7887 10567
rect 8273 10553 8287 10567
rect 8953 10553 8967 10567
rect 9713 10553 9727 10567
rect 10933 10453 10947 10467
rect 11013 10453 11027 10467
rect 6233 10413 6247 10427
rect 6273 10413 6287 10427
rect 4733 10093 4747 10107
rect 9753 10093 9767 10107
rect 5733 10073 5747 10087
rect 5873 10073 5887 10087
rect 773 10053 787 10067
rect 8453 9973 8467 9987
rect 8513 9973 8527 9987
rect 2613 9873 2627 9887
rect 2753 9873 2767 9887
rect 7493 9613 7507 9627
rect 293 9573 307 9587
rect 2013 9593 2027 9607
rect 7993 9593 8007 9607
rect 8733 9593 8747 9607
rect 9873 9593 9887 9607
rect 4013 9493 4027 9507
rect 4073 9493 4087 9507
rect 2973 9433 2987 9447
rect 3073 9433 3087 9447
rect 5333 9433 5347 9447
rect 5493 9433 5507 9447
rect 5813 9433 5827 9447
rect 5893 9433 5907 9447
rect 10573 9433 10587 9447
rect 10633 9433 10647 9447
rect 3753 9293 3767 9307
rect 3853 9293 3867 9307
rect 6773 9293 6787 9307
rect 6833 9293 6847 9307
rect 93 9113 107 9127
rect 153 9113 167 9127
rect 773 9113 787 9127
rect 3613 9113 3627 9127
rect 5673 9093 5687 9107
rect 5713 9093 5727 9107
rect 8813 9053 8827 9067
rect 8853 9053 8867 9067
rect 2113 9013 2127 9027
rect 2213 9013 2227 9027
rect 4493 8933 4507 8947
rect 4533 8933 4547 8947
rect 5553 8793 5567 8807
rect 5653 8793 5667 8807
rect 2133 8753 2147 8767
rect 2213 8753 2227 8767
rect 3113 8653 3127 8667
rect 73 8613 87 8627
rect 333 8633 347 8647
rect 6833 8633 6847 8647
rect 7293 8633 7307 8647
rect 6233 8573 6247 8587
rect 6293 8573 6307 8587
rect 5933 8493 5947 8507
rect 6033 8493 6047 8507
rect 6533 8493 6547 8507
rect 6613 8493 6627 8507
rect 9353 8473 9367 8487
rect 9413 8473 9427 8487
rect 6913 8373 6927 8387
rect 7013 8373 7027 8387
rect 3593 8313 3607 8327
rect 3673 8313 3687 8327
rect 633 8153 647 8167
rect 6093 8093 6107 8107
rect 6193 8093 6207 8107
rect 6213 8073 6227 8087
rect 6273 8073 6287 8087
rect 5893 8053 5907 8067
rect 5953 8053 5967 8067
rect 5373 7993 5387 8007
rect 5413 7993 5427 8007
rect 5433 7993 5447 8007
rect 6113 7993 6127 8007
rect 6293 7993 6307 8007
rect 4713 7973 4727 7987
rect 4813 7973 4827 7987
rect 5193 7953 5207 7967
rect 5273 7953 5287 7967
rect 6493 7873 6507 7887
rect 6553 7873 6567 7887
rect 7193 7873 7207 7887
rect 7313 7873 7327 7887
rect 2433 7853 2447 7867
rect 2533 7853 2547 7867
rect 4073 7853 4087 7867
rect 4173 7853 4187 7867
rect 7953 7853 7967 7867
rect 8073 7853 8087 7867
rect 4773 7773 4787 7787
rect 4913 7773 4927 7787
rect 5913 7753 5927 7767
rect 6013 7753 6027 7767
rect 73 7713 87 7727
rect 93 7713 107 7727
rect 6653 7673 6667 7687
rect 8593 7673 8607 7687
rect 5713 7573 5727 7587
rect 5773 7573 5787 7587
rect 733 7533 747 7547
rect 893 7533 907 7547
rect 7413 7613 7427 7627
rect 7413 7533 7427 7547
rect 7513 7513 7527 7527
rect 7593 7513 7607 7527
rect 5513 7413 5527 7427
rect 5573 7413 5587 7427
rect 3733 7373 3747 7387
rect 3893 7373 3907 7387
rect 1833 7353 1847 7367
rect 7713 7333 7727 7347
rect 7873 7333 7887 7347
rect 7973 7313 7987 7327
rect 8033 7313 8047 7327
rect 2153 7293 2167 7307
rect 2313 7293 2327 7307
rect 1833 7273 1847 7287
rect 173 7213 187 7227
rect 10013 7213 10027 7227
rect 1133 7193 1147 7207
rect 4813 7133 4827 7147
rect 4953 7133 4967 7147
rect 5813 7033 5827 7047
rect 5953 7033 5967 7047
rect 5313 6993 5327 7007
rect 5433 6993 5447 7007
rect 8553 6913 8567 6927
rect 8593 6913 8607 6927
rect 4113 6873 4127 6887
rect 4293 6873 4307 6887
rect 7993 6873 8007 6887
rect 8053 6873 8067 6887
rect 1853 6853 1867 6867
rect 1893 6853 1907 6867
rect 4693 6833 4707 6847
rect 4813 6833 4827 6847
rect 3413 6813 3427 6827
rect 3533 6813 3547 6827
rect 773 6793 787 6807
rect 813 6793 827 6807
rect 553 6753 567 6767
rect 633 6753 647 6767
rect 2833 6713 2847 6727
rect 4553 6713 4567 6727
rect 6393 6713 6407 6727
rect 9513 6713 9527 6727
rect 10533 6713 10547 6727
rect 6753 6613 6767 6627
rect 6793 6613 6807 6627
rect 273 6427 287 6441
rect 433 6413 447 6427
rect 8333 6333 8347 6347
rect 8393 6333 8407 6347
rect 2193 6253 2207 6267
rect 2453 6253 2467 6267
rect 413 6233 427 6247
rect 1253 6233 1267 6247
rect 3973 6213 3987 6227
rect 4933 6233 4947 6247
rect 6733 6233 6747 6247
rect 6873 6233 6887 6247
rect 10873 6233 10887 6247
rect 10933 6233 10947 6247
rect 6953 6173 6967 6187
rect 7133 6173 7147 6187
rect 1273 6153 1287 6167
rect 1393 6153 1407 6167
rect 8073 6133 8087 6147
rect 8153 6133 8167 6147
rect 993 6093 1007 6107
rect 1093 6093 1107 6107
rect 5333 5973 5347 5987
rect 5373 5973 5387 5987
rect 11173 5893 11187 5907
rect 11213 5893 11227 5907
rect 1913 5793 1927 5807
rect 773 5753 787 5767
rect 933 5753 947 5767
rect 4293 5753 4307 5767
rect 6493 5753 6507 5767
rect 6773 5753 6787 5767
rect 7493 5753 7507 5767
rect 6113 5653 6127 5667
rect 6193 5653 6207 5667
rect 1633 5633 1647 5647
rect 1713 5633 1727 5647
rect 3033 5613 3047 5627
rect 3073 5613 3087 5627
rect 6473 5593 6487 5607
rect 6633 5593 6647 5607
rect 10033 5593 10047 5607
rect 10113 5593 10127 5607
rect 2993 5493 3007 5507
rect 3113 5493 3127 5507
rect 9853 5433 9867 5447
rect 9993 5433 10007 5447
rect 6133 5413 6147 5427
rect 6253 5413 6267 5427
rect 2733 5393 2747 5407
rect 2773 5393 2787 5407
rect 8893 5393 8907 5407
rect 8973 5393 8987 5407
rect 2313 5313 2327 5327
rect 73 5253 87 5267
rect 413 5273 427 5287
rect 3613 5273 3627 5287
rect 4933 5273 4947 5287
rect 5193 5273 5207 5287
rect 8253 5253 8267 5267
rect 8333 5253 8347 5267
rect 7773 5193 7787 5207
rect 7813 5193 7827 5207
rect 9673 5133 9687 5147
rect 9773 5133 9787 5147
rect 6853 5093 6867 5107
rect 6893 5093 6907 5107
rect 8433 4953 8447 4967
rect 8553 4953 8567 4967
rect 913 4813 927 4827
rect 1173 4813 1187 4827
rect 4073 4813 4087 4827
rect 73 4793 87 4807
rect 11093 4633 11107 4647
rect 11193 4633 11207 4647
rect 7773 4473 7787 4487
rect 7833 4473 7847 4487
rect 9213 4473 9227 4487
rect 9413 4493 9427 4507
rect 4173 4433 4187 4447
rect 4393 4433 4407 4447
rect 4733 4433 4747 4447
rect 4773 4433 4787 4447
rect 9613 4413 9627 4427
rect 9673 4413 9687 4427
rect 73 4313 87 4327
rect 873 4313 887 4327
rect 2153 4313 2167 4327
rect 2533 4313 2547 4327
rect 3333 4313 3347 4327
rect 3833 4313 3847 4327
rect 4653 4313 4667 4327
rect 5253 4313 5267 4327
rect 6213 4293 6227 4307
rect 3773 4173 3787 4187
rect 3953 4173 3967 4187
rect 5533 4153 5547 4167
rect 5573 4153 5587 4167
rect 9313 4153 9327 4167
rect 9353 4153 9367 4167
rect 6753 4053 6767 4067
rect 6813 4053 6827 4067
rect 11113 4013 11127 4027
rect 11173 4013 11187 4027
rect 7633 3953 7647 3967
rect 7753 3953 7767 3967
rect 10473 3933 10487 3947
rect 10513 3933 10527 3947
rect 5833 3893 5847 3907
rect 5873 3893 5887 3907
rect 73 3833 87 3847
rect 3273 3833 3287 3847
rect 1833 3813 1847 3827
rect 9113 3733 9127 3747
rect 9193 3733 9207 3747
rect 6673 3713 6687 3727
rect 6773 3713 6787 3727
rect 8553 3673 8567 3687
rect 8713 3673 8727 3687
rect 9273 3653 9287 3667
rect 9313 3653 9327 3667
rect 9013 3633 9027 3647
rect 9113 3633 9127 3647
rect 10133 3533 10147 3547
rect 10253 3533 10267 3547
rect 1133 3353 1147 3367
rect 1473 3353 1487 3367
rect 2453 3353 2467 3367
rect 673 3253 687 3267
rect 813 3253 827 3267
rect 6313 3253 6327 3267
rect 6353 3253 6367 3267
rect 6273 3213 6287 3227
rect 6373 3213 6387 3227
rect 10153 3213 10167 3227
rect 10233 3213 10247 3227
rect 10293 3193 10307 3207
rect 10353 3193 10367 3207
rect 7813 3073 7827 3087
rect 7893 3073 7907 3087
rect 6393 3053 6407 3067
rect 6433 3053 6447 3067
rect 8053 3053 8067 3067
rect 8133 3053 8147 3067
rect 10613 3053 10627 3067
rect 10793 3053 10807 3067
rect 3093 3013 3107 3027
rect 3193 3013 3207 3027
rect 9973 2993 9987 3007
rect 10093 2993 10107 3007
rect 10053 2973 10067 2987
rect 10093 2973 10107 2987
rect 10493 2953 10507 2967
rect 10553 2953 10567 2967
rect 1013 2873 1027 2887
rect 2553 2873 2567 2887
rect 3433 2873 3447 2887
rect 4873 2873 4887 2887
rect 5133 2873 5147 2887
rect 8587 2713 8601 2727
rect 8673 2713 8687 2727
rect 11093 2593 11107 2607
rect 11133 2593 11147 2607
rect 3113 2573 3127 2587
rect 3273 2573 3287 2587
rect 6353 2573 6367 2587
rect 6413 2573 6427 2587
rect 6653 2573 6667 2587
rect 6693 2573 6707 2587
rect 2073 2513 2087 2527
rect 2153 2513 2167 2527
rect 10633 2513 10647 2527
rect 10753 2513 10767 2527
rect 9933 2473 9947 2487
rect 9993 2473 10007 2487
rect 1753 2433 1767 2447
rect 573 2393 587 2407
rect 713 2393 727 2407
rect 3813 2393 3827 2407
rect 4033 2393 4047 2407
rect 9133 2213 9147 2227
rect 9253 2213 9267 2227
rect 2733 2093 2747 2107
rect 2793 2093 2807 2107
rect 6893 2093 6907 2107
rect 6953 2093 6967 2107
rect 8193 2093 8207 2107
rect 8353 2093 8367 2107
rect 9673 2093 9687 2107
rect 9713 2093 9727 2107
rect 10713 2093 10727 2107
rect 10773 2093 10787 2107
rect 11053 2093 11067 2107
rect 11133 2093 11147 2107
rect 9773 2013 9787 2027
rect 9853 2013 9867 2027
rect 493 1913 507 1927
rect 873 1913 887 1927
rect 2373 1913 2387 1927
rect 3913 1913 3927 1927
rect 4353 1913 4367 1927
rect 5193 1913 5207 1927
rect 8733 1793 8747 1807
rect 8873 1773 8887 1787
rect 5233 1433 5247 1447
rect 2953 1353 2967 1367
rect 3053 1353 3067 1367
rect 2333 1153 2347 1167
rect 2413 1153 2427 1167
rect 5773 1133 5787 1147
rect 5873 1133 5887 1147
rect 5913 1133 5927 1147
rect 6093 1133 6107 1147
rect 6293 1133 6307 1147
rect 6333 1133 6347 1147
rect 6533 1133 6547 1147
rect 6593 1133 6607 1147
rect 7673 1133 7687 1147
rect 7873 1133 7887 1147
rect 8273 1133 8287 1147
rect 8453 1133 8467 1147
rect 9493 1113 9507 1127
rect 9613 1113 9627 1127
rect 7413 953 7427 967
rect 9713 953 9727 967
rect 10233 953 10247 967
rect 8393 853 8407 867
rect 8593 813 8607 827
rect 8633 813 8647 827
rect 6347 793 6361 807
rect 6453 793 6467 807
rect 8393 793 8407 807
rect 10193 793 10207 807
rect 10253 793 10267 807
rect 8693 653 8707 667
rect 8853 653 8867 667
rect 9533 573 9547 587
rect 9593 573 9607 587
rect 10513 493 10527 507
rect 5833 473 5847 487
rect 9133 473 9147 487
rect 9713 473 9727 487
rect 8353 313 8367 327
rect 8513 313 8527 327
rect 5813 153 5827 167
rect 6013 153 6027 167
rect 10573 113 10587 127
rect 10633 113 10647 127
<< metal2 >>
rect 3936 11336 3963 11343
rect 1196 11216 1223 11223
rect 36 10936 63 10943
rect 56 10507 63 10936
rect 196 10927 203 11183
rect 336 11147 343 11183
rect 616 11163 623 11213
rect 936 11187 943 11213
rect 1196 11187 1203 11216
rect 2456 11216 2483 11223
rect 596 11156 623 11163
rect 76 10907 83 10923
rect 456 10916 483 10923
rect 476 10867 483 10916
rect 536 10907 543 11033
rect 176 10716 203 10723
rect 236 10716 243 10733
rect 176 10687 183 10716
rect 16 10207 23 10233
rect 56 9987 63 10493
rect 176 10436 203 10443
rect 176 10407 183 10436
rect 36 9187 43 9243
rect 56 9187 63 9973
rect 156 9943 163 10353
rect 216 10347 223 10403
rect 196 10236 203 10273
rect 236 10236 263 10243
rect 256 10167 263 10236
rect 156 9936 183 9943
rect 216 9887 223 9943
rect 156 9487 163 9733
rect 236 9723 243 10153
rect 276 9927 283 10233
rect 176 9647 183 9723
rect 216 9716 243 9723
rect 76 9256 103 9263
rect 96 9127 103 9256
rect 156 9007 163 9113
rect 176 8763 183 9633
rect 236 9476 243 9633
rect 296 9587 303 9963
rect 316 9867 323 10733
rect 456 10716 463 10733
rect 516 10667 523 10713
rect 376 10436 383 10533
rect 436 10283 443 10423
rect 416 10276 443 10283
rect 216 9363 223 9463
rect 196 9356 223 9363
rect 196 9296 203 9356
rect 276 9023 283 9173
rect 356 9163 363 9853
rect 336 9156 363 9163
rect 276 9016 303 9023
rect 236 8867 243 8983
rect 256 8763 263 8813
rect 296 8763 303 9016
rect 336 8827 343 9156
rect 396 9103 403 10273
rect 416 10227 423 10276
rect 456 10263 463 10453
rect 516 10447 523 10653
rect 436 10256 463 10263
rect 436 10236 443 10256
rect 516 10247 523 10433
rect 496 10127 503 10223
rect 536 10207 543 10733
rect 556 9727 563 9873
rect 416 9647 423 9723
rect 436 9523 443 9693
rect 416 9516 443 9523
rect 416 9483 423 9516
rect 416 9476 443 9483
rect 476 9476 483 9633
rect 516 9463 523 9473
rect 456 9303 463 9463
rect 496 9456 523 9463
rect 436 9296 463 9303
rect 396 9096 423 9103
rect 416 8823 423 9096
rect 436 9007 443 9296
rect 476 9263 483 9313
rect 456 9256 483 9263
rect 576 9107 583 11133
rect 596 10827 603 11156
rect 636 10903 643 11173
rect 956 11167 963 11183
rect 636 10896 663 10903
rect 676 10716 683 10873
rect 656 10687 663 10703
rect 716 10687 723 10903
rect 616 10427 623 10443
rect 636 10347 643 10463
rect 696 10447 703 10513
rect 736 10507 743 10953
rect 736 10456 743 10493
rect 756 10427 763 10933
rect 876 10683 883 10853
rect 896 10827 903 10903
rect 936 10887 943 10903
rect 916 10727 923 10883
rect 956 10787 963 11153
rect 996 10887 1003 11173
rect 1056 10847 1063 10913
rect 876 10676 903 10683
rect 696 10236 723 10243
rect 736 10236 743 10313
rect 596 10047 603 10233
rect 616 10167 623 10233
rect 596 9267 603 9953
rect 636 9947 643 10113
rect 676 9956 703 9963
rect 636 9743 643 9933
rect 696 9847 703 9956
rect 676 9776 683 9833
rect 716 9767 723 10236
rect 636 9736 663 9743
rect 636 9296 643 9313
rect 656 9307 663 9736
rect 676 9287 683 9453
rect 716 9347 723 9443
rect 676 9263 683 9273
rect 656 9256 683 9263
rect 616 8987 623 9003
rect 696 8996 703 9333
rect 716 9187 723 9243
rect 736 9143 743 10193
rect 776 10067 783 10443
rect 876 10267 883 10676
rect 936 10667 943 10683
rect 1056 10443 1063 10833
rect 1176 10696 1183 10773
rect 1196 10747 1203 10903
rect 1336 10827 1343 11213
rect 1356 10923 1363 11213
rect 1436 11196 1443 11213
rect 1496 11196 1523 11203
rect 1356 10916 1383 10923
rect 1396 10807 1403 10903
rect 1216 10696 1223 10713
rect 1396 10696 1403 10713
rect 1436 10696 1443 10773
rect 1456 10747 1463 10913
rect 1156 10547 1163 10683
rect 1416 10676 1423 10693
rect 1056 10436 1083 10443
rect 1156 10436 1163 10493
rect 896 10387 903 10403
rect 976 10256 983 10333
rect 936 10236 963 10243
rect 996 10236 1023 10243
rect 916 9907 923 9943
rect 936 9927 943 10236
rect 1016 9987 1023 10236
rect 1076 9967 1083 10436
rect 1176 10236 1183 10273
rect 1236 10236 1243 10453
rect 1376 10447 1383 10673
rect 1456 10447 1463 10683
rect 1496 10407 1503 10693
rect 1516 10667 1523 11196
rect 1556 10907 1563 11033
rect 1616 10923 1623 11213
rect 1736 11196 1763 11203
rect 1796 11196 1803 11213
rect 1736 11187 1743 11196
rect 1816 11176 1823 11193
rect 1876 10967 1883 11153
rect 1736 10936 1743 10953
rect 1616 10916 1643 10923
rect 1396 10236 1423 10243
rect 1456 10236 1483 10243
rect 1116 9976 1143 9983
rect 1176 9976 1183 10033
rect 1116 9807 1123 9976
rect 1196 9967 1203 10203
rect 1396 10187 1403 10236
rect 1476 10067 1483 10236
rect 916 9723 923 9753
rect 856 9647 863 9723
rect 896 9716 923 9723
rect 896 9483 903 9693
rect 896 9476 923 9483
rect 956 9476 963 9633
rect 856 9447 863 9473
rect 936 9367 943 9463
rect 876 9296 883 9353
rect 756 9256 783 9263
rect 716 9136 743 9143
rect 416 8816 443 8823
rect 616 8783 623 8973
rect 716 8807 723 9136
rect 776 9127 783 9256
rect 316 8776 343 8783
rect 176 8756 203 8763
rect 236 8756 263 8763
rect 276 8756 303 8763
rect 76 8296 83 8613
rect 176 8523 183 8733
rect 196 8567 203 8756
rect 176 8516 203 8523
rect 236 8516 243 8553
rect 276 8507 283 8756
rect 336 8647 343 8776
rect 596 8776 623 8783
rect 216 8403 223 8503
rect 256 8427 263 8503
rect 496 8487 503 8503
rect 196 8396 223 8403
rect 196 8336 203 8396
rect 376 8296 383 8313
rect 476 8303 483 8333
rect 456 8296 483 8303
rect 36 8087 43 8283
rect 36 8056 43 8073
rect 56 7583 63 8073
rect 396 8043 403 8053
rect 76 7727 83 8043
rect 376 8036 403 8043
rect 456 8036 483 8043
rect 196 7836 203 8003
rect 216 7767 223 7823
rect 36 7576 63 7583
rect 56 7107 63 7576
rect 96 7563 103 7713
rect 76 7556 103 7563
rect 256 7356 283 7363
rect 36 7096 53 7103
rect 56 6763 63 7093
rect 96 7047 103 7353
rect 236 7327 243 7343
rect 276 7307 283 7356
rect 296 7327 303 7353
rect 176 7087 183 7213
rect 256 6843 263 6893
rect 36 6756 63 6763
rect 36 6616 43 6756
rect 196 6747 203 6843
rect 236 6836 263 6843
rect 76 6247 83 6603
rect 196 6396 203 6563
rect 76 5896 83 6233
rect 236 6116 243 6173
rect 176 5943 183 6103
rect 256 6087 263 6113
rect 216 6067 223 6083
rect 276 6067 283 6413
rect 176 5936 203 5943
rect 36 5663 43 5873
rect 36 5656 63 5663
rect 16 4967 23 5013
rect 56 4923 63 5656
rect 76 5267 83 5643
rect 356 5627 363 8013
rect 396 7563 403 8036
rect 476 8003 483 8036
rect 496 8027 503 8473
rect 596 8327 603 8776
rect 676 8536 683 8553
rect 716 8536 723 8793
rect 736 8787 743 8893
rect 676 8303 683 8413
rect 656 8296 683 8303
rect 636 8167 643 8293
rect 636 8047 643 8153
rect 676 8036 683 8093
rect 716 8087 723 8283
rect 776 8107 783 9093
rect 856 8803 863 9293
rect 1036 9256 1063 9263
rect 896 8907 903 8963
rect 856 8796 883 8803
rect 896 8767 903 8783
rect 956 8767 963 9013
rect 1036 8987 1043 9256
rect 1076 9007 1083 9793
rect 1096 9736 1103 9773
rect 1136 9303 1143 9733
rect 1196 9427 1203 9443
rect 1116 9296 1143 9303
rect 1116 9027 1123 9296
rect 1196 9267 1203 9413
rect 1116 8996 1123 9013
rect 1076 8983 1083 8993
rect 1156 8987 1163 9003
rect 1076 8976 1103 8983
rect 1136 8827 1143 8983
rect 1156 8796 1163 8933
rect 1216 8927 1223 9973
rect 1136 8767 1143 8783
rect 956 8516 963 8553
rect 1156 8516 1163 8533
rect 1196 8507 1203 8523
rect 936 8407 943 8503
rect 976 8407 983 8503
rect 1136 8427 1143 8503
rect 876 8336 883 8393
rect 1056 8307 1063 8313
rect 1096 8287 1103 8333
rect 1156 8303 1163 8333
rect 1136 8296 1163 8303
rect 476 7996 503 8003
rect 376 7556 403 7563
rect 396 7087 403 7556
rect 416 7703 423 7833
rect 436 7703 443 7793
rect 416 7696 443 7703
rect 416 7307 423 7696
rect 476 7643 483 7803
rect 496 7643 503 7996
rect 636 7836 643 8013
rect 716 7987 723 8073
rect 816 8036 823 8053
rect 676 7836 683 7973
rect 476 7636 503 7643
rect 496 7567 503 7636
rect 716 7576 743 7583
rect 456 7556 483 7563
rect 476 7543 483 7556
rect 476 7536 503 7543
rect 436 7307 443 7323
rect 476 7303 483 7323
rect 456 7296 483 7303
rect 376 7076 393 7083
rect 456 7083 463 7296
rect 496 7263 503 7536
rect 436 7076 463 7083
rect 476 7256 503 7263
rect 396 6603 403 7073
rect 436 7043 443 7076
rect 436 7036 463 7043
rect 456 6883 463 7036
rect 476 6907 483 7256
rect 496 6887 503 7113
rect 456 6876 483 6883
rect 436 6856 443 6873
rect 476 6856 483 6876
rect 416 6607 423 6843
rect 536 6663 543 7293
rect 556 7127 563 7533
rect 556 6767 563 7083
rect 576 6987 583 7333
rect 636 7203 643 7573
rect 696 7547 703 7563
rect 736 7547 743 7576
rect 676 7356 683 7513
rect 696 7307 703 7343
rect 636 7196 663 7203
rect 536 6656 563 6663
rect 376 6596 403 6603
rect 376 6567 383 6596
rect 456 6596 483 6603
rect 376 5927 383 6553
rect 476 6427 483 6596
rect 436 6396 443 6413
rect 476 6396 483 6413
rect 407 6236 413 6243
rect 496 6103 503 6393
rect 436 6067 443 6103
rect 476 6096 503 6103
rect 376 5896 383 5913
rect 396 5643 403 5913
rect 376 5636 403 5643
rect 176 5596 203 5603
rect 176 5436 183 5596
rect 436 5487 443 6053
rect 476 5903 483 6096
rect 456 5896 483 5903
rect 536 5703 543 6133
rect 516 5696 543 5703
rect 456 5636 463 5653
rect 216 5456 223 5473
rect 276 5427 283 5453
rect 436 5436 443 5473
rect 476 5436 483 5653
rect 236 5416 263 5423
rect 76 4936 83 5253
rect 176 5147 183 5163
rect 256 5143 263 5416
rect 196 4976 203 5143
rect 236 5136 263 5143
rect 236 5047 243 5136
rect 356 4936 383 4943
rect 36 4916 63 4923
rect 76 4456 83 4793
rect 216 4676 223 4793
rect 196 4496 203 4663
rect 356 4647 363 4936
rect 396 4707 403 5153
rect 416 5127 423 5273
rect 516 5167 523 5696
rect 556 5467 563 6656
rect 616 6627 623 6853
rect 656 6847 663 7196
rect 676 7027 683 7043
rect 676 6856 683 6893
rect 696 6876 703 6973
rect 816 6807 823 7093
rect 636 6587 643 6753
rect 716 6616 723 6653
rect 776 6616 783 6793
rect 696 6583 703 6603
rect 816 6587 823 6603
rect 696 6576 723 6583
rect 676 6396 683 6413
rect 716 6396 723 6576
rect 756 6396 763 6413
rect 696 6367 703 6383
rect 656 6087 663 6123
rect 696 6116 703 6133
rect 736 6087 743 6383
rect 576 5907 583 6073
rect 776 5936 783 6033
rect 596 5896 603 5913
rect 776 5767 783 5893
rect 536 5176 543 5273
rect 416 4807 423 5033
rect 436 4967 443 5163
rect 496 5067 503 5143
rect 476 4943 483 4953
rect 456 4936 483 4943
rect 416 4696 443 4703
rect 476 4696 483 4713
rect 356 4463 363 4633
rect 356 4456 383 4463
rect 56 3963 63 4433
rect 76 3976 83 4313
rect 196 4187 203 4203
rect 216 4083 223 4183
rect 256 4127 263 4183
rect 356 4147 363 4456
rect 396 4207 403 4693
rect 416 4667 423 4696
rect 516 4687 523 5153
rect 576 5127 583 5163
rect 416 4427 423 4653
rect 516 4487 523 4673
rect 456 4163 463 4203
rect 496 4196 503 4473
rect 536 4183 543 5053
rect 556 4467 563 4713
rect 596 4667 603 5453
rect 656 5443 663 5643
rect 656 5436 683 5443
rect 636 5416 663 5423
rect 636 5267 643 5416
rect 676 5396 683 5436
rect 796 5407 803 6273
rect 836 6267 843 8093
rect 876 8056 883 8073
rect 936 7747 943 7803
rect 856 6967 863 7073
rect 876 6847 883 7553
rect 896 7547 903 7563
rect 916 7336 923 7583
rect 956 7576 963 7653
rect 1016 7576 1023 8073
rect 1196 8043 1203 8293
rect 1236 8207 1243 9833
rect 1256 9747 1263 9993
rect 1356 9807 1363 9943
rect 1396 9907 1403 9943
rect 1496 9927 1503 10393
rect 1396 9776 1403 9793
rect 1356 9756 1363 9773
rect 1376 9727 1383 9743
rect 1376 9476 1383 9493
rect 1336 9463 1343 9473
rect 1336 9456 1363 9463
rect 1316 9243 1323 9433
rect 1336 9276 1343 9456
rect 1376 9276 1383 9293
rect 1316 9236 1343 9243
rect 1196 8036 1223 8043
rect 1036 7947 1043 8003
rect 1216 7987 1223 8036
rect 1256 8027 1263 8773
rect 1276 8527 1283 8993
rect 1316 8787 1323 9213
rect 1336 8796 1343 9236
rect 1356 9227 1363 9263
rect 1436 9007 1443 9733
rect 1456 9487 1463 9513
rect 1476 9467 1483 9713
rect 1416 8887 1423 8963
rect 1076 7836 1103 7843
rect 1136 7836 1143 7933
rect 1316 7867 1323 8753
rect 1356 8647 1363 8773
rect 1476 8516 1483 8953
rect 1376 8303 1383 8393
rect 1456 8327 1463 8483
rect 1356 8296 1383 8303
rect 1496 8036 1503 8993
rect 1536 8987 1543 10893
rect 1656 10867 1663 10903
rect 1696 10767 1703 10903
rect 1716 10887 1723 10913
rect 1636 10487 1643 10713
rect 1656 10443 1663 10753
rect 1736 10727 1743 10793
rect 1716 10667 1723 10703
rect 1716 10487 1723 10653
rect 1636 10436 1663 10443
rect 1616 9756 1623 9853
rect 1636 9736 1663 9743
rect 1596 9487 1603 9493
rect 1636 9487 1643 9553
rect 1656 9507 1663 9736
rect 1596 8547 1603 9473
rect 1676 9467 1683 9483
rect 1616 9447 1623 9463
rect 1636 9296 1643 9433
rect 1616 9276 1623 9293
rect 1656 9276 1663 9293
rect 1696 9007 1703 9713
rect 1616 8963 1623 9003
rect 1616 8956 1643 8963
rect 1636 8816 1643 8956
rect 1676 8947 1683 8983
rect 1676 8607 1683 8933
rect 1696 8727 1703 8993
rect 1716 8963 1723 9933
rect 1756 9787 1763 10913
rect 1776 10907 1783 10923
rect 1796 10443 1803 10473
rect 1856 10447 1863 10713
rect 1876 10467 1883 10953
rect 1896 10927 1903 11213
rect 2456 11187 2463 11216
rect 2716 11196 2723 11213
rect 2216 11176 2243 11183
rect 2196 11047 2203 11173
rect 2236 11147 2243 11176
rect 2736 11176 2743 11233
rect 2936 11216 2963 11223
rect 1896 10867 1903 10883
rect 1916 10736 1923 10813
rect 2056 10727 2063 10873
rect 2076 10847 2083 10923
rect 1936 10716 1963 10723
rect 1796 10436 1823 10443
rect 1896 10407 1903 10433
rect 1856 10256 1863 10393
rect 1736 8987 1743 9253
rect 1716 8956 1743 8963
rect 1576 8447 1583 8513
rect 1656 8507 1663 8523
rect 1696 8516 1703 8713
rect 1676 8467 1683 8503
rect 1556 8316 1563 8413
rect 1576 8336 1583 8433
rect 1596 8316 1603 8373
rect 1076 7807 1083 7836
rect 1356 7836 1363 7853
rect 1436 7836 1443 7853
rect 1116 7787 1123 7823
rect 896 7087 903 7323
rect 936 6876 943 6973
rect 956 6856 963 7073
rect 976 7007 983 7353
rect 1056 7193 1063 7563
rect 1076 7347 1083 7773
rect 1336 7767 1343 7833
rect 1376 7807 1383 7823
rect 1456 7807 1463 7833
rect 1176 7356 1183 7523
rect 916 6507 923 6833
rect 936 6527 943 6563
rect 976 6396 983 6493
rect 1016 6396 1023 6413
rect 956 6367 963 6383
rect 996 6167 1003 6383
rect 936 6047 943 6103
rect 976 6096 993 6103
rect 956 5947 963 6033
rect 936 5863 943 5873
rect 916 5856 943 5863
rect 916 5623 923 5856
rect 936 5647 943 5753
rect 1016 5667 1023 6353
rect 896 5616 923 5623
rect 636 4987 643 5073
rect 676 4956 683 5353
rect 656 4883 663 4943
rect 636 4876 663 4883
rect 636 4463 643 4876
rect 656 4867 663 4876
rect 676 4696 683 4913
rect 696 4487 703 4683
rect 716 4607 723 4703
rect 736 4467 743 4683
rect 636 4456 663 4463
rect 656 4247 663 4456
rect 516 4176 543 4183
rect 456 4156 483 4163
rect 196 4076 223 4083
rect 196 4016 203 4076
rect 356 3983 363 4133
rect 356 3976 383 3983
rect 36 3956 63 3963
rect 56 3483 63 3956
rect 76 3496 83 3833
rect 236 3716 243 3773
rect 176 3623 183 3703
rect 256 3687 263 3713
rect 216 3667 223 3683
rect 176 3616 203 3623
rect 196 3536 203 3616
rect 356 3503 363 3976
rect 396 3787 403 4113
rect 476 3987 483 4156
rect 656 4047 663 4233
rect 716 4227 723 4433
rect 716 4183 723 4213
rect 756 4183 763 4713
rect 776 4676 783 4933
rect 816 4387 823 4913
rect 836 4407 843 4953
rect 856 4907 863 5613
rect 916 5527 923 5616
rect 916 5436 923 5453
rect 856 4727 863 4893
rect 856 4647 863 4683
rect 876 4647 883 5153
rect 896 5127 903 5433
rect 936 5407 943 5423
rect 956 5156 963 5353
rect 1016 5287 1023 5513
rect 996 5067 1003 5253
rect 1016 5176 1023 5273
rect 956 4956 963 4973
rect 996 4956 1003 5053
rect 976 4927 983 4943
rect 1036 4927 1043 6493
rect 1096 6387 1103 6993
rect 1116 6927 1123 7333
rect 1136 7047 1143 7179
rect 1196 7087 1203 7293
rect 1156 6987 1163 7083
rect 1176 7027 1183 7063
rect 1127 6876 1143 6883
rect 1116 6783 1123 6873
rect 1196 6856 1203 6933
rect 1236 6867 1243 7073
rect 1276 7067 1283 7173
rect 1116 6776 1143 6783
rect 1116 6567 1123 6603
rect 1136 6407 1143 6776
rect 1156 6507 1163 6853
rect 1096 6107 1103 6373
rect 1136 5916 1143 6393
rect 1216 6247 1223 6383
rect 1256 6376 1263 6593
rect 1176 6147 1183 6233
rect 1176 6116 1183 6133
rect 1236 6123 1243 6153
rect 1216 6116 1243 6123
rect 1096 5587 1103 5913
rect 1156 5883 1163 6093
rect 1256 5896 1263 6233
rect 1276 6187 1283 7053
rect 1296 7047 1303 7083
rect 1316 6587 1323 7373
rect 1336 7187 1343 7753
rect 1476 7747 1483 8033
rect 1576 8007 1583 8033
rect 1656 8027 1663 8393
rect 1476 7567 1483 7733
rect 1356 7307 1363 7563
rect 1436 7556 1463 7563
rect 1456 7387 1463 7556
rect 1376 7376 1423 7383
rect 1376 7347 1383 7376
rect 1436 7356 1443 7373
rect 1396 6967 1403 7293
rect 1496 7187 1503 7353
rect 1516 7307 1523 8003
rect 1616 7836 1643 7843
rect 1616 7807 1623 7836
rect 1676 7576 1703 7583
rect 1656 7547 1663 7553
rect 1416 6983 1423 7043
rect 1416 6976 1443 6983
rect 1436 6876 1443 6976
rect 1596 6967 1603 7083
rect 1416 6856 1423 6873
rect 1456 6687 1463 6853
rect 1376 6367 1383 6613
rect 1456 6596 1463 6613
rect 1396 6567 1403 6583
rect 1396 6427 1403 6553
rect 1436 6547 1443 6583
rect 1476 6396 1483 6513
rect 1516 6487 1523 6913
rect 1516 6396 1523 6473
rect 1456 6376 1463 6393
rect 1276 6167 1283 6173
rect 1276 5907 1283 6133
rect 1356 5887 1363 6133
rect 1396 6103 1403 6153
rect 1496 6127 1503 6383
rect 1536 6347 1543 6873
rect 1576 6547 1583 6873
rect 1476 6107 1483 6123
rect 1536 6116 1543 6153
rect 1596 6123 1603 6953
rect 1616 6747 1623 7313
rect 1636 6407 1643 7173
rect 1656 7083 1663 7323
rect 1656 7076 1683 7083
rect 1656 6947 1663 7076
rect 1696 6907 1703 7576
rect 1716 6967 1723 8503
rect 1736 8467 1743 8956
rect 1756 8767 1763 9773
rect 1756 8407 1763 8533
rect 1776 8467 1783 10253
rect 1816 10236 1843 10243
rect 1876 10236 1883 10273
rect 1816 10227 1823 10236
rect 1796 9127 1803 9933
rect 1816 9767 1823 10213
rect 1836 9867 1843 9963
rect 1876 9956 1883 9993
rect 1856 9887 1863 9943
rect 1916 9927 1923 10413
rect 1876 9756 1883 9913
rect 1816 9363 1823 9753
rect 1836 9736 1863 9743
rect 1836 9447 1843 9736
rect 1896 9727 1903 9743
rect 1936 9723 1943 10453
rect 1956 10427 1963 10716
rect 1976 9747 1983 9833
rect 1996 9767 2003 10593
rect 2056 10443 2063 10713
rect 2036 10436 2063 10443
rect 2036 9947 2043 10436
rect 2076 10367 2083 10403
rect 2056 10236 2083 10243
rect 2056 10207 2063 10236
rect 2076 9976 2083 10053
rect 2096 10027 2103 10833
rect 2116 10367 2123 10913
rect 2216 10767 2223 10873
rect 2236 10847 2243 11133
rect 2376 10887 2383 10923
rect 2176 10716 2203 10723
rect 2196 10287 2203 10716
rect 2216 10423 2223 10753
rect 2296 10436 2303 10453
rect 2216 10416 2243 10423
rect 2276 10387 2283 10423
rect 2116 10236 2143 10243
rect 2136 9947 2143 10236
rect 1996 9736 2023 9743
rect 1936 9716 1963 9723
rect 2016 9607 2023 9736
rect 1876 9476 1883 9493
rect 2156 9476 2163 9493
rect 1816 9356 1843 9363
rect 1816 9107 1823 9333
rect 1836 9276 1843 9356
rect 1856 9347 1863 9463
rect 1936 9447 1943 9463
rect 1876 9276 1883 9293
rect 1856 9127 1863 9263
rect 1836 8796 1843 9113
rect 1856 9016 1863 9093
rect 1876 8823 1883 9003
rect 1876 8816 1893 8823
rect 1856 8767 1863 8783
rect 1896 8776 1903 8813
rect 1916 8767 1923 9113
rect 1936 8967 1943 9433
rect 1976 8787 1983 9473
rect 2076 9427 2083 9453
rect 2216 9447 2223 9463
rect 2076 9243 2083 9413
rect 2076 9236 2103 9243
rect 2136 9027 2143 9243
rect 2116 8996 2123 9013
rect 2136 8847 2143 8963
rect 2196 8947 2203 9253
rect 2156 8816 2163 8833
rect 2136 8767 2143 8783
rect 1756 8036 1763 8393
rect 1776 8307 1783 8333
rect 1796 8316 1803 8333
rect 1836 8316 1843 8533
rect 1976 8487 1983 8503
rect 2076 8347 2083 8573
rect 2136 8503 2143 8753
rect 2176 8667 2183 8773
rect 2216 8767 2223 9013
rect 2236 9007 2243 9473
rect 2256 9467 2263 9513
rect 2136 8496 2163 8503
rect 2156 8367 2163 8496
rect 2196 8447 2203 8503
rect 2076 8316 2083 8333
rect 2156 8316 2183 8323
rect 1816 8287 1823 8303
rect 1856 8287 1863 8303
rect 1816 8043 1823 8053
rect 1796 8036 1823 8043
rect 1776 8007 1783 8023
rect 1736 7087 1743 7553
rect 1756 7507 1763 7793
rect 1656 6856 1663 6893
rect 1696 6856 1703 6873
rect 1676 6836 1683 6853
rect 1736 6843 1743 6973
rect 1716 6836 1743 6843
rect 1776 6627 1783 7973
rect 1796 7107 1803 7573
rect 1836 7567 1843 7853
rect 1856 7836 1863 8033
rect 1936 7787 1943 8313
rect 2136 8287 2143 8293
rect 1816 7103 1823 7353
rect 1836 7336 1843 7353
rect 1876 7336 1883 7353
rect 1856 7316 1863 7333
rect 1836 7127 1843 7273
rect 1916 7147 1923 7543
rect 1956 7507 1963 7543
rect 1976 7527 1983 7553
rect 1996 7347 2003 8003
rect 2176 7987 2183 8316
rect 2236 8247 2243 8993
rect 2256 8307 2263 8833
rect 2276 8727 2283 10353
rect 2336 10267 2343 10433
rect 2396 10427 2403 10903
rect 2416 10527 2423 10703
rect 2436 10687 2443 10903
rect 2456 10747 2463 10913
rect 2776 10907 2783 11193
rect 2936 11183 2943 11216
rect 3676 11216 3703 11223
rect 3956 11216 3963 11336
rect 4136 11307 4143 11343
rect 4376 11307 4383 11343
rect 2816 11176 2843 11183
rect 2936 11176 2963 11183
rect 2816 11047 2823 11176
rect 2636 10867 2643 10903
rect 2456 10716 2463 10733
rect 2516 10716 2543 10723
rect 2536 10687 2543 10716
rect 2516 10423 2523 10453
rect 2596 10436 2603 10853
rect 2676 10707 2683 10903
rect 2736 10736 2743 10853
rect 2716 10716 2723 10733
rect 2756 10716 2763 10753
rect 2616 10467 2623 10493
rect 2516 10416 2543 10423
rect 2296 10236 2303 10253
rect 2316 10207 2323 10223
rect 2296 9736 2303 10013
rect 2316 10007 2323 10193
rect 2376 10067 2383 10233
rect 2356 9967 2363 9973
rect 2336 9787 2343 9943
rect 2376 9867 2383 9943
rect 2396 9647 2403 9953
rect 2396 9327 2403 9473
rect 2416 9427 2423 9493
rect 2496 9427 2503 9463
rect 2036 7856 2063 7863
rect 2036 7807 2043 7856
rect 2076 7836 2083 7873
rect 2236 7867 2243 8003
rect 2276 7887 2283 8653
rect 2296 8387 2303 9193
rect 2396 9016 2403 9313
rect 2436 9187 2443 9263
rect 2496 9027 2503 9413
rect 2376 8796 2383 8913
rect 2396 8747 2403 8783
rect 2396 8503 2403 8633
rect 2436 8516 2443 8573
rect 2396 8496 2423 8503
rect 2296 8027 2303 8373
rect 2356 8347 2363 8393
rect 2356 8316 2363 8333
rect 2316 8027 2323 8053
rect 2436 7867 2443 8353
rect 2456 8023 2463 8773
rect 2476 8167 2483 8793
rect 2496 8056 2503 8313
rect 2516 8307 2523 9473
rect 2536 9287 2543 10253
rect 2576 10236 2583 10253
rect 2616 10223 2623 10453
rect 2676 10407 2683 10693
rect 2736 10436 2763 10443
rect 2736 10287 2743 10436
rect 2796 10423 2803 10913
rect 2836 10887 2843 10933
rect 2916 10916 2923 10933
rect 2956 10907 2963 11176
rect 3116 11176 3143 11183
rect 3116 11147 3123 11176
rect 3156 10947 3163 11113
rect 3196 10927 3203 11033
rect 2856 10867 2863 10893
rect 2936 10847 2943 10903
rect 3096 10887 3103 10913
rect 3096 10747 3103 10873
rect 3116 10767 3123 10903
rect 3176 10867 3183 10923
rect 3196 10847 3203 10873
rect 3216 10867 3223 11183
rect 3236 10936 3263 10943
rect 2816 10436 2823 10693
rect 2916 10687 2923 10713
rect 2996 10696 3023 10703
rect 2776 10416 2803 10423
rect 2776 10347 2783 10416
rect 2836 10327 2843 10423
rect 2596 10216 2623 10223
rect 2556 9956 2563 10213
rect 2576 9916 2603 9923
rect 2596 9736 2603 9916
rect 2616 9887 2623 10216
rect 2736 10167 2743 10273
rect 2836 10236 2843 10293
rect 2916 10227 2923 10413
rect 3016 10407 3023 10696
rect 3116 10567 3123 10753
rect 3216 10736 3243 10743
rect 3196 10587 3203 10703
rect 3236 10607 3243 10736
rect 3036 10403 3043 10433
rect 3096 10407 3103 10423
rect 3136 10407 3143 10423
rect 3036 10396 3063 10403
rect 2756 10216 2783 10223
rect 2576 9467 2583 9723
rect 2636 9547 2643 9853
rect 2656 9727 2663 9753
rect 2636 9463 2643 9533
rect 2676 9476 2683 9553
rect 2716 9467 2723 9483
rect 2636 9456 2663 9463
rect 2696 9443 2703 9463
rect 2736 9443 2743 9953
rect 2756 9943 2763 10216
rect 2816 10207 2823 10223
rect 2816 9967 2823 10193
rect 2836 9956 2863 9963
rect 2756 9936 2783 9943
rect 2696 9436 2743 9443
rect 2576 9267 2583 9293
rect 2656 9276 2663 9393
rect 2556 8787 2563 8853
rect 2576 8767 2583 8993
rect 2596 8867 2603 9023
rect 2636 9016 2643 9263
rect 2676 9247 2683 9253
rect 2616 8987 2623 9003
rect 2596 8796 2603 8853
rect 2656 8796 2663 8993
rect 2576 8296 2583 8713
rect 2616 8516 2623 8553
rect 2596 8447 2603 8483
rect 2636 8407 2643 8753
rect 2596 8316 2603 8373
rect 2636 8316 2663 8323
rect 2456 8016 2483 8023
rect 2336 7836 2363 7843
rect 2336 7827 2343 7836
rect 2096 7376 2103 7533
rect 2176 7527 2183 7543
rect 2116 7356 2123 7453
rect 2156 7307 2163 7513
rect 2116 7187 2123 7293
rect 1816 7096 1843 7103
rect 1716 6596 1723 6613
rect 1816 6596 1823 6633
rect 1696 6467 1703 6583
rect 1776 6567 1783 6583
rect 1716 6407 1723 6433
rect 1756 6396 1763 6453
rect 1596 6116 1623 6123
rect 1396 6096 1423 6103
rect 1456 6087 1463 6103
rect 1136 5876 1163 5883
rect 1136 5623 1143 5876
rect 1196 5656 1203 5873
rect 1516 5867 1523 6113
rect 1556 5896 1563 5953
rect 1116 5616 1143 5623
rect 1116 5267 1123 5616
rect 1156 5587 1163 5623
rect 1216 5403 1223 5453
rect 1156 5367 1163 5403
rect 1196 5396 1223 5403
rect 1216 5387 1223 5396
rect 1056 4827 1063 5163
rect 1256 5047 1263 5053
rect 927 4816 933 4823
rect 1136 4647 1143 4953
rect 1196 4936 1203 4973
rect 1256 4956 1263 5033
rect 1176 4683 1183 4813
rect 1196 4696 1223 4703
rect 1156 4676 1183 4683
rect 1216 4627 1223 4696
rect 856 4463 863 4593
rect 1216 4507 1223 4613
rect 856 4456 883 4463
rect 916 4456 923 4473
rect 696 4176 723 4183
rect 736 4176 763 4183
rect 496 3707 503 3993
rect 416 3507 423 3693
rect 456 3687 463 3703
rect 456 3667 463 3673
rect 356 3496 383 3503
rect 36 3476 63 3483
rect 356 3387 363 3496
rect 176 3267 183 3293
rect 176 3236 183 3253
rect 316 3236 323 3373
rect 216 3016 223 3233
rect 196 2767 203 3003
rect 236 2787 243 2993
rect 176 2527 183 2743
rect 216 2727 223 2743
rect 276 2547 283 3013
rect 376 2763 383 3453
rect 536 3247 543 3713
rect 396 3027 403 3213
rect 416 3027 423 3233
rect 436 3016 443 3053
rect 476 3003 483 3173
rect 456 2996 483 3003
rect 456 2776 463 2953
rect 376 2756 403 2763
rect 396 2587 403 2756
rect 596 2727 603 3753
rect 616 3067 623 4013
rect 636 3227 643 3953
rect 656 3667 663 4033
rect 696 3976 703 4153
rect 716 3707 723 3953
rect 736 3767 743 4176
rect 816 4167 823 4373
rect 836 3923 843 4393
rect 856 4067 863 4456
rect 936 4427 943 4443
rect 876 4187 883 4313
rect 936 4247 943 4413
rect 916 4216 923 4233
rect 956 4216 963 4433
rect 1056 4227 1063 4493
rect 1236 4467 1243 4943
rect 1316 4487 1323 5073
rect 1336 4667 1343 5573
rect 1356 5547 1363 5603
rect 1416 5436 1423 5533
rect 1456 5467 1463 5473
rect 1476 5407 1483 5423
rect 1436 5156 1463 5163
rect 1356 5107 1363 5153
rect 1456 5147 1463 5156
rect 1416 4967 1423 4973
rect 1496 4956 1503 5113
rect 1416 4483 1423 4953
rect 1516 4947 1523 4973
rect 1436 4927 1443 4943
rect 1536 4923 1543 5153
rect 1516 4916 1543 4923
rect 1436 4507 1443 4653
rect 1416 4476 1443 4483
rect 1156 4407 1163 4443
rect 1036 4187 1043 4203
rect 856 3967 863 4053
rect 996 3996 1003 4033
rect 836 3916 863 3923
rect 736 3696 763 3703
rect 656 3516 683 3523
rect 716 3516 723 3653
rect 756 3523 763 3696
rect 756 3516 773 3523
rect 656 3247 663 3516
rect 696 3383 703 3503
rect 776 3483 783 3513
rect 796 3507 803 3733
rect 756 3476 783 3483
rect 696 3376 723 3383
rect 616 2767 623 3053
rect 676 3036 683 3253
rect 696 3016 703 3213
rect 716 3207 723 3376
rect 696 2776 703 2973
rect 36 2303 43 2513
rect 276 2367 283 2533
rect 36 2296 63 2303
rect 56 2043 63 2296
rect 76 2227 83 2283
rect 76 2056 83 2073
rect 36 2036 63 2043
rect 36 1816 43 2036
rect 96 1707 103 2233
rect 176 2096 203 2103
rect 136 827 143 1553
rect 156 1267 163 1713
rect 176 1347 183 2096
rect 196 1727 203 1763
rect 216 1576 223 1693
rect 196 1316 203 1333
rect 176 1287 183 1303
rect 216 1116 223 1253
rect 256 1116 263 1353
rect 356 1287 363 2353
rect 376 2267 383 2283
rect 376 2063 383 2253
rect 396 2083 403 2573
rect 596 2536 603 2593
rect 396 2076 423 2083
rect 416 2067 423 2076
rect 376 2056 403 2063
rect 396 1803 403 2056
rect 496 1927 503 2073
rect 496 1807 503 1913
rect 376 1796 403 1803
rect 436 1796 463 1803
rect 436 1616 443 1796
rect 416 1367 423 1573
rect 407 1336 423 1343
rect 456 1336 483 1343
rect 396 1107 403 1333
rect 476 1307 483 1336
rect 476 1116 483 1153
rect 176 1096 203 1103
rect 176 823 183 1096
rect 176 816 203 823
rect 176 616 183 733
rect 196 636 203 816
rect 256 627 263 823
rect 216 387 223 613
rect 176 356 203 363
rect 176 307 183 356
rect 276 343 283 893
rect 416 867 423 1093
rect 496 1087 503 1103
rect 416 823 423 853
rect 416 816 443 823
rect 436 747 443 816
rect 436 616 443 713
rect 496 667 503 1073
rect 536 827 543 1693
rect 556 1587 563 2433
rect 576 2407 583 2533
rect 596 2087 603 2293
rect 616 2267 623 2593
rect 616 2063 623 2253
rect 636 2243 643 2763
rect 656 2287 663 2553
rect 676 2507 683 2543
rect 676 2307 683 2473
rect 676 2276 683 2293
rect 696 2267 703 2573
rect 716 2487 723 3033
rect 736 2567 743 3253
rect 756 2987 763 3476
rect 776 3247 783 3313
rect 816 3236 823 3253
rect 856 3223 863 3916
rect 936 3907 943 3983
rect 896 3467 903 3703
rect 956 3667 963 3723
rect 976 3516 983 3893
rect 1016 3687 1023 3993
rect 1016 3516 1023 3653
rect 1056 3507 1063 4213
rect 1136 3747 1143 4233
rect 1176 4003 1183 4093
rect 1236 4007 1243 4073
rect 1316 4007 1323 4473
rect 1356 4447 1363 4463
rect 1336 4147 1343 4203
rect 1156 3996 1183 4003
rect 1156 3907 1163 3996
rect 1176 3767 1183 3773
rect 1116 3687 1123 3713
rect 1136 3703 1143 3733
rect 1176 3716 1183 3753
rect 1256 3707 1263 3993
rect 1136 3696 1163 3703
rect 1196 3587 1203 3703
rect 1336 3607 1343 4133
rect 1356 3967 1363 4433
rect 1396 4167 1403 4473
rect 1416 4196 1423 4213
rect 1436 4087 1443 4476
rect 1516 4107 1523 4916
rect 1556 4707 1563 5853
rect 1576 5407 1583 5973
rect 1596 5647 1603 6116
rect 1636 6027 1643 6393
rect 1796 6127 1803 6593
rect 1836 6587 1843 7096
rect 1916 7096 1923 7113
rect 1856 6887 1863 7083
rect 1816 6027 1823 6553
rect 1856 6367 1863 6853
rect 1876 6583 1883 7093
rect 2116 7076 2123 7173
rect 1896 6867 1903 7073
rect 2176 7007 2183 7063
rect 2196 6867 2203 7353
rect 2216 7047 2223 7813
rect 2276 7087 2283 7333
rect 2296 7327 2303 7673
rect 2456 7543 2463 7773
rect 2476 7547 2483 7793
rect 2436 7536 2463 7543
rect 2376 7327 2383 7493
rect 2316 7307 2323 7323
rect 2396 7103 2403 7453
rect 2376 7096 2403 7103
rect 2376 7076 2383 7096
rect 2296 6847 2303 6873
rect 2356 6867 2363 7063
rect 2396 7047 2403 7063
rect 2436 6907 2443 7536
rect 2516 7307 2523 8293
rect 2656 8287 2663 8316
rect 2536 8003 2543 8023
rect 2536 7996 2563 8003
rect 2556 7856 2563 7996
rect 2536 7836 2543 7853
rect 2576 7836 2583 7853
rect 2616 7467 2623 7523
rect 2556 7327 2563 7343
rect 2676 7327 2683 9233
rect 2756 8547 2763 9873
rect 2816 9867 2823 9923
rect 2856 9847 2863 9956
rect 2816 9756 2823 9833
rect 2796 9507 2803 9713
rect 2836 9607 2843 9743
rect 2876 9727 2883 9743
rect 2796 9447 2803 9493
rect 2776 8047 2783 8893
rect 2796 8107 2803 9433
rect 2916 9407 2923 10213
rect 2976 9667 2983 9953
rect 2996 9943 3003 10333
rect 3056 10236 3063 10396
rect 3096 10236 3103 10253
rect 3076 10167 3083 10213
rect 2996 9936 3023 9943
rect 2816 9047 2823 9253
rect 2856 9243 2863 9293
rect 2856 9236 2883 9243
rect 2876 9016 2883 9213
rect 2936 9207 2943 9463
rect 2976 9447 2983 9463
rect 2816 8987 2823 9003
rect 2816 8807 2823 8973
rect 2916 8847 2923 9093
rect 2916 8816 2923 8833
rect 2956 8783 2963 9373
rect 2996 9227 3003 9913
rect 3036 9776 3063 9783
rect 3016 9387 3023 9753
rect 3036 9747 3043 9776
rect 2996 8787 3003 9013
rect 2856 8467 2863 8503
rect 2816 8296 2823 8453
rect 2896 8367 2903 8783
rect 2936 8776 2963 8783
rect 2936 8363 2943 8776
rect 2916 8356 2943 8363
rect 2876 8316 2903 8323
rect 2796 8036 2803 8093
rect 2716 7867 2723 8033
rect 2816 8027 2823 8193
rect 2856 8087 2863 8293
rect 2896 8287 2903 8316
rect 2896 8007 2903 8273
rect 2776 7987 2783 8003
rect 2756 7347 2763 7553
rect 2776 7507 2783 7873
rect 2796 7836 2803 7993
rect 2916 7767 2923 8356
rect 2776 7336 2783 7493
rect 2856 7467 2863 7563
rect 2796 7356 2803 7373
rect 2836 7356 2843 7373
rect 2916 7367 2923 7543
rect 2696 7076 2723 7083
rect 2616 7043 2623 7073
rect 2716 7047 2723 7076
rect 2616 7036 2643 7043
rect 2636 6876 2643 7036
rect 2676 7027 2683 7043
rect 2676 6876 2683 7013
rect 2716 6867 2723 7033
rect 2736 7027 2743 7073
rect 1916 6647 1923 6843
rect 1956 6747 1963 6843
rect 1876 6576 1903 6583
rect 1636 5807 1643 5903
rect 1656 5647 1663 5653
rect 1616 5636 1633 5643
rect 1616 5447 1623 5453
rect 1616 4967 1623 5433
rect 1636 5427 1643 5453
rect 1656 5403 1663 5633
rect 1676 5447 1683 6013
rect 1716 5447 1723 5633
rect 1756 5567 1763 6013
rect 1896 6007 1903 6576
rect 2076 6507 2083 6563
rect 1956 6416 1963 6433
rect 1916 6387 1923 6413
rect 1936 6347 1943 6383
rect 1836 5916 1843 5973
rect 1876 5916 1883 5933
rect 1856 5867 1863 5903
rect 1896 5896 1903 5913
rect 1916 5807 1923 6123
rect 1816 5636 1823 5793
rect 1936 5783 1943 5993
rect 1916 5776 1943 5783
rect 1796 5567 1803 5623
rect 1656 5396 1683 5403
rect 1676 5167 1683 5396
rect 1756 5143 1763 5553
rect 1876 5447 1883 5623
rect 1876 5416 1903 5423
rect 1736 5136 1763 5143
rect 1656 4963 1663 5133
rect 1656 4956 1683 4963
rect 1576 4503 1583 4713
rect 1556 4496 1583 4503
rect 1556 4483 1563 4496
rect 1536 4476 1563 4483
rect 1416 3927 1423 3973
rect 1456 3956 1463 4053
rect 1476 3976 1483 3993
rect 1436 3763 1443 3933
rect 1536 3767 1543 4476
rect 1616 4456 1623 4473
rect 1636 4216 1643 4393
rect 1616 3967 1623 4203
rect 1696 4067 1703 4933
rect 1736 4867 1743 5136
rect 1776 4967 1783 5013
rect 1656 3927 1663 3993
rect 1716 3976 1723 3993
rect 1756 3963 1763 4853
rect 1796 4687 1803 5153
rect 1836 4947 1843 5393
rect 1856 5087 1863 5413
rect 1876 5367 1883 5416
rect 1916 5407 1923 5776
rect 1976 5427 1983 6353
rect 2016 6116 2023 6453
rect 2056 6387 2063 6493
rect 1996 5967 2003 6093
rect 2056 5967 2063 6113
rect 2076 6087 2083 6393
rect 2096 6187 2103 6733
rect 2196 6267 2203 6603
rect 2216 6376 2223 6633
rect 2296 6596 2303 6833
rect 2416 6767 2423 6843
rect 2276 6396 2303 6403
rect 2256 6227 2263 6373
rect 2096 6107 2103 6123
rect 1996 5643 2003 5953
rect 2296 5947 2303 6396
rect 2316 6387 2323 6673
rect 2376 6107 2383 6593
rect 2556 6507 2563 6563
rect 2496 6396 2503 6493
rect 2536 6396 2543 6473
rect 2476 6376 2483 6393
rect 2576 6387 2583 6853
rect 2656 6407 2663 6753
rect 2756 6396 2763 6493
rect 2456 6127 2463 6253
rect 2156 5916 2163 5933
rect 2316 5916 2323 5933
rect 2076 5896 2103 5903
rect 2076 5807 2083 5896
rect 2376 5896 2383 5953
rect 2356 5656 2363 5693
rect 1996 5636 2023 5643
rect 2016 5407 2023 5593
rect 2036 5407 2043 5633
rect 2196 5567 2203 5603
rect 2136 5283 2143 5393
rect 2176 5387 2183 5403
rect 2116 5276 2143 5283
rect 1956 5143 1963 5163
rect 1936 5136 1963 5143
rect 1936 5087 1943 5136
rect 1956 4976 1963 5013
rect 1976 4947 1983 5183
rect 2116 5167 2123 5276
rect 2136 5163 2143 5173
rect 2136 5156 2163 5163
rect 2176 5143 2183 5183
rect 2216 5176 2223 5213
rect 2196 5147 2203 5163
rect 2156 5136 2183 5143
rect 1936 4727 1943 4943
rect 1896 4667 1903 4683
rect 1936 4676 1943 4693
rect 1976 4667 1983 4913
rect 1916 4647 1923 4663
rect 1796 4476 1803 4493
rect 1816 4387 1823 4463
rect 1856 4456 1883 4463
rect 1876 4227 1883 4456
rect 1856 4196 1883 4203
rect 1836 4127 1843 4163
rect 1876 4107 1883 4196
rect 1736 3956 1763 3963
rect 1436 3756 1463 3763
rect 1456 3743 1463 3756
rect 1456 3736 1483 3743
rect 1236 3536 1243 3573
rect 956 3227 963 3493
rect 836 3216 863 3223
rect 796 2967 803 3193
rect 876 3036 903 3043
rect 956 3036 963 3153
rect 756 2527 763 2933
rect 876 2787 883 3036
rect 956 2747 963 2993
rect 936 2736 953 2743
rect 636 2236 663 2243
rect 636 2067 643 2236
rect 716 2227 723 2393
rect 736 2167 743 2513
rect 796 2447 803 2733
rect 976 2727 983 3433
rect 996 3187 1003 3503
rect 1116 3496 1143 3503
rect 1416 3496 1423 3593
rect 1056 3483 1063 3493
rect 1056 3476 1083 3483
rect 1136 3367 1143 3496
rect 1116 3236 1123 3253
rect 1356 3207 1363 3233
rect 1016 3016 1043 3023
rect 996 2947 1003 3003
rect 1016 2887 1023 3016
rect 1136 2807 1143 3193
rect 1336 3167 1343 3203
rect 1356 3023 1363 3193
rect 1336 3016 1363 3023
rect 1076 2607 1083 2773
rect 1136 2756 1143 2793
rect 1356 2787 1363 3016
rect 1376 2787 1383 3053
rect 876 2576 903 2583
rect 596 2056 623 2063
rect 616 1627 623 2033
rect 676 1707 683 1783
rect 776 1687 783 2053
rect 616 1596 643 1603
rect 676 1596 683 1673
rect 716 1596 723 1613
rect 796 1607 803 2273
rect 876 2227 883 2576
rect 1076 2536 1083 2593
rect 896 2087 903 2263
rect 876 2056 903 2063
rect 876 1927 883 2056
rect 916 2043 923 2153
rect 936 2107 943 2263
rect 1116 2247 1123 2283
rect 1176 2207 1183 2263
rect 1196 2247 1203 2613
rect 916 2036 943 2043
rect 936 1847 943 2036
rect 616 1327 623 1596
rect 496 636 523 643
rect 516 427 523 636
rect 256 336 283 343
rect 176 143 183 293
rect 396 156 403 313
rect 456 307 463 363
rect 496 356 503 413
rect 536 367 543 633
rect 556 627 563 653
rect 516 327 523 343
rect 176 136 203 143
rect 616 123 623 1133
rect 636 347 643 1313
rect 656 1287 663 1583
rect 676 1087 683 1253
rect 696 1116 703 1153
rect 716 1136 723 1273
rect 736 1267 743 1293
rect 656 767 663 843
rect 696 836 703 893
rect 736 823 743 853
rect 716 816 743 823
rect 756 787 763 1093
rect 776 827 783 1113
rect 656 627 663 753
rect 696 636 703 773
rect 736 247 743 323
rect 656 136 663 153
rect 816 127 823 1613
rect 856 1587 863 1773
rect 916 1747 923 1783
rect 976 1783 983 2073
rect 967 1776 983 1783
rect 936 1623 943 1753
rect 936 1616 963 1623
rect 956 1596 963 1616
rect 936 1316 943 1583
rect 1016 1367 1023 1733
rect 1076 1647 1083 2093
rect 1136 2076 1163 2083
rect 1196 2076 1203 2213
rect 1096 1327 1103 1793
rect 956 1267 963 1283
rect 916 1083 923 1133
rect 916 1076 943 1083
rect 996 887 1003 1253
rect 1116 1247 1123 2053
rect 1136 2047 1143 2076
rect 1136 1747 1143 1763
rect 1196 1616 1203 2033
rect 1276 1807 1283 2733
rect 1296 1887 1303 2573
rect 1336 2543 1343 2713
rect 1336 2536 1363 2543
rect 1396 2307 1403 2573
rect 1436 2547 1443 3573
rect 1476 3503 1483 3736
rect 1636 3736 1663 3743
rect 1476 3496 1503 3503
rect 1476 3227 1483 3353
rect 1456 2767 1463 3033
rect 1516 2727 1523 2953
rect 1416 2063 1423 2193
rect 1416 2056 1443 2063
rect 1296 1767 1303 1873
rect 1156 1596 1183 1603
rect 1216 1596 1243 1603
rect 1156 1347 1163 1596
rect 1196 1316 1203 1353
rect 1236 1307 1243 1596
rect 1336 1347 1343 1783
rect 1376 1743 1383 1783
rect 1396 1747 1403 1753
rect 1356 1736 1383 1743
rect 1136 1287 1143 1293
rect 1216 1283 1223 1303
rect 1316 1287 1323 1313
rect 1216 1276 1243 1283
rect 1016 1087 1023 1213
rect 1156 1136 1163 1233
rect 1176 1116 1183 1153
rect 1236 1127 1243 1276
rect 936 836 943 873
rect 956 807 963 823
rect 856 136 863 773
rect 996 636 1003 693
rect 916 616 943 623
rect 916 587 923 616
rect 916 367 923 573
rect 976 567 983 623
rect 876 156 883 233
rect 916 156 923 193
rect 956 167 963 323
rect 1016 167 1023 793
rect 1116 323 1123 893
rect 1156 747 1163 843
rect 1176 636 1183 793
rect 1216 787 1223 823
rect 1236 807 1243 1113
rect 1196 567 1203 623
rect 1256 387 1263 1093
rect 1356 907 1363 1736
rect 1376 1323 1383 1573
rect 1396 1563 1403 1733
rect 1476 1563 1483 2273
rect 1536 2087 1543 3713
rect 1636 3667 1643 3736
rect 1676 3687 1683 3723
rect 1716 3716 1743 3723
rect 1616 3027 1623 3633
rect 1676 3516 1703 3523
rect 1676 3327 1683 3516
rect 1716 3467 1723 3483
rect 1736 3467 1743 3716
rect 1756 3516 1763 3733
rect 1836 3496 1843 3813
rect 1916 3727 1923 4533
rect 2016 4467 2023 4693
rect 2036 4407 2043 4913
rect 2056 4683 2063 5093
rect 2156 4936 2163 5136
rect 2176 4767 2183 4923
rect 2056 4676 2083 4683
rect 2076 4507 2083 4676
rect 2056 4476 2063 4493
rect 2096 4476 2103 4673
rect 2116 4467 2123 4733
rect 2076 4387 2083 4463
rect 2096 4196 2103 4233
rect 1976 3996 1983 4073
rect 2116 3716 2123 4373
rect 2156 4327 2163 4553
rect 2256 4456 2263 4493
rect 2276 4423 2283 5393
rect 2316 5327 2323 5643
rect 2416 5436 2423 5553
rect 2456 5447 2463 6073
rect 2376 5387 2383 5433
rect 2336 5127 2343 5143
rect 2376 5107 2383 5143
rect 2376 4956 2403 4963
rect 2376 4907 2383 4956
rect 2476 4927 2483 6173
rect 2516 6167 2523 6373
rect 2556 6347 2563 6353
rect 2556 5923 2563 6333
rect 2636 6087 2643 6393
rect 2736 6367 2743 6383
rect 2656 6027 2663 6083
rect 2556 5916 2583 5923
rect 2616 5916 2623 6013
rect 2596 5867 2603 5903
rect 2636 5896 2643 5913
rect 2496 5427 2503 5713
rect 2616 5656 2623 5753
rect 2556 5607 2563 5643
rect 2596 5627 2603 5643
rect 2696 5456 2703 5593
rect 2376 4807 2383 4893
rect 2396 4696 2423 4703
rect 2376 4567 2383 4683
rect 2396 4627 2403 4696
rect 2256 4416 2283 4423
rect 2256 4187 2263 4416
rect 2356 4203 2363 4273
rect 2336 4196 2363 4203
rect 2316 4167 2323 4183
rect 2156 3716 2163 3753
rect 1896 3587 1903 3673
rect 1956 3536 1963 3553
rect 2136 3496 2143 3593
rect 2196 3503 2203 3793
rect 2216 3747 2223 3983
rect 2196 3496 2223 3503
rect 1776 3483 1783 3493
rect 1776 3476 1803 3483
rect 1656 3236 1663 3293
rect 1676 3047 1683 3273
rect 1696 3256 1723 3263
rect 1696 3247 1703 3256
rect 1656 3007 1663 3023
rect 1556 2556 1563 2593
rect 1576 2587 1583 2893
rect 1596 2763 1603 2873
rect 1656 2787 1663 2993
rect 1696 2947 1703 3233
rect 1756 3227 1763 3243
rect 2056 3207 2063 3243
rect 2136 3236 2143 3253
rect 1876 3187 1883 3203
rect 1716 2776 1723 2933
rect 1596 2756 1623 2763
rect 1656 2756 1663 2773
rect 1596 2556 1603 2633
rect 1616 2507 1623 2756
rect 1736 2747 1743 3033
rect 1876 3016 1883 3053
rect 1856 2907 1863 3003
rect 2036 2763 2043 3193
rect 2116 3036 2123 3173
rect 2196 3047 2203 3473
rect 2156 3036 2183 3043
rect 2176 3027 2183 3036
rect 1636 2627 1643 2743
rect 1636 2276 1643 2593
rect 1596 1627 1603 1783
rect 1616 1667 1623 2263
rect 1696 2103 1703 2113
rect 1676 2096 1703 2103
rect 1696 1967 1703 2096
rect 1656 1616 1663 1953
rect 1396 1556 1423 1563
rect 1456 1556 1483 1563
rect 1616 1596 1643 1603
rect 1676 1596 1703 1603
rect 1616 1563 1623 1596
rect 1696 1567 1703 1596
rect 1616 1556 1643 1563
rect 1376 1316 1403 1323
rect 1416 1116 1423 1153
rect 1436 1087 1443 1133
rect 1116 316 1143 323
rect 1296 187 1303 733
rect 1416 667 1423 823
rect 1456 647 1463 1153
rect 1476 807 1483 1556
rect 1496 1147 1503 1353
rect 1636 1336 1643 1556
rect 1716 1323 1723 2473
rect 1736 2287 1743 2633
rect 1756 2447 1763 2763
rect 2036 2756 2063 2763
rect 1776 2543 1783 2713
rect 1876 2687 1883 2723
rect 1816 2556 1823 2673
rect 2096 2667 2103 3023
rect 2136 2983 2143 3023
rect 2116 2976 2143 2983
rect 1856 2556 1863 2573
rect 1776 2536 1803 2543
rect 1736 1607 1743 2273
rect 1756 2067 1763 2413
rect 1776 2267 1783 2513
rect 1836 2427 1843 2543
rect 1876 2263 1883 2653
rect 2096 2576 2103 2613
rect 2116 2587 2123 2976
rect 2036 2547 2043 2573
rect 2116 2536 2143 2543
rect 2076 2276 2083 2513
rect 1856 2256 1883 2263
rect 1656 1316 1683 1323
rect 1596 1127 1603 1293
rect 1656 1116 1663 1133
rect 1576 1096 1603 1103
rect 1576 767 1583 1096
rect 1616 723 1623 823
rect 1656 747 1663 823
rect 1596 716 1623 723
rect 1376 407 1383 633
rect 1436 607 1443 623
rect 1456 363 1463 393
rect 1596 367 1603 716
rect 1636 656 1643 733
rect 1676 587 1683 1316
rect 1696 1316 1723 1323
rect 1696 1007 1703 1316
rect 1736 1247 1743 1593
rect 1736 1167 1743 1233
rect 1696 707 1703 993
rect 1756 867 1763 2033
rect 1776 1827 1783 2253
rect 1816 2087 1823 2243
rect 1896 2076 1903 2273
rect 2136 2147 2143 2536
rect 2156 2527 2163 2613
rect 2196 2567 2203 3033
rect 2156 2507 2163 2513
rect 2136 2096 2143 2133
rect 1936 2076 1963 2083
rect 1756 827 1763 853
rect 1776 627 1783 1813
rect 1816 1787 1823 2073
rect 1956 2067 1963 2076
rect 2156 2076 2163 2113
rect 1916 2047 1923 2063
rect 1796 1767 1803 1783
rect 1896 1576 1903 1593
rect 1936 1587 1943 1793
rect 1956 1627 1963 2053
rect 2176 1787 2183 2293
rect 2056 1707 2063 1783
rect 2056 1687 2063 1693
rect 1976 1567 1983 1653
rect 2116 1616 2123 1753
rect 2196 1627 2203 2533
rect 2096 1607 2103 1613
rect 2136 1596 2143 1613
rect 1436 356 1463 363
rect 616 116 643 123
rect 1296 123 1303 173
rect 1336 136 1343 353
rect 1376 123 1383 173
rect 1556 156 1563 293
rect 1596 156 1603 353
rect 1636 347 1643 363
rect 1676 347 1683 363
rect 1796 327 1803 1133
rect 1836 1067 1843 1083
rect 1836 687 1843 1053
rect 1876 887 1883 1073
rect 1896 1067 1903 1133
rect 1936 967 1943 1333
rect 1896 816 1923 823
rect 1896 656 1903 673
rect 1856 647 1863 653
rect 1856 623 1863 633
rect 1856 616 1883 623
rect 1796 156 1803 313
rect 1916 307 1923 816
rect 1936 567 1943 953
rect 2016 867 2023 1313
rect 1956 607 1963 633
rect 1936 387 1943 553
rect 1976 367 1983 813
rect 1996 807 2003 833
rect 1836 143 1843 173
rect 1816 136 1843 143
rect 1976 127 1983 353
rect 2016 187 2023 793
rect 2036 787 2043 1313
rect 2076 1127 2083 1553
rect 2156 1387 2163 1613
rect 2096 1336 2103 1373
rect 2136 1336 2163 1343
rect 2116 1267 2123 1323
rect 2156 1267 2163 1336
rect 2096 1136 2103 1213
rect 2056 1047 2063 1113
rect 2056 836 2063 853
rect 2116 767 2123 823
rect 2116 656 2123 673
rect 2096 636 2103 653
rect 2136 636 2143 953
rect 2156 847 2163 893
rect 2216 747 2223 3093
rect 2156 627 2163 653
rect 2056 343 2063 373
rect 2056 336 2083 343
rect 2056 327 2063 336
rect 2156 327 2163 613
rect 2036 156 2043 293
rect 2216 207 2223 733
rect 2236 387 2243 4013
rect 2256 3996 2263 4073
rect 2256 3007 2263 3313
rect 2256 1287 2263 2993
rect 2276 2647 2283 2993
rect 2296 2987 2303 4153
rect 2316 3996 2343 4003
rect 2336 3447 2343 3996
rect 2356 3487 2363 4133
rect 2376 3987 2383 4313
rect 2456 4287 2463 4873
rect 2496 4667 2503 5413
rect 2536 4456 2563 4463
rect 2536 4327 2543 4456
rect 2376 3523 2383 3773
rect 2396 3736 2403 3773
rect 2436 3736 2443 3793
rect 2416 3547 2423 3723
rect 2376 3516 2403 3523
rect 2436 3516 2443 3553
rect 2456 3547 2463 4253
rect 2536 4207 2543 4273
rect 2576 4267 2583 5433
rect 2716 5407 2723 5423
rect 2736 5407 2743 6013
rect 2796 5907 2803 6153
rect 2816 6027 2823 7313
rect 2936 6867 2943 7833
rect 2836 6847 2843 6863
rect 2836 6827 2843 6833
rect 2836 6607 2843 6713
rect 2836 6107 2843 6113
rect 2856 5916 2863 5933
rect 2876 5707 2883 6613
rect 2896 6596 2923 6603
rect 2896 6367 2903 6596
rect 2896 6116 2923 6123
rect 2896 5967 2903 6116
rect 2956 6003 2963 8593
rect 2996 8507 3003 8773
rect 3016 8587 3023 9273
rect 3036 8527 3043 9653
rect 3056 9527 3063 9733
rect 3076 9547 3083 9743
rect 3056 9267 3063 9513
rect 3076 9447 3083 9533
rect 3096 9023 3103 9633
rect 3136 9327 3143 10393
rect 3156 10387 3163 10433
rect 3196 9807 3203 10573
rect 3256 10007 3263 10936
rect 3376 10883 3383 11213
rect 3456 11196 3463 11213
rect 3436 11167 3443 11183
rect 3476 11127 3483 11183
rect 3556 10923 3563 11133
rect 3676 10923 3683 11216
rect 4176 11207 4183 11293
rect 4116 11196 4143 11203
rect 3716 11167 3723 11183
rect 3556 10916 3583 10923
rect 3656 10916 3683 10923
rect 3376 10876 3403 10883
rect 3476 10716 3503 10723
rect 3456 10647 3463 10703
rect 3496 10667 3503 10716
rect 3536 10703 3543 10773
rect 3516 10696 3543 10703
rect 3336 10427 3343 10443
rect 3376 10427 3383 10553
rect 3576 10527 3583 10916
rect 3276 10236 3283 10253
rect 3376 10227 3383 10253
rect 3256 9667 3263 9993
rect 3396 9927 3403 10253
rect 3296 9916 3323 9923
rect 3276 9723 3283 9773
rect 3316 9736 3323 9916
rect 3276 9716 3303 9723
rect 3156 9496 3203 9503
rect 3156 9447 3163 9496
rect 3196 9476 3203 9496
rect 3236 9476 3243 9493
rect 3156 9407 3163 9433
rect 3216 9347 3223 9443
rect 3196 9276 3203 9333
rect 3176 9107 3183 9263
rect 3296 9027 3303 9653
rect 3336 9467 3343 9723
rect 3416 9507 3423 9953
rect 3436 9507 3443 10513
rect 3516 10236 3523 10253
rect 3556 10236 3563 10353
rect 3576 10267 3583 10443
rect 3596 10236 3603 10273
rect 3636 10227 3643 10423
rect 3656 10287 3663 10433
rect 3456 9947 3463 9973
rect 3536 9956 3543 10013
rect 3476 9927 3483 9943
rect 3396 9427 3403 9463
rect 3396 9387 3403 9413
rect 3336 9256 3363 9263
rect 3336 9227 3343 9256
rect 3376 9236 3383 9273
rect 3396 9256 3403 9293
rect 3096 9016 3123 9023
rect 3076 8787 3083 9003
rect 3116 8687 3123 9016
rect 3156 8796 3163 8833
rect 3176 8687 3183 8783
rect 3127 8656 3133 8663
rect 3156 8536 3163 8653
rect 3056 8487 3063 8523
rect 3216 8523 3223 9013
rect 3276 8623 3283 8773
rect 3296 8747 3303 8953
rect 3316 8847 3323 8963
rect 3276 8616 3303 8623
rect 3196 8516 3223 8523
rect 3096 8336 3103 8473
rect 3056 8316 3083 8323
rect 3036 8127 3043 8313
rect 3056 8287 3063 8316
rect 3136 8187 3143 8513
rect 3196 8467 3203 8516
rect 3296 8343 3303 8616
rect 3316 8527 3323 8813
rect 3456 8767 3463 9033
rect 3476 9003 3483 9493
rect 3496 9047 3503 9373
rect 3476 8996 3503 9003
rect 3276 8336 3303 8343
rect 3256 8307 3263 8333
rect 3276 8316 3283 8336
rect 2976 8027 2983 8043
rect 3016 8036 3023 8073
rect 3036 8007 3043 8023
rect 3056 7827 3063 8153
rect 2976 7327 2983 7373
rect 2976 6127 2983 6383
rect 2976 6107 2983 6113
rect 2956 5996 2983 6003
rect 2896 5916 2923 5923
rect 2776 5567 2783 5633
rect 2796 5527 2803 5623
rect 2656 4947 2663 5133
rect 2676 4956 2683 5163
rect 2696 5127 2703 5143
rect 2696 4887 2703 4943
rect 2736 4747 2743 5143
rect 2656 4676 2663 4693
rect 2616 4443 2623 4613
rect 2636 4507 2643 4663
rect 2596 4436 2623 4443
rect 2596 4196 2603 4373
rect 2616 4307 2623 4436
rect 2576 4027 2583 4183
rect 2616 4027 2623 4183
rect 2376 3287 2383 3516
rect 2416 3483 2423 3503
rect 2456 3496 2463 3513
rect 2396 3476 2423 3483
rect 2316 3056 2323 3253
rect 2316 2743 2323 2773
rect 2316 2736 2343 2743
rect 2316 2536 2323 2693
rect 2356 2487 2363 3223
rect 2376 2687 2383 2743
rect 2276 2296 2303 2303
rect 2276 2247 2283 2296
rect 2396 2267 2403 3476
rect 2416 3207 2423 3223
rect 2436 3027 2443 3413
rect 2456 3227 2463 3353
rect 2296 2047 2303 2073
rect 2296 1796 2303 2033
rect 2276 1087 2283 1753
rect 2336 1667 2343 2253
rect 2376 2096 2383 2233
rect 2387 1916 2393 1923
rect 2336 1596 2343 1653
rect 2376 1596 2403 1603
rect 2396 1567 2403 1596
rect 2416 1347 2423 2593
rect 2436 1787 2443 2533
rect 2316 1167 2323 1293
rect 2356 1267 2363 1283
rect 2336 1116 2343 1153
rect 2356 947 2363 1253
rect 2376 1127 2383 1293
rect 2416 1167 2423 1333
rect 2436 1267 2443 1593
rect 2356 767 2363 803
rect 2396 767 2403 1073
rect 2296 636 2343 643
rect 2296 427 2303 636
rect 2336 616 2343 636
rect 2376 603 2383 673
rect 2456 607 2463 2253
rect 2476 827 2483 3993
rect 2636 3967 2643 4473
rect 2656 4207 2663 4233
rect 2496 3947 2503 3963
rect 2496 2527 2503 3813
rect 2516 3707 2523 3893
rect 2536 3707 2543 3953
rect 2516 2607 2523 3553
rect 2536 3007 2543 3533
rect 2576 3223 2583 3913
rect 2596 3723 2603 3933
rect 2676 3743 2683 4553
rect 2716 4207 2723 4493
rect 2716 4027 2723 4193
rect 2756 4127 2763 5473
rect 2776 5427 2783 5493
rect 2776 4447 2783 5393
rect 2796 4967 2803 5513
rect 2836 4587 2843 5573
rect 2856 5427 2863 5633
rect 2916 5587 2923 5916
rect 2936 5647 2943 5923
rect 2976 5607 2983 5996
rect 2996 5507 3003 7813
rect 3016 7807 3023 7823
rect 3156 7627 3163 8233
rect 3216 8036 3223 8073
rect 3196 8007 3203 8023
rect 3196 7843 3203 7973
rect 3236 7947 3243 8023
rect 3196 7836 3223 7843
rect 3256 7836 3283 7843
rect 3156 7543 3163 7613
rect 3096 7507 3103 7543
rect 3136 7536 3163 7543
rect 3056 7147 3063 7323
rect 3036 6607 3043 7133
rect 3096 6856 3103 7453
rect 3116 7096 3123 7333
rect 3196 7147 3203 7836
rect 3276 7787 3283 7836
rect 3296 7587 3303 7853
rect 3247 7556 3263 7563
rect 3256 7387 3263 7556
rect 3336 7527 3343 7563
rect 3376 7547 3383 7563
rect 3256 7356 3263 7373
rect 3136 7047 3143 7083
rect 3056 6527 3063 6853
rect 3116 6707 3123 6843
rect 3196 6827 3203 7093
rect 3176 6607 3183 6813
rect 3216 6583 3223 6953
rect 3156 6567 3163 6583
rect 3196 6576 3223 6583
rect 3116 6267 3123 6383
rect 3036 5916 3063 5923
rect 2896 5407 2903 5433
rect 2916 5416 2923 5453
rect 2936 5436 2943 5493
rect 2896 5187 2903 5393
rect 2936 5123 2943 5153
rect 3016 5147 3023 5633
rect 3036 5627 3043 5916
rect 3116 5667 3123 6253
rect 3136 6136 3143 6173
rect 3156 5687 3163 6123
rect 3196 5987 3203 6576
rect 3056 5636 3083 5643
rect 3056 5627 3063 5636
rect 3087 5616 3103 5623
rect 3136 5607 3143 5623
rect 3156 5616 3183 5623
rect 3036 5427 3043 5553
rect 2916 5116 2943 5123
rect 2916 4976 2923 5116
rect 2896 4967 2903 4973
rect 2936 4956 2963 4963
rect 2876 4696 2883 4933
rect 2956 4887 2963 4956
rect 2976 4947 2983 5133
rect 3036 5107 3043 5143
rect 2916 4696 2943 4703
rect 2816 4456 2823 4513
rect 2936 4507 2943 4696
rect 2876 4476 2883 4493
rect 2916 4207 2923 4253
rect 2936 4227 2943 4473
rect 2996 4467 3003 4953
rect 2716 3996 2723 4013
rect 2736 3967 2743 3983
rect 2776 3976 2783 3993
rect 2816 3767 2823 3973
rect 2656 3736 2683 3743
rect 2656 3727 2663 3736
rect 2596 3716 2623 3723
rect 2596 3487 2603 3716
rect 2696 3707 2703 3753
rect 2596 3267 2603 3473
rect 2636 3327 2643 3703
rect 2676 3256 2703 3263
rect 2576 3216 2603 3223
rect 2556 3036 2563 3053
rect 2596 3036 2603 3216
rect 2616 3107 2623 3243
rect 2656 3207 2663 3253
rect 2676 3247 2683 3256
rect 2636 3036 2643 3113
rect 2536 2307 2543 2973
rect 2576 2967 2583 3023
rect 2616 2987 2623 3023
rect 2556 2667 2563 2873
rect 2596 2727 2603 2743
rect 2596 2556 2603 2593
rect 2636 2556 2643 2693
rect 2716 2683 2723 3513
rect 2736 3487 2743 3713
rect 2736 3227 2743 3243
rect 2696 2676 2723 2683
rect 2656 2587 2663 2633
rect 2656 2547 2663 2573
rect 2676 2347 2683 2523
rect 2656 2296 2663 2333
rect 2696 2323 2703 2676
rect 2716 2536 2723 2653
rect 2756 2627 2763 3573
rect 2816 3527 2823 3753
rect 2836 3267 2843 4053
rect 2916 3716 2923 4033
rect 2936 3967 2943 4193
rect 2996 4016 3003 4093
rect 3016 4067 3023 4993
rect 3056 4707 3063 5553
rect 3116 4967 3123 5493
rect 3156 5487 3163 5616
rect 3236 5587 3243 5913
rect 3256 5663 3263 7253
rect 3296 6847 3303 7353
rect 3356 7027 3363 7063
rect 3296 6403 3303 6833
rect 3316 6807 3323 6843
rect 3296 6396 3323 6403
rect 3356 6396 3363 6813
rect 3396 6623 3403 6853
rect 3416 6827 3423 8293
rect 3456 8043 3463 8533
rect 3476 8523 3483 8996
rect 3476 8516 3503 8523
rect 3516 8267 3523 9913
rect 3536 9787 3543 9913
rect 3576 9467 3583 10213
rect 3596 9907 3603 9953
rect 3656 9947 3663 10253
rect 3636 9847 3643 9933
rect 3556 8996 3583 9003
rect 3556 8827 3563 8996
rect 3576 8516 3583 8533
rect 3596 8327 3603 9793
rect 3616 9247 3623 9713
rect 3636 9627 3643 9833
rect 3676 9707 3683 10916
rect 3716 10307 3723 11153
rect 3756 10716 3763 11193
rect 4116 11187 4123 11196
rect 3896 10867 3903 10883
rect 3836 10703 3843 10753
rect 3816 10696 3843 10703
rect 3716 10207 3723 10293
rect 3776 10267 3783 10693
rect 3807 10456 3823 10463
rect 3796 10187 3803 10453
rect 3836 10387 3843 10443
rect 3836 10256 3843 10273
rect 3876 10267 3883 10613
rect 3816 10247 3823 10253
rect 3696 9507 3703 9773
rect 3736 9747 3743 9773
rect 3756 9756 3763 9963
rect 3836 9943 3843 10193
rect 3816 9936 3843 9943
rect 3836 9807 3843 9853
rect 3836 9743 3843 9793
rect 3776 9727 3783 9743
rect 3816 9736 3843 9743
rect 3656 9296 3663 9483
rect 3696 9476 3703 9493
rect 3616 9007 3623 9113
rect 3636 8947 3643 9213
rect 3716 9067 3723 9463
rect 3636 8787 3643 8833
rect 3676 8767 3683 8813
rect 3616 8427 3623 8733
rect 3576 8296 3583 8313
rect 3616 8296 3623 8413
rect 3456 8036 3483 8043
rect 3516 8036 3523 8073
rect 3496 7967 3503 8023
rect 3536 7887 3543 8023
rect 3476 7836 3483 7873
rect 3436 6827 3443 7373
rect 3456 7356 3463 7413
rect 3476 7376 3483 7533
rect 3556 7427 3563 8253
rect 3496 7356 3503 7393
rect 3516 7123 3523 7353
rect 3496 7116 3523 7123
rect 3396 6616 3413 6623
rect 3396 6407 3403 6583
rect 3296 6027 3303 6396
rect 3436 6387 3443 6813
rect 3456 6567 3463 6583
rect 3476 6387 3483 7073
rect 3376 6376 3403 6383
rect 3396 6247 3403 6376
rect 3376 6116 3383 6213
rect 3476 6127 3483 6133
rect 3296 5916 3303 5993
rect 3336 5916 3343 6073
rect 3356 5947 3363 6103
rect 3256 5656 3283 5663
rect 3256 5587 3263 5623
rect 3156 5416 3163 5473
rect 3176 5436 3183 5533
rect 3216 5436 3223 5513
rect 3156 5136 3183 5143
rect 3156 4956 3163 5093
rect 3176 5047 3183 5136
rect 3176 4936 3183 4953
rect 3136 4767 3143 4933
rect 3196 4887 3203 5413
rect 3136 4676 3143 4733
rect 3176 4663 3183 4693
rect 3116 4567 3123 4663
rect 3156 4656 3183 4663
rect 3156 4507 3163 4656
rect 3076 4447 3083 4463
rect 3036 4187 3043 4203
rect 2956 3967 2963 4013
rect 2976 3967 2983 3983
rect 2956 3703 2963 3953
rect 3056 3823 3063 4433
rect 3076 4216 3083 4293
rect 3056 3816 3083 3823
rect 2896 3587 2903 3703
rect 2936 3696 2963 3703
rect 3076 3703 3083 3816
rect 3096 3747 3103 3993
rect 3176 3947 3183 4553
rect 3196 3987 3203 4433
rect 3236 4016 3243 4213
rect 3256 4047 3263 5493
rect 3276 4207 3283 5656
rect 3296 5147 3303 5573
rect 3316 5567 3323 5893
rect 3296 4243 3303 5113
rect 3316 4567 3323 5453
rect 3336 4727 3343 5153
rect 3356 5143 3363 5773
rect 3376 5467 3383 5953
rect 3396 5907 3403 6103
rect 3396 5436 3403 5513
rect 3436 5436 3443 5593
rect 3416 5387 3423 5413
rect 3476 5267 3483 5653
rect 3456 5156 3463 5173
rect 3356 5136 3383 5143
rect 3376 4943 3383 5033
rect 3456 4956 3463 4973
rect 3376 4936 3403 4943
rect 3376 4696 3383 4936
rect 3436 4887 3443 4943
rect 3356 4527 3363 4683
rect 3336 4463 3343 4493
rect 3316 4456 3343 4463
rect 3316 4267 3323 4456
rect 3296 4236 3323 4243
rect 3276 4147 3283 4163
rect 3216 3967 3223 3983
rect 3176 3723 3183 3733
rect 3156 3716 3183 3723
rect 3076 3696 3103 3703
rect 2896 3536 2903 3553
rect 2876 3516 2883 3533
rect 2916 3516 2923 3553
rect 2796 3056 2823 3063
rect 2796 2787 2803 3056
rect 2856 2743 2863 3053
rect 2996 2807 3003 3273
rect 3036 3227 3043 3243
rect 3036 3187 3043 3213
rect 2836 2736 2863 2743
rect 2836 2647 2843 2736
rect 2676 2316 2703 2323
rect 2596 2276 2603 2293
rect 2636 2263 2643 2293
rect 2576 2247 2583 2263
rect 2616 2256 2643 2263
rect 2676 2127 2683 2316
rect 2816 2283 2823 2613
rect 2836 2576 2843 2593
rect 3016 2563 3023 3173
rect 3056 3127 3063 3593
rect 3076 3287 3083 3696
rect 3136 3687 3143 3703
rect 3196 3587 3203 3713
rect 3196 3527 3203 3533
rect 3136 3496 3143 3513
rect 3056 3016 3063 3093
rect 3096 3027 3103 3493
rect 3116 3236 3143 3243
rect 3136 3187 3143 3236
rect 3056 2776 3063 2793
rect 3096 2776 3103 2993
rect 3076 2747 3083 2763
rect 2996 2556 3023 2563
rect 2996 2323 3003 2556
rect 2516 1827 2523 2113
rect 2556 2076 2563 2113
rect 2596 2076 2623 2083
rect 2616 2047 2623 2076
rect 2596 1816 2603 1833
rect 2496 1587 2503 1793
rect 2556 1767 2563 1783
rect 2556 1727 2563 1753
rect 2576 1647 2583 1653
rect 2576 1596 2583 1633
rect 2616 1607 2623 2033
rect 2696 1927 2703 2283
rect 2796 2276 2823 2283
rect 2976 2316 3003 2323
rect 2976 2283 2983 2316
rect 2976 2276 3003 2283
rect 2796 2107 2803 2276
rect 2656 1803 2663 1913
rect 2636 1796 2663 1803
rect 2736 1787 2743 2093
rect 2756 1807 2763 2073
rect 2776 2067 2783 2093
rect 2896 2076 2903 2093
rect 2876 2047 2883 2063
rect 2976 1807 2983 2276
rect 3016 1807 3023 2113
rect 2736 1756 2763 1763
rect 2736 1707 2743 1756
rect 2496 1307 2503 1573
rect 2356 596 2383 603
rect 2476 407 2483 813
rect 2496 647 2503 1293
rect 2556 1247 2563 1323
rect 2536 1116 2543 1233
rect 2576 1227 2583 1343
rect 2616 1336 2623 1493
rect 2596 1096 2603 1273
rect 2556 856 2563 913
rect 2616 907 2623 1133
rect 2616 863 2623 893
rect 2756 867 2763 1733
rect 2856 1596 2863 1693
rect 2836 1507 2843 1583
rect 2876 1576 2883 1613
rect 2816 1276 2843 1283
rect 2796 927 2803 1233
rect 2836 1107 2843 1276
rect 2896 1187 2903 1793
rect 2856 1007 2863 1083
rect 2596 856 2623 863
rect 2576 616 2583 713
rect 2556 587 2563 603
rect 2476 327 2483 393
rect 2576 376 2583 393
rect 1296 116 1323 123
rect 1356 116 1383 123
rect 2216 107 2223 193
rect 2276 136 2283 193
rect 2316 123 2323 313
rect 2556 167 2563 363
rect 2596 147 2603 593
rect 2756 383 2763 853
rect 2796 656 2803 913
rect 2816 856 2823 953
rect 2836 827 2843 843
rect 2876 607 2883 1073
rect 2936 847 2943 1693
rect 3036 1667 3043 2733
rect 3116 2543 3123 2573
rect 3096 2536 3123 2543
rect 3076 2276 3103 2283
rect 3096 2247 3103 2276
rect 3096 2076 3103 2213
rect 3136 2127 3143 3113
rect 3136 2076 3163 2083
rect 3076 2056 3083 2073
rect 3056 1596 3063 1793
rect 3116 1747 3123 2063
rect 3156 2047 3163 2076
rect 3096 1596 3103 1613
rect 3136 1596 3143 1873
rect 3176 1787 3183 3473
rect 3196 1767 3203 3013
rect 3216 2727 3223 3713
rect 3236 3527 3243 3973
rect 3256 3483 3263 3933
rect 3316 3927 3323 4236
rect 3336 4187 3343 4313
rect 3276 3496 3283 3833
rect 3236 3476 3263 3483
rect 3236 3027 3243 3373
rect 3296 3147 3303 3733
rect 3396 3563 3403 4713
rect 3436 3607 3443 4713
rect 3476 4463 3483 5253
rect 3456 4456 3483 4463
rect 3456 3607 3463 4456
rect 3496 4447 3503 7116
rect 3516 5927 3523 7093
rect 3556 7063 3563 7413
rect 3576 7107 3583 8033
rect 3596 7567 3603 7893
rect 3636 7647 3643 8673
rect 3616 7107 3623 7533
rect 3636 7063 3643 7073
rect 3556 7056 3583 7063
rect 3616 7056 3643 7063
rect 3536 6843 3543 6893
rect 3616 6843 3623 6913
rect 3636 6867 3643 7056
rect 3536 6836 3563 6843
rect 3596 6836 3623 6843
rect 3516 5507 3523 5913
rect 3536 5807 3543 6813
rect 3656 6767 3663 8273
rect 3596 6583 3603 6613
rect 3596 6576 3623 6583
rect 3656 6567 3663 6583
rect 3556 6107 3563 6123
rect 3576 5916 3583 6413
rect 3636 6396 3643 6563
rect 3676 6507 3683 8313
rect 3696 7907 3703 9033
rect 3736 8967 3743 9493
rect 3716 8047 3723 8773
rect 3736 8687 3743 8873
rect 3756 8507 3763 9293
rect 3736 8267 3743 8373
rect 3756 8023 3763 8333
rect 3736 8016 3763 8023
rect 3776 8323 3783 9613
rect 3796 9247 3803 9253
rect 3796 9016 3803 9233
rect 3816 9047 3823 9736
rect 3836 9267 3843 9313
rect 3856 9307 3863 9813
rect 3876 9647 3883 10253
rect 3896 9887 3903 10853
rect 3916 10347 3923 10913
rect 3936 10867 3943 11183
rect 4116 10963 4123 11173
rect 4116 10956 4143 10963
rect 4136 10923 4143 10956
rect 4116 10916 4143 10923
rect 4296 10923 4303 11173
rect 4336 11163 4343 11293
rect 4616 11196 4643 11203
rect 4616 11167 4623 11196
rect 4336 11156 4363 11163
rect 4296 10916 4323 10923
rect 3916 10167 3923 10333
rect 3876 9476 3903 9483
rect 3876 9307 3883 9476
rect 3916 9407 3923 9443
rect 3856 9276 3863 9293
rect 3936 9283 3943 10833
rect 4036 10807 4043 10913
rect 4396 10903 4403 11153
rect 4056 10827 4063 10903
rect 4096 10887 4103 10903
rect 4336 10867 4343 10903
rect 4376 10896 4403 10903
rect 4036 10747 4043 10753
rect 3996 10707 4003 10733
rect 4016 10676 4023 10713
rect 4036 10696 4043 10733
rect 4076 10683 4083 10793
rect 4056 10676 4083 10683
rect 4096 10587 4103 10793
rect 4116 10507 4123 10813
rect 4116 10436 4123 10493
rect 4096 10367 4103 10423
rect 4156 10267 4163 10423
rect 4076 10187 4083 10203
rect 4036 9976 4053 9983
rect 4016 9947 4023 9963
rect 3996 9776 4003 9933
rect 3956 9756 3983 9763
rect 3956 9447 3963 9756
rect 4016 9507 4023 9693
rect 4056 9667 4063 9973
rect 4076 9767 4083 10173
rect 3936 9276 3963 9283
rect 3876 9127 3883 9263
rect 3916 9256 3943 9263
rect 3836 9007 3843 9023
rect 3816 8907 3823 9003
rect 3856 8947 3863 9003
rect 3856 8776 3863 8893
rect 3836 8747 3843 8763
rect 3836 8587 3843 8733
rect 3796 8487 3803 8503
rect 3836 8467 3843 8573
rect 3776 8316 3803 8323
rect 3696 7816 3703 7853
rect 3716 7836 3723 7913
rect 3756 7836 3763 7873
rect 3696 7356 3703 7573
rect 3776 7447 3783 8316
rect 3836 7567 3843 8273
rect 3856 8107 3863 8303
rect 3736 7356 3743 7373
rect 3756 7227 3763 7373
rect 3736 6127 3743 7093
rect 3756 6587 3763 6873
rect 3776 6863 3783 7393
rect 3796 7267 3803 7553
rect 3816 7427 3823 7523
rect 3856 7467 3863 8093
rect 3876 8047 3883 8073
rect 3876 7827 3883 8033
rect 3896 7867 3903 8713
rect 3916 8327 3923 9033
rect 3936 8847 3943 9256
rect 3956 8307 3963 9276
rect 3976 8307 3983 8533
rect 4016 8503 4023 9493
rect 4076 9476 4083 9493
rect 4056 9407 4063 9473
rect 4156 9443 4163 9953
rect 4136 9436 4163 9443
rect 4096 9327 4103 9433
rect 4116 9147 4123 9293
rect 4136 9183 4143 9436
rect 4136 9176 4163 9183
rect 4036 9016 4043 9033
rect 4076 9016 4083 9093
rect 4076 8796 4083 8853
rect 4116 8796 4123 8833
rect 4096 8767 4103 8783
rect 4116 8503 4123 8593
rect 4016 8496 4043 8503
rect 3956 8107 3963 8293
rect 3916 7907 3923 8013
rect 3936 7887 3943 8023
rect 3936 7836 3943 7873
rect 3976 7867 3983 8023
rect 3996 7816 4003 8013
rect 3956 7803 3963 7813
rect 3936 7796 3963 7803
rect 3836 6947 3843 7043
rect 3856 6927 3863 7373
rect 3896 7343 3903 7373
rect 3896 7336 3923 7343
rect 3856 6876 3863 6893
rect 3776 6856 3803 6863
rect 3756 6407 3763 6573
rect 3776 6467 3783 6856
rect 3876 6627 3883 7013
rect 3816 6583 3823 6613
rect 3816 6576 3843 6583
rect 3876 6567 3883 6583
rect 3896 6383 3903 6593
rect 3916 6387 3923 6413
rect 3876 6376 3903 6383
rect 3896 6367 3903 6376
rect 3596 5727 3603 5903
rect 3656 5887 3663 5903
rect 3576 5547 3583 5643
rect 3596 5447 3603 5573
rect 3516 5427 3523 5443
rect 3636 5436 3643 5453
rect 3516 5147 3523 5413
rect 3556 4987 3563 5033
rect 3556 4663 3563 4973
rect 3596 4967 3603 5173
rect 3616 5167 3623 5273
rect 3676 5176 3683 5193
rect 3656 5023 3663 5163
rect 3696 5027 3703 5913
rect 3636 5016 3663 5023
rect 3636 4936 3643 5016
rect 3656 4956 3663 4993
rect 3596 4676 3603 4873
rect 3556 4656 3583 4663
rect 3636 4503 3643 4683
rect 3616 4496 3643 4503
rect 3696 4496 3703 4913
rect 3476 3947 3483 4293
rect 3516 4196 3523 4213
rect 3516 4016 3543 4023
rect 3536 3967 3543 4016
rect 3556 3703 3563 4233
rect 3616 4167 3623 4496
rect 3716 4463 3723 6013
rect 3736 5687 3743 5693
rect 3736 5407 3743 5673
rect 3756 5587 3763 6153
rect 3896 6143 3903 6293
rect 3896 6136 3923 6143
rect 3836 5943 3843 6113
rect 3816 5936 3843 5943
rect 3816 5923 3823 5936
rect 3796 5916 3823 5923
rect 3796 5667 3803 5916
rect 3836 5887 3843 5903
rect 3876 5896 3883 5913
rect 3796 5627 3803 5653
rect 3816 5607 3823 5643
rect 3896 5623 3903 5973
rect 3916 5883 3923 6136
rect 3936 6063 3943 7796
rect 3956 7387 3963 7753
rect 3956 7356 3963 7373
rect 3996 7063 4003 7553
rect 4016 7387 4023 8313
rect 4036 8047 4043 8496
rect 4056 8447 4063 8503
rect 4096 8496 4123 8503
rect 4056 8296 4063 8373
rect 4116 8363 4123 8496
rect 4116 8356 4143 8363
rect 4116 8316 4123 8333
rect 4096 8227 4103 8303
rect 4036 7727 4043 7853
rect 4056 7627 4063 7853
rect 4076 7583 4083 7853
rect 4096 7827 4103 8213
rect 4076 7576 4103 7583
rect 4056 7127 4063 7563
rect 3996 7056 4023 7063
rect 3996 6383 4003 7056
rect 4036 7027 4043 7043
rect 4056 6947 4063 7063
rect 4076 6927 4083 7373
rect 4096 7347 4103 7576
rect 4116 7167 4123 7833
rect 4136 7747 4143 8356
rect 4156 8027 4163 9176
rect 4136 7047 4143 7613
rect 4156 7587 4163 7873
rect 4176 7867 4183 10853
rect 4336 10847 4343 10853
rect 4396 10767 4403 10896
rect 4236 10716 4283 10723
rect 4196 10247 4203 10713
rect 4236 10707 4243 10716
rect 4476 10716 4503 10723
rect 4536 10716 4553 10723
rect 4236 10687 4243 10693
rect 4296 10627 4303 10703
rect 4336 10683 4343 10693
rect 4316 10676 4343 10683
rect 4216 10443 4223 10453
rect 4276 10443 4283 10513
rect 4216 10436 4243 10443
rect 4276 10436 4303 10443
rect 4216 9943 4223 10233
rect 4236 10163 4243 10436
rect 4296 10287 4303 10436
rect 4316 10407 4323 10676
rect 4476 10647 4483 10716
rect 4556 10667 4563 10713
rect 4576 10407 4583 10713
rect 4296 10236 4303 10253
rect 4256 10187 4263 10233
rect 4236 10156 4263 10163
rect 4256 9967 4263 10156
rect 4216 9936 4243 9943
rect 4216 9827 4223 9936
rect 4216 9736 4223 9753
rect 4196 9467 4203 9713
rect 4216 9367 4223 9593
rect 4296 9467 4303 9733
rect 4316 9727 4323 10223
rect 4356 9963 4363 10273
rect 4556 10203 4563 10233
rect 4496 10167 4503 10203
rect 4536 10196 4563 10203
rect 4616 10167 4623 10713
rect 4356 9956 4383 9963
rect 4496 9747 4503 9793
rect 4556 9756 4563 9813
rect 4536 9667 4543 9743
rect 4336 9476 4343 9513
rect 4236 9247 4243 9273
rect 4256 8976 4283 8983
rect 4256 8847 4263 8976
rect 4276 8816 4283 8853
rect 4296 8607 4303 8783
rect 4316 8767 4323 8973
rect 4336 8787 4343 9353
rect 4356 8747 4363 9433
rect 4416 9427 4423 9473
rect 4376 8887 4383 9273
rect 4396 9187 4403 9273
rect 4436 8987 4443 9653
rect 4476 9307 4483 9313
rect 4496 9276 4523 9283
rect 4516 9267 4523 9276
rect 4496 8947 4503 9233
rect 4516 8987 4523 9253
rect 4536 9087 4543 9633
rect 4576 9507 4583 9953
rect 4656 9747 4663 11233
rect 6116 11227 6123 11233
rect 5296 11216 5323 11223
rect 4676 10387 4683 11193
rect 5296 11187 5303 11216
rect 5816 11216 5843 11223
rect 4716 11176 4743 11183
rect 5016 11176 5043 11183
rect 4696 10947 4703 11163
rect 4716 11047 4723 11176
rect 5016 11087 5023 11176
rect 4756 10936 4783 10943
rect 4696 10467 4703 10933
rect 4736 10847 4743 10893
rect 4756 10827 4763 10936
rect 4956 10927 4963 11073
rect 4836 10916 4863 10923
rect 4736 10716 4743 10753
rect 4796 10747 4803 10903
rect 4836 10887 4843 10916
rect 5116 10867 5123 10883
rect 4816 10716 4823 10773
rect 4836 10707 4843 10733
rect 4896 10707 4903 10813
rect 5236 10743 5243 10923
rect 4996 10736 5023 10743
rect 5216 10736 5243 10743
rect 4996 10687 5003 10736
rect 5216 10687 5223 10736
rect 5276 10716 5283 10773
rect 5216 10563 5223 10673
rect 5256 10667 5263 10703
rect 5296 10696 5303 10753
rect 5316 10667 5323 10833
rect 5216 10556 5233 10563
rect 4716 10007 4723 10453
rect 4736 10447 4743 10553
rect 4776 10236 4783 10493
rect 4856 10456 4863 10473
rect 4876 10427 4883 10443
rect 4896 10407 4903 10463
rect 5316 10456 5323 10653
rect 5356 10467 5363 10753
rect 5376 10687 5383 10923
rect 5396 10723 5403 11213
rect 5496 11196 5523 11203
rect 5556 11196 5563 11213
rect 5496 11123 5503 11196
rect 5836 11183 5843 11216
rect 6136 11187 6143 11233
rect 6436 11196 6463 11203
rect 6496 11196 6503 11213
rect 6736 11207 6743 11343
rect 5476 11116 5503 11123
rect 5476 10767 5483 11116
rect 5496 10807 5503 10883
rect 5556 10727 5563 10733
rect 5396 10716 5423 10723
rect 4916 10307 4923 10443
rect 5096 10367 5103 10423
rect 5016 10236 5023 10313
rect 5076 10236 5103 10243
rect 5036 10187 5043 10193
rect 5096 10187 5103 10236
rect 4716 9976 4723 9993
rect 4736 9967 4743 10093
rect 4676 9767 4683 9873
rect 4836 9756 4843 9773
rect 4576 9476 4583 9493
rect 4556 9247 4563 9473
rect 4536 9016 4543 9073
rect 4556 8967 4563 9003
rect 4576 8947 4583 9023
rect 4616 9003 4623 9193
rect 4596 8996 4623 9003
rect 4336 8587 4343 8633
rect 4336 8516 4343 8573
rect 4196 8227 4203 8513
rect 4316 8467 4323 8503
rect 4296 8387 4303 8453
rect 4236 8147 4243 8313
rect 4216 8036 4243 8043
rect 4236 7987 4243 8036
rect 4256 7887 4263 8313
rect 4276 8047 4283 8153
rect 4296 8087 4303 8373
rect 4316 8296 4323 8353
rect 4336 8316 4343 8393
rect 4276 7836 4283 8033
rect 4196 7816 4223 7823
rect 4196 7807 4203 7816
rect 4156 7343 4163 7573
rect 4256 7563 4263 7773
rect 4296 7627 4303 8073
rect 4316 7767 4323 7993
rect 4356 7807 4363 8053
rect 4256 7556 4283 7563
rect 4196 7367 4203 7473
rect 4296 7367 4303 7543
rect 4236 7356 4263 7363
rect 4156 7336 4183 7343
rect 4036 6876 4063 6883
rect 4036 6827 4043 6876
rect 4116 6807 4123 6873
rect 4036 6383 4043 6573
rect 4096 6427 4103 6583
rect 4136 6447 4143 6573
rect 4116 6396 4143 6403
rect 3996 6376 4023 6383
rect 4036 6376 4063 6383
rect 3976 6127 3983 6213
rect 3936 6056 3963 6063
rect 3916 5876 3943 5883
rect 3916 5687 3923 5876
rect 3956 5727 3963 6056
rect 3976 5896 3983 6113
rect 3996 5887 4003 6353
rect 4016 6187 4023 6376
rect 4136 6116 4143 6396
rect 4156 6127 4163 7336
rect 4176 6167 4183 6773
rect 4176 6116 4183 6153
rect 4096 5947 4103 6033
rect 4116 6007 4123 6103
rect 4196 6047 4203 7213
rect 4256 7007 4263 7356
rect 4276 7027 4283 7063
rect 3736 5183 3743 5393
rect 3756 5207 3763 5573
rect 3836 5467 3843 5623
rect 3876 5616 3903 5623
rect 3896 5436 3903 5513
rect 3936 5436 3943 5533
rect 3956 5427 3963 5613
rect 3996 5447 4003 5623
rect 3996 5427 4003 5433
rect 3736 5176 3763 5183
rect 3756 4707 3763 5176
rect 3796 4927 3803 5413
rect 3916 5387 3923 5423
rect 4056 5087 4063 5713
rect 3696 4456 3723 4463
rect 3696 4127 3703 4456
rect 3736 4196 3743 4273
rect 3756 4176 3773 4183
rect 3656 3996 3683 4003
rect 3716 3996 3723 4013
rect 3596 3727 3603 3913
rect 3636 3827 3643 3993
rect 3656 3987 3663 3996
rect 3696 3927 3703 3983
rect 3736 3976 3743 3993
rect 3796 3947 3803 3963
rect 3636 3716 3643 3813
rect 3556 3696 3583 3703
rect 3387 3556 3403 3563
rect 3376 3507 3383 3553
rect 3616 3547 3623 3703
rect 3676 3503 3683 3553
rect 3576 3496 3603 3503
rect 3656 3496 3683 3503
rect 3336 3107 3343 3243
rect 3596 3227 3603 3496
rect 3356 3207 3363 3223
rect 3396 3147 3403 3223
rect 3556 3187 3563 3203
rect 3616 3187 3623 3233
rect 3636 3227 3643 3453
rect 3796 3307 3803 3593
rect 3816 3587 3823 5073
rect 4076 4987 4083 5163
rect 4116 5067 4123 5433
rect 4136 5007 4143 5473
rect 4156 5416 4163 5553
rect 4196 5387 4203 5423
rect 4156 5156 4163 5233
rect 4216 5047 4223 5313
rect 3896 4976 3923 4983
rect 3916 4947 3923 4976
rect 4156 4956 4163 5033
rect 3876 4767 3883 4913
rect 3836 4667 3843 4683
rect 3876 4676 3883 4753
rect 3836 4507 3843 4633
rect 3836 4476 3843 4493
rect 3856 4487 3863 4663
rect 3916 4447 3923 4483
rect 3836 3976 3843 4313
rect 3836 3743 3843 3853
rect 3856 3767 3863 4193
rect 3876 4187 3883 4253
rect 3916 4167 3923 4433
rect 3956 4187 3963 4613
rect 3996 4487 4003 4953
rect 4196 4947 4203 4963
rect 4136 4887 4143 4943
rect 4076 4687 4083 4813
rect 4236 4807 4243 5693
rect 4256 5447 4263 6913
rect 4276 5967 4283 7013
rect 4336 6927 4343 7543
rect 4356 6907 4363 7633
rect 4307 6876 4323 6883
rect 4336 6827 4343 6863
rect 4336 6583 4343 6733
rect 4316 6576 4343 6583
rect 4296 6087 4303 6413
rect 4316 6396 4323 6513
rect 4296 6067 4303 6073
rect 4276 5896 4303 5903
rect 4296 5863 4303 5896
rect 4276 5856 4303 5863
rect 4276 5427 4283 5856
rect 4296 5416 4303 5753
rect 4336 5707 4343 6576
rect 4356 6396 4363 6413
rect 4376 6267 4383 8093
rect 4396 7547 4403 8093
rect 4416 8036 4423 8493
rect 4436 8067 4443 8853
rect 4476 8287 4483 8793
rect 4516 8787 4523 8933
rect 4536 8796 4543 8933
rect 4596 8767 4603 8996
rect 4556 8647 4563 8753
rect 4676 8727 4683 9753
rect 4776 9543 4783 9743
rect 4776 9536 4803 9543
rect 4736 9276 4743 9413
rect 4776 9276 4783 9473
rect 4796 9307 4803 9536
rect 4816 9507 4823 9733
rect 4856 9427 4863 9443
rect 4856 9347 4863 9413
rect 4696 9256 4723 9263
rect 4696 9247 4703 9256
rect 4756 9227 4763 9263
rect 4756 9027 4763 9213
rect 4796 9007 4803 9273
rect 4516 8367 4523 8593
rect 4556 8527 4563 8633
rect 4496 8327 4503 8353
rect 4536 8307 4543 8503
rect 4596 8296 4603 8523
rect 4676 8467 4683 8593
rect 4696 8487 4703 8973
rect 4376 6116 4383 6233
rect 4376 5903 4383 5953
rect 4356 5896 4383 5903
rect 4396 5867 4403 7053
rect 4416 6867 4423 7973
rect 4436 7647 4443 7793
rect 4436 7507 4443 7633
rect 4476 7567 4483 7803
rect 4456 7356 4463 7533
rect 4436 6967 4443 7323
rect 4316 5547 4323 5643
rect 4396 5623 4403 5673
rect 4376 5616 4403 5623
rect 4416 5487 4423 6853
rect 4436 5847 4443 6893
rect 4456 5527 4463 6993
rect 4476 6727 4483 7553
rect 4516 7107 4523 7993
rect 4556 7587 4563 8173
rect 4576 8087 4583 8283
rect 4636 8267 4643 8293
rect 4636 8036 4643 8073
rect 4616 7687 4623 8003
rect 4536 7547 4543 7563
rect 4576 7556 4583 7573
rect 4596 7527 4603 7543
rect 4496 7007 4503 7043
rect 4496 6867 4503 6933
rect 4476 6587 4483 6613
rect 4496 6587 4503 6853
rect 4516 6843 4523 6873
rect 4516 6836 4543 6843
rect 4516 6607 4523 6836
rect 4576 6807 4583 6843
rect 4596 6807 4603 7433
rect 4616 6887 4623 7593
rect 4636 7067 4643 7993
rect 4656 6847 4663 8273
rect 4676 7487 4683 8253
rect 4696 8007 4703 8473
rect 4716 8267 4723 8993
rect 4796 8783 4803 8953
rect 4776 8776 4803 8783
rect 4736 8287 4743 8753
rect 4716 7816 4723 7973
rect 4736 7707 4743 7803
rect 4696 7527 4703 7613
rect 4736 7563 4743 7673
rect 4756 7607 4763 8713
rect 4816 8567 4823 8813
rect 4836 8787 4843 8993
rect 4836 8747 4843 8773
rect 4776 8527 4783 8553
rect 4876 8547 4883 10013
rect 4896 9387 4903 9773
rect 4916 9467 4923 10173
rect 4936 9947 4943 9963
rect 4976 9956 4983 9973
rect 5016 9943 5023 9953
rect 4956 9927 4963 9943
rect 4996 9936 5023 9943
rect 5016 9756 5023 9833
rect 4996 9727 5003 9753
rect 5136 9687 5143 10423
rect 5296 10187 5303 10203
rect 5116 9476 5143 9483
rect 4896 9167 4903 9373
rect 4776 7567 4783 7773
rect 4796 7607 4803 8533
rect 4836 8487 4843 8503
rect 4876 8496 4903 8503
rect 4836 8316 4843 8453
rect 4876 8316 4883 8353
rect 4856 8267 4863 8303
rect 4896 8167 4903 8496
rect 4916 8367 4923 8793
rect 4936 8507 4943 9173
rect 4956 8987 4963 9193
rect 4976 9127 4983 9263
rect 4996 8823 5003 9473
rect 5136 9467 5143 9476
rect 5036 8996 5043 9013
rect 5016 8967 5023 8983
rect 5076 8963 5083 8993
rect 5056 8956 5083 8963
rect 4996 8816 5023 8823
rect 4936 8307 4943 8393
rect 4956 8227 4963 8513
rect 4816 7987 4823 8003
rect 4736 7556 4763 7563
rect 4776 7507 4783 7523
rect 4676 7356 4683 7453
rect 4716 7356 4743 7363
rect 4736 7307 4743 7356
rect 4696 6847 4703 7073
rect 4536 6707 4543 6793
rect 4476 6307 4483 6573
rect 4536 6387 4543 6693
rect 4556 6567 4563 6713
rect 4616 6707 4623 6813
rect 4576 6587 4583 6603
rect 4616 6596 4623 6693
rect 4596 6507 4603 6583
rect 4556 6396 4563 6493
rect 4596 6396 4603 6473
rect 4576 6367 4583 6383
rect 4616 6376 4643 6383
rect 4576 6167 4583 6353
rect 4636 6227 4643 6376
rect 4536 5936 4543 5953
rect 4576 5947 4583 6123
rect 4596 5907 4603 6143
rect 4616 5763 4623 6053
rect 4596 5756 4623 5763
rect 4556 5656 4563 5673
rect 4596 5656 4603 5756
rect 4576 5567 4583 5643
rect 4396 5456 4423 5463
rect 4256 4963 4263 4973
rect 4276 4963 4283 5413
rect 4256 4956 4283 4963
rect 4256 4647 4263 4956
rect 4296 4827 4303 5133
rect 4316 5047 4323 5433
rect 4396 5423 4403 5456
rect 4396 5416 4423 5423
rect 4416 5127 4423 5416
rect 4316 4956 4323 5013
rect 4276 4647 4283 4683
rect 4096 4627 4103 4643
rect 4036 4183 4043 4593
rect 4116 4447 4123 4463
rect 4156 4456 4163 4553
rect 4176 4447 4183 4473
rect 4016 4176 4043 4183
rect 3936 3763 3943 4173
rect 3976 4167 3983 4173
rect 4136 3976 4143 4213
rect 3936 3756 3963 3763
rect 3836 3736 3863 3743
rect 3896 3736 3903 3753
rect 3876 3707 3883 3723
rect 3796 3236 3803 3293
rect 3316 3036 3323 3053
rect 3296 2987 3303 3023
rect 3316 2763 3323 2833
rect 3296 2756 3323 2763
rect 3276 2587 3283 2723
rect 3316 2707 3323 2756
rect 3336 2727 3343 3093
rect 3356 3027 3363 3073
rect 3396 3007 3403 3133
rect 3716 3023 3723 3233
rect 3816 3023 3823 3053
rect 3416 3016 3443 3023
rect 3716 3016 3743 3023
rect 3796 3016 3823 3023
rect 3376 2787 3383 3003
rect 3316 2556 3323 2633
rect 3236 2287 3243 2533
rect 3296 2487 3303 2543
rect 3336 2536 3343 2613
rect 3376 2523 3383 2773
rect 3376 2516 3403 2523
rect 3296 2307 3303 2453
rect 3396 2347 3403 2516
rect 3296 2276 3303 2293
rect 3276 1796 3283 1833
rect 2956 1547 2963 1553
rect 2956 1367 2963 1533
rect 2956 627 2963 1353
rect 2976 567 2983 1113
rect 2736 376 2763 383
rect 2716 136 2723 173
rect 2736 163 2743 376
rect 2996 376 3003 1253
rect 3016 1247 3023 1553
rect 3116 1447 3123 1583
rect 3056 1336 3063 1353
rect 3016 1116 3023 1233
rect 3056 1116 3063 1133
rect 3076 1127 3083 1323
rect 3136 1087 3143 1093
rect 3016 807 3023 1053
rect 3016 603 3023 693
rect 3036 643 3043 793
rect 3036 636 3063 643
rect 3056 616 3063 636
rect 3016 596 3043 603
rect 3076 596 3083 633
rect 3096 616 3103 873
rect 3056 383 3063 393
rect 3036 376 3063 383
rect 2776 347 2783 363
rect 2936 207 2943 373
rect 2736 156 2763 163
rect 2936 156 2943 193
rect 2956 176 2963 213
rect 2976 156 2983 173
rect 2756 123 2763 156
rect 2296 116 2323 123
rect 2696 107 2703 123
rect 2736 116 2763 123
rect 3056 107 3063 376
rect 3116 167 3123 813
rect 3136 387 3143 1073
rect 3156 787 3163 1433
rect 3196 1347 3203 1733
rect 3216 1367 3223 1763
rect 3236 1627 3243 1773
rect 3176 1207 3183 1333
rect 3176 807 3183 833
rect 3196 827 3203 1333
rect 3296 1307 3303 2113
rect 3316 2107 3323 2293
rect 3356 2276 3363 2293
rect 3396 2076 3403 2133
rect 3416 2047 3423 2973
rect 3436 2887 3443 3016
rect 3436 2767 3443 2873
rect 3736 2767 3743 3016
rect 3436 2536 3443 2753
rect 3536 2727 3543 2743
rect 3516 2627 3523 2723
rect 3556 2576 3563 2593
rect 3436 2107 3443 2273
rect 3356 1787 3363 2033
rect 3356 1576 3363 1593
rect 3396 1563 3403 1753
rect 3376 1556 3403 1563
rect 3276 1287 3283 1303
rect 3236 1107 3243 1213
rect 3336 1116 3343 1273
rect 3396 1107 3403 1556
rect 3216 647 3223 913
rect 3236 823 3243 1093
rect 3316 1047 3323 1103
rect 3396 967 3403 1093
rect 3236 816 3263 823
rect 3256 807 3263 816
rect 3336 787 3343 823
rect 3276 636 3283 653
rect 3296 607 3303 623
rect 3336 616 3343 653
rect 3176 176 3183 413
rect 3256 356 3263 373
rect 3276 307 3283 343
rect 3456 187 3463 2573
rect 3616 2227 3623 2243
rect 3616 2056 3623 2193
rect 3536 1796 3563 1803
rect 3496 1307 3503 1593
rect 3516 1447 3523 1763
rect 3556 1727 3563 1796
rect 3576 1647 3583 2033
rect 3596 1887 3603 2043
rect 3576 1616 3583 1633
rect 3556 1596 3563 1613
rect 3516 1227 3523 1333
rect 3536 1267 3543 1303
rect 3556 1227 3563 1283
rect 3576 1187 3583 1293
rect 3496 643 3503 1153
rect 3556 1136 3563 1173
rect 3516 1116 3543 1123
rect 3516 1087 3523 1116
rect 3616 1107 3623 1433
rect 3536 827 3543 1073
rect 3556 1027 3563 1093
rect 3556 856 3563 1013
rect 3516 807 3523 823
rect 3576 787 3583 823
rect 3496 636 3523 643
rect 3476 387 3483 633
rect 3636 627 3643 1313
rect 3536 343 3543 613
rect 3156 156 3163 173
rect 3376 156 3403 163
rect 3416 156 3423 173
rect 3476 167 3483 343
rect 3516 336 3543 343
rect 3396 -17 3403 156
rect 3616 156 3643 163
rect 3656 156 3663 1873
rect 3716 1843 3723 2613
rect 3736 2547 3743 2753
rect 3756 2267 3763 2723
rect 3816 2527 3823 2543
rect 3776 2296 3783 2333
rect 3796 2047 3803 2333
rect 3816 2287 3823 2393
rect 3816 2076 3823 2113
rect 3856 2076 3863 2213
rect 3876 2207 3883 2533
rect 3896 2076 3903 2313
rect 3916 2307 3923 3533
rect 3956 2687 3963 3756
rect 3976 2567 3983 3453
rect 4036 3087 4043 3813
rect 4036 3023 4043 3073
rect 4016 3016 4043 3023
rect 3976 2367 3983 2553
rect 3996 2307 4003 3013
rect 4016 2756 4023 2793
rect 4056 2556 4063 2593
rect 4076 2587 4083 3833
rect 4116 3716 4123 3753
rect 4096 3667 4103 3703
rect 4156 3687 4163 3723
rect 4176 3707 4183 4033
rect 4096 3516 4103 3533
rect 4156 3487 4163 3653
rect 4096 2767 4103 3473
rect 4196 3467 4203 4473
rect 4236 4183 4243 4553
rect 4256 4227 4263 4633
rect 4216 4176 4243 4183
rect 4216 3967 4223 3983
rect 4216 3527 4223 3953
rect 4236 3747 4243 4176
rect 4116 3223 4123 3253
rect 4116 3216 4143 3223
rect 4156 3167 4163 3203
rect 4176 3167 4183 3223
rect 4256 3207 4263 4183
rect 4276 3787 4283 4213
rect 4296 3987 4303 4813
rect 4316 3847 4323 4773
rect 4276 3063 4283 3773
rect 4336 3767 4343 4993
rect 4356 4676 4383 4683
rect 4376 4647 4383 4676
rect 4416 4667 4423 4893
rect 4416 4527 4423 4653
rect 4376 4496 4383 4513
rect 4396 4447 4403 4463
rect 4436 4287 4443 4873
rect 4456 4247 4463 5093
rect 4476 4467 4483 5073
rect 4396 4183 4403 4213
rect 4396 4176 4423 4183
rect 4356 3736 4363 4133
rect 4476 3963 4483 3993
rect 4456 3956 4483 3963
rect 4416 3867 4423 3953
rect 4396 3736 4423 3743
rect 4316 3496 4323 3733
rect 4416 3687 4423 3736
rect 4456 3707 4463 3956
rect 4496 3887 4503 5033
rect 4296 3127 4303 3483
rect 4336 3447 4343 3483
rect 4376 3236 4383 3673
rect 4416 3507 4423 3673
rect 4276 3056 4303 3063
rect 4296 3036 4303 3056
rect 4216 3016 4233 3023
rect 4216 2807 4223 3016
rect 4096 2556 4103 2753
rect 4276 2747 4283 3023
rect 4256 2587 4263 2723
rect 4256 2527 4263 2573
rect 4296 2556 4303 2633
rect 4336 2556 4343 3073
rect 4376 2556 4383 3113
rect 4396 3067 4403 3203
rect 4416 2687 4423 2743
rect 4416 2627 4423 2673
rect 4316 2507 4323 2543
rect 4036 2287 4043 2393
rect 4076 2307 4083 2333
rect 3936 2247 3943 2273
rect 3956 2087 3963 2263
rect 3716 1836 3743 1843
rect 3676 1816 3703 1823
rect 3736 1816 3743 1836
rect 3676 1627 3683 1816
rect 3876 1807 3883 2063
rect 3916 1927 3923 2053
rect 3996 2023 4003 2233
rect 4236 2227 4243 2243
rect 4276 2107 4283 2173
rect 3976 2016 4003 2023
rect 4076 2096 4103 2103
rect 3976 1807 3983 2016
rect 3716 1787 3723 1803
rect 4016 1796 4023 1813
rect 3676 1167 3683 1613
rect 3736 603 3743 993
rect 3756 867 3763 1633
rect 3856 1596 3863 1653
rect 3876 1607 3883 1793
rect 3816 1336 3843 1343
rect 3796 1096 3803 1113
rect 3776 887 3783 1083
rect 3836 1067 3843 1336
rect 3936 1327 3943 1793
rect 4056 1783 4063 1853
rect 4076 1787 4083 2096
rect 4276 2056 4283 2093
rect 4376 2063 4383 2093
rect 4356 2056 4383 2063
rect 4296 1803 4303 1913
rect 4276 1796 4303 1803
rect 4036 1776 4063 1783
rect 3956 1747 3963 1773
rect 4196 1707 4203 1793
rect 3996 1303 4003 1653
rect 4056 1596 4063 1613
rect 4216 1607 4223 1783
rect 4356 1767 4363 1913
rect 4396 1827 4403 2533
rect 4436 2467 4443 3433
rect 4496 3016 4503 3713
rect 4516 3567 4523 5033
rect 4576 4987 4583 5513
rect 4616 5387 4623 5756
rect 4636 5447 4643 6073
rect 4616 5207 4623 5373
rect 4596 5087 4603 5123
rect 4596 4956 4603 5013
rect 4576 4936 4583 4953
rect 4616 4927 4623 4943
rect 4596 4683 4603 4833
rect 4656 4747 4663 6813
rect 4676 6616 4683 6633
rect 4676 5907 4683 6493
rect 4696 5967 4703 6693
rect 4716 6687 4723 6853
rect 4716 6667 4723 6673
rect 4716 6567 4723 6603
rect 4576 4676 4603 4683
rect 4536 3967 4543 4453
rect 4596 4267 4603 4676
rect 4616 4476 4623 4533
rect 4676 4323 4683 4683
rect 4696 4607 4703 5853
rect 4716 4907 4723 6533
rect 4736 6007 4743 7033
rect 4756 7027 4763 7063
rect 4796 6896 4803 7493
rect 4816 7147 4823 7543
rect 4856 7407 4863 8153
rect 4976 7867 4983 8533
rect 5016 8507 5023 8816
rect 5056 8647 5063 8956
rect 5096 8867 5103 9443
rect 5096 8767 5103 8853
rect 5056 8523 5063 8633
rect 5116 8587 5123 9013
rect 5136 9007 5143 9233
rect 5056 8516 5083 8523
rect 5116 8516 5123 8573
rect 4996 8207 5003 8433
rect 5016 7987 5023 8393
rect 5076 8367 5083 8516
rect 5116 8316 5123 8433
rect 5156 8316 5163 9953
rect 5176 9747 5183 9923
rect 5296 9847 5303 10173
rect 5316 9987 5323 10013
rect 5256 9787 5263 9813
rect 5256 9756 5263 9773
rect 5276 9727 5283 9743
rect 5316 9736 5323 9973
rect 5396 9943 5403 10693
rect 5416 9987 5423 10716
rect 5456 10187 5463 10673
rect 5476 10207 5483 10713
rect 5556 10696 5563 10713
rect 5496 10647 5503 10683
rect 5516 10423 5523 10453
rect 5556 10436 5563 10453
rect 5636 10423 5643 10713
rect 5516 10416 5543 10423
rect 5436 9956 5443 9973
rect 5396 9936 5423 9943
rect 5436 9916 5463 9923
rect 5276 9667 5283 9713
rect 5256 9227 5263 9253
rect 5296 9127 5303 9453
rect 5336 9447 5343 9463
rect 5336 9247 5343 9433
rect 5176 8667 5183 9113
rect 5276 8996 5283 9113
rect 5356 8983 5363 9733
rect 5376 9027 5383 9773
rect 5436 9487 5443 9916
rect 5456 9276 5463 9793
rect 5496 9503 5503 10413
rect 5576 10407 5583 10423
rect 5616 10416 5643 10423
rect 5656 10463 5663 10933
rect 5696 10923 5703 11153
rect 5796 11127 5803 11183
rect 5836 11176 5863 11183
rect 5916 11176 5943 11183
rect 5916 11167 5923 11176
rect 6216 11176 6243 11183
rect 6216 11047 6223 11176
rect 5687 10916 5703 10923
rect 5656 10456 5683 10463
rect 5536 10216 5543 10353
rect 5516 10187 5523 10203
rect 5516 9807 5523 10173
rect 5556 10083 5563 10193
rect 5536 10076 5563 10083
rect 5536 9756 5543 10076
rect 5576 9787 5583 10253
rect 5596 9967 5603 10233
rect 5576 9756 5583 9773
rect 5556 9723 5563 9743
rect 5556 9716 5583 9723
rect 5476 9496 5503 9503
rect 5476 9303 5483 9496
rect 5556 9467 5563 9483
rect 5496 9447 5503 9463
rect 5476 9296 5503 9303
rect 5496 9287 5503 9296
rect 5416 9256 5443 9263
rect 5336 8976 5363 8983
rect 5216 8796 5223 8853
rect 5036 8247 5043 8313
rect 5096 8227 5103 8303
rect 5136 8287 5143 8303
rect 4976 7807 4983 7853
rect 4916 7787 4923 7803
rect 4956 7796 4973 7803
rect 5056 7707 5063 7833
rect 4816 7087 4823 7113
rect 4836 6903 4843 7353
rect 4856 7047 4863 7393
rect 4876 7047 4883 7593
rect 4936 7527 4943 7633
rect 4976 7447 4983 7573
rect 4996 7543 5003 7693
rect 5076 7587 5083 8023
rect 5136 8003 5143 8273
rect 5116 7996 5143 8003
rect 4996 7536 5023 7543
rect 4976 7347 4983 7433
rect 4896 7067 4903 7273
rect 4836 6896 4863 6903
rect 4856 6867 4863 6896
rect 4756 5987 4763 6453
rect 4776 6087 4783 6453
rect 4796 6416 4803 6433
rect 4816 6427 4823 6833
rect 4876 6787 4883 7033
rect 4916 6707 4923 7293
rect 4936 7287 4943 7313
rect 4936 7007 4943 7113
rect 4956 6787 4963 7133
rect 4996 7087 5003 7333
rect 5076 7327 5083 7373
rect 5096 7367 5103 7973
rect 5016 7096 5023 7193
rect 4976 7027 4983 7063
rect 5056 6867 5063 7133
rect 5076 7067 5083 7193
rect 5116 7027 5123 7996
rect 5176 7843 5183 8333
rect 5196 7967 5203 8033
rect 5156 7836 5183 7843
rect 5196 7836 5203 7853
rect 5136 7356 5143 7733
rect 5156 7387 5163 7836
rect 5176 7687 5183 7803
rect 5176 7356 5183 7533
rect 5196 7447 5203 7633
rect 5216 7503 5223 8553
rect 5236 7523 5243 8493
rect 5256 7947 5263 8173
rect 5276 8167 5283 8473
rect 5276 8047 5283 8113
rect 5256 7556 5263 7653
rect 5276 7647 5283 7953
rect 5296 7787 5303 8963
rect 5316 8503 5323 8953
rect 5376 8847 5383 9013
rect 5356 8516 5363 8593
rect 5396 8527 5403 9113
rect 5416 8967 5423 9256
rect 5476 8987 5483 9253
rect 5476 8816 5503 8823
rect 5316 8496 5343 8503
rect 5376 8476 5403 8483
rect 5356 8296 5363 8473
rect 5316 8283 5323 8293
rect 5316 8276 5343 8283
rect 5356 8047 5363 8253
rect 5316 7823 5323 7933
rect 5336 7847 5343 8023
rect 5376 8007 5383 8023
rect 5396 8007 5403 8476
rect 5416 8007 5423 8793
rect 5436 8783 5443 8793
rect 5436 8776 5463 8783
rect 5496 8627 5503 8816
rect 5496 8547 5503 8613
rect 5436 8027 5443 8513
rect 5516 8487 5523 9393
rect 5536 9307 5543 9463
rect 5576 9267 5583 9716
rect 5596 9527 5603 9953
rect 5596 9447 5603 9513
rect 5616 9407 5623 10193
rect 5656 10007 5663 10456
rect 5696 10427 5703 10916
rect 5756 10916 5783 10923
rect 5716 10083 5723 10443
rect 5736 10267 5743 10913
rect 5776 10867 5783 10916
rect 6016 10916 6023 10933
rect 6056 10907 6063 10933
rect 5956 10767 5963 10903
rect 5996 10827 6003 10903
rect 6036 10847 6043 10903
rect 6216 10887 6223 11033
rect 6336 10943 6343 11153
rect 6436 11147 6443 11196
rect 6776 11187 6783 11233
rect 6976 11207 6983 11343
rect 6476 11127 6483 11183
rect 6716 11147 6723 11163
rect 6956 11147 6963 11163
rect 6336 10936 6363 10943
rect 6236 10767 6243 10923
rect 6276 10916 6283 10933
rect 6296 10896 6323 10903
rect 6036 10707 6043 10713
rect 5776 10687 5783 10703
rect 6076 10696 6083 10733
rect 6016 10667 6023 10683
rect 5976 10407 5983 10453
rect 6016 10427 6023 10443
rect 6016 10347 6023 10413
rect 5716 10076 5733 10083
rect 5776 9987 5783 10153
rect 5636 9507 5643 9943
rect 5716 9727 5723 9973
rect 5776 9763 5783 9973
rect 5816 9967 5823 10213
rect 5756 9756 5783 9763
rect 5576 9227 5583 9253
rect 5556 8996 5563 9193
rect 5616 9023 5623 9273
rect 5636 9207 5643 9493
rect 5616 9016 5643 9023
rect 5576 8947 5583 8963
rect 5556 8487 5563 8793
rect 5576 8587 5583 8933
rect 5616 8787 5623 8993
rect 5596 8516 5603 8773
rect 5636 8567 5643 9016
rect 5656 8987 5663 9713
rect 5696 9276 5703 9713
rect 5776 9667 5783 9756
rect 5716 9107 5723 9253
rect 5756 9247 5763 9263
rect 5776 9207 5783 9463
rect 5796 9436 5813 9443
rect 5676 8796 5683 9093
rect 5656 8776 5663 8793
rect 5576 8407 5583 8503
rect 5316 7816 5343 7823
rect 5296 7556 5303 7573
rect 5236 7516 5263 7523
rect 5216 7496 5243 7503
rect 5156 7307 5163 7343
rect 5196 7327 5203 7343
rect 5236 7287 5243 7496
rect 5256 7367 5263 7516
rect 5276 7507 5283 7523
rect 5076 6876 5083 7013
rect 5116 6876 5123 6913
rect 4996 6467 5003 6853
rect 5096 6727 5103 6863
rect 5016 6587 5023 6603
rect 5096 6596 5103 6633
rect 5136 6487 5143 7093
rect 5156 6647 5163 7273
rect 5256 7227 5263 7353
rect 5276 7287 5283 7493
rect 5316 7487 5323 7543
rect 5336 7527 5343 7816
rect 5196 7063 5203 7173
rect 5276 7076 5283 7093
rect 5196 7056 5223 7063
rect 5196 6963 5203 7056
rect 5316 7007 5323 7373
rect 5336 7187 5343 7313
rect 5356 7147 5363 7993
rect 5396 7856 5403 7893
rect 5176 6956 5203 6963
rect 4816 6107 4823 6383
rect 4876 6307 4883 6363
rect 4836 6067 4843 6103
rect 4756 5916 4763 5973
rect 4856 5907 4863 6083
rect 4876 5927 4883 6033
rect 4796 5643 4803 5693
rect 4776 5636 4803 5643
rect 4736 5167 4743 5373
rect 4756 4867 4763 5493
rect 4776 4727 4783 5636
rect 4816 5567 4823 5603
rect 4816 5247 4823 5553
rect 4836 5183 4843 5473
rect 4856 5427 4863 5873
rect 4876 5463 4883 5913
rect 4896 5487 4903 6433
rect 5036 6416 5043 6453
rect 4916 6376 4943 6383
rect 4936 6247 4943 6376
rect 5036 5916 5043 6373
rect 5176 6363 5183 6956
rect 5296 6887 5303 6933
rect 5336 6876 5343 6953
rect 5356 6923 5363 7053
rect 5376 6943 5383 7453
rect 5396 7347 5403 7573
rect 5416 7356 5423 7593
rect 5436 7467 5443 7993
rect 5456 7947 5463 8273
rect 5456 7547 5463 7833
rect 5456 7356 5463 7513
rect 5476 7387 5483 8373
rect 5516 8307 5523 8313
rect 5516 8127 5523 8293
rect 5536 8107 5543 8313
rect 5576 8283 5583 8353
rect 5596 8316 5603 8473
rect 5636 8387 5643 8473
rect 5636 8336 5643 8373
rect 5616 8287 5623 8303
rect 5576 8276 5603 8283
rect 5556 8047 5563 8173
rect 5576 8036 5583 8173
rect 5496 7607 5503 8013
rect 5536 7807 5543 8033
rect 5516 7607 5523 7793
rect 5556 7667 5563 8003
rect 5576 7667 5583 7913
rect 5516 7447 5523 7563
rect 5556 7556 5563 7573
rect 5596 7543 5603 8276
rect 5616 7783 5623 8113
rect 5636 7907 5643 8113
rect 5656 8027 5663 8303
rect 5676 8287 5683 8533
rect 5676 8247 5683 8273
rect 5696 7967 5703 8733
rect 5716 7987 5723 8553
rect 5736 7987 5743 9013
rect 5756 8787 5763 9033
rect 5776 8867 5783 9193
rect 5756 8567 5763 8673
rect 5676 7907 5683 7953
rect 5716 7927 5723 7973
rect 5636 7816 5643 7873
rect 5716 7843 5723 7913
rect 5696 7836 5723 7843
rect 5736 7827 5743 7853
rect 5676 7803 5683 7823
rect 5676 7796 5703 7803
rect 5616 7776 5643 7783
rect 5616 7547 5623 7673
rect 5576 7536 5603 7543
rect 5436 7327 5443 7343
rect 5516 7287 5523 7413
rect 5536 7327 5543 7413
rect 5396 6967 5403 7253
rect 5376 6936 5403 6943
rect 5356 6916 5383 6923
rect 5376 6887 5383 6916
rect 5196 6447 5203 6873
rect 5236 6587 5243 6773
rect 5216 6407 5223 6573
rect 5216 6376 5223 6393
rect 5176 6356 5203 6363
rect 5096 6123 5103 6253
rect 5096 6116 5123 6123
rect 5036 5876 5063 5883
rect 4996 5643 5003 5713
rect 4976 5636 5003 5643
rect 4876 5456 4903 5463
rect 4896 5436 4903 5456
rect 4916 5427 4923 5473
rect 4956 5436 4963 5633
rect 4816 5176 4843 5183
rect 4816 4976 4823 5176
rect 4856 5156 4863 5353
rect 4936 5347 4943 5423
rect 4876 5147 4883 5333
rect 4896 5187 4903 5293
rect 4836 4787 4843 4943
rect 4936 4936 4943 5273
rect 4896 4867 4903 4923
rect 4956 4867 4963 5393
rect 4976 5247 4983 5636
rect 5036 5603 5043 5876
rect 5076 5687 5083 6103
rect 5116 5947 5123 6116
rect 5096 5916 5123 5923
rect 5116 5887 5123 5916
rect 5196 5827 5203 6356
rect 5236 6207 5243 6573
rect 5256 6123 5263 6873
rect 5276 6787 5283 6833
rect 5356 6647 5363 6863
rect 5316 6596 5323 6613
rect 5336 6567 5343 6583
rect 5276 6383 5283 6473
rect 5336 6427 5343 6453
rect 5276 6376 5303 6383
rect 5296 6347 5303 6376
rect 5236 6116 5263 6123
rect 5236 5787 5243 6116
rect 5276 6007 5283 6103
rect 5316 6087 5323 6413
rect 5336 5987 5343 6393
rect 5376 6027 5383 6693
rect 5396 6467 5403 6936
rect 5416 6907 5423 7273
rect 5416 6667 5423 6713
rect 5436 6567 5443 6993
rect 5476 6747 5483 7233
rect 5516 7076 5523 7213
rect 5536 6707 5543 7043
rect 5556 6647 5563 7473
rect 5576 7427 5583 7536
rect 5576 6827 5583 7393
rect 5616 7307 5623 7333
rect 5596 6947 5603 7193
rect 5616 6947 5623 7293
rect 5616 6896 5623 6933
rect 5596 6847 5603 6853
rect 5636 6643 5643 7776
rect 5656 7527 5663 7593
rect 5616 6636 5643 6643
rect 5536 6616 5543 6633
rect 5587 6616 5603 6623
rect 5436 6547 5443 6553
rect 5276 5896 5283 5953
rect 5296 5727 5303 5883
rect 5056 5656 5083 5663
rect 5016 5596 5043 5603
rect 4976 5107 4983 5233
rect 5016 5047 5023 5596
rect 4696 4427 4703 4473
rect 4776 4447 4783 4693
rect 4667 4316 4683 4323
rect 4676 3996 4683 4293
rect 4736 4216 4743 4433
rect 4796 4187 4803 4643
rect 4856 4476 4863 4493
rect 4896 4476 4903 4573
rect 4876 4407 4883 4463
rect 4916 4456 4923 4553
rect 4916 4196 4923 4413
rect 4896 4147 4903 4163
rect 4656 3967 4663 3983
rect 4556 3723 4563 3753
rect 4556 3716 4583 3723
rect 4636 3667 4643 3703
rect 4516 3447 4523 3483
rect 4536 3003 4543 3053
rect 4456 2547 4463 2733
rect 4476 2523 4483 3003
rect 4516 2996 4543 3003
rect 4456 2516 4483 2523
rect 4416 2187 4423 2283
rect 4436 1787 4443 2233
rect 4456 1867 4463 2516
rect 3996 1296 4023 1303
rect 4056 1247 4063 1303
rect 3996 1083 4003 1193
rect 4036 1096 4043 1133
rect 3996 1076 4023 1083
rect 3756 823 3763 853
rect 3796 836 3803 933
rect 3756 816 3783 823
rect 3776 647 3783 653
rect 3776 616 3783 633
rect 3736 596 3763 603
rect 3796 387 3803 603
rect 3816 343 3823 823
rect 3836 807 3843 833
rect 3736 207 3743 343
rect 3796 336 3823 343
rect 3836 327 3843 793
rect 3856 227 3863 1073
rect 4056 927 4063 1083
rect 4016 703 4023 823
rect 4036 787 4043 803
rect 4016 696 4043 703
rect 3976 656 3983 673
rect 4016 636 4023 673
rect 3956 376 3963 393
rect 3976 347 3983 363
rect 4036 347 4043 696
rect 4056 367 4063 813
rect 4076 627 4083 773
rect 4196 687 4203 1313
rect 4216 1307 4223 1593
rect 4276 1576 4283 1653
rect 4476 1647 4483 2353
rect 4516 1887 4523 2913
rect 4576 2747 4583 3653
rect 4596 3407 4603 3573
rect 4556 2556 4563 2593
rect 4596 2583 4603 3243
rect 4676 3227 4683 3253
rect 4636 2587 4643 3033
rect 4696 2783 4703 3713
rect 4716 3483 4723 4113
rect 4916 3996 4923 4033
rect 4856 3907 4863 3993
rect 4936 3967 4943 3983
rect 4856 3716 4863 3773
rect 4896 3716 4903 3733
rect 4936 3703 4943 3833
rect 4836 3687 4843 3703
rect 4876 3687 4883 3703
rect 4916 3696 4943 3703
rect 4716 3476 4743 3483
rect 4736 3327 4743 3476
rect 4776 3467 4783 3483
rect 4816 3467 4823 3513
rect 4716 3167 4723 3233
rect 4756 3036 4783 3043
rect 4776 3027 4783 3036
rect 4676 2776 4703 2783
rect 4656 2727 4663 2743
rect 4596 2576 4623 2583
rect 4616 2563 4623 2576
rect 4616 2556 4643 2563
rect 4576 1867 4583 2063
rect 4516 1796 4523 1833
rect 4556 1796 4563 1813
rect 4596 1807 4603 2373
rect 4616 1816 4623 2033
rect 4596 1783 4603 1793
rect 4496 1747 4503 1783
rect 4536 1747 4543 1783
rect 4576 1776 4603 1783
rect 4496 1707 4503 1733
rect 4256 1547 4263 1563
rect 4296 1447 4303 1563
rect 4296 1267 4303 1303
rect 4316 1287 4323 1323
rect 4236 1147 4243 1153
rect 4216 787 4223 833
rect 4236 803 4243 823
rect 4236 796 4263 803
rect 4256 623 4263 796
rect 4236 616 4263 623
rect 4276 363 4283 653
rect 4356 387 4363 1633
rect 4376 407 4383 1593
rect 4476 1567 4483 1613
rect 4536 1596 4543 1633
rect 4396 687 4403 1113
rect 4416 983 4423 1233
rect 4436 1083 4443 1533
rect 4516 1327 4523 1433
rect 4636 1323 4643 2556
rect 4676 2287 4683 2776
rect 4716 2276 4723 2313
rect 4676 2243 4683 2273
rect 4676 2236 4703 2243
rect 4656 1767 4663 1803
rect 4676 1667 4683 2073
rect 4736 2067 4743 2553
rect 4776 2547 4783 2553
rect 4796 2547 4803 3233
rect 4816 3203 4823 3453
rect 4816 3196 4843 3203
rect 4856 3016 4883 3023
rect 4816 2747 4823 3003
rect 4876 2887 4883 3016
rect 4816 2647 4823 2733
rect 4816 2556 4823 2573
rect 4776 2276 4783 2533
rect 4796 2076 4803 2213
rect 4776 1847 4783 2063
rect 4836 2047 4843 2393
rect 4876 2283 4883 2853
rect 4956 2783 4963 4793
rect 4976 4667 4983 4683
rect 4976 3996 4983 4013
rect 4996 3967 5003 3983
rect 5016 3727 5023 4753
rect 5036 4627 5043 5413
rect 5056 5367 5063 5593
rect 5076 5407 5083 5656
rect 5096 5287 5103 5643
rect 5196 5627 5203 5653
rect 5376 5643 5383 5973
rect 5376 5636 5403 5643
rect 5156 5456 5163 5473
rect 5196 5436 5203 5513
rect 5396 5503 5403 5636
rect 5396 5496 5423 5503
rect 5187 5276 5193 5283
rect 5216 5187 5223 5413
rect 5136 5047 5143 5143
rect 5176 5136 5203 5143
rect 5056 4976 5063 5033
rect 5196 4947 5203 5136
rect 5216 5087 5223 5153
rect 5236 4943 5243 5173
rect 5336 4943 5343 4993
rect 5216 4936 5243 4943
rect 5316 4936 5343 4943
rect 5056 4676 5063 4693
rect 5216 4667 5223 4936
rect 5016 3516 5023 3653
rect 5036 3647 5043 4593
rect 5056 4456 5063 4633
rect 5076 4307 5083 4493
rect 5096 4427 5103 4613
rect 5256 4607 5263 4663
rect 5296 4627 5303 4663
rect 5356 4487 5363 5193
rect 5396 5143 5403 5423
rect 5416 5187 5423 5496
rect 5436 5387 5443 6493
rect 5476 6396 5483 6433
rect 5516 6396 5523 6413
rect 5496 6367 5503 6383
rect 5596 6367 5603 6616
rect 5496 5936 5503 6193
rect 5096 4183 5103 4213
rect 5096 4176 5123 4183
rect 5056 3767 5063 4033
rect 4996 3467 5003 3503
rect 5056 3243 5063 3733
rect 5076 3387 5083 3973
rect 5116 3667 5123 3703
rect 5156 3607 5163 4183
rect 5176 4007 5183 4333
rect 5256 4327 5263 4453
rect 5216 3996 5223 4293
rect 5376 4227 5383 5143
rect 5396 5136 5423 5143
rect 5416 4747 5423 4853
rect 5416 4443 5423 4733
rect 5396 4436 5423 4443
rect 5436 4307 5443 5133
rect 5456 4587 5463 5933
rect 5516 5803 5523 5903
rect 5496 5796 5523 5803
rect 5476 5636 5483 5653
rect 5496 5083 5503 5796
rect 5516 5347 5523 5773
rect 5476 5076 5503 5083
rect 5256 3996 5263 4013
rect 5196 3723 5203 3953
rect 5236 3947 5243 3983
rect 5196 3716 5223 3723
rect 5036 3236 5063 3243
rect 5036 3127 5043 3236
rect 5096 3203 5103 3513
rect 5176 3507 5183 3633
rect 5216 3563 5223 3716
rect 5196 3556 5223 3563
rect 5076 3196 5103 3203
rect 5096 3123 5103 3196
rect 5096 3116 5123 3123
rect 4976 3056 4983 3073
rect 5116 3027 5123 3116
rect 5136 2907 5143 3473
rect 5176 3047 5183 3493
rect 5156 3016 5183 3023
rect 4956 2776 4983 2783
rect 4936 2743 4943 2773
rect 4976 2743 4983 2776
rect 4916 2736 4943 2743
rect 4956 2736 4983 2743
rect 4916 2407 4923 2736
rect 4956 2727 4963 2736
rect 5056 2587 5063 2893
rect 5116 2767 5123 2793
rect 5136 2747 5143 2873
rect 5176 2867 5183 3016
rect 5196 2807 5203 3556
rect 5256 3536 5263 3873
rect 5276 3547 5283 4013
rect 5316 3547 5323 4213
rect 5336 4167 5343 4183
rect 5396 3996 5423 4003
rect 5456 3996 5463 4533
rect 5476 4007 5483 5076
rect 5496 4647 5503 5053
rect 5536 5027 5543 6173
rect 5556 5467 5563 6293
rect 5576 5667 5583 5713
rect 5576 5463 5583 5653
rect 5596 5607 5603 5733
rect 5616 5667 5623 6636
rect 5576 5456 5603 5463
rect 5516 4976 5523 4993
rect 5576 4927 5583 5456
rect 5616 5307 5623 5423
rect 5616 5156 5623 5173
rect 5516 4696 5523 4913
rect 5567 4696 5583 4703
rect 5516 4387 5523 4573
rect 5216 2783 5223 3533
rect 5296 3516 5323 3523
rect 5276 3487 5283 3503
rect 5316 3467 5323 3516
rect 5236 3256 5263 3263
rect 5296 3256 5303 3273
rect 5236 3187 5243 3256
rect 5196 2776 5223 2783
rect 5196 2767 5203 2776
rect 5016 2536 5043 2543
rect 5016 2387 5023 2536
rect 5056 2516 5063 2573
rect 5116 2523 5123 2573
rect 5176 2547 5183 2743
rect 5096 2516 5123 2523
rect 5196 2307 5203 2633
rect 5216 2467 5223 2743
rect 4856 2276 4883 2283
rect 4856 2187 4863 2276
rect 5036 2227 5043 2243
rect 4716 1607 4723 1673
rect 4756 1607 4763 1813
rect 4936 1803 4943 2173
rect 5156 2167 5163 2283
rect 5196 2147 5203 2153
rect 5016 2096 5043 2103
rect 4936 1796 4963 1803
rect 4776 1747 4783 1763
rect 4636 1316 4663 1323
rect 4476 1096 4483 1113
rect 4436 1076 4463 1083
rect 4496 1027 4503 1083
rect 4416 976 4443 983
rect 4416 827 4423 933
rect 4436 636 4443 976
rect 4456 656 4463 833
rect 4476 643 4483 1013
rect 4516 847 4523 1313
rect 4636 1303 4643 1316
rect 4536 1087 4543 1293
rect 4576 1287 4583 1303
rect 4616 1296 4643 1303
rect 4496 767 4503 823
rect 4476 636 4503 643
rect 4496 407 4503 636
rect 4536 607 4543 813
rect 4676 767 4683 1593
rect 4936 1327 4943 1796
rect 4976 1596 4983 1693
rect 5016 1596 5023 2096
rect 5196 2067 5203 2133
rect 5216 2056 5223 2173
rect 5196 1927 5203 2053
rect 5036 1796 5063 1803
rect 5056 1767 5063 1796
rect 4996 1547 5003 1583
rect 5076 1343 5083 1813
rect 5096 1607 5103 1893
rect 5196 1787 5203 1913
rect 5236 1847 5243 2853
rect 5276 1867 5283 2753
rect 5296 2747 5303 2763
rect 5316 2727 5323 3033
rect 5336 2927 5343 3993
rect 5396 3987 5403 3996
rect 5476 3976 5503 3983
rect 5496 3947 5503 3976
rect 5496 3767 5503 3933
rect 5376 3716 5383 3733
rect 5356 3563 5363 3713
rect 5516 3707 5523 4373
rect 5536 4167 5543 4653
rect 5576 4647 5583 4696
rect 5556 3987 5563 4573
rect 5596 4207 5603 4993
rect 5616 4476 5623 5073
rect 5636 4907 5643 6113
rect 5656 5387 5663 7093
rect 5676 7047 5683 7553
rect 5696 7487 5703 7796
rect 5716 7607 5723 7813
rect 5716 7523 5723 7573
rect 5756 7567 5763 8553
rect 5796 8507 5803 9373
rect 5836 8543 5843 9773
rect 5856 9487 5863 10233
rect 5896 10216 5903 10333
rect 6196 10216 6203 10533
rect 6236 10427 6243 10753
rect 6276 10736 6283 10833
rect 6256 10716 6263 10733
rect 6316 10707 6323 10896
rect 6356 10687 6363 10936
rect 6376 10887 6383 10923
rect 6396 10487 6403 10933
rect 6476 10887 6483 10913
rect 6676 10907 6683 10923
rect 6496 10827 6503 10883
rect 6276 10427 6283 10443
rect 6236 10147 6243 10203
rect 5876 9967 5883 10073
rect 5856 9047 5863 9473
rect 5896 9447 5903 9963
rect 5936 9956 5943 9973
rect 5956 9767 5963 9943
rect 5956 9727 5963 9753
rect 5956 9276 5963 9673
rect 5976 9387 5983 10113
rect 5996 10007 6003 10133
rect 5996 9976 6003 9993
rect 6016 9667 6023 9743
rect 6056 9736 6063 9773
rect 5996 9276 6003 9453
rect 5976 9207 5983 9263
rect 5936 9027 5943 9153
rect 5996 9127 6003 9153
rect 5876 8996 5883 9013
rect 5936 8983 5943 9013
rect 5956 9007 5963 9053
rect 5916 8976 5943 8983
rect 5856 8647 5863 8973
rect 5936 8796 5943 8893
rect 5976 8796 5983 8813
rect 5996 8807 6003 9113
rect 6096 9087 6103 9473
rect 5816 8536 5843 8543
rect 5796 8147 5803 8253
rect 5816 8147 5823 8536
rect 5856 8516 5863 8533
rect 5916 8467 5923 8773
rect 5856 8363 5863 8453
rect 5836 8356 5863 8363
rect 5836 8316 5843 8356
rect 5876 8316 5903 8323
rect 5776 7747 5783 8093
rect 5836 8067 5843 8273
rect 5876 8023 5883 8133
rect 5896 8067 5903 8316
rect 5916 8027 5923 8053
rect 5936 8027 5943 8493
rect 5956 8487 5963 8783
rect 5976 8487 5983 8533
rect 5856 8016 5883 8023
rect 5796 7587 5803 8013
rect 5776 7556 5783 7573
rect 5716 7516 5743 7523
rect 5696 7356 5703 7373
rect 5736 7356 5743 7516
rect 5776 7356 5783 7393
rect 5716 7187 5723 7343
rect 5796 7323 5803 7353
rect 5776 7316 5803 7323
rect 5676 6927 5683 7033
rect 5696 6867 5703 7173
rect 5776 7107 5783 7316
rect 5776 7076 5783 7093
rect 5716 6927 5723 7013
rect 5676 6307 5683 6633
rect 5736 6407 5743 6973
rect 5796 6887 5803 7063
rect 5816 7047 5823 7973
rect 5836 7627 5843 7853
rect 5856 7836 5863 7873
rect 5876 7867 5883 8016
rect 5936 8007 5943 8013
rect 5956 8007 5963 8053
rect 5996 7987 6003 8453
rect 5876 7807 5883 7823
rect 5856 7783 5863 7793
rect 5856 7776 5883 7783
rect 5856 7427 5863 7513
rect 5756 6583 5763 6873
rect 5816 6827 5823 6853
rect 5836 6727 5843 7273
rect 5856 6847 5863 7073
rect 5756 6576 5783 6583
rect 5796 6547 5803 6563
rect 5816 6427 5823 6583
rect 5836 6547 5843 6613
rect 5736 6347 5743 6363
rect 5776 6107 5783 6353
rect 5716 5947 5723 6103
rect 5816 5987 5823 6393
rect 5736 5916 5743 5973
rect 5756 5747 5763 5903
rect 5676 5607 5683 5623
rect 5676 4667 5683 5553
rect 5716 5127 5723 5633
rect 5696 4956 5723 4963
rect 5696 4807 5703 4956
rect 5696 4463 5703 4713
rect 5636 4347 5643 4463
rect 5676 4456 5703 4463
rect 5636 4187 5643 4273
rect 5576 4167 5583 4183
rect 5436 3687 5443 3703
rect 5356 3556 5383 3563
rect 5356 2867 5363 3533
rect 5376 3027 5383 3556
rect 5536 3516 5543 3913
rect 5556 3787 5563 3973
rect 5556 3627 5563 3773
rect 5576 3647 5583 4153
rect 5596 4147 5603 4163
rect 5596 3747 5603 4133
rect 5676 4027 5683 4456
rect 5616 3687 5623 3973
rect 5676 3807 5683 3983
rect 5636 3736 5663 3743
rect 5696 3736 5703 3873
rect 5636 3687 5643 3736
rect 5576 3516 5583 3533
rect 5596 3507 5603 3633
rect 5556 3447 5563 3503
rect 5456 3203 5463 3273
rect 5536 3236 5543 3253
rect 5456 3196 5483 3203
rect 5496 3187 5503 3223
rect 5396 3036 5423 3043
rect 5396 3007 5403 3036
rect 5396 2687 5403 2993
rect 5616 2763 5623 3553
rect 5596 2756 5623 2763
rect 5356 2556 5363 2673
rect 5556 2627 5563 2653
rect 5556 2556 5563 2613
rect 5616 2587 5623 2756
rect 5636 2647 5643 3593
rect 5716 3427 5723 4793
rect 5736 4727 5743 5473
rect 5756 5156 5763 5273
rect 5776 5047 5783 5873
rect 5756 4956 5783 4963
rect 5776 4747 5783 4956
rect 5796 4887 5803 5793
rect 5816 5567 5823 5893
rect 5836 5887 5843 6153
rect 5856 5767 5863 6533
rect 5876 5647 5883 7776
rect 5896 7687 5903 7733
rect 5876 5403 5883 5453
rect 5816 5087 5823 5403
rect 5856 5396 5883 5403
rect 5876 5187 5883 5353
rect 5776 4676 5783 4713
rect 5756 3996 5763 4663
rect 5796 4647 5803 4663
rect 5796 4527 5803 4633
rect 5296 2487 5303 2543
rect 5296 2147 5303 2283
rect 5596 2187 5603 2283
rect 5656 2103 5663 3353
rect 5736 3287 5743 3983
rect 5776 3587 5783 4473
rect 5816 4267 5823 5033
rect 5836 4707 5843 4973
rect 5836 4676 5843 4693
rect 5876 4687 5883 5173
rect 5896 4947 5903 7413
rect 5916 6527 5923 7753
rect 5936 7207 5943 7553
rect 5976 7507 5983 7833
rect 6016 7767 6023 8513
rect 6036 8507 6043 9033
rect 6116 8567 6123 9833
rect 6136 9487 6143 9953
rect 6316 9947 6323 10443
rect 6356 9963 6363 10413
rect 6336 9956 6363 9963
rect 6156 9827 6163 9923
rect 6376 9903 6383 10273
rect 6396 9956 6423 9963
rect 6396 9947 6403 9956
rect 6356 9896 6383 9903
rect 6316 9756 6323 9813
rect 6356 9787 6363 9896
rect 6356 9756 6363 9773
rect 6216 9476 6223 9493
rect 6236 9447 6243 9463
rect 6236 9303 6243 9433
rect 6236 9296 6263 9303
rect 6136 8907 6143 9003
rect 6176 8996 6183 9213
rect 6196 8967 6203 8983
rect 6216 8943 6223 9053
rect 6196 8936 6223 8943
rect 6156 8796 6163 8833
rect 6196 8796 6203 8936
rect 6236 8803 6243 9253
rect 6276 9087 6283 9263
rect 6236 8796 6263 8803
rect 6176 8763 6183 8783
rect 6176 8756 6203 8763
rect 6196 8707 6203 8756
rect 6076 8516 6083 8533
rect 6047 8496 6063 8503
rect 6136 8496 6163 8503
rect 6036 8327 6043 8373
rect 6056 8316 6063 8353
rect 6096 8316 6103 8453
rect 6136 8316 6143 8353
rect 6076 8147 6083 8293
rect 6116 8287 6123 8303
rect 6096 8107 6103 8273
rect 6076 8007 6083 8023
rect 5996 7383 6003 7573
rect 6036 7407 6043 7933
rect 6076 7643 6083 7773
rect 6096 7767 6103 8043
rect 6116 8007 6123 8273
rect 6136 7867 6143 8133
rect 6156 8107 6163 8496
rect 6176 8287 6183 8533
rect 6196 8527 6203 8693
rect 6216 8547 6223 8783
rect 6196 8307 6203 8513
rect 6176 8083 6183 8133
rect 6207 8096 6213 8103
rect 6156 8076 6183 8083
rect 6116 7836 6123 7853
rect 6156 7836 6163 8076
rect 6216 8007 6223 8073
rect 6196 7836 6223 7843
rect 6136 7807 6143 7823
rect 6116 7647 6123 7793
rect 6076 7636 6103 7643
rect 5996 7376 6023 7383
rect 5956 7343 5963 7373
rect 5956 7336 5983 7343
rect 5936 6507 5943 7173
rect 5956 7067 5963 7213
rect 6016 7207 6023 7376
rect 6056 7247 6063 7543
rect 6076 7327 6083 7613
rect 5996 7076 6003 7113
rect 6076 7087 6083 7313
rect 5976 7047 5983 7063
rect 5956 6447 5963 7033
rect 6076 6876 6083 6953
rect 6016 6787 6023 6853
rect 6056 6847 6063 6863
rect 5976 6487 5983 6753
rect 6036 6647 6043 6793
rect 5976 6376 5983 6413
rect 6016 6363 6023 6473
rect 6056 6367 6063 6413
rect 5996 6356 6023 6363
rect 5956 6116 5963 6293
rect 5976 6047 5983 6103
rect 6016 5943 6023 6233
rect 6036 6107 6043 6133
rect 6056 6067 6063 6353
rect 5996 5936 6023 5943
rect 6036 5916 6063 5923
rect 5976 5767 5983 5893
rect 5936 5647 5943 5673
rect 5956 5636 5963 5653
rect 5916 5307 5923 5633
rect 5996 5623 6003 5893
rect 6016 5867 6023 5903
rect 6056 5867 6063 5916
rect 6036 5707 6043 5773
rect 5976 5616 6003 5623
rect 5936 5587 5943 5603
rect 5976 5367 5983 5616
rect 6016 5287 6023 5673
rect 6076 5507 6083 6773
rect 6096 5987 6103 7636
rect 6116 7107 6123 7633
rect 6156 7547 6163 7633
rect 6216 7527 6223 7836
rect 6196 7356 6203 7433
rect 6236 7407 6243 8573
rect 6256 7887 6263 8796
rect 6276 8087 6283 8813
rect 6296 8587 6303 9233
rect 6316 8727 6323 9693
rect 6336 9267 6343 9733
rect 6396 9247 6403 9933
rect 6416 9467 6423 9493
rect 6436 9367 6443 10753
rect 6576 10607 6583 10713
rect 6456 10216 6463 10453
rect 6556 10407 6563 10423
rect 6476 10236 6483 10253
rect 6516 10236 6523 10273
rect 6456 9687 6463 10153
rect 6536 9776 6543 9933
rect 6576 9823 6583 10593
rect 6676 10427 6683 10893
rect 6976 10887 6983 10903
rect 6736 10487 6743 10703
rect 6796 10436 6803 10733
rect 6916 10716 6943 10723
rect 6916 10683 6923 10716
rect 6996 10696 7003 10913
rect 7016 10707 7023 11293
rect 7136 11167 7143 11343
rect 7176 11307 7183 11343
rect 7276 11187 7283 11213
rect 7436 11207 7443 11343
rect 8156 11307 8163 11343
rect 8156 11196 8163 11213
rect 7556 11176 7583 11183
rect 7236 11147 7243 11153
rect 7256 10927 7263 11173
rect 7416 10907 7423 11153
rect 7176 10867 7183 10903
rect 7216 10747 7223 10753
rect 7396 10707 7403 10893
rect 7416 10887 7423 10893
rect 7456 10747 7463 10903
rect 7496 10703 7503 10733
rect 7476 10696 7503 10703
rect 6916 10676 6943 10683
rect 6856 10436 6883 10443
rect 6676 10236 6703 10243
rect 6736 10236 6743 10253
rect 6676 10207 6683 10236
rect 6676 10007 6683 10193
rect 6596 9967 6603 9973
rect 6576 9816 6603 9823
rect 6456 9496 6463 9653
rect 6576 9507 6583 9793
rect 6456 9367 6463 9413
rect 6476 9387 6483 9483
rect 6516 9407 6523 9483
rect 6456 9296 6463 9353
rect 6436 9167 6443 9263
rect 6476 9187 6483 9263
rect 6396 8987 6403 9033
rect 6416 9016 6423 9113
rect 6516 9087 6523 9373
rect 6516 8987 6523 9073
rect 6296 8507 6303 8553
rect 6316 8507 6323 8673
rect 6336 8523 6343 8913
rect 6416 8747 6423 8783
rect 6336 8516 6363 8523
rect 6296 8063 6303 8353
rect 6356 8316 6363 8373
rect 6376 8287 6383 8303
rect 6276 8056 6303 8063
rect 6276 8023 6283 8056
rect 6356 8036 6383 8043
rect 6276 8016 6303 8023
rect 6256 7687 6263 7853
rect 6296 7807 6303 7993
rect 6336 7827 6343 8023
rect 6296 7707 6303 7753
rect 6296 7556 6303 7693
rect 6276 7527 6283 7543
rect 6276 7343 6283 7393
rect 6216 7267 6223 7343
rect 6256 7336 6283 7343
rect 6296 7227 6303 7493
rect 6116 6807 6123 6853
rect 6116 6187 6123 6713
rect 6136 6427 6143 6933
rect 6156 6407 6163 7033
rect 6176 6856 6203 6863
rect 6176 6767 6183 6856
rect 6156 6307 6163 6393
rect 6176 6167 6183 6693
rect 6216 6667 6223 7113
rect 6276 7096 6283 7213
rect 6316 7187 6323 7543
rect 6356 7487 6363 8013
rect 6376 7907 6383 8036
rect 6416 7947 6423 8493
rect 6436 8467 6443 8693
rect 6456 8507 6463 8833
rect 6496 8783 6503 8813
rect 6476 8776 6503 8783
rect 6456 8163 6463 8473
rect 6476 8183 6483 8776
rect 6496 8487 6503 8753
rect 6516 8327 6523 8893
rect 6536 8507 6543 9133
rect 6596 8847 6603 9816
rect 6616 9447 6623 9913
rect 6676 9827 6683 9953
rect 6716 9947 6723 10223
rect 6756 10127 6763 10213
rect 6656 9467 6663 9753
rect 6676 9427 6683 9813
rect 6816 9743 6823 10433
rect 6836 10407 6843 10423
rect 6876 10167 6883 10436
rect 6896 10267 6903 10413
rect 6936 10047 6943 10676
rect 7036 10567 7043 10693
rect 7056 10487 7063 10673
rect 7516 10487 7523 11163
rect 7576 11047 7583 11176
rect 7836 11176 7863 11183
rect 7676 10747 7683 10883
rect 7836 10727 7843 11176
rect 7936 11107 7943 11183
rect 8136 11127 8143 11183
rect 8196 11167 8203 11293
rect 8156 10936 8163 11153
rect 8196 10947 8203 10953
rect 8116 10907 8123 10933
rect 8216 10927 8223 11173
rect 8336 10947 8343 11343
rect 11256 11216 11283 11223
rect 8456 11196 8483 11203
rect 8376 11183 8383 11193
rect 8376 11176 8403 11183
rect 8376 10967 8383 11176
rect 8376 10936 8383 10953
rect 7816 10467 7823 10703
rect 7836 10463 7843 10473
rect 7836 10456 7863 10463
rect 7496 10427 7503 10443
rect 7116 10407 7123 10423
rect 7096 10307 7103 10403
rect 6967 10236 6983 10243
rect 6856 9956 6863 9973
rect 6776 9527 6783 9743
rect 6816 9736 6843 9743
rect 6716 9476 6723 9513
rect 6616 8987 6623 9033
rect 6636 8983 6643 9413
rect 6676 9047 6683 9373
rect 6736 9307 6743 9393
rect 6836 9387 6843 9736
rect 6916 9467 6923 9773
rect 6736 9276 6743 9293
rect 6776 9276 6783 9293
rect 6716 9256 6723 9273
rect 6756 9227 6763 9263
rect 6676 8996 6683 9033
rect 6816 8987 6823 9233
rect 6836 9187 6843 9293
rect 6636 8976 6663 8983
rect 6656 8907 6663 8976
rect 6816 8867 6823 8953
rect 6736 8816 6743 8833
rect 6836 8827 6843 9173
rect 6916 9127 6923 9253
rect 6916 8983 6923 9113
rect 6936 8987 6943 10033
rect 6956 9947 6963 10233
rect 6996 9463 7003 9953
rect 7076 9923 7083 10213
rect 7116 10167 7123 10393
rect 7196 10236 7203 10413
rect 7316 10387 7323 10423
rect 7256 10227 7263 10273
rect 7216 10167 7223 10223
rect 7116 9956 7143 9963
rect 7076 9916 7103 9923
rect 7016 9756 7023 9773
rect 7056 9756 7063 9793
rect 7096 9756 7123 9763
rect 7116 9747 7123 9756
rect 7036 9727 7043 9743
rect 7136 9727 7143 9956
rect 7276 9776 7283 9993
rect 7296 9943 7303 10233
rect 7356 10227 7363 10423
rect 7816 10423 7823 10453
rect 7796 10416 7823 10423
rect 7676 10347 7683 10403
rect 7336 9956 7343 9973
rect 7416 9943 7423 10213
rect 7436 9947 7443 9973
rect 7476 9967 7483 10223
rect 7296 9936 7323 9943
rect 6976 9456 7003 9463
rect 6996 9347 7003 9456
rect 6996 9256 7003 9293
rect 6896 8976 6923 8983
rect 6876 8947 6883 8963
rect 6896 8907 6903 8976
rect 6596 8747 6603 8813
rect 6836 8776 6863 8783
rect 6556 8407 6563 8493
rect 6476 8176 6503 8183
rect 6456 8156 6483 8163
rect 6436 7856 6443 7873
rect 6376 7836 6403 7843
rect 6376 7587 6383 7836
rect 6356 7447 6363 7473
rect 6336 7347 6343 7373
rect 6376 6896 6383 6953
rect 6416 6947 6423 7453
rect 6436 7387 6443 7733
rect 6476 7587 6483 8156
rect 6496 7887 6503 8176
rect 6496 7827 6503 7853
rect 6516 7747 6523 8313
rect 6536 8207 6543 8313
rect 6556 8247 6563 8333
rect 6576 8227 6583 8513
rect 6616 8507 6623 8523
rect 6636 8467 6643 8503
rect 6596 8316 6603 8393
rect 6616 8267 6623 8303
rect 6676 8227 6683 8333
rect 6716 8327 6723 8513
rect 6736 8287 6743 8433
rect 6756 8423 6763 8753
rect 6836 8647 6843 8776
rect 6836 8516 6863 8523
rect 6796 8447 6803 8493
rect 6756 8416 6783 8423
rect 6576 8187 6583 8213
rect 6536 8036 6563 8043
rect 6596 8036 6603 8053
rect 6536 7787 6543 8036
rect 6576 7887 6583 8003
rect 6556 7583 6563 7873
rect 6536 7576 6563 7583
rect 6496 7356 6503 7393
rect 6536 7356 6543 7576
rect 6556 7467 6563 7553
rect 6576 7407 6583 7713
rect 6476 7247 6483 7343
rect 6456 7047 6463 7073
rect 6476 6987 6483 7233
rect 6516 7187 6523 7333
rect 6556 7307 6563 7393
rect 6496 7007 6503 7113
rect 6536 7076 6543 7213
rect 6576 7076 6583 7113
rect 6516 7007 6523 7063
rect 6496 6987 6503 6993
rect 6196 6483 6203 6613
rect 6216 6503 6223 6653
rect 6256 6596 6283 6603
rect 6236 6527 6243 6563
rect 6276 6507 6283 6596
rect 6216 6496 6243 6503
rect 6196 6476 6223 6483
rect 6216 6416 6223 6476
rect 6236 6403 6243 6496
rect 6236 6396 6263 6403
rect 6256 6367 6263 6396
rect 6316 6247 6323 6753
rect 6396 6727 6403 6853
rect 6176 6136 6183 6153
rect 6276 6116 6283 6153
rect 6116 5903 6123 6073
rect 6176 5907 6183 6093
rect 6336 6007 6343 6713
rect 6356 6407 6363 6633
rect 6496 6596 6503 6813
rect 6516 6727 6523 6993
rect 6556 6907 6563 7043
rect 6416 6427 6423 6593
rect 6436 6567 6443 6583
rect 6516 6507 6523 6583
rect 6476 6267 6483 6383
rect 6536 6307 6543 6843
rect 6356 6107 6363 6123
rect 6376 6107 6383 6233
rect 6556 6227 6563 6513
rect 6596 6407 6603 7993
rect 6616 7836 6623 7913
rect 6656 7836 6663 7893
rect 6676 7867 6683 8213
rect 6716 8107 6723 8253
rect 6716 7843 6723 8093
rect 6696 7836 6723 7843
rect 6636 7803 6643 7823
rect 6627 7796 6643 7803
rect 6576 6376 6603 6383
rect 6576 6247 6583 6376
rect 6616 6283 6623 7793
rect 6636 6367 6643 7573
rect 6656 7507 6663 7673
rect 6676 7547 6683 7813
rect 6736 7707 6743 8033
rect 6756 7927 6763 8333
rect 6716 7556 6723 7593
rect 6736 7567 6743 7693
rect 6756 7627 6763 7913
rect 6776 7647 6783 8416
rect 6796 8067 6803 8413
rect 6816 8347 6823 8493
rect 6836 8483 6843 8516
rect 6916 8487 6923 8503
rect 6836 8476 6863 8483
rect 6856 8347 6863 8476
rect 6876 8427 6883 8473
rect 6916 8387 6923 8433
rect 6936 8367 6943 8793
rect 6876 8316 6883 8333
rect 6856 8287 6863 8303
rect 6816 8027 6823 8043
rect 6836 8007 6843 8023
rect 6816 7807 6823 7873
rect 6756 7556 6763 7593
rect 6696 7503 6703 7543
rect 6676 7496 6703 7503
rect 6676 7287 6683 7496
rect 6736 7487 6743 7513
rect 6696 7367 6703 7473
rect 6776 7423 6783 7593
rect 6796 7576 6803 7633
rect 6796 7503 6803 7533
rect 6816 7527 6823 7793
rect 6836 7627 6843 7853
rect 6836 7507 6843 7563
rect 6796 7496 6823 7503
rect 6776 7416 6803 7423
rect 6696 7067 6703 7353
rect 6736 7336 6743 7353
rect 6776 7336 6783 7393
rect 6776 7247 6783 7293
rect 6796 7147 6803 7416
rect 6816 7147 6823 7496
rect 6676 6547 6683 6593
rect 6696 6547 6703 7053
rect 6716 6627 6723 7093
rect 6796 7076 6803 7093
rect 6836 7063 6843 7373
rect 6776 6883 6783 7063
rect 6816 7056 6843 7063
rect 6776 6876 6803 6883
rect 6776 6807 6783 6843
rect 6796 6627 6803 6876
rect 6756 6596 6763 6613
rect 6736 6527 6743 6583
rect 6816 6567 6823 6893
rect 6856 6667 6863 7833
rect 6876 7767 6883 8023
rect 6916 7847 6923 8353
rect 6976 7943 6983 9033
rect 7016 8967 7023 9073
rect 6996 8487 7003 8513
rect 7016 8507 7023 8913
rect 7036 8807 7043 9333
rect 7016 8387 7023 8473
rect 7016 8247 7023 8293
rect 6976 7936 7003 7943
rect 6976 7803 6983 7913
rect 6956 7796 6983 7803
rect 6996 7687 7003 7936
rect 7016 7667 7023 7793
rect 7036 7747 7043 8773
rect 7056 8767 7063 9493
rect 7116 9467 7123 9483
rect 7136 9227 7143 9593
rect 7356 9587 7363 9943
rect 7396 9936 7423 9943
rect 7316 9443 7323 9573
rect 7296 9436 7323 9443
rect 7396 9303 7403 9936
rect 7416 9907 7423 9936
rect 7576 9827 7583 9973
rect 7716 9947 7723 10333
rect 7576 9756 7583 9813
rect 7636 9767 7643 9923
rect 7496 9487 7503 9613
rect 7516 9507 7523 9673
rect 7556 9607 7563 9743
rect 7736 9687 7743 10113
rect 7756 9767 7763 10253
rect 7776 9903 7783 9953
rect 7796 9927 7803 10416
rect 7856 10127 7863 10456
rect 7876 10447 7883 10553
rect 7896 10387 7903 10903
rect 8176 10783 8183 10923
rect 8156 10776 8183 10783
rect 7956 10696 7963 10713
rect 7876 10236 7883 10273
rect 7956 10223 7963 10253
rect 7936 10216 7963 10223
rect 7836 9956 7843 9973
rect 7816 9907 7823 9943
rect 7916 9943 7923 10193
rect 7896 9936 7923 9943
rect 7936 9923 7943 10173
rect 7916 9916 7943 9923
rect 7776 9896 7803 9903
rect 7776 9776 7783 9873
rect 7796 9756 7803 9896
rect 7396 9296 7423 9303
rect 7196 9276 7203 9293
rect 7236 9276 7263 9283
rect 7096 8943 7103 8973
rect 7076 8936 7103 8943
rect 7076 8743 7083 8936
rect 7116 8827 7123 8993
rect 7056 8736 7083 8743
rect 7056 7667 7063 8736
rect 7096 8507 7103 8813
rect 7116 8796 7123 8813
rect 7156 8796 7163 9033
rect 7176 8847 7183 9273
rect 7256 9087 7263 9276
rect 7376 9267 7383 9293
rect 7396 9227 7403 9296
rect 7416 9276 7423 9296
rect 7436 9187 7443 9263
rect 7196 8807 7203 8853
rect 7136 8747 7143 8783
rect 7136 8516 7143 8733
rect 7176 8547 7183 8783
rect 7176 8516 7183 8533
rect 7116 8487 7123 8503
rect 7156 8487 7163 8503
rect 7076 8107 7083 8393
rect 7096 8367 7103 8413
rect 7116 8316 7123 8393
rect 7156 8316 7183 8323
rect 7136 8207 7143 8303
rect 7116 8047 7123 8173
rect 7176 8067 7183 8316
rect 7096 7847 7103 8023
rect 7136 8003 7143 8013
rect 7116 7996 7143 8003
rect 6876 7347 6883 7393
rect 6896 6767 6903 7353
rect 6916 7347 6923 7473
rect 6916 7007 6923 7093
rect 6936 6727 6943 7613
rect 7056 7427 7063 7453
rect 6956 7356 6963 7413
rect 6996 7287 7003 7313
rect 6956 7067 6963 7113
rect 6956 6847 6963 7053
rect 6976 7047 6983 7233
rect 7016 7076 7023 7093
rect 7056 7047 7063 7083
rect 6996 6876 7003 6953
rect 7016 6847 7023 6863
rect 6956 6563 6963 6813
rect 6976 6607 6983 6793
rect 6956 6556 6983 6563
rect 6776 6416 6783 6453
rect 6616 6276 6643 6283
rect 6556 6147 6563 6153
rect 6536 6047 6543 6083
rect 6096 5896 6123 5903
rect 6356 5727 6363 5893
rect 6096 5436 6103 5573
rect 6116 5527 6123 5653
rect 6136 5636 6163 5643
rect 6196 5636 6203 5653
rect 6136 5487 6143 5636
rect 6136 5427 6143 5473
rect 5976 5156 5983 5173
rect 5956 5107 5963 5143
rect 5976 4976 5983 5053
rect 6016 4956 6023 5153
rect 6056 5147 6063 5393
rect 6076 5167 6083 5423
rect 6156 5367 6163 5413
rect 6096 5147 6103 5173
rect 6056 4947 6063 5113
rect 5856 4496 5863 4533
rect 5896 4507 5903 4913
rect 5896 4463 5903 4493
rect 5876 4456 5903 4463
rect 5796 3567 5803 4233
rect 5816 3647 5823 4053
rect 5756 3516 5783 3523
rect 5816 3516 5823 3613
rect 5756 3287 5763 3516
rect 5716 3256 5743 3263
rect 5716 3247 5723 3256
rect 5716 2767 5723 2993
rect 5756 2787 5763 3243
rect 5636 2096 5663 2103
rect 5696 2096 5703 2473
rect 5716 2307 5723 2553
rect 5316 2063 5323 2093
rect 5296 2056 5323 2063
rect 5316 1827 5323 2033
rect 5496 1907 5503 2053
rect 5216 1587 5223 1613
rect 5236 1596 5243 1653
rect 5276 1596 5283 1693
rect 5256 1547 5263 1583
rect 5296 1576 5303 1613
rect 5076 1336 5103 1343
rect 4696 1247 4703 1313
rect 4916 1267 4923 1283
rect 4736 1116 4743 1153
rect 4776 856 4803 863
rect 4716 827 4723 843
rect 4736 823 4743 853
rect 4736 816 4763 823
rect 4676 603 4683 633
rect 4676 596 4703 603
rect 4356 367 4363 373
rect 4256 356 4283 363
rect 4416 343 4423 393
rect 4536 367 4543 593
rect 4696 376 4703 413
rect 4736 376 4743 433
rect 4756 427 4763 816
rect 4796 787 4803 856
rect 4416 336 4443 343
rect 3976 307 3983 333
rect 4476 247 4483 343
rect 3856 156 3863 213
rect 3896 156 3903 233
rect 4716 227 4723 363
rect 3636 -17 3643 156
rect 4036 127 4043 173
rect 4136 156 4143 213
rect 4816 203 4823 1113
rect 4876 847 4883 1133
rect 4896 1116 4903 1153
rect 4936 1116 4943 1173
rect 4876 447 4883 833
rect 4916 636 4923 893
rect 4956 843 4963 873
rect 4956 836 4983 843
rect 5016 827 5023 843
rect 5056 827 5063 1133
rect 4996 636 5023 643
rect 4976 607 4983 623
rect 5016 607 5023 636
rect 4976 427 4983 593
rect 5096 587 5103 1336
rect 5116 1116 5143 1123
rect 5176 1116 5203 1123
rect 5116 767 5123 1116
rect 5196 887 5203 1116
rect 5216 1107 5223 1333
rect 5236 1327 5243 1433
rect 5256 1327 5263 1533
rect 5336 1363 5343 1833
rect 5356 1787 5363 1803
rect 5476 1707 5483 1763
rect 5456 1587 5463 1633
rect 5476 1596 5503 1603
rect 5476 1567 5483 1596
rect 5636 1587 5643 2096
rect 5656 2076 5683 2083
rect 5716 2076 5723 2293
rect 5656 2027 5663 2076
rect 5656 1787 5663 1803
rect 5756 1787 5763 2573
rect 5776 2067 5783 2693
rect 5796 2567 5803 3193
rect 5816 2287 5823 3273
rect 5836 2603 5843 3893
rect 5856 3007 5863 4153
rect 5876 3907 5883 4253
rect 5916 4007 5923 4473
rect 5936 4467 5943 4933
rect 5956 4827 5963 4943
rect 5996 4927 6003 4943
rect 6196 4727 6203 5573
rect 6216 5467 6223 5623
rect 6216 5067 6223 5143
rect 6236 4983 6243 5653
rect 6296 5436 6303 5553
rect 6336 5436 6343 5533
rect 6376 5463 6383 5993
rect 6456 5683 6463 5973
rect 6476 5896 6503 5903
rect 6496 5767 6503 5896
rect 6516 5767 6523 5883
rect 6436 5676 6463 5683
rect 6436 5656 6443 5676
rect 6476 5656 6483 5753
rect 6356 5456 6383 5463
rect 6267 5416 6283 5423
rect 6256 5287 6263 5413
rect 6316 5367 6323 5423
rect 6216 4976 6243 4983
rect 6216 4967 6223 4976
rect 5956 4207 5963 4553
rect 5936 3996 5943 4193
rect 5976 3996 5983 4373
rect 5956 3927 5963 3983
rect 5896 3716 5903 3733
rect 5936 3727 5943 3753
rect 5876 3487 5883 3703
rect 5916 3627 5923 3683
rect 5916 3016 5923 3493
rect 5876 2647 5883 2743
rect 5896 2707 5903 3003
rect 5956 2947 5963 3613
rect 5916 2607 5923 2743
rect 5836 2596 5863 2603
rect 5836 2556 5843 2573
rect 5836 1803 5843 2493
rect 5856 1823 5863 2596
rect 5916 2527 5923 2593
rect 5916 2276 5923 2293
rect 5956 2263 5963 2513
rect 5976 2407 5983 3733
rect 6016 3367 6023 4553
rect 6076 4476 6083 4513
rect 6076 4196 6083 4253
rect 6056 3516 6063 4113
rect 6156 3747 6163 4593
rect 6116 3663 6123 3703
rect 6116 3656 6143 3663
rect 6096 3516 6103 3553
rect 6076 3487 6083 3503
rect 5996 3147 6003 3243
rect 6036 3236 6043 3293
rect 6016 3167 6023 3223
rect 6056 3187 6063 3223
rect 5896 1927 5903 2263
rect 5936 2256 5963 2263
rect 5976 2096 5983 2373
rect 5996 2063 6003 2293
rect 5856 1816 5883 1823
rect 5836 1796 5863 1803
rect 5476 1367 5483 1553
rect 5336 1356 5363 1363
rect 5316 1336 5333 1343
rect 5336 1067 5343 1333
rect 5196 843 5203 873
rect 5196 836 5223 843
rect 5236 807 5243 863
rect 5276 856 5283 993
rect 4936 387 4943 393
rect 4936 356 4943 373
rect 4996 356 5003 393
rect 4796 196 4823 203
rect 4316 167 4323 173
rect 4556 156 4563 173
rect 4316 123 4323 153
rect 4356 136 4363 153
rect 4796 127 4803 196
rect 4816 156 4823 173
rect 4856 156 4863 353
rect 5016 327 5023 343
rect 5176 323 5183 793
rect 5196 616 5203 693
rect 5256 687 5263 753
rect 5216 636 5223 653
rect 5256 636 5263 673
rect 5236 603 5243 623
rect 5216 596 5243 603
rect 5216 356 5223 596
rect 5316 347 5323 653
rect 5176 316 5203 323
rect 5076 136 5083 173
rect 4316 116 4343 123
rect 5096 116 5103 193
rect 5336 176 5343 213
rect 3376 -24 3403 -17
rect 3616 -24 3643 -17
rect 5356 -17 5363 1356
rect 5476 1336 5503 1343
rect 5476 1227 5483 1336
rect 5396 1136 5403 1213
rect 5456 1107 5463 1133
rect 5376 1067 5383 1103
rect 5436 887 5443 1013
rect 5436 843 5443 873
rect 5436 836 5463 843
rect 5476 827 5483 863
rect 5516 856 5523 873
rect 5416 603 5423 813
rect 5496 807 5503 843
rect 5496 603 5503 793
rect 5576 747 5583 833
rect 5596 827 5603 1233
rect 5616 1116 5643 1123
rect 5676 1116 5693 1123
rect 5416 596 5443 603
rect 5476 596 5503 603
rect 5396 363 5403 413
rect 5476 376 5483 413
rect 5616 387 5623 1116
rect 5696 727 5703 1113
rect 5716 747 5723 1773
rect 5756 1596 5763 1633
rect 5796 1596 5803 1753
rect 5836 1607 5843 1773
rect 5856 1587 5863 1796
rect 5776 1447 5783 1583
rect 5736 1336 5743 1353
rect 5776 1336 5803 1343
rect 5756 1267 5763 1323
rect 5796 1307 5803 1336
rect 5876 1147 5883 1816
rect 5916 1247 5923 2063
rect 5976 2056 6003 2063
rect 5976 1967 5983 2056
rect 5976 1796 5983 1953
rect 5956 1627 5963 1783
rect 6016 1727 6023 2553
rect 6036 2247 6043 2993
rect 6056 2747 6063 3173
rect 6116 3167 6123 3573
rect 6136 3467 6143 3656
rect 6076 2576 6083 3093
rect 6136 3056 6143 3133
rect 6156 3107 6163 3553
rect 6056 2267 6063 2543
rect 6096 2287 6103 2733
rect 6116 2307 6123 2723
rect 6136 2487 6143 2743
rect 6156 2507 6163 3023
rect 6176 3007 6183 4413
rect 6196 4016 6203 4473
rect 6216 4307 6223 4683
rect 6236 4507 6243 4933
rect 6296 4903 6303 5133
rect 6276 4896 6303 4903
rect 6256 4696 6263 4733
rect 6216 3267 6223 3983
rect 6236 3967 6243 4493
rect 6236 3247 6243 3653
rect 6276 3607 6283 4896
rect 6316 4667 6323 5353
rect 6336 4607 6343 5393
rect 6316 4443 6323 4513
rect 6356 4487 6363 5456
rect 6376 5387 6383 5423
rect 6376 4627 6383 5193
rect 6316 4436 6343 4443
rect 6296 4216 6303 4253
rect 6376 4167 6383 4433
rect 6336 3736 6343 4133
rect 6376 3736 6383 3793
rect 6276 3496 6283 3573
rect 6356 3487 6363 3723
rect 6336 3467 6343 3483
rect 6356 3267 6363 3473
rect 6096 2256 6123 2263
rect 6096 1807 6103 2256
rect 6156 2103 6163 2253
rect 6176 2127 6183 2553
rect 6196 2367 6203 3233
rect 6276 3227 6283 3243
rect 6216 3187 6223 3223
rect 6216 2527 6223 3033
rect 6296 2567 6303 3253
rect 6196 2107 6203 2353
rect 6236 2287 6243 2513
rect 6136 2096 6163 2103
rect 5976 1207 5983 1593
rect 6016 1316 6023 1433
rect 6116 1327 6123 1813
rect 5896 1136 5913 1143
rect 5736 787 5743 843
rect 5776 836 5783 1133
rect 5916 1116 5943 1123
rect 5736 636 5743 713
rect 5756 687 5763 823
rect 5796 807 5803 823
rect 5936 767 5943 1116
rect 6036 927 6043 1303
rect 6136 1167 6143 2096
rect 6216 2103 6223 2273
rect 6216 2096 6243 2103
rect 6236 2076 6243 2096
rect 6156 2063 6163 2073
rect 6156 2056 6183 2063
rect 6156 2007 6163 2056
rect 6056 836 6063 1153
rect 6136 1136 6163 1143
rect 6096 1127 6103 1133
rect 5996 767 6003 813
rect 6076 807 6083 823
rect 5716 567 5723 623
rect 5396 356 5423 363
rect 5456 327 5463 363
rect 5756 347 5763 633
rect 5816 616 5843 623
rect 5776 587 5783 603
rect 5836 487 5843 616
rect 5736 336 5753 343
rect 5696 327 5703 333
rect 5496 136 5503 193
rect 5716 187 5723 323
rect 5516 116 5523 173
rect 5756 167 5763 213
rect 5796 156 5803 173
rect 6016 167 6023 473
rect 6096 387 6103 833
rect 6116 727 6123 733
rect 6116 616 6123 713
rect 6156 707 6163 1136
rect 6176 623 6183 2013
rect 6216 1787 6223 1973
rect 6196 1307 6203 1773
rect 6256 1643 6263 2113
rect 6236 1636 6263 1643
rect 6196 1047 6203 1133
rect 6176 616 6203 623
rect 6196 547 6203 616
rect 6136 376 6143 393
rect 5536 136 5543 153
rect 5776 127 5783 143
rect 5816 136 5823 153
rect 6016 136 6023 153
rect 6036 116 6043 233
rect 6156 167 6163 363
rect 6236 347 6243 1636
rect 6276 1623 6283 2393
rect 6296 2267 6303 2533
rect 6256 1616 6283 1623
rect 6276 1303 6283 1583
rect 6256 1296 6283 1303
rect 6296 1163 6303 1303
rect 6276 1156 6303 1163
rect 6276 907 6283 1156
rect 6296 1107 6303 1133
rect 6256 843 6263 853
rect 6256 836 6283 843
rect 6316 836 6323 3253
rect 6356 3036 6363 3233
rect 6376 3227 6383 3473
rect 6396 3067 6403 5513
rect 6416 4447 6423 5533
rect 6456 5443 6463 5643
rect 6436 5436 6463 5443
rect 6436 5167 6443 5436
rect 6476 5207 6483 5593
rect 6496 5407 6503 5733
rect 6536 5607 6543 5913
rect 6556 5667 6563 6133
rect 6576 5527 6583 5993
rect 6616 5627 6623 5653
rect 6616 5527 6623 5613
rect 6636 5607 6643 6276
rect 6676 6247 6683 6273
rect 6696 6147 6703 6293
rect 6676 6136 6693 6143
rect 6656 5987 6663 6093
rect 6676 5767 6683 6136
rect 6736 6127 6743 6233
rect 6696 5747 6703 5953
rect 6756 5916 6763 6253
rect 6776 5947 6783 6353
rect 6796 6283 6803 6533
rect 6876 6376 6903 6383
rect 6796 6276 6823 6283
rect 6796 5916 6803 5933
rect 6716 5747 6723 5773
rect 6696 5663 6703 5733
rect 6676 5656 6703 5663
rect 6676 5636 6683 5656
rect 6696 5507 6703 5623
rect 6716 5607 6723 5643
rect 6636 5456 6643 5493
rect 6736 5387 6743 5773
rect 6776 5627 6783 5753
rect 6796 5647 6803 5813
rect 6756 5416 6763 5613
rect 6816 5567 6823 6276
rect 6876 6247 6883 6376
rect 6916 6307 6923 6473
rect 6916 6116 6923 6293
rect 6936 6147 6943 6363
rect 6956 6347 6963 6556
rect 6956 6187 6963 6333
rect 6856 6027 6863 6093
rect 6936 6047 6943 6103
rect 6456 5127 6463 5143
rect 6456 5007 6463 5113
rect 6496 5107 6503 5143
rect 6516 5107 6523 5163
rect 6536 4987 6543 5273
rect 6456 4676 6463 4973
rect 6516 4956 6543 4963
rect 6536 4907 6543 4956
rect 6696 4936 6703 5193
rect 6776 5143 6783 5393
rect 6796 5387 6803 5403
rect 6756 5136 6783 5143
rect 6436 4607 6443 4663
rect 6476 4647 6483 4663
rect 6436 4127 6443 4593
rect 6456 4107 6463 4613
rect 6516 4287 6523 4653
rect 6536 4627 6543 4893
rect 6576 4467 6583 4493
rect 6596 4476 6603 4933
rect 6736 4923 6743 4933
rect 6656 4607 6663 4713
rect 6636 4476 6643 4493
rect 6616 4427 6623 4463
rect 6416 4016 6423 4033
rect 6436 3727 6443 3983
rect 6436 3203 6443 3573
rect 6456 3247 6463 4093
rect 6476 3427 6483 4213
rect 6556 4196 6563 4273
rect 6596 4183 6603 4213
rect 6616 4187 6623 4273
rect 6676 4227 6683 4923
rect 6716 4916 6743 4923
rect 6796 4747 6803 5373
rect 6816 5167 6823 5333
rect 6836 5207 6843 5513
rect 6856 5107 6863 6013
rect 6736 4696 6743 4713
rect 6876 4667 6883 5933
rect 6896 5487 6903 5933
rect 6976 5787 6983 6533
rect 6996 6427 7003 6583
rect 7016 6563 7023 6833
rect 7016 6556 7043 6563
rect 6996 6367 7003 6373
rect 6996 6127 7003 6353
rect 7016 5967 7023 6513
rect 7036 6167 7043 6556
rect 7056 6267 7063 6753
rect 7056 6107 7063 6193
rect 7016 5867 7023 5903
rect 7056 5867 7063 5903
rect 7036 5807 7043 5853
rect 6956 5656 6963 5773
rect 6976 5663 6983 5753
rect 6976 5656 7003 5663
rect 6936 5607 6943 5643
rect 6896 5127 6903 5473
rect 6956 5407 6963 5553
rect 6976 5387 6983 5656
rect 7016 5567 7023 5773
rect 7036 5627 7043 5643
rect 7056 5436 7063 5833
rect 7076 5787 7083 7453
rect 7096 6547 7103 7613
rect 7116 7227 7123 7996
rect 7196 7887 7203 8493
rect 7216 8027 7223 8813
rect 7256 8807 7263 8973
rect 7336 8947 7343 8983
rect 7376 8823 7383 8983
rect 7416 8967 7423 8983
rect 7376 8816 7403 8823
rect 7216 7803 7223 7853
rect 7196 7796 7223 7803
rect 7236 7747 7243 8573
rect 7256 8443 7263 8793
rect 7276 8776 7303 8783
rect 7296 8647 7303 8776
rect 7276 8467 7283 8613
rect 7256 8436 7283 8443
rect 7256 7947 7263 8033
rect 7156 7587 7163 7733
rect 7256 7723 7263 7813
rect 7236 7716 7263 7723
rect 7156 7563 7163 7573
rect 7136 7556 7163 7563
rect 7136 7487 7143 7533
rect 7136 7347 7143 7473
rect 7156 7207 7163 7533
rect 7176 7067 7183 7513
rect 7196 7356 7203 7673
rect 7236 7356 7243 7716
rect 7256 7527 7263 7593
rect 7276 7507 7283 8436
rect 7296 7627 7303 8353
rect 7316 8327 7323 8533
rect 7316 8047 7323 8313
rect 7336 8207 7343 8513
rect 7396 8507 7403 8523
rect 7456 8483 7463 8503
rect 7436 8476 7463 8483
rect 7356 8296 7363 8333
rect 7376 8316 7383 8333
rect 7436 8323 7443 8476
rect 7416 8316 7443 8323
rect 7396 8167 7403 8303
rect 7356 8036 7363 8153
rect 7276 7356 7283 7373
rect 7316 7367 7323 7873
rect 7336 7787 7343 8003
rect 7216 7187 7223 7343
rect 7256 7247 7263 7343
rect 7296 7327 7303 7353
rect 7216 7007 7223 7173
rect 7256 7096 7263 7193
rect 7296 7096 7303 7113
rect 7276 7047 7283 7083
rect 7236 6896 7263 6903
rect 7256 6807 7263 6896
rect 7196 6547 7203 6713
rect 7256 6547 7263 6563
rect 7096 6327 7103 6413
rect 7116 5903 7123 6213
rect 7096 5896 7123 5903
rect 6996 5347 7003 5423
rect 7036 5407 7043 5423
rect 6536 3987 6543 4183
rect 6576 4176 6603 4183
rect 6616 3996 6623 4173
rect 6496 3227 6503 3513
rect 6436 3196 6463 3203
rect 6336 2747 6343 2763
rect 6336 1787 6343 2633
rect 6356 2587 6363 2743
rect 6396 2587 6403 2743
rect 6416 2727 6423 3053
rect 6356 2527 6363 2553
rect 6396 2527 6403 2573
rect 6356 2276 6383 2283
rect 6336 1287 6343 1773
rect 6356 1167 6363 2276
rect 6416 2107 6423 2573
rect 6436 2247 6443 3053
rect 6396 1803 6403 2033
rect 6416 1987 6423 2063
rect 6456 1827 6463 3053
rect 6496 2536 6503 2573
rect 6516 2567 6523 3853
rect 6536 3683 6543 3953
rect 6556 3736 6583 3743
rect 6556 3707 6563 3736
rect 6596 3707 6603 3723
rect 6656 3707 6663 3753
rect 6676 3747 6683 4013
rect 6536 3676 6563 3683
rect 6556 3536 6563 3676
rect 6576 3516 6583 3533
rect 6476 2507 6483 2523
rect 6496 2076 6503 2333
rect 6536 2087 6543 3233
rect 6556 2307 6563 3253
rect 6576 3036 6583 3413
rect 6676 3236 6683 3713
rect 6696 3687 6703 3993
rect 6596 3007 6603 3023
rect 6656 2807 6663 3033
rect 6616 2756 6623 2793
rect 6656 2756 6663 2773
rect 6696 2587 6703 3673
rect 6716 3287 6723 3973
rect 6736 3267 6743 4653
rect 6856 4496 6863 4593
rect 6816 4476 6843 4483
rect 6876 4476 6883 4553
rect 6776 4196 6783 4353
rect 6756 4156 6773 4163
rect 6756 3703 6763 4053
rect 6776 3727 6783 4153
rect 6756 3696 6783 3703
rect 6756 2767 6763 3633
rect 6776 3607 6783 3696
rect 6776 3536 6783 3593
rect 6796 3547 6803 4253
rect 6816 4067 6823 4476
rect 6816 3703 6823 4013
rect 6896 3996 6903 5093
rect 6916 4923 6923 5333
rect 6976 5107 6983 5143
rect 6916 4916 6943 4923
rect 6936 4663 6943 4893
rect 6976 4707 6983 4913
rect 7016 4667 7023 5133
rect 7036 5007 7043 5153
rect 7076 4927 7083 5453
rect 6936 4656 6963 4663
rect 6936 4027 6943 4656
rect 6976 4447 6983 4643
rect 7036 4427 7043 4693
rect 7096 4476 7103 5013
rect 6996 4167 7003 4183
rect 7036 4127 7043 4183
rect 6856 3976 6883 3983
rect 6856 3847 6863 3976
rect 6916 3947 6923 3983
rect 6816 3696 6843 3703
rect 6596 2327 6603 2373
rect 6596 2276 6603 2313
rect 6556 2263 6563 2273
rect 6636 2267 6643 2283
rect 6556 2256 6583 2263
rect 6476 1827 6483 2063
rect 6396 1796 6423 1803
rect 6496 1787 6503 1993
rect 6536 1807 6543 2073
rect 6436 1547 6443 1783
rect 6476 1547 6483 1563
rect 6416 1147 6423 1293
rect 6336 1116 6343 1133
rect 6416 1116 6423 1133
rect 6356 1027 6363 1103
rect 6396 1087 6403 1103
rect 6356 987 6363 1013
rect 6367 897 6383 904
rect 6296 787 6303 823
rect 6336 807 6343 823
rect 6376 756 6383 897
rect 6356 749 6383 756
rect 6076 87 6083 123
rect 6276 107 6283 143
rect 6356 27 6363 749
rect 6436 643 6443 1153
rect 6456 807 6463 1293
rect 6536 1287 6543 1303
rect 6596 1187 6603 2093
rect 6616 2087 6623 2263
rect 6616 1707 6623 2073
rect 6636 1767 6643 1783
rect 6636 1567 6643 1753
rect 6656 1167 6663 2573
rect 6676 2556 6703 2563
rect 6676 2527 6683 2556
rect 6756 2536 6763 2573
rect 6676 2267 6683 2513
rect 6696 2287 6703 2513
rect 6756 2076 6763 2133
rect 6696 1227 6703 1783
rect 6756 1307 6763 1773
rect 6776 1647 6783 2793
rect 6796 2547 6803 3113
rect 6816 3036 6823 3073
rect 6836 3067 6843 3593
rect 6856 3307 6863 3613
rect 6856 3036 6863 3293
rect 6896 3247 6903 3753
rect 6916 3667 6923 3933
rect 6956 3707 6963 3993
rect 6996 3536 7003 4013
rect 6876 2347 6883 3053
rect 6836 2276 6843 2293
rect 6876 2267 6883 2283
rect 6816 1343 6823 2173
rect 6856 1387 6863 2263
rect 6896 2107 6903 2553
rect 6916 2547 6923 3273
rect 6956 3207 6963 3223
rect 6936 2127 6943 3093
rect 6996 3087 7003 3223
rect 7016 2967 7023 3233
rect 6976 2576 6983 2793
rect 7036 2783 7043 3533
rect 7056 3107 7063 4433
rect 7076 4167 7083 4413
rect 7116 3867 7123 5553
rect 7136 5127 7143 6173
rect 7156 6136 7163 6213
rect 7176 6167 7183 6363
rect 7196 6136 7203 6153
rect 7176 5896 7183 5973
rect 7196 5807 7203 6013
rect 7216 5867 7223 6513
rect 7316 6327 7323 7253
rect 7336 6867 7343 7593
rect 7356 6027 7363 7553
rect 7376 7467 7383 7933
rect 7396 7827 7403 8033
rect 7436 7927 7443 8316
rect 7396 6527 7403 7793
rect 7416 7627 7423 7823
rect 7456 7607 7463 8153
rect 7416 7547 7423 7563
rect 7456 7556 7463 7593
rect 7476 7507 7483 7543
rect 7496 7507 7503 8053
rect 7516 7807 7523 8613
rect 7536 8527 7543 8673
rect 7556 8327 7563 9353
rect 7576 8787 7583 9453
rect 7596 9016 7623 9023
rect 7656 9016 7663 9033
rect 7596 8947 7603 9016
rect 7576 8507 7583 8673
rect 7596 8427 7603 8933
rect 7636 8787 7643 9003
rect 7656 8607 7663 8783
rect 7676 8627 7683 9443
rect 7836 9387 7843 9913
rect 7876 9887 7883 9913
rect 7856 9687 7863 9723
rect 7856 9467 7863 9483
rect 7716 9256 7723 9273
rect 7696 9227 7703 9243
rect 7616 8516 7623 8533
rect 7636 8467 7643 8483
rect 7576 8207 7583 8393
rect 7596 8296 7603 8373
rect 7616 8347 7623 8393
rect 7616 8276 7623 8333
rect 7636 8296 7643 8413
rect 7676 8283 7683 8333
rect 7656 8276 7683 8283
rect 7576 8027 7583 8043
rect 7616 8036 7623 8073
rect 7616 7867 7623 7973
rect 7636 7927 7643 8023
rect 7516 7527 7523 7753
rect 7416 7127 7423 7493
rect 7507 7376 7523 7383
rect 7456 7063 7463 7353
rect 7516 7247 7523 7376
rect 7456 7056 7483 7063
rect 7416 6787 7423 6863
rect 7456 6583 7463 6653
rect 7496 6627 7503 7033
rect 7516 6903 7523 7063
rect 7536 7027 7543 7083
rect 7516 6896 7543 6903
rect 7516 6647 7523 6873
rect 7536 6867 7543 6896
rect 7496 6596 7503 6613
rect 7536 6587 7543 6603
rect 7456 6576 7483 6583
rect 7356 5936 7363 5973
rect 7316 5623 7323 5793
rect 7316 5616 7343 5623
rect 7156 5447 7163 5603
rect 7296 5456 7303 5553
rect 7276 5436 7283 5453
rect 7196 5156 7203 5193
rect 7216 5127 7223 5143
rect 7136 4447 7143 4953
rect 7176 4936 7183 5113
rect 7156 4423 7163 4923
rect 7196 4887 7203 4913
rect 7216 4656 7243 4663
rect 7136 4416 7163 4423
rect 7136 4027 7143 4416
rect 7076 3747 7083 3773
rect 7136 3767 7143 3983
rect 7096 3707 7103 3723
rect 7136 3587 7143 3713
rect 7116 3527 7123 3573
rect 7056 3036 7063 3073
rect 7076 3067 7083 3493
rect 7096 3467 7103 3513
rect 7096 3047 7103 3293
rect 7016 2776 7043 2783
rect 6996 2747 7003 2773
rect 7016 2583 7023 2776
rect 7056 2687 7063 2723
rect 7016 2576 7043 2583
rect 6956 2527 6963 2543
rect 6896 2067 6903 2093
rect 6936 2047 6943 2093
rect 6956 2076 6963 2093
rect 6996 2076 7003 2133
rect 6896 1727 6903 1783
rect 6956 1596 6963 1673
rect 6996 1596 7003 1633
rect 6796 1336 6823 1343
rect 6796 1316 6803 1336
rect 6836 1316 6843 1333
rect 6767 1296 6783 1303
rect 6536 1107 6543 1133
rect 6596 1116 6603 1133
rect 6676 1116 6683 1133
rect 6556 1027 6563 1093
rect 6576 1067 6583 1113
rect 6696 1107 6703 1153
rect 6496 836 6523 843
rect 6496 807 6503 836
rect 6556 803 6563 1013
rect 6616 987 6623 1103
rect 6536 796 6563 803
rect 6396 636 6423 643
rect 6436 636 6463 643
rect 6376 -17 6383 343
rect 5356 -24 5383 -17
rect 6356 -24 6383 -17
rect 6396 -24 6403 636
rect 6636 343 6643 753
rect 6656 636 6663 673
rect 6676 623 6683 773
rect 6716 643 6723 1173
rect 6816 1167 6823 1303
rect 6856 1223 6863 1303
rect 6836 1216 6863 1223
rect 6816 1047 6823 1113
rect 6736 807 6743 823
rect 6776 787 6783 823
rect 6836 767 6843 1216
rect 6936 1116 6943 1133
rect 6876 987 6883 1103
rect 6996 867 7003 1333
rect 7016 1107 7023 2113
rect 7036 1087 7043 2576
rect 7056 1407 7063 2553
rect 7076 1767 7083 2533
rect 7116 2527 7123 2753
rect 7136 2547 7143 3033
rect 7156 2727 7163 3973
rect 7176 3587 7183 4513
rect 7196 3767 7203 4473
rect 7176 3007 7183 3573
rect 7196 3567 7203 3753
rect 7216 3607 7223 4656
rect 7236 4216 7243 4253
rect 7256 4247 7263 5353
rect 7276 5147 7283 5293
rect 7296 4476 7323 4483
rect 7276 4447 7283 4463
rect 7236 3667 7243 3733
rect 7256 3647 7263 4193
rect 7316 4107 7323 4476
rect 7336 4447 7343 5616
rect 7356 5167 7363 5773
rect 7376 5567 7383 6433
rect 7416 6396 7423 6453
rect 7456 6396 7483 6403
rect 7436 6367 7443 6383
rect 7476 6167 7483 6396
rect 7476 6103 7483 6153
rect 7496 6127 7503 6393
rect 7516 6387 7523 6583
rect 7556 6567 7563 6893
rect 7416 5987 7423 6103
rect 7456 6096 7483 6103
rect 7496 6007 7503 6113
rect 7476 5896 7503 5903
rect 7496 5767 7503 5896
rect 7516 5767 7523 5883
rect 7396 5636 7423 5643
rect 7396 5607 7403 5636
rect 7436 5587 7443 5633
rect 7436 5227 7443 5513
rect 7456 5367 7463 5653
rect 7376 4467 7383 5053
rect 7416 4976 7423 5153
rect 7436 4956 7443 5033
rect 7396 4667 7403 4693
rect 7356 3996 7363 4013
rect 7376 3987 7383 4453
rect 7336 3783 7343 3983
rect 7336 3776 7363 3783
rect 7216 3496 7223 3513
rect 7256 3496 7263 3553
rect 7276 3467 7283 3483
rect 7196 3187 7203 3223
rect 7176 2747 7183 2993
rect 7136 2276 7143 2333
rect 7176 2127 7183 2553
rect 7196 2267 7203 3173
rect 7296 3127 7303 3553
rect 7316 3227 7323 3593
rect 7356 3247 7363 3776
rect 7376 3527 7383 3913
rect 7376 3247 7383 3513
rect 7396 3256 7403 4293
rect 7436 4287 7443 4633
rect 7416 3367 7423 4213
rect 7436 3283 7443 4213
rect 7456 3947 7463 4653
rect 7476 4227 7483 5273
rect 7496 4607 7503 5713
rect 7536 5527 7543 6333
rect 7576 6087 7583 7733
rect 7596 7567 7603 7813
rect 7696 7707 7703 9093
rect 7716 8007 7723 9153
rect 7736 7747 7743 8453
rect 7756 8227 7763 9333
rect 7636 7547 7643 7593
rect 7676 7563 7683 7693
rect 7676 7556 7703 7563
rect 7516 5407 7523 5423
rect 7556 5187 7563 5993
rect 7576 5447 7583 5973
rect 7596 5647 7603 7513
rect 7656 7376 7683 7383
rect 7656 7327 7663 7376
rect 7736 7347 7743 7553
rect 7696 7336 7713 7343
rect 7616 6147 7623 6933
rect 7636 6227 7643 7133
rect 7736 7076 7743 7333
rect 7756 7043 7763 7953
rect 7736 7036 7763 7043
rect 7676 6687 7683 7033
rect 7696 6876 7703 7013
rect 7696 6416 7703 6553
rect 7736 6543 7743 7036
rect 7776 7027 7783 8873
rect 7756 6567 7763 6583
rect 7736 6536 7763 6543
rect 7716 6347 7723 6383
rect 7636 6116 7643 6153
rect 7616 5987 7623 6103
rect 7616 5907 7623 5933
rect 7656 5627 7663 6073
rect 7696 5923 7703 5953
rect 7716 5947 7723 6313
rect 7676 5916 7703 5923
rect 7676 5747 7683 5916
rect 7696 5607 7703 5873
rect 7756 5807 7763 6536
rect 7796 5863 7803 9373
rect 7876 9247 7883 9853
rect 7916 9347 7923 9916
rect 7956 9907 7963 10216
rect 7976 10167 7983 10273
rect 8156 10263 8163 10776
rect 8176 10436 8183 10453
rect 8136 10256 8163 10263
rect 7976 9867 7983 10153
rect 8016 9847 8023 10233
rect 8136 10216 8143 10256
rect 8196 10236 8203 10253
rect 8116 9956 8123 9973
rect 8096 9867 8103 9923
rect 8016 9776 8023 9833
rect 8216 9747 8223 10433
rect 8196 9736 8213 9743
rect 7956 9276 7963 9633
rect 7996 9607 8003 9733
rect 8016 9276 8023 9473
rect 7816 9016 7843 9023
rect 7876 9016 7883 9073
rect 7816 8987 7823 9016
rect 7896 8776 7903 8973
rect 7936 8763 7943 9033
rect 7916 8756 7943 8763
rect 7876 8516 7883 8533
rect 7856 8447 7863 8513
rect 7956 8503 7963 8613
rect 7936 8496 7963 8503
rect 7896 8327 7903 8483
rect 7876 8263 7883 8283
rect 7876 8256 7903 8263
rect 7816 7987 7823 8003
rect 7816 6947 7823 7513
rect 7836 6747 7843 7993
rect 7876 7867 7883 8173
rect 7896 7867 7903 8256
rect 7916 8247 7923 8283
rect 7936 8027 7943 8213
rect 7856 7207 7863 7853
rect 7896 7836 7903 7853
rect 7936 7836 7943 7913
rect 7956 7867 7963 8313
rect 7976 8267 7983 9263
rect 7996 8323 8003 9013
rect 8036 8967 8043 9263
rect 8076 9047 8083 9513
rect 8176 9047 8183 9443
rect 8036 8727 8043 8953
rect 8076 8796 8083 9033
rect 8136 9016 8163 9023
rect 8116 8796 8123 8973
rect 8156 8867 8163 9016
rect 8196 9007 8203 9653
rect 8216 9467 8223 9733
rect 8236 9647 8243 10933
rect 8356 10727 8363 10753
rect 8256 10696 8283 10703
rect 8276 10567 8283 10696
rect 8296 10507 8303 10683
rect 8316 10467 8323 10693
rect 8216 9276 8223 9293
rect 8236 9087 8243 9263
rect 8256 8987 8263 9833
rect 8296 9743 8303 9753
rect 8276 9736 8303 9743
rect 8276 9276 8283 9493
rect 8276 8987 8283 9033
rect 8156 8796 8183 8803
rect 8096 8763 8103 8783
rect 8176 8767 8183 8796
rect 8087 8756 8103 8763
rect 7996 8316 8023 8323
rect 7876 7816 7883 7833
rect 7916 7807 7923 7823
rect 7916 7547 7923 7563
rect 7976 7527 7983 7543
rect 7876 7427 7883 7473
rect 7916 7356 7923 7393
rect 7956 7367 7963 7493
rect 7887 7336 7903 7343
rect 7976 7327 7983 7513
rect 7816 6527 7823 6593
rect 7816 6507 7823 6513
rect 7776 5856 7803 5863
rect 7576 5247 7583 5433
rect 7536 4496 7543 4913
rect 7576 4687 7583 5233
rect 7516 4476 7523 4493
rect 7476 4027 7483 4183
rect 7516 4107 7523 4183
rect 7536 4167 7543 4453
rect 7576 4147 7583 4553
rect 7596 4283 7603 5473
rect 7736 5416 7743 5793
rect 7776 5687 7783 5856
rect 7616 4387 7623 5353
rect 7636 4936 7643 5213
rect 7696 5176 7703 5393
rect 7676 5067 7683 5163
rect 7656 4916 7663 5013
rect 7636 4647 7643 4853
rect 7696 4703 7703 4923
rect 7696 4696 7723 4703
rect 7656 4487 7663 4663
rect 7696 4627 7703 4663
rect 7596 4276 7623 4283
rect 7456 3487 7463 3793
rect 7476 3483 7483 3973
rect 7516 3967 7523 4013
rect 7547 3996 7563 4003
rect 7596 3996 7603 4033
rect 7516 3687 7523 3853
rect 7536 3807 7543 3993
rect 7576 3967 7583 3983
rect 7616 3976 7623 4276
rect 7636 3987 7643 4253
rect 7656 3967 7663 4413
rect 7516 3496 7523 3573
rect 7476 3476 7503 3483
rect 7436 3276 7463 3283
rect 7376 3036 7383 3073
rect 7296 3016 7323 3023
rect 7296 3003 7303 3016
rect 7276 2996 7303 3003
rect 7276 2767 7283 2996
rect 7356 2967 7363 3023
rect 7316 2756 7343 2763
rect 7216 2556 7223 2613
rect 7276 2536 7303 2543
rect 7296 2287 7303 2536
rect 7316 2147 7323 2756
rect 7356 2727 7363 2743
rect 7396 2276 7403 2353
rect 7416 2327 7423 3243
rect 7416 2247 7423 2263
rect 7216 2096 7223 2113
rect 7256 2063 7263 2113
rect 7456 2087 7463 3276
rect 7476 3267 7483 3476
rect 7556 3347 7563 3393
rect 7576 3187 7583 3953
rect 7536 3027 7543 3153
rect 7576 3036 7583 3093
rect 7556 3016 7563 3033
rect 7636 2867 7643 3953
rect 7676 3607 7683 4473
rect 7696 4287 7703 4613
rect 7716 4327 7723 4696
rect 7736 4647 7743 4933
rect 7756 4887 7763 4953
rect 7736 4507 7743 4633
rect 7756 4527 7763 4673
rect 7776 4487 7783 5193
rect 7796 4767 7803 5733
rect 7816 5207 7823 6353
rect 7836 5947 7843 6633
rect 7856 6347 7863 7033
rect 7896 6587 7903 7113
rect 7936 7076 7943 7313
rect 7916 6967 7923 7043
rect 7936 6876 7943 6893
rect 7996 6887 8003 8253
rect 7956 6827 7963 6863
rect 8016 6767 8023 8316
rect 8036 7667 8043 8593
rect 8076 8307 8083 8753
rect 8176 8587 8183 8753
rect 8096 8307 8103 8573
rect 8156 8507 8163 8523
rect 8116 8316 8123 8333
rect 8196 8316 8203 8353
rect 8216 8307 8223 8373
rect 8096 8036 8103 8073
rect 8076 8007 8083 8023
rect 7976 6596 7983 6613
rect 7956 6416 7963 6553
rect 7996 6407 8003 6583
rect 8016 6567 8023 6603
rect 8036 6543 8043 7313
rect 8076 7287 8083 7853
rect 8136 7816 8143 8113
rect 8156 7836 8163 7873
rect 8196 7847 8203 8013
rect 8096 7327 8103 7813
rect 8016 6536 8043 6543
rect 7896 6396 7923 6403
rect 7896 6367 7903 6396
rect 7976 6247 7983 6373
rect 7856 6067 7863 6113
rect 7836 5887 7843 5913
rect 7836 5507 7843 5873
rect 7856 5727 7863 6053
rect 7876 6047 7883 6123
rect 7936 6083 7943 6103
rect 7916 6076 7943 6083
rect 7916 5827 7923 6076
rect 7936 6067 7943 6076
rect 7956 5936 7963 6073
rect 7936 5867 7943 5903
rect 7916 5636 7923 5653
rect 7896 5527 7903 5603
rect 7836 5183 7843 5433
rect 7876 5427 7883 5453
rect 7816 5176 7843 5183
rect 7796 4667 7803 4733
rect 7816 4707 7823 5176
rect 7856 5107 7863 5173
rect 7856 4927 7863 5093
rect 7876 4903 7883 5413
rect 7896 5387 7903 5493
rect 7936 5487 7943 5833
rect 7936 5416 7943 5473
rect 7956 5436 7963 5613
rect 7996 5547 8003 6233
rect 8016 5927 8023 6536
rect 8036 6063 8043 6153
rect 8056 6087 8063 6873
rect 8076 6867 8083 7273
rect 8096 6427 8103 6893
rect 8116 6807 8123 7793
rect 8136 7387 8143 7653
rect 8216 7567 8223 8033
rect 8236 7987 8243 8633
rect 8256 7827 8263 8513
rect 8276 8487 8283 8973
rect 8316 8187 8323 10453
rect 8356 10447 8363 10713
rect 8456 10707 8463 11153
rect 8476 11147 8483 11196
rect 8856 11196 8883 11203
rect 8916 11196 8933 11203
rect 8696 11167 8703 11183
rect 8576 10847 8583 11093
rect 8636 10916 8643 11113
rect 8616 10847 8623 10883
rect 8516 10716 8523 10733
rect 8476 10696 8503 10703
rect 8476 10603 8483 10696
rect 8476 10596 8503 10603
rect 8416 10456 8443 10463
rect 8396 10427 8403 10443
rect 8336 9956 8343 10213
rect 8436 10207 8443 10456
rect 8456 10436 8483 10443
rect 8356 10187 8363 10203
rect 8456 10187 8463 10436
rect 8496 10427 8503 10596
rect 8576 10327 8583 10833
rect 8696 10687 8703 11153
rect 8856 11147 8863 11196
rect 8896 11147 8903 11183
rect 8956 11147 8963 11213
rect 9196 11196 9223 11203
rect 8856 10916 8863 11133
rect 8816 10883 8823 10913
rect 8816 10876 8843 10883
rect 8756 10687 8763 10703
rect 8836 10687 8843 10876
rect 8976 10707 8983 11193
rect 8996 10727 9003 11173
rect 9136 11147 9143 11193
rect 9216 11167 9223 11196
rect 9616 11187 9623 11193
rect 10056 11176 10083 11183
rect 10116 11176 10123 11193
rect 9616 11163 9623 11173
rect 9696 11163 9703 11173
rect 9376 10916 9383 11163
rect 9416 11147 9423 11163
rect 9616 11156 9643 11163
rect 9676 11156 9703 11163
rect 9076 10747 9083 10903
rect 9076 10703 9083 10733
rect 8736 10347 8743 10403
rect 8636 10236 8643 10333
rect 8576 10207 8583 10233
rect 8576 9983 8583 10193
rect 8527 9976 8543 9983
rect 8576 9976 8603 9983
rect 8356 9767 8363 9923
rect 8416 9747 8423 9893
rect 8336 9707 8343 9743
rect 8376 9247 8383 9443
rect 8396 9427 8403 9463
rect 8396 9267 8403 9413
rect 8416 9187 8423 9273
rect 8356 8967 8363 9003
rect 8356 8947 8363 8953
rect 8376 8947 8383 9023
rect 8396 8987 8403 9003
rect 8416 8947 8423 9173
rect 8436 8927 8443 9973
rect 8456 9707 8463 9973
rect 8596 9947 8603 9976
rect 8356 8827 8363 8873
rect 8396 8796 8403 8853
rect 8456 8807 8463 9293
rect 8496 9247 8503 9263
rect 8536 9256 8543 9333
rect 8576 9247 8583 9463
rect 8576 9107 8583 9233
rect 8476 8787 8483 9093
rect 8516 8987 8523 9013
rect 8356 8287 8363 8773
rect 8456 8523 8463 8613
rect 8436 8516 8463 8523
rect 8276 8043 8283 8093
rect 8276 8036 8303 8043
rect 8376 8023 8383 8493
rect 8396 8316 8403 8333
rect 8436 8316 8443 8453
rect 8476 8316 8483 8573
rect 8316 8007 8323 8023
rect 8356 8016 8383 8023
rect 8356 7927 8363 8016
rect 8156 7507 8163 7533
rect 8176 7487 8183 7563
rect 8196 7467 8203 7543
rect 8236 7387 8243 7533
rect 8136 7147 8143 7373
rect 8236 7367 8243 7373
rect 8256 7347 8263 7613
rect 8276 7547 8283 7833
rect 8296 7523 8303 7553
rect 8276 7516 8303 7523
rect 8156 7127 8163 7343
rect 8136 6867 8143 6993
rect 8176 6876 8183 7133
rect 8216 6876 8223 7053
rect 8256 6883 8263 7233
rect 8276 7087 8283 7516
rect 8316 7443 8323 7573
rect 8356 7527 8363 7913
rect 8436 7827 8443 8273
rect 8436 7647 8443 7813
rect 8416 7576 8423 7613
rect 8296 7436 8323 7443
rect 8296 7336 8303 7436
rect 8256 6876 8283 6883
rect 8076 6107 8083 6133
rect 8096 6127 8103 6413
rect 8136 6247 8143 6833
rect 8196 6727 8203 6853
rect 8236 6847 8243 6863
rect 8236 6596 8243 6793
rect 8196 6556 8223 6563
rect 8156 6396 8163 6553
rect 8196 6387 8203 6556
rect 8176 6147 8183 6363
rect 8156 6116 8163 6133
rect 8176 6087 8183 6103
rect 8036 6056 8063 6063
rect 8016 5407 8023 5653
rect 7896 5083 7903 5373
rect 7916 5107 7923 5163
rect 7896 5076 7923 5083
rect 7916 4936 7923 5076
rect 7856 4896 7883 4903
rect 7796 4456 7823 4463
rect 7816 4407 7823 4456
rect 7696 4207 7703 4233
rect 7696 3407 7703 3993
rect 7716 3627 7723 4173
rect 7736 3967 7743 4073
rect 7756 3967 7763 4273
rect 7776 3927 7783 4393
rect 7756 3716 7763 3753
rect 7796 3716 7803 3933
rect 7736 3687 7743 3693
rect 7816 3687 7823 4193
rect 7836 4007 7843 4473
rect 7856 4427 7863 4896
rect 7936 4727 7943 4913
rect 7976 4763 7983 5143
rect 7976 4756 8003 4763
rect 7876 4663 7883 4693
rect 7916 4676 7923 4693
rect 7876 4656 7903 4663
rect 7936 4656 7963 4663
rect 7896 4183 7903 4613
rect 7936 4207 7943 4513
rect 7956 4496 7963 4656
rect 7976 4527 7983 4713
rect 7956 4427 7963 4453
rect 7976 4447 7983 4453
rect 7996 4327 8003 4756
rect 8016 4707 8023 5373
rect 8036 4707 8043 5693
rect 8056 5387 8063 6056
rect 8136 6047 8143 6083
rect 8076 5687 8083 5713
rect 8156 5707 8163 5903
rect 8096 5656 8103 5673
rect 8136 5656 8163 5663
rect 8116 5607 8123 5643
rect 8056 4927 8063 5153
rect 8016 4647 8023 4693
rect 8016 4447 8023 4473
rect 8036 4367 8043 4673
rect 7896 4176 7923 4183
rect 7896 4167 7903 4176
rect 7956 4167 7963 4183
rect 7876 3956 7883 4033
rect 7956 4007 7963 4153
rect 7896 3976 7903 3993
rect 7696 3367 7703 3373
rect 7696 3256 7703 3353
rect 7716 3067 7723 3593
rect 7736 3567 7743 3593
rect 7756 3536 7763 3653
rect 7736 3516 7743 3533
rect 7836 3527 7843 3893
rect 7916 3787 7923 3973
rect 7756 3283 7763 3493
rect 7736 3276 7763 3283
rect 7496 2536 7503 2753
rect 7476 2507 7483 2523
rect 7476 2287 7483 2493
rect 7236 2056 7263 2063
rect 7136 1796 7143 1853
rect 7156 1687 7163 1783
rect 7156 1547 7163 1613
rect 7076 1267 7083 1323
rect 7096 1267 7103 1343
rect 7176 1327 7183 1803
rect 7196 1596 7203 1613
rect 7276 1567 7283 1673
rect 7296 1336 7303 1773
rect 7336 1336 7343 1873
rect 7356 1367 7363 2073
rect 7396 2043 7403 2073
rect 7396 2036 7423 2043
rect 7376 1767 7383 1783
rect 7416 1747 7423 1783
rect 7556 1767 7563 1813
rect 7576 1787 7583 2743
rect 7616 2507 7623 2743
rect 7656 2527 7663 3053
rect 7736 2767 7743 3276
rect 7756 3027 7763 3253
rect 7696 2563 7703 2633
rect 7696 2556 7723 2563
rect 7736 2556 7743 2733
rect 7596 2267 7603 2283
rect 7636 2276 7643 2513
rect 7716 2367 7723 2556
rect 7616 2167 7623 2263
rect 7576 1607 7583 1773
rect 7496 1303 7503 1393
rect 7556 1347 7563 1373
rect 7496 1296 7523 1303
rect 6956 787 6963 823
rect 6716 636 6743 643
rect 6676 616 6703 623
rect 6736 347 6743 636
rect 6756 387 6763 623
rect 6976 407 6983 803
rect 6996 687 7003 823
rect 7036 647 7043 853
rect 7056 667 7063 1153
rect 7116 1116 7123 1193
rect 6996 347 7003 623
rect 7116 587 7123 893
rect 7136 867 7143 1133
rect 7176 1116 7183 1133
rect 7156 1067 7163 1083
rect 7156 807 7163 833
rect 7176 827 7183 843
rect 7196 747 7203 863
rect 7236 856 7263 863
rect 7256 767 7263 856
rect 7336 707 7343 1213
rect 7376 1096 7383 1233
rect 7356 1007 7363 1073
rect 7356 867 7363 913
rect 7376 847 7383 933
rect 7396 787 7403 873
rect 7416 827 7423 953
rect 7436 927 7443 1083
rect 7456 1047 7463 1093
rect 7256 656 7263 693
rect 7276 636 7283 653
rect 7316 363 7323 693
rect 7476 636 7483 653
rect 7536 647 7543 913
rect 7556 856 7563 893
rect 7576 847 7583 1303
rect 7596 1147 7603 2053
rect 7616 1816 7623 2093
rect 7676 2076 7683 2193
rect 7716 2083 7723 2293
rect 7696 2076 7723 2083
rect 7636 1607 7643 1803
rect 7696 1727 7703 2076
rect 7716 1616 7723 1633
rect 7676 1147 7683 1553
rect 7756 1323 7763 2153
rect 7776 1387 7783 3393
rect 7816 3227 7823 3253
rect 7816 3056 7823 3073
rect 7796 3007 7803 3023
rect 7796 2247 7803 2973
rect 7816 2756 7823 3013
rect 7836 2987 7843 3513
rect 7836 2647 7843 2723
rect 7856 2307 7863 3733
rect 7916 3283 7923 3553
rect 7976 3527 7983 4193
rect 7996 3887 8003 4073
rect 8036 3767 8043 3993
rect 8056 3747 8063 4713
rect 8076 4007 8083 4693
rect 8096 4007 8103 5413
rect 8116 5227 8123 5593
rect 8156 5527 8163 5656
rect 8176 5436 8183 5913
rect 8196 5403 8203 6213
rect 8216 6087 8223 6133
rect 8176 5396 8203 5403
rect 8176 5176 8183 5396
rect 8256 5267 8263 6713
rect 8276 6027 8283 6876
rect 8296 6607 8303 7213
rect 8316 7187 8323 7436
rect 8476 7376 8483 7473
rect 8296 6067 8303 6593
rect 8336 6347 8343 7193
rect 8416 7096 8423 7193
rect 8376 6367 8383 6813
rect 8416 6583 8423 7013
rect 8436 6896 8463 6903
rect 8436 6787 8443 6896
rect 8496 6623 8503 8653
rect 8516 8507 8523 8933
rect 8536 8547 8543 9073
rect 8636 9047 8643 9633
rect 8636 8996 8643 9033
rect 8556 8947 8563 8993
rect 8556 8767 8563 8933
rect 8656 8867 8663 8983
rect 8576 8307 8583 8813
rect 8596 8767 8603 8853
rect 8636 8816 8643 8853
rect 8596 8707 8603 8753
rect 8656 8667 8663 8853
rect 8596 8367 8603 8653
rect 8656 8516 8663 8533
rect 8636 8407 8643 8483
rect 8556 8036 8563 8293
rect 8576 7827 8583 8233
rect 8596 8087 8603 8353
rect 8676 8316 8683 9453
rect 8696 8747 8703 10313
rect 8756 9943 8763 10673
rect 8896 10456 8903 10493
rect 8816 9956 8823 10013
rect 8756 9936 8783 9943
rect 8716 9736 8743 9743
rect 8736 9607 8743 9736
rect 8756 9687 8763 9723
rect 8776 9447 8783 9936
rect 8796 9787 8803 9943
rect 8816 9507 8823 9733
rect 8876 9667 8883 10253
rect 8816 9476 8823 9493
rect 8796 9447 8803 9463
rect 8796 9427 8803 9433
rect 8736 9276 8763 9283
rect 8796 9276 8803 9393
rect 8836 9287 8843 9333
rect 8736 8987 8743 9276
rect 8816 9167 8823 9263
rect 8716 8316 8723 8353
rect 8636 8296 8663 8303
rect 8636 8263 8643 8296
rect 8636 8256 8663 8263
rect 8596 7836 8603 8073
rect 8516 7527 8523 7573
rect 8516 7107 8523 7153
rect 8536 6827 8543 7233
rect 8556 6927 8563 7213
rect 8576 6847 8583 7793
rect 8596 7336 8603 7673
rect 8616 7227 8623 7813
rect 8636 7407 8643 8173
rect 8656 7807 8663 8256
rect 8756 8247 8763 8793
rect 8776 8547 8783 9153
rect 8856 9067 8863 9483
rect 8896 9407 8903 10033
rect 8916 9347 8923 10373
rect 8936 9947 8943 10693
rect 9016 10687 9023 10703
rect 9056 10696 9083 10703
rect 8956 10447 8963 10553
rect 9016 10147 9023 10673
rect 9056 10203 9063 10696
rect 9136 10467 9143 10873
rect 9156 10707 9163 10903
rect 9176 10887 9183 10913
rect 9176 10716 9203 10723
rect 9236 10716 9243 10853
rect 9096 10407 9103 10423
rect 9156 10387 9163 10443
rect 9176 10407 9183 10716
rect 9216 10447 9223 10703
rect 9316 10687 9323 10703
rect 9336 10663 9343 10913
rect 9396 10907 9403 11113
rect 9616 10916 9643 10923
rect 9616 10907 9623 10916
rect 9356 10867 9363 10903
rect 9396 10696 9403 10753
rect 9416 10707 9423 10893
rect 9576 10736 9603 10743
rect 9316 10656 9343 10663
rect 9096 10216 9103 10253
rect 9116 10207 9123 10373
rect 9287 10236 9303 10243
rect 9136 10216 9163 10223
rect 9056 10196 9083 10203
rect 8936 9776 8963 9783
rect 8936 9527 8943 9776
rect 8996 9487 9003 9953
rect 9016 9847 9023 9943
rect 9076 9927 9083 9963
rect 9096 9947 9103 10133
rect 9156 9927 9163 10216
rect 8816 8887 8823 9053
rect 8836 9016 8863 9023
rect 8896 9016 8923 9023
rect 8836 8796 8843 9016
rect 8916 8987 8923 9016
rect 8856 8776 8863 8793
rect 8896 8787 8903 8933
rect 8896 8707 8903 8773
rect 8836 8387 8843 8483
rect 8736 8056 8763 8063
rect 8796 8056 8803 8073
rect 8736 8047 8743 8056
rect 8736 7807 8743 8033
rect 8676 7556 8683 7653
rect 8656 7527 8663 7543
rect 8696 7487 8703 7543
rect 8636 7247 8643 7323
rect 8656 7096 8683 7103
rect 8636 7067 8643 7083
rect 8676 7047 8683 7096
rect 8496 6616 8523 6623
rect 8416 6576 8443 6583
rect 8516 6467 8523 6616
rect 8416 6376 8423 6393
rect 8396 6347 8403 6363
rect 8276 5467 8283 5933
rect 8156 4976 8163 5113
rect 8196 5087 8203 5163
rect 8236 5067 8243 5163
rect 8116 4956 8143 4963
rect 8116 4867 8123 4956
rect 8156 4696 8183 4703
rect 8116 4167 8123 4693
rect 8156 4667 8163 4696
rect 8276 4647 8283 5073
rect 8156 4427 8163 4473
rect 8196 4456 8203 4473
rect 8216 4436 8223 4513
rect 8136 4207 8143 4373
rect 8076 3867 8083 3973
rect 8136 3956 8143 4013
rect 8156 3976 8163 4013
rect 7996 3707 8003 3723
rect 8056 3667 8063 3703
rect 7936 3487 7943 3513
rect 7947 3476 7963 3483
rect 7916 3276 7943 3283
rect 7876 3207 7883 3223
rect 7876 3047 7883 3193
rect 7896 3087 7903 3203
rect 7876 2747 7883 3033
rect 7856 2227 7863 2263
rect 7896 2207 7903 2533
rect 7916 2163 7923 3093
rect 7936 2187 7943 3276
rect 7956 3227 7963 3273
rect 7956 2647 7963 3033
rect 7956 2547 7963 2593
rect 7976 2587 7983 3293
rect 7996 3036 8003 3073
rect 8056 3067 8063 3653
rect 8016 2747 8023 2763
rect 8056 2756 8063 3033
rect 8076 2787 8083 3753
rect 8096 3627 8103 3713
rect 8116 3687 8123 3733
rect 8096 3307 8103 3613
rect 8176 3363 8183 4393
rect 8196 4216 8203 4313
rect 8236 4216 8243 4293
rect 8216 4187 8223 4203
rect 8216 3567 8223 4173
rect 8256 3967 8263 4633
rect 8296 3963 8303 5453
rect 8316 4807 8323 6053
rect 8336 5327 8343 6113
rect 8396 6047 8403 6333
rect 8416 6116 8423 6333
rect 8356 5916 8363 5953
rect 8396 5916 8403 6013
rect 8436 5907 8443 6173
rect 8376 5887 8383 5903
rect 8356 5636 8363 5713
rect 8376 5607 8383 5873
rect 8436 5687 8443 5713
rect 8316 4267 8323 4593
rect 8316 3996 8323 4193
rect 8336 4107 8343 5253
rect 8356 4227 8363 5033
rect 8376 4956 8383 5233
rect 8436 5167 8443 5673
rect 8456 5287 8463 6393
rect 8536 6347 8543 6813
rect 8476 5447 8483 5913
rect 8496 5647 8503 5773
rect 8496 5163 8503 5513
rect 8476 5156 8503 5163
rect 8416 5107 8423 5143
rect 8396 4987 8403 5073
rect 8396 4167 8403 4943
rect 8436 4936 8443 4953
rect 8476 4627 8483 5156
rect 8436 4456 8443 4493
rect 8416 4367 8423 4443
rect 8456 4436 8463 4473
rect 8476 4456 8483 4513
rect 8496 4167 8503 5133
rect 8516 4947 8523 5153
rect 8536 4687 8543 6113
rect 8556 5367 8563 6833
rect 8576 5567 8583 6413
rect 8596 6027 8603 6913
rect 8696 6856 8703 7353
rect 8756 6967 8763 7973
rect 8776 7827 8783 8043
rect 8836 7803 8843 7893
rect 8856 7836 8863 7853
rect 8816 7796 8843 7803
rect 8716 6747 8723 6843
rect 8676 6616 8683 6733
rect 8696 6387 8703 6593
rect 8716 6567 8723 6623
rect 8756 6607 8763 6913
rect 8616 6187 8623 6273
rect 8696 6207 8703 6373
rect 8616 6123 8623 6173
rect 8616 6116 8643 6123
rect 8696 6087 8703 6103
rect 8636 5936 8643 6033
rect 8656 5916 8663 5933
rect 8636 5547 8643 5893
rect 8716 5827 8723 6553
rect 8736 5707 8743 6593
rect 8696 5656 8723 5663
rect 8596 5436 8623 5443
rect 8556 4967 8563 5153
rect 8596 5107 8603 5436
rect 8636 5163 8643 5533
rect 8696 5527 8703 5656
rect 8736 5547 8743 5643
rect 8636 5156 8663 5163
rect 8676 5147 8683 5183
rect 8516 4447 8523 4653
rect 8556 4287 8563 4953
rect 8576 4507 8583 5033
rect 8596 5003 8603 5093
rect 8596 4996 8623 5003
rect 8616 4956 8623 4996
rect 8656 4956 8663 5013
rect 8676 4967 8683 5133
rect 8696 5127 8703 5163
rect 8636 4903 8643 4933
rect 8616 4896 8643 4903
rect 8356 3996 8383 4003
rect 8296 3956 8323 3963
rect 8196 3407 8203 3483
rect 8196 3387 8203 3393
rect 8176 3356 8203 3363
rect 8016 2556 8023 2713
rect 7896 2156 7923 2163
rect 7896 1847 7903 2156
rect 7936 2096 7943 2133
rect 8036 2127 8043 2743
rect 8076 2627 8083 2743
rect 8096 2347 8103 3233
rect 8116 3167 8123 3223
rect 8176 3207 8183 3243
rect 7916 1807 7923 2063
rect 7836 1767 7843 1783
rect 7756 1316 7783 1323
rect 7776 1147 7783 1316
rect 7636 1116 7643 1133
rect 7676 1116 7683 1133
rect 7756 1007 7763 1133
rect 7856 943 7863 1763
rect 7936 1596 7963 1603
rect 7956 1567 7963 1596
rect 7876 1116 7883 1133
rect 7856 936 7883 943
rect 7596 827 7603 843
rect 7716 767 7723 803
rect 7736 656 7743 693
rect 7396 376 7423 383
rect 7316 356 7343 363
rect 6616 336 6643 343
rect 6516 176 6523 213
rect 6596 207 6603 323
rect 6496 156 6503 173
rect 6536 156 6563 163
rect 6556 127 6563 156
rect 6736 136 6743 253
rect 6756 116 6763 153
rect 6876 127 6883 323
rect 6996 176 7003 273
rect 7136 167 7143 323
rect 7156 307 7163 343
rect 7196 136 7203 153
rect 7376 127 7383 363
rect 7416 327 7423 376
rect 7536 187 7543 633
rect 7876 587 7883 936
rect 7896 927 7903 1373
rect 7936 1116 7943 1333
rect 7916 1087 7923 1103
rect 7976 943 7983 1103
rect 7996 1087 8003 1813
rect 7956 936 7983 943
rect 7896 727 7903 843
rect 7936 656 7943 913
rect 7636 376 7643 393
rect 7916 387 7923 623
rect 7616 267 7623 343
rect 7876 343 7883 373
rect 7956 347 7963 936
rect 7976 836 7983 913
rect 7996 827 8003 1073
rect 8016 347 8023 1853
rect 8036 967 8043 2073
rect 8076 1767 8083 2243
rect 8096 2207 8103 2263
rect 8096 2067 8103 2193
rect 8116 1867 8123 2773
rect 8136 2087 8143 3053
rect 8196 2847 8203 3356
rect 8256 3047 8263 3633
rect 8296 3047 8303 3153
rect 8316 3067 8323 3956
rect 8256 2756 8263 2853
rect 8296 2747 8303 2763
rect 8156 2127 8163 2693
rect 8236 2607 8243 2743
rect 8276 2707 8283 2743
rect 8256 2556 8263 2593
rect 8176 2536 8203 2543
rect 8176 2527 8183 2536
rect 8216 2187 8223 2473
rect 8156 2096 8193 2103
rect 8156 2076 8163 2096
rect 8216 2067 8223 2173
rect 8116 1607 8123 1793
rect 8116 1547 8123 1573
rect 8176 1556 8183 1593
rect 8196 1576 8203 1593
rect 8236 1343 8243 2513
rect 8276 2343 8283 2613
rect 8316 2547 8323 3053
rect 8256 2336 8283 2343
rect 8256 2287 8263 2336
rect 8256 2263 8263 2273
rect 8336 2263 8343 3713
rect 8376 3707 8383 3996
rect 8396 3927 8403 4153
rect 8416 3547 8423 4013
rect 8576 4007 8583 4273
rect 8516 3996 8543 4003
rect 8456 3647 8463 3993
rect 8516 3867 8523 3996
rect 8516 3807 8523 3853
rect 8496 3627 8503 3723
rect 8547 3676 8553 3683
rect 8356 2267 8363 3493
rect 8436 3367 8443 3573
rect 8456 3527 8463 3613
rect 8476 3487 8483 3503
rect 8396 3227 8403 3243
rect 8436 3236 8443 3353
rect 8256 2256 8283 2263
rect 8316 2256 8343 2263
rect 8256 1807 8263 2113
rect 8296 1387 8303 2243
rect 8356 2087 8363 2093
rect 8376 1847 8383 3173
rect 8396 2076 8403 2133
rect 8416 2083 8423 3223
rect 8456 3207 8463 3223
rect 8496 3147 8503 3613
rect 8556 3407 8563 3633
rect 8576 3243 8583 3953
rect 8596 3287 8603 4753
rect 8616 4507 8623 4896
rect 8676 4696 8703 4703
rect 8696 4607 8703 4696
rect 8616 4307 8623 4493
rect 8676 4456 8683 4493
rect 8736 4476 8743 4613
rect 8756 4467 8763 4933
rect 8776 4727 8783 7053
rect 8796 6107 8803 7793
rect 8816 6387 8823 7693
rect 8876 7487 8883 8493
rect 8896 7827 8903 8693
rect 8936 8507 8943 9433
rect 8936 8267 8943 8303
rect 8876 7376 8883 7413
rect 8916 7067 8923 7613
rect 8936 7587 8943 7833
rect 8956 7627 8963 9333
rect 9036 9256 9043 9913
rect 9156 9756 9183 9763
rect 9216 9756 9223 10193
rect 9236 9787 9243 9953
rect 9156 9667 9163 9756
rect 9056 9496 9083 9503
rect 9116 9496 9143 9503
rect 9056 9467 9063 9496
rect 9136 9287 9143 9496
rect 9016 9187 9023 9243
rect 9076 9007 9083 9253
rect 9116 8996 9123 9233
rect 8976 7687 8983 8893
rect 9136 8827 9143 8963
rect 9136 8796 9143 8813
rect 9176 8767 9183 9613
rect 9216 9163 9223 9713
rect 9256 9276 9263 9993
rect 9276 9727 9283 10233
rect 9316 10047 9323 10656
rect 9416 10467 9423 10673
rect 9336 10387 9343 10453
rect 9336 10236 9343 10373
rect 9356 9967 9363 10433
rect 9396 9987 9403 10193
rect 9396 9956 9403 9973
rect 9296 9663 9303 9773
rect 9276 9656 9303 9663
rect 9276 9467 9283 9656
rect 9336 9527 9343 9923
rect 9316 9476 9323 9513
rect 9296 9447 9303 9463
rect 9376 9447 9383 9953
rect 9416 9923 9423 10153
rect 9396 9916 9423 9923
rect 9336 9287 9343 9313
rect 9216 9156 9243 9163
rect 9196 8787 9203 8993
rect 9016 7867 9023 8013
rect 8976 7576 9003 7583
rect 8996 7507 9003 7576
rect 9016 7567 9023 7833
rect 8936 6887 8943 7433
rect 8996 7327 9003 7473
rect 8996 6867 9003 7313
rect 9016 7047 9023 7373
rect 8916 6727 8923 6863
rect 8916 6547 8923 6603
rect 8836 6396 8843 6533
rect 8936 6387 8943 6583
rect 8856 6047 8863 6373
rect 8976 6127 8983 6413
rect 8876 6067 8883 6103
rect 8876 5916 8883 6013
rect 8756 4427 8763 4453
rect 8796 4407 8803 5913
rect 8896 5907 8903 6033
rect 8656 4187 8663 4203
rect 8696 4196 8703 4273
rect 8676 4167 8683 4183
rect 8616 4027 8623 4093
rect 8616 3267 8623 3793
rect 8636 3667 8643 4093
rect 8736 4067 8743 4253
rect 8816 4247 8823 5693
rect 8836 4547 8843 5653
rect 8856 5263 8863 5423
rect 8876 5263 8883 5433
rect 8896 5407 8903 5423
rect 8916 5383 8923 6053
rect 8936 6047 8943 6123
rect 8936 5947 8943 5973
rect 8956 5636 8963 5933
rect 8976 5927 8983 6113
rect 8976 5407 8983 5613
rect 9016 5607 9023 7033
rect 9036 6847 9043 8733
rect 9076 8527 9083 8733
rect 9056 8047 9063 8493
rect 9136 8327 9143 8473
rect 9216 8323 9223 8793
rect 9196 8316 9223 8323
rect 9136 8296 9143 8313
rect 9176 8147 9183 8303
rect 9216 8087 9223 8316
rect 9136 7836 9143 7893
rect 9156 7847 9163 8073
rect 9196 8036 9203 8053
rect 9236 8047 9243 9156
rect 9336 8983 9343 9273
rect 9356 9016 9363 9053
rect 9316 8967 9323 8983
rect 9336 8976 9363 8983
rect 9256 8727 9263 8873
rect 9256 8067 9263 8713
rect 9356 8587 9363 8976
rect 9376 8767 9383 8953
rect 9356 8547 9363 8573
rect 9296 8536 9323 8543
rect 9296 8507 9303 8536
rect 9156 7827 9163 7833
rect 9076 7356 9083 7393
rect 9116 7356 9123 7373
rect 9136 7347 9143 7573
rect 9156 7367 9163 7563
rect 9196 7556 9203 7793
rect 9176 7427 9183 7543
rect 9216 7487 9223 7543
rect 9096 7327 9103 7343
rect 9236 7287 9243 7773
rect 9256 7127 9263 8053
rect 9276 7547 9283 8033
rect 9296 7747 9303 8373
rect 9336 8347 9343 8523
rect 9376 8507 9383 8753
rect 9356 7816 9363 8473
rect 9396 8467 9403 9916
rect 9416 9476 9443 9483
rect 9416 8487 9423 9413
rect 9436 8387 9443 9476
rect 9456 9367 9463 10453
rect 9476 10227 9483 10453
rect 9596 10427 9603 10736
rect 9676 10707 9683 11133
rect 9856 11127 9863 11163
rect 9896 11143 9903 11163
rect 9896 11136 9923 11143
rect 9836 10916 9843 10933
rect 9796 10903 9803 10913
rect 9796 10896 9823 10903
rect 9876 10827 9883 10923
rect 9896 10887 9903 10933
rect 9916 10907 9923 11136
rect 10056 10923 10063 11176
rect 10056 10916 10083 10923
rect 10116 10916 10123 11113
rect 9696 10696 9723 10703
rect 9676 10483 9683 10693
rect 9716 10567 9723 10696
rect 9736 10507 9743 10683
rect 9896 10667 9903 10873
rect 9936 10747 9943 10913
rect 10076 10827 10083 10916
rect 10136 10887 10143 10903
rect 9936 10696 9943 10733
rect 9956 10716 9963 10813
rect 10196 10736 10203 10873
rect 10007 10716 10023 10723
rect 9976 10667 9983 10703
rect 9656 10476 9683 10483
rect 9656 10436 9663 10476
rect 9676 10387 9683 10423
rect 9576 10203 9583 10373
rect 9556 10196 9583 10203
rect 9476 9907 9483 9963
rect 9676 9923 9683 10233
rect 9736 10147 9743 10493
rect 9876 10407 9883 10423
rect 9836 10236 9843 10373
rect 9876 10207 9883 10393
rect 9756 9963 9763 10093
rect 9816 9987 9823 10133
rect 9756 9956 9783 9963
rect 9656 9916 9683 9923
rect 9476 9483 9483 9893
rect 9696 9756 9723 9763
rect 9516 9487 9523 9733
rect 9676 9647 9683 9743
rect 9716 9707 9723 9756
rect 9836 9647 9843 9773
rect 9856 9687 9863 9973
rect 9936 9756 9943 10653
rect 9876 9707 9883 9743
rect 9976 9727 9983 10193
rect 9996 9967 10003 10413
rect 10016 10407 10023 10716
rect 10156 10716 10183 10723
rect 10216 10716 10223 10733
rect 10156 10667 10163 10716
rect 10016 10307 10023 10393
rect 10036 10216 10043 10393
rect 10236 10227 10243 11173
rect 10416 11163 10423 11173
rect 10396 11156 10423 11163
rect 10596 11143 10603 11163
rect 10596 11136 10623 11143
rect 10296 10883 10303 11133
rect 10556 10887 10563 10893
rect 10616 10887 10623 11136
rect 10636 10947 10643 11163
rect 10636 10927 10643 10933
rect 10296 10876 10323 10883
rect 10316 10627 10323 10876
rect 10576 10767 10583 10883
rect 10396 10736 10423 10743
rect 10256 10407 10263 10613
rect 10356 10427 10363 10443
rect 10396 10427 10403 10736
rect 10456 10703 10463 10733
rect 10696 10716 10703 10753
rect 10716 10727 10723 10893
rect 10716 10707 10723 10713
rect 10436 10696 10463 10703
rect 10276 10216 10283 10413
rect 10296 10403 10303 10423
rect 10336 10407 10343 10423
rect 10296 10396 10323 10403
rect 10256 10167 10263 10203
rect 10296 9987 10303 10193
rect 10316 10167 10323 10396
rect 10476 10256 10483 10693
rect 10596 10447 10603 10453
rect 10556 10347 10563 10443
rect 9996 9943 10003 9953
rect 9996 9936 10023 9943
rect 9996 9707 10003 9936
rect 9856 9503 9863 9673
rect 9836 9496 9863 9503
rect 9476 9476 9503 9483
rect 9636 9283 9643 9293
rect 9636 9276 9663 9283
rect 9596 9023 9603 9253
rect 9636 9087 9643 9276
rect 9716 9256 9723 9313
rect 9576 9016 9603 9023
rect 9636 9016 9643 9073
rect 9576 8987 9583 9016
rect 9616 8987 9623 9003
rect 9536 8807 9543 8953
rect 9616 8783 9623 8833
rect 9596 8776 9623 8783
rect 9456 8316 9483 8323
rect 9396 8296 9403 8313
rect 9296 7507 9303 7573
rect 9336 7527 9343 7803
rect 9376 7747 9383 7803
rect 9296 7356 9303 7493
rect 9336 7356 9343 7473
rect 9396 7447 9403 7533
rect 9356 7336 9363 7353
rect 9416 7327 9423 8073
rect 9456 8027 9463 8233
rect 9476 8147 9483 8316
rect 9496 8307 9503 8573
rect 9556 8567 9563 8773
rect 9556 8536 9563 8553
rect 9516 8247 9523 8493
rect 9536 8467 9543 8533
rect 9616 8487 9623 8776
rect 9656 8296 9663 8473
rect 9696 8287 9703 9233
rect 9856 9227 9863 9496
rect 9876 9487 9883 9593
rect 9936 9256 9943 9293
rect 9896 8996 9903 9053
rect 9716 8707 9723 8993
rect 9916 8867 9923 8983
rect 9776 8796 9803 8803
rect 9756 8767 9763 8793
rect 9776 8567 9783 8796
rect 9876 8796 9883 8853
rect 9816 8707 9823 8783
rect 9776 8536 9793 8543
rect 9776 8507 9783 8536
rect 9836 8543 9843 8673
rect 9836 8536 9863 8543
rect 9856 8507 9863 8536
rect 9836 8327 9843 8433
rect 9476 8056 9483 8133
rect 9516 7827 9523 8133
rect 9636 7803 9643 8273
rect 9676 8227 9683 8283
rect 9836 8283 9843 8313
rect 9916 8283 9923 8313
rect 9836 8276 9863 8283
rect 9896 8276 9923 8283
rect 9696 8087 9703 8213
rect 9896 8147 9903 8276
rect 9696 8056 9703 8073
rect 9736 8056 9753 8063
rect 9716 7847 9723 8043
rect 9756 8027 9763 8053
rect 9836 7836 9843 8133
rect 9916 8027 9923 8073
rect 9796 7816 9823 7823
rect 9636 7796 9663 7803
rect 9436 7527 9443 7543
rect 9436 7327 9443 7513
rect 9056 6807 9063 7093
rect 9116 7076 9123 7093
rect 9096 7027 9103 7063
rect 9136 7047 9143 7063
rect 9096 6747 9103 6973
rect 9096 6416 9103 6733
rect 9116 6627 9123 6853
rect 9136 6447 9143 6833
rect 9176 6747 9183 6843
rect 9196 6616 9223 6623
rect 9176 6587 9183 6603
rect 9116 6396 9123 6413
rect 8856 5256 8883 5263
rect 8876 4687 8883 5256
rect 8896 5376 8923 5383
rect 8896 5083 8903 5376
rect 8976 5147 8983 5393
rect 8916 5107 8923 5143
rect 8956 5127 8963 5143
rect 8896 5076 8923 5083
rect 8916 4956 8923 5076
rect 8936 5067 8943 5123
rect 8976 4963 8983 5133
rect 8996 5107 9003 5473
rect 8956 4956 8983 4963
rect 8896 4936 8903 4953
rect 8936 4907 8943 4943
rect 8936 4807 8943 4893
rect 8876 4663 8883 4673
rect 8976 4667 8983 4956
rect 8856 4656 8883 4663
rect 8776 3976 8783 4033
rect 8756 3947 8763 3963
rect 8776 3736 8803 3743
rect 8656 3687 8663 3713
rect 8716 3687 8723 3713
rect 8756 3547 8763 3723
rect 8796 3647 8803 3736
rect 8676 3263 8683 3503
rect 8656 3256 8683 3263
rect 8556 3236 8583 3243
rect 8436 2787 8443 3053
rect 8496 3036 8503 3073
rect 8536 3036 8543 3053
rect 8436 2556 8443 2773
rect 8456 2587 8463 2653
rect 8476 2567 8483 2613
rect 8496 2147 8503 2953
rect 8556 2767 8563 3236
rect 8616 3223 8623 3253
rect 8616 3216 8643 3223
rect 8516 2667 8523 2763
rect 8607 2757 8621 2764
rect 8576 2727 8583 2743
rect 8614 2705 8621 2757
rect 8636 2747 8643 3193
rect 8656 2807 8663 3256
rect 8676 3047 8683 3223
rect 8656 2767 8663 2793
rect 8676 2727 8683 3033
rect 8596 2698 8621 2705
rect 8516 2607 8523 2653
rect 8516 2167 8523 2283
rect 8556 2267 8563 2283
rect 8416 2076 8443 2083
rect 8236 1336 8263 1343
rect 8296 1336 8303 1353
rect 8076 1167 8083 1283
rect 8196 1147 8203 1173
rect 8276 1147 8283 1323
rect 8176 1067 8183 1113
rect 8196 1096 8203 1133
rect 8216 1087 8223 1093
rect 8036 927 8043 953
rect 7856 336 7883 343
rect 7896 247 7903 343
rect 7616 207 7623 233
rect 7416 127 7423 143
rect 7616 136 7623 193
rect 7696 123 7703 173
rect 8036 127 8043 893
rect 8156 856 8183 863
rect 8076 467 8083 853
rect 8156 667 8163 856
rect 8196 787 8203 843
rect 8096 567 8103 653
rect 8176 603 8183 693
rect 8116 587 8123 603
rect 8156 596 8183 603
rect 7676 116 7703 123
rect 6436 -24 6443 13
rect 8116 -17 8123 343
rect 8196 307 8203 653
rect 8096 -24 8123 -17
rect 8136 -24 8143 233
rect 8196 176 8203 293
rect 8236 143 8243 373
rect 8256 167 8263 1083
rect 8276 1007 8283 1093
rect 8316 867 8323 1633
rect 8376 1616 8383 1693
rect 8396 1667 8403 1783
rect 8396 1407 8403 1583
rect 8436 1307 8443 2076
rect 8476 2047 8483 2073
rect 8556 1787 8563 2253
rect 8596 2187 8603 2698
rect 8616 2123 8623 2293
rect 8596 2116 8623 2123
rect 8456 1167 8463 1333
rect 8476 1327 8483 1593
rect 8536 1307 8543 1343
rect 8456 1116 8463 1133
rect 8496 1116 8503 1153
rect 8556 1147 8563 1323
rect 8536 1087 8543 1133
rect 8376 787 8383 893
rect 8407 856 8423 863
rect 8496 843 8503 893
rect 8576 867 8583 1613
rect 8456 836 8503 843
rect 8396 823 8403 833
rect 8456 823 8463 836
rect 8596 827 8603 2116
rect 8656 2107 8663 2593
rect 8676 2556 8683 2593
rect 8696 2576 8703 3253
rect 8796 3207 8803 3513
rect 8776 3016 8783 3193
rect 8816 3067 8823 4213
rect 8836 3647 8843 4533
rect 8856 4167 8863 4553
rect 8856 3907 8863 4033
rect 8856 3527 8863 3853
rect 8876 3827 8883 4633
rect 8896 4467 8903 4663
rect 8996 4567 9003 5093
rect 9036 4647 9043 6393
rect 9116 6067 9123 6103
rect 9136 6067 9143 6083
rect 9176 6067 9183 6513
rect 9216 6387 9223 6616
rect 9116 5927 9123 5953
rect 9056 5896 9083 5903
rect 9116 5896 9123 5913
rect 9056 5847 9063 5896
rect 9156 5863 9163 5913
rect 9136 5856 9163 5863
rect 9076 5427 9083 5853
rect 9116 5443 9123 5513
rect 9096 5436 9123 5443
rect 8956 4476 8963 4513
rect 8996 4476 9013 4483
rect 8896 4387 8903 4453
rect 8976 4427 8983 4463
rect 9016 4207 9023 4473
rect 8896 3587 8903 4153
rect 8916 3987 8923 4173
rect 8916 3707 8923 3973
rect 8936 3907 8943 4183
rect 8976 3967 8983 4193
rect 8936 3807 8943 3893
rect 8927 3696 8943 3703
rect 8976 3687 8983 3703
rect 8956 3587 8963 3683
rect 8936 3516 8943 3553
rect 8816 2763 8823 3033
rect 8796 2756 8823 2763
rect 8716 2556 8743 2563
rect 8736 2487 8743 2556
rect 8616 2076 8623 2093
rect 8676 2056 8683 2113
rect 8696 2067 8703 2133
rect 8756 2087 8763 2353
rect 8776 2327 8783 2743
rect 8816 2276 8823 2613
rect 8836 2487 8843 3233
rect 8856 3223 8863 3513
rect 8976 3447 8983 3673
rect 8996 3527 9003 4133
rect 9036 4016 9043 4453
rect 9056 4167 9063 5213
rect 9116 4963 9123 5436
rect 9136 5227 9143 5856
rect 9156 5587 9163 5613
rect 9196 5607 9203 5623
rect 9176 5127 9183 5143
rect 9136 5067 9143 5073
rect 9096 4956 9123 4963
rect 9096 4923 9103 4956
rect 9136 4936 9143 5053
rect 9096 4916 9113 4923
rect 9156 4907 9163 4923
rect 9196 4767 9203 5153
rect 9216 4747 9223 5613
rect 9236 5607 9243 6953
rect 9256 6127 9263 6873
rect 9316 6416 9323 7313
rect 9336 6887 9343 7063
rect 9336 6547 9343 6873
rect 9356 6856 9363 6953
rect 9376 6876 9383 6893
rect 9416 6887 9423 7113
rect 9396 6787 9403 6863
rect 9456 6827 9463 6843
rect 9436 6623 9443 6753
rect 9376 6616 9403 6623
rect 9436 6616 9463 6623
rect 9376 6587 9383 6616
rect 9276 6396 9303 6403
rect 9336 6396 9343 6413
rect 9416 6407 9423 6603
rect 9156 4247 9163 4633
rect 9216 4567 9223 4733
rect 9216 4436 9223 4473
rect 9236 4456 9243 4513
rect 9156 4187 9163 4203
rect 9096 4167 9103 4183
rect 9136 4127 9143 4183
rect 9176 4167 9183 4213
rect 9156 4103 9163 4133
rect 9136 4096 9163 4103
rect 9056 3996 9063 4033
rect 9076 4027 9083 4053
rect 9016 3667 9023 3953
rect 8856 3216 8883 3223
rect 8936 3207 8943 3243
rect 8996 3207 9003 3453
rect 9016 3227 9023 3633
rect 8856 2263 8863 2653
rect 8836 2256 8863 2263
rect 8616 1787 8623 1803
rect 8656 1796 8663 1813
rect 8696 1783 8703 1793
rect 8636 1647 8643 1783
rect 8676 1776 8703 1783
rect 8616 1576 8623 1613
rect 8676 1596 8703 1603
rect 8696 1587 8703 1596
rect 8656 1567 8663 1583
rect 8696 1307 8703 1573
rect 8716 1567 8723 1813
rect 8736 1787 8743 1793
rect 8756 1303 8763 2073
rect 8816 1787 8823 2093
rect 8836 1807 8843 2256
rect 8876 1887 8883 3053
rect 8976 3036 8983 3073
rect 8896 2607 8903 3033
rect 9036 2783 9043 3913
rect 9056 3507 9063 3853
rect 9076 3787 9083 3993
rect 9076 3267 9083 3773
rect 9096 3567 9103 4013
rect 9116 3647 9123 3733
rect 9096 3107 9103 3553
rect 9136 3536 9143 4096
rect 9156 3947 9163 4033
rect 9196 3967 9203 4193
rect 9256 3996 9263 5893
rect 9276 4847 9283 6396
rect 9396 6116 9403 6153
rect 9376 6067 9383 6103
rect 9416 6083 9423 6103
rect 9407 6076 9423 6083
rect 9296 5647 9303 6033
rect 9316 5916 9323 5933
rect 9296 5436 9303 5493
rect 9336 5436 9343 5473
rect 9396 5367 9403 6073
rect 9456 5887 9463 6616
rect 9476 6367 9483 7673
rect 9656 7583 9663 7796
rect 9656 7576 9673 7583
rect 9536 7096 9543 7573
rect 9596 7287 9603 7323
rect 9576 7096 9583 7113
rect 9556 6967 9563 7083
rect 9636 7076 9643 7273
rect 9676 6987 9683 7573
rect 9776 7363 9783 7633
rect 9796 7567 9803 7816
rect 9856 7807 9863 7823
rect 9836 7556 9843 7573
rect 9776 7356 9803 7363
rect 9856 7363 9863 7533
rect 9936 7523 9943 9213
rect 9956 8687 9963 9243
rect 9976 8967 9983 9673
rect 9996 9247 10003 9693
rect 9996 8527 10003 8793
rect 10016 8747 10023 9773
rect 10056 9767 10063 9943
rect 10156 9787 10163 9953
rect 10196 9756 10203 9973
rect 10276 9956 10283 9973
rect 10056 9687 10063 9753
rect 10136 9727 10143 9743
rect 10136 9547 10143 9713
rect 10176 9667 10183 9733
rect 10036 9427 10043 9483
rect 10056 9447 10063 9463
rect 10176 9447 10183 9653
rect 10336 9527 10343 10013
rect 10076 8987 10083 9253
rect 10096 9003 10103 9433
rect 10196 9276 10203 9413
rect 10216 9256 10223 9293
rect 10096 8996 10123 9003
rect 10156 8996 10163 9053
rect 10116 8847 10123 8996
rect 10176 8967 10183 8983
rect 10196 8787 10203 9013
rect 10296 8887 10303 9483
rect 10336 9476 10343 9513
rect 10356 9447 10363 9463
rect 10376 9267 10383 9973
rect 10496 9956 10503 9973
rect 10436 9756 10443 9953
rect 10476 9923 10483 9943
rect 10476 9916 10503 9923
rect 10496 9747 10503 9916
rect 10456 9627 10463 9733
rect 10576 9503 10583 10423
rect 10636 9723 10643 10653
rect 10736 10447 10743 11173
rect 10876 11163 10883 11173
rect 10816 11127 10823 11163
rect 10856 11156 10883 11163
rect 10756 10887 10763 10903
rect 10756 10707 10763 10873
rect 10896 10736 10903 10933
rect 10936 10767 10943 11153
rect 11096 11147 11103 11163
rect 10936 10716 10943 10753
rect 10816 10456 10823 10673
rect 10856 10456 10883 10463
rect 10836 10427 10843 10443
rect 10736 10216 10743 10253
rect 10756 10236 10763 10333
rect 10796 10236 10823 10243
rect 10676 9747 10683 10213
rect 10776 10187 10783 10223
rect 10816 10007 10823 10236
rect 10756 9976 10763 9993
rect 10796 9976 10823 9983
rect 10776 9927 10783 9963
rect 10816 9947 10823 9976
rect 10876 9783 10883 10456
rect 10856 9776 10883 9783
rect 10636 9716 10663 9723
rect 10576 9496 10603 9503
rect 10516 9443 10523 9473
rect 10596 9467 10603 9496
rect 10576 9447 10583 9463
rect 10516 9436 10563 9443
rect 10616 9287 10623 9533
rect 10636 9447 10643 9473
rect 10656 9276 10663 9716
rect 10696 9547 10703 9743
rect 10316 8983 10323 9053
rect 10356 9027 10363 9253
rect 10456 9243 10463 9273
rect 10436 9236 10463 9243
rect 10356 8996 10363 9013
rect 10316 8976 10343 8983
rect 10096 8776 10123 8783
rect 10056 8587 10063 8773
rect 10116 8767 10123 8776
rect 10276 8763 10283 8793
rect 10316 8776 10323 8873
rect 10356 8763 10363 8813
rect 10516 8803 10523 9273
rect 10696 9263 10703 9493
rect 10636 9247 10643 9263
rect 10676 9256 10703 9263
rect 10696 9247 10703 9256
rect 10276 8756 10303 8763
rect 10336 8756 10363 8763
rect 10036 8516 10043 8533
rect 10076 8467 10083 8523
rect 9996 8036 10003 8053
rect 10036 8047 10043 8453
rect 10056 8307 10063 8333
rect 10256 8267 10263 8533
rect 10336 8487 10343 8523
rect 10356 8507 10363 8756
rect 10496 8796 10523 8803
rect 10556 8796 10563 8953
rect 10376 8367 10383 8473
rect 10296 8283 10303 8313
rect 10296 8276 10323 8283
rect 10256 8067 10263 8253
rect 9956 7547 9963 8033
rect 9976 7847 9983 8023
rect 10136 7823 10143 7893
rect 10156 7867 10163 8053
rect 10256 8036 10263 8053
rect 10376 8047 10383 8353
rect 10396 8347 10403 8513
rect 10496 8487 10503 8796
rect 10576 8787 10583 8793
rect 10536 8767 10543 8783
rect 10636 8767 10643 9233
rect 10696 8987 10703 9233
rect 10536 8547 10543 8753
rect 10556 8447 10563 8523
rect 10596 8516 10603 8533
rect 10616 8487 10623 8503
rect 10456 8056 10463 8293
rect 10496 8067 10503 8353
rect 10556 8327 10563 8333
rect 10656 8307 10663 8793
rect 10616 8296 10643 8303
rect 10576 8287 10583 8293
rect 10636 8267 10643 8296
rect 10116 7816 10143 7823
rect 9936 7516 9963 7523
rect 9847 7356 9863 7363
rect 9696 7083 9703 7173
rect 9696 7076 9723 7083
rect 9716 6967 9723 7076
rect 9916 7043 9923 7353
rect 9956 7287 9963 7516
rect 10056 7427 10063 7563
rect 10096 7556 10103 7613
rect 10116 7527 10123 7543
rect 9996 7216 10013 7223
rect 9996 7083 10003 7216
rect 10036 7103 10043 7273
rect 10036 7096 10063 7103
rect 9996 7076 10023 7083
rect 9896 7036 9923 7043
rect 9496 6856 9523 6863
rect 9796 6856 9803 6953
rect 9896 6863 9903 6893
rect 9876 6856 9903 6863
rect 9496 6587 9503 6773
rect 9516 6727 9523 6856
rect 10036 6827 10043 7096
rect 9656 6623 9663 6733
rect 9656 6616 9683 6623
rect 9596 6396 9603 6433
rect 9656 6427 9663 6616
rect 9696 6447 9703 6583
rect 9956 6583 9963 6613
rect 10076 6587 10083 6863
rect 9936 6576 9963 6583
rect 9596 5903 9603 6093
rect 9616 6047 9623 6083
rect 9636 6067 9643 6103
rect 9576 5896 9603 5903
rect 9416 5587 9423 5623
rect 9456 5607 9463 5623
rect 9496 5587 9503 5623
rect 9436 5207 9443 5573
rect 9416 5156 9443 5163
rect 9376 4936 9383 5153
rect 9396 5116 9423 5123
rect 9416 5007 9423 5116
rect 9416 4903 9423 4993
rect 9436 4947 9443 5156
rect 9396 4896 9423 4903
rect 9276 4147 9283 4753
rect 9296 4467 9303 4653
rect 9296 4027 9303 4453
rect 9316 4387 9323 4893
rect 9336 4647 9343 4663
rect 9316 4327 9323 4373
rect 9316 4167 9323 4233
rect 9216 3976 9243 3983
rect 9156 3716 9163 3933
rect 9216 3867 9223 3976
rect 9196 3716 9203 3733
rect 9236 3703 9243 3773
rect 9216 3696 9243 3703
rect 9176 3667 9183 3683
rect 9156 3516 9183 3523
rect 9176 3483 9183 3516
rect 9156 3476 9183 3483
rect 9156 3243 9163 3476
rect 9156 3236 9183 3243
rect 9096 3087 9103 3093
rect 9016 2776 9043 2783
rect 9016 2756 9023 2776
rect 8916 2327 8923 2523
rect 8916 2247 8923 2313
rect 8956 2127 8963 2513
rect 8896 2076 8903 2113
rect 8916 1796 8923 1833
rect 8887 1776 8903 1783
rect 8816 1327 8823 1653
rect 8836 1596 8843 1773
rect 8876 1596 8883 1613
rect 8956 1587 8963 2113
rect 8976 1827 8983 2713
rect 8996 2567 9003 2743
rect 9036 2343 9043 2743
rect 9056 2667 9063 2763
rect 9156 2556 9163 3173
rect 9176 2627 9183 3236
rect 9196 3167 9203 3513
rect 9256 3043 9263 3953
rect 9276 3927 9283 3983
rect 9316 3667 9323 4013
rect 9336 4007 9343 4553
rect 9376 4307 9383 4493
rect 9396 4427 9403 4896
rect 9456 4647 9463 5393
rect 9496 5127 9503 5173
rect 9476 4547 9483 4813
rect 9427 4496 9433 4503
rect 9456 4476 9463 4493
rect 9436 4447 9443 4463
rect 9476 4456 9483 4533
rect 9376 4196 9383 4293
rect 9356 4167 9363 4183
rect 9356 3767 9363 4153
rect 9236 3036 9263 3043
rect 9256 3027 9263 3036
rect 9276 2756 9283 3653
rect 9296 2987 9303 3633
rect 9016 2336 9043 2343
rect 9116 2536 9143 2543
rect 8856 1567 8863 1583
rect 8996 1567 9003 2333
rect 9016 2287 9023 2336
rect 9036 2296 9043 2313
rect 9096 2063 9103 2113
rect 9116 2087 9123 2536
rect 9176 2487 9183 2543
rect 9136 2076 9143 2213
rect 9176 2083 9183 2293
rect 9176 2076 9193 2083
rect 9096 2056 9123 2063
rect 9096 1687 9103 2056
rect 9156 1967 9163 2053
rect 9196 1787 9203 2073
rect 9116 1727 9123 1783
rect 9116 1596 9123 1613
rect 9136 1567 9143 1583
rect 8736 1296 8763 1303
rect 8776 1167 8783 1293
rect 8716 1096 8723 1113
rect 8916 1107 8923 1353
rect 8936 1347 8943 1393
rect 9016 1336 9043 1343
rect 8956 1287 8963 1323
rect 9036 1307 9043 1336
rect 8936 1127 8943 1133
rect 8936 1096 8943 1113
rect 8396 816 8463 823
rect 8647 816 8663 823
rect 8276 167 8283 713
rect 8396 683 8403 793
rect 8396 676 8423 683
rect 8416 636 8423 676
rect 8296 343 8303 613
rect 8376 343 8383 453
rect 8296 336 8323 343
rect 8356 336 8383 343
rect 8336 316 8353 323
rect 8476 227 8483 273
rect 8476 156 8483 213
rect 8496 176 8503 773
rect 8676 767 8683 803
rect 8596 616 8603 653
rect 8576 567 8583 613
rect 8616 596 8623 613
rect 8676 603 8683 693
rect 8736 667 8743 1083
rect 8956 1076 8963 1173
rect 9016 1083 9023 1253
rect 9176 1107 9183 1373
rect 9196 1103 9203 1613
rect 9216 1607 9223 2553
rect 9236 1807 9243 2613
rect 9256 2227 9263 2263
rect 9296 1627 9303 2253
rect 9316 2247 9323 2763
rect 9336 2347 9343 3553
rect 9376 3536 9383 3693
rect 9396 3687 9403 4153
rect 9436 3867 9443 4413
rect 9496 4267 9503 5073
rect 9516 4447 9523 5353
rect 9496 3996 9503 4253
rect 9516 4107 9523 4433
rect 9536 4027 9543 5193
rect 9556 5187 9563 5403
rect 9556 4907 9563 5153
rect 9556 4167 9563 4633
rect 9576 4003 9583 5633
rect 9656 5207 9663 6393
rect 9676 5947 9683 6433
rect 9916 6407 9923 6563
rect 9936 6427 9943 6576
rect 9876 6376 9883 6393
rect 9796 6107 9803 6373
rect 9856 6136 9883 6143
rect 9816 6047 9823 6133
rect 9876 6047 9883 6136
rect 9796 5916 9803 5953
rect 9836 5903 9843 5913
rect 9816 5896 9843 5903
rect 9676 5587 9683 5653
rect 9716 5636 9723 5653
rect 9776 5643 9783 5693
rect 9756 5636 9783 5643
rect 9696 5247 9703 5613
rect 9596 4956 9603 5133
rect 9616 5127 9623 5143
rect 9656 5136 9673 5143
rect 9616 4923 9623 4943
rect 9596 4916 9623 4923
rect 9596 4887 9603 4916
rect 9596 4507 9603 4663
rect 9536 3996 9583 4003
rect 9456 3976 9483 3983
rect 9456 3927 9463 3976
rect 9456 3847 9463 3913
rect 9456 3647 9463 3703
rect 9376 3467 9383 3493
rect 9416 3236 9423 3453
rect 9356 2727 9363 3203
rect 9376 3187 9383 3223
rect 9436 3056 9443 3333
rect 9476 2707 9483 3673
rect 9496 3547 9503 3703
rect 9516 3607 9523 3833
rect 9516 3187 9523 3513
rect 9536 3227 9543 3953
rect 9556 3887 9563 3996
rect 9356 2267 9363 2573
rect 9416 2556 9423 2573
rect 9456 2556 9483 2563
rect 9476 2527 9483 2556
rect 9496 2547 9503 3133
rect 9516 2687 9523 2723
rect 9356 2087 9363 2093
rect 9396 2076 9403 2113
rect 9416 2056 9423 2073
rect 9336 1727 9343 1783
rect 9396 1763 9403 1803
rect 9376 1756 9403 1763
rect 9336 1587 9343 1713
rect 9376 1596 9383 1756
rect 9416 1607 9423 1653
rect 9236 1147 9243 1283
rect 9256 1267 9263 1303
rect 9276 1267 9283 1333
rect 9276 1167 9283 1253
rect 9276 1116 9283 1153
rect 9196 1096 9223 1103
rect 8996 1076 9023 1083
rect 8696 627 8703 653
rect 8656 596 8683 603
rect 8596 376 8623 383
rect 8516 356 8543 363
rect 8516 327 8523 356
rect 8616 347 8623 376
rect 8636 176 8663 183
rect 8636 147 8643 176
rect 8716 147 8723 613
rect 8216 136 8243 143
rect 8756 143 8763 1053
rect 8776 147 8783 953
rect 8796 847 8803 993
rect 9256 947 9263 1093
rect 9156 827 9163 843
rect 8936 807 8943 823
rect 8916 747 8923 803
rect 8836 643 8843 673
rect 8867 656 8883 663
rect 8836 636 8863 643
rect 8896 636 8903 713
rect 8856 327 8863 343
rect 8836 307 8843 323
rect 8736 136 8763 143
rect 8816 136 8823 153
rect 9016 87 9023 333
rect 9036 307 9043 633
rect 9116 616 9123 633
rect 9156 616 9163 673
rect 9056 247 9063 363
rect 9096 356 9103 603
rect 9136 596 9143 613
rect 9296 487 9303 1293
rect 9316 647 9323 873
rect 9396 856 9403 873
rect 9336 767 9343 843
rect 9356 827 9363 853
rect 9416 847 9423 893
rect 9356 656 9363 673
rect 9336 636 9343 653
rect 9076 287 9083 343
rect 9136 323 9143 473
rect 9316 383 9323 633
rect 9396 587 9403 673
rect 9436 567 9443 2233
rect 9456 1647 9463 2473
rect 9496 2067 9503 2243
rect 9516 2227 9523 2263
rect 9496 1767 9503 2053
rect 9456 1587 9463 1633
rect 9476 1247 9483 1323
rect 9476 1096 9483 1133
rect 9456 727 9463 1083
rect 9496 1076 9503 1113
rect 9516 1107 9523 1773
rect 9536 587 9543 2693
rect 9556 2227 9563 3853
rect 9596 3607 9603 4493
rect 9616 4427 9623 4893
rect 9636 4403 9643 4913
rect 9656 4787 9663 4943
rect 9656 4707 9663 4773
rect 9656 4427 9663 4693
rect 9676 4547 9683 4793
rect 9696 4667 9703 5233
rect 9716 4807 9723 5573
rect 9736 5507 9743 5623
rect 9736 5427 9743 5433
rect 9716 4487 9723 4673
rect 9716 4427 9723 4443
rect 9636 4396 9663 4403
rect 9636 4196 9643 4213
rect 9656 4207 9663 4396
rect 9616 3647 9623 4153
rect 9596 3536 9603 3573
rect 9636 3287 9643 4133
rect 9656 3687 9663 4193
rect 9676 4167 9683 4413
rect 9696 4147 9703 4393
rect 9716 4187 9723 4413
rect 9716 4047 9723 4173
rect 9736 4167 9743 5413
rect 9776 5147 9783 5403
rect 9816 5127 9823 5403
rect 9836 5087 9843 5896
rect 9856 5347 9863 5433
rect 9896 5187 9903 6103
rect 9936 5687 9943 6413
rect 9956 5643 9963 6453
rect 10076 6396 10083 6433
rect 10096 6416 10103 6453
rect 10116 6136 10143 6143
rect 10136 6107 10143 6136
rect 10156 6127 10163 7853
rect 10176 7647 10183 7833
rect 10236 7827 10243 8023
rect 10276 7907 10283 8023
rect 10296 7836 10323 7843
rect 10376 7836 10383 7893
rect 10176 7527 10183 7633
rect 10176 7507 10183 7513
rect 10276 7356 10283 7433
rect 10236 6867 10243 7113
rect 10256 7096 10263 7113
rect 10296 7103 10303 7836
rect 10316 7547 10323 7563
rect 10356 7556 10363 7633
rect 10476 7567 10483 8043
rect 10576 7816 10583 8053
rect 10596 7867 10603 8253
rect 10536 7587 10543 7813
rect 10596 7796 10603 7853
rect 10336 7527 10343 7543
rect 10376 7427 10383 7543
rect 10476 7347 10483 7553
rect 10536 7527 10543 7573
rect 10296 7096 10323 7103
rect 10056 5916 10063 6093
rect 10256 6067 10263 6873
rect 10276 6856 10283 7083
rect 10316 7067 10323 7096
rect 10476 7087 10483 7113
rect 10516 7107 10523 7343
rect 10536 7147 10543 7373
rect 10556 7356 10563 7373
rect 10616 7127 10623 7543
rect 10636 7387 10643 7833
rect 10656 7827 10663 8293
rect 10676 7567 10683 8073
rect 10696 8056 10703 8313
rect 10716 8087 10723 9733
rect 10816 9476 10823 9493
rect 10696 7667 10703 7933
rect 10716 7907 10723 8043
rect 10696 7527 10703 7653
rect 10736 7567 10743 7913
rect 10636 7107 10643 7373
rect 10276 6396 10283 6433
rect 10356 6423 10363 6563
rect 10376 6447 10383 6583
rect 10336 6416 10363 6423
rect 10336 6376 10343 6416
rect 10296 5936 10303 6353
rect 10316 6136 10323 6353
rect 10356 6136 10363 6393
rect 10336 6007 10343 6123
rect 10396 6116 10403 6933
rect 10516 6896 10523 6933
rect 10536 6903 10543 7063
rect 10536 6896 10563 6903
rect 10556 6867 10563 6896
rect 10536 6747 10543 6863
rect 10576 6747 10583 6873
rect 10536 6607 10543 6713
rect 10576 6623 10583 6733
rect 10656 6623 10663 6813
rect 10556 6616 10583 6623
rect 10616 6616 10643 6623
rect 10656 6616 10683 6623
rect 10476 6387 10483 6573
rect 10096 5916 10103 5933
rect 10036 5747 10043 5903
rect 10076 5887 10083 5903
rect 9956 5636 9983 5643
rect 10116 5627 10123 5913
rect 9916 5143 9923 5173
rect 9856 5063 9863 5143
rect 9896 5136 9923 5143
rect 9836 5056 9863 5063
rect 9776 4927 9783 4953
rect 9796 4767 9803 4933
rect 9836 4923 9843 5056
rect 9876 4947 9883 4993
rect 9956 4947 9963 5613
rect 10036 5607 10043 5623
rect 9976 4987 9983 5593
rect 10007 5436 10023 5443
rect 10056 5436 10063 5453
rect 10036 5407 10043 5423
rect 10116 5387 10123 5593
rect 9836 4916 9863 4923
rect 9756 4607 9763 4663
rect 9756 4503 9763 4593
rect 9756 4496 9783 4503
rect 9756 4407 9763 4473
rect 9756 4227 9763 4353
rect 9736 4016 9743 4133
rect 9756 4007 9763 4213
rect 9676 3467 9683 3993
rect 9776 3807 9783 4496
rect 9796 3967 9803 4393
rect 9836 4227 9843 4793
rect 9856 4687 9863 4893
rect 9936 4707 9943 4913
rect 9936 4667 9943 4693
rect 9956 4667 9963 4933
rect 9876 4447 9883 4473
rect 9896 4443 9903 4613
rect 9936 4456 9943 4513
rect 9896 4436 9923 4443
rect 9836 4196 9843 4213
rect 9876 4207 9883 4273
rect 9716 3736 9723 3773
rect 9736 3747 9743 3773
rect 9556 1347 9563 1793
rect 9576 867 9583 1873
rect 9596 1807 9603 3273
rect 9656 3256 9663 3333
rect 9616 2247 9623 3213
rect 9636 3207 9643 3243
rect 9636 3036 9643 3093
rect 9696 2787 9703 3593
rect 9656 2287 9663 2313
rect 9616 2107 9623 2153
rect 9676 2107 9683 2753
rect 9696 2556 9703 2773
rect 9716 2523 9723 3673
rect 9696 2516 9723 2523
rect 9616 2056 9623 2093
rect 9696 2043 9703 2516
rect 9736 2347 9743 3593
rect 9756 3587 9763 3703
rect 9816 3523 9823 4173
rect 9856 4167 9863 4183
rect 9836 3707 9843 4153
rect 9896 4147 9903 4183
rect 9876 3527 9883 3993
rect 9796 3516 9823 3523
rect 9756 2307 9763 3493
rect 9796 3247 9803 3516
rect 9836 3447 9843 3503
rect 9836 2747 9843 3033
rect 9816 2727 9823 2743
rect 9816 2367 9823 2553
rect 9796 2283 9803 2313
rect 9776 2276 9803 2283
rect 9716 2167 9723 2263
rect 9756 2183 9763 2263
rect 9736 2176 9763 2183
rect 9676 2036 9703 2043
rect 9596 1596 9603 1613
rect 9616 1127 9623 1573
rect 9656 1567 9663 1773
rect 9596 856 9603 1013
rect 9636 927 9643 1273
rect 9636 856 9643 913
rect 9616 787 9623 843
rect 9616 616 9623 733
rect 9576 603 9583 613
rect 9576 596 9603 603
rect 9636 587 9643 603
rect 9316 376 9343 383
rect 9336 347 9343 376
rect 9316 327 9323 343
rect 9116 316 9143 323
rect 9116 136 9123 316
rect 9296 307 9303 323
rect 9376 156 9383 553
rect 9496 323 9503 453
rect 9536 356 9543 373
rect 9496 316 9523 323
rect 9596 156 9603 573
rect 9656 503 9663 1373
rect 9676 1283 9683 2036
rect 9716 1316 9723 2093
rect 9736 1607 9743 2176
rect 9756 2147 9763 2153
rect 9756 2067 9763 2133
rect 9776 1727 9783 2013
rect 9816 1867 9823 2333
rect 9836 2267 9843 2733
rect 9856 2727 9863 3433
rect 9896 3307 9903 4093
rect 9916 3987 9923 4213
rect 9936 4187 9943 4213
rect 9936 3996 9943 4133
rect 9976 4107 9983 4973
rect 10056 4947 10063 5373
rect 10136 5347 10143 5873
rect 10156 5627 10163 5813
rect 10116 5167 10123 5183
rect 10096 5047 10103 5163
rect 10116 4956 10123 4973
rect 10056 4827 10063 4933
rect 10176 4927 10183 5933
rect 10256 5916 10283 5923
rect 10256 5907 10263 5916
rect 10196 5023 10203 5673
rect 10236 5636 10243 5713
rect 10316 5647 10323 5653
rect 10336 5647 10343 5693
rect 10216 5527 10223 5623
rect 10296 5607 10303 5623
rect 10236 5416 10243 5473
rect 10256 5396 10263 5493
rect 10276 5416 10283 5433
rect 10196 5016 10223 5023
rect 10056 4676 10063 4773
rect 9976 3996 9983 4053
rect 9936 3447 9943 3703
rect 9956 3567 9963 3973
rect 10016 3947 10023 4673
rect 10076 4447 10083 4663
rect 10076 4407 10083 4433
rect 9976 3667 9983 3713
rect 9876 3256 9883 3293
rect 9896 3067 9903 3243
rect 9936 3027 9943 3053
rect 9896 3003 9903 3023
rect 9896 2996 9923 3003
rect 9856 2523 9863 2593
rect 9876 2567 9883 2993
rect 9896 2536 9903 2973
rect 9916 2707 9923 2996
rect 9856 2516 9883 2523
rect 9856 2287 9863 2353
rect 9836 2087 9843 2253
rect 9836 1827 9843 2053
rect 9856 2027 9863 2043
rect 9796 1727 9803 1783
rect 9836 1747 9843 1783
rect 9836 1596 9843 1733
rect 9756 1316 9783 1323
rect 9776 1307 9783 1316
rect 9876 1287 9883 1853
rect 9676 1276 9703 1283
rect 9636 496 9663 503
rect 9636 123 9643 496
rect 9656 156 9663 473
rect 9676 407 9683 603
rect 9676 127 9683 393
rect 9696 247 9703 1276
rect 9736 1096 9743 1193
rect 9916 1147 9923 2293
rect 9716 987 9723 1083
rect 9716 616 9723 953
rect 9776 823 9783 973
rect 9776 816 9803 823
rect 9836 807 9843 823
rect 9716 347 9723 473
rect 9776 376 9803 383
rect 9756 327 9763 363
rect 9796 307 9803 376
rect 9816 207 9823 803
rect 9936 767 9943 2473
rect 9956 1367 9963 3193
rect 9976 3183 9983 3653
rect 9996 3207 10003 3513
rect 9976 3176 10003 3183
rect 9976 2807 9983 2993
rect 9976 2487 9983 2793
rect 9996 2487 10003 3176
rect 10036 3147 10043 3973
rect 10056 3267 10063 4293
rect 10096 4167 10103 4183
rect 10076 3987 10083 4163
rect 10076 3767 10083 3853
rect 10076 3527 10083 3753
rect 10096 3516 10103 3913
rect 10116 3827 10123 4653
rect 10136 4196 10143 4913
rect 10196 4687 10203 4933
rect 10176 4456 10183 4493
rect 10156 4407 10163 4443
rect 10216 4423 10223 5016
rect 10196 4416 10223 4423
rect 10176 3743 10183 4133
rect 10196 4007 10203 4416
rect 10256 4287 10263 5333
rect 10276 4696 10283 5133
rect 10316 4947 10323 5633
rect 10356 5156 10363 5453
rect 10416 5447 10423 6133
rect 10496 6123 10503 6573
rect 10536 6396 10543 6433
rect 10556 6427 10563 6616
rect 10596 6567 10603 6603
rect 10636 6507 10643 6616
rect 10596 6376 10603 6453
rect 10676 6367 10683 6616
rect 10716 6227 10723 7373
rect 10736 7363 10743 7553
rect 10756 7387 10763 9273
rect 10796 9027 10803 9463
rect 10836 9427 10843 9463
rect 10856 9227 10863 9776
rect 10896 9256 10903 9293
rect 10916 9287 10923 10453
rect 10936 9927 10943 10453
rect 10936 9243 10943 9413
rect 10916 9236 10943 9243
rect 10816 8827 10823 8983
rect 10876 8887 10883 9003
rect 10776 8796 10783 8813
rect 10836 8767 10843 8783
rect 10776 8483 10783 8493
rect 10776 8476 10803 8483
rect 10836 8087 10843 8303
rect 10776 7927 10783 8053
rect 10776 7816 10803 7823
rect 10776 7783 10783 7816
rect 10776 7776 10803 7783
rect 10776 7527 10783 7573
rect 10736 7356 10763 7363
rect 10796 7356 10803 7776
rect 10836 7356 10843 7413
rect 10736 6927 10743 7333
rect 10776 7327 10783 7343
rect 10856 7327 10863 7373
rect 10756 7096 10763 7133
rect 10736 6876 10743 6913
rect 10816 6603 10823 6873
rect 10896 6827 10903 9213
rect 10916 8087 10923 8533
rect 10956 8087 10963 10773
rect 11016 10747 11023 10903
rect 11076 10787 11083 10913
rect 11096 10907 11103 11113
rect 11196 10887 11203 11133
rect 11016 10707 11023 10733
rect 11076 10467 11083 10753
rect 11116 10716 11123 10733
rect 11196 10703 11203 10873
rect 11176 10696 11203 10703
rect 11027 10456 11043 10463
rect 10996 10236 11003 10273
rect 11056 10267 11063 10443
rect 10916 8056 10923 8073
rect 10936 7847 10943 8043
rect 10976 7627 10983 9773
rect 10996 9527 11003 10193
rect 11056 9747 11063 9973
rect 11096 9787 11103 10293
rect 11196 9947 11203 10696
rect 11216 9907 11223 10453
rect 10996 9267 11003 9513
rect 11236 9476 11243 10933
rect 11256 10667 11263 11216
rect 11296 10947 11303 11183
rect 11296 10456 11303 10713
rect 11316 10287 11323 10443
rect 11316 10256 11343 10263
rect 11276 10236 11303 10243
rect 11276 10203 11283 10236
rect 11276 10196 11303 10203
rect 11276 10187 11283 10196
rect 11296 9967 11303 10196
rect 11336 10007 11343 10256
rect 11256 9927 11263 9963
rect 11336 9943 11343 9993
rect 11316 9936 11343 9943
rect 11116 9276 11123 9433
rect 11216 9427 11223 9463
rect 11256 9447 11263 9463
rect 11276 9307 11283 9483
rect 10976 7447 10983 7613
rect 10996 7527 11003 9013
rect 11036 8563 11043 8813
rect 11056 8807 11063 9273
rect 11176 9256 11183 9293
rect 11096 8887 11103 9003
rect 11136 8996 11143 9013
rect 11116 8827 11123 8983
rect 11056 8763 11063 8793
rect 11056 8756 11083 8763
rect 11036 8556 11063 8563
rect 11056 8536 11063 8556
rect 11036 8367 11043 8523
rect 11016 8316 11043 8323
rect 11076 8316 11103 8323
rect 11016 8207 11023 8316
rect 11096 8287 11103 8316
rect 10996 7383 11003 7493
rect 11036 7467 11043 7543
rect 10976 7376 11003 7383
rect 10956 7087 10963 7333
rect 10976 7063 10983 7376
rect 11016 7356 11023 7433
rect 11036 7103 11043 7413
rect 11056 7387 11063 7823
rect 11096 7543 11103 7573
rect 11076 7536 11103 7543
rect 11016 7096 11043 7103
rect 11016 7076 11023 7096
rect 10976 7056 11003 7063
rect 11036 6887 11043 7063
rect 11056 6843 11063 6913
rect 10996 6647 11003 6843
rect 11036 6836 11063 6843
rect 10796 6596 10823 6603
rect 10796 6563 10803 6596
rect 10996 6587 11003 6603
rect 10796 6556 10823 6563
rect 10816 6416 10823 6433
rect 10796 6396 10803 6413
rect 10836 6396 10843 6493
rect 10476 6116 10503 6123
rect 10336 4936 10343 4993
rect 10356 4916 10363 4973
rect 10376 4936 10383 4993
rect 10416 4923 10423 5123
rect 10396 4916 10423 4923
rect 10296 4667 10303 4683
rect 10216 3996 10223 4073
rect 10256 3996 10263 4273
rect 10196 3976 10203 3993
rect 10236 3843 10243 3973
rect 10216 3836 10243 3843
rect 10176 3736 10203 3743
rect 10196 3703 10203 3736
rect 10136 3667 10143 3703
rect 10176 3696 10203 3703
rect 10136 3516 10143 3533
rect 10076 3496 10083 3513
rect 10116 3467 10123 3503
rect 10036 2827 10043 3033
rect 10056 2987 10063 3033
rect 10016 2707 10023 2743
rect 10016 2327 10023 2493
rect 10016 2296 10023 2313
rect 9996 2227 10003 2283
rect 9976 1387 9983 2113
rect 10016 1767 10023 2093
rect 10036 2047 10043 2713
rect 10076 2507 10083 3453
rect 10156 3287 10163 3673
rect 10096 3007 10103 3223
rect 10156 3056 10163 3213
rect 10176 3187 10183 3653
rect 10196 3487 10203 3533
rect 10096 2727 10103 2973
rect 10116 2867 10123 3053
rect 10176 3043 10183 3053
rect 10196 3043 10203 3273
rect 10216 3227 10223 3836
rect 10236 3227 10243 3813
rect 10256 3347 10263 3533
rect 10176 3036 10203 3043
rect 10116 2536 10123 2793
rect 10076 1827 10083 2333
rect 10096 2307 10103 2513
rect 10096 2247 10103 2293
rect 10116 2056 10123 2493
rect 10156 1883 10163 2793
rect 10136 1876 10163 1883
rect 10056 1667 10063 1783
rect 10016 1387 10023 1613
rect 10036 1596 10043 1653
rect 10076 1596 10083 1633
rect 9996 1296 10023 1303
rect 9996 1167 10003 1296
rect 9996 1096 10003 1153
rect 9976 1047 9983 1083
rect 10016 1076 10023 1273
rect 10036 1096 10043 1333
rect 10096 1287 10103 1783
rect 10056 856 10063 933
rect 10096 856 10103 1253
rect 9836 656 9843 693
rect 10116 623 10123 1353
rect 9996 616 10023 623
rect 10096 616 10123 623
rect 9836 376 9843 393
rect 9836 176 9843 233
rect 9856 227 9863 373
rect 9876 347 9883 363
rect 9896 347 9903 393
rect 9996 367 10003 616
rect 10136 487 10143 1876
rect 10156 267 10163 1813
rect 10176 407 10183 2253
rect 10196 1303 10203 3013
rect 10216 2727 10223 3153
rect 10256 3087 10263 3333
rect 10276 3327 10283 3993
rect 10296 3727 10303 4593
rect 10316 3687 10323 4653
rect 10416 4476 10423 4673
rect 10436 4667 10443 6093
rect 10476 5787 10483 6116
rect 10516 6023 10523 6173
rect 10656 6067 10663 6083
rect 10516 6016 10543 6023
rect 10536 5936 10543 6016
rect 10516 5916 10523 5933
rect 10556 5916 10583 5923
rect 10576 5887 10583 5916
rect 10456 5656 10483 5663
rect 10456 5527 10463 5656
rect 10656 5607 10663 5673
rect 10496 5436 10523 5443
rect 10576 5436 10583 5473
rect 10456 4503 10463 5173
rect 10496 5167 10503 5436
rect 10536 5207 10543 5403
rect 10676 5207 10683 6213
rect 10436 4496 10463 4503
rect 10436 4467 10443 4496
rect 10396 4447 10403 4463
rect 10396 4367 10403 4433
rect 10336 4196 10343 4293
rect 10376 4196 10383 4213
rect 10456 4047 10463 4473
rect 10476 4007 10483 5133
rect 10536 5027 10543 5193
rect 10636 5176 10643 5193
rect 10696 5143 10703 5933
rect 10716 5896 10743 5903
rect 10716 5647 10723 5896
rect 10756 5876 10763 6193
rect 10816 6136 10823 6353
rect 10776 5656 10783 5713
rect 10816 5647 10823 5893
rect 10816 5627 10823 5633
rect 10776 5436 10783 5493
rect 10836 5436 10843 5473
rect 10616 5007 10623 5143
rect 10676 5136 10703 5143
rect 10556 4976 10583 4983
rect 10536 4647 10543 4663
rect 10496 4527 10503 4533
rect 10336 3847 10343 3973
rect 10336 3736 10363 3743
rect 10396 3736 10403 3953
rect 10416 3747 10423 3993
rect 10476 3947 10483 3963
rect 10336 3547 10343 3736
rect 10376 3627 10383 3723
rect 10376 3483 10383 3553
rect 10316 3463 10323 3483
rect 10356 3476 10383 3483
rect 10356 3467 10363 3476
rect 10316 3456 10343 3463
rect 10236 2947 10243 3033
rect 10216 1347 10223 2353
rect 10236 2347 10243 2933
rect 10276 2767 10283 3313
rect 10296 3207 10303 3233
rect 10336 3067 10343 3456
rect 10396 3207 10403 3223
rect 10316 3003 10323 3053
rect 10356 3027 10363 3193
rect 10376 3067 10383 3203
rect 10316 2996 10343 3003
rect 10336 2987 10343 2996
rect 10256 2647 10263 2743
rect 10256 2507 10263 2633
rect 10236 2227 10243 2263
rect 10296 1627 10303 2553
rect 10316 2527 10323 2713
rect 10336 2567 10343 2753
rect 10356 2707 10363 2953
rect 10356 2536 10363 2693
rect 10316 2267 10323 2293
rect 10336 2056 10343 2493
rect 10356 2227 10363 2333
rect 10376 2327 10383 2523
rect 10376 2207 10383 2313
rect 10376 2047 10383 2193
rect 10396 2167 10403 3173
rect 10416 2887 10423 3713
rect 10436 3507 10443 3833
rect 10436 3007 10443 3073
rect 10476 2947 10483 3913
rect 10496 2967 10503 4513
rect 10516 3947 10523 4453
rect 10536 4227 10543 4633
rect 10556 4567 10563 4976
rect 10596 4907 10603 4943
rect 10676 4927 10683 5136
rect 10556 4063 10563 4553
rect 10576 4507 10583 4663
rect 10676 4587 10683 4913
rect 10596 4183 10603 4453
rect 10636 4407 10643 4443
rect 10676 4427 10683 4443
rect 10576 4167 10583 4183
rect 10596 4176 10623 4183
rect 10576 4147 10583 4153
rect 10536 4056 10563 4063
rect 10536 3967 10543 4056
rect 10356 2027 10363 2043
rect 10336 1796 10343 1853
rect 10316 1767 10323 1783
rect 10276 1616 10293 1623
rect 10256 1567 10263 1613
rect 10196 1296 10223 1303
rect 10236 1247 10243 1283
rect 10256 1267 10263 1303
rect 10196 807 10203 1113
rect 10276 1087 10283 1103
rect 9816 156 9823 173
rect 9856 156 9863 193
rect 10056 136 10063 253
rect 10176 167 10183 353
rect 10196 327 10203 753
rect 10216 127 10223 893
rect 10236 847 10243 953
rect 10296 887 10303 1333
rect 10316 1127 10323 1753
rect 10336 1307 10343 1583
rect 10336 1107 10343 1293
rect 10356 927 10363 1783
rect 10376 1067 10383 1593
rect 10416 1587 10423 2873
rect 10436 2776 10463 2783
rect 10436 2727 10443 2776
rect 10476 2296 10483 2333
rect 10456 1827 10463 2233
rect 10416 1127 10423 1303
rect 10456 1227 10463 1293
rect 10476 1147 10483 2093
rect 10496 1187 10503 2733
rect 10516 2127 10523 3733
rect 10536 3707 10543 3873
rect 10536 2967 10543 3693
rect 10556 3227 10563 4033
rect 10576 3847 10583 4113
rect 10596 3867 10603 3973
rect 10616 3907 10623 4176
rect 10636 3767 10643 3993
rect 10576 3683 10583 3723
rect 10576 3676 10603 3683
rect 10596 3516 10603 3676
rect 10636 3516 10643 3553
rect 10576 3496 10583 3513
rect 10616 3256 10643 3263
rect 10596 3147 10603 3243
rect 10636 3067 10643 3256
rect 10576 3016 10583 3033
rect 10556 2987 10563 3003
rect 10536 2747 10543 2933
rect 10556 2767 10563 2953
rect 10576 2743 10583 2973
rect 10556 2736 10583 2743
rect 10536 2107 10543 2573
rect 10556 2247 10563 2736
rect 10576 2556 10583 2593
rect 10596 2576 10603 2713
rect 10616 2587 10623 3053
rect 10636 3007 10643 3053
rect 10656 2807 10663 4213
rect 10696 4127 10703 5113
rect 10676 3996 10683 4053
rect 10716 4027 10723 5193
rect 10796 5147 10803 5403
rect 10856 5207 10863 6473
rect 10916 6376 10943 6383
rect 10936 6247 10943 6376
rect 11016 6283 11023 6813
rect 11076 6596 11083 6613
rect 11096 6527 11103 6893
rect 11036 6416 11043 6513
rect 11116 6487 11123 8073
rect 11156 8007 11163 8023
rect 11176 6327 11183 8973
rect 11276 8816 11283 8973
rect 11256 8536 11263 8773
rect 11296 8767 11303 8783
rect 11236 8316 11263 8323
rect 11216 8023 11223 8313
rect 11236 8187 11243 8316
rect 11196 8016 11223 8023
rect 11276 7947 11283 8523
rect 11296 8316 11303 8353
rect 11236 7836 11243 7873
rect 11276 7836 11303 7843
rect 11296 7807 11303 7836
rect 11236 7543 11243 7593
rect 11236 7536 11263 7543
rect 10996 6276 11023 6283
rect 10876 6127 10883 6233
rect 10896 5607 10903 5713
rect 10916 5267 10923 5913
rect 10976 5647 10983 6053
rect 10996 6043 11003 6276
rect 11016 6067 11023 6103
rect 11036 6047 11043 6083
rect 10996 6036 11023 6043
rect 11016 5936 11023 6036
rect 11036 5916 11043 5933
rect 11016 5636 11023 5673
rect 10956 5487 10963 5623
rect 10856 5123 10863 5143
rect 10856 5116 10883 5123
rect 10856 4963 10863 5093
rect 10776 4956 10803 4963
rect 10836 4956 10863 4963
rect 10736 4607 10743 4933
rect 10776 4687 10783 4956
rect 10856 4923 10863 4956
rect 10836 4916 10863 4923
rect 10756 4607 10763 4663
rect 10756 4543 10763 4593
rect 10776 4567 10783 4643
rect 10736 4536 10763 4543
rect 10736 4407 10743 4536
rect 10736 4123 10743 4193
rect 10776 4187 10783 4473
rect 10796 4427 10803 4653
rect 10816 4227 10823 4693
rect 10836 4207 10843 4916
rect 10876 4627 10883 5116
rect 10916 4907 10923 5163
rect 10936 5067 10943 5413
rect 10996 5403 11003 5453
rect 11036 5416 11043 5433
rect 10996 5396 11023 5403
rect 10896 4496 10903 4573
rect 10916 4527 10923 4673
rect 10856 4476 10883 4483
rect 10856 4443 10863 4476
rect 10856 4436 10883 4443
rect 10796 4127 10803 4203
rect 10856 4167 10863 4183
rect 10736 4116 10763 4123
rect 10696 3927 10703 3983
rect 10676 3607 10683 3733
rect 10616 2556 10643 2563
rect 10636 2547 10643 2556
rect 10656 2527 10663 2773
rect 10676 2767 10683 3513
rect 10696 3507 10703 3533
rect 10716 2987 10723 3953
rect 10736 3167 10743 3933
rect 10756 3527 10763 4116
rect 10756 3047 10763 3213
rect 10636 2287 10643 2513
rect 10516 2067 10523 2073
rect 10556 2056 10563 2173
rect 10656 2107 10663 2513
rect 10676 2247 10683 2263
rect 10696 2247 10703 2553
rect 10756 2527 10763 3033
rect 10516 2043 10523 2053
rect 10516 2036 10543 2043
rect 10536 1836 10603 1843
rect 10516 1767 10523 1813
rect 10536 1767 10543 1836
rect 10596 1816 10603 1836
rect 10696 1807 10703 2233
rect 10736 2207 10743 2263
rect 10576 1596 10583 1753
rect 10616 1596 10623 1613
rect 10696 1607 10703 1793
rect 10536 1576 10563 1583
rect 10536 1567 10543 1576
rect 10716 1367 10723 2093
rect 10756 2063 10763 2273
rect 10776 2107 10783 4013
rect 10796 3067 10803 4033
rect 10816 3787 10823 4053
rect 10816 3667 10823 3773
rect 10836 3727 10843 4013
rect 10876 3947 10883 4436
rect 10936 4167 10943 4193
rect 10916 3703 10923 4153
rect 10956 4047 10963 5193
rect 10976 4067 10983 5153
rect 11076 4956 11083 5373
rect 11096 5127 11103 5893
rect 11116 4983 11123 5633
rect 11136 5187 11143 5653
rect 11136 5156 11143 5173
rect 11156 5167 11163 5653
rect 11156 5107 11163 5123
rect 11116 4976 11143 4983
rect 10996 4647 11003 4663
rect 11056 4587 11063 4683
rect 10996 4003 11003 4553
rect 11056 4196 11063 4273
rect 10976 3996 11003 4003
rect 10896 3696 10923 3703
rect 10856 3516 10863 3533
rect 10916 3227 10923 3513
rect 10836 3087 10843 3203
rect 10796 2567 10803 2953
rect 10816 2576 10823 2773
rect 10836 2607 10843 2773
rect 10856 2563 10863 2993
rect 10836 2556 10863 2563
rect 10856 2547 10863 2556
rect 10736 2056 10763 2063
rect 10796 2056 10803 2153
rect 10516 1163 10523 1193
rect 10496 1156 10523 1163
rect 10276 836 10283 853
rect 10256 807 10263 823
rect 10256 647 10263 793
rect 10296 663 10303 793
rect 10316 727 10323 843
rect 10276 656 10303 663
rect 10276 547 10283 656
rect 10316 607 10323 613
rect 10256 356 10263 393
rect 10276 176 10283 393
rect 10316 376 10323 493
rect 10336 347 10343 853
rect 10396 807 10403 1113
rect 10436 463 10443 1133
rect 10496 1116 10503 1156
rect 10516 1096 10523 1113
rect 10536 907 10543 1353
rect 10736 1347 10743 2056
rect 10776 2027 10783 2043
rect 10756 1747 10763 1813
rect 10776 1727 10783 2013
rect 10796 1767 10803 2013
rect 10816 1827 10823 2033
rect 10836 2027 10843 2513
rect 10856 2307 10863 2533
rect 10876 2527 10883 3033
rect 10856 1816 10863 2093
rect 10836 1787 10843 1803
rect 10796 1616 10803 1733
rect 10596 1287 10603 1313
rect 10756 1303 10763 1553
rect 10656 1247 10663 1303
rect 10696 1247 10703 1303
rect 10736 1296 10763 1303
rect 10656 1127 10663 1233
rect 10536 747 10543 803
rect 10556 636 10563 713
rect 10516 607 10523 633
rect 10536 616 10543 633
rect 10576 587 10583 623
rect 10616 587 10623 633
rect 10507 496 10513 503
rect 10436 456 10463 463
rect 10356 347 10363 363
rect 9616 116 9643 123
rect 10036 107 10043 123
rect 10456 107 10463 456
rect 10476 287 10483 323
rect 10536 136 10543 153
rect 10636 127 10643 433
rect 10696 307 10703 1173
rect 10716 1127 10723 1253
rect 10736 1136 10743 1273
rect 10756 1116 10763 1213
rect 10716 367 10723 843
rect 10796 836 10803 1413
rect 10776 616 10783 653
rect 10736 356 10743 433
rect 10716 156 10723 193
rect 10736 176 10743 293
rect 10816 127 10823 1333
rect 10836 167 10843 1753
rect 10856 147 10863 1773
rect 10876 1287 10883 2293
rect 10896 443 10903 3013
rect 10916 2807 10923 3213
rect 10936 3207 10943 3793
rect 10956 3687 10963 3973
rect 10956 2807 10963 3673
rect 10976 3547 10983 3693
rect 10976 2987 10983 3533
rect 10996 2803 11003 3753
rect 10976 2796 11003 2803
rect 10936 2287 10943 2593
rect 10936 1767 10943 2213
rect 10956 1867 10963 2573
rect 10976 2147 10983 2796
rect 10976 1787 10983 2113
rect 10996 1827 11003 2773
rect 11016 2727 11023 4033
rect 11036 3047 11043 3993
rect 11076 3716 11083 4913
rect 11096 4667 11103 4943
rect 11096 4227 11103 4633
rect 11116 4476 11123 4633
rect 11136 4567 11143 4976
rect 11156 4476 11163 4513
rect 11096 4027 11103 4183
rect 11076 3536 11083 3653
rect 11096 3527 11103 4013
rect 11056 3187 11063 3223
rect 11056 3027 11063 3173
rect 11036 2787 11043 3003
rect 11056 2547 11063 2973
rect 11076 2967 11083 3003
rect 11076 2747 11083 2813
rect 11096 2607 11103 3213
rect 11036 2507 11043 2523
rect 11016 2267 11023 2313
rect 11016 2076 11023 2253
rect 11056 2107 11063 2333
rect 11076 2307 11083 2493
rect 11076 2083 11083 2293
rect 11056 2076 11083 2083
rect 11076 2043 11083 2076
rect 11056 2036 11083 2043
rect 11056 1796 11063 2036
rect 11096 1883 11103 2533
rect 11076 1876 11103 1883
rect 10916 1367 10923 1573
rect 10936 1427 10943 1753
rect 10936 1247 10943 1343
rect 10996 1267 11003 1563
rect 11016 1327 11023 1373
rect 10976 1136 10983 1153
rect 10996 1116 11003 1133
rect 10876 436 10903 443
rect 10876 187 10883 436
rect 10896 347 10903 413
rect 10916 187 10923 853
rect 11036 836 11043 1333
rect 11056 843 11063 1153
rect 11076 867 11083 1876
rect 11056 836 11083 843
rect 11016 687 11023 823
rect 10976 427 10983 673
rect 10996 636 11003 653
rect 11016 387 11023 413
rect 11036 367 11043 413
rect 10996 347 11003 363
rect 10956 176 10963 313
rect 11096 187 11103 1853
rect 11116 387 11123 4013
rect 11136 3767 11143 4213
rect 11136 2787 11143 3733
rect 11156 3687 11163 4183
rect 11176 4027 11183 5893
rect 11196 4647 11203 7513
rect 11256 7356 11263 7393
rect 11296 7356 11323 7363
rect 11316 7327 11323 7356
rect 11256 7027 11263 7063
rect 11216 6876 11223 6913
rect 11256 6876 11263 6893
rect 11276 6856 11303 6863
rect 11296 6647 11303 6856
rect 11256 6616 11283 6623
rect 11316 6616 11323 6913
rect 11216 6376 11223 6573
rect 11256 6507 11263 6616
rect 11256 6387 11263 6493
rect 11216 5907 11223 6313
rect 11256 6087 11263 6103
rect 11276 6067 11283 6083
rect 11296 5987 11303 6103
rect 11316 5883 11323 6293
rect 11296 5876 11323 5883
rect 11216 5807 11223 5873
rect 11276 5687 11283 5853
rect 11256 5623 11263 5653
rect 11236 5616 11263 5623
rect 11196 4016 11203 4613
rect 11216 4047 11223 5153
rect 11216 3996 11223 4013
rect 11156 3227 11163 3513
rect 11176 3207 11183 3293
rect 11196 3167 11203 3973
rect 11236 3963 11243 5616
rect 11256 5436 11263 5453
rect 11276 5427 11283 5643
rect 11296 5436 11323 5443
rect 11316 5407 11323 5436
rect 11336 5387 11343 9893
rect 11256 3967 11263 5373
rect 11296 4707 11303 4943
rect 11307 4696 11323 4703
rect 11276 4587 11283 4683
rect 11316 4676 11323 4696
rect 11216 3956 11243 3963
rect 11216 3203 11223 3956
rect 11276 3536 11283 4373
rect 11296 3747 11303 4663
rect 11336 4607 11343 4663
rect 11336 3743 11343 4493
rect 11356 3987 11363 8533
rect 11336 3736 11363 3743
rect 11336 3687 11343 3703
rect 11316 3567 11323 3683
rect 11236 3516 11263 3523
rect 11236 3227 11243 3516
rect 11216 3196 11243 3203
rect 11176 2727 11183 2743
rect 11136 2287 11143 2593
rect 11156 2367 11163 2723
rect 11196 2347 11203 2773
rect 11196 2296 11203 2313
rect 11136 1147 11143 2093
rect 11136 807 11143 833
rect 11156 407 11163 2133
rect 11216 1903 11223 2793
rect 11196 1896 11223 1903
rect 11176 1607 11183 1813
rect 11176 1543 11183 1593
rect 11196 1567 11203 1896
rect 11236 1883 11243 3196
rect 11276 3016 11283 3213
rect 11256 2967 11263 3003
rect 11316 2983 11323 3223
rect 11336 3187 11343 3673
rect 11296 2976 11323 2983
rect 11296 2547 11303 2976
rect 11256 2227 11263 2493
rect 11256 2076 11263 2213
rect 11276 2127 11283 2513
rect 11316 2507 11323 2523
rect 11296 2076 11303 2113
rect 11216 1876 11243 1883
rect 11216 1763 11223 1876
rect 11296 1816 11303 1833
rect 11236 1787 11243 1803
rect 11256 1796 11283 1803
rect 11216 1756 11243 1763
rect 11176 1536 11203 1543
rect 11196 1316 11203 1536
rect 11176 447 11183 1273
rect 11236 1103 11243 1756
rect 11256 1727 11263 1796
rect 11256 1596 11263 1713
rect 11296 1563 11303 1753
rect 11316 1596 11323 2313
rect 11276 1556 11303 1563
rect 11196 647 11203 1103
rect 11216 1096 11243 1103
rect 11196 376 11203 393
rect 10976 156 10983 173
rect 11216 147 11223 1096
rect 11236 803 11243 873
rect 11236 796 11263 803
rect 11256 427 11263 623
rect 11336 367 11343 3153
rect 11356 2587 11363 3736
rect 11356 207 11363 2533
rect 10556 116 10573 123
<< m3contact >>
rect 2733 11233 2747 11247
rect 613 11213 627 11227
rect 793 11213 807 11227
rect 933 11213 947 11227
rect 973 11213 987 11227
rect 573 11173 587 11187
rect 553 11153 567 11167
rect 1013 11193 1027 11207
rect 1353 11213 1367 11227
rect 1613 11213 1627 11227
rect 1793 11213 1807 11227
rect 1893 11213 1907 11227
rect 2033 11213 2047 11227
rect 633 11173 647 11187
rect 773 11173 787 11187
rect 933 11173 947 11187
rect 333 11133 347 11147
rect 573 11133 587 11147
rect 193 10913 207 10927
rect 373 10913 387 10927
rect 73 10893 87 10907
rect 193 10873 207 10887
rect 533 10893 547 10907
rect 473 10853 487 10867
rect 233 10733 247 10747
rect 313 10733 327 10747
rect 453 10733 467 10747
rect 533 10733 547 10747
rect 173 10673 187 10687
rect 53 10493 67 10507
rect 13 10233 27 10247
rect 13 10193 27 10207
rect 173 10393 187 10407
rect 153 10353 167 10367
rect 53 9973 67 9987
rect 213 10333 227 10347
rect 193 10273 207 10287
rect 273 10233 287 10247
rect 233 10153 247 10167
rect 253 10153 267 10167
rect 213 9873 227 9887
rect 153 9733 167 9747
rect 193 9733 207 9747
rect 253 9973 267 9987
rect 273 9913 287 9927
rect 173 9633 187 9647
rect 233 9633 247 9647
rect 153 9473 167 9487
rect 33 9173 47 9187
rect 53 9173 67 9187
rect 153 8993 167 9007
rect 193 9473 207 9487
rect 413 10713 427 10727
rect 513 10713 527 10727
rect 513 10653 527 10667
rect 373 10533 387 10547
rect 453 10453 467 10467
rect 413 10433 427 10447
rect 393 10393 407 10407
rect 393 10273 407 10287
rect 313 9853 327 9867
rect 353 9853 367 9867
rect 253 9453 267 9467
rect 273 9173 287 9187
rect 373 9253 387 9267
rect 193 8973 207 8987
rect 233 8853 247 8867
rect 253 8813 267 8827
rect 213 8773 227 8787
rect 313 8993 327 9007
rect 513 10433 527 10447
rect 473 10233 487 10247
rect 513 10233 527 10247
rect 413 10213 427 10227
rect 453 10213 467 10227
rect 533 10193 547 10207
rect 493 10113 507 10127
rect 413 9913 427 9927
rect 553 9873 567 9887
rect 433 9733 447 9747
rect 453 9713 467 9727
rect 553 9713 567 9727
rect 433 9693 447 9707
rect 413 9633 427 9647
rect 473 9633 487 9647
rect 513 9473 527 9487
rect 473 9313 487 9327
rect 333 8813 347 8827
rect 993 11173 1007 11187
rect 1193 11173 1207 11187
rect 1233 11173 1247 11187
rect 953 11153 967 11167
rect 733 10953 747 10967
rect 693 10933 707 10947
rect 673 10873 687 10887
rect 593 10813 607 10827
rect 633 10713 647 10727
rect 693 10693 707 10707
rect 653 10673 667 10687
rect 713 10673 727 10687
rect 693 10513 707 10527
rect 613 10413 627 10427
rect 673 10453 687 10467
rect 753 10933 767 10947
rect 733 10493 747 10507
rect 653 10433 667 10447
rect 693 10433 707 10447
rect 873 10853 887 10867
rect 893 10813 907 10827
rect 933 10873 947 10887
rect 1053 10913 1067 10927
rect 993 10873 1007 10887
rect 1153 10893 1167 10907
rect 1173 10873 1187 10887
rect 1053 10833 1067 10847
rect 953 10773 967 10787
rect 913 10713 927 10727
rect 913 10693 927 10707
rect 753 10413 767 10427
rect 633 10333 647 10347
rect 733 10313 747 10327
rect 593 10233 607 10247
rect 613 10233 627 10247
rect 613 10153 627 10167
rect 633 10113 647 10127
rect 593 10033 607 10047
rect 593 9953 607 9967
rect 633 9933 647 9947
rect 673 9833 687 9847
rect 693 9833 707 9847
rect 733 10193 747 10207
rect 713 9753 727 9767
rect 633 9313 647 9327
rect 693 9473 707 9487
rect 673 9453 687 9467
rect 653 9293 667 9307
rect 693 9333 707 9347
rect 713 9333 727 9347
rect 673 9273 687 9287
rect 593 9253 607 9267
rect 573 9093 587 9107
rect 433 8993 447 9007
rect 713 9173 727 9187
rect 933 10653 947 10667
rect 1173 10773 1187 10787
rect 1473 11173 1487 11187
rect 1413 10913 1427 10927
rect 1453 10913 1467 10927
rect 1333 10813 1347 10827
rect 1433 10893 1447 10907
rect 1393 10793 1407 10807
rect 1433 10773 1447 10787
rect 1193 10733 1207 10747
rect 1213 10713 1227 10727
rect 1393 10713 1407 10727
rect 1413 10693 1427 10707
rect 1453 10733 1467 10747
rect 1493 10693 1507 10707
rect 1193 10673 1207 10687
rect 1373 10673 1387 10687
rect 1153 10533 1167 10547
rect 1153 10493 1167 10507
rect 1233 10453 1247 10467
rect 893 10373 907 10387
rect 973 10333 987 10347
rect 873 10253 887 10267
rect 873 9933 887 9947
rect 893 9913 907 9927
rect 1013 9973 1027 9987
rect 1173 10273 1187 10287
rect 1373 10433 1387 10447
rect 1453 10433 1467 10447
rect 1533 11173 1547 11187
rect 1813 11193 1827 11207
rect 1733 11173 1747 11187
rect 1773 11173 1787 11187
rect 1873 11153 1887 11167
rect 1733 10953 1747 10967
rect 1873 10953 1887 10967
rect 1673 10913 1687 10927
rect 1713 10913 1727 10927
rect 1753 10913 1767 10927
rect 1533 10893 1547 10907
rect 1553 10893 1567 10907
rect 1513 10653 1527 10667
rect 1393 10393 1407 10407
rect 1493 10393 1507 10407
rect 1173 10033 1187 10047
rect 1073 9953 1087 9967
rect 933 9913 947 9927
rect 913 9893 927 9907
rect 1393 10173 1407 10187
rect 1473 10053 1487 10067
rect 1253 9993 1267 10007
rect 1213 9973 1227 9987
rect 1153 9953 1167 9967
rect 1193 9953 1207 9967
rect 1073 9793 1087 9807
rect 1113 9793 1127 9807
rect 913 9753 927 9767
rect 873 9733 887 9747
rect 893 9693 907 9707
rect 853 9633 867 9647
rect 853 9473 867 9487
rect 953 9633 967 9647
rect 853 9433 867 9447
rect 973 9453 987 9467
rect 873 9353 887 9367
rect 933 9353 947 9367
rect 853 9293 867 9307
rect 613 8973 627 8987
rect 433 8953 447 8967
rect 773 9093 787 9107
rect 733 8893 747 8907
rect 713 8793 727 8807
rect 173 8733 187 8747
rect 193 8553 207 8567
rect 233 8553 247 8567
rect 273 8493 287 8507
rect 453 8493 467 8507
rect 493 8473 507 8487
rect 253 8413 267 8427
rect 473 8333 487 8347
rect 373 8313 387 8327
rect 33 8073 47 8087
rect 53 8073 67 8087
rect 393 8053 407 8067
rect 353 8013 367 8027
rect 233 7833 247 7847
rect 173 7813 187 7827
rect 213 7753 227 7767
rect 193 7513 207 7527
rect 93 7353 107 7367
rect 213 7353 227 7367
rect 53 7093 67 7107
rect 73 7073 87 7087
rect 193 7333 207 7347
rect 233 7313 247 7327
rect 293 7353 307 7367
rect 293 7313 307 7327
rect 273 7293 287 7307
rect 173 7073 187 7087
rect 93 7033 107 7047
rect 193 7033 207 7047
rect 253 6893 267 6907
rect 213 6853 227 6867
rect 193 6733 207 6747
rect 233 6413 247 6427
rect 273 6413 287 6427
rect 213 6373 227 6387
rect 253 6373 267 6387
rect 73 6233 87 6247
rect 233 6173 247 6187
rect 193 6113 207 6127
rect 253 6113 267 6127
rect 253 6073 267 6087
rect 213 6053 227 6067
rect 273 6053 287 6067
rect 33 5873 47 5887
rect 13 5013 27 5027
rect 13 4953 27 4967
rect 693 8773 707 8787
rect 673 8553 687 8567
rect 733 8773 747 8787
rect 693 8513 707 8527
rect 673 8413 687 8427
rect 633 8333 647 8347
rect 593 8313 607 8327
rect 633 8293 647 8307
rect 753 8293 767 8307
rect 673 8093 687 8107
rect 633 8033 647 8047
rect 953 9013 967 9027
rect 913 8993 927 9007
rect 893 8893 907 8907
rect 913 8793 927 8807
rect 933 8773 947 8787
rect 1093 9773 1107 9787
rect 1113 9753 1127 9767
rect 1153 9753 1167 9767
rect 1133 9733 1147 9747
rect 1173 9473 1187 9487
rect 1193 9413 1207 9427
rect 1133 9253 1147 9267
rect 1193 9253 1207 9267
rect 1113 9013 1127 9027
rect 1073 8993 1087 9007
rect 1033 8973 1047 8987
rect 1153 8973 1167 8987
rect 1153 8933 1167 8947
rect 1133 8813 1147 8827
rect 1233 9833 1247 9847
rect 1213 8913 1227 8927
rect 893 8753 907 8767
rect 953 8753 967 8767
rect 1133 8753 1147 8767
rect 953 8553 967 8567
rect 913 8513 927 8527
rect 1153 8533 1167 8547
rect 1173 8493 1187 8507
rect 1193 8493 1207 8507
rect 1133 8413 1147 8427
rect 873 8393 887 8407
rect 933 8393 947 8407
rect 973 8393 987 8407
rect 1093 8333 1107 8347
rect 1153 8333 1167 8347
rect 1053 8313 1067 8327
rect 1053 8293 1067 8307
rect 1193 8293 1207 8307
rect 1093 8273 1107 8287
rect 773 8093 787 8107
rect 833 8093 847 8107
rect 713 8073 727 8087
rect 493 8013 507 8027
rect 633 8013 647 8027
rect 413 7833 427 7847
rect 453 7813 467 7827
rect 433 7793 447 7807
rect 813 8053 827 8067
rect 673 7973 687 7987
rect 713 7973 727 7987
rect 633 7573 647 7587
rect 673 7573 687 7587
rect 493 7553 507 7567
rect 453 7333 467 7347
rect 413 7293 427 7307
rect 433 7293 447 7307
rect 393 7073 407 7087
rect 553 7533 567 7547
rect 533 7293 547 7307
rect 433 6873 447 6887
rect 493 7113 507 7127
rect 473 6893 487 6907
rect 513 7093 527 7107
rect 493 6873 507 6887
rect 453 6833 467 6847
rect 573 7333 587 7347
rect 553 7113 567 7127
rect 653 7553 667 7567
rect 693 7533 707 7547
rect 673 7513 687 7527
rect 713 7353 727 7367
rect 653 7333 667 7347
rect 693 7293 707 7307
rect 573 6973 587 6987
rect 613 6853 627 6867
rect 413 6593 427 6607
rect 373 6553 387 6567
rect 453 6413 467 6427
rect 473 6413 487 6427
rect 493 6393 507 6407
rect 393 6233 407 6247
rect 533 6133 547 6147
rect 453 6073 467 6087
rect 433 6053 447 6067
rect 373 5913 387 5927
rect 393 5913 407 5927
rect 353 5613 367 5627
rect 513 5893 527 5907
rect 453 5653 467 5667
rect 473 5653 487 5667
rect 213 5473 227 5487
rect 433 5473 447 5487
rect 273 5453 287 5467
rect 453 5453 467 5467
rect 193 5413 207 5427
rect 213 5153 227 5167
rect 173 5133 187 5147
rect 273 5413 287 5427
rect 393 5153 407 5167
rect 233 5033 247 5047
rect 213 4793 227 4807
rect 173 4673 187 4687
rect 233 4653 247 4667
rect 813 7093 827 7107
rect 673 7013 687 7027
rect 693 6973 707 6987
rect 673 6893 687 6907
rect 733 6873 747 6887
rect 713 6853 727 6867
rect 653 6833 667 6847
rect 613 6613 627 6627
rect 713 6653 727 6667
rect 673 6613 687 6627
rect 653 6593 667 6607
rect 633 6573 647 6587
rect 673 6413 687 6427
rect 813 6573 827 6587
rect 753 6413 767 6427
rect 693 6353 707 6367
rect 693 6133 707 6147
rect 673 6093 687 6107
rect 713 6093 727 6107
rect 793 6273 807 6287
rect 573 6073 587 6087
rect 653 6073 667 6087
rect 733 6073 747 6087
rect 773 6033 787 6047
rect 593 5913 607 5927
rect 573 5893 587 5907
rect 773 5893 787 5907
rect 633 5653 647 5667
rect 673 5653 687 5667
rect 553 5453 567 5467
rect 593 5453 607 5467
rect 533 5273 547 5287
rect 413 5113 427 5127
rect 413 5033 427 5047
rect 473 5153 487 5167
rect 513 5153 527 5167
rect 453 5133 467 5147
rect 493 5053 507 5067
rect 433 4953 447 4967
rect 473 4953 487 4967
rect 413 4793 427 4807
rect 473 4713 487 4727
rect 393 4693 407 4707
rect 353 4633 367 4647
rect 33 4433 47 4447
rect 53 4433 67 4447
rect 233 4193 247 4207
rect 193 4173 207 4187
rect 573 5113 587 5127
rect 533 5053 547 5067
rect 453 4673 467 4687
rect 513 4673 527 4687
rect 413 4653 427 4667
rect 493 4473 507 4487
rect 513 4473 527 4487
rect 453 4453 467 4467
rect 413 4413 427 4427
rect 393 4193 407 4207
rect 473 4173 487 4187
rect 553 4713 567 4727
rect 693 5413 707 5427
rect 873 8073 887 8087
rect 1013 8073 1027 8087
rect 913 8033 927 8047
rect 913 7813 927 7827
rect 893 7793 907 7807
rect 933 7733 947 7747
rect 953 7653 967 7667
rect 873 7553 887 7567
rect 853 7073 867 7087
rect 853 6953 867 6967
rect 1373 9913 1387 9927
rect 1493 9913 1507 9927
rect 1393 9893 1407 9907
rect 1353 9793 1367 9807
rect 1393 9793 1407 9807
rect 1353 9773 1367 9787
rect 1253 9733 1267 9747
rect 1413 9733 1427 9747
rect 1433 9733 1447 9747
rect 1373 9713 1387 9727
rect 1373 9493 1387 9507
rect 1333 9473 1347 9487
rect 1413 9473 1427 9487
rect 1313 9433 1327 9447
rect 1393 9453 1407 9467
rect 1373 9293 1387 9307
rect 1313 9213 1327 9227
rect 1273 8993 1287 9007
rect 1253 8773 1267 8787
rect 1233 8193 1247 8207
rect 1393 9253 1407 9267
rect 1353 9213 1367 9227
rect 1473 9713 1487 9727
rect 1453 9513 1467 9527
rect 1453 9473 1467 9487
rect 1473 9453 1487 9467
rect 1393 8993 1407 9007
rect 1433 8993 1447 9007
rect 1493 8993 1507 9007
rect 1373 8973 1387 8987
rect 1473 8953 1487 8967
rect 1413 8873 1427 8887
rect 1373 8793 1387 8807
rect 1313 8773 1327 8787
rect 1353 8773 1367 8787
rect 1393 8773 1407 8787
rect 1313 8753 1327 8767
rect 1273 8513 1287 8527
rect 1293 8033 1307 8047
rect 1253 8013 1267 8027
rect 1213 7973 1227 7987
rect 1033 7933 1047 7947
rect 1133 7933 1147 7947
rect 1353 8633 1367 8647
rect 1433 8513 1447 8527
rect 1413 8493 1427 8507
rect 1373 8393 1387 8407
rect 1333 8333 1347 8347
rect 1453 8313 1467 8327
rect 1473 8033 1487 8047
rect 1653 10853 1667 10867
rect 1713 10873 1727 10887
rect 1733 10793 1747 10807
rect 1653 10753 1667 10767
rect 1693 10753 1707 10767
rect 1633 10713 1647 10727
rect 1633 10473 1647 10487
rect 1573 10453 1587 10467
rect 1613 10453 1627 10467
rect 1593 10433 1607 10447
rect 1693 10713 1707 10727
rect 1733 10713 1747 10727
rect 1673 10693 1687 10707
rect 1713 10653 1727 10667
rect 1713 10473 1727 10487
rect 1653 10253 1667 10267
rect 1633 10213 1647 10227
rect 1613 9933 1627 9947
rect 1653 9933 1667 9947
rect 1713 9933 1727 9947
rect 1633 9913 1647 9927
rect 1613 9853 1627 9867
rect 1653 9773 1667 9787
rect 1633 9553 1647 9567
rect 1593 9493 1607 9507
rect 1673 9733 1687 9747
rect 1693 9713 1707 9727
rect 1653 9493 1667 9507
rect 1593 9473 1607 9487
rect 1633 9473 1647 9487
rect 1533 8973 1547 8987
rect 1653 9453 1667 9467
rect 1673 9453 1687 9467
rect 1613 9433 1627 9447
rect 1633 9433 1647 9447
rect 1613 9293 1627 9307
rect 1653 9293 1667 9307
rect 1653 8993 1667 9007
rect 1693 8993 1707 9007
rect 1633 8973 1647 8987
rect 1673 8933 1687 8947
rect 1613 8793 1627 8807
rect 1653 8793 1667 8807
rect 1773 10893 1787 10907
rect 1853 10713 1867 10727
rect 1793 10473 1807 10487
rect 2713 11213 2727 11227
rect 2673 11193 2687 11207
rect 1913 11173 1927 11187
rect 2193 11173 2207 11187
rect 2293 11173 2307 11187
rect 2453 11173 2467 11187
rect 2493 11173 2507 11187
rect 2693 11173 2707 11187
rect 2773 11193 2787 11207
rect 2233 11133 2247 11147
rect 1893 10913 1907 10927
rect 2053 10873 2067 10887
rect 1893 10853 1907 10867
rect 1913 10813 1927 10827
rect 2113 10913 2127 10927
rect 2153 10913 2167 10927
rect 2073 10833 2087 10847
rect 2093 10833 2107 10847
rect 1893 10713 1907 10727
rect 1873 10453 1887 10467
rect 1933 10453 1947 10467
rect 1853 10433 1867 10447
rect 1893 10433 1907 10447
rect 1833 10413 1847 10427
rect 1873 10413 1887 10427
rect 1913 10413 1927 10427
rect 1853 10393 1867 10407
rect 1893 10393 1907 10407
rect 1773 10253 1787 10267
rect 1873 10273 1887 10287
rect 1753 9773 1767 9787
rect 1733 9253 1747 9267
rect 1733 8973 1747 8987
rect 1693 8713 1707 8727
rect 1673 8593 1687 8607
rect 1593 8533 1607 8547
rect 1573 8513 1587 8527
rect 1653 8493 1667 8507
rect 1673 8453 1687 8467
rect 1573 8433 1587 8447
rect 1553 8413 1567 8427
rect 1653 8393 1667 8407
rect 1593 8373 1607 8387
rect 1533 8033 1547 8047
rect 1573 8033 1587 8047
rect 1313 7853 1327 7867
rect 1353 7853 1367 7867
rect 1433 7853 1447 7867
rect 1333 7833 1347 7847
rect 1393 7833 1407 7847
rect 1453 7833 1467 7847
rect 1073 7793 1087 7807
rect 1153 7813 1167 7827
rect 1073 7773 1087 7787
rect 1113 7773 1127 7787
rect 933 7553 947 7567
rect 973 7353 987 7367
rect 933 7313 947 7327
rect 893 7073 907 7087
rect 933 7073 947 7087
rect 953 7073 967 7087
rect 933 6973 947 6987
rect 893 6873 907 6887
rect 913 6853 927 6867
rect 1413 7813 1427 7827
rect 1373 7793 1387 7807
rect 1453 7793 1467 7807
rect 1333 7753 1347 7767
rect 1133 7373 1147 7387
rect 1313 7373 1327 7387
rect 1073 7333 1087 7347
rect 1113 7333 1127 7347
rect 1153 7333 1167 7347
rect 1053 7179 1067 7193
rect 973 6993 987 7007
rect 1093 6993 1107 7007
rect 873 6833 887 6847
rect 913 6833 927 6847
rect 933 6513 947 6527
rect 913 6493 927 6507
rect 973 6493 987 6507
rect 1033 6493 1047 6507
rect 933 6393 947 6407
rect 1013 6413 1027 6427
rect 953 6353 967 6367
rect 833 6253 847 6267
rect 1013 6353 1027 6367
rect 993 6153 1007 6167
rect 913 6113 927 6127
rect 953 6113 967 6127
rect 933 6033 947 6047
rect 953 6033 967 6047
rect 953 5933 967 5947
rect 893 5893 907 5907
rect 933 5873 947 5887
rect 853 5613 867 5627
rect 1013 5653 1027 5667
rect 933 5633 947 5647
rect 713 5393 727 5407
rect 793 5393 807 5407
rect 673 5353 687 5367
rect 633 5253 647 5267
rect 633 5073 647 5087
rect 633 4973 647 4987
rect 633 4953 647 4967
rect 693 5113 707 5127
rect 713 4953 727 4967
rect 833 4953 847 4967
rect 693 4933 707 4947
rect 773 4933 787 4947
rect 673 4913 687 4927
rect 593 4653 607 4667
rect 553 4453 567 4467
rect 653 4853 667 4867
rect 753 4713 767 4727
rect 713 4593 727 4607
rect 673 4473 687 4487
rect 693 4473 707 4487
rect 733 4453 747 4467
rect 713 4433 727 4447
rect 653 4233 667 4247
rect 353 4133 367 4147
rect 253 4113 267 4127
rect 393 4113 407 4127
rect 233 3773 247 3787
rect 193 3713 207 3727
rect 253 3713 267 3727
rect 253 3673 267 3687
rect 213 3653 227 3667
rect 713 4213 727 4227
rect 813 4913 827 4927
rect 913 5513 927 5527
rect 1013 5513 1027 5527
rect 913 5453 927 5467
rect 893 5433 907 5447
rect 953 5433 967 5447
rect 873 5153 887 5167
rect 853 4893 867 4907
rect 853 4713 867 4727
rect 973 5413 987 5427
rect 933 5393 947 5407
rect 953 5353 967 5367
rect 1013 5273 1027 5287
rect 993 5253 1007 5267
rect 893 5113 907 5127
rect 993 5053 1007 5067
rect 953 4973 967 4987
rect 933 4933 947 4947
rect 1193 7293 1207 7307
rect 1133 7179 1147 7193
rect 1273 7173 1287 7187
rect 1253 7093 1267 7107
rect 1133 7033 1147 7047
rect 1193 7073 1207 7087
rect 1233 7073 1247 7087
rect 1213 7053 1227 7067
rect 1173 7013 1187 7027
rect 1153 6973 1167 6987
rect 1193 6933 1207 6947
rect 1113 6913 1127 6927
rect 1113 6873 1127 6887
rect 1173 6873 1187 6887
rect 1153 6853 1167 6867
rect 1273 7053 1287 7067
rect 1233 6853 1247 6867
rect 1113 6553 1127 6567
rect 1193 6593 1207 6607
rect 1253 6593 1267 6607
rect 1153 6493 1167 6507
rect 1133 6393 1147 6407
rect 1193 6393 1207 6407
rect 1233 6393 1247 6407
rect 1093 6373 1107 6387
rect 1093 5913 1107 5927
rect 1173 6233 1187 6247
rect 1213 6233 1227 6247
rect 1233 6153 1247 6167
rect 1173 6133 1187 6147
rect 1153 6093 1167 6107
rect 1193 6093 1207 6107
rect 1173 5913 1187 5927
rect 1293 7033 1307 7047
rect 1553 8013 1567 8027
rect 1653 8013 1667 8027
rect 1473 7733 1487 7747
rect 1473 7553 1487 7567
rect 1433 7373 1447 7387
rect 1453 7373 1467 7387
rect 1393 7353 1407 7367
rect 1493 7353 1507 7367
rect 1373 7333 1387 7347
rect 1353 7293 1367 7307
rect 1393 7293 1407 7307
rect 1333 7173 1347 7187
rect 1573 7993 1587 8007
rect 1653 7853 1667 7867
rect 1673 7833 1687 7847
rect 1613 7793 1627 7807
rect 1633 7573 1647 7587
rect 1613 7553 1627 7567
rect 1653 7553 1667 7567
rect 1653 7533 1667 7547
rect 1633 7333 1647 7347
rect 1613 7313 1627 7327
rect 1513 7293 1527 7307
rect 1493 7173 1507 7187
rect 1393 6953 1407 6967
rect 1413 6873 1427 6887
rect 1593 6953 1607 6967
rect 1513 6913 1527 6927
rect 1473 6873 1487 6887
rect 1453 6853 1467 6867
rect 1453 6673 1467 6687
rect 1373 6613 1387 6627
rect 1453 6613 1467 6627
rect 1313 6573 1327 6587
rect 1413 6593 1427 6607
rect 1393 6553 1407 6567
rect 1473 6573 1487 6587
rect 1433 6533 1447 6547
rect 1473 6513 1487 6527
rect 1393 6413 1407 6427
rect 1453 6393 1467 6407
rect 1533 6873 1547 6887
rect 1573 6873 1587 6887
rect 1513 6473 1527 6487
rect 1373 6353 1387 6367
rect 1273 6173 1287 6187
rect 1273 6133 1287 6147
rect 1353 6133 1367 6147
rect 1273 5893 1287 5907
rect 1573 6533 1587 6547
rect 1533 6333 1547 6347
rect 1533 6153 1547 6167
rect 1433 6113 1447 6127
rect 1493 6113 1507 6127
rect 1513 6113 1527 6127
rect 1633 7173 1647 7187
rect 1613 6733 1627 6747
rect 1653 6933 1667 6947
rect 1753 8753 1767 8767
rect 1753 8533 1767 8547
rect 1733 8453 1747 8467
rect 1813 10213 1827 10227
rect 1793 9933 1807 9947
rect 1873 9993 1887 10007
rect 1893 9933 1907 9947
rect 1873 9913 1887 9927
rect 1913 9913 1927 9927
rect 1853 9873 1867 9887
rect 1833 9853 1847 9867
rect 1813 9753 1827 9767
rect 1913 9753 1927 9767
rect 1893 9713 1907 9727
rect 2053 10713 2067 10727
rect 1993 10593 2007 10607
rect 1953 10413 1967 10427
rect 1973 9833 1987 9847
rect 2073 10353 2087 10367
rect 2053 10193 2067 10207
rect 2073 10053 2087 10067
rect 2213 10873 2227 10887
rect 2413 10913 2427 10927
rect 2453 10913 2467 10927
rect 2373 10873 2387 10887
rect 2233 10833 2247 10847
rect 2213 10753 2227 10767
rect 2153 10733 2167 10747
rect 2133 10713 2147 10727
rect 2113 10353 2127 10367
rect 2293 10453 2307 10467
rect 2253 10433 2267 10447
rect 2333 10433 2347 10447
rect 2313 10413 2327 10427
rect 2273 10373 2287 10387
rect 2273 10353 2287 10367
rect 2193 10273 2207 10287
rect 2093 10013 2107 10027
rect 2113 9973 2127 9987
rect 2093 9953 2107 9967
rect 2033 9933 2047 9947
rect 2133 9933 2147 9947
rect 2113 9773 2127 9787
rect 1993 9753 2007 9767
rect 1973 9733 1987 9747
rect 2253 9513 2267 9527
rect 1873 9493 1887 9507
rect 2153 9493 2167 9507
rect 1913 9473 1927 9487
rect 1973 9473 1987 9487
rect 2193 9473 2207 9487
rect 2233 9473 2247 9487
rect 1833 9433 1847 9447
rect 1813 9333 1827 9347
rect 1793 9113 1807 9127
rect 1893 9453 1907 9467
rect 1933 9433 1947 9447
rect 1853 9333 1867 9347
rect 1873 9293 1887 9307
rect 1893 9253 1907 9267
rect 1833 9113 1847 9127
rect 1853 9113 1867 9127
rect 1913 9113 1927 9127
rect 1813 9093 1827 9107
rect 1853 9093 1867 9107
rect 1893 9013 1907 9027
rect 1893 8813 1907 8827
rect 1873 8793 1887 8807
rect 1933 8953 1947 8967
rect 2073 9453 2087 9467
rect 2133 9453 2147 9467
rect 2173 9453 2187 9467
rect 2213 9433 2227 9447
rect 2073 9413 2087 9427
rect 2113 9253 2127 9267
rect 2193 9253 2207 9267
rect 2133 9013 2147 9027
rect 2153 8993 2167 9007
rect 2093 8973 2107 8987
rect 2193 8933 2207 8947
rect 2133 8833 2147 8847
rect 2153 8833 2167 8847
rect 2113 8793 2127 8807
rect 1973 8773 1987 8787
rect 2173 8773 2187 8787
rect 1853 8753 1867 8767
rect 1913 8753 1927 8767
rect 2073 8573 2087 8587
rect 1833 8533 1847 8547
rect 1933 8533 1947 8547
rect 1773 8453 1787 8467
rect 1753 8393 1767 8407
rect 1773 8333 1787 8347
rect 1793 8333 1807 8347
rect 1913 8493 1927 8507
rect 1973 8473 1987 8487
rect 2253 9453 2267 9467
rect 2233 8993 2247 9007
rect 2173 8653 2187 8667
rect 2173 8473 2187 8487
rect 2193 8433 2207 8447
rect 2153 8353 2167 8367
rect 2073 8333 2087 8347
rect 1873 8313 1887 8327
rect 1933 8313 1947 8327
rect 2113 8313 2127 8327
rect 1773 8293 1787 8307
rect 1813 8273 1827 8287
rect 1853 8273 1867 8287
rect 1813 8053 1827 8067
rect 1853 8033 1867 8047
rect 1733 8013 1747 8027
rect 1773 7993 1787 8007
rect 1773 7973 1787 7987
rect 1753 7793 1767 7807
rect 1733 7553 1747 7567
rect 1753 7493 1767 7507
rect 1733 7073 1747 7087
rect 1733 6973 1747 6987
rect 1713 6953 1727 6967
rect 1653 6893 1667 6907
rect 1693 6893 1707 6907
rect 1693 6873 1707 6887
rect 1673 6853 1687 6867
rect 1833 7853 1847 7867
rect 1793 7573 1807 7587
rect 1873 7853 1887 7867
rect 1893 7833 1907 7847
rect 2093 8293 2107 8307
rect 2133 8293 2147 8307
rect 2133 8273 2147 8287
rect 2013 8033 2027 8047
rect 1933 7773 1947 7787
rect 1833 7553 1847 7567
rect 1893 7553 1907 7567
rect 1933 7553 1947 7567
rect 1973 7553 1987 7567
rect 1813 7353 1827 7367
rect 1873 7353 1887 7367
rect 1793 7093 1807 7107
rect 1853 7333 1867 7347
rect 1893 7313 1907 7327
rect 1973 7513 1987 7527
rect 1953 7493 1967 7507
rect 2253 8833 2267 8847
rect 3373 11213 3387 11227
rect 3453 11213 3467 11227
rect 4133 11293 4147 11307
rect 4173 11293 4187 11307
rect 4333 11293 4347 11307
rect 4373 11293 4387 11307
rect 2793 11153 2807 11167
rect 2833 10933 2847 10947
rect 2913 10933 2927 10947
rect 2793 10913 2807 10927
rect 2653 10873 2667 10887
rect 2593 10853 2607 10867
rect 2633 10853 2647 10867
rect 2453 10733 2467 10747
rect 2473 10693 2487 10707
rect 2433 10673 2447 10687
rect 2533 10673 2547 10687
rect 2413 10513 2427 10527
rect 2513 10453 2527 10467
rect 2393 10413 2407 10427
rect 2553 10433 2567 10447
rect 2773 10893 2787 10907
rect 2733 10853 2747 10867
rect 2713 10733 2727 10747
rect 2753 10753 2767 10767
rect 2673 10693 2687 10707
rect 2613 10493 2627 10507
rect 2613 10453 2627 10467
rect 2573 10393 2587 10407
rect 2293 10253 2307 10267
rect 2333 10253 2347 10267
rect 2533 10253 2547 10267
rect 2573 10253 2587 10267
rect 2333 10233 2347 10247
rect 2373 10233 2387 10247
rect 2353 10213 2367 10227
rect 2313 10193 2327 10207
rect 2293 10013 2307 10027
rect 2373 10053 2387 10067
rect 2313 9993 2327 10007
rect 2353 9973 2367 9987
rect 2313 9953 2327 9967
rect 2353 9953 2367 9967
rect 2393 9953 2407 9967
rect 2373 9853 2387 9867
rect 2333 9773 2347 9787
rect 2373 9733 2387 9747
rect 2393 9633 2407 9647
rect 2413 9493 2427 9507
rect 2393 9473 2407 9487
rect 2433 9473 2447 9487
rect 2473 9473 2487 9487
rect 2513 9473 2527 9487
rect 2453 9453 2467 9467
rect 2413 9413 2427 9427
rect 2493 9413 2507 9427
rect 2393 9313 2407 9327
rect 2353 9273 2367 9287
rect 2373 9253 2387 9267
rect 2293 9193 2307 9207
rect 2273 8713 2287 8727
rect 2273 8653 2287 8667
rect 2253 8293 2267 8307
rect 2233 8233 2247 8247
rect 2213 8013 2227 8027
rect 2253 8013 2267 8027
rect 2173 7973 2187 7987
rect 2073 7873 2087 7887
rect 2353 9013 2367 9027
rect 2413 9273 2427 9287
rect 2433 9173 2447 9187
rect 2493 9013 2507 9027
rect 2373 8993 2387 9007
rect 2373 8913 2387 8927
rect 2413 8793 2427 8807
rect 2473 8793 2487 8807
rect 2353 8773 2367 8787
rect 2453 8773 2467 8787
rect 2393 8733 2407 8747
rect 2393 8633 2407 8647
rect 2433 8573 2447 8587
rect 2353 8393 2367 8407
rect 2293 8373 2307 8387
rect 2433 8353 2447 8367
rect 2353 8333 2367 8347
rect 2333 8293 2347 8307
rect 2313 8053 2327 8067
rect 2293 8013 2307 8027
rect 2313 8013 2327 8027
rect 2273 7873 2287 7887
rect 2493 8313 2507 8327
rect 2473 8153 2487 8167
rect 2553 10213 2567 10227
rect 2673 10393 2687 10407
rect 2873 10913 2887 10927
rect 3113 11133 3127 11147
rect 3153 11113 3167 11127
rect 3153 10933 3167 10947
rect 3093 10913 3107 10927
rect 3133 10913 3147 10927
rect 2853 10893 2867 10907
rect 2893 10893 2907 10907
rect 2833 10873 2847 10887
rect 2853 10853 2867 10867
rect 2953 10893 2967 10907
rect 3093 10873 3107 10887
rect 2933 10833 2947 10847
rect 3153 10893 3167 10907
rect 3193 10913 3207 10927
rect 3193 10873 3207 10887
rect 3173 10853 3187 10867
rect 3213 10853 3227 10867
rect 3193 10833 3207 10847
rect 3113 10753 3127 10767
rect 3093 10733 3107 10747
rect 2913 10713 2927 10727
rect 2813 10693 2827 10707
rect 2953 10693 2967 10707
rect 2913 10673 2927 10687
rect 2933 10673 2947 10687
rect 2973 10673 2987 10687
rect 2773 10333 2787 10347
rect 2913 10413 2927 10427
rect 2833 10313 2847 10327
rect 2833 10293 2847 10307
rect 2733 10273 2747 10287
rect 2793 10233 2807 10247
rect 3233 10593 3247 10607
rect 3193 10573 3207 10587
rect 3113 10553 3127 10567
rect 3033 10433 3047 10447
rect 3073 10433 3087 10447
rect 3113 10433 3127 10447
rect 3153 10433 3167 10447
rect 3013 10393 3027 10407
rect 3053 10413 3067 10427
rect 2993 10333 3007 10347
rect 2733 10153 2747 10167
rect 2733 9953 2747 9967
rect 2633 9853 2647 9867
rect 2613 9713 2627 9727
rect 2653 9753 2667 9767
rect 2653 9713 2667 9727
rect 2673 9553 2687 9567
rect 2633 9533 2647 9547
rect 2573 9453 2587 9467
rect 2713 9453 2727 9467
rect 2913 10213 2927 10227
rect 2813 10193 2827 10207
rect 2793 9953 2807 9967
rect 2813 9953 2827 9967
rect 2653 9393 2667 9407
rect 2573 9293 2587 9307
rect 2613 9293 2627 9307
rect 2533 9273 2547 9287
rect 2573 9253 2587 9267
rect 2593 9253 2607 9267
rect 2573 8993 2587 9007
rect 2553 8853 2567 8867
rect 2553 8773 2567 8787
rect 2673 9253 2687 9267
rect 2673 9233 2687 9247
rect 2653 8993 2667 9007
rect 2613 8973 2627 8987
rect 2593 8853 2607 8867
rect 2573 8753 2587 8767
rect 2633 8753 2647 8767
rect 2573 8713 2587 8727
rect 2513 8293 2527 8307
rect 2613 8553 2627 8567
rect 2593 8433 2607 8447
rect 2633 8393 2647 8407
rect 2593 8373 2607 8387
rect 2613 8293 2627 8307
rect 2233 7853 2247 7867
rect 2313 7833 2327 7847
rect 2113 7813 2127 7827
rect 2213 7813 2227 7827
rect 2333 7813 2347 7827
rect 2033 7793 2047 7807
rect 2093 7533 2107 7547
rect 2133 7533 2147 7547
rect 2153 7513 2167 7527
rect 2173 7513 2187 7527
rect 2113 7453 2127 7467
rect 2073 7353 2087 7367
rect 1993 7333 2007 7347
rect 2193 7353 2207 7367
rect 2113 7293 2127 7307
rect 2113 7173 2127 7187
rect 1913 7133 1927 7147
rect 1833 7113 1847 7127
rect 1913 7113 1927 7127
rect 1813 6633 1827 6647
rect 1713 6613 1727 6627
rect 1773 6613 1787 6627
rect 1753 6593 1767 6607
rect 1793 6593 1807 6607
rect 1733 6573 1747 6587
rect 1773 6553 1787 6567
rect 1693 6453 1707 6467
rect 1753 6453 1767 6467
rect 1713 6433 1727 6447
rect 1733 6413 1747 6427
rect 1633 6393 1647 6407
rect 1713 6393 1727 6407
rect 1473 6093 1487 6107
rect 1453 6073 1467 6087
rect 1373 5933 1387 5947
rect 1193 5873 1207 5887
rect 1213 5873 1227 5887
rect 1353 5873 1367 5887
rect 1573 5973 1587 5987
rect 1553 5953 1567 5967
rect 1513 5853 1527 5867
rect 1553 5853 1567 5867
rect 1233 5633 1247 5647
rect 1533 5633 1547 5647
rect 1093 5573 1107 5587
rect 1153 5573 1167 5587
rect 1333 5573 1347 5587
rect 1213 5453 1227 5467
rect 1173 5413 1187 5427
rect 1213 5373 1227 5387
rect 1153 5353 1167 5367
rect 1113 5253 1127 5267
rect 973 4913 987 4927
rect 1033 4913 1047 4927
rect 1173 5113 1187 5127
rect 1313 5073 1327 5087
rect 1253 5053 1267 5067
rect 1253 5033 1267 5047
rect 1193 4973 1207 4987
rect 1133 4953 1147 4967
rect 933 4813 947 4827
rect 1053 4813 1067 4827
rect 1213 4953 1227 4967
rect 853 4633 867 4647
rect 873 4633 887 4647
rect 1033 4633 1047 4647
rect 1133 4633 1147 4647
rect 1213 4613 1227 4627
rect 853 4593 867 4607
rect 1053 4493 1067 4507
rect 1213 4493 1227 4507
rect 913 4473 927 4487
rect 833 4393 847 4407
rect 813 4373 827 4387
rect 693 4153 707 4167
rect 653 4033 667 4047
rect 613 4013 627 4027
rect 493 3993 507 4007
rect 453 3973 467 3987
rect 473 3973 487 3987
rect 393 3773 407 3787
rect 593 3753 607 3767
rect 533 3713 547 3727
rect 413 3693 427 3707
rect 493 3693 507 3707
rect 433 3673 447 3687
rect 453 3673 467 3687
rect 453 3653 467 3667
rect 413 3493 427 3507
rect 453 3493 467 3507
rect 373 3453 387 3467
rect 313 3373 327 3387
rect 353 3373 367 3387
rect 173 3293 187 3307
rect 173 3253 187 3267
rect 213 3233 227 3247
rect 273 3013 287 3027
rect 233 2993 247 3007
rect 233 2773 247 2787
rect 193 2753 207 2767
rect 213 2713 227 2727
rect 213 2573 227 2587
rect 413 3233 427 3247
rect 533 3233 547 3247
rect 573 3233 587 3247
rect 393 3213 407 3227
rect 513 3213 527 3227
rect 553 3213 567 3227
rect 473 3173 487 3187
rect 433 3053 447 3067
rect 393 3013 407 3027
rect 413 3013 427 3027
rect 413 2993 427 3007
rect 453 2953 467 2967
rect 413 2773 427 2787
rect 433 2753 447 2767
rect 633 3953 647 3967
rect 673 3953 687 3967
rect 713 3953 727 3967
rect 693 3733 707 3747
rect 813 4153 827 4167
rect 893 4433 907 4447
rect 953 4433 967 4447
rect 933 4413 947 4427
rect 913 4233 927 4247
rect 933 4233 947 4247
rect 1353 5533 1367 5547
rect 1413 5533 1427 5547
rect 1453 5473 1467 5487
rect 1453 5453 1467 5467
rect 1433 5413 1447 5427
rect 1473 5393 1487 5407
rect 1353 5153 1367 5167
rect 1533 5153 1547 5167
rect 1453 5133 1467 5147
rect 1493 5113 1507 5127
rect 1353 5093 1367 5107
rect 1413 4973 1427 4987
rect 1453 4973 1467 4987
rect 1413 4953 1427 4967
rect 1513 4973 1527 4987
rect 1333 4653 1347 4667
rect 1393 4653 1407 4667
rect 1373 4493 1387 4507
rect 1313 4473 1327 4487
rect 1393 4473 1407 4487
rect 1473 4933 1487 4947
rect 1513 4933 1527 4947
rect 1433 4913 1447 4927
rect 1433 4653 1447 4667
rect 1433 4493 1447 4507
rect 1133 4453 1147 4467
rect 1233 4453 1247 4467
rect 1113 4433 1127 4447
rect 1153 4393 1167 4407
rect 1133 4233 1147 4247
rect 993 4213 1007 4227
rect 1053 4213 1067 4227
rect 933 4193 947 4207
rect 873 4173 887 4187
rect 1033 4173 1047 4187
rect 853 4053 867 4067
rect 993 4033 1007 4047
rect 913 3993 927 4007
rect 953 3993 967 4007
rect 1013 3993 1027 4007
rect 853 3953 867 3967
rect 733 3753 747 3767
rect 793 3733 807 3747
rect 673 3693 687 3707
rect 713 3693 727 3707
rect 653 3653 667 3667
rect 713 3653 727 3667
rect 773 3513 787 3527
rect 733 3493 747 3507
rect 793 3493 807 3507
rect 653 3233 667 3247
rect 633 3213 647 3227
rect 613 3053 627 3067
rect 633 3033 647 3047
rect 693 3213 707 3227
rect 653 3013 667 3027
rect 733 3253 747 3267
rect 713 3193 727 3207
rect 713 3033 727 3047
rect 693 2973 707 2987
rect 653 2773 667 2787
rect 613 2753 627 2767
rect 593 2713 607 2727
rect 593 2593 607 2607
rect 613 2593 627 2607
rect 393 2573 407 2587
rect 413 2573 427 2587
rect 193 2533 207 2547
rect 273 2533 287 2547
rect 293 2533 307 2547
rect 33 2513 47 2527
rect 173 2513 187 2527
rect 253 2513 267 2527
rect 273 2353 287 2367
rect 353 2353 367 2367
rect 93 2233 107 2247
rect 193 2233 207 2247
rect 73 2213 87 2227
rect 73 2073 87 2087
rect 73 1793 87 1807
rect 153 1713 167 1727
rect 93 1693 107 1707
rect 133 1553 147 1567
rect 193 1713 207 1727
rect 213 1693 227 1707
rect 193 1553 207 1567
rect 233 1553 247 1567
rect 253 1353 267 1367
rect 173 1333 187 1347
rect 193 1333 207 1347
rect 233 1313 247 1327
rect 213 1293 227 1307
rect 173 1273 187 1287
rect 153 1253 167 1267
rect 213 1253 227 1267
rect 373 2253 387 2267
rect 573 2533 587 2547
rect 553 2433 567 2447
rect 453 2273 467 2287
rect 493 2073 507 2087
rect 413 2053 427 2067
rect 453 2053 467 2067
rect 513 2053 527 2067
rect 493 1793 507 1807
rect 533 1693 547 1707
rect 413 1573 427 1587
rect 413 1353 427 1367
rect 393 1333 407 1347
rect 353 1273 367 1287
rect 433 1313 447 1327
rect 473 1293 487 1307
rect 473 1153 487 1167
rect 513 1113 527 1127
rect 133 813 147 827
rect 233 1093 247 1107
rect 393 1093 407 1107
rect 413 1093 427 1107
rect 453 1093 467 1107
rect 273 893 287 907
rect 193 833 207 847
rect 233 833 247 847
rect 173 733 187 747
rect 213 813 227 827
rect 233 633 247 647
rect 213 613 227 627
rect 253 613 267 627
rect 213 373 227 387
rect 233 353 247 367
rect 213 333 227 347
rect 493 1073 507 1087
rect 413 853 427 867
rect 473 813 487 827
rect 433 733 447 747
rect 433 713 447 727
rect 593 2293 607 2307
rect 613 2253 627 2267
rect 593 2073 607 2087
rect 673 2753 687 2767
rect 693 2573 707 2587
rect 653 2553 667 2567
rect 673 2493 687 2507
rect 673 2473 687 2487
rect 673 2293 687 2307
rect 653 2273 667 2287
rect 773 3313 787 3327
rect 773 3233 787 3247
rect 973 3973 987 3987
rect 933 3893 947 3907
rect 973 3893 987 3907
rect 913 3713 927 3727
rect 933 3693 947 3707
rect 953 3653 967 3667
rect 933 3513 947 3527
rect 1013 3673 1027 3687
rect 1013 3653 1027 3667
rect 1153 4153 1167 4167
rect 1173 4093 1187 4107
rect 1233 4073 1247 4087
rect 1353 4433 1367 4447
rect 1333 4133 1347 4147
rect 1233 3993 1247 4007
rect 1253 3993 1267 4007
rect 1313 3993 1327 4007
rect 1213 3953 1227 3967
rect 1153 3893 1167 3907
rect 1173 3773 1187 3787
rect 1173 3753 1187 3767
rect 1133 3733 1147 3747
rect 1113 3713 1127 3727
rect 1213 3713 1227 3727
rect 1113 3673 1127 3687
rect 1253 3693 1267 3707
rect 1413 4213 1427 4227
rect 1393 4153 1407 4167
rect 1873 7093 1887 7107
rect 1853 6873 1867 6887
rect 1833 6573 1847 6587
rect 1813 6553 1827 6567
rect 1793 6113 1807 6127
rect 1793 6073 1807 6087
rect 1893 7073 1907 7087
rect 2153 7073 2167 7087
rect 2133 7033 2147 7047
rect 2173 6993 2187 7007
rect 2153 6893 2167 6907
rect 2473 7793 2487 7807
rect 2453 7773 2467 7787
rect 2293 7673 2307 7687
rect 2273 7333 2287 7347
rect 2393 7533 2407 7547
rect 2413 7513 2427 7527
rect 2373 7493 2387 7507
rect 2333 7333 2347 7347
rect 2393 7453 2407 7467
rect 2293 7313 2307 7327
rect 2353 7313 2367 7327
rect 2373 7313 2387 7327
rect 2273 7073 2287 7087
rect 2413 7073 2427 7087
rect 2213 7033 2227 7047
rect 2293 6873 2307 6887
rect 1933 6853 1947 6867
rect 2173 6853 2187 6867
rect 2193 6853 2207 6867
rect 2393 7033 2407 7047
rect 2473 7533 2487 7547
rect 2653 8273 2667 8287
rect 2573 7853 2587 7867
rect 2633 7553 2647 7567
rect 2613 7453 2627 7467
rect 2573 7373 2587 7387
rect 2813 9853 2827 9867
rect 2813 9833 2827 9847
rect 2853 9833 2867 9847
rect 2853 9753 2867 9767
rect 2893 9753 2907 9767
rect 2793 9713 2807 9727
rect 2873 9713 2887 9727
rect 2833 9593 2847 9607
rect 2793 9493 2807 9507
rect 2793 9433 2807 9447
rect 2773 8893 2787 8907
rect 2753 8533 2767 8547
rect 2973 9953 2987 9967
rect 3093 10393 3107 10407
rect 3133 10393 3147 10407
rect 3093 10253 3107 10267
rect 3033 10213 3047 10227
rect 3073 10213 3087 10227
rect 3073 10153 3087 10167
rect 3033 9953 3047 9967
rect 3073 9953 3087 9967
rect 3053 9933 3067 9947
rect 2993 9913 3007 9927
rect 2973 9653 2987 9667
rect 2913 9393 2927 9407
rect 2853 9293 2867 9307
rect 2813 9253 2827 9267
rect 2893 9253 2907 9267
rect 2913 9233 2927 9247
rect 2873 9213 2887 9227
rect 2813 9033 2827 9047
rect 2833 9013 2847 9027
rect 2953 9433 2967 9447
rect 2953 9373 2967 9387
rect 2933 9193 2947 9207
rect 2913 9093 2927 9107
rect 2853 8993 2867 9007
rect 2813 8973 2827 8987
rect 2913 8833 2927 8847
rect 2813 8793 2827 8807
rect 2873 8793 2887 8807
rect 3013 9753 3027 9767
rect 3033 9733 3047 9747
rect 3053 9733 3067 9747
rect 3033 9653 3047 9667
rect 3013 9373 3027 9387
rect 3013 9273 3027 9287
rect 2993 9213 3007 9227
rect 2993 9013 3007 9027
rect 2813 8493 2827 8507
rect 2813 8453 2827 8467
rect 2853 8453 2867 8467
rect 2893 8353 2907 8367
rect 2993 8773 3007 8787
rect 2953 8593 2967 8607
rect 2833 8313 2847 8327
rect 2853 8293 2867 8307
rect 2813 8193 2827 8207
rect 2793 8093 2807 8107
rect 2713 8033 2727 8047
rect 2753 8033 2767 8047
rect 2773 8033 2787 8047
rect 2893 8273 2907 8287
rect 2853 8073 2867 8087
rect 2733 8013 2747 8027
rect 2813 8013 2827 8027
rect 2793 7993 2807 8007
rect 2893 7993 2907 8007
rect 2773 7973 2787 7987
rect 2773 7873 2787 7887
rect 2713 7853 2727 7867
rect 2753 7553 2767 7567
rect 2833 7833 2847 7847
rect 2933 7833 2947 7847
rect 2913 7753 2927 7767
rect 2773 7493 2787 7507
rect 2753 7333 2767 7347
rect 2893 7553 2907 7567
rect 2873 7533 2887 7547
rect 2853 7453 2867 7467
rect 2793 7373 2807 7387
rect 2833 7373 2847 7387
rect 2913 7353 2927 7367
rect 2813 7333 2827 7347
rect 2553 7313 2567 7327
rect 2673 7313 2687 7327
rect 2813 7313 2827 7327
rect 2513 7293 2527 7307
rect 2613 7073 2627 7087
rect 2653 7073 2667 7087
rect 2633 7053 2647 7067
rect 2733 7073 2747 7087
rect 2433 6893 2447 6907
rect 2713 7033 2727 7047
rect 2673 7013 2687 7027
rect 2733 7013 2747 7027
rect 2353 6853 2367 6867
rect 2393 6853 2407 6867
rect 2573 6853 2587 6867
rect 2613 6853 2627 6867
rect 2653 6853 2667 6867
rect 2713 6853 2727 6867
rect 2293 6833 2307 6847
rect 2373 6833 2387 6847
rect 1953 6733 1967 6747
rect 2093 6733 2107 6747
rect 1913 6633 1927 6647
rect 1893 6593 1907 6607
rect 1853 6353 1867 6367
rect 1633 6013 1647 6027
rect 1673 6013 1687 6027
rect 1753 6013 1767 6027
rect 1813 6013 1827 6027
rect 1633 5793 1647 5807
rect 1653 5653 1667 5667
rect 1593 5633 1607 5647
rect 1653 5633 1667 5647
rect 1613 5453 1627 5467
rect 1633 5453 1647 5467
rect 1613 5433 1627 5447
rect 1573 5393 1587 5407
rect 1633 5413 1647 5427
rect 1693 5453 1707 5467
rect 2053 6493 2067 6507
rect 2073 6493 2087 6507
rect 2013 6453 2027 6467
rect 1953 6433 1967 6447
rect 1913 6413 1927 6427
rect 1993 6393 2007 6407
rect 1913 6373 1927 6387
rect 1973 6373 1987 6387
rect 1973 6353 1987 6367
rect 1933 6333 1947 6347
rect 1953 6133 1967 6147
rect 1893 5993 1907 6007
rect 1833 5973 1847 5987
rect 1873 5933 1887 5947
rect 1893 5913 1907 5927
rect 1853 5853 1867 5867
rect 1933 5993 1947 6007
rect 1813 5793 1827 5807
rect 1853 5633 1867 5647
rect 1833 5613 1847 5627
rect 1753 5553 1767 5567
rect 1793 5553 1807 5567
rect 1673 5433 1687 5447
rect 1713 5433 1727 5447
rect 1673 5153 1687 5167
rect 1713 5153 1727 5167
rect 1653 5133 1667 5147
rect 1693 5133 1707 5147
rect 1873 5433 1887 5447
rect 1853 5413 1867 5427
rect 1833 5393 1847 5407
rect 1793 5153 1807 5167
rect 1613 4953 1627 4967
rect 1693 4973 1707 4987
rect 1713 4953 1727 4967
rect 1693 4933 1707 4947
rect 1573 4713 1587 4727
rect 1553 4693 1567 4707
rect 1633 4673 1647 4687
rect 1673 4673 1687 4687
rect 1613 4653 1627 4667
rect 1653 4653 1667 4667
rect 1513 4093 1527 4107
rect 1433 4073 1447 4087
rect 1453 4053 1467 4067
rect 1413 3973 1427 3987
rect 1433 3973 1447 3987
rect 1353 3953 1367 3967
rect 1473 3993 1487 4007
rect 1493 3953 1507 3967
rect 1433 3933 1447 3947
rect 1413 3913 1427 3927
rect 1593 4473 1607 4487
rect 1613 4473 1627 4487
rect 1573 4453 1587 4467
rect 1633 4393 1647 4407
rect 1593 4213 1607 4227
rect 1773 5013 1787 5027
rect 1773 4953 1787 4967
rect 1733 4853 1747 4867
rect 1753 4853 1767 4867
rect 1693 4053 1707 4067
rect 1653 3993 1667 4007
rect 1713 3993 1727 4007
rect 1613 3953 1627 3967
rect 1673 3973 1687 3987
rect 1693 3953 1707 3967
rect 1933 5633 1947 5647
rect 2073 6393 2087 6407
rect 2053 6373 2067 6387
rect 2053 6113 2067 6127
rect 1993 6093 2007 6107
rect 2213 6633 2227 6647
rect 2233 6613 2247 6627
rect 2413 6753 2427 6767
rect 2313 6673 2327 6687
rect 2233 6393 2247 6407
rect 2253 6373 2267 6387
rect 2253 6213 2267 6227
rect 2093 6173 2107 6187
rect 2093 6093 2107 6107
rect 2073 6073 2087 6087
rect 2273 6073 2287 6087
rect 1993 5953 2007 5967
rect 2053 5953 2067 5967
rect 2373 6593 2387 6607
rect 2313 6373 2327 6387
rect 2493 6493 2507 6507
rect 2553 6493 2567 6507
rect 2473 6393 2487 6407
rect 2533 6473 2547 6487
rect 2653 6753 2667 6767
rect 2713 6613 2727 6627
rect 2673 6593 2687 6607
rect 2753 6493 2767 6507
rect 2633 6393 2647 6407
rect 2653 6393 2667 6407
rect 2713 6393 2727 6407
rect 2513 6373 2527 6387
rect 2573 6373 2587 6387
rect 2433 6133 2447 6147
rect 2473 6173 2487 6187
rect 2393 6113 2407 6127
rect 2453 6113 2467 6127
rect 2373 6093 2387 6107
rect 2453 6073 2467 6087
rect 2373 5953 2387 5967
rect 2153 5933 2167 5947
rect 2293 5933 2307 5947
rect 2313 5933 2327 5947
rect 2113 5913 2127 5927
rect 2353 5913 2367 5927
rect 2133 5893 2147 5907
rect 2333 5893 2347 5907
rect 2073 5793 2087 5807
rect 2353 5693 2367 5707
rect 2033 5633 2047 5647
rect 2013 5593 2027 5607
rect 1933 5413 1947 5427
rect 1973 5413 1987 5427
rect 2193 5553 2207 5567
rect 2153 5413 2167 5427
rect 1913 5393 1927 5407
rect 1953 5393 1967 5407
rect 2013 5393 2027 5407
rect 2033 5393 2047 5407
rect 2133 5393 2147 5407
rect 1873 5353 1887 5367
rect 2273 5393 2287 5407
rect 2173 5373 2187 5387
rect 1933 5173 1947 5187
rect 1853 5073 1867 5087
rect 1933 5073 1947 5087
rect 1953 5013 1967 5027
rect 2213 5213 2227 5227
rect 2133 5173 2147 5187
rect 1993 5153 2007 5167
rect 2113 5153 2127 5167
rect 2053 5093 2067 5107
rect 1833 4933 1847 4947
rect 1973 4933 1987 4947
rect 1973 4913 1987 4927
rect 2033 4913 2047 4927
rect 1933 4713 1947 4727
rect 1933 4693 1947 4707
rect 1793 4673 1807 4687
rect 2013 4693 2027 4707
rect 1993 4673 2007 4687
rect 1893 4653 1907 4667
rect 1953 4653 1967 4667
rect 1973 4653 1987 4667
rect 1913 4633 1927 4647
rect 1913 4533 1927 4547
rect 1793 4493 1807 4507
rect 1833 4473 1847 4487
rect 1813 4373 1827 4387
rect 1873 4213 1887 4227
rect 1833 4113 1847 4127
rect 1873 4093 1887 4107
rect 1653 3913 1667 3927
rect 1413 3733 1427 3747
rect 1533 3753 1547 3767
rect 1433 3713 1447 3727
rect 1333 3593 1347 3607
rect 1413 3593 1427 3607
rect 1193 3573 1207 3587
rect 1233 3573 1247 3587
rect 953 3493 967 3507
rect 893 3453 907 3467
rect 973 3433 987 3447
rect 953 3213 967 3227
rect 793 3193 807 3207
rect 753 2973 767 2987
rect 953 3153 967 3167
rect 793 2953 807 2967
rect 753 2933 767 2947
rect 733 2553 747 2567
rect 913 2993 927 3007
rect 953 2993 967 3007
rect 873 2773 887 2787
rect 793 2733 807 2747
rect 893 2733 907 2747
rect 953 2733 967 2747
rect 773 2533 787 2547
rect 733 2513 747 2527
rect 753 2513 767 2527
rect 713 2473 727 2487
rect 693 2253 707 2267
rect 713 2213 727 2227
rect 1053 3493 1067 3507
rect 1433 3573 1447 3587
rect 1113 3253 1127 3267
rect 1073 3233 1087 3247
rect 1313 3233 1327 3247
rect 1353 3233 1367 3247
rect 1053 3213 1067 3227
rect 1093 3193 1107 3207
rect 1133 3193 1147 3207
rect 993 3173 1007 3187
rect 993 2933 1007 2947
rect 1353 3193 1367 3207
rect 1333 3153 1347 3167
rect 1153 3053 1167 3067
rect 1373 3053 1387 3067
rect 1133 2793 1147 2807
rect 1073 2773 1087 2787
rect 913 2713 927 2727
rect 973 2713 987 2727
rect 1413 3013 1427 3027
rect 1353 2773 1367 2787
rect 1373 2773 1387 2787
rect 1353 2753 1367 2767
rect 1393 2753 1407 2767
rect 1273 2733 1287 2747
rect 1333 2733 1347 2747
rect 1373 2733 1387 2747
rect 1113 2713 1127 2727
rect 1193 2613 1207 2627
rect 1073 2593 1087 2607
rect 793 2433 807 2447
rect 793 2273 807 2287
rect 733 2153 747 2167
rect 773 2093 787 2107
rect 633 2053 647 2067
rect 773 2053 787 2067
rect 613 2033 627 2047
rect 713 1773 727 1787
rect 673 1693 687 1707
rect 673 1673 687 1687
rect 773 1673 787 1687
rect 613 1613 627 1627
rect 713 1613 727 1627
rect 1153 2533 1167 2547
rect 873 2213 887 2227
rect 913 2153 927 2167
rect 893 2073 907 2087
rect 1153 2273 1167 2287
rect 1133 2253 1147 2267
rect 1113 2233 1127 2247
rect 1193 2233 1207 2247
rect 1193 2213 1207 2227
rect 1173 2193 1187 2207
rect 933 2093 947 2107
rect 1073 2093 1087 2107
rect 973 2073 987 2087
rect 933 1833 947 1847
rect 853 1773 867 1787
rect 813 1613 827 1627
rect 553 1573 567 1587
rect 793 1593 807 1607
rect 613 1313 627 1327
rect 633 1313 647 1327
rect 613 1133 627 1147
rect 533 813 547 827
rect 493 653 507 667
rect 553 653 567 667
rect 453 633 467 647
rect 473 613 487 627
rect 533 633 547 647
rect 493 413 507 427
rect 513 413 527 427
rect 393 313 407 327
rect 173 293 187 307
rect 213 173 227 187
rect 553 613 567 627
rect 533 353 547 367
rect 473 333 487 347
rect 513 313 527 327
rect 453 293 467 307
rect 413 173 427 187
rect 433 153 447 167
rect 693 1573 707 1587
rect 673 1313 687 1327
rect 713 1313 727 1327
rect 693 1293 707 1307
rect 733 1293 747 1307
rect 653 1273 667 1287
rect 713 1273 727 1287
rect 673 1253 687 1267
rect 693 1153 707 1167
rect 733 1253 747 1267
rect 733 1113 747 1127
rect 773 1113 787 1127
rect 753 1093 767 1107
rect 673 1073 687 1087
rect 693 893 707 907
rect 733 853 747 867
rect 673 813 687 827
rect 773 813 787 827
rect 693 773 707 787
rect 753 773 767 787
rect 653 753 667 767
rect 673 653 687 667
rect 653 613 667 627
rect 733 613 747 627
rect 713 353 727 367
rect 753 353 767 367
rect 633 333 647 347
rect 693 333 707 347
rect 733 233 747 247
rect 653 153 667 167
rect 953 1773 967 1787
rect 933 1753 947 1767
rect 913 1733 927 1747
rect 1013 1733 1027 1747
rect 873 1593 887 1607
rect 913 1593 927 1607
rect 853 1573 867 1587
rect 893 1573 907 1587
rect 1113 2053 1127 2067
rect 1093 1793 1107 1807
rect 1073 1633 1087 1647
rect 1013 1353 1027 1367
rect 1093 1313 1107 1327
rect 953 1253 967 1267
rect 993 1253 1007 1267
rect 913 1133 927 1147
rect 953 1093 967 1107
rect 973 1073 987 1087
rect 1233 2073 1247 2087
rect 1173 2053 1187 2067
rect 1213 2053 1227 2067
rect 1133 2033 1147 2047
rect 1193 2033 1207 2047
rect 1153 1793 1167 1807
rect 1133 1733 1147 1747
rect 1333 2713 1347 2727
rect 1293 2573 1307 2587
rect 1373 2573 1387 2587
rect 1393 2573 1407 2587
rect 1533 3713 1547 3727
rect 1513 3233 1527 3247
rect 1473 3213 1487 3227
rect 1453 3033 1467 3047
rect 1513 2953 1527 2967
rect 1453 2753 1467 2767
rect 1513 2713 1527 2727
rect 1433 2533 1447 2547
rect 1393 2293 1407 2307
rect 1373 2273 1387 2287
rect 1413 2273 1427 2287
rect 1473 2273 1487 2287
rect 1393 2253 1407 2267
rect 1433 2253 1447 2267
rect 1413 2193 1427 2207
rect 1453 2093 1467 2107
rect 1293 1873 1307 1887
rect 1273 1793 1287 1807
rect 1293 1753 1307 1767
rect 1193 1353 1207 1367
rect 1153 1333 1167 1347
rect 1153 1313 1167 1327
rect 1353 1753 1367 1767
rect 1393 1753 1407 1767
rect 1333 1333 1347 1347
rect 1313 1313 1327 1327
rect 1133 1293 1147 1307
rect 1173 1293 1187 1307
rect 1133 1273 1147 1287
rect 1233 1293 1247 1307
rect 1113 1233 1127 1247
rect 1153 1233 1167 1247
rect 1013 1213 1027 1227
rect 1173 1153 1187 1167
rect 1133 1113 1147 1127
rect 1313 1273 1327 1287
rect 1233 1113 1247 1127
rect 1013 1073 1027 1087
rect 1113 893 1127 907
rect 933 873 947 887
rect 993 873 1007 887
rect 893 833 907 847
rect 913 813 927 827
rect 953 793 967 807
rect 1013 793 1027 807
rect 853 773 867 787
rect 993 693 1007 707
rect 953 633 967 647
rect 913 573 927 587
rect 973 553 987 567
rect 913 353 927 367
rect 933 353 947 367
rect 873 233 887 247
rect 913 193 927 207
rect 1193 833 1207 847
rect 1173 813 1187 827
rect 1173 793 1187 807
rect 1153 733 1167 747
rect 1253 1093 1267 1107
rect 1233 793 1247 807
rect 1213 773 1227 787
rect 1193 553 1207 567
rect 1393 1733 1407 1747
rect 1373 1573 1387 1587
rect 1433 1573 1447 1587
rect 1693 3733 1707 3747
rect 1753 3733 1767 3747
rect 1673 3673 1687 3687
rect 1633 3653 1647 3667
rect 1613 3633 1627 3647
rect 1773 3493 1787 3507
rect 2013 4453 2027 4467
rect 2193 5133 2207 5147
rect 2133 4913 2147 4927
rect 2173 4753 2187 4767
rect 2113 4733 2127 4747
rect 2093 4673 2107 4687
rect 2053 4493 2067 4507
rect 2073 4493 2087 4507
rect 2253 4633 2267 4647
rect 2153 4553 2167 4567
rect 2033 4393 2047 4407
rect 2113 4453 2127 4467
rect 2073 4373 2087 4387
rect 2113 4373 2127 4387
rect 2093 4233 2107 4247
rect 2073 4173 2087 4187
rect 1973 4073 1987 4087
rect 1953 4013 1967 4027
rect 1933 3993 1947 4007
rect 1913 3713 1927 3727
rect 2253 4493 2267 4507
rect 2173 4453 2187 4467
rect 2413 5553 2427 5567
rect 2373 5433 2387 5447
rect 2453 5433 2467 5447
rect 2393 5413 2407 5427
rect 2433 5413 2447 5427
rect 2373 5373 2387 5387
rect 2333 5113 2347 5127
rect 2453 5133 2467 5147
rect 2373 5093 2387 5107
rect 2433 4953 2447 4967
rect 2553 6353 2567 6367
rect 2553 6333 2567 6347
rect 2513 6153 2527 6167
rect 2493 6133 2507 6147
rect 2533 6113 2547 6127
rect 2773 6373 2787 6387
rect 2733 6353 2747 6367
rect 2793 6153 2807 6167
rect 2633 6073 2647 6087
rect 2613 6013 2627 6027
rect 2653 6013 2667 6027
rect 2733 6013 2747 6027
rect 2633 5913 2647 5927
rect 2593 5853 2607 5867
rect 2613 5753 2627 5767
rect 2493 5713 2507 5727
rect 2573 5653 2587 5667
rect 2593 5613 2607 5627
rect 2553 5593 2567 5607
rect 2693 5593 2707 5607
rect 2573 5433 2587 5447
rect 2653 5433 2667 5447
rect 2493 5413 2507 5427
rect 2473 4913 2487 4927
rect 2373 4893 2387 4907
rect 2453 4873 2467 4887
rect 2373 4793 2387 4807
rect 2393 4613 2407 4627
rect 2373 4553 2387 4567
rect 2433 4493 2447 4507
rect 2373 4313 2387 4327
rect 2353 4273 2367 4287
rect 2293 4193 2307 4207
rect 2253 4173 2267 4187
rect 2273 4173 2287 4187
rect 2293 4153 2307 4167
rect 2313 4153 2327 4167
rect 2253 4073 2267 4087
rect 2233 4013 2247 4027
rect 2193 3793 2207 3807
rect 2153 3753 2167 3767
rect 2173 3693 2187 3707
rect 1893 3673 1907 3687
rect 2133 3673 2147 3687
rect 2133 3593 2147 3607
rect 1893 3573 1907 3587
rect 1953 3553 1967 3567
rect 2213 3733 2227 3747
rect 2193 3473 2207 3487
rect 1713 3453 1727 3467
rect 1733 3453 1747 3467
rect 1673 3313 1687 3327
rect 1653 3293 1667 3307
rect 1673 3273 1687 3287
rect 2133 3253 2147 3267
rect 1693 3233 1707 3247
rect 1633 3033 1647 3047
rect 1673 3033 1687 3047
rect 1613 3013 1627 3027
rect 1653 2993 1667 3007
rect 1573 2893 1587 2907
rect 1553 2593 1567 2607
rect 1593 2873 1607 2887
rect 1753 3213 1767 3227
rect 2033 3193 2047 3207
rect 2053 3193 2067 3207
rect 1873 3173 1887 3187
rect 1873 3053 1887 3067
rect 1733 3033 1747 3047
rect 1693 2933 1707 2947
rect 1713 2933 1727 2947
rect 1653 2773 1667 2787
rect 1593 2633 1607 2647
rect 1573 2573 1587 2587
rect 1893 2993 1907 3007
rect 1853 2893 1867 2907
rect 2113 3173 2127 3187
rect 2073 3033 2087 3047
rect 2213 3093 2227 3107
rect 2193 3033 2207 3047
rect 1673 2733 1687 2747
rect 1733 2733 1747 2747
rect 1733 2633 1747 2647
rect 1633 2613 1647 2627
rect 1633 2593 1647 2607
rect 1613 2493 1627 2507
rect 1713 2473 1727 2487
rect 1533 2073 1547 2087
rect 1573 1793 1587 1807
rect 1693 2113 1707 2127
rect 1653 2053 1667 2067
rect 1653 1953 1667 1967
rect 1693 1953 1707 1967
rect 1613 1653 1627 1667
rect 1593 1613 1607 1627
rect 1433 1313 1447 1327
rect 1413 1293 1427 1307
rect 1453 1293 1467 1307
rect 1413 1153 1427 1167
rect 1453 1153 1467 1167
rect 1393 1133 1407 1147
rect 1373 1113 1387 1127
rect 1433 1133 1447 1147
rect 1433 1073 1447 1087
rect 1353 893 1367 907
rect 1433 833 1447 847
rect 1293 733 1307 747
rect 1253 373 1267 387
rect 1153 353 1167 367
rect 1413 653 1427 667
rect 1493 1353 1507 1367
rect 1693 1553 1707 1567
rect 1673 1333 1687 1347
rect 1773 2713 1787 2727
rect 1813 2673 1827 2687
rect 1873 2673 1887 2687
rect 2173 3013 2187 3027
rect 1873 2653 1887 2667
rect 2093 2653 2107 2667
rect 1853 2573 1867 2587
rect 1773 2513 1787 2527
rect 1753 2413 1767 2427
rect 1733 2273 1747 2287
rect 1833 2413 1847 2427
rect 1793 2273 1807 2287
rect 1833 2273 1847 2287
rect 1773 2253 1787 2267
rect 2093 2613 2107 2627
rect 2033 2573 2047 2587
rect 2133 2753 2147 2767
rect 2153 2613 2167 2627
rect 2113 2573 2127 2587
rect 2053 2553 2067 2567
rect 2033 2533 2047 2547
rect 2073 2533 2087 2547
rect 1893 2273 1907 2287
rect 1753 2053 1767 2067
rect 1753 2033 1767 2047
rect 1733 1593 1747 1607
rect 1593 1293 1607 1307
rect 1493 1133 1507 1147
rect 1653 1133 1667 1147
rect 1593 1113 1607 1127
rect 1613 1113 1627 1127
rect 1473 793 1487 807
rect 1633 1093 1647 1107
rect 1573 753 1587 767
rect 1633 793 1647 807
rect 1633 733 1647 747
rect 1653 733 1667 747
rect 1373 633 1387 647
rect 1413 633 1427 647
rect 1453 633 1467 647
rect 1393 613 1407 627
rect 1433 593 1447 607
rect 1373 393 1387 407
rect 1453 393 1467 407
rect 1373 373 1387 387
rect 1413 373 1427 387
rect 1333 353 1347 367
rect 1393 353 1407 367
rect 1613 633 1627 647
rect 1653 633 1667 647
rect 1733 1233 1747 1247
rect 1733 1153 1747 1167
rect 1693 993 1707 1007
rect 1813 2073 1827 2087
rect 2093 2233 2107 2247
rect 2193 2553 2207 2567
rect 2193 2533 2207 2547
rect 2153 2493 2167 2507
rect 2173 2293 2187 2307
rect 2133 2133 2147 2147
rect 2153 2113 2167 2127
rect 1773 1813 1787 1827
rect 1753 853 1767 867
rect 1753 813 1767 827
rect 1693 693 1707 707
rect 2113 2073 2127 2087
rect 1873 2053 1887 2067
rect 1953 2053 1967 2067
rect 1913 2033 1927 2047
rect 1833 1813 1847 1827
rect 1933 1793 1947 1807
rect 1813 1773 1827 1787
rect 1853 1773 1867 1787
rect 1793 1753 1807 1767
rect 1893 1593 1907 1607
rect 2093 1773 2107 1787
rect 2173 1773 2187 1787
rect 2113 1753 2127 1767
rect 2053 1693 2067 1707
rect 2053 1673 2067 1687
rect 1973 1653 1987 1667
rect 1953 1613 1967 1627
rect 1933 1573 1947 1587
rect 2093 1613 2107 1627
rect 2133 1613 2147 1627
rect 2153 1613 2167 1627
rect 2193 1613 2207 1627
rect 2093 1593 2107 1607
rect 1873 1553 1887 1567
rect 1913 1553 1927 1567
rect 1973 1553 1987 1567
rect 2073 1553 2087 1567
rect 1933 1333 1947 1347
rect 1893 1313 1907 1327
rect 1913 1273 1927 1287
rect 1793 1133 1807 1147
rect 1893 1133 1907 1147
rect 1773 613 1787 627
rect 1673 573 1687 587
rect 1613 373 1627 387
rect 1653 373 1667 387
rect 1593 353 1607 367
rect 1133 173 1147 187
rect 1293 173 1307 187
rect 953 153 967 167
rect 1013 153 1027 167
rect 893 133 907 147
rect 1113 133 1127 147
rect 673 113 687 127
rect 813 113 827 127
rect 1553 293 1567 307
rect 1373 173 1387 187
rect 1573 173 1587 187
rect 1633 333 1647 347
rect 1673 333 1687 347
rect 1853 1093 1867 1107
rect 1873 1073 1887 1087
rect 1833 1053 1847 1067
rect 1893 1053 1907 1067
rect 2013 1313 2027 1327
rect 2033 1313 2047 1327
rect 1933 953 1947 967
rect 1873 873 1887 887
rect 1853 813 1867 827
rect 1873 793 1887 807
rect 1833 673 1847 687
rect 1893 673 1907 687
rect 1853 653 1867 667
rect 1853 633 1867 647
rect 1873 353 1887 367
rect 1793 313 1807 327
rect 1893 313 1907 327
rect 2013 853 2027 867
rect 1993 833 2007 847
rect 1973 813 1987 827
rect 1953 633 1967 647
rect 1953 593 1967 607
rect 1933 553 1947 567
rect 1933 373 1947 387
rect 1993 793 2007 807
rect 2013 793 2027 807
rect 1973 353 1987 367
rect 1913 293 1927 307
rect 1833 173 1847 187
rect 2093 1373 2107 1387
rect 2153 1373 2167 1387
rect 2113 1253 2127 1267
rect 2153 1253 2167 1267
rect 2093 1213 2107 1227
rect 2053 1113 2067 1127
rect 2073 1113 2087 1127
rect 2113 1113 2127 1127
rect 2053 1033 2067 1047
rect 2133 953 2147 967
rect 2053 853 2067 867
rect 2093 833 2107 847
rect 2073 793 2087 807
rect 2033 773 2047 787
rect 2113 753 2127 767
rect 2113 673 2127 687
rect 2093 653 2107 667
rect 2153 893 2167 907
rect 2153 833 2167 847
rect 2213 733 2227 747
rect 2153 653 2167 667
rect 2153 613 2167 627
rect 2053 373 2067 387
rect 2113 333 2127 347
rect 2053 313 2067 327
rect 2093 313 2107 327
rect 2153 313 2167 327
rect 2033 293 2047 307
rect 2013 173 2027 187
rect 1993 153 2007 167
rect 2273 3973 2287 3987
rect 2253 3313 2267 3327
rect 2253 2993 2267 3007
rect 2273 2993 2287 3007
rect 2353 4133 2367 4147
rect 2493 4653 2507 4667
rect 2453 4273 2467 4287
rect 2533 4273 2547 4287
rect 2453 4253 2467 4267
rect 2373 3973 2387 3987
rect 2433 3793 2447 3807
rect 2373 3773 2387 3787
rect 2393 3773 2407 3787
rect 2433 3553 2447 3567
rect 2413 3533 2427 3547
rect 2673 5413 2687 5427
rect 2893 7073 2907 7087
rect 2873 7033 2887 7047
rect 2873 6853 2887 6867
rect 2933 6853 2947 6867
rect 2833 6833 2847 6847
rect 2833 6813 2847 6827
rect 2873 6613 2887 6627
rect 2833 6593 2847 6607
rect 2833 6113 2847 6127
rect 2833 6093 2847 6107
rect 2813 6013 2827 6027
rect 2853 5933 2867 5947
rect 2793 5893 2807 5907
rect 2933 6553 2947 6567
rect 2893 6353 2907 6367
rect 3013 8573 3027 8587
rect 3093 9633 3107 9647
rect 3073 9533 3087 9547
rect 3053 9513 3067 9527
rect 3053 9253 3067 9267
rect 3053 9013 3067 9027
rect 3153 10373 3167 10387
rect 3273 10913 3287 10927
rect 3413 11193 3427 11207
rect 3493 11193 3507 11207
rect 3433 11153 3447 11167
rect 3553 11133 3567 11147
rect 3473 11113 3487 11127
rect 3753 11193 3767 11207
rect 3713 11153 3727 11167
rect 3533 10773 3547 10787
rect 3413 10713 3427 10727
rect 3493 10653 3507 10667
rect 3453 10633 3467 10647
rect 3373 10553 3387 10567
rect 3313 10453 3327 10467
rect 3353 10453 3367 10467
rect 3433 10513 3447 10527
rect 3573 10513 3587 10527
rect 3333 10413 3347 10427
rect 3373 10413 3387 10427
rect 3273 10253 3287 10267
rect 3293 10253 3307 10267
rect 3373 10253 3387 10267
rect 3393 10253 3407 10267
rect 3313 10233 3327 10247
rect 3373 10213 3387 10227
rect 3253 9993 3267 10007
rect 3193 9793 3207 9807
rect 3273 9953 3287 9967
rect 3413 9953 3427 9967
rect 3273 9773 3287 9787
rect 3393 9913 3407 9927
rect 3253 9653 3267 9667
rect 3293 9653 3307 9667
rect 3233 9493 3247 9507
rect 3173 9453 3187 9467
rect 3153 9433 3167 9447
rect 3153 9393 3167 9407
rect 3193 9333 3207 9347
rect 3213 9333 3227 9347
rect 3133 9313 3147 9327
rect 3113 9273 3127 9287
rect 3153 9273 3167 9287
rect 3133 9253 3147 9267
rect 3173 9093 3187 9107
rect 3553 10353 3567 10367
rect 3513 10253 3527 10267
rect 3613 10433 3627 10447
rect 3653 10433 3667 10447
rect 3593 10413 3607 10427
rect 3593 10273 3607 10287
rect 3573 10253 3587 10267
rect 3653 10273 3667 10287
rect 3653 10253 3667 10267
rect 3533 10213 3547 10227
rect 3573 10213 3587 10227
rect 3633 10213 3647 10227
rect 3533 10013 3547 10027
rect 3453 9973 3467 9987
rect 3493 9953 3507 9967
rect 3453 9933 3467 9947
rect 3513 9933 3527 9947
rect 3553 9933 3567 9947
rect 3473 9913 3487 9927
rect 3513 9913 3527 9927
rect 3533 9913 3547 9927
rect 3413 9493 3427 9507
rect 3433 9493 3447 9507
rect 3473 9493 3487 9507
rect 3413 9473 3427 9487
rect 3453 9473 3467 9487
rect 3333 9453 3347 9467
rect 3433 9453 3447 9467
rect 3393 9413 3407 9427
rect 3393 9373 3407 9387
rect 3393 9293 3407 9307
rect 3373 9273 3387 9287
rect 3413 9233 3427 9247
rect 3333 9213 3347 9227
rect 3453 9033 3467 9047
rect 3073 8773 3087 8787
rect 3153 9013 3167 9027
rect 3213 9013 3227 9027
rect 3293 9013 3307 9027
rect 3193 8993 3207 9007
rect 3153 8833 3167 8847
rect 3193 8793 3207 8807
rect 3133 8773 3147 8787
rect 3113 8673 3127 8687
rect 3173 8673 3187 8687
rect 3133 8653 3147 8667
rect 3153 8653 3167 8667
rect 3033 8513 3047 8527
rect 2993 8493 3007 8507
rect 3093 8513 3107 8527
rect 3133 8513 3147 8527
rect 3293 8953 3307 8967
rect 3273 8773 3287 8787
rect 3313 8833 3327 8847
rect 3313 8813 3327 8827
rect 3413 8813 3427 8827
rect 3293 8733 3307 8747
rect 3073 8493 3087 8507
rect 3113 8493 3127 8507
rect 3053 8473 3067 8487
rect 3093 8473 3107 8487
rect 3033 8313 3047 8327
rect 3113 8313 3127 8327
rect 3053 8273 3067 8287
rect 3193 8453 3207 8467
rect 3253 8333 3267 8347
rect 3393 8773 3407 8787
rect 3493 9373 3507 9387
rect 3493 9033 3507 9047
rect 3453 8753 3467 8767
rect 3453 8533 3467 8547
rect 3313 8513 3327 8527
rect 3313 8473 3327 8487
rect 3313 8313 3327 8327
rect 3253 8293 3267 8307
rect 3293 8293 3307 8307
rect 3333 8293 3347 8307
rect 3413 8293 3427 8307
rect 3153 8233 3167 8247
rect 3133 8173 3147 8187
rect 3053 8153 3067 8167
rect 3033 8113 3047 8127
rect 3013 8073 3027 8087
rect 2973 8013 2987 8027
rect 2993 8013 3007 8027
rect 3033 7993 3047 8007
rect 2993 7853 3007 7867
rect 2993 7813 3007 7827
rect 2973 7373 2987 7387
rect 2973 7313 2987 7327
rect 2973 6113 2987 6127
rect 2973 6093 2987 6107
rect 2893 5953 2907 5967
rect 2873 5693 2887 5707
rect 2773 5633 2787 5647
rect 2813 5633 2827 5647
rect 2853 5633 2867 5647
rect 2773 5553 2787 5567
rect 2833 5613 2847 5627
rect 2833 5573 2847 5587
rect 2793 5513 2807 5527
rect 2773 5493 2787 5507
rect 2753 5473 2767 5487
rect 2713 5393 2727 5407
rect 2653 5133 2667 5147
rect 2713 5153 2727 5167
rect 2693 5113 2707 5127
rect 2713 4953 2727 4967
rect 2653 4933 2667 4947
rect 2693 4873 2707 4887
rect 2733 4733 2747 4747
rect 2653 4693 2667 4707
rect 2613 4673 2627 4687
rect 2613 4613 2627 4627
rect 2673 4653 2687 4667
rect 2673 4553 2687 4567
rect 2633 4493 2647 4507
rect 2633 4473 2647 4487
rect 2593 4373 2607 4387
rect 2573 4253 2587 4267
rect 2533 4193 2547 4207
rect 2553 4193 2567 4207
rect 2613 4293 2627 4307
rect 2573 4013 2587 4027
rect 2613 4013 2627 4027
rect 2473 3993 2487 4007
rect 2453 3533 2467 3547
rect 2353 3473 2367 3487
rect 2333 3433 2347 3447
rect 2453 3513 2467 3527
rect 2373 3273 2387 3287
rect 2313 3253 2327 3267
rect 2373 3253 2387 3267
rect 2333 3013 2347 3027
rect 2293 2973 2307 2987
rect 2313 2773 2327 2787
rect 2313 2693 2327 2707
rect 2273 2633 2287 2647
rect 2273 2533 2287 2547
rect 2293 2513 2307 2527
rect 2333 2513 2347 2527
rect 2373 2673 2387 2687
rect 2353 2473 2367 2487
rect 2333 2293 2347 2307
rect 2313 2273 2327 2287
rect 2433 3413 2447 3427
rect 2413 3193 2427 3207
rect 2453 3213 2467 3227
rect 2433 3013 2447 3027
rect 2413 2593 2427 2607
rect 2333 2253 2347 2267
rect 2393 2253 2407 2267
rect 2273 2233 2287 2247
rect 2293 2073 2307 2087
rect 2293 2033 2307 2047
rect 2273 1753 2287 1767
rect 2253 1273 2267 1287
rect 2373 2233 2387 2247
rect 2353 2073 2367 2087
rect 2393 2073 2407 2087
rect 2393 1913 2407 1927
rect 2333 1653 2347 1667
rect 2353 1613 2367 1627
rect 2393 1553 2407 1567
rect 2433 2533 2447 2547
rect 2453 2253 2467 2267
rect 2433 1773 2447 1787
rect 2433 1593 2447 1607
rect 2413 1333 2427 1347
rect 2313 1293 2327 1307
rect 2333 1293 2347 1307
rect 2373 1293 2387 1307
rect 2353 1253 2367 1267
rect 2313 1153 2327 1167
rect 2313 1133 2327 1147
rect 2293 1113 2307 1127
rect 2273 1073 2287 1087
rect 2433 1253 2447 1267
rect 2373 1113 2387 1127
rect 2393 1073 2407 1087
rect 2353 933 2367 947
rect 2333 813 2347 827
rect 2373 813 2387 827
rect 2353 753 2367 767
rect 2393 753 2407 767
rect 2373 673 2387 687
rect 2313 593 2327 607
rect 2513 3973 2527 3987
rect 2653 4233 2667 4247
rect 2653 4193 2667 4207
rect 2533 3953 2547 3967
rect 2633 3953 2647 3967
rect 2493 3933 2507 3947
rect 2513 3893 2527 3907
rect 2493 3813 2507 3827
rect 2593 3933 2607 3947
rect 2573 3913 2587 3927
rect 2513 3693 2527 3707
rect 2533 3693 2547 3707
rect 2513 3553 2527 3567
rect 2533 3533 2547 3547
rect 2713 4493 2727 4507
rect 2713 4193 2727 4207
rect 2733 4193 2747 4207
rect 2773 5413 2787 5427
rect 2793 4953 2807 4967
rect 2933 5633 2947 5647
rect 2973 5593 2987 5607
rect 2913 5573 2927 5587
rect 3053 7813 3067 7827
rect 3013 7793 3027 7807
rect 3213 8073 3227 8087
rect 3253 8033 3267 8047
rect 3193 7993 3207 8007
rect 3193 7973 3207 7987
rect 3233 7933 3247 7947
rect 3233 7853 3247 7867
rect 3293 7853 3307 7867
rect 3153 7613 3167 7627
rect 3113 7513 3127 7527
rect 3093 7493 3107 7507
rect 3093 7453 3107 7467
rect 3033 7333 3047 7347
rect 3013 7313 3027 7327
rect 3033 7133 3047 7147
rect 3053 7133 3067 7147
rect 3053 6853 3067 6867
rect 3113 7333 3127 7347
rect 3273 7773 3287 7787
rect 3293 7573 3307 7587
rect 3353 7573 3367 7587
rect 3393 7573 3407 7587
rect 3233 7553 3247 7567
rect 3373 7533 3387 7547
rect 3333 7513 3347 7527
rect 3233 7373 3247 7387
rect 3253 7373 3267 7387
rect 3213 7353 3227 7367
rect 3293 7353 3307 7367
rect 3253 7253 3267 7267
rect 3193 7133 3207 7147
rect 3153 7093 3167 7107
rect 3193 7093 3207 7107
rect 3133 7033 3147 7047
rect 3033 6593 3047 6607
rect 3073 6833 3087 6847
rect 3213 6953 3227 6967
rect 3173 6813 3187 6827
rect 3193 6813 3207 6827
rect 3113 6693 3127 6707
rect 3133 6593 3147 6607
rect 3173 6593 3187 6607
rect 3153 6553 3167 6567
rect 3053 6513 3067 6527
rect 3113 6253 3127 6267
rect 3013 5913 3027 5927
rect 3013 5633 3027 5647
rect 2933 5493 2947 5507
rect 2913 5453 2927 5467
rect 2893 5433 2907 5447
rect 2853 5413 2867 5427
rect 2973 5433 2987 5447
rect 2953 5413 2967 5427
rect 2893 5393 2907 5407
rect 2893 5173 2907 5187
rect 2893 5153 2907 5167
rect 2933 5153 2947 5167
rect 2913 5133 2927 5147
rect 3133 6173 3147 6187
rect 3173 6133 3187 6147
rect 3193 5973 3207 5987
rect 3233 5913 3247 5927
rect 3153 5673 3167 5687
rect 3113 5653 3127 5667
rect 3113 5633 3127 5647
rect 3053 5613 3067 5627
rect 3133 5593 3147 5607
rect 3033 5553 3047 5567
rect 3053 5553 3067 5567
rect 3033 5413 3047 5427
rect 2973 5133 2987 5147
rect 3013 5133 3027 5147
rect 2893 4973 2907 4987
rect 2893 4953 2907 4967
rect 2873 4933 2887 4947
rect 3033 5093 3047 5107
rect 3013 4993 3027 5007
rect 2993 4953 3007 4967
rect 2973 4933 2987 4947
rect 2953 4873 2967 4887
rect 2893 4673 2907 4687
rect 2833 4573 2847 4587
rect 2813 4513 2827 4527
rect 2873 4493 2887 4507
rect 2933 4493 2947 4507
rect 2833 4473 2847 4487
rect 2933 4473 2947 4487
rect 2853 4453 2867 4467
rect 2773 4433 2787 4447
rect 2913 4253 2927 4267
rect 2993 4453 3007 4467
rect 2933 4213 2947 4227
rect 2913 4193 2927 4207
rect 2933 4193 2947 4207
rect 2913 4153 2927 4167
rect 2753 4113 2767 4127
rect 2833 4053 2847 4067
rect 2713 4013 2727 4027
rect 2753 3993 2767 4007
rect 2773 3993 2787 4007
rect 2813 3973 2827 3987
rect 2733 3953 2747 3967
rect 2693 3753 2707 3767
rect 2813 3753 2827 3767
rect 2653 3713 2667 3727
rect 2733 3713 2747 3727
rect 2593 3473 2607 3487
rect 2673 3693 2687 3707
rect 2693 3693 2707 3707
rect 2713 3513 2727 3527
rect 2673 3493 2687 3507
rect 2653 3473 2667 3487
rect 2693 3473 2707 3487
rect 2633 3313 2647 3327
rect 2593 3253 2607 3267
rect 2633 3253 2647 3267
rect 2653 3253 2667 3267
rect 2553 3053 2567 3067
rect 2673 3233 2687 3247
rect 2653 3193 2667 3207
rect 2633 3113 2647 3127
rect 2613 3093 2627 3107
rect 2533 2993 2547 3007
rect 2533 2973 2547 2987
rect 2513 2593 2527 2607
rect 2493 2513 2507 2527
rect 2613 2973 2627 2987
rect 2573 2953 2587 2967
rect 2573 2753 2587 2767
rect 2613 2753 2627 2767
rect 2633 2733 2647 2747
rect 2593 2713 2607 2727
rect 2633 2693 2647 2707
rect 2553 2653 2567 2667
rect 2593 2593 2607 2607
rect 2553 2553 2567 2567
rect 2753 3573 2767 3587
rect 2733 3473 2747 3487
rect 2733 3213 2747 3227
rect 2653 2633 2667 2647
rect 2653 2573 2667 2587
rect 2573 2533 2587 2547
rect 2613 2533 2627 2547
rect 2653 2533 2667 2547
rect 2653 2333 2667 2347
rect 2673 2333 2687 2347
rect 2533 2293 2547 2307
rect 2593 2293 2607 2307
rect 2633 2293 2647 2307
rect 2713 2653 2727 2667
rect 2813 3513 2827 3527
rect 2913 4033 2927 4047
rect 2873 3713 2887 3727
rect 2993 4093 3007 4107
rect 2953 4013 2967 4027
rect 3073 5133 3087 5147
rect 3393 7073 3407 7087
rect 3333 7033 3347 7047
rect 3353 7013 3367 7027
rect 3333 6853 3347 6867
rect 3393 6853 3407 6867
rect 3293 6833 3307 6847
rect 3353 6833 3367 6847
rect 3353 6813 3367 6827
rect 3313 6793 3327 6807
rect 3533 9773 3547 9787
rect 3553 9773 3567 9787
rect 3533 9733 3547 9747
rect 3593 9953 3607 9967
rect 3633 9933 3647 9947
rect 3653 9933 3667 9947
rect 3593 9893 3607 9907
rect 3633 9833 3647 9847
rect 3593 9793 3607 9807
rect 3573 9453 3587 9467
rect 3553 8813 3567 8827
rect 3573 8533 3587 8547
rect 3613 9713 3627 9727
rect 4173 11193 4187 11207
rect 3873 10913 3887 10927
rect 3913 10913 3927 10927
rect 3893 10853 3907 10867
rect 3833 10753 3847 10767
rect 3793 10733 3807 10747
rect 3773 10693 3787 10707
rect 3713 10293 3727 10307
rect 3873 10613 3887 10627
rect 3793 10453 3807 10467
rect 3853 10453 3867 10467
rect 3773 10253 3787 10267
rect 3713 10193 3727 10207
rect 3833 10373 3847 10387
rect 3833 10273 3847 10287
rect 3813 10253 3827 10267
rect 3873 10253 3887 10267
rect 3813 10233 3827 10247
rect 3853 10233 3867 10247
rect 3833 10193 3847 10207
rect 3793 10173 3807 10187
rect 3693 9773 3707 9787
rect 3733 9773 3747 9787
rect 3673 9693 3687 9707
rect 3633 9613 3647 9627
rect 3793 9953 3807 9967
rect 3773 9933 3787 9947
rect 3833 9853 3847 9867
rect 3853 9813 3867 9827
rect 3833 9793 3847 9807
rect 3793 9773 3807 9787
rect 3733 9733 3747 9747
rect 3773 9713 3787 9727
rect 3773 9613 3787 9627
rect 3693 9493 3707 9507
rect 3733 9493 3747 9507
rect 3673 9453 3687 9467
rect 3633 9273 3647 9287
rect 3673 9273 3687 9287
rect 3613 9233 3627 9247
rect 3633 9213 3647 9227
rect 3613 8993 3627 9007
rect 3713 9053 3727 9067
rect 3693 9033 3707 9047
rect 3633 8933 3647 8947
rect 3633 8833 3647 8847
rect 3673 8813 3687 8827
rect 3633 8773 3647 8787
rect 3613 8753 3627 8767
rect 3653 8753 3667 8767
rect 3673 8753 3687 8767
rect 3613 8733 3627 8747
rect 3633 8673 3647 8687
rect 3613 8413 3627 8427
rect 3573 8313 3587 8327
rect 3553 8273 3567 8287
rect 3593 8273 3607 8287
rect 3513 8253 3527 8267
rect 3553 8253 3567 8267
rect 3513 8073 3527 8087
rect 3493 7953 3507 7967
rect 3473 7873 3487 7887
rect 3533 7873 3547 7887
rect 3433 7833 3447 7847
rect 3473 7533 3487 7547
rect 3453 7413 3467 7427
rect 3433 7373 3447 7387
rect 3573 8033 3587 8047
rect 3553 7413 3567 7427
rect 3493 7393 3507 7407
rect 3513 7353 3527 7367
rect 3473 7073 3487 7087
rect 3433 6813 3447 6827
rect 3413 6613 3427 6627
rect 3393 6393 3407 6407
rect 3453 6553 3467 6567
rect 3333 6373 3347 6387
rect 3433 6373 3447 6387
rect 3473 6373 3487 6387
rect 3393 6233 3407 6247
rect 3373 6213 3387 6227
rect 3473 6133 3487 6147
rect 3413 6113 3427 6127
rect 3473 6113 3487 6127
rect 3333 6073 3347 6087
rect 3293 6013 3307 6027
rect 3293 5993 3307 6007
rect 3373 5953 3387 5967
rect 3353 5933 3367 5947
rect 3313 5893 3327 5907
rect 3353 5893 3367 5907
rect 3233 5573 3247 5587
rect 3253 5573 3267 5587
rect 3173 5533 3187 5547
rect 3153 5473 3167 5487
rect 3213 5513 3227 5527
rect 3253 5493 3267 5507
rect 3193 5413 3207 5427
rect 3153 5093 3167 5107
rect 3113 4953 3127 4967
rect 3173 5033 3187 5047
rect 3173 4953 3187 4967
rect 3133 4933 3147 4947
rect 3193 4873 3207 4887
rect 3133 4753 3147 4767
rect 3133 4733 3147 4747
rect 3053 4693 3067 4707
rect 3093 4673 3107 4687
rect 3173 4693 3187 4707
rect 3113 4553 3127 4567
rect 3173 4553 3187 4567
rect 3093 4493 3107 4507
rect 3153 4493 3167 4507
rect 3053 4473 3067 4487
rect 3113 4453 3127 4467
rect 3053 4433 3067 4447
rect 3073 4433 3087 4447
rect 3033 4173 3047 4187
rect 3013 4053 3027 4067
rect 3033 3993 3047 4007
rect 3013 3973 3027 3987
rect 2933 3953 2947 3967
rect 2953 3953 2967 3967
rect 2973 3953 2987 3967
rect 3073 4293 3087 4307
rect 3093 3993 3107 4007
rect 3193 4433 3207 4447
rect 3233 4213 3247 4227
rect 3293 5613 3307 5627
rect 3293 5573 3307 5587
rect 3353 5773 3367 5787
rect 3313 5553 3327 5567
rect 3313 5453 3327 5467
rect 3293 5133 3307 5147
rect 3293 5113 3307 5127
rect 3333 5153 3347 5167
rect 3393 5893 3407 5907
rect 3473 5653 3487 5667
rect 3433 5593 3447 5607
rect 3393 5513 3407 5527
rect 3373 5453 3387 5467
rect 3413 5413 3427 5427
rect 3453 5413 3467 5427
rect 3413 5373 3427 5387
rect 3473 5253 3487 5267
rect 3453 5173 3467 5187
rect 3393 5153 3407 5167
rect 3433 5133 3447 5147
rect 3373 5033 3387 5047
rect 3453 4973 3467 4987
rect 3413 4953 3427 4967
rect 3333 4713 3347 4727
rect 3333 4693 3347 4707
rect 3433 4873 3447 4887
rect 3393 4713 3407 4727
rect 3433 4713 3447 4727
rect 3313 4553 3327 4567
rect 3353 4513 3367 4527
rect 3333 4493 3347 4507
rect 3313 4253 3327 4267
rect 3273 4193 3287 4207
rect 3293 4193 3307 4207
rect 3273 4133 3287 4147
rect 3253 4033 3267 4047
rect 3273 3993 3287 4007
rect 3193 3973 3207 3987
rect 3233 3973 3247 3987
rect 3253 3973 3267 3987
rect 3213 3953 3227 3967
rect 3173 3933 3187 3947
rect 3093 3733 3107 3747
rect 3173 3733 3187 3747
rect 3113 3713 3127 3727
rect 3193 3713 3207 3727
rect 3213 3713 3227 3727
rect 3053 3593 3067 3607
rect 2893 3573 2907 3587
rect 2893 3553 2907 3567
rect 2913 3553 2927 3567
rect 2873 3533 2887 3547
rect 2993 3273 3007 3287
rect 2833 3253 2847 3267
rect 2853 3193 2867 3207
rect 2853 3053 2867 3067
rect 2833 3013 2847 3027
rect 2793 2773 2807 2787
rect 2793 2733 2807 2747
rect 3033 3213 3047 3227
rect 3013 3173 3027 3187
rect 3033 3173 3047 3187
rect 2993 2793 3007 2807
rect 2833 2633 2847 2647
rect 2753 2613 2767 2627
rect 2813 2613 2827 2627
rect 2553 2273 2567 2287
rect 2533 2253 2547 2267
rect 2573 2233 2587 2247
rect 2833 2593 2847 2607
rect 3133 3673 3147 3687
rect 3193 3573 3207 3587
rect 3193 3533 3207 3547
rect 3133 3513 3147 3527
rect 3153 3513 3167 3527
rect 3193 3513 3207 3527
rect 3093 3493 3107 3507
rect 3173 3493 3187 3507
rect 3073 3273 3087 3287
rect 3053 3113 3067 3127
rect 3053 3093 3067 3107
rect 3173 3473 3187 3487
rect 3133 3173 3147 3187
rect 3133 3113 3147 3127
rect 3033 2993 3047 3007
rect 3073 2993 3087 3007
rect 3093 2993 3107 3007
rect 3053 2793 3067 2807
rect 3033 2733 3047 2747
rect 3073 2733 3087 2747
rect 3013 2533 3027 2547
rect 2513 2113 2527 2127
rect 2553 2113 2567 2127
rect 2673 2113 2687 2127
rect 2573 2093 2587 2107
rect 2613 2033 2627 2047
rect 2593 1833 2607 1847
rect 2513 1813 2527 1827
rect 2493 1793 2507 1807
rect 2533 1793 2547 1807
rect 2513 1773 2527 1787
rect 2553 1753 2567 1767
rect 2553 1713 2567 1727
rect 2573 1653 2587 1667
rect 2573 1633 2587 1647
rect 2813 2233 2827 2247
rect 2773 2093 2787 2107
rect 2893 2093 2907 2107
rect 2653 1913 2667 1927
rect 2693 1913 2707 1927
rect 2753 2073 2767 2087
rect 2813 2073 2827 2087
rect 2853 2073 2867 2087
rect 2773 2053 2787 2067
rect 2833 2053 2847 2067
rect 2873 2033 2887 2047
rect 3013 2113 3027 2127
rect 2753 1793 2767 1807
rect 2893 1793 2907 1807
rect 2933 1793 2947 1807
rect 2973 1793 2987 1807
rect 3013 1793 3027 1807
rect 2733 1773 2747 1787
rect 2753 1733 2767 1747
rect 2733 1693 2747 1707
rect 2613 1593 2627 1607
rect 2493 1573 2507 1587
rect 2613 1493 2627 1507
rect 2493 1293 2507 1307
rect 2473 813 2487 827
rect 2453 593 2467 607
rect 2293 413 2307 427
rect 2533 1233 2547 1247
rect 2553 1233 2567 1247
rect 2593 1313 2607 1327
rect 2593 1273 2607 1287
rect 2573 1213 2587 1227
rect 2573 1113 2587 1127
rect 2553 1093 2567 1107
rect 2613 1133 2627 1147
rect 2553 913 2567 927
rect 2613 893 2627 907
rect 2853 1693 2867 1707
rect 2813 1593 2827 1607
rect 2873 1613 2887 1627
rect 2833 1493 2847 1507
rect 2833 1313 2847 1327
rect 2793 1233 2807 1247
rect 2933 1693 2947 1707
rect 2893 1173 2907 1187
rect 2833 1093 2847 1107
rect 2813 1073 2827 1087
rect 2873 1073 2887 1087
rect 2853 993 2867 1007
rect 2813 953 2827 967
rect 2793 913 2807 927
rect 2753 853 2767 867
rect 2573 833 2587 847
rect 2573 713 2587 727
rect 2493 633 2507 647
rect 2593 593 2607 607
rect 2553 573 2567 587
rect 2473 393 2487 407
rect 2573 393 2587 407
rect 2233 373 2247 387
rect 2313 353 2327 367
rect 2533 373 2547 387
rect 2293 313 2307 327
rect 2313 313 2327 327
rect 2473 313 2487 327
rect 2213 193 2227 207
rect 2273 193 2287 207
rect 1973 113 1987 127
rect 2253 113 2267 127
rect 2493 173 2507 187
rect 2553 153 2567 167
rect 2853 853 2867 867
rect 2833 813 2847 827
rect 2813 613 2827 627
rect 3093 2233 3107 2247
rect 3093 2213 3107 2227
rect 3073 2073 3087 2087
rect 3133 2113 3147 2127
rect 3053 1793 3067 1807
rect 3033 1653 3047 1667
rect 3153 2033 3167 2047
rect 3133 1873 3147 1887
rect 3113 1733 3127 1747
rect 3093 1613 3107 1627
rect 3173 1773 3187 1787
rect 3253 3933 3267 3947
rect 3233 3513 3247 3527
rect 3333 4173 3347 4187
rect 3313 3913 3327 3927
rect 3293 3733 3307 3747
rect 3233 3373 3247 3387
rect 3373 3713 3387 3727
rect 3353 3673 3367 3687
rect 3373 3553 3387 3567
rect 3513 7093 3527 7107
rect 3593 7893 3607 7907
rect 3653 8273 3667 8287
rect 3633 7633 3647 7647
rect 3593 7553 3607 7567
rect 3613 7533 3627 7547
rect 3573 7093 3587 7107
rect 3613 7093 3627 7107
rect 3633 7073 3647 7087
rect 3593 7033 3607 7047
rect 3613 6913 3627 6927
rect 3533 6893 3547 6907
rect 3573 6853 3587 6867
rect 3633 6853 3647 6867
rect 3513 5913 3527 5927
rect 3653 6753 3667 6767
rect 3593 6613 3607 6627
rect 3573 6413 3587 6427
rect 3613 6413 3627 6427
rect 3553 6093 3567 6107
rect 3593 6393 3607 6407
rect 3653 6553 3667 6567
rect 3733 8953 3747 8967
rect 3733 8873 3747 8887
rect 3713 8773 3727 8787
rect 3733 8673 3747 8687
rect 3753 8493 3767 8507
rect 3733 8373 3747 8387
rect 3753 8333 3767 8347
rect 3733 8253 3747 8267
rect 3713 8033 3727 8047
rect 3793 9253 3807 9267
rect 3793 9233 3807 9247
rect 3833 9313 3847 9327
rect 4113 11173 4127 11187
rect 4293 11173 4307 11187
rect 4033 10913 4047 10927
rect 4073 10913 4087 10927
rect 4653 11233 4667 11247
rect 6113 11233 6127 11247
rect 6133 11233 6147 11247
rect 4593 11193 4607 11207
rect 4373 11173 4387 11187
rect 4393 11153 4407 11167
rect 4613 11153 4627 11167
rect 4353 10913 4367 10927
rect 3933 10853 3947 10867
rect 3933 10833 3947 10847
rect 3913 10333 3927 10347
rect 3913 10153 3927 10167
rect 3893 9873 3907 9887
rect 3873 9633 3887 9647
rect 3913 9393 3927 9407
rect 3873 9293 3887 9307
rect 3893 9273 3907 9287
rect 4553 10913 4567 10927
rect 4093 10873 4107 10887
rect 4173 10853 4187 10867
rect 4333 10853 4347 10867
rect 4053 10813 4067 10827
rect 4113 10813 4127 10827
rect 4033 10793 4047 10807
rect 4073 10793 4087 10807
rect 4093 10793 4107 10807
rect 4033 10753 4047 10767
rect 3993 10733 4007 10747
rect 4033 10733 4047 10747
rect 4013 10713 4027 10727
rect 3993 10693 4007 10707
rect 4093 10573 4107 10587
rect 4113 10493 4127 10507
rect 4053 10433 4067 10447
rect 4093 10353 4107 10367
rect 4153 10253 4167 10267
rect 4053 10213 4067 10227
rect 4033 10193 4047 10207
rect 4073 10173 4087 10187
rect 3993 9973 4007 9987
rect 4053 9973 4067 9987
rect 3993 9933 4007 9947
rect 4013 9933 4027 9947
rect 4013 9753 4027 9767
rect 4013 9693 4027 9707
rect 4153 9953 4167 9967
rect 4073 9753 4087 9767
rect 4053 9653 4067 9667
rect 3953 9433 3967 9447
rect 3833 9253 3847 9267
rect 3873 9113 3887 9127
rect 3813 9033 3827 9047
rect 3913 9033 3927 9047
rect 3833 8993 3847 9007
rect 3853 8933 3867 8947
rect 3813 8893 3827 8907
rect 3853 8893 3867 8907
rect 3873 8753 3887 8767
rect 3833 8733 3847 8747
rect 3893 8713 3907 8727
rect 3833 8573 3847 8587
rect 3813 8533 3827 8547
rect 3793 8473 3807 8487
rect 3853 8493 3867 8507
rect 3833 8453 3847 8467
rect 3713 7913 3727 7927
rect 3693 7893 3707 7907
rect 3693 7853 3707 7867
rect 3753 7873 3767 7887
rect 3733 7813 3747 7827
rect 3693 7573 3707 7587
rect 3833 8313 3847 8327
rect 3873 8313 3887 8327
rect 3813 8293 3827 8307
rect 3833 8273 3847 8287
rect 3853 8093 3867 8107
rect 3793 7553 3807 7567
rect 3833 7553 3847 7567
rect 3773 7433 3787 7447
rect 3773 7393 3787 7407
rect 3713 7373 3727 7387
rect 3753 7373 3767 7387
rect 3753 7213 3767 7227
rect 3733 7093 3747 7107
rect 3673 6493 3687 6507
rect 3753 6873 3767 6887
rect 3873 8073 3887 8087
rect 3873 8033 3887 8047
rect 3933 8833 3947 8847
rect 3913 8313 3927 8327
rect 3973 8533 3987 8547
rect 4053 9473 4067 9487
rect 4113 9473 4127 9487
rect 4133 9453 4147 9467
rect 4093 9433 4107 9447
rect 4053 9393 4067 9407
rect 4093 9313 4107 9327
rect 4113 9293 4127 9307
rect 4153 9253 4167 9267
rect 4113 9133 4127 9147
rect 4073 9093 4087 9107
rect 4033 9033 4047 9047
rect 4053 8993 4067 9007
rect 4073 8853 4087 8867
rect 4113 8833 4127 8847
rect 4053 8773 4067 8787
rect 4093 8753 4107 8767
rect 4113 8593 4127 8607
rect 4033 8513 4047 8527
rect 4073 8513 4087 8527
rect 4013 8313 4027 8327
rect 3953 8293 3967 8307
rect 3973 8293 3987 8307
rect 3953 8093 3967 8107
rect 3953 8033 3967 8047
rect 3993 8033 4007 8047
rect 3913 8013 3927 8027
rect 3913 7893 3927 7907
rect 3933 7873 3947 7887
rect 3893 7853 3907 7867
rect 3993 8013 4007 8027
rect 3973 7853 3987 7867
rect 3973 7833 3987 7847
rect 3873 7813 3887 7827
rect 3953 7813 3967 7827
rect 3853 7453 3867 7467
rect 3813 7413 3827 7427
rect 3853 7373 3867 7387
rect 3793 7253 3807 7267
rect 3813 7073 3827 7087
rect 3833 6933 3847 6947
rect 3873 7013 3887 7027
rect 3853 6913 3867 6927
rect 3853 6893 3867 6907
rect 3813 6873 3827 6887
rect 3753 6573 3767 6587
rect 3833 6853 3847 6867
rect 3813 6613 3827 6627
rect 3873 6613 3887 6627
rect 3893 6593 3907 6607
rect 3853 6553 3867 6567
rect 3873 6553 3887 6567
rect 3773 6453 3787 6467
rect 3753 6393 3767 6407
rect 3813 6393 3827 6407
rect 3853 6393 3867 6407
rect 3833 6373 3847 6387
rect 3913 6413 3927 6427
rect 3913 6373 3927 6387
rect 3893 6353 3907 6367
rect 3893 6293 3907 6307
rect 3753 6153 3767 6167
rect 3733 6113 3747 6127
rect 3733 6073 3747 6087
rect 3713 6013 3727 6027
rect 3633 5913 3647 5927
rect 3693 5913 3707 5927
rect 3533 5793 3547 5807
rect 3653 5873 3667 5887
rect 3593 5713 3607 5727
rect 3613 5633 3627 5647
rect 3593 5613 3607 5627
rect 3633 5613 3647 5627
rect 3593 5573 3607 5587
rect 3573 5533 3587 5547
rect 3513 5493 3527 5507
rect 3633 5453 3647 5467
rect 3593 5433 3607 5447
rect 3513 5413 3527 5427
rect 3593 5173 3607 5187
rect 3513 5133 3527 5147
rect 3553 5033 3567 5047
rect 3553 4973 3567 4987
rect 3673 5193 3687 5207
rect 3633 5173 3647 5187
rect 3613 5153 3627 5167
rect 3593 4953 3607 4967
rect 3693 5013 3707 5027
rect 3653 4993 3667 5007
rect 3693 4953 3707 4967
rect 3673 4933 3687 4947
rect 3693 4913 3707 4927
rect 3593 4873 3607 4887
rect 3613 4653 3627 4667
rect 3493 4433 3507 4447
rect 3473 4293 3487 4307
rect 3553 4233 3567 4247
rect 3513 4213 3527 4227
rect 3533 4153 3547 4167
rect 3493 3973 3507 3987
rect 3533 3953 3547 3967
rect 3473 3933 3487 3947
rect 3673 4453 3687 4467
rect 3733 5693 3747 5707
rect 3733 5673 3747 5687
rect 3833 6113 3847 6127
rect 3853 6113 3867 6127
rect 3893 5973 3907 5987
rect 3853 5913 3867 5927
rect 3873 5913 3887 5927
rect 3833 5873 3847 5887
rect 3793 5653 3807 5667
rect 3793 5613 3807 5627
rect 3853 5633 3867 5647
rect 3953 7753 3967 7767
rect 3993 7553 4007 7567
rect 3953 7373 3967 7387
rect 3973 7373 3987 7387
rect 4053 8433 4067 8447
rect 4053 8373 4067 8387
rect 4113 8333 4127 8347
rect 4073 8313 4087 8327
rect 4093 8213 4107 8227
rect 4033 8033 4047 8047
rect 4033 7853 4047 7867
rect 4053 7853 4067 7867
rect 4033 7713 4047 7727
rect 4053 7613 4067 7627
rect 4033 7573 4047 7587
rect 4113 7833 4127 7847
rect 4093 7813 4107 7827
rect 4013 7373 4027 7387
rect 4073 7373 4087 7387
rect 4053 7113 4067 7127
rect 4033 7013 4047 7027
rect 4053 6933 4067 6947
rect 4093 7333 4107 7347
rect 4153 8013 4167 8027
rect 4153 7873 4167 7887
rect 4133 7733 4147 7747
rect 4133 7613 4147 7627
rect 4113 7153 4127 7167
rect 4333 10833 4347 10847
rect 4573 10873 4587 10887
rect 4393 10753 4407 10767
rect 4513 10733 4527 10747
rect 4193 10713 4207 10727
rect 4313 10713 4327 10727
rect 4233 10693 4247 10707
rect 4253 10693 4267 10707
rect 4233 10673 4247 10687
rect 4333 10693 4347 10707
rect 4293 10613 4307 10627
rect 4273 10513 4287 10527
rect 4213 10453 4227 10467
rect 4193 10233 4207 10247
rect 4213 10233 4227 10247
rect 4573 10713 4587 10727
rect 4553 10653 4567 10667
rect 4473 10633 4487 10647
rect 4593 10433 4607 10447
rect 4313 10393 4327 10407
rect 4473 10393 4487 10407
rect 4573 10393 4587 10407
rect 4293 10273 4307 10287
rect 4353 10273 4367 10287
rect 4293 10253 4307 10267
rect 4253 10233 4267 10247
rect 4333 10233 4347 10247
rect 4273 10213 4287 10227
rect 4253 10173 4267 10187
rect 4253 9953 4267 9967
rect 4293 9953 4307 9967
rect 4213 9813 4227 9827
rect 4213 9753 4227 9767
rect 4253 9733 4267 9747
rect 4293 9733 4307 9747
rect 4193 9713 4207 9727
rect 4233 9713 4247 9727
rect 4273 9713 4287 9727
rect 4213 9593 4227 9607
rect 4193 9453 4207 9467
rect 4553 10233 4567 10247
rect 4513 10213 4527 10227
rect 4633 10453 4647 10467
rect 4493 10153 4507 10167
rect 4613 10153 4627 10167
rect 4573 9953 4587 9967
rect 4553 9913 4567 9927
rect 4553 9813 4567 9827
rect 4493 9793 4507 9807
rect 4513 9753 4527 9767
rect 4493 9733 4507 9747
rect 4313 9713 4327 9727
rect 4433 9653 4447 9667
rect 4533 9653 4547 9667
rect 4333 9513 4347 9527
rect 4373 9473 4387 9487
rect 4413 9473 4427 9487
rect 4293 9453 4307 9467
rect 4393 9453 4407 9467
rect 4353 9433 4367 9447
rect 4213 9353 4227 9367
rect 4333 9353 4347 9367
rect 4193 9273 4207 9287
rect 4233 9273 4247 9287
rect 4253 9273 4267 9287
rect 4213 9253 4227 9267
rect 4233 9233 4247 9247
rect 4313 8973 4327 8987
rect 4293 8953 4307 8967
rect 4273 8853 4287 8867
rect 4253 8833 4267 8847
rect 4333 8773 4347 8787
rect 4313 8753 4327 8767
rect 4413 9413 4427 9427
rect 4373 9273 4387 9287
rect 4393 9273 4407 9287
rect 4393 9173 4407 9187
rect 4533 9633 4547 9647
rect 4473 9313 4487 9327
rect 4473 9293 4487 9307
rect 4453 9273 4467 9287
rect 4513 9253 4527 9267
rect 4493 9233 4507 9247
rect 4433 8973 4447 8987
rect 4853 11213 4867 11227
rect 4673 11193 4687 11207
rect 5393 11213 5407 11227
rect 5553 11213 5567 11227
rect 5113 11173 5127 11187
rect 5293 11173 5307 11187
rect 5333 11173 5347 11187
rect 4953 11073 4967 11087
rect 5013 11073 5027 11087
rect 4693 10933 4707 10947
rect 4733 10893 4747 10907
rect 4733 10833 4747 10847
rect 5273 10933 5287 10947
rect 5333 10933 5347 10947
rect 4753 10813 4767 10827
rect 4733 10753 4747 10767
rect 4933 10913 4947 10927
rect 4953 10913 4967 10927
rect 4833 10873 4847 10887
rect 5113 10853 5127 10867
rect 4893 10813 4907 10827
rect 4813 10773 4827 10787
rect 4793 10733 4807 10747
rect 4773 10713 4787 10727
rect 4833 10733 4847 10747
rect 5313 10833 5327 10847
rect 5273 10773 5287 10787
rect 4753 10693 4767 10707
rect 4793 10693 4807 10707
rect 4833 10693 4847 10707
rect 4893 10693 4907 10707
rect 5033 10693 5047 10707
rect 5233 10713 5247 10727
rect 5293 10753 5307 10767
rect 4993 10673 5007 10687
rect 5213 10673 5227 10687
rect 5353 10753 5367 10767
rect 5253 10653 5267 10667
rect 5313 10653 5327 10667
rect 4693 10453 4707 10467
rect 4713 10453 4727 10467
rect 4673 10373 4687 10387
rect 4773 10493 4787 10507
rect 4733 10433 4747 10447
rect 4853 10473 4867 10487
rect 4873 10413 4887 10427
rect 5533 11173 5547 11187
rect 5573 11173 5587 11187
rect 6113 11213 6127 11227
rect 6493 11213 6507 11227
rect 6773 11233 6787 11247
rect 5693 11153 5707 11167
rect 5653 10933 5667 10947
rect 5493 10793 5507 10807
rect 5473 10753 5487 10767
rect 5553 10733 5567 10747
rect 5393 10693 5407 10707
rect 5373 10673 5387 10687
rect 5353 10453 5367 10467
rect 4893 10393 4907 10407
rect 5333 10433 5347 10447
rect 5113 10393 5127 10407
rect 5093 10353 5107 10367
rect 5013 10313 5027 10327
rect 4913 10293 4927 10307
rect 4813 10233 4827 10247
rect 4753 10213 4767 10227
rect 4793 10213 4807 10227
rect 5033 10193 5047 10207
rect 4913 10173 4927 10187
rect 5033 10173 5047 10187
rect 5093 10173 5107 10187
rect 4713 9993 4727 10007
rect 4873 10013 4887 10027
rect 4673 9953 4687 9967
rect 4733 9953 4747 9967
rect 4673 9873 4687 9887
rect 4833 9773 4847 9787
rect 4673 9753 4687 9767
rect 4753 9753 4767 9767
rect 4793 9753 4807 9767
rect 4653 9733 4667 9747
rect 4573 9493 4587 9507
rect 4553 9473 4567 9487
rect 4613 9473 4627 9487
rect 4633 9453 4647 9467
rect 4593 9433 4607 9447
rect 4553 9233 4567 9247
rect 4613 9193 4627 9207
rect 4533 9073 4547 9087
rect 4513 8973 4527 8987
rect 4553 8953 4567 8967
rect 4513 8933 4527 8947
rect 4573 8933 4587 8947
rect 4373 8873 4387 8887
rect 4433 8853 4447 8867
rect 4353 8733 4367 8747
rect 4333 8633 4347 8647
rect 4293 8593 4307 8607
rect 4333 8573 4347 8587
rect 4193 8513 4207 8527
rect 4293 8513 4307 8527
rect 4353 8493 4367 8507
rect 4413 8493 4427 8507
rect 4293 8453 4307 8467
rect 4313 8453 4327 8467
rect 4333 8393 4347 8407
rect 4293 8373 4307 8387
rect 4233 8313 4247 8327
rect 4253 8313 4267 8327
rect 4193 8213 4207 8227
rect 4233 8133 4247 8147
rect 4193 7993 4207 8007
rect 4233 7973 4247 7987
rect 4273 8153 4287 8167
rect 4313 8353 4327 8367
rect 4373 8313 4387 8327
rect 4353 8293 4367 8307
rect 4373 8093 4387 8107
rect 4393 8093 4407 8107
rect 4293 8073 4307 8087
rect 4273 8033 4287 8047
rect 4253 7873 4267 7887
rect 4233 7833 4247 7847
rect 4253 7813 4267 7827
rect 4193 7793 4207 7807
rect 4253 7773 4267 7787
rect 4153 7573 4167 7587
rect 4353 8053 4367 8067
rect 4313 7993 4327 8007
rect 4353 7793 4367 7807
rect 4313 7753 4327 7767
rect 4353 7633 4367 7647
rect 4293 7613 4307 7627
rect 4313 7553 4327 7567
rect 4193 7473 4207 7487
rect 4193 7353 4207 7367
rect 4133 7033 4147 7047
rect 4073 6913 4087 6927
rect 4073 6893 4087 6907
rect 4093 6873 4107 6887
rect 4033 6813 4047 6827
rect 4113 6793 4127 6807
rect 4033 6573 4047 6587
rect 4133 6573 4147 6587
rect 4113 6553 4127 6567
rect 4133 6433 4147 6447
rect 4073 6413 4087 6427
rect 4093 6413 4107 6427
rect 3993 6353 4007 6367
rect 3973 6113 3987 6127
rect 4093 6373 4107 6387
rect 4013 6173 4027 6187
rect 4213 7333 4227 7347
rect 4193 7213 4207 7227
rect 4173 6773 4187 6787
rect 4173 6153 4187 6167
rect 4153 6113 4167 6127
rect 4093 6033 4107 6047
rect 4153 6073 4167 6087
rect 4293 7353 4307 7367
rect 4313 7053 4327 7067
rect 4293 7033 4307 7047
rect 4273 7013 4287 7027
rect 4253 6993 4267 7007
rect 4253 6913 4267 6927
rect 4193 6033 4207 6047
rect 4113 5993 4127 6007
rect 4093 5933 4107 5947
rect 3993 5873 4007 5887
rect 3953 5713 3967 5727
rect 4053 5713 4067 5727
rect 3913 5673 3927 5687
rect 3813 5593 3827 5607
rect 3753 5573 3767 5587
rect 3733 5393 3747 5407
rect 3913 5613 3927 5627
rect 3953 5613 3967 5627
rect 3933 5533 3947 5547
rect 3893 5513 3907 5527
rect 3833 5453 3847 5467
rect 4033 5613 4047 5627
rect 3993 5433 4007 5447
rect 3793 5413 3807 5427
rect 3753 5193 3767 5207
rect 3773 5153 3787 5167
rect 3953 5413 3967 5427
rect 3993 5413 4007 5427
rect 3913 5373 3927 5387
rect 3893 5113 3907 5127
rect 4233 5693 4247 5707
rect 4153 5553 4167 5567
rect 4133 5473 4147 5487
rect 4113 5433 4127 5447
rect 3813 5073 3827 5087
rect 4053 5073 4067 5087
rect 3793 4913 3807 4927
rect 3753 4693 3767 4707
rect 3793 4473 3807 4487
rect 3613 4153 3627 4167
rect 3733 4273 3747 4287
rect 3773 4193 3787 4207
rect 3713 4173 3727 4187
rect 3693 4113 3707 4127
rect 3713 4013 3727 4027
rect 3633 3993 3647 4007
rect 3593 3913 3607 3927
rect 3733 3993 3747 4007
rect 3653 3973 3667 3987
rect 3793 3933 3807 3947
rect 3693 3913 3707 3927
rect 3633 3813 3647 3827
rect 3593 3713 3607 3727
rect 3433 3593 3447 3607
rect 3453 3593 3467 3607
rect 3653 3693 3667 3707
rect 3793 3593 3807 3607
rect 3673 3553 3687 3567
rect 3393 3533 3407 3547
rect 3613 3533 3627 3547
rect 3373 3493 3387 3507
rect 3293 3133 3307 3147
rect 3373 3233 3387 3247
rect 3573 3233 3587 3247
rect 3633 3453 3647 3467
rect 3613 3233 3627 3247
rect 3353 3193 3367 3207
rect 3593 3213 3607 3227
rect 4113 5053 4127 5067
rect 4173 5433 4187 5447
rect 4213 5433 4227 5447
rect 4193 5373 4207 5387
rect 4213 5313 4227 5327
rect 4153 5233 4167 5247
rect 4153 5033 4167 5047
rect 4213 5033 4227 5047
rect 4133 4993 4147 5007
rect 4073 4973 4087 4987
rect 3993 4953 4007 4967
rect 4113 4953 4127 4967
rect 3873 4933 3887 4947
rect 3913 4933 3927 4947
rect 3873 4913 3887 4927
rect 3873 4753 3887 4767
rect 3933 4693 3947 4707
rect 3973 4673 3987 4687
rect 3833 4653 3847 4667
rect 3833 4633 3847 4647
rect 3833 4493 3847 4507
rect 3893 4653 3907 4667
rect 3953 4613 3967 4627
rect 3853 4473 3867 4487
rect 3913 4433 3927 4447
rect 3873 4253 3887 4267
rect 3853 4193 3867 4207
rect 3833 3853 3847 3867
rect 3873 4173 3887 4187
rect 4093 4933 4107 4947
rect 4193 4933 4207 4947
rect 4133 4873 4147 4887
rect 4333 6913 4347 6927
rect 4353 6893 4367 6907
rect 4353 6873 4367 6887
rect 4293 6853 4307 6867
rect 4333 6813 4347 6827
rect 4333 6733 4347 6747
rect 4313 6513 4327 6527
rect 4293 6413 4307 6427
rect 4293 6073 4307 6087
rect 4293 6053 4307 6067
rect 4273 5953 4287 5967
rect 4253 5433 4267 5447
rect 4273 5413 4287 5427
rect 4353 6573 4367 6587
rect 4353 6413 4367 6427
rect 4473 8793 4487 8807
rect 4573 8793 4587 8807
rect 4513 8773 4527 8787
rect 4553 8773 4567 8787
rect 4553 8753 4567 8767
rect 4593 8753 4607 8767
rect 4813 9733 4827 9747
rect 4773 9473 4787 9487
rect 4733 9413 4747 9427
rect 4813 9493 4827 9507
rect 4833 9473 4847 9487
rect 4853 9413 4867 9427
rect 4853 9333 4867 9347
rect 4793 9293 4807 9307
rect 4793 9273 4807 9287
rect 4693 9233 4707 9247
rect 4753 9213 4767 9227
rect 4753 9013 4767 9027
rect 4713 8993 4727 9007
rect 4793 8993 4807 9007
rect 4833 8993 4847 9007
rect 4693 8973 4707 8987
rect 4673 8713 4687 8727
rect 4553 8633 4567 8647
rect 4513 8593 4527 8607
rect 4673 8593 4687 8607
rect 4553 8513 4567 8527
rect 4493 8353 4507 8367
rect 4513 8353 4527 8367
rect 4493 8313 4507 8327
rect 4573 8493 4587 8507
rect 4533 8293 4547 8307
rect 4693 8473 4707 8487
rect 4673 8453 4687 8467
rect 4633 8293 4647 8307
rect 4473 8273 4487 8287
rect 4553 8173 4567 8187
rect 4433 8053 4447 8067
rect 4433 7993 4447 8007
rect 4513 7993 4527 8007
rect 4413 7973 4427 7987
rect 4393 7533 4407 7547
rect 4393 7353 4407 7367
rect 4393 7053 4407 7067
rect 4373 6253 4387 6267
rect 4373 6233 4387 6247
rect 4353 6073 4367 6087
rect 4373 5953 4387 5967
rect 4453 7813 4467 7827
rect 4433 7793 4447 7807
rect 4433 7633 4447 7647
rect 4473 7553 4487 7567
rect 4453 7533 4467 7547
rect 4433 7493 4447 7507
rect 4453 6993 4467 7007
rect 4433 6953 4447 6967
rect 4433 6893 4447 6907
rect 4413 6853 4427 6867
rect 4393 5853 4407 5867
rect 4333 5693 4347 5707
rect 4393 5673 4407 5687
rect 4353 5633 4367 5647
rect 4333 5613 4347 5627
rect 4313 5533 4327 5547
rect 4433 5833 4447 5847
rect 4613 8273 4627 8287
rect 4653 8273 4667 8287
rect 4633 8253 4647 8267
rect 4573 8073 4587 8087
rect 4633 8073 4647 8087
rect 4633 7993 4647 8007
rect 4613 7673 4627 7687
rect 4613 7593 4627 7607
rect 4553 7573 4567 7587
rect 4573 7573 4587 7587
rect 4533 7533 4547 7547
rect 4553 7533 4567 7547
rect 4593 7513 4607 7527
rect 4593 7433 4607 7447
rect 4513 7093 4527 7107
rect 4513 7073 4527 7087
rect 4493 6993 4507 7007
rect 4493 6933 4507 6947
rect 4513 6873 4527 6887
rect 4493 6853 4507 6867
rect 4473 6713 4487 6727
rect 4473 6613 4487 6627
rect 4553 6853 4567 6867
rect 4633 7053 4647 7067
rect 4613 6873 4627 6887
rect 4673 8253 4687 8267
rect 4773 8973 4787 8987
rect 4813 8973 4827 8987
rect 4793 8953 4807 8967
rect 4753 8813 4767 8827
rect 4813 8813 4827 8827
rect 4733 8753 4747 8767
rect 4753 8713 4767 8727
rect 4733 8273 4747 8287
rect 4713 8253 4727 8267
rect 4693 7993 4707 8007
rect 4693 7793 4707 7807
rect 4733 7693 4747 7707
rect 4733 7673 4747 7687
rect 4693 7613 4707 7627
rect 4833 8773 4847 8787
rect 4833 8733 4847 8747
rect 4773 8553 4787 8567
rect 4813 8553 4827 8567
rect 4893 9773 4907 9787
rect 4973 9973 4987 9987
rect 5013 9953 5027 9967
rect 4933 9933 4947 9947
rect 4953 9913 4967 9927
rect 5013 9833 5027 9847
rect 4993 9753 5007 9767
rect 5073 9753 5087 9767
rect 4993 9713 5007 9727
rect 5033 9713 5047 9727
rect 5273 10213 5287 10227
rect 5253 10193 5267 10207
rect 5293 10173 5307 10187
rect 5153 9953 5167 9967
rect 5193 9953 5207 9967
rect 5133 9673 5147 9687
rect 4993 9473 5007 9487
rect 5073 9473 5087 9487
rect 4913 9453 4927 9467
rect 4893 9373 4907 9387
rect 4953 9293 4967 9307
rect 4953 9193 4967 9207
rect 4933 9173 4947 9187
rect 4893 9153 4907 9167
rect 4913 8793 4927 8807
rect 4793 8533 4807 8547
rect 4873 8533 4887 8547
rect 4773 8513 4787 8527
rect 4753 7593 4767 7607
rect 4813 8513 4827 8527
rect 4853 8513 4867 8527
rect 4833 8473 4847 8487
rect 4833 8453 4847 8467
rect 4873 8353 4887 8367
rect 4813 8293 4827 8307
rect 4853 8253 4867 8267
rect 4973 9113 4987 9127
rect 4953 8973 4967 8987
rect 5053 9453 5067 9467
rect 5133 9453 5147 9467
rect 5033 9013 5047 9027
rect 5073 8993 5087 9007
rect 5053 8973 5067 8987
rect 5013 8953 5027 8967
rect 4973 8773 4987 8787
rect 4973 8533 4987 8547
rect 4953 8513 4967 8527
rect 4933 8493 4947 8507
rect 4933 8393 4947 8407
rect 4913 8353 4927 8367
rect 4933 8293 4947 8307
rect 4953 8213 4967 8227
rect 4853 8153 4867 8167
rect 4893 8153 4907 8167
rect 4833 8033 4847 8047
rect 4793 7593 4807 7607
rect 4773 7553 4787 7567
rect 4793 7553 4807 7567
rect 4693 7513 4707 7527
rect 4773 7493 4787 7507
rect 4793 7493 4807 7507
rect 4673 7473 4687 7487
rect 4673 7453 4687 7467
rect 4693 7373 4707 7387
rect 4733 7293 4747 7307
rect 4693 7073 4707 7087
rect 4733 7073 4747 7087
rect 4773 7073 4787 7087
rect 4713 7053 4727 7067
rect 4733 7033 4747 7047
rect 4713 6853 4727 6867
rect 4653 6833 4667 6847
rect 4613 6813 4627 6827
rect 4653 6813 4667 6827
rect 4533 6793 4547 6807
rect 4573 6793 4587 6807
rect 4593 6793 4607 6807
rect 4533 6693 4547 6707
rect 4513 6593 4527 6607
rect 4473 6573 4487 6587
rect 4493 6573 4507 6587
rect 4613 6693 4627 6707
rect 4573 6573 4587 6587
rect 4553 6553 4567 6567
rect 4633 6573 4647 6587
rect 4553 6493 4567 6507
rect 4593 6493 4607 6507
rect 4593 6473 4607 6487
rect 4533 6373 4547 6387
rect 4573 6353 4587 6367
rect 4473 6293 4487 6307
rect 4633 6213 4647 6227
rect 4573 6153 4587 6167
rect 4533 5953 4547 5967
rect 4573 5933 4587 5947
rect 4633 6133 4647 6147
rect 4613 6113 4627 6127
rect 4633 6073 4647 6087
rect 4613 6053 4627 6067
rect 4553 5893 4567 5907
rect 4593 5893 4607 5907
rect 4553 5673 4567 5687
rect 4573 5553 4587 5567
rect 4453 5513 4467 5527
rect 4573 5513 4587 5527
rect 4413 5473 4427 5487
rect 4313 5433 4327 5447
rect 4253 5393 4267 5407
rect 4253 4973 4267 4987
rect 4293 5133 4307 5147
rect 4233 4793 4247 4807
rect 4073 4673 4087 4687
rect 4353 5133 4367 5147
rect 4393 5133 4407 5147
rect 4373 5113 4387 5127
rect 4413 5113 4427 5127
rect 4453 5093 4467 5107
rect 4313 5033 4327 5047
rect 4313 5013 4327 5027
rect 4333 4993 4347 5007
rect 4293 4813 4307 4827
rect 4253 4633 4267 4647
rect 4273 4633 4287 4647
rect 4093 4613 4107 4627
rect 4033 4593 4047 4607
rect 3993 4473 4007 4487
rect 3933 4173 3947 4187
rect 3973 4173 3987 4187
rect 4153 4553 4167 4567
rect 4233 4553 4247 4567
rect 4093 4473 4107 4487
rect 4133 4473 4147 4487
rect 4173 4473 4187 4487
rect 4193 4473 4207 4487
rect 4113 4433 4127 4447
rect 4133 4213 4147 4227
rect 3913 4153 3927 4167
rect 3853 3753 3867 3767
rect 3893 3753 3907 3767
rect 3973 4153 3987 4167
rect 3953 4013 3967 4027
rect 4173 4033 4187 4047
rect 4073 3833 4087 3847
rect 4033 3813 4047 3827
rect 3873 3693 3887 3707
rect 3813 3573 3827 3587
rect 3853 3533 3867 3547
rect 3913 3533 3927 3547
rect 3873 3493 3887 3507
rect 3793 3293 3807 3307
rect 3713 3233 3727 3247
rect 3633 3213 3647 3227
rect 3553 3173 3567 3187
rect 3613 3173 3627 3187
rect 3393 3133 3407 3147
rect 3333 3093 3347 3107
rect 3273 3053 3287 3067
rect 3313 3053 3327 3067
rect 3233 3013 3247 3027
rect 3253 3013 3267 3027
rect 3293 2973 3307 2987
rect 3313 2833 3327 2847
rect 3213 2713 3227 2727
rect 3353 3073 3367 3087
rect 3353 3013 3367 3027
rect 3533 3053 3547 3067
rect 3813 3053 3827 3067
rect 3393 2993 3407 3007
rect 3413 2973 3427 2987
rect 3373 2773 3387 2787
rect 3333 2713 3347 2727
rect 3313 2693 3327 2707
rect 3313 2633 3327 2647
rect 3273 2553 3287 2567
rect 3333 2613 3347 2627
rect 3233 2533 3247 2547
rect 3293 2473 3307 2487
rect 3293 2453 3307 2467
rect 3393 2333 3407 2347
rect 3293 2293 3307 2307
rect 3313 2293 3327 2307
rect 3353 2293 3367 2307
rect 3233 2273 3247 2287
rect 3273 2233 3287 2247
rect 3293 2113 3307 2127
rect 3273 1833 3287 1847
rect 3233 1773 3247 1787
rect 3193 1753 3207 1767
rect 3193 1733 3207 1747
rect 3073 1573 3087 1587
rect 2953 1553 2967 1567
rect 3013 1553 3027 1567
rect 2953 1533 2967 1547
rect 2933 833 2947 847
rect 2993 1253 3007 1267
rect 2973 1113 2987 1127
rect 2953 613 2967 627
rect 2873 593 2887 607
rect 2973 553 2987 567
rect 2713 173 2727 187
rect 2473 133 2487 147
rect 2593 133 2607 147
rect 2793 373 2807 387
rect 2933 373 2947 387
rect 3113 1433 3127 1447
rect 3153 1433 3167 1447
rect 3093 1333 3107 1347
rect 3013 1233 3027 1247
rect 3053 1133 3067 1147
rect 3073 1113 3087 1127
rect 3033 1093 3047 1107
rect 3073 1093 3087 1107
rect 3133 1093 3147 1107
rect 3133 1073 3147 1087
rect 3013 1053 3027 1067
rect 3093 873 3107 887
rect 3033 813 3047 827
rect 3073 813 3087 827
rect 3013 793 3027 807
rect 3033 793 3047 807
rect 3053 793 3067 807
rect 3013 693 3027 707
rect 3073 633 3087 647
rect 3113 813 3127 827
rect 3053 393 3067 407
rect 2773 333 2787 347
rect 3013 353 3027 367
rect 2953 213 2967 227
rect 2933 193 2947 207
rect 2973 173 2987 187
rect 3233 1613 3247 1627
rect 3213 1353 3227 1367
rect 3173 1333 3187 1347
rect 3193 1333 3207 1347
rect 3173 1193 3187 1207
rect 3173 833 3187 847
rect 3393 2133 3407 2147
rect 3313 2093 3327 2107
rect 3333 2073 3347 2087
rect 3593 2773 3607 2787
rect 3433 2753 3447 2767
rect 3633 2753 3647 2767
rect 3733 2753 3747 2767
rect 3493 2733 3507 2747
rect 3533 2713 3547 2727
rect 3513 2613 3527 2627
rect 3713 2613 3727 2627
rect 3553 2593 3567 2607
rect 3453 2573 3467 2587
rect 3433 2273 3447 2287
rect 3433 2093 3447 2107
rect 3353 2033 3367 2047
rect 3413 2033 3427 2047
rect 3353 1773 3367 1787
rect 3393 1753 3407 1767
rect 3353 1593 3367 1607
rect 3333 1553 3347 1567
rect 3313 1333 3327 1347
rect 3293 1293 3307 1307
rect 3333 1293 3347 1307
rect 3273 1273 3287 1287
rect 3333 1273 3347 1287
rect 3233 1213 3247 1227
rect 3293 1133 3307 1147
rect 3233 1093 3247 1107
rect 3273 1093 3287 1107
rect 3213 913 3227 927
rect 3193 813 3207 827
rect 3173 793 3187 807
rect 3153 773 3167 787
rect 3393 1093 3407 1107
rect 3313 1033 3327 1047
rect 3393 953 3407 967
rect 3273 833 3287 847
rect 3313 833 3327 847
rect 3293 813 3307 827
rect 3253 793 3267 807
rect 3333 773 3347 787
rect 3273 653 3287 667
rect 3333 653 3347 667
rect 3213 633 3227 647
rect 3313 633 3327 647
rect 3293 593 3307 607
rect 3173 413 3187 427
rect 3133 373 3147 387
rect 3153 173 3167 187
rect 3253 373 3267 387
rect 3213 353 3227 367
rect 3193 333 3207 347
rect 3233 333 3247 347
rect 3273 293 3287 307
rect 3613 2213 3627 2227
rect 3613 2193 3627 2207
rect 3573 2033 3587 2047
rect 3493 1793 3507 1807
rect 3473 1773 3487 1787
rect 3493 1593 3507 1607
rect 3553 1713 3567 1727
rect 3633 2033 3647 2047
rect 3593 1873 3607 1887
rect 3653 1873 3667 1887
rect 3573 1633 3587 1647
rect 3553 1613 3567 1627
rect 3593 1593 3607 1607
rect 3513 1433 3527 1447
rect 3613 1433 3627 1447
rect 3513 1333 3527 1347
rect 3493 1293 3507 1307
rect 3573 1293 3587 1307
rect 3533 1253 3547 1267
rect 3513 1213 3527 1227
rect 3553 1213 3567 1227
rect 3553 1173 3567 1187
rect 3573 1173 3587 1187
rect 3493 1153 3507 1167
rect 3473 633 3487 647
rect 3573 1113 3587 1127
rect 3633 1313 3647 1327
rect 3553 1093 3567 1107
rect 3613 1093 3627 1107
rect 3513 1073 3527 1087
rect 3533 1073 3547 1087
rect 3553 1013 3567 1027
rect 3533 813 3547 827
rect 3513 793 3527 807
rect 3573 773 3587 787
rect 3533 653 3547 667
rect 3553 633 3567 647
rect 3533 613 3547 627
rect 3633 613 3647 627
rect 3473 373 3487 387
rect 3413 173 3427 187
rect 3453 173 3467 187
rect 3113 153 3127 167
rect 3193 153 3207 167
rect 3493 313 3507 327
rect 2213 93 2227 107
rect 2693 93 2707 107
rect 3053 93 3067 107
rect 3473 153 3487 167
rect 3733 2533 3747 2547
rect 3733 2273 3747 2287
rect 3873 2533 3887 2547
rect 3813 2513 3827 2527
rect 3773 2333 3787 2347
rect 3793 2333 3807 2347
rect 3753 2253 3767 2267
rect 3813 2273 3827 2287
rect 3853 2213 3867 2227
rect 3813 2113 3827 2127
rect 3893 2313 3907 2327
rect 3873 2193 3887 2207
rect 3933 3233 3947 3247
rect 3933 2753 3947 2767
rect 3973 3453 3987 3467
rect 3953 2673 3967 2687
rect 4033 3073 4047 3087
rect 3993 3053 4007 3067
rect 3993 3013 4007 3027
rect 3973 2553 3987 2567
rect 3973 2353 3987 2367
rect 4013 2793 4027 2807
rect 4053 2593 4067 2607
rect 4113 3753 4127 3767
rect 4133 3693 4147 3707
rect 4173 3693 4187 3707
rect 4153 3673 4167 3687
rect 4093 3653 4107 3667
rect 4153 3653 4167 3667
rect 4093 3533 4107 3547
rect 4113 3533 4127 3547
rect 4133 3513 4147 3527
rect 4093 3473 4107 3487
rect 4153 3473 4167 3487
rect 4253 4213 4267 4227
rect 4273 4213 4287 4227
rect 4213 3953 4227 3967
rect 4233 3733 4247 3747
rect 4213 3513 4227 3527
rect 4193 3453 4207 3467
rect 4113 3253 4127 3267
rect 4313 4773 4327 4787
rect 4293 3973 4307 3987
rect 4313 3833 4327 3847
rect 4273 3773 4287 3787
rect 4253 3193 4267 3207
rect 4153 3153 4167 3167
rect 4173 3153 4187 3167
rect 4413 4893 4427 4907
rect 4433 4873 4447 4887
rect 4413 4653 4427 4667
rect 4373 4633 4387 4647
rect 4373 4513 4387 4527
rect 4413 4513 4427 4527
rect 4413 4473 4427 4487
rect 4353 4453 4367 4467
rect 4433 4273 4447 4287
rect 4473 5073 4487 5087
rect 4493 5033 4507 5047
rect 4513 5033 4527 5047
rect 4473 4453 4487 4467
rect 4453 4233 4467 4247
rect 4393 4213 4407 4227
rect 4433 4193 4447 4207
rect 4473 4193 4487 4207
rect 4453 4173 4467 4187
rect 4353 4133 4367 4147
rect 4333 3753 4347 3767
rect 4313 3733 4327 3747
rect 4473 3993 4487 4007
rect 4433 3973 4447 3987
rect 4413 3953 4427 3967
rect 4413 3853 4427 3867
rect 4373 3713 4387 3727
rect 4493 3873 4507 3887
rect 4493 3713 4507 3727
rect 4453 3693 4467 3707
rect 4373 3673 4387 3687
rect 4413 3673 4427 3687
rect 4333 3433 4347 3447
rect 4413 3493 4427 3507
rect 4433 3433 4447 3447
rect 4293 3113 4307 3127
rect 4373 3113 4387 3127
rect 4333 3073 4347 3087
rect 4253 3033 4267 3047
rect 4233 3013 4247 3027
rect 4213 2793 4227 2807
rect 4093 2753 4107 2767
rect 4233 2753 4247 2767
rect 4073 2573 4087 2587
rect 4273 2733 4287 2747
rect 4293 2633 4307 2647
rect 4253 2573 4267 2587
rect 4033 2533 4047 2547
rect 4073 2533 4087 2547
rect 4393 3053 4407 3067
rect 4413 2673 4427 2687
rect 4413 2613 4427 2627
rect 4253 2513 4267 2527
rect 4353 2533 4367 2547
rect 4393 2533 4407 2547
rect 4313 2493 4327 2507
rect 3913 2293 3927 2307
rect 3993 2293 4007 2307
rect 4073 2333 4087 2347
rect 4073 2293 4087 2307
rect 3933 2273 3947 2287
rect 3973 2273 3987 2287
rect 4013 2273 4027 2287
rect 4033 2273 4047 2287
rect 4113 2273 4127 2287
rect 3933 2233 3947 2247
rect 3993 2253 4007 2267
rect 3993 2233 4007 2247
rect 3953 2073 3967 2087
rect 3833 2053 3847 2067
rect 3793 2033 3807 2047
rect 3913 2053 3927 2067
rect 3973 2053 3987 2067
rect 3933 2033 3947 2047
rect 4233 2213 4247 2227
rect 4273 2173 4287 2187
rect 4053 1853 4067 1867
rect 4013 1813 4027 1827
rect 3873 1793 3887 1807
rect 3933 1793 3947 1807
rect 3973 1793 3987 1807
rect 3713 1773 3727 1787
rect 3853 1653 3867 1667
rect 3753 1633 3767 1647
rect 3673 1613 3687 1627
rect 3673 1153 3687 1167
rect 3733 993 3747 1007
rect 3813 1593 3827 1607
rect 3873 1593 3887 1607
rect 3773 1333 3787 1347
rect 3793 1313 3807 1327
rect 3793 1113 3807 1127
rect 3813 1073 3827 1087
rect 3953 1773 3967 1787
rect 3993 1773 4007 1787
rect 4273 2093 4287 2107
rect 4373 2093 4387 2107
rect 4293 1913 4307 1927
rect 4193 1793 4207 1807
rect 4233 1793 4247 1807
rect 4073 1773 4087 1787
rect 3953 1733 3967 1747
rect 4193 1693 4207 1707
rect 3993 1653 4007 1667
rect 3933 1313 3947 1327
rect 4053 1613 4067 1627
rect 4073 1613 4087 1627
rect 4253 1773 4267 1787
rect 4593 5413 4607 5427
rect 4633 5433 4647 5447
rect 4613 5373 4627 5387
rect 4613 5193 4627 5207
rect 4613 5153 4627 5167
rect 4593 5073 4607 5087
rect 4593 5013 4607 5027
rect 4573 4973 4587 4987
rect 4573 4953 4587 4967
rect 4633 4953 4647 4967
rect 4613 4913 4627 4927
rect 4593 4833 4607 4847
rect 4693 6693 4707 6707
rect 4673 6633 4687 6647
rect 4673 6493 4687 6507
rect 4713 6673 4727 6687
rect 4713 6653 4727 6667
rect 4713 6553 4727 6567
rect 4713 6533 4727 6547
rect 4693 5953 4707 5967
rect 4673 5893 4687 5907
rect 4693 5853 4707 5867
rect 4673 5413 4687 5427
rect 4653 4733 4667 4747
rect 4633 4693 4647 4707
rect 4553 4633 4567 4647
rect 4533 4453 4547 4467
rect 4613 4533 4627 4547
rect 4633 4493 4647 4507
rect 4653 4473 4667 4487
rect 4753 7013 4767 7027
rect 5133 9233 5147 9247
rect 5113 9013 5127 9027
rect 5093 8853 5107 8867
rect 5093 8753 5107 8767
rect 5053 8633 5067 8647
rect 5133 8993 5147 9007
rect 5113 8573 5127 8587
rect 5013 8493 5027 8507
rect 4993 8433 5007 8447
rect 5013 8393 5027 8407
rect 4993 8193 5007 8207
rect 5093 8493 5107 8507
rect 5133 8493 5147 8507
rect 5113 8433 5127 8447
rect 5073 8353 5087 8367
rect 5033 8313 5047 8327
rect 5073 8313 5087 8327
rect 5313 10013 5327 10027
rect 5313 9973 5327 9987
rect 5293 9833 5307 9847
rect 5253 9813 5267 9827
rect 5253 9773 5267 9787
rect 5293 9753 5307 9767
rect 5173 9733 5187 9747
rect 5473 10713 5487 10727
rect 5553 10713 5567 10727
rect 5633 10713 5647 10727
rect 5453 10673 5467 10687
rect 5513 10693 5527 10707
rect 5533 10673 5547 10687
rect 5493 10633 5507 10647
rect 5513 10453 5527 10467
rect 5553 10453 5567 10467
rect 5493 10413 5507 10427
rect 5593 10433 5607 10447
rect 5473 10193 5487 10207
rect 5453 10173 5467 10187
rect 5413 9973 5427 9987
rect 5433 9973 5447 9987
rect 5473 9953 5487 9967
rect 5373 9773 5387 9787
rect 5353 9733 5367 9747
rect 5273 9713 5287 9727
rect 5273 9653 5287 9667
rect 5293 9453 5307 9467
rect 5173 9253 5187 9267
rect 5213 9253 5227 9267
rect 5253 9253 5267 9267
rect 5193 9233 5207 9247
rect 5233 9233 5247 9247
rect 5253 9213 5267 9227
rect 5313 9433 5327 9447
rect 5333 9233 5347 9247
rect 5173 9113 5187 9127
rect 5273 9113 5287 9127
rect 5293 9113 5307 9127
rect 5313 8993 5327 9007
rect 5453 9793 5467 9807
rect 5433 9473 5447 9487
rect 5673 10913 5687 10927
rect 6133 11173 6147 11187
rect 5913 11153 5927 11167
rect 5793 11113 5807 11127
rect 6273 11153 6287 11167
rect 6333 11153 6347 11167
rect 6013 10933 6027 10947
rect 6053 10933 6067 10947
rect 5573 10393 5587 10407
rect 5533 10353 5547 10367
rect 5573 10253 5587 10267
rect 5553 10193 5567 10207
rect 5513 10173 5527 10187
rect 5513 9793 5527 9807
rect 5593 10233 5607 10247
rect 5613 10193 5627 10207
rect 5593 9953 5607 9967
rect 5573 9773 5587 9787
rect 5513 9733 5527 9747
rect 5513 9473 5527 9487
rect 5513 9393 5527 9407
rect 5493 9273 5507 9287
rect 5393 9113 5407 9127
rect 5373 9013 5387 9027
rect 5213 8853 5227 8867
rect 5253 8793 5267 8807
rect 5193 8773 5207 8787
rect 5233 8773 5247 8787
rect 5173 8653 5187 8667
rect 5213 8553 5227 8567
rect 5173 8333 5187 8347
rect 5033 8233 5047 8247
rect 5133 8273 5147 8287
rect 5093 8213 5107 8227
rect 5053 8033 5067 8047
rect 5093 8033 5107 8047
rect 5013 7973 5027 7987
rect 4973 7853 4987 7867
rect 4933 7813 4947 7827
rect 5053 7833 5067 7847
rect 4973 7793 4987 7807
rect 4993 7693 5007 7707
rect 5053 7693 5067 7707
rect 4933 7633 4947 7647
rect 4873 7593 4887 7607
rect 4853 7393 4867 7407
rect 4833 7353 4847 7367
rect 4813 7113 4827 7127
rect 4813 7073 4827 7087
rect 4973 7573 4987 7587
rect 4933 7513 4947 7527
rect 5113 8013 5127 8027
rect 5093 7973 5107 7987
rect 5073 7573 5087 7587
rect 5033 7553 5047 7567
rect 5073 7553 5087 7567
rect 5053 7513 5067 7527
rect 4973 7433 4987 7447
rect 4913 7353 4927 7367
rect 4953 7353 4967 7367
rect 5073 7373 5087 7387
rect 4893 7333 4907 7347
rect 4933 7333 4947 7347
rect 4973 7333 4987 7347
rect 4993 7333 5007 7347
rect 4933 7313 4947 7327
rect 4913 7293 4927 7307
rect 4893 7273 4907 7287
rect 4893 7053 4907 7067
rect 4853 7033 4867 7047
rect 4873 7033 4887 7047
rect 4833 6873 4847 6887
rect 4773 6853 4787 6867
rect 4813 6853 4827 6867
rect 4853 6853 4867 6867
rect 4753 6453 4767 6467
rect 4773 6453 4787 6467
rect 4733 5993 4747 6007
rect 4793 6433 4807 6447
rect 4873 6773 4887 6787
rect 4933 7273 4947 7287
rect 4933 7113 4947 7127
rect 4933 6993 4947 7007
rect 5093 7353 5107 7367
rect 5073 7313 5087 7327
rect 5013 7193 5027 7207
rect 5073 7193 5087 7207
rect 5053 7133 5067 7147
rect 4993 7073 5007 7087
rect 5033 7053 5047 7067
rect 4973 7013 4987 7027
rect 5073 7053 5087 7067
rect 5133 7833 5147 7847
rect 5193 8033 5207 8047
rect 5193 7853 5207 7867
rect 5133 7733 5147 7747
rect 5173 7673 5187 7687
rect 5193 7633 5207 7647
rect 5173 7533 5187 7547
rect 5153 7373 5167 7387
rect 5233 8493 5247 8507
rect 5273 8473 5287 8487
rect 5253 8173 5267 8187
rect 5273 8153 5287 8167
rect 5273 8113 5287 8127
rect 5273 8033 5287 8047
rect 5253 7933 5267 7947
rect 5253 7653 5267 7667
rect 5313 8953 5327 8967
rect 5373 8833 5387 8847
rect 5353 8593 5367 8607
rect 5473 9253 5487 9267
rect 5473 8973 5487 8987
rect 5413 8953 5427 8967
rect 5413 8793 5427 8807
rect 5433 8793 5447 8807
rect 5393 8513 5407 8527
rect 5353 8473 5367 8487
rect 5313 8293 5327 8307
rect 5373 8273 5387 8287
rect 5353 8253 5367 8267
rect 5313 8033 5327 8047
rect 5353 8033 5367 8047
rect 5313 7933 5327 7947
rect 5493 8613 5507 8627
rect 5493 8533 5507 8547
rect 5433 8513 5447 8527
rect 5553 9453 5567 9467
rect 5533 9293 5547 9307
rect 5593 9513 5607 9527
rect 5593 9433 5607 9447
rect 5733 10913 5747 10927
rect 5693 10413 5707 10427
rect 5973 10913 5987 10927
rect 5773 10853 5787 10867
rect 6053 10893 6067 10907
rect 6273 10933 6287 10947
rect 6733 11193 6747 11207
rect 7013 11293 7027 11307
rect 6973 11193 6987 11207
rect 6433 11133 6447 11147
rect 6513 11173 6527 11187
rect 6733 11173 6747 11187
rect 6773 11173 6787 11187
rect 6973 11173 6987 11187
rect 6753 11153 6767 11167
rect 6993 11153 7007 11167
rect 6713 11133 6727 11147
rect 6953 11133 6967 11147
rect 6473 11113 6487 11127
rect 6213 10873 6227 10887
rect 6033 10833 6047 10847
rect 5993 10813 6007 10827
rect 6253 10893 6267 10907
rect 6273 10833 6287 10847
rect 5953 10753 5967 10767
rect 6233 10753 6247 10767
rect 5793 10733 5807 10747
rect 6073 10733 6087 10747
rect 5753 10713 5767 10727
rect 6033 10713 6047 10727
rect 5813 10693 5827 10707
rect 6033 10693 6047 10707
rect 5773 10673 5787 10687
rect 6053 10673 6067 10687
rect 6013 10653 6027 10667
rect 5973 10453 5987 10467
rect 6093 10433 6107 10447
rect 6013 10413 6027 10427
rect 5833 10393 5847 10407
rect 5973 10393 5987 10407
rect 5893 10333 5907 10347
rect 6013 10333 6027 10347
rect 5733 10253 5747 10267
rect 5753 10233 5767 10247
rect 5853 10233 5867 10247
rect 5733 10213 5747 10227
rect 5813 10213 5827 10227
rect 5773 10153 5787 10167
rect 5653 9993 5667 10007
rect 5713 9973 5727 9987
rect 5773 9973 5787 9987
rect 5653 9953 5667 9967
rect 5693 9953 5707 9967
rect 5673 9933 5687 9947
rect 5813 9953 5827 9967
rect 5833 9773 5847 9787
rect 5653 9713 5667 9727
rect 5693 9713 5707 9727
rect 5713 9713 5727 9727
rect 5633 9493 5647 9507
rect 5613 9393 5627 9407
rect 5613 9273 5627 9287
rect 5573 9253 5587 9267
rect 5573 9213 5587 9227
rect 5553 9193 5567 9207
rect 5633 9193 5647 9207
rect 5593 8993 5607 9007
rect 5613 8993 5627 9007
rect 5533 8973 5547 8987
rect 5573 8933 5587 8947
rect 5593 8773 5607 8787
rect 5613 8773 5627 8787
rect 5573 8573 5587 8587
rect 5813 9753 5827 9767
rect 5793 9713 5807 9727
rect 5773 9653 5787 9667
rect 5733 9293 5747 9307
rect 5713 9253 5727 9267
rect 5753 9233 5767 9247
rect 5813 9453 5827 9467
rect 5793 9373 5807 9387
rect 5773 9193 5787 9207
rect 5653 8973 5667 8987
rect 5753 9033 5767 9047
rect 5733 9013 5747 9027
rect 5713 8793 5727 8807
rect 5693 8773 5707 8787
rect 5693 8733 5707 8747
rect 5633 8553 5647 8567
rect 5673 8533 5687 8547
rect 5633 8513 5647 8527
rect 5513 8473 5527 8487
rect 5553 8473 5567 8487
rect 5613 8493 5627 8507
rect 5593 8473 5607 8487
rect 5633 8473 5647 8487
rect 5573 8393 5587 8407
rect 5473 8373 5487 8387
rect 5453 8273 5467 8287
rect 5433 8013 5447 8027
rect 5353 7993 5367 8007
rect 5393 7993 5407 8007
rect 5333 7833 5347 7847
rect 5293 7773 5307 7787
rect 5273 7633 5287 7647
rect 5293 7573 5307 7587
rect 5193 7433 5207 7447
rect 5213 7353 5227 7367
rect 5193 7313 5207 7327
rect 5153 7293 5167 7307
rect 5273 7493 5287 7507
rect 5253 7353 5267 7367
rect 5153 7273 5167 7287
rect 5233 7273 5247 7287
rect 5133 7093 5147 7107
rect 5073 7013 5087 7027
rect 5113 7013 5127 7027
rect 5113 6913 5127 6927
rect 4993 6853 5007 6867
rect 5053 6853 5067 6867
rect 4953 6773 4967 6787
rect 4913 6693 4927 6707
rect 4833 6553 4847 6567
rect 5093 6713 5107 6727
rect 5093 6633 5107 6647
rect 5013 6573 5027 6587
rect 5333 7513 5347 7527
rect 5313 7473 5327 7487
rect 5313 7373 5327 7387
rect 5273 7273 5287 7287
rect 5253 7213 5267 7227
rect 5193 7173 5207 7187
rect 5273 7093 5287 7107
rect 5233 7073 5247 7087
rect 5253 7053 5267 7067
rect 5293 7053 5307 7067
rect 5333 7313 5347 7327
rect 5333 7173 5347 7187
rect 5393 7893 5407 7907
rect 5373 7833 5387 7847
rect 5413 7833 5427 7847
rect 5413 7593 5427 7607
rect 5393 7573 5407 7587
rect 5373 7453 5387 7467
rect 5353 7133 5367 7147
rect 5353 7053 5367 7067
rect 5153 6633 5167 6647
rect 5133 6473 5147 6487
rect 4993 6453 5007 6467
rect 5033 6453 5047 6467
rect 4893 6433 4907 6447
rect 4813 6413 4827 6427
rect 4873 6293 4887 6307
rect 4813 6093 4827 6107
rect 4773 6073 4787 6087
rect 4873 6093 4887 6107
rect 4833 6053 4847 6067
rect 4753 5973 4767 5987
rect 4793 5913 4807 5927
rect 4873 6033 4887 6047
rect 4873 5913 4887 5927
rect 4773 5893 4787 5907
rect 4813 5893 4827 5907
rect 4853 5893 4867 5907
rect 4853 5873 4867 5887
rect 4793 5693 4807 5707
rect 4753 5493 4767 5507
rect 4733 5373 4747 5387
rect 4733 5153 4747 5167
rect 4713 4893 4727 4907
rect 4753 4853 4767 4867
rect 4813 5553 4827 5567
rect 4833 5473 4847 5487
rect 4813 5233 4827 5247
rect 5033 6373 5047 6387
rect 5333 6953 5347 6967
rect 5293 6933 5307 6947
rect 5193 6873 5207 6887
rect 5253 6873 5267 6887
rect 5293 6873 5307 6887
rect 5453 7933 5467 7947
rect 5453 7833 5467 7847
rect 5453 7533 5467 7547
rect 5453 7513 5467 7527
rect 5433 7453 5447 7467
rect 5573 8353 5587 8367
rect 5513 8313 5527 8327
rect 5533 8313 5547 8327
rect 5513 8293 5527 8307
rect 5513 8113 5527 8127
rect 5633 8373 5647 8387
rect 5553 8173 5567 8187
rect 5573 8173 5587 8187
rect 5533 8093 5547 8107
rect 5533 8033 5547 8047
rect 5553 8033 5567 8047
rect 5493 8013 5507 8027
rect 5513 7793 5527 7807
rect 5533 7793 5547 7807
rect 5573 7913 5587 7927
rect 5553 7653 5567 7667
rect 5573 7653 5587 7667
rect 5493 7593 5507 7607
rect 5513 7593 5527 7607
rect 5553 7573 5567 7587
rect 5533 7533 5547 7547
rect 5613 8273 5627 8287
rect 5613 8113 5627 8127
rect 5633 8113 5647 8127
rect 5673 8273 5687 8287
rect 5673 8233 5687 8247
rect 5653 8013 5667 8027
rect 5713 8553 5727 8567
rect 5773 8853 5787 8867
rect 5753 8773 5767 8787
rect 5753 8673 5767 8687
rect 5753 8553 5767 8567
rect 5713 7973 5727 7987
rect 5733 7973 5747 7987
rect 5673 7953 5687 7967
rect 5693 7953 5707 7967
rect 5713 7913 5727 7927
rect 5633 7893 5647 7907
rect 5673 7893 5687 7907
rect 5633 7873 5647 7887
rect 5653 7833 5667 7847
rect 5733 7853 5747 7867
rect 5713 7813 5727 7827
rect 5733 7813 5747 7827
rect 5613 7673 5627 7687
rect 5553 7473 5567 7487
rect 5513 7433 5527 7447
rect 5533 7413 5547 7427
rect 5473 7373 5487 7387
rect 5493 7353 5507 7367
rect 5393 7333 5407 7347
rect 5473 7333 5487 7347
rect 5433 7313 5447 7327
rect 5533 7313 5547 7327
rect 5413 7273 5427 7287
rect 5513 7273 5527 7287
rect 5393 7253 5407 7267
rect 5393 6953 5407 6967
rect 5373 6873 5387 6887
rect 5233 6773 5247 6787
rect 5213 6573 5227 6587
rect 5233 6573 5247 6587
rect 5193 6433 5207 6447
rect 5213 6393 5227 6407
rect 5093 6253 5107 6267
rect 4993 5713 5007 5727
rect 4953 5633 4967 5647
rect 4893 5473 4907 5487
rect 4913 5473 4927 5487
rect 4853 5413 4867 5427
rect 4873 5413 4887 5427
rect 4913 5413 4927 5427
rect 4853 5353 4867 5367
rect 4953 5393 4967 5407
rect 4873 5333 4887 5347
rect 4933 5333 4947 5347
rect 4893 5293 4907 5307
rect 4893 5173 4907 5187
rect 4913 5153 4927 5167
rect 4833 5133 4847 5147
rect 4873 5133 4887 5147
rect 4893 5133 4907 5147
rect 5113 5933 5127 5947
rect 5113 5873 5127 5887
rect 5233 6193 5247 6207
rect 5313 6853 5327 6867
rect 5273 6833 5287 6847
rect 5273 6773 5287 6787
rect 5373 6693 5387 6707
rect 5353 6633 5367 6647
rect 5313 6613 5327 6627
rect 5353 6593 5367 6607
rect 5293 6573 5307 6587
rect 5333 6553 5347 6567
rect 5273 6473 5287 6487
rect 5333 6453 5347 6467
rect 5313 6413 5327 6427
rect 5333 6413 5347 6427
rect 5293 6333 5307 6347
rect 5193 5813 5207 5827
rect 5333 6393 5347 6407
rect 5313 6073 5327 6087
rect 5273 5993 5287 6007
rect 5473 7233 5487 7247
rect 5413 6893 5427 6907
rect 5413 6713 5427 6727
rect 5413 6653 5427 6667
rect 5513 7213 5527 7227
rect 5473 6733 5487 6747
rect 5533 6693 5547 6707
rect 5613 7533 5627 7547
rect 5573 7393 5587 7407
rect 5613 7333 5627 7347
rect 5613 7293 5627 7307
rect 5593 7193 5607 7207
rect 5593 6933 5607 6947
rect 5613 6933 5627 6947
rect 5593 6853 5607 6867
rect 5593 6833 5607 6847
rect 5573 6813 5587 6827
rect 5533 6633 5547 6647
rect 5553 6633 5567 6647
rect 5653 7593 5667 7607
rect 5673 7553 5687 7567
rect 5653 7513 5667 7527
rect 5653 7093 5667 7107
rect 5573 6613 5587 6627
rect 5553 6593 5567 6607
rect 5433 6553 5447 6567
rect 5433 6533 5447 6547
rect 5433 6493 5447 6507
rect 5393 6453 5407 6467
rect 5373 6013 5387 6027
rect 5273 5953 5287 5967
rect 5253 5873 5267 5887
rect 5233 5773 5247 5787
rect 5293 5713 5307 5727
rect 5073 5673 5087 5687
rect 4973 5233 4987 5247
rect 4973 5093 4987 5107
rect 5053 5593 5067 5607
rect 5033 5413 5047 5427
rect 5013 5033 5027 5047
rect 4893 4853 4907 4867
rect 4953 4853 4967 4867
rect 4953 4793 4967 4807
rect 4833 4773 4847 4787
rect 4773 4713 4787 4727
rect 4773 4693 4787 4707
rect 4693 4593 4707 4607
rect 4693 4473 4707 4487
rect 4693 4413 4707 4427
rect 4673 4293 4687 4307
rect 4593 4253 4607 4267
rect 4633 3993 4647 4007
rect 4693 4213 4707 4227
rect 4713 4193 4727 4207
rect 4893 4573 4907 4587
rect 4853 4493 4867 4507
rect 4913 4553 4927 4567
rect 4913 4413 4927 4427
rect 4873 4393 4887 4407
rect 4793 4173 4807 4187
rect 4893 4133 4907 4147
rect 4713 4113 4727 4127
rect 4693 3973 4707 3987
rect 4533 3953 4547 3967
rect 4653 3953 4667 3967
rect 4553 3753 4567 3767
rect 4613 3713 4627 3727
rect 4693 3713 4707 3727
rect 4593 3693 4607 3707
rect 4573 3653 4587 3667
rect 4633 3653 4647 3667
rect 4513 3553 4527 3567
rect 4533 3493 4547 3507
rect 4553 3473 4567 3487
rect 4513 3433 4527 3447
rect 4533 3053 4547 3067
rect 4453 2733 4467 2747
rect 4453 2533 4467 2547
rect 4513 2913 4527 2927
rect 4433 2453 4447 2467
rect 4433 2233 4447 2247
rect 4413 2173 4427 2187
rect 4393 1813 4407 1827
rect 4473 2353 4487 2367
rect 4453 1853 4467 1867
rect 4433 1773 4447 1787
rect 4353 1753 4367 1767
rect 4273 1653 4287 1667
rect 4093 1593 4107 1607
rect 4213 1593 4227 1607
rect 4193 1313 4207 1327
rect 4053 1233 4067 1247
rect 3993 1193 4007 1207
rect 3853 1073 3867 1087
rect 4033 1133 4047 1147
rect 3833 1053 3847 1067
rect 3793 933 3807 947
rect 3773 873 3787 887
rect 3753 853 3767 867
rect 3833 833 3847 847
rect 3773 653 3787 667
rect 3773 633 3787 647
rect 3753 373 3767 387
rect 3793 373 3807 387
rect 3833 793 3847 807
rect 3833 313 3847 327
rect 4053 913 4067 927
rect 4053 813 4067 827
rect 4033 773 4047 787
rect 3973 673 3987 687
rect 4013 673 4027 687
rect 3953 613 3967 627
rect 3993 613 4007 627
rect 3953 393 3967 407
rect 3993 373 4007 387
rect 4073 773 4087 787
rect 4493 2273 4507 2287
rect 4593 3573 4607 3587
rect 4593 3393 4607 3407
rect 4673 3253 4687 3267
rect 4573 2733 4587 2747
rect 4553 2593 4567 2607
rect 4633 3233 4647 3247
rect 4613 3213 4627 3227
rect 4653 3213 4667 3227
rect 4673 3213 4687 3227
rect 4633 3033 4647 3047
rect 4913 4033 4927 4047
rect 4853 3993 4867 4007
rect 4933 3953 4947 3967
rect 4853 3893 4867 3907
rect 4933 3833 4947 3847
rect 4853 3773 4867 3787
rect 4893 3733 4907 3747
rect 4833 3673 4847 3687
rect 4873 3673 4887 3687
rect 4813 3513 4827 3527
rect 4753 3493 4767 3507
rect 4773 3453 4787 3467
rect 4813 3453 4827 3467
rect 4733 3313 4747 3327
rect 4713 3233 4727 3247
rect 4793 3233 4807 3247
rect 4713 3153 4727 3167
rect 4733 3053 4747 3067
rect 4713 3033 4727 3047
rect 4773 3013 4787 3027
rect 4653 2713 4667 2727
rect 4593 2553 4607 2567
rect 4633 2573 4647 2587
rect 4573 2533 4587 2547
rect 4613 2533 4627 2547
rect 4593 2373 4607 2387
rect 4553 2093 4567 2107
rect 4513 1873 4527 1887
rect 4573 1853 4587 1867
rect 4513 1833 4527 1847
rect 4553 1813 4567 1827
rect 4613 2033 4627 2047
rect 4593 1793 4607 1807
rect 4493 1733 4507 1747
rect 4533 1733 4547 1747
rect 4493 1693 4507 1707
rect 4353 1633 4367 1647
rect 4473 1633 4487 1647
rect 4533 1633 4547 1647
rect 4253 1533 4267 1547
rect 4293 1433 4307 1447
rect 4273 1313 4287 1327
rect 4213 1293 4227 1307
rect 4253 1293 4267 1307
rect 4313 1273 4327 1287
rect 4293 1253 4307 1267
rect 4233 1153 4247 1167
rect 4233 1133 4247 1147
rect 4253 1093 4267 1107
rect 4213 833 4227 847
rect 4253 833 4267 847
rect 4293 833 4307 847
rect 4273 813 4287 827
rect 4213 773 4227 787
rect 4193 673 4207 687
rect 4213 653 4227 667
rect 4073 613 4087 627
rect 4273 653 4287 667
rect 4053 353 4067 367
rect 4213 353 4227 367
rect 4473 1613 4487 1627
rect 4513 1613 4527 1627
rect 4373 1593 4387 1607
rect 4493 1593 4507 1607
rect 4473 1553 4487 1567
rect 4433 1533 4447 1547
rect 4413 1233 4427 1247
rect 4393 1113 4407 1127
rect 4513 1433 4527 1447
rect 4513 1313 4527 1327
rect 4553 1313 4567 1327
rect 4593 1313 4607 1327
rect 4693 2733 4707 2747
rect 4733 2553 4747 2567
rect 4773 2553 4787 2567
rect 4713 2313 4727 2327
rect 4673 2273 4687 2287
rect 4673 2073 4687 2087
rect 4653 1753 4667 1767
rect 4853 3233 4867 3247
rect 4873 2853 4887 2867
rect 4813 2733 4827 2747
rect 4813 2633 4827 2647
rect 4813 2573 4827 2587
rect 4833 2573 4847 2587
rect 4853 2553 4867 2567
rect 4773 2533 4787 2547
rect 4793 2533 4807 2547
rect 4833 2393 4847 2407
rect 4793 2213 4807 2227
rect 4753 2073 4767 2087
rect 4733 2053 4747 2067
rect 4813 2053 4827 2067
rect 4933 2773 4947 2787
rect 5013 4753 5027 4767
rect 4973 4653 4987 4667
rect 4973 4453 4987 4467
rect 4973 4013 4987 4027
rect 4993 3953 5007 3967
rect 5193 5653 5207 5667
rect 5073 5393 5087 5407
rect 5053 5353 5067 5367
rect 5193 5613 5207 5627
rect 5213 5593 5227 5607
rect 5193 5513 5207 5527
rect 5153 5473 5167 5487
rect 5373 5453 5387 5467
rect 5133 5413 5147 5427
rect 5173 5413 5187 5427
rect 5213 5413 5227 5427
rect 5093 5273 5107 5287
rect 5173 5273 5187 5287
rect 5353 5193 5367 5207
rect 5213 5173 5227 5187
rect 5233 5173 5247 5187
rect 5113 5153 5127 5167
rect 5153 5153 5167 5167
rect 5213 5153 5227 5167
rect 5053 5033 5067 5047
rect 5133 5033 5147 5047
rect 5213 5073 5227 5087
rect 5193 4933 5207 4947
rect 5333 4993 5347 5007
rect 5053 4693 5067 4707
rect 5213 4653 5227 4667
rect 5053 4633 5067 4647
rect 5033 4613 5047 4627
rect 5033 4593 5047 4607
rect 5013 3713 5027 3727
rect 5013 3653 5027 3667
rect 4973 3513 4987 3527
rect 5093 4613 5107 4627
rect 5073 4493 5087 4507
rect 5273 4633 5287 4647
rect 5293 4613 5307 4627
rect 5253 4593 5267 4607
rect 5233 4493 5247 4507
rect 5473 6433 5487 6447
rect 5513 6413 5527 6427
rect 5533 6373 5547 6387
rect 5493 6353 5507 6367
rect 5593 6353 5607 6367
rect 5553 6293 5567 6307
rect 5493 6193 5507 6207
rect 5473 6113 5487 6127
rect 5453 6073 5467 6087
rect 5453 5933 5467 5947
rect 5533 6173 5547 6187
rect 5433 5373 5447 5387
rect 5413 5173 5427 5187
rect 5353 4473 5367 4487
rect 5253 4453 5267 4467
rect 5353 4453 5367 4467
rect 5093 4413 5107 4427
rect 5173 4333 5187 4347
rect 5073 4293 5087 4307
rect 5093 4213 5107 4227
rect 5053 4033 5067 4047
rect 5073 3973 5087 3987
rect 5053 3753 5067 3767
rect 5053 3733 5067 3747
rect 5033 3633 5047 3647
rect 5033 3493 5047 3507
rect 4993 3453 5007 3467
rect 5133 3713 5147 3727
rect 5113 3653 5127 3667
rect 5213 4293 5227 4307
rect 5173 3993 5187 4007
rect 5433 5133 5447 5147
rect 5413 4853 5427 4867
rect 5413 4733 5427 4747
rect 5473 5653 5487 5667
rect 5513 5773 5527 5787
rect 5513 5333 5527 5347
rect 5453 4573 5467 4587
rect 5453 4533 5467 4547
rect 5433 4293 5447 4307
rect 5313 4213 5327 4227
rect 5373 4213 5387 4227
rect 5253 4013 5267 4027
rect 5273 4013 5287 4027
rect 5193 3973 5207 3987
rect 5193 3953 5207 3967
rect 5233 3933 5247 3947
rect 5253 3873 5267 3887
rect 5173 3693 5187 3707
rect 5173 3633 5187 3647
rect 5153 3593 5167 3607
rect 5093 3513 5107 3527
rect 5073 3373 5087 3387
rect 5173 3493 5187 3507
rect 5133 3473 5147 3487
rect 5033 3113 5047 3127
rect 4973 3073 4987 3087
rect 5113 3013 5127 3027
rect 5173 3033 5187 3047
rect 5053 2893 5067 2907
rect 5133 2893 5147 2907
rect 4953 2713 4967 2727
rect 5113 2793 5127 2807
rect 5113 2753 5127 2767
rect 5173 2853 5187 2867
rect 5213 3533 5227 3547
rect 5373 4173 5387 4187
rect 5333 4153 5347 4167
rect 5333 3993 5347 4007
rect 5493 5053 5507 5067
rect 5593 5733 5607 5747
rect 5573 5713 5587 5727
rect 5573 5653 5587 5667
rect 5553 5453 5567 5467
rect 5633 6113 5647 6127
rect 5613 5653 5627 5667
rect 5593 5593 5607 5607
rect 5533 5013 5547 5027
rect 5513 4993 5527 5007
rect 5533 4933 5547 4947
rect 5613 5293 5627 5307
rect 5613 5173 5627 5187
rect 5613 5073 5627 5087
rect 5593 4993 5607 5007
rect 5513 4913 5527 4927
rect 5573 4913 5587 4927
rect 5553 4693 5567 4707
rect 5533 4673 5547 4687
rect 5533 4653 5547 4667
rect 5493 4633 5507 4647
rect 5513 4573 5527 4587
rect 5513 4373 5527 4387
rect 5273 3533 5287 3547
rect 5313 3533 5327 3547
rect 5193 2793 5207 2807
rect 5233 3493 5247 3507
rect 5273 3473 5287 3487
rect 5313 3453 5327 3467
rect 5293 3273 5307 3287
rect 5273 3233 5287 3247
rect 5233 3173 5247 3187
rect 5313 3033 5327 3047
rect 5233 3013 5247 3027
rect 5233 2853 5247 2867
rect 5153 2753 5167 2767
rect 5193 2753 5207 2767
rect 5133 2733 5147 2747
rect 5053 2573 5067 2587
rect 5113 2573 5127 2587
rect 4913 2393 4927 2407
rect 5073 2533 5087 2547
rect 5193 2633 5207 2647
rect 5173 2533 5187 2547
rect 5013 2373 5027 2387
rect 5213 2453 5227 2467
rect 5193 2293 5207 2307
rect 5033 2213 5047 2227
rect 4853 2173 4867 2187
rect 4933 2173 4947 2187
rect 4913 2053 4927 2067
rect 4833 2033 4847 2047
rect 4873 2033 4887 2047
rect 4773 1833 4787 1847
rect 4753 1813 4767 1827
rect 4713 1673 4727 1687
rect 4673 1653 4687 1667
rect 5213 2173 5227 2187
rect 5153 2153 5167 2167
rect 5193 2153 5207 2167
rect 5193 2133 5207 2147
rect 4773 1733 4787 1747
rect 4673 1593 4687 1607
rect 4713 1593 4727 1607
rect 4753 1593 4767 1607
rect 4473 1113 4487 1127
rect 4473 1013 4487 1027
rect 4493 1013 4507 1027
rect 4413 933 4427 947
rect 4413 813 4427 827
rect 4393 673 4407 687
rect 4453 833 4467 847
rect 4533 1293 4547 1307
rect 4573 1273 4587 1287
rect 4533 1073 4547 1087
rect 4513 833 4527 847
rect 4533 813 4547 827
rect 4493 753 4507 767
rect 4973 1693 4987 1707
rect 5193 2053 5207 2067
rect 5093 1893 5107 1907
rect 5073 1813 5087 1827
rect 5053 1753 5067 1767
rect 5053 1593 5067 1607
rect 5033 1573 5047 1587
rect 4993 1533 5007 1547
rect 5253 2773 5267 2787
rect 5273 2753 5287 2767
rect 5253 2293 5267 2307
rect 5293 2733 5307 2747
rect 5473 3993 5487 4007
rect 5393 3973 5407 3987
rect 5433 3973 5447 3987
rect 5493 3933 5507 3947
rect 5493 3753 5507 3767
rect 5373 3733 5387 3747
rect 5353 3713 5367 3727
rect 5413 3713 5427 3727
rect 5573 4633 5587 4647
rect 5553 4573 5567 4587
rect 5713 7593 5727 7607
rect 5813 8993 5827 9007
rect 6073 10253 6087 10267
rect 6253 10733 6267 10747
rect 6293 10713 6307 10727
rect 6313 10693 6327 10707
rect 6393 10933 6407 10947
rect 6373 10873 6387 10887
rect 6353 10673 6367 10687
rect 6473 10913 6487 10927
rect 6753 10913 6767 10927
rect 6953 10913 6967 10927
rect 6993 10913 7007 10927
rect 6673 10893 6687 10907
rect 6473 10873 6487 10887
rect 6493 10813 6507 10827
rect 6433 10753 6447 10767
rect 6393 10473 6407 10487
rect 6293 10453 6307 10467
rect 6333 10453 6347 10467
rect 5993 10133 6007 10147
rect 6233 10133 6247 10147
rect 5973 10113 5987 10127
rect 5933 9973 5947 9987
rect 5873 9953 5887 9967
rect 5853 9473 5867 9487
rect 5913 9933 5927 9947
rect 5953 9753 5967 9767
rect 5953 9713 5967 9727
rect 5953 9673 5967 9687
rect 5913 9273 5927 9287
rect 5993 9993 6007 10007
rect 6033 9953 6047 9967
rect 6133 9953 6147 9967
rect 6113 9833 6127 9847
rect 6053 9773 6067 9787
rect 5993 9753 6007 9767
rect 6033 9753 6047 9767
rect 6013 9653 6027 9667
rect 6013 9473 6027 9487
rect 6053 9473 6067 9487
rect 6093 9473 6107 9487
rect 5993 9453 6007 9467
rect 5973 9373 5987 9387
rect 6033 9433 6047 9447
rect 5933 9253 5947 9267
rect 5973 9193 5987 9207
rect 5933 9153 5947 9167
rect 5993 9153 6007 9167
rect 5853 9033 5867 9047
rect 5993 9113 6007 9127
rect 5953 9053 5967 9067
rect 5873 9013 5887 9027
rect 5933 9013 5947 9027
rect 5853 8973 5867 8987
rect 5953 8993 5967 9007
rect 5933 8893 5947 8907
rect 5893 8793 5907 8807
rect 5973 8813 5987 8827
rect 6093 9073 6107 9087
rect 6033 9033 6047 9047
rect 5993 8793 6007 8807
rect 5913 8773 5927 8787
rect 5853 8633 5867 8647
rect 5793 8493 5807 8507
rect 5793 8253 5807 8267
rect 5853 8533 5867 8547
rect 5893 8513 5907 8527
rect 5833 8493 5847 8507
rect 5873 8473 5887 8487
rect 5853 8453 5867 8467
rect 5913 8453 5927 8467
rect 5853 8333 5867 8347
rect 5833 8273 5847 8287
rect 5793 8133 5807 8147
rect 5813 8133 5827 8147
rect 5773 8093 5787 8107
rect 5873 8133 5887 8147
rect 5833 8053 5847 8067
rect 5793 8033 5807 8047
rect 5833 8033 5847 8047
rect 5793 8013 5807 8027
rect 5813 8013 5827 8027
rect 5913 8053 5927 8067
rect 5973 8533 5987 8547
rect 6013 8513 6027 8527
rect 5953 8473 5967 8487
rect 5973 8473 5987 8487
rect 5993 8453 6007 8467
rect 5773 7733 5787 7747
rect 5813 7973 5827 7987
rect 5793 7573 5807 7587
rect 5733 7553 5747 7567
rect 5753 7553 5767 7567
rect 5793 7533 5807 7547
rect 5693 7473 5707 7487
rect 5693 7373 5707 7387
rect 5753 7513 5767 7527
rect 5773 7393 5787 7407
rect 5793 7353 5807 7367
rect 5753 7333 5767 7347
rect 5693 7173 5707 7187
rect 5713 7173 5727 7187
rect 5673 7033 5687 7047
rect 5673 6913 5687 6927
rect 5773 7093 5787 7107
rect 5733 7073 5747 7087
rect 5713 7053 5727 7067
rect 5753 7053 5767 7067
rect 5713 7013 5727 7027
rect 5733 6973 5747 6987
rect 5713 6913 5727 6927
rect 5693 6853 5707 6867
rect 5673 6633 5687 6647
rect 5853 7873 5867 7887
rect 5833 7853 5847 7867
rect 5913 8013 5927 8027
rect 5933 8013 5947 8027
rect 5933 7993 5947 8007
rect 5953 7993 5967 8007
rect 5993 7973 6007 7987
rect 5873 7853 5887 7867
rect 5893 7833 5907 7847
rect 5973 7833 5987 7847
rect 5913 7813 5927 7827
rect 5853 7793 5867 7807
rect 5873 7793 5887 7807
rect 5833 7613 5847 7627
rect 5853 7513 5867 7527
rect 5853 7413 5867 7427
rect 5833 7273 5847 7287
rect 5753 6873 5767 6887
rect 5793 6873 5807 6887
rect 5813 6853 5827 6867
rect 5813 6813 5827 6827
rect 5853 7073 5867 7087
rect 5853 6833 5867 6847
rect 5833 6713 5847 6727
rect 5833 6613 5847 6627
rect 5793 6533 5807 6547
rect 5833 6533 5847 6547
rect 5853 6533 5867 6547
rect 5813 6413 5827 6427
rect 5733 6393 5747 6407
rect 5813 6393 5827 6407
rect 5753 6373 5767 6387
rect 5773 6353 5787 6367
rect 5733 6333 5747 6347
rect 5673 6293 5687 6307
rect 5693 6113 5707 6127
rect 5733 6113 5747 6127
rect 5673 6093 5687 6107
rect 5773 6093 5787 6107
rect 5833 6153 5847 6167
rect 5733 5973 5747 5987
rect 5813 5973 5827 5987
rect 5713 5933 5727 5947
rect 5793 5913 5807 5927
rect 5813 5893 5827 5907
rect 5773 5873 5787 5887
rect 5753 5733 5767 5747
rect 5693 5633 5707 5647
rect 5713 5633 5727 5647
rect 5753 5633 5767 5647
rect 5673 5593 5687 5607
rect 5673 5553 5687 5567
rect 5653 5373 5667 5387
rect 5633 4893 5647 4907
rect 5733 5613 5747 5627
rect 5733 5473 5747 5487
rect 5713 5113 5727 5127
rect 5693 4793 5707 4807
rect 5713 4793 5727 4807
rect 5693 4713 5707 4727
rect 5673 4653 5687 4667
rect 5653 4493 5667 4507
rect 5633 4333 5647 4347
rect 5633 4273 5647 4287
rect 5593 4193 5607 4207
rect 5613 4173 5627 4187
rect 5633 4173 5647 4187
rect 5553 3973 5567 3987
rect 5533 3913 5547 3927
rect 5513 3693 5527 3707
rect 5393 3673 5407 3687
rect 5433 3673 5447 3687
rect 5353 3533 5367 3547
rect 5333 2913 5347 2927
rect 5493 3513 5507 3527
rect 5553 3773 5567 3787
rect 5593 4133 5607 4147
rect 5673 4013 5687 4027
rect 5693 3993 5707 4007
rect 5613 3973 5627 3987
rect 5593 3733 5607 3747
rect 5693 3873 5707 3887
rect 5673 3793 5687 3807
rect 5673 3713 5687 3727
rect 5613 3673 5627 3687
rect 5633 3673 5647 3687
rect 5573 3633 5587 3647
rect 5593 3633 5607 3647
rect 5553 3613 5567 3627
rect 5573 3533 5587 3547
rect 5633 3593 5647 3607
rect 5613 3553 5627 3567
rect 5513 3493 5527 3507
rect 5593 3493 5607 3507
rect 5553 3433 5567 3447
rect 5453 3273 5467 3287
rect 5533 3253 5547 3267
rect 5493 3173 5507 3187
rect 5373 3013 5387 3027
rect 5453 3033 5467 3047
rect 5433 3013 5447 3027
rect 5473 3013 5487 3027
rect 5393 2993 5407 3007
rect 5353 2853 5367 2867
rect 5313 2713 5327 2727
rect 5413 2713 5427 2727
rect 5353 2673 5367 2687
rect 5393 2673 5407 2687
rect 5313 2573 5327 2587
rect 5553 2653 5567 2667
rect 5553 2613 5567 2627
rect 5753 5273 5767 5287
rect 5793 5793 5807 5807
rect 5773 5033 5787 5047
rect 5833 5873 5847 5887
rect 5853 5753 5867 5767
rect 5893 7733 5907 7747
rect 5893 7673 5907 7687
rect 5893 7413 5907 7427
rect 5873 5633 5887 5647
rect 5813 5553 5827 5567
rect 5873 5453 5887 5467
rect 5833 5413 5847 5427
rect 5873 5353 5887 5367
rect 5873 5173 5887 5187
rect 5813 5073 5827 5087
rect 5813 5033 5827 5047
rect 5793 4873 5807 4887
rect 5773 4733 5787 4747
rect 5733 4713 5747 4727
rect 5773 4713 5787 4727
rect 5733 4673 5747 4687
rect 5793 4633 5807 4647
rect 5793 4513 5807 4527
rect 5773 4473 5787 4487
rect 5713 3413 5727 3427
rect 5653 3353 5667 3367
rect 5633 2633 5647 2647
rect 5613 2573 5627 2587
rect 5593 2553 5607 2567
rect 5333 2533 5347 2547
rect 5293 2473 5307 2487
rect 5413 2233 5427 2247
rect 5593 2173 5607 2187
rect 5293 2133 5307 2147
rect 5313 2093 5327 2107
rect 5473 2093 5487 2107
rect 5833 4973 5847 4987
rect 5833 4693 5847 4707
rect 5933 7553 5947 7567
rect 6353 10413 6367 10427
rect 6373 10273 6387 10287
rect 6313 9933 6327 9947
rect 6393 9933 6407 9947
rect 6153 9813 6167 9827
rect 6313 9813 6327 9827
rect 6273 9753 6287 9767
rect 6353 9773 6367 9787
rect 6293 9733 6307 9747
rect 6333 9733 6347 9747
rect 6313 9693 6327 9707
rect 6213 9493 6227 9507
rect 6133 9473 6147 9487
rect 6233 9433 6247 9447
rect 6213 9273 6227 9287
rect 6233 9253 6247 9267
rect 6173 9213 6187 9227
rect 6213 9053 6227 9067
rect 6153 8973 6167 8987
rect 6193 8953 6207 8967
rect 6133 8893 6147 8907
rect 6153 8833 6167 8847
rect 6293 9233 6307 9247
rect 6273 9073 6287 9087
rect 6273 8813 6287 8827
rect 6193 8693 6207 8707
rect 6113 8553 6127 8567
rect 6073 8533 6087 8547
rect 6173 8533 6187 8547
rect 6113 8513 6127 8527
rect 6093 8493 6107 8507
rect 6093 8453 6107 8467
rect 6033 8373 6047 8387
rect 6053 8353 6067 8367
rect 6033 8313 6047 8327
rect 6133 8353 6147 8367
rect 6073 8293 6087 8307
rect 6093 8273 6107 8287
rect 6113 8273 6127 8287
rect 6073 8133 6087 8147
rect 6053 8033 6067 8047
rect 6033 8013 6047 8027
rect 6073 7993 6087 8007
rect 6033 7933 6047 7947
rect 5993 7573 6007 7587
rect 5973 7493 5987 7507
rect 5953 7373 5967 7387
rect 6013 7533 6027 7547
rect 6073 7773 6087 7787
rect 6133 8133 6147 8147
rect 6213 8533 6227 8547
rect 6193 8513 6207 8527
rect 6193 8293 6207 8307
rect 6173 8273 6187 8287
rect 6173 8133 6187 8147
rect 6153 8093 6167 8107
rect 6213 8093 6227 8107
rect 6113 7853 6127 7867
rect 6133 7853 6147 7867
rect 6213 7993 6227 8007
rect 6173 7813 6187 7827
rect 6113 7793 6127 7807
rect 6133 7793 6147 7807
rect 6093 7753 6107 7767
rect 6073 7613 6087 7627
rect 6033 7393 6047 7407
rect 5953 7213 5967 7227
rect 5933 7193 5947 7207
rect 5933 7173 5947 7187
rect 5913 6513 5927 6527
rect 6073 7313 6087 7327
rect 6053 7233 6067 7247
rect 6013 7193 6027 7207
rect 5993 7113 6007 7127
rect 6033 7073 6047 7087
rect 6073 7073 6087 7087
rect 5953 7053 5967 7067
rect 6013 7053 6027 7067
rect 5973 7033 5987 7047
rect 5933 6493 5947 6507
rect 6073 6953 6087 6967
rect 5993 6873 6007 6887
rect 6033 6873 6047 6887
rect 6013 6853 6027 6867
rect 6053 6833 6067 6847
rect 6033 6793 6047 6807
rect 6013 6773 6027 6787
rect 5973 6753 5987 6767
rect 6073 6773 6087 6787
rect 6033 6633 6047 6647
rect 5993 6613 6007 6627
rect 6033 6613 6047 6627
rect 6013 6593 6027 6607
rect 5973 6473 5987 6487
rect 6013 6473 6027 6487
rect 5953 6433 5967 6447
rect 5973 6413 5987 6427
rect 5953 6353 5967 6367
rect 6053 6413 6067 6427
rect 6053 6353 6067 6367
rect 5953 6293 5967 6307
rect 6013 6233 6027 6247
rect 5993 6113 6007 6127
rect 5933 6093 5947 6107
rect 5973 6033 5987 6047
rect 6033 6133 6047 6147
rect 6033 6093 6047 6107
rect 6053 6053 6067 6067
rect 5973 5893 5987 5907
rect 5993 5893 6007 5907
rect 5973 5753 5987 5767
rect 5933 5673 5947 5687
rect 5953 5653 5967 5667
rect 5913 5633 5927 5647
rect 5933 5633 5947 5647
rect 6013 5853 6027 5867
rect 6053 5853 6067 5867
rect 6033 5773 6047 5787
rect 6033 5693 6047 5707
rect 6013 5673 6027 5687
rect 5933 5573 5947 5587
rect 5973 5353 5987 5367
rect 5913 5293 5927 5307
rect 6113 7633 6127 7647
rect 6153 7633 6167 7647
rect 6153 7533 6167 7547
rect 6213 7513 6227 7527
rect 6193 7433 6207 7447
rect 6333 9253 6347 9267
rect 6413 9493 6427 9507
rect 6413 9453 6427 9467
rect 6493 10733 6507 10747
rect 6573 10713 6587 10727
rect 6513 10693 6527 10707
rect 6573 10593 6587 10607
rect 6453 10453 6467 10467
rect 6533 10433 6547 10447
rect 6553 10393 6567 10407
rect 6513 10273 6527 10287
rect 6473 10253 6487 10267
rect 6493 10213 6507 10227
rect 6453 10153 6467 10167
rect 6533 9933 6547 9947
rect 6973 10873 6987 10887
rect 6713 10733 6727 10747
rect 6793 10733 6807 10747
rect 6733 10473 6747 10487
rect 6973 10713 6987 10727
rect 6953 10693 6967 10707
rect 7173 11293 7187 11307
rect 7273 11213 7287 11227
rect 8153 11293 8167 11307
rect 8193 11293 8207 11307
rect 7673 11213 7687 11227
rect 8153 11213 8167 11227
rect 7433 11193 7447 11207
rect 8113 11193 8127 11207
rect 7213 11173 7227 11187
rect 7253 11173 7267 11187
rect 7273 11173 7287 11187
rect 7433 11173 7447 11187
rect 7133 11153 7147 11167
rect 7193 11153 7207 11167
rect 7233 11153 7247 11167
rect 7233 11133 7247 11147
rect 7413 11153 7427 11167
rect 7453 11153 7467 11167
rect 7213 10913 7227 10927
rect 7253 10913 7267 10927
rect 7433 10913 7447 10927
rect 7473 10913 7487 10927
rect 7153 10873 7167 10887
rect 7393 10893 7407 10907
rect 7413 10893 7427 10907
rect 7173 10853 7187 10867
rect 7213 10753 7227 10767
rect 7213 10733 7227 10747
rect 7413 10873 7427 10887
rect 7493 10893 7507 10907
rect 7453 10733 7467 10747
rect 7493 10733 7507 10747
rect 7013 10693 7027 10707
rect 7033 10693 7047 10707
rect 7093 10693 7107 10707
rect 7393 10693 7407 10707
rect 6813 10433 6827 10447
rect 6673 10413 6687 10427
rect 6733 10253 6747 10267
rect 6773 10233 6787 10247
rect 6673 10193 6687 10207
rect 6673 9993 6687 10007
rect 6593 9973 6607 9987
rect 6593 9953 6607 9967
rect 6633 9953 6647 9967
rect 6673 9953 6687 9967
rect 6653 9933 6667 9947
rect 6613 9913 6627 9927
rect 6573 9793 6587 9807
rect 6553 9733 6567 9747
rect 6453 9673 6467 9687
rect 6453 9653 6467 9667
rect 6493 9493 6507 9507
rect 6573 9493 6587 9507
rect 6453 9413 6467 9427
rect 6513 9393 6527 9407
rect 6473 9373 6487 9387
rect 6513 9373 6527 9387
rect 6433 9353 6447 9367
rect 6453 9353 6467 9367
rect 6493 9273 6507 9287
rect 6393 9233 6407 9247
rect 6473 9173 6487 9187
rect 6433 9153 6447 9167
rect 6413 9113 6427 9127
rect 6393 9033 6407 9047
rect 6533 9133 6547 9147
rect 6513 9073 6527 9087
rect 6373 8973 6387 8987
rect 6393 8973 6407 8987
rect 6433 8973 6447 8987
rect 6513 8973 6527 8987
rect 6333 8913 6347 8927
rect 6313 8713 6327 8727
rect 6313 8673 6327 8687
rect 6293 8553 6307 8567
rect 6513 8893 6527 8907
rect 6453 8833 6467 8847
rect 6433 8813 6447 8827
rect 6413 8733 6427 8747
rect 6433 8693 6447 8707
rect 6393 8513 6407 8527
rect 6293 8493 6307 8507
rect 6313 8493 6327 8507
rect 6373 8493 6387 8507
rect 6413 8493 6427 8507
rect 6353 8373 6367 8387
rect 6293 8353 6307 8367
rect 6313 8313 6327 8327
rect 6393 8313 6407 8327
rect 6333 8293 6347 8307
rect 6373 8273 6387 8287
rect 6313 8033 6327 8047
rect 6253 7873 6267 7887
rect 6253 7853 6267 7867
rect 6353 8013 6367 8027
rect 6333 7813 6347 7827
rect 6293 7793 6307 7807
rect 6293 7753 6307 7767
rect 6293 7693 6307 7707
rect 6253 7673 6267 7687
rect 6253 7553 6267 7567
rect 6273 7513 6287 7527
rect 6293 7493 6307 7507
rect 6233 7393 6247 7407
rect 6273 7393 6287 7407
rect 6233 7373 6247 7387
rect 6213 7253 6227 7267
rect 6273 7213 6287 7227
rect 6293 7213 6307 7227
rect 6213 7113 6227 7127
rect 6113 7093 6127 7107
rect 6153 7033 6167 7047
rect 6133 6933 6147 6947
rect 6113 6853 6127 6867
rect 6113 6793 6127 6807
rect 6113 6713 6127 6727
rect 6133 6413 6147 6427
rect 6173 6753 6187 6767
rect 6173 6693 6187 6707
rect 6153 6393 6167 6407
rect 6153 6293 6167 6307
rect 6113 6173 6127 6187
rect 6493 8813 6507 8827
rect 6453 8493 6467 8507
rect 6453 8473 6467 8487
rect 6433 8453 6447 8467
rect 6493 8753 6507 8767
rect 6493 8473 6507 8487
rect 6753 10213 6767 10227
rect 6753 10113 6767 10127
rect 6713 9933 6727 9947
rect 6673 9813 6687 9827
rect 6653 9753 6667 9767
rect 6653 9453 6667 9467
rect 6613 9433 6627 9447
rect 6753 9753 6767 9767
rect 6793 9753 6807 9767
rect 6833 10393 6847 10407
rect 6893 10413 6907 10427
rect 6893 10253 6907 10267
rect 6873 10153 6887 10167
rect 7053 10673 7067 10687
rect 7693 10913 7707 10927
rect 7673 10733 7687 10747
rect 8173 11173 8187 11187
rect 8213 11173 8227 11187
rect 8153 11153 8167 11167
rect 8193 11153 8207 11167
rect 8133 11113 8147 11127
rect 7933 11093 7947 11107
rect 8113 10933 8127 10947
rect 8193 10953 8207 10967
rect 8193 10933 8207 10947
rect 8953 11213 8967 11227
rect 9173 11213 9187 11227
rect 8373 11193 8387 11207
rect 8413 11193 8427 11207
rect 8433 11173 8447 11187
rect 8453 11153 8467 11167
rect 8373 10953 8387 10967
rect 8233 10933 8247 10947
rect 8333 10933 8347 10947
rect 8413 10933 8427 10947
rect 7833 10713 7847 10727
rect 7673 10693 7687 10707
rect 7053 10473 7067 10487
rect 7513 10473 7527 10487
rect 7873 10693 7887 10707
rect 7833 10473 7847 10487
rect 7813 10453 7827 10467
rect 7413 10433 7427 10447
rect 7793 10433 7807 10447
rect 7073 10413 7087 10427
rect 7193 10413 7207 10427
rect 7113 10393 7127 10407
rect 7093 10293 7107 10307
rect 6993 10253 7007 10267
rect 6953 10233 6967 10247
rect 7013 10233 7027 10247
rect 6933 10033 6947 10047
rect 6853 9973 6867 9987
rect 6893 9953 6907 9967
rect 6913 9933 6927 9947
rect 6873 9913 6887 9927
rect 6913 9773 6927 9787
rect 6713 9513 6727 9527
rect 6773 9513 6787 9527
rect 6753 9473 6767 9487
rect 6693 9453 6707 9467
rect 6733 9453 6747 9467
rect 6633 9413 6647 9427
rect 6673 9413 6687 9427
rect 6613 9033 6627 9047
rect 6613 8973 6627 8987
rect 6733 9393 6747 9407
rect 6673 9373 6687 9387
rect 6913 9453 6927 9467
rect 6833 9373 6847 9387
rect 6733 9293 6747 9307
rect 6713 9273 6727 9287
rect 6813 9233 6827 9247
rect 6753 9213 6767 9227
rect 6673 9033 6687 9047
rect 6913 9253 6927 9267
rect 6833 9173 6847 9187
rect 6813 8973 6827 8987
rect 6813 8953 6827 8967
rect 6653 8893 6667 8907
rect 6813 8853 6827 8867
rect 6593 8833 6607 8847
rect 6733 8833 6747 8847
rect 6593 8813 6607 8827
rect 6913 9113 6927 9127
rect 6853 8973 6867 8987
rect 7073 10213 7087 10227
rect 6993 9953 7007 9967
rect 6953 9933 6967 9947
rect 6953 9473 6967 9487
rect 7313 10373 7327 10387
rect 7253 10273 7267 10287
rect 7233 10233 7247 10247
rect 7293 10233 7307 10247
rect 7253 10213 7267 10227
rect 7113 10153 7127 10167
rect 7213 10153 7227 10167
rect 7273 9993 7287 10007
rect 7053 9793 7067 9807
rect 7013 9773 7027 9787
rect 7073 9733 7087 9747
rect 7113 9733 7127 9747
rect 7493 10413 7507 10427
rect 7673 10333 7687 10347
rect 7713 10333 7727 10347
rect 7453 10253 7467 10267
rect 7693 10253 7707 10267
rect 7353 10213 7367 10227
rect 7413 10213 7427 10227
rect 7333 9973 7347 9987
rect 7373 9953 7387 9967
rect 7433 9973 7447 9987
rect 7673 10213 7687 10227
rect 7573 9973 7587 9987
rect 7473 9953 7487 9967
rect 7293 9733 7307 9747
rect 7033 9713 7047 9727
rect 7133 9713 7147 9727
rect 7133 9593 7147 9607
rect 7053 9493 7067 9507
rect 7033 9473 7047 9487
rect 6993 9333 7007 9347
rect 7033 9333 7047 9347
rect 6993 9293 7007 9307
rect 6953 9253 6967 9267
rect 6973 9233 6987 9247
rect 7013 9233 7027 9247
rect 7013 9073 7027 9087
rect 6973 9033 6987 9047
rect 6873 8933 6887 8947
rect 6933 8973 6947 8987
rect 6893 8893 6907 8907
rect 6833 8813 6847 8827
rect 6553 8773 6567 8787
rect 6933 8793 6947 8807
rect 6753 8753 6767 8767
rect 6593 8733 6607 8747
rect 6573 8513 6587 8527
rect 6553 8493 6567 8507
rect 6553 8393 6567 8407
rect 6553 8333 6567 8347
rect 6513 8313 6527 8327
rect 6533 8313 6547 8327
rect 6413 7933 6427 7947
rect 6373 7893 6387 7907
rect 6433 7873 6447 7887
rect 6413 7813 6427 7827
rect 6453 7813 6467 7827
rect 6433 7733 6447 7747
rect 6373 7573 6387 7587
rect 6353 7473 6367 7487
rect 6413 7453 6427 7467
rect 6353 7433 6367 7447
rect 6333 7373 6347 7387
rect 6333 7333 6347 7347
rect 6313 7173 6327 7187
rect 6233 7053 6247 7067
rect 6293 7053 6307 7067
rect 6373 6953 6387 6967
rect 6493 7853 6507 7867
rect 6493 7813 6507 7827
rect 6553 8233 6567 8247
rect 6653 8513 6667 8527
rect 6713 8513 6727 8527
rect 6673 8493 6687 8507
rect 6633 8453 6647 8467
rect 6593 8393 6607 8407
rect 6633 8333 6647 8347
rect 6673 8333 6687 8347
rect 6653 8293 6667 8307
rect 6613 8253 6627 8267
rect 6733 8433 6747 8447
rect 6713 8313 6727 8327
rect 6893 8753 6907 8767
rect 6793 8493 6807 8507
rect 6813 8493 6827 8507
rect 6793 8433 6807 8447
rect 6753 8333 6767 8347
rect 6733 8273 6747 8287
rect 6713 8253 6727 8267
rect 6573 8213 6587 8227
rect 6673 8213 6687 8227
rect 6533 8193 6547 8207
rect 6573 8173 6587 8187
rect 6593 8053 6607 8067
rect 6613 8013 6627 8027
rect 6593 7993 6607 8007
rect 6573 7873 6587 7887
rect 6533 7773 6547 7787
rect 6513 7733 6527 7747
rect 6473 7573 6487 7587
rect 6573 7713 6587 7727
rect 6493 7553 6507 7567
rect 6513 7513 6527 7527
rect 6493 7393 6507 7407
rect 6433 7373 6447 7387
rect 6453 7353 6467 7367
rect 6553 7553 6567 7567
rect 6553 7453 6567 7467
rect 6553 7393 6567 7407
rect 6573 7393 6587 7407
rect 6513 7333 6527 7347
rect 6473 7233 6487 7247
rect 6453 7073 6467 7087
rect 6453 7033 6467 7047
rect 6553 7293 6567 7307
rect 6533 7213 6547 7227
rect 6513 7173 6527 7187
rect 6493 7113 6507 7127
rect 6573 7113 6587 7127
rect 6493 6993 6507 7007
rect 6513 6993 6527 7007
rect 6473 6973 6487 6987
rect 6493 6973 6507 6987
rect 6413 6933 6427 6947
rect 6393 6853 6407 6867
rect 6493 6853 6507 6867
rect 6313 6753 6327 6767
rect 6213 6653 6227 6667
rect 6193 6613 6207 6627
rect 6233 6513 6247 6527
rect 6193 6393 6207 6407
rect 6273 6493 6287 6507
rect 6253 6353 6267 6367
rect 6493 6813 6507 6827
rect 6333 6713 6347 6727
rect 6313 6233 6327 6247
rect 6173 6153 6187 6167
rect 6273 6153 6287 6167
rect 6213 6133 6227 6147
rect 6193 6113 6207 6127
rect 6173 6093 6187 6107
rect 6113 6073 6127 6087
rect 6093 5973 6107 5987
rect 6353 6633 6367 6647
rect 6413 6593 6427 6607
rect 6453 6593 6467 6607
rect 6553 6893 6567 6907
rect 6513 6713 6527 6727
rect 6473 6573 6487 6587
rect 6433 6553 6447 6567
rect 6513 6493 6527 6507
rect 6413 6413 6427 6427
rect 6353 6393 6367 6407
rect 6453 6393 6467 6407
rect 6513 6373 6527 6387
rect 6553 6513 6567 6527
rect 6533 6293 6547 6307
rect 6473 6253 6487 6267
rect 6373 6233 6387 6247
rect 6613 7913 6627 7927
rect 6653 7893 6667 7907
rect 6713 8093 6727 8107
rect 6673 7853 6687 7867
rect 6733 8033 6747 8047
rect 6613 7793 6627 7807
rect 6673 7813 6687 7827
rect 6593 6393 6607 6407
rect 6633 7573 6647 7587
rect 6753 7913 6767 7927
rect 6733 7693 6747 7707
rect 6713 7593 6727 7607
rect 6793 8413 6807 8427
rect 6893 8513 6907 8527
rect 6873 8473 6887 8487
rect 6913 8473 6927 8487
rect 6913 8433 6927 8447
rect 6873 8413 6887 8427
rect 6913 8353 6927 8367
rect 6933 8353 6947 8367
rect 6813 8333 6827 8347
rect 6833 8333 6847 8347
rect 6853 8333 6867 8347
rect 6873 8333 6887 8347
rect 6813 8293 6827 8307
rect 6853 8273 6867 8287
rect 6793 8053 6807 8067
rect 6853 8033 6867 8047
rect 6813 8013 6827 8027
rect 6833 7993 6847 8007
rect 6813 7873 6827 7887
rect 6833 7853 6847 7867
rect 6813 7793 6827 7807
rect 6773 7633 6787 7647
rect 6793 7633 6807 7647
rect 6753 7613 6767 7627
rect 6753 7593 6767 7607
rect 6773 7593 6787 7607
rect 6733 7553 6747 7567
rect 6673 7533 6687 7547
rect 6653 7493 6667 7507
rect 6733 7513 6747 7527
rect 6693 7473 6707 7487
rect 6733 7473 6747 7487
rect 6793 7533 6807 7547
rect 6853 7833 6867 7847
rect 6833 7613 6847 7627
rect 6813 7513 6827 7527
rect 6773 7393 6787 7407
rect 6693 7353 6707 7367
rect 6733 7353 6747 7367
rect 6673 7273 6687 7287
rect 6713 7313 6727 7327
rect 6753 7313 6767 7327
rect 6773 7293 6787 7307
rect 6773 7233 6787 7247
rect 6833 7493 6847 7507
rect 6833 7373 6847 7387
rect 6793 7133 6807 7147
rect 6813 7133 6827 7147
rect 6713 7093 6727 7107
rect 6793 7093 6807 7107
rect 6693 7053 6707 7067
rect 6673 6593 6687 6607
rect 6753 7073 6767 7087
rect 6813 6893 6827 6907
rect 6753 6853 6767 6867
rect 6733 6833 6747 6847
rect 6773 6793 6787 6807
rect 6713 6613 6727 6627
rect 6793 6593 6807 6607
rect 6673 6533 6687 6547
rect 6693 6533 6707 6547
rect 7013 8953 7027 8967
rect 7013 8913 7027 8927
rect 6993 8513 7007 8527
rect 7033 8793 7047 8807
rect 7033 8773 7047 8787
rect 7013 8493 7027 8507
rect 6993 8473 7007 8487
rect 7013 8473 7027 8487
rect 7013 8293 7027 8307
rect 7013 8233 7027 8247
rect 6973 7913 6987 7927
rect 6913 7833 6927 7847
rect 6933 7813 6947 7827
rect 6913 7793 6927 7807
rect 6873 7753 6887 7767
rect 7013 7793 7027 7807
rect 6993 7673 7007 7687
rect 7113 9453 7127 9467
rect 7313 9573 7327 9587
rect 7353 9573 7367 9587
rect 7193 9293 7207 9307
rect 7213 9293 7227 9307
rect 7373 9293 7387 9307
rect 7433 9933 7447 9947
rect 7413 9893 7427 9907
rect 7613 9953 7627 9967
rect 7653 9953 7667 9967
rect 7753 10253 7767 10267
rect 7733 10113 7747 10127
rect 7593 9933 7607 9947
rect 7713 9933 7727 9947
rect 7573 9813 7587 9827
rect 7533 9753 7547 9767
rect 7633 9753 7647 9767
rect 7513 9733 7527 9747
rect 7513 9673 7527 9687
rect 7453 9493 7467 9507
rect 7773 9953 7787 9967
rect 7873 10433 7887 10447
rect 7933 10893 7947 10907
rect 8113 10893 8127 10907
rect 8213 10913 8227 10927
rect 8133 10733 8147 10747
rect 7953 10713 7967 10727
rect 8033 10433 8047 10447
rect 7893 10373 7907 10387
rect 7873 10273 7887 10287
rect 7973 10273 7987 10287
rect 7953 10253 7967 10267
rect 7913 10233 7927 10247
rect 7893 10213 7907 10227
rect 7913 10193 7927 10207
rect 7853 10113 7867 10127
rect 7833 9973 7847 9987
rect 7873 9953 7887 9967
rect 7793 9913 7807 9927
rect 7853 9933 7867 9947
rect 7933 10173 7947 10187
rect 7833 9913 7847 9927
rect 7873 9913 7887 9927
rect 7773 9873 7787 9887
rect 7753 9753 7767 9767
rect 7813 9893 7827 9907
rect 7733 9673 7747 9687
rect 7553 9593 7567 9607
rect 7513 9493 7527 9507
rect 7413 9473 7427 9487
rect 7493 9473 7507 9487
rect 7553 9473 7567 9487
rect 7573 9453 7587 9467
rect 7553 9353 7567 9367
rect 7173 9273 7187 9287
rect 7133 9213 7147 9227
rect 7153 9033 7167 9047
rect 7113 8993 7127 9007
rect 7133 8993 7147 9007
rect 7093 8973 7107 8987
rect 7073 8953 7087 8967
rect 7053 8753 7067 8767
rect 7093 8813 7107 8827
rect 7113 8813 7127 8827
rect 7033 7733 7047 7747
rect 7373 9253 7387 9267
rect 7453 9273 7467 9287
rect 7493 9273 7507 9287
rect 7393 9213 7407 9227
rect 7473 9253 7487 9267
rect 7433 9173 7447 9187
rect 7253 9073 7267 9087
rect 7353 8993 7367 9007
rect 7393 8993 7407 9007
rect 7253 8973 7267 8987
rect 7193 8853 7207 8867
rect 7173 8833 7187 8847
rect 7213 8813 7227 8827
rect 7193 8793 7207 8807
rect 7133 8733 7147 8747
rect 7173 8533 7187 8547
rect 7093 8493 7107 8507
rect 7193 8493 7207 8507
rect 7113 8473 7127 8487
rect 7153 8473 7167 8487
rect 7093 8413 7107 8427
rect 7073 8393 7087 8407
rect 7113 8393 7127 8407
rect 7093 8353 7107 8367
rect 7093 8293 7107 8307
rect 7133 8193 7147 8207
rect 7113 8173 7127 8187
rect 7073 8093 7087 8107
rect 7173 8053 7187 8067
rect 7073 8033 7087 8047
rect 7113 8033 7127 8047
rect 7133 8013 7147 8027
rect 7093 7833 7107 7847
rect 7013 7653 7027 7667
rect 7053 7653 7067 7667
rect 6933 7613 6947 7627
rect 7093 7613 7107 7627
rect 6913 7473 6927 7487
rect 6873 7393 6887 7407
rect 6893 7353 6907 7367
rect 6873 7333 6887 7347
rect 6913 7333 6927 7347
rect 6913 7093 6927 7107
rect 6913 6993 6927 7007
rect 6893 6753 6907 6767
rect 6953 7513 6967 7527
rect 7053 7453 7067 7467
rect 7073 7453 7087 7467
rect 6953 7413 6967 7427
rect 7053 7413 7067 7427
rect 6993 7353 7007 7367
rect 6973 7333 6987 7347
rect 7013 7333 7027 7347
rect 6993 7313 7007 7327
rect 6993 7273 7007 7287
rect 6973 7233 6987 7247
rect 6953 7113 6967 7127
rect 6953 7053 6967 7067
rect 7013 7093 7027 7107
rect 6993 7053 7007 7067
rect 7033 7053 7047 7067
rect 6973 7033 6987 7047
rect 7053 7033 7067 7047
rect 6993 6953 7007 6967
rect 7033 6873 7047 6887
rect 6973 6853 6987 6867
rect 6953 6833 6967 6847
rect 7013 6833 7027 6847
rect 6953 6813 6967 6827
rect 6933 6713 6947 6727
rect 6853 6653 6867 6667
rect 6773 6553 6787 6567
rect 6813 6553 6827 6567
rect 6973 6793 6987 6807
rect 6973 6593 6987 6607
rect 6793 6533 6807 6547
rect 6733 6513 6747 6527
rect 6773 6453 6787 6467
rect 6633 6353 6647 6367
rect 6773 6353 6787 6367
rect 6693 6293 6707 6307
rect 6573 6233 6587 6247
rect 6553 6213 6567 6227
rect 6553 6153 6567 6167
rect 6553 6133 6567 6147
rect 6353 6093 6367 6107
rect 6373 6093 6387 6107
rect 6533 6033 6547 6047
rect 6333 5993 6347 6007
rect 6373 5993 6387 6007
rect 6353 5933 6367 5947
rect 6173 5893 6187 5907
rect 6353 5893 6367 5907
rect 6353 5713 6367 5727
rect 6233 5653 6247 5667
rect 6093 5573 6107 5587
rect 6073 5493 6087 5507
rect 6053 5433 6067 5447
rect 6113 5513 6127 5527
rect 6173 5593 6187 5607
rect 6193 5573 6207 5587
rect 6133 5473 6147 5487
rect 6033 5413 6047 5427
rect 6053 5393 6067 5407
rect 6013 5273 6027 5287
rect 5973 5173 5987 5187
rect 6013 5153 6027 5167
rect 5993 5133 6007 5147
rect 5953 5093 5967 5107
rect 5973 5053 5987 5067
rect 6153 5413 6167 5427
rect 6153 5353 6167 5367
rect 6093 5173 6107 5187
rect 6073 5153 6087 5167
rect 6053 5133 6067 5147
rect 6093 5133 6107 5147
rect 6053 5113 6067 5127
rect 5893 4933 5907 4947
rect 5933 4933 5947 4947
rect 5893 4913 5907 4927
rect 5873 4673 5887 4687
rect 5853 4533 5867 4547
rect 5913 4673 5927 4687
rect 5893 4493 5907 4507
rect 5913 4473 5927 4487
rect 5813 4253 5827 4267
rect 5873 4253 5887 4267
rect 5793 4233 5807 4247
rect 5773 3573 5787 3587
rect 5833 4193 5847 4207
rect 5853 4153 5867 4167
rect 5813 4053 5827 4067
rect 5813 3633 5827 3647
rect 5813 3613 5827 3627
rect 5793 3553 5807 3567
rect 5793 3533 5807 3547
rect 5733 3273 5747 3287
rect 5753 3273 5767 3287
rect 5813 3273 5827 3287
rect 5773 3253 5787 3267
rect 5713 3233 5727 3247
rect 5693 3013 5707 3027
rect 5673 2993 5687 3007
rect 5713 2993 5727 3007
rect 5793 3193 5807 3207
rect 5753 2773 5767 2787
rect 5673 2753 5687 2767
rect 5713 2753 5727 2767
rect 5773 2693 5787 2707
rect 5753 2573 5767 2587
rect 5713 2553 5727 2567
rect 5693 2473 5707 2487
rect 5673 2273 5687 2287
rect 5713 2293 5727 2307
rect 5493 2053 5507 2067
rect 5313 2033 5327 2047
rect 5273 1853 5287 1867
rect 5233 1833 5247 1847
rect 5493 1893 5507 1907
rect 5333 1833 5347 1847
rect 5313 1813 5327 1827
rect 5253 1793 5267 1807
rect 5193 1773 5207 1787
rect 5233 1753 5247 1767
rect 5273 1693 5287 1707
rect 5233 1653 5247 1667
rect 5213 1613 5227 1627
rect 5093 1593 5107 1607
rect 5293 1613 5307 1627
rect 5213 1573 5227 1587
rect 5253 1533 5267 1547
rect 4693 1313 4707 1327
rect 4733 1313 4747 1327
rect 4933 1313 4947 1327
rect 5033 1313 5047 1327
rect 4913 1253 4927 1267
rect 4693 1233 4707 1247
rect 4933 1173 4947 1187
rect 4733 1153 4747 1167
rect 4893 1153 4907 1167
rect 4713 1133 4727 1147
rect 4693 1113 4707 1127
rect 4873 1133 4887 1147
rect 4813 1113 4827 1127
rect 4733 853 4747 867
rect 4713 813 4727 827
rect 4753 833 4767 847
rect 4673 753 4687 767
rect 4673 633 4687 647
rect 4533 593 4547 607
rect 4713 613 4727 627
rect 4733 593 4747 607
rect 4373 393 4387 407
rect 4413 393 4427 407
rect 4493 393 4507 407
rect 4353 373 4367 387
rect 4353 353 4367 367
rect 3973 333 3987 347
rect 4033 333 4047 347
rect 4193 333 4207 347
rect 4233 333 4247 347
rect 4733 433 4747 447
rect 4693 413 4707 427
rect 4793 773 4807 787
rect 4753 413 4767 427
rect 4453 353 4467 367
rect 4493 353 4507 367
rect 4533 353 4547 367
rect 3973 293 3987 307
rect 3893 233 3907 247
rect 4473 233 4487 247
rect 3853 213 3867 227
rect 3733 193 3747 207
rect 3873 173 3887 187
rect 4133 213 4147 227
rect 4713 213 4727 227
rect 4033 173 4047 187
rect 4073 153 4087 167
rect 4913 1133 4927 1147
rect 5053 1133 5067 1147
rect 4913 893 4927 907
rect 4873 833 4887 847
rect 4953 873 4967 887
rect 4993 853 5007 867
rect 5033 853 5047 867
rect 5013 813 5027 827
rect 5053 813 5067 827
rect 4953 633 4967 647
rect 4933 613 4947 627
rect 4973 593 4987 607
rect 5013 593 5027 607
rect 4873 433 4887 447
rect 5213 1333 5227 1347
rect 5353 1773 5367 1787
rect 5473 1693 5487 1707
rect 5453 1633 5467 1647
rect 5453 1573 5467 1587
rect 5533 1593 5547 1607
rect 5573 1593 5587 1607
rect 5653 2013 5667 2027
rect 5733 1793 5747 1807
rect 5793 2553 5807 2567
rect 6053 4933 6067 4947
rect 5993 4913 6007 4927
rect 5953 4813 5967 4827
rect 6213 5453 6227 5467
rect 6213 5053 6227 5067
rect 6293 5553 6307 5567
rect 6333 5533 6347 5547
rect 6453 5973 6467 5987
rect 6533 5913 6547 5927
rect 6473 5753 6487 5767
rect 6513 5753 6527 5767
rect 6493 5733 6507 5747
rect 6413 5533 6427 5547
rect 6393 5513 6407 5527
rect 6333 5393 6347 5407
rect 6313 5353 6327 5367
rect 6253 5273 6267 5287
rect 6253 5173 6267 5187
rect 6273 5133 6287 5147
rect 6293 5133 6307 5147
rect 6213 4953 6227 4967
rect 6253 4953 6267 4967
rect 6233 4933 6247 4947
rect 6273 4933 6287 4947
rect 6193 4713 6207 4727
rect 6093 4633 6107 4647
rect 6153 4593 6167 4607
rect 5953 4553 5967 4567
rect 6013 4553 6027 4567
rect 5933 4453 5947 4467
rect 5973 4373 5987 4387
rect 5933 4193 5947 4207
rect 5953 4193 5967 4207
rect 5913 3993 5927 4007
rect 5993 3973 6007 3987
rect 5953 3913 5967 3927
rect 5933 3753 5947 3767
rect 5893 3733 5907 3747
rect 5973 3733 5987 3747
rect 5933 3713 5947 3727
rect 5913 3613 5927 3627
rect 5953 3613 5967 3627
rect 5913 3493 5927 3507
rect 5873 3473 5887 3487
rect 5853 2993 5867 3007
rect 5933 2993 5947 3007
rect 5953 2933 5967 2947
rect 5893 2693 5907 2707
rect 5873 2633 5887 2647
rect 5833 2573 5847 2587
rect 5833 2493 5847 2507
rect 5813 2273 5827 2287
rect 5773 2053 5787 2067
rect 5913 2593 5927 2607
rect 5913 2513 5927 2527
rect 5953 2513 5967 2527
rect 5913 2293 5927 2307
rect 5873 2273 5887 2287
rect 6073 4513 6087 4527
rect 6113 4473 6127 4487
rect 6093 4453 6107 4467
rect 6133 4453 6147 4467
rect 6073 4253 6087 4267
rect 6033 4193 6047 4207
rect 6053 4173 6067 4187
rect 6093 4173 6107 4187
rect 6053 4113 6067 4127
rect 6193 4473 6207 4487
rect 6173 4413 6187 4427
rect 6153 3733 6167 3747
rect 6153 3693 6167 3707
rect 6133 3673 6147 3687
rect 6113 3573 6127 3587
rect 6093 3553 6107 3567
rect 6033 3493 6047 3507
rect 6073 3473 6087 3487
rect 6013 3353 6027 3367
rect 6033 3293 6047 3307
rect 6053 3173 6067 3187
rect 6013 3153 6027 3167
rect 5993 3133 6007 3147
rect 6033 2993 6047 3007
rect 6013 2553 6027 2567
rect 5973 2393 5987 2407
rect 5973 2373 5987 2387
rect 5993 2293 6007 2307
rect 5953 2073 5967 2087
rect 5893 1913 5907 1927
rect 5653 1773 5667 1787
rect 5713 1773 5727 1787
rect 5753 1773 5767 1787
rect 5833 1773 5847 1787
rect 5513 1573 5527 1587
rect 5553 1573 5567 1587
rect 5633 1573 5647 1587
rect 5473 1553 5487 1567
rect 5273 1333 5287 1347
rect 5333 1333 5347 1347
rect 5233 1313 5247 1327
rect 5253 1313 5267 1327
rect 5293 1313 5307 1327
rect 5213 1093 5227 1107
rect 5333 1053 5347 1067
rect 5273 993 5287 1007
rect 5193 873 5207 887
rect 5253 833 5267 847
rect 5173 793 5187 807
rect 5233 793 5247 807
rect 5113 753 5127 767
rect 5093 573 5107 587
rect 4973 413 4987 427
rect 4933 393 4947 407
rect 4993 393 5007 407
rect 4933 373 4947 387
rect 4853 353 4867 367
rect 4313 173 4327 187
rect 4553 173 4567 187
rect 4313 153 4327 167
rect 4353 153 4367 167
rect 4613 153 4627 167
rect 4033 113 4047 127
rect 4093 113 4107 127
rect 4813 173 4827 187
rect 4833 173 4847 187
rect 4953 333 4967 347
rect 5013 313 5027 327
rect 5253 753 5267 767
rect 5193 693 5207 707
rect 5253 673 5267 687
rect 5213 653 5227 667
rect 5313 653 5327 667
rect 5313 333 5327 347
rect 5333 213 5347 227
rect 5093 193 5107 207
rect 5073 173 5087 187
rect 4373 113 4387 127
rect 4593 113 4607 127
rect 4793 113 4807 127
rect 5053 113 5067 127
rect 5113 133 5127 147
rect 5313 133 5327 147
rect 5473 1353 5487 1367
rect 5533 1333 5547 1347
rect 5513 1313 5527 1327
rect 5593 1233 5607 1247
rect 5393 1213 5407 1227
rect 5473 1213 5487 1227
rect 5453 1133 5467 1147
rect 5433 1113 5447 1127
rect 5413 1093 5427 1107
rect 5453 1093 5467 1107
rect 5373 1053 5387 1067
rect 5433 1013 5447 1027
rect 5433 873 5447 887
rect 5513 873 5527 887
rect 5413 813 5427 827
rect 5473 813 5487 827
rect 5573 833 5587 847
rect 5493 793 5507 807
rect 5453 613 5467 627
rect 5653 1133 5667 1147
rect 5593 813 5607 827
rect 5573 733 5587 747
rect 5393 413 5407 427
rect 5473 413 5487 427
rect 5433 373 5447 387
rect 5693 1113 5707 1127
rect 5793 1753 5807 1767
rect 5753 1633 5767 1647
rect 5833 1593 5847 1607
rect 5813 1573 5827 1587
rect 5853 1573 5867 1587
rect 5773 1433 5787 1447
rect 5733 1353 5747 1367
rect 5793 1293 5807 1307
rect 5753 1253 5767 1267
rect 5973 1953 5987 1967
rect 5933 1793 5947 1807
rect 5993 1773 6007 1787
rect 6153 3553 6167 3567
rect 6133 3453 6147 3467
rect 6113 3153 6127 3167
rect 6133 3133 6147 3147
rect 6073 3093 6087 3107
rect 6053 2733 6067 2747
rect 6153 3093 6167 3107
rect 6093 2733 6107 2747
rect 6253 4733 6267 4747
rect 6233 4493 6247 4507
rect 6233 3953 6247 3967
rect 6233 3653 6247 3667
rect 6213 3253 6227 3267
rect 6313 4653 6327 4667
rect 6333 4593 6347 4607
rect 6313 4513 6327 4527
rect 6373 5373 6387 5387
rect 6373 5193 6387 5207
rect 6373 4613 6387 4627
rect 6353 4473 6367 4487
rect 6353 4453 6367 4467
rect 6373 4433 6387 4447
rect 6293 4253 6307 4267
rect 6333 4213 6347 4227
rect 6313 4193 6327 4207
rect 6373 4153 6387 4167
rect 6333 4133 6347 4147
rect 6373 3793 6387 3807
rect 6273 3593 6287 3607
rect 6273 3573 6287 3587
rect 6313 3493 6327 3507
rect 6293 3473 6307 3487
rect 6353 3473 6367 3487
rect 6373 3473 6387 3487
rect 6333 3453 6347 3467
rect 6293 3253 6307 3267
rect 6193 3233 6207 3247
rect 6233 3233 6247 3247
rect 6173 2993 6187 3007
rect 6173 2553 6187 2567
rect 6153 2493 6167 2507
rect 6133 2473 6147 2487
rect 6113 2293 6127 2307
rect 6093 2273 6107 2287
rect 6053 2253 6067 2267
rect 6033 2233 6047 2247
rect 6153 2253 6167 2267
rect 6133 2233 6147 2247
rect 6253 3213 6267 3227
rect 6213 3173 6227 3187
rect 6213 3033 6227 3047
rect 6293 2553 6307 2567
rect 6253 2533 6267 2547
rect 6293 2533 6307 2547
rect 6213 2513 6227 2527
rect 6233 2513 6247 2527
rect 6273 2513 6287 2527
rect 6193 2353 6207 2367
rect 6173 2113 6187 2127
rect 6273 2393 6287 2407
rect 6213 2273 6227 2287
rect 6233 2273 6247 2287
rect 6113 1813 6127 1827
rect 6093 1793 6107 1807
rect 6013 1713 6027 1727
rect 5953 1613 5967 1627
rect 5973 1593 5987 1607
rect 6033 1593 6047 1607
rect 6093 1593 6107 1607
rect 5913 1233 5927 1247
rect 6053 1553 6067 1567
rect 6013 1433 6027 1447
rect 6053 1313 6067 1327
rect 6113 1313 6127 1327
rect 5993 1293 6007 1307
rect 5973 1193 5987 1207
rect 5873 1113 5887 1127
rect 5733 773 5747 787
rect 5713 733 5727 747
rect 5693 713 5707 727
rect 5733 713 5747 727
rect 5693 633 5707 647
rect 5793 793 5807 807
rect 6073 1293 6087 1307
rect 6193 2093 6207 2107
rect 6253 2113 6267 2127
rect 6153 2073 6167 2087
rect 6193 2073 6207 2087
rect 6213 2053 6227 2067
rect 6173 2013 6187 2027
rect 6153 1993 6167 2007
rect 6053 1153 6067 1167
rect 6133 1153 6147 1167
rect 6033 913 6047 927
rect 6013 833 6027 847
rect 6093 1113 6107 1127
rect 6113 1093 6127 1107
rect 6093 833 6107 847
rect 5993 813 6007 827
rect 6033 813 6047 827
rect 6073 793 6087 807
rect 5933 753 5947 767
rect 5993 753 6007 767
rect 5753 673 5767 687
rect 5933 653 5947 667
rect 5753 633 5767 647
rect 5673 613 5687 627
rect 5713 553 5727 567
rect 5613 373 5627 387
rect 5773 573 5787 587
rect 6013 473 6027 487
rect 5953 353 5967 367
rect 5693 333 5707 347
rect 5753 333 5767 347
rect 5913 333 5927 347
rect 5453 313 5467 327
rect 5693 313 5707 327
rect 5493 193 5507 207
rect 5893 313 5907 327
rect 5753 213 5767 227
rect 5513 173 5527 187
rect 5713 173 5727 187
rect 5793 173 5807 187
rect 5533 153 5547 167
rect 5753 153 5767 167
rect 6113 733 6127 747
rect 6113 713 6127 727
rect 6153 693 6167 707
rect 6213 1973 6227 1987
rect 6193 1773 6207 1787
rect 6213 1773 6227 1787
rect 6233 1773 6247 1787
rect 6193 1293 6207 1307
rect 6193 1133 6207 1147
rect 6193 1033 6207 1047
rect 6193 533 6207 547
rect 6133 393 6147 407
rect 6093 373 6107 387
rect 6173 373 6187 387
rect 6033 233 6047 247
rect 5553 113 5567 127
rect 5773 113 5787 127
rect 6293 2253 6307 2267
rect 6293 1093 6307 1107
rect 6273 893 6287 907
rect 6253 853 6267 867
rect 6353 3233 6367 3247
rect 6453 5413 6467 5427
rect 6573 5993 6587 6007
rect 6553 5653 6567 5667
rect 6533 5593 6547 5607
rect 6613 5653 6627 5667
rect 6613 5613 6627 5627
rect 6673 6273 6687 6287
rect 6673 6233 6687 6247
rect 6753 6253 6767 6267
rect 6653 6113 6667 6127
rect 6653 6093 6667 6107
rect 6653 5973 6667 5987
rect 6693 6133 6707 6147
rect 6733 6113 6747 6127
rect 6693 5953 6707 5967
rect 6673 5753 6687 5767
rect 6913 6473 6927 6487
rect 6773 5933 6787 5947
rect 6793 5933 6807 5947
rect 6733 5893 6747 5907
rect 6773 5893 6787 5907
rect 6793 5813 6807 5827
rect 6713 5773 6727 5787
rect 6733 5773 6747 5787
rect 6693 5733 6707 5747
rect 6713 5733 6727 5747
rect 6653 5613 6667 5627
rect 6573 5513 6587 5527
rect 6613 5513 6627 5527
rect 6713 5593 6727 5607
rect 6633 5493 6647 5507
rect 6693 5493 6707 5507
rect 6493 5393 6507 5407
rect 6793 5633 6807 5647
rect 6753 5613 6767 5627
rect 6773 5613 6787 5627
rect 6913 6293 6927 6307
rect 6973 6533 6987 6547
rect 6953 6333 6967 6347
rect 6933 6133 6947 6147
rect 6953 6113 6967 6127
rect 6853 6093 6867 6107
rect 6893 6093 6907 6107
rect 6933 6033 6947 6047
rect 6853 6013 6867 6027
rect 6813 5553 6827 5567
rect 6833 5513 6847 5527
rect 6773 5393 6787 5407
rect 6733 5373 6747 5387
rect 6533 5273 6547 5287
rect 6473 5193 6487 5207
rect 6433 5153 6447 5167
rect 6473 5153 6487 5167
rect 6453 5113 6467 5127
rect 6493 5093 6507 5107
rect 6513 5093 6527 5107
rect 6453 4993 6467 5007
rect 6693 5193 6707 5207
rect 6453 4973 6467 4987
rect 6493 4973 6507 4987
rect 6533 4973 6547 4987
rect 6473 4953 6487 4967
rect 6593 4933 6607 4947
rect 6713 5133 6727 5147
rect 6793 5373 6807 5387
rect 6733 4933 6747 4947
rect 6533 4893 6547 4907
rect 6493 4673 6507 4687
rect 6513 4653 6527 4667
rect 6473 4633 6487 4647
rect 6453 4613 6467 4627
rect 6433 4593 6447 4607
rect 6413 4433 6427 4447
rect 6433 4113 6447 4127
rect 6533 4613 6547 4627
rect 6573 4493 6587 4507
rect 6653 4713 6667 4727
rect 6653 4593 6667 4607
rect 6633 4493 6647 4507
rect 6573 4453 6587 4467
rect 6613 4413 6627 4427
rect 6513 4273 6527 4287
rect 6553 4273 6567 4287
rect 6613 4273 6627 4287
rect 6473 4213 6487 4227
rect 6453 4093 6467 4107
rect 6413 4033 6427 4047
rect 6433 3713 6447 3727
rect 6433 3573 6447 3587
rect 6513 4193 6527 4207
rect 6593 4213 6607 4227
rect 6813 5333 6827 5347
rect 6833 5193 6847 5207
rect 6813 5153 6827 5167
rect 6873 5933 6887 5947
rect 6893 5933 6907 5947
rect 6793 4733 6807 4747
rect 6733 4713 6747 4727
rect 6693 4693 6707 4707
rect 6713 4673 6727 4687
rect 7053 6753 7067 6767
rect 7033 6593 7047 6607
rect 7013 6513 7027 6527
rect 6993 6413 7007 6427
rect 6993 6373 7007 6387
rect 6993 6353 7007 6367
rect 6993 6113 7007 6127
rect 7053 6253 7067 6267
rect 7053 6193 7067 6207
rect 7033 6153 7047 6167
rect 7053 6093 7067 6107
rect 7013 5953 7027 5967
rect 7033 5933 7047 5947
rect 6993 5913 7007 5927
rect 7013 5853 7027 5867
rect 7033 5853 7047 5867
rect 7053 5853 7067 5867
rect 7053 5833 7067 5847
rect 7033 5793 7047 5807
rect 6953 5773 6967 5787
rect 6973 5773 6987 5787
rect 7013 5773 7027 5787
rect 6913 5653 6927 5667
rect 6973 5753 6987 5767
rect 6933 5593 6947 5607
rect 6953 5553 6967 5567
rect 6893 5473 6907 5487
rect 6953 5393 6967 5407
rect 7033 5613 7047 5627
rect 7013 5553 7027 5567
rect 7013 5453 7027 5467
rect 7333 8933 7347 8947
rect 7413 8953 7427 8967
rect 7253 8793 7267 8807
rect 7233 8753 7247 8767
rect 7233 8573 7247 8587
rect 7213 8013 7227 8027
rect 7213 7853 7227 7867
rect 7133 7813 7147 7827
rect 7173 7813 7187 7827
rect 7153 7793 7167 7807
rect 7533 8673 7547 8687
rect 7273 8613 7287 8627
rect 7513 8613 7527 8627
rect 7313 8533 7327 8547
rect 7273 8453 7287 8467
rect 7253 8033 7267 8047
rect 7253 7933 7267 7947
rect 7253 7813 7267 7827
rect 7153 7733 7167 7747
rect 7233 7733 7247 7747
rect 7193 7673 7207 7687
rect 7153 7573 7167 7587
rect 7133 7533 7147 7547
rect 7153 7533 7167 7547
rect 7133 7473 7147 7487
rect 7133 7333 7147 7347
rect 7113 7213 7127 7227
rect 7173 7513 7187 7527
rect 7153 7193 7167 7207
rect 7213 7553 7227 7567
rect 7253 7593 7267 7607
rect 7253 7513 7267 7527
rect 7293 8353 7307 8367
rect 7333 8513 7347 8527
rect 7313 8313 7327 8327
rect 7433 8513 7447 8527
rect 7393 8493 7407 8507
rect 7413 8493 7427 8507
rect 7353 8333 7367 8347
rect 7373 8333 7387 8347
rect 7333 8193 7347 8207
rect 7353 8153 7367 8167
rect 7393 8153 7407 8167
rect 7313 8033 7327 8047
rect 7393 8033 7407 8047
rect 7373 8013 7387 8027
rect 7293 7613 7307 7627
rect 7273 7493 7287 7507
rect 7273 7373 7287 7387
rect 7373 7933 7387 7947
rect 7333 7773 7347 7787
rect 7333 7593 7347 7607
rect 7293 7353 7307 7367
rect 7313 7353 7327 7367
rect 7293 7313 7307 7327
rect 7313 7253 7327 7267
rect 7253 7233 7267 7247
rect 7253 7193 7267 7207
rect 7213 7173 7227 7187
rect 7173 7053 7187 7067
rect 7293 7113 7307 7127
rect 7273 7033 7287 7047
rect 7213 6993 7227 7007
rect 7213 6853 7227 6867
rect 7253 6793 7267 6807
rect 7193 6713 7207 6727
rect 7233 6593 7247 6607
rect 7273 6593 7287 6607
rect 7293 6573 7307 6587
rect 7093 6533 7107 6547
rect 7193 6533 7207 6547
rect 7253 6533 7267 6547
rect 7213 6513 7227 6527
rect 7093 6413 7107 6427
rect 7153 6373 7167 6387
rect 7133 6353 7147 6367
rect 7093 6313 7107 6327
rect 7113 6213 7127 6227
rect 7153 6213 7167 6227
rect 7073 5773 7087 5787
rect 7113 5553 7127 5567
rect 7073 5453 7087 5467
rect 6973 5373 6987 5387
rect 7033 5393 7047 5407
rect 6913 5333 6927 5347
rect 6993 5333 7007 5347
rect 6893 5113 6907 5127
rect 6733 4653 6747 4667
rect 6873 4653 6887 4667
rect 6673 4213 6687 4227
rect 6613 4173 6627 4187
rect 6633 4013 6647 4027
rect 6673 4013 6687 4027
rect 6653 3993 6667 4007
rect 6533 3973 6547 3987
rect 6533 3953 6547 3967
rect 6513 3853 6527 3867
rect 6493 3513 6507 3527
rect 6473 3413 6487 3427
rect 6453 3233 6467 3247
rect 6473 3233 6487 3247
rect 6493 3213 6507 3227
rect 6373 3053 6387 3067
rect 6413 3053 6427 3067
rect 6453 3053 6467 3067
rect 6393 3033 6407 3047
rect 6373 2753 6387 2767
rect 6333 2733 6347 2747
rect 6333 2633 6347 2647
rect 6413 2713 6427 2727
rect 6393 2573 6407 2587
rect 6353 2553 6367 2567
rect 6353 2513 6367 2527
rect 6393 2513 6407 2527
rect 6333 1773 6347 1787
rect 6333 1273 6347 1287
rect 6393 2233 6407 2247
rect 6433 2233 6447 2247
rect 6413 2093 6427 2107
rect 6433 2073 6447 2087
rect 6393 2033 6407 2047
rect 6413 1973 6427 1987
rect 6493 2573 6507 2587
rect 6653 3753 6667 3767
rect 6613 3733 6627 3747
rect 6633 3713 6647 3727
rect 6693 3993 6707 4007
rect 6673 3733 6687 3747
rect 6553 3693 6567 3707
rect 6593 3693 6607 3707
rect 6653 3693 6667 3707
rect 6573 3533 6587 3547
rect 6533 3513 6547 3527
rect 6573 3413 6587 3427
rect 6553 3253 6567 3267
rect 6533 3233 6547 3247
rect 6513 2553 6527 2567
rect 6513 2513 6527 2527
rect 6473 2493 6487 2507
rect 6493 2333 6507 2347
rect 6713 3973 6727 3987
rect 6693 3673 6707 3687
rect 6613 3033 6627 3047
rect 6653 3033 6667 3047
rect 6633 3013 6647 3027
rect 6593 2993 6607 3007
rect 6613 2793 6627 2807
rect 6653 2793 6667 2807
rect 6653 2773 6667 2787
rect 6593 2733 6607 2747
rect 6633 2713 6647 2727
rect 6713 3273 6727 3287
rect 6853 4593 6867 4607
rect 6873 4553 6887 4567
rect 6773 4353 6787 4367
rect 6793 4253 6807 4267
rect 6773 4153 6787 4167
rect 6753 3633 6767 3647
rect 6733 3253 6747 3267
rect 6713 3213 6727 3227
rect 6733 3193 6747 3207
rect 6773 3593 6787 3607
rect 6813 4013 6827 4027
rect 6953 5153 6967 5167
rect 6993 5153 7007 5167
rect 7033 5153 7047 5167
rect 7013 5133 7027 5147
rect 6973 5093 6987 5107
rect 6953 4933 6967 4947
rect 6973 4913 6987 4927
rect 6933 4893 6947 4907
rect 6973 4693 6987 4707
rect 7033 4993 7047 5007
rect 7093 5013 7107 5027
rect 7073 4913 7087 4927
rect 7033 4693 7047 4707
rect 6993 4653 7007 4667
rect 7013 4653 7027 4667
rect 6973 4433 6987 4447
rect 7073 4493 7087 4507
rect 7053 4473 7067 4487
rect 7053 4433 7067 4447
rect 7033 4413 7047 4427
rect 6993 4153 7007 4167
rect 7013 4153 7027 4167
rect 7033 4113 7047 4127
rect 6933 4013 6947 4027
rect 6993 4013 7007 4027
rect 6933 3993 6947 4007
rect 6953 3993 6967 4007
rect 6913 3933 6927 3947
rect 6853 3833 6867 3847
rect 6893 3753 6907 3767
rect 6873 3693 6887 3707
rect 6853 3673 6867 3687
rect 6853 3613 6867 3627
rect 6833 3593 6847 3607
rect 6793 3533 6807 3547
rect 6793 3493 6807 3507
rect 6793 3113 6807 3127
rect 6773 2793 6787 2807
rect 6753 2753 6767 2767
rect 6753 2573 6767 2587
rect 6593 2373 6607 2387
rect 6593 2313 6607 2327
rect 6553 2293 6567 2307
rect 6553 2273 6567 2287
rect 6593 2093 6607 2107
rect 6533 2073 6547 2087
rect 6493 1993 6507 2007
rect 6453 1813 6467 1827
rect 6473 1813 6487 1827
rect 6453 1793 6467 1807
rect 6533 1793 6547 1807
rect 6473 1773 6487 1787
rect 6493 1773 6507 1787
rect 6493 1573 6507 1587
rect 6513 1553 6527 1567
rect 6433 1533 6447 1547
rect 6473 1533 6487 1547
rect 6413 1293 6427 1307
rect 6453 1293 6467 1307
rect 6353 1153 6367 1167
rect 6433 1153 6447 1167
rect 6413 1133 6427 1147
rect 6373 1113 6387 1127
rect 6393 1073 6407 1087
rect 6353 1013 6367 1027
rect 6353 973 6367 987
rect 6353 893 6367 907
rect 6333 793 6347 807
rect 6293 773 6307 787
rect 6233 333 6247 347
rect 6253 173 6267 187
rect 6153 153 6167 167
rect 6053 133 6067 147
rect 6273 93 6287 107
rect 6073 73 6087 87
rect 6573 1293 6587 1307
rect 6533 1273 6547 1287
rect 6633 2253 6647 2267
rect 6613 2073 6627 2087
rect 6633 1753 6647 1767
rect 6613 1693 6627 1707
rect 6633 1553 6647 1567
rect 6593 1173 6607 1187
rect 6733 2553 6747 2567
rect 6713 2533 6727 2547
rect 6673 2513 6687 2527
rect 6693 2513 6707 2527
rect 6693 2273 6707 2287
rect 6673 2253 6687 2267
rect 6753 2133 6767 2147
rect 6733 2093 6747 2107
rect 6713 2073 6727 2087
rect 6673 1813 6687 1827
rect 6753 1773 6767 1787
rect 6713 1593 6727 1607
rect 6733 1553 6747 1567
rect 6813 3073 6827 3087
rect 6853 3293 6867 3307
rect 6833 3053 6847 3067
rect 6953 3693 6967 3707
rect 6913 3653 6927 3667
rect 7033 3533 7047 3547
rect 6973 3513 6987 3527
rect 7013 3513 7027 3527
rect 6913 3273 6927 3287
rect 6893 3233 6907 3247
rect 6873 3053 6887 3067
rect 6833 2753 6847 2767
rect 6813 2713 6827 2727
rect 6793 2533 6807 2547
rect 6893 2553 6907 2567
rect 6873 2333 6887 2347
rect 6833 2293 6847 2307
rect 6813 2253 6827 2267
rect 6813 2173 6827 2187
rect 6773 1633 6787 1647
rect 6773 1593 6787 1607
rect 6873 2253 6887 2267
rect 6933 3233 6947 3247
rect 6973 3233 6987 3247
rect 7013 3233 7027 3247
rect 6953 3193 6967 3207
rect 6933 3093 6947 3107
rect 6913 2533 6927 2547
rect 6993 3073 7007 3087
rect 7013 2953 7027 2967
rect 6973 2793 6987 2807
rect 6993 2773 7007 2787
rect 7073 4413 7087 4427
rect 7073 4153 7087 4167
rect 7173 6153 7187 6167
rect 7193 6153 7207 6167
rect 7173 6113 7187 6127
rect 7193 6013 7207 6027
rect 7173 5973 7187 5987
rect 7353 7553 7367 7567
rect 7333 6853 7347 6867
rect 7313 6313 7327 6327
rect 7453 8153 7467 8167
rect 7433 7913 7447 7927
rect 7433 7853 7447 7867
rect 7393 7813 7407 7827
rect 7393 7793 7407 7807
rect 7373 7453 7387 7467
rect 7493 8053 7507 8067
rect 7453 7593 7467 7607
rect 7433 7533 7447 7547
rect 7533 8513 7547 8527
rect 7653 9033 7667 9047
rect 7593 8933 7607 8947
rect 7573 8773 7587 8787
rect 7573 8673 7587 8687
rect 7573 8493 7587 8507
rect 7633 8773 7647 8787
rect 7873 9873 7887 9887
rect 7873 9853 7887 9867
rect 7853 9673 7867 9687
rect 7853 9453 7867 9467
rect 7793 9373 7807 9387
rect 7833 9373 7847 9387
rect 7753 9333 7767 9347
rect 7713 9273 7727 9287
rect 7733 9233 7747 9247
rect 7693 9213 7707 9227
rect 7713 9153 7727 9167
rect 7693 9093 7707 9107
rect 7673 8613 7687 8627
rect 7653 8593 7667 8607
rect 7613 8533 7627 8547
rect 7653 8513 7667 8527
rect 7673 8493 7687 8507
rect 7633 8453 7647 8467
rect 7593 8413 7607 8427
rect 7633 8413 7647 8427
rect 7573 8393 7587 8407
rect 7613 8393 7627 8407
rect 7553 8313 7567 8327
rect 7593 8373 7607 8387
rect 7613 8333 7627 8347
rect 7673 8333 7687 8347
rect 7573 8193 7587 8207
rect 7613 8073 7627 8087
rect 7573 8013 7587 8027
rect 7593 8013 7607 8027
rect 7613 7973 7627 7987
rect 7633 7913 7647 7927
rect 7613 7853 7627 7867
rect 7653 7833 7667 7847
rect 7593 7813 7607 7827
rect 7633 7813 7647 7827
rect 7513 7793 7527 7807
rect 7513 7753 7527 7767
rect 7573 7733 7587 7747
rect 7413 7493 7427 7507
rect 7473 7493 7487 7507
rect 7493 7493 7507 7507
rect 7493 7373 7507 7387
rect 7453 7353 7467 7367
rect 7413 7113 7427 7127
rect 7473 7333 7487 7347
rect 7513 7233 7527 7247
rect 7493 7073 7507 7087
rect 7493 7033 7507 7047
rect 7433 6893 7447 6907
rect 7473 6873 7487 6887
rect 7453 6853 7467 6867
rect 7413 6773 7427 6787
rect 7453 6653 7467 6667
rect 7533 7013 7547 7027
rect 7513 6873 7527 6887
rect 7553 6893 7567 6907
rect 7533 6853 7547 6867
rect 7513 6633 7527 6647
rect 7493 6613 7507 6627
rect 7393 6513 7407 6527
rect 7413 6453 7427 6467
rect 7373 6433 7387 6447
rect 7353 6013 7367 6027
rect 7353 5973 7367 5987
rect 7213 5853 7227 5867
rect 7193 5793 7207 5807
rect 7313 5793 7327 5807
rect 7353 5773 7367 5787
rect 7333 5633 7347 5647
rect 7293 5553 7307 5567
rect 7273 5453 7287 5467
rect 7153 5433 7167 5447
rect 7313 5433 7327 5447
rect 7253 5353 7267 5367
rect 7193 5193 7207 5207
rect 7233 5153 7247 5167
rect 7173 5133 7187 5147
rect 7133 5113 7147 5127
rect 7173 5113 7187 5127
rect 7213 5113 7227 5127
rect 7133 4953 7147 4967
rect 7133 4433 7147 4447
rect 7193 4913 7207 4927
rect 7193 4873 7207 4887
rect 7193 4653 7207 4667
rect 7173 4513 7187 4527
rect 7133 4013 7147 4027
rect 7153 4013 7167 4027
rect 7113 3853 7127 3867
rect 7073 3773 7087 3787
rect 7153 3973 7167 3987
rect 7133 3753 7147 3767
rect 7073 3733 7087 3747
rect 7113 3733 7127 3747
rect 7133 3713 7147 3727
rect 7093 3693 7107 3707
rect 7113 3573 7127 3587
rect 7133 3573 7147 3587
rect 7093 3513 7107 3527
rect 7113 3513 7127 3527
rect 7073 3493 7087 3507
rect 7053 3093 7067 3107
rect 7053 3073 7067 3087
rect 7093 3453 7107 3467
rect 7093 3293 7107 3307
rect 7073 3053 7087 3067
rect 7093 3033 7107 3047
rect 7133 3033 7147 3047
rect 6993 2733 7007 2747
rect 7113 2753 7127 2767
rect 7033 2733 7047 2747
rect 7073 2733 7087 2747
rect 7053 2673 7067 2687
rect 7013 2553 7027 2567
rect 6993 2533 7007 2547
rect 6953 2513 6967 2527
rect 6993 2133 7007 2147
rect 6933 2113 6947 2127
rect 6933 2093 6947 2107
rect 6973 2093 6987 2107
rect 6893 2053 6907 2067
rect 7013 2113 7027 2127
rect 6933 2033 6947 2047
rect 6933 1773 6947 1787
rect 6893 1713 6907 1727
rect 6953 1673 6967 1687
rect 6993 1633 7007 1647
rect 6973 1613 6987 1627
rect 6853 1373 6867 1387
rect 6833 1333 6847 1347
rect 6993 1333 7007 1347
rect 6753 1293 6767 1307
rect 6693 1213 6707 1227
rect 6713 1173 6727 1187
rect 6653 1153 6667 1167
rect 6693 1153 6707 1167
rect 6673 1133 6687 1147
rect 6573 1113 6587 1127
rect 6633 1113 6647 1127
rect 6533 1093 6547 1107
rect 6553 1093 6567 1107
rect 6573 1053 6587 1067
rect 6553 1013 6567 1027
rect 6493 793 6507 807
rect 6653 1093 6667 1107
rect 6693 1093 6707 1107
rect 6613 973 6627 987
rect 6673 773 6687 787
rect 6633 753 6647 767
rect 6353 13 6367 27
rect 6413 333 6427 347
rect 6653 673 6667 687
rect 6813 1153 6827 1167
rect 6813 1113 6827 1127
rect 6813 1033 6827 1047
rect 6733 793 6747 807
rect 6753 793 6767 807
rect 6773 773 6787 787
rect 6933 1133 6947 1147
rect 6853 1113 6867 1127
rect 6893 1113 6907 1127
rect 6913 1093 6927 1107
rect 6873 973 6887 987
rect 7013 1093 7027 1107
rect 7053 2553 7067 2567
rect 7073 2533 7087 2547
rect 7193 4473 7207 4487
rect 7193 3753 7207 3767
rect 7173 3573 7187 3587
rect 7233 4253 7247 4267
rect 7273 5293 7287 5307
rect 7273 5133 7287 5147
rect 7273 4433 7287 4447
rect 7253 4233 7267 4247
rect 7273 4213 7287 4227
rect 7253 4193 7267 4207
rect 7233 3733 7247 3747
rect 7233 3653 7247 3667
rect 7393 6373 7407 6387
rect 7433 6353 7447 6367
rect 7493 6393 7507 6407
rect 7473 6153 7487 6167
rect 7393 6113 7407 6127
rect 7433 6113 7447 6127
rect 7533 6573 7547 6587
rect 7553 6553 7567 6567
rect 7513 6373 7527 6387
rect 7533 6333 7547 6347
rect 7493 6113 7507 6127
rect 7493 5993 7507 6007
rect 7413 5973 7427 5987
rect 7513 5753 7527 5767
rect 7493 5713 7507 5727
rect 7453 5653 7467 5667
rect 7433 5633 7447 5647
rect 7393 5593 7407 5607
rect 7433 5573 7447 5587
rect 7373 5553 7387 5567
rect 7433 5513 7447 5527
rect 7453 5353 7467 5367
rect 7473 5273 7487 5287
rect 7433 5213 7447 5227
rect 7353 5153 7367 5167
rect 7413 5153 7427 5167
rect 7453 5153 7467 5167
rect 7373 5053 7387 5067
rect 7433 5113 7447 5127
rect 7433 5033 7447 5047
rect 7393 4953 7407 4967
rect 7393 4693 7407 4707
rect 7393 4653 7407 4667
rect 7413 4653 7427 4667
rect 7453 4653 7467 4667
rect 7433 4633 7447 4647
rect 7373 4453 7387 4467
rect 7333 4433 7347 4447
rect 7313 4093 7327 4107
rect 7353 4013 7367 4027
rect 7313 3993 7327 4007
rect 7393 4293 7407 4307
rect 7373 3973 7387 3987
rect 7373 3913 7387 3927
rect 7293 3693 7307 3707
rect 7333 3693 7347 3707
rect 7313 3673 7327 3687
rect 7253 3633 7267 3647
rect 7213 3593 7227 3607
rect 7313 3593 7327 3607
rect 7193 3553 7207 3567
rect 7253 3553 7267 3567
rect 7293 3553 7307 3567
rect 7213 3513 7227 3527
rect 7233 3473 7247 3487
rect 7273 3453 7287 3467
rect 7233 3213 7247 3227
rect 7193 3173 7207 3187
rect 7173 2993 7187 3007
rect 7173 2733 7187 2747
rect 7153 2713 7167 2727
rect 7173 2553 7187 2567
rect 7133 2533 7147 2547
rect 7113 2513 7127 2527
rect 7133 2333 7147 2347
rect 7093 2273 7107 2287
rect 7113 2253 7127 2267
rect 7153 2253 7167 2267
rect 7373 3513 7387 3527
rect 7433 4273 7447 4287
rect 7413 4213 7427 4227
rect 7433 4213 7447 4227
rect 7413 3353 7427 3367
rect 7733 8453 7747 8467
rect 7713 7993 7727 8007
rect 7773 8873 7787 8887
rect 7753 8213 7767 8227
rect 7753 7953 7767 7967
rect 7733 7733 7747 7747
rect 7673 7693 7687 7707
rect 7693 7693 7707 7707
rect 7633 7593 7647 7607
rect 7593 7553 7607 7567
rect 7653 7553 7667 7567
rect 7733 7553 7747 7567
rect 7633 7533 7647 7547
rect 7713 7533 7727 7547
rect 7673 7513 7687 7527
rect 7573 6073 7587 6087
rect 7553 5993 7567 6007
rect 7533 5513 7547 5527
rect 7533 5453 7547 5467
rect 7513 5393 7527 5407
rect 7573 5973 7587 5987
rect 7733 7333 7747 7347
rect 7653 7313 7667 7327
rect 7633 7133 7647 7147
rect 7613 6933 7627 6947
rect 7673 7033 7687 7047
rect 7713 7033 7727 7047
rect 7693 7013 7707 7027
rect 7713 6833 7727 6847
rect 7673 6673 7687 6687
rect 7693 6553 7707 6567
rect 7773 7013 7787 7027
rect 7753 6873 7767 6887
rect 7773 6593 7787 6607
rect 7753 6553 7767 6567
rect 7653 6393 7667 6407
rect 7673 6373 7687 6387
rect 7713 6333 7727 6347
rect 7713 6313 7727 6327
rect 7633 6213 7647 6227
rect 7633 6153 7647 6167
rect 7613 6133 7627 6147
rect 7673 6113 7687 6127
rect 7653 6093 7667 6107
rect 7653 6073 7667 6087
rect 7613 5973 7627 5987
rect 7613 5933 7627 5947
rect 7613 5893 7627 5907
rect 7593 5633 7607 5647
rect 7633 5633 7647 5647
rect 7693 5953 7707 5967
rect 7713 5933 7727 5947
rect 7733 5913 7747 5927
rect 7693 5873 7707 5887
rect 7673 5733 7687 5747
rect 7653 5613 7667 5627
rect 7893 9733 7907 9747
rect 8173 10453 8187 10467
rect 8213 10433 8227 10447
rect 8013 10233 8027 10247
rect 7973 10153 7987 10167
rect 7953 9893 7967 9907
rect 7973 9853 7987 9867
rect 8193 10253 8207 10267
rect 8153 10233 8167 10247
rect 8173 10213 8187 10227
rect 8113 9973 8127 9987
rect 8093 9853 8107 9867
rect 8013 9833 8027 9847
rect 7993 9733 8007 9747
rect 8213 9733 8227 9747
rect 7953 9633 7967 9647
rect 7933 9473 7947 9487
rect 7913 9333 7927 9347
rect 8193 9653 8207 9667
rect 8073 9513 8087 9527
rect 8013 9473 8027 9487
rect 7873 9233 7887 9247
rect 7873 9073 7887 9087
rect 7933 9033 7947 9047
rect 7853 8993 7867 9007
rect 7813 8973 7827 8987
rect 7893 8973 7907 8987
rect 7873 8753 7887 8767
rect 7953 8613 7967 8627
rect 7873 8533 7887 8547
rect 7853 8513 7867 8527
rect 7913 8513 7927 8527
rect 7853 8433 7867 8447
rect 7893 8313 7907 8327
rect 7953 8313 7967 8327
rect 7893 8293 7907 8307
rect 7873 8173 7887 8187
rect 7833 8033 7847 8047
rect 7833 7993 7847 8007
rect 7813 7973 7827 7987
rect 7813 7513 7827 7527
rect 7813 6933 7827 6947
rect 7913 8233 7927 8247
rect 7933 8213 7947 8227
rect 7933 8013 7947 8027
rect 7933 7913 7947 7927
rect 7853 7853 7867 7867
rect 7873 7853 7887 7867
rect 7893 7853 7907 7867
rect 7873 7833 7887 7847
rect 7993 9013 8007 9027
rect 8153 9473 8167 9487
rect 8073 9033 8087 9047
rect 8173 9033 8187 9047
rect 8033 8953 8047 8967
rect 8093 9013 8107 9027
rect 8113 8993 8127 9007
rect 8113 8973 8127 8987
rect 8393 10913 8407 10927
rect 8353 10753 8367 10767
rect 8353 10713 8367 10727
rect 8313 10693 8327 10707
rect 8293 10493 8307 10507
rect 8313 10453 8327 10467
rect 8253 9833 8267 9847
rect 8233 9633 8247 9647
rect 8213 9453 8227 9467
rect 8213 9293 8227 9307
rect 8233 9073 8247 9087
rect 8193 8993 8207 9007
rect 8293 9753 8307 9767
rect 8273 9493 8287 9507
rect 8293 9253 8307 9267
rect 8273 9033 8287 9047
rect 8253 8973 8267 8987
rect 8273 8973 8287 8987
rect 8153 8853 8167 8867
rect 8073 8753 8087 8767
rect 8133 8773 8147 8787
rect 8173 8753 8187 8767
rect 8033 8713 8047 8727
rect 8033 8593 8047 8607
rect 7973 8253 7987 8267
rect 7993 8253 8007 8267
rect 7913 7793 7927 7807
rect 7953 7553 7967 7567
rect 7913 7533 7927 7547
rect 7933 7533 7947 7547
rect 7973 7513 7987 7527
rect 7953 7493 7967 7507
rect 7873 7473 7887 7487
rect 7873 7413 7887 7427
rect 7913 7393 7927 7407
rect 7953 7353 7967 7367
rect 7933 7333 7947 7347
rect 7933 7313 7947 7327
rect 7853 7193 7867 7207
rect 7893 7113 7907 7127
rect 7853 7033 7867 7047
rect 7833 6733 7847 6747
rect 7833 6633 7847 6647
rect 7813 6593 7827 6607
rect 7813 6513 7827 6527
rect 7813 6493 7827 6507
rect 7813 6353 7827 6367
rect 7733 5793 7747 5807
rect 7753 5793 7767 5807
rect 7613 5593 7627 5607
rect 7693 5593 7707 5607
rect 7593 5473 7607 5487
rect 7573 5433 7587 5447
rect 7573 5233 7587 5247
rect 7553 5173 7567 5187
rect 7533 4913 7547 4927
rect 7493 4593 7507 4607
rect 7513 4493 7527 4507
rect 7573 4673 7587 4687
rect 7573 4553 7587 4567
rect 7553 4473 7567 4487
rect 7533 4453 7547 4467
rect 7473 4213 7487 4227
rect 7493 4153 7507 4167
rect 7533 4153 7547 4167
rect 7793 5733 7807 5747
rect 7773 5673 7787 5687
rect 7693 5393 7707 5407
rect 7713 5393 7727 5407
rect 7753 5393 7767 5407
rect 7613 5353 7627 5367
rect 7633 5213 7647 5227
rect 7653 5173 7667 5187
rect 7673 5053 7687 5067
rect 7653 5013 7667 5027
rect 7753 4953 7767 4967
rect 7673 4933 7687 4947
rect 7733 4933 7747 4947
rect 7633 4853 7647 4867
rect 7633 4633 7647 4647
rect 7673 4633 7687 4647
rect 7693 4613 7707 4627
rect 7653 4473 7667 4487
rect 7673 4473 7687 4487
rect 7653 4413 7667 4427
rect 7613 4373 7627 4387
rect 7573 4133 7587 4147
rect 7513 4093 7527 4107
rect 7593 4033 7607 4047
rect 7473 4013 7487 4027
rect 7513 4013 7527 4027
rect 7473 3973 7487 3987
rect 7453 3933 7467 3947
rect 7453 3793 7467 3807
rect 7453 3473 7467 3487
rect 7533 3993 7547 4007
rect 7513 3953 7527 3967
rect 7513 3853 7527 3867
rect 7633 4253 7647 4267
rect 7633 3973 7647 3987
rect 7573 3953 7587 3967
rect 7653 3953 7667 3967
rect 7533 3793 7547 3807
rect 7533 3713 7547 3727
rect 7513 3673 7527 3687
rect 7553 3673 7567 3687
rect 7513 3573 7527 3587
rect 7433 3253 7447 3267
rect 7353 3233 7367 3247
rect 7373 3233 7387 3247
rect 7313 3213 7327 3227
rect 7293 3113 7307 3127
rect 7373 3073 7387 3087
rect 7333 3033 7347 3047
rect 7353 2953 7367 2967
rect 7273 2753 7287 2767
rect 7293 2733 7307 2747
rect 7213 2613 7227 2627
rect 7253 2553 7267 2567
rect 7233 2533 7247 2547
rect 7293 2273 7307 2287
rect 7193 2253 7207 2267
rect 7353 2713 7367 2727
rect 7393 2353 7407 2367
rect 7353 2273 7367 2287
rect 7413 2313 7427 2327
rect 7373 2253 7387 2267
rect 7413 2233 7427 2247
rect 7313 2133 7327 2147
rect 7173 2113 7187 2127
rect 7213 2113 7227 2127
rect 7253 2113 7267 2127
rect 7173 2073 7187 2087
rect 7193 2053 7207 2067
rect 7533 3473 7547 3487
rect 7553 3393 7567 3407
rect 7553 3333 7567 3347
rect 7473 3253 7487 3267
rect 7573 3173 7587 3187
rect 7533 3153 7547 3167
rect 7573 3093 7587 3107
rect 7553 3033 7567 3047
rect 7613 3033 7627 3047
rect 7533 3013 7547 3027
rect 7593 3013 7607 3027
rect 7753 4873 7767 4887
rect 7753 4673 7767 4687
rect 7733 4633 7747 4647
rect 7753 4513 7767 4527
rect 7733 4493 7747 4507
rect 7913 6953 7927 6967
rect 7933 6893 7947 6907
rect 7973 6873 7987 6887
rect 7993 6853 8007 6867
rect 7953 6813 7967 6827
rect 8233 8633 8247 8647
rect 8093 8573 8107 8587
rect 8173 8573 8187 8587
rect 8193 8513 8207 8527
rect 8153 8493 8167 8507
rect 8173 8493 8187 8507
rect 8213 8493 8227 8507
rect 8213 8373 8227 8387
rect 8193 8353 8207 8367
rect 8113 8333 8127 8347
rect 8153 8313 8167 8327
rect 8073 8293 8087 8307
rect 8093 8293 8107 8307
rect 8133 8293 8147 8307
rect 8173 8293 8187 8307
rect 8213 8293 8227 8307
rect 8133 8113 8147 8127
rect 8093 8073 8107 8087
rect 8053 8033 8067 8047
rect 8113 8013 8127 8027
rect 8073 7993 8087 8007
rect 8033 7653 8047 7667
rect 8013 6753 8027 6767
rect 7973 6613 7987 6627
rect 7893 6573 7907 6587
rect 7953 6573 7967 6587
rect 7953 6553 7967 6567
rect 8013 6553 8027 6567
rect 8093 7813 8107 7827
rect 8213 8033 8227 8047
rect 8193 8013 8207 8027
rect 8153 7873 8167 7887
rect 8193 7833 8207 7847
rect 8173 7813 8187 7827
rect 8113 7793 8127 7807
rect 8093 7313 8107 7327
rect 8073 7273 8087 7287
rect 7993 6393 8007 6407
rect 7933 6373 7947 6387
rect 7973 6373 7987 6387
rect 7893 6353 7907 6367
rect 7853 6333 7867 6347
rect 7973 6233 7987 6247
rect 7993 6233 8007 6247
rect 7853 6113 7867 6127
rect 7853 6053 7867 6067
rect 7833 5933 7847 5947
rect 7833 5913 7847 5927
rect 7833 5873 7847 5887
rect 7913 6113 7927 6127
rect 7893 6093 7907 6107
rect 7873 6033 7887 6047
rect 7953 6073 7967 6087
rect 7933 6053 7947 6067
rect 7933 5853 7947 5867
rect 7933 5833 7947 5847
rect 7913 5813 7927 5827
rect 7853 5713 7867 5727
rect 7913 5653 7927 5667
rect 7873 5633 7887 5647
rect 7853 5613 7867 5627
rect 7893 5513 7907 5527
rect 7833 5493 7847 5507
rect 7893 5493 7907 5507
rect 7873 5453 7887 5467
rect 7833 5433 7847 5447
rect 7873 5413 7887 5427
rect 7793 4753 7807 4767
rect 7793 4733 7807 4747
rect 7853 5173 7867 5187
rect 7853 5093 7867 5107
rect 7853 4913 7867 4927
rect 7953 5613 7967 5627
rect 7933 5473 7947 5487
rect 8033 6153 8047 6167
rect 8093 6893 8107 6907
rect 8073 6853 8087 6867
rect 8133 7653 8147 7667
rect 8253 8513 8267 8527
rect 8233 7973 8247 7987
rect 8273 8473 8287 8487
rect 8673 11193 8687 11207
rect 8713 11193 8727 11207
rect 8653 11173 8667 11187
rect 8693 11153 8707 11167
rect 8473 11133 8487 11147
rect 8633 11113 8647 11127
rect 8573 11093 8587 11107
rect 8573 10833 8587 10847
rect 8613 10833 8627 10847
rect 8513 10733 8527 10747
rect 8553 10713 8567 10727
rect 8453 10693 8467 10707
rect 8533 10693 8547 10707
rect 8373 10453 8387 10467
rect 8353 10433 8367 10447
rect 8393 10413 8407 10427
rect 8333 10213 8347 10227
rect 8373 10213 8387 10227
rect 8393 10193 8407 10207
rect 8433 10193 8447 10207
rect 8553 10433 8567 10447
rect 8493 10413 8507 10427
rect 8933 11173 8947 11187
rect 8973 11193 8987 11207
rect 9153 11193 9167 11207
rect 8853 11133 8867 11147
rect 8893 11133 8907 11147
rect 8953 11133 8967 11147
rect 8813 10913 8827 10927
rect 8773 10733 8787 10747
rect 8733 10713 8747 10727
rect 8793 10693 8807 10707
rect 8993 11173 9007 11187
rect 9613 11193 9627 11207
rect 10113 11193 10127 11207
rect 9393 11173 9407 11187
rect 9613 11173 9627 11187
rect 9653 11173 9667 11187
rect 9693 11173 9707 11187
rect 9873 11173 9887 11187
rect 9213 11153 9227 11167
rect 9133 11133 9147 11147
rect 9093 10913 9107 10927
rect 9133 10913 9147 10927
rect 9173 10913 9187 10927
rect 9333 10913 9347 10927
rect 9413 11133 9427 11147
rect 9673 11133 9687 11147
rect 9393 11113 9407 11127
rect 9113 10893 9127 10907
rect 9133 10873 9147 10887
rect 9073 10733 9087 10747
rect 8993 10713 9007 10727
rect 9033 10713 9047 10727
rect 8933 10693 8947 10707
rect 8973 10693 8987 10707
rect 8693 10673 8707 10687
rect 8633 10333 8647 10347
rect 8733 10333 8747 10347
rect 8573 10313 8587 10327
rect 8573 10233 8587 10247
rect 8693 10313 8707 10327
rect 8673 10233 8687 10247
rect 8613 10213 8627 10227
rect 8653 10213 8667 10227
rect 8573 10193 8587 10207
rect 8353 10173 8367 10187
rect 8453 10173 8467 10187
rect 8433 9973 8447 9987
rect 8413 9893 8427 9907
rect 8353 9753 8367 9767
rect 8413 9733 8427 9747
rect 8333 9693 8347 9707
rect 8353 9453 8367 9467
rect 8393 9413 8407 9427
rect 8413 9273 8427 9287
rect 8393 9253 8407 9267
rect 8373 9233 8387 9247
rect 8413 9173 8427 9187
rect 8333 9013 8347 9027
rect 8353 8953 8367 8967
rect 8393 8973 8407 8987
rect 8353 8933 8367 8947
rect 8373 8933 8387 8947
rect 8413 8933 8427 8947
rect 8553 9953 8567 9967
rect 8593 9933 8607 9947
rect 8593 9773 8607 9787
rect 8453 9693 8467 9707
rect 8633 9633 8647 9647
rect 8533 9333 8547 9347
rect 8453 9293 8467 9307
rect 8433 8913 8447 8927
rect 8353 8873 8367 8887
rect 8393 8853 8407 8867
rect 8353 8813 8367 8827
rect 8473 9273 8487 9287
rect 8513 9273 8527 9287
rect 8613 9453 8627 9467
rect 8593 9433 8607 9447
rect 8493 9233 8507 9247
rect 8573 9233 8587 9247
rect 8473 9093 8487 9107
rect 8573 9093 8587 9107
rect 8453 8793 8467 8807
rect 8533 9073 8547 9087
rect 8513 9013 8527 9027
rect 8513 8973 8527 8987
rect 8513 8933 8527 8947
rect 8333 8773 8347 8787
rect 8353 8773 8367 8787
rect 8373 8773 8387 8787
rect 8473 8773 8487 8787
rect 8493 8653 8507 8667
rect 8453 8613 8467 8627
rect 8393 8513 8407 8527
rect 8473 8573 8487 8587
rect 8373 8493 8387 8507
rect 8413 8493 8427 8507
rect 8353 8273 8367 8287
rect 8313 8173 8327 8187
rect 8273 8093 8287 8107
rect 8333 8033 8347 8047
rect 8433 8453 8447 8467
rect 8393 8333 8407 8347
rect 8413 8293 8427 8307
rect 8453 8293 8467 8307
rect 8433 8273 8447 8287
rect 8313 7993 8327 8007
rect 8353 7913 8367 7927
rect 8273 7833 8287 7847
rect 8253 7813 8267 7827
rect 8253 7613 8267 7627
rect 8153 7533 8167 7547
rect 8153 7493 8167 7507
rect 8213 7553 8227 7567
rect 8173 7473 8187 7487
rect 8233 7533 8247 7547
rect 8193 7453 8207 7467
rect 8133 7373 8147 7387
rect 8173 7373 8187 7387
rect 8233 7373 8247 7387
rect 8233 7353 8247 7367
rect 8313 7573 8327 7587
rect 8293 7553 8307 7567
rect 8273 7533 8287 7547
rect 8133 7133 8147 7147
rect 8213 7333 8227 7347
rect 8253 7333 8267 7347
rect 8253 7233 8267 7247
rect 8173 7133 8187 7147
rect 8153 7113 8167 7127
rect 8153 7073 8167 7087
rect 8133 7033 8147 7047
rect 8133 6993 8147 7007
rect 8213 7053 8227 7067
rect 8413 7853 8427 7867
rect 8393 7813 8407 7827
rect 8433 7813 8447 7827
rect 8433 7633 8447 7647
rect 8413 7613 8427 7627
rect 8453 7573 8467 7587
rect 8433 7553 8447 7567
rect 8353 7513 8367 7527
rect 8473 7473 8487 7487
rect 8293 7213 8307 7227
rect 8273 7073 8287 7087
rect 8133 6853 8147 6867
rect 8193 6853 8207 6867
rect 8133 6833 8147 6847
rect 8113 6793 8127 6807
rect 8093 6413 8107 6427
rect 8233 6833 8247 6847
rect 8233 6793 8247 6807
rect 8193 6713 8207 6727
rect 8253 6713 8267 6727
rect 8153 6553 8167 6567
rect 8213 6393 8227 6407
rect 8193 6373 8207 6387
rect 8133 6233 8147 6247
rect 8193 6213 8207 6227
rect 8173 6133 8187 6147
rect 8093 6113 8107 6127
rect 8113 6113 8127 6127
rect 8073 6093 8087 6107
rect 8053 6073 8067 6087
rect 8013 5913 8027 5927
rect 8033 5693 8047 5707
rect 8013 5653 8027 5667
rect 7993 5533 8007 5547
rect 7993 5433 8007 5447
rect 7973 5413 7987 5427
rect 8013 5393 8027 5407
rect 7893 5373 7907 5387
rect 8013 5373 8027 5387
rect 7953 5153 7967 5167
rect 7933 5133 7947 5147
rect 7913 5093 7927 5107
rect 7893 4913 7907 4927
rect 7933 4913 7947 4927
rect 7813 4693 7827 4707
rect 7793 4653 7807 4667
rect 7753 4453 7767 4467
rect 7733 4433 7747 4447
rect 7773 4433 7787 4447
rect 7773 4393 7787 4407
rect 7813 4393 7827 4407
rect 7713 4313 7727 4327
rect 7693 4273 7707 4287
rect 7753 4273 7767 4287
rect 7693 4233 7707 4247
rect 7693 4193 7707 4207
rect 7733 4193 7747 4207
rect 7713 4173 7727 4187
rect 7693 3993 7707 4007
rect 7673 3593 7687 3607
rect 7733 4073 7747 4087
rect 7733 3953 7747 3967
rect 7813 4193 7827 4207
rect 7793 3933 7807 3947
rect 7773 3913 7787 3927
rect 7753 3753 7767 3767
rect 7733 3693 7747 3707
rect 7933 4713 7947 4727
rect 7973 4713 7987 4727
rect 7873 4693 7887 4707
rect 7913 4693 7927 4707
rect 7953 4673 7967 4687
rect 7893 4613 7907 4627
rect 7853 4413 7867 4427
rect 7933 4513 7947 4527
rect 7973 4513 7987 4527
rect 7953 4453 7967 4467
rect 7973 4453 7987 4467
rect 7973 4433 7987 4447
rect 7953 4413 7967 4427
rect 8173 6073 8187 6087
rect 8133 6033 8147 6047
rect 8133 5933 8147 5947
rect 8173 5913 8187 5927
rect 8073 5713 8087 5727
rect 8153 5693 8167 5707
rect 8073 5673 8087 5687
rect 8093 5673 8107 5687
rect 8113 5593 8127 5607
rect 8093 5413 8107 5427
rect 8053 5373 8067 5387
rect 8053 5153 8067 5167
rect 8053 4913 8067 4927
rect 8053 4713 8067 4727
rect 8013 4693 8027 4707
rect 8033 4693 8047 4707
rect 8033 4673 8047 4687
rect 8013 4633 8027 4647
rect 8013 4473 8027 4487
rect 8013 4433 8027 4447
rect 8033 4353 8047 4367
rect 7993 4313 8007 4327
rect 7933 4193 7947 4207
rect 7973 4193 7987 4207
rect 7893 4153 7907 4167
rect 7953 4153 7967 4167
rect 7873 4033 7887 4047
rect 7833 3993 7847 4007
rect 7853 3973 7867 3987
rect 7833 3953 7847 3967
rect 7893 3993 7907 4007
rect 7953 3993 7967 4007
rect 7913 3973 7927 3987
rect 7833 3893 7847 3907
rect 7733 3673 7747 3687
rect 7773 3673 7787 3687
rect 7813 3673 7827 3687
rect 7753 3653 7767 3667
rect 7713 3613 7727 3627
rect 7713 3593 7727 3607
rect 7733 3593 7747 3607
rect 7693 3393 7707 3407
rect 7693 3373 7707 3387
rect 7693 3353 7707 3367
rect 7653 3253 7667 3267
rect 7673 3233 7687 3247
rect 7733 3553 7747 3567
rect 7733 3533 7747 3547
rect 7913 3773 7927 3787
rect 7853 3733 7867 3747
rect 7773 3513 7787 3527
rect 7833 3513 7847 3527
rect 7753 3493 7767 3507
rect 7773 3393 7787 3407
rect 7653 3053 7667 3067
rect 7713 3053 7727 3067
rect 7633 2853 7647 2867
rect 7493 2753 7507 2767
rect 7553 2753 7567 2767
rect 7593 2753 7607 2767
rect 7513 2513 7527 2527
rect 7473 2493 7487 2507
rect 7473 2273 7487 2287
rect 7353 2073 7367 2087
rect 7393 2073 7407 2087
rect 7453 2073 7467 2087
rect 7333 1873 7347 1887
rect 7133 1853 7147 1867
rect 7113 1773 7127 1787
rect 7073 1753 7087 1767
rect 7153 1673 7167 1687
rect 7153 1613 7167 1627
rect 7153 1533 7167 1547
rect 7053 1393 7067 1407
rect 7053 1333 7067 1347
rect 7293 1773 7307 1787
rect 7273 1673 7287 1687
rect 7193 1613 7207 1627
rect 7253 1593 7267 1607
rect 7233 1553 7247 1567
rect 7273 1553 7287 1567
rect 7433 2053 7447 2067
rect 7453 2033 7467 2047
rect 7553 1813 7567 1827
rect 7373 1753 7387 1767
rect 7393 1753 7407 1767
rect 7753 3253 7767 3267
rect 7753 3013 7767 3027
rect 7733 2753 7747 2767
rect 7733 2733 7747 2747
rect 7693 2633 7707 2647
rect 7633 2513 7647 2527
rect 7653 2513 7667 2527
rect 7613 2493 7627 2507
rect 7713 2353 7727 2367
rect 7713 2293 7727 2307
rect 7593 2253 7607 2267
rect 7653 2253 7667 2267
rect 7673 2193 7687 2207
rect 7613 2153 7627 2167
rect 7613 2093 7627 2107
rect 7593 2053 7607 2067
rect 7573 1773 7587 1787
rect 7553 1753 7567 1767
rect 7413 1733 7427 1747
rect 7473 1613 7487 1627
rect 7453 1593 7467 1607
rect 7493 1593 7507 1607
rect 7573 1593 7587 1607
rect 7493 1393 7507 1407
rect 7353 1353 7367 1367
rect 7113 1313 7127 1327
rect 7173 1313 7187 1327
rect 7313 1313 7327 1327
rect 7553 1373 7567 1387
rect 7553 1333 7567 1347
rect 7073 1253 7087 1267
rect 7093 1253 7107 1267
rect 7373 1233 7387 1247
rect 7333 1213 7347 1227
rect 7113 1193 7127 1207
rect 7053 1153 7067 1167
rect 7033 1073 7047 1087
rect 6993 853 7007 867
rect 7033 853 7047 867
rect 6953 773 6967 787
rect 6833 753 6847 767
rect 6653 353 6667 367
rect 6993 673 7007 687
rect 7133 1133 7147 1147
rect 7173 1133 7187 1147
rect 7113 893 7127 907
rect 7053 653 7067 667
rect 7033 633 7047 647
rect 6973 393 6987 407
rect 6753 373 6767 387
rect 7153 1053 7167 1067
rect 7133 853 7147 867
rect 7153 833 7167 847
rect 7173 813 7187 827
rect 7153 793 7167 807
rect 7213 833 7227 847
rect 7253 753 7267 767
rect 7193 733 7207 747
rect 7413 1093 7427 1107
rect 7453 1093 7467 1107
rect 7353 1073 7367 1087
rect 7393 1073 7407 1087
rect 7353 993 7367 1007
rect 7373 933 7387 947
rect 7353 913 7367 927
rect 7353 853 7367 867
rect 7393 873 7407 887
rect 7373 833 7387 847
rect 7453 1033 7467 1047
rect 7433 913 7447 927
rect 7533 913 7547 927
rect 7453 853 7467 867
rect 7493 853 7507 867
rect 7433 833 7447 847
rect 7473 833 7487 847
rect 7413 813 7427 827
rect 7393 773 7407 787
rect 7253 693 7267 707
rect 7313 693 7327 707
rect 7333 693 7347 707
rect 7273 653 7287 667
rect 7233 633 7247 647
rect 7113 573 7127 587
rect 7473 653 7487 667
rect 7493 653 7507 667
rect 7553 893 7567 907
rect 7753 2153 7767 2167
rect 7653 1813 7667 1827
rect 7693 1713 7707 1727
rect 7713 1633 7727 1647
rect 7633 1593 7647 1607
rect 7693 1573 7707 1587
rect 7673 1553 7687 1567
rect 7813 3253 7827 3267
rect 7813 3213 7827 3227
rect 7813 3013 7827 3027
rect 7793 2993 7807 3007
rect 7793 2973 7807 2987
rect 7833 2973 7847 2987
rect 7833 2633 7847 2647
rect 7913 3553 7927 3567
rect 7993 4073 8007 4087
rect 8033 3993 8047 4007
rect 7993 3873 8007 3887
rect 8033 3753 8047 3767
rect 8073 4693 8087 4707
rect 8153 5513 8167 5527
rect 8153 5413 8167 5427
rect 8213 6133 8227 6147
rect 8213 6073 8227 6087
rect 8113 5213 8127 5227
rect 8333 7193 8347 7207
rect 8413 7193 8427 7207
rect 8313 7173 8327 7187
rect 8293 6593 8307 6607
rect 8373 7093 8387 7107
rect 8393 7073 8407 7087
rect 8413 7013 8427 7027
rect 8373 6813 8387 6827
rect 8473 6853 8487 6867
rect 8433 6773 8447 6787
rect 8673 9453 8687 9467
rect 8633 9033 8647 9047
rect 8553 8993 8567 9007
rect 8593 8993 8607 9007
rect 8573 8973 8587 8987
rect 8613 8973 8627 8987
rect 8553 8933 8567 8947
rect 8593 8853 8607 8867
rect 8633 8853 8647 8867
rect 8653 8853 8667 8867
rect 8573 8813 8587 8827
rect 8553 8753 8567 8767
rect 8533 8533 8547 8547
rect 8513 8493 8527 8507
rect 8613 8773 8627 8787
rect 8593 8753 8607 8767
rect 8593 8693 8607 8707
rect 8593 8653 8607 8667
rect 8653 8653 8667 8667
rect 8653 8533 8667 8547
rect 8633 8393 8647 8407
rect 8593 8353 8607 8367
rect 8553 8293 8567 8307
rect 8573 8293 8587 8307
rect 8573 8233 8587 8247
rect 8533 7993 8547 8007
rect 8893 10493 8907 10507
rect 8853 10433 8867 10447
rect 8913 10373 8927 10387
rect 8873 10253 8887 10267
rect 8853 10233 8867 10247
rect 8813 10013 8827 10027
rect 8773 9953 8787 9967
rect 8753 9673 8767 9687
rect 8833 9933 8847 9947
rect 8793 9773 8807 9787
rect 8813 9733 8827 9747
rect 8893 10233 8907 10247
rect 8893 10033 8907 10047
rect 8873 9653 8887 9667
rect 8813 9493 8827 9507
rect 8833 9453 8847 9467
rect 8773 9433 8787 9447
rect 8793 9433 8807 9447
rect 8793 9413 8807 9427
rect 8793 9393 8807 9407
rect 8833 9333 8847 9347
rect 8833 9273 8847 9287
rect 8773 9253 8787 9267
rect 8773 9153 8787 9167
rect 8813 9153 8827 9167
rect 8733 8973 8747 8987
rect 8753 8793 8767 8807
rect 8693 8733 8707 8747
rect 8713 8353 8727 8367
rect 8693 8293 8707 8307
rect 8633 8173 8647 8187
rect 8593 8073 8607 8087
rect 8573 7813 8587 7827
rect 8613 7813 8627 7827
rect 8573 7793 8587 7807
rect 8513 7573 8527 7587
rect 8513 7513 8527 7527
rect 8533 7233 8547 7247
rect 8513 7153 8527 7167
rect 8513 7093 8527 7107
rect 8553 7213 8567 7227
rect 8893 9393 8907 9407
rect 9013 10673 9027 10687
rect 8953 10433 8967 10447
rect 9173 10873 9187 10887
rect 9233 10853 9247 10867
rect 9153 10693 9167 10707
rect 9133 10453 9147 10467
rect 9113 10433 9127 10447
rect 9133 10413 9147 10427
rect 9093 10393 9107 10407
rect 9253 10693 9267 10707
rect 9313 10673 9327 10687
rect 9433 10913 9447 10927
rect 9393 10893 9407 10907
rect 9413 10893 9427 10907
rect 9613 10893 9627 10907
rect 9353 10853 9367 10867
rect 9393 10753 9407 10767
rect 9653 10873 9667 10887
rect 9413 10693 9427 10707
rect 9413 10673 9427 10687
rect 9213 10433 9227 10447
rect 9173 10393 9187 10407
rect 9113 10373 9127 10387
rect 9153 10373 9167 10387
rect 9093 10253 9107 10267
rect 9273 10233 9287 10247
rect 9113 10193 9127 10207
rect 9013 10133 9027 10147
rect 9093 10133 9107 10147
rect 8993 9953 9007 9967
rect 9033 9953 9047 9967
rect 8933 9933 8947 9947
rect 8973 9733 8987 9747
rect 8933 9513 8947 9527
rect 9053 9933 9067 9947
rect 9093 9933 9107 9947
rect 9213 10193 9227 10207
rect 9033 9913 9047 9927
rect 9073 9913 9087 9927
rect 9153 9913 9167 9927
rect 9013 9833 9027 9847
rect 8993 9473 9007 9487
rect 8933 9433 8947 9447
rect 8913 9333 8927 9347
rect 8813 8873 8827 8887
rect 8793 8793 8807 8807
rect 8873 8993 8887 9007
rect 8913 8973 8927 8987
rect 8893 8933 8907 8947
rect 8853 8793 8867 8807
rect 8813 8773 8827 8787
rect 8893 8773 8907 8787
rect 8893 8693 8907 8707
rect 8773 8533 8787 8547
rect 8853 8513 8867 8527
rect 8873 8493 8887 8507
rect 8833 8373 8847 8387
rect 8753 8233 8767 8247
rect 8793 8073 8807 8087
rect 8733 8033 8747 8047
rect 8753 7973 8767 7987
rect 8653 7793 8667 7807
rect 8733 7793 8747 7807
rect 8673 7653 8687 7667
rect 8713 7553 8727 7567
rect 8653 7513 8667 7527
rect 8693 7473 8707 7487
rect 8633 7393 8647 7407
rect 8693 7353 8707 7367
rect 8633 7233 8647 7247
rect 8613 7213 8627 7227
rect 8613 7093 8627 7107
rect 8593 7073 8607 7087
rect 8633 7053 8647 7067
rect 8673 7033 8687 7047
rect 8553 6833 8567 6847
rect 8573 6833 8587 6847
rect 8533 6813 8547 6827
rect 8453 6593 8467 6607
rect 8493 6593 8507 6607
rect 8473 6553 8487 6567
rect 8513 6453 8527 6467
rect 8413 6393 8427 6407
rect 8453 6393 8467 6407
rect 8373 6353 8387 6367
rect 8433 6353 8447 6367
rect 8413 6333 8427 6347
rect 8333 6113 8347 6127
rect 8373 6113 8387 6127
rect 8293 6053 8307 6067
rect 8313 6053 8327 6067
rect 8273 6013 8287 6027
rect 8273 5933 8287 5947
rect 8273 5453 8287 5467
rect 8293 5453 8307 5467
rect 8213 5173 8227 5187
rect 8153 5113 8167 5127
rect 8193 5073 8207 5087
rect 8273 5073 8287 5087
rect 8233 5053 8247 5067
rect 8173 4953 8187 4967
rect 8113 4853 8127 4867
rect 8113 4693 8127 4707
rect 8213 4693 8227 4707
rect 8193 4673 8207 4687
rect 8233 4673 8247 4687
rect 8153 4653 8167 4667
rect 8253 4633 8267 4647
rect 8273 4633 8287 4647
rect 8213 4513 8227 4527
rect 8153 4473 8167 4487
rect 8193 4473 8207 4487
rect 8173 4433 8187 4447
rect 8233 4453 8247 4467
rect 8153 4413 8167 4427
rect 8173 4393 8187 4407
rect 8133 4373 8147 4387
rect 8133 4193 8147 4207
rect 8113 4153 8127 4167
rect 8133 4013 8147 4027
rect 8153 4013 8167 4027
rect 8073 3993 8087 4007
rect 8093 3993 8107 4007
rect 8073 3973 8087 3987
rect 8113 3973 8127 3987
rect 8093 3953 8107 3967
rect 8073 3853 8087 3867
rect 8073 3753 8087 3767
rect 8053 3733 8067 3747
rect 8033 3713 8047 3727
rect 7993 3693 8007 3707
rect 8013 3693 8027 3707
rect 8053 3653 8067 3667
rect 7933 3513 7947 3527
rect 7973 3513 7987 3527
rect 7973 3493 7987 3507
rect 7933 3473 7947 3487
rect 7993 3473 8007 3487
rect 7973 3293 7987 3307
rect 7913 3213 7927 3227
rect 7873 3193 7887 3207
rect 7913 3093 7927 3107
rect 7873 3033 7887 3047
rect 7873 2733 7887 2747
rect 7893 2533 7907 2547
rect 7853 2293 7867 2307
rect 7813 2253 7827 2267
rect 7793 2233 7807 2247
rect 7833 2233 7847 2247
rect 7853 2213 7867 2227
rect 7893 2193 7907 2207
rect 7953 3273 7967 3287
rect 7953 3213 7967 3227
rect 7953 3033 7967 3047
rect 7953 2633 7967 2647
rect 7953 2593 7967 2607
rect 7993 3073 8007 3087
rect 8013 3053 8027 3067
rect 8033 3033 8047 3047
rect 8053 3033 8067 3047
rect 8113 3733 8127 3747
rect 8093 3713 8107 3727
rect 8113 3673 8127 3687
rect 8093 3613 8107 3627
rect 8193 4313 8207 4327
rect 8233 4293 8247 4307
rect 8213 4173 8227 4187
rect 8253 3953 8267 3967
rect 8433 6173 8447 6187
rect 8393 6033 8407 6047
rect 8393 6013 8407 6027
rect 8353 5953 8367 5967
rect 8413 5893 8427 5907
rect 8433 5893 8447 5907
rect 8373 5873 8387 5887
rect 8353 5713 8367 5727
rect 8433 5713 8447 5727
rect 8433 5673 8447 5687
rect 8373 5593 8387 5607
rect 8373 5453 8387 5467
rect 8393 5413 8407 5427
rect 8333 5313 8347 5327
rect 8313 4793 8327 4807
rect 8313 4593 8327 4607
rect 8313 4253 8327 4267
rect 8313 4193 8327 4207
rect 8373 5233 8387 5247
rect 8353 5033 8367 5047
rect 8533 6333 8547 6347
rect 8533 6113 8547 6127
rect 8473 5913 8487 5927
rect 8493 5773 8507 5787
rect 8493 5633 8507 5647
rect 8493 5513 8507 5527
rect 8473 5433 8487 5447
rect 8453 5273 8467 5287
rect 8433 5153 8447 5167
rect 8453 5133 8467 5147
rect 8413 5093 8427 5107
rect 8393 5073 8407 5087
rect 8393 4973 8407 4987
rect 8413 4953 8427 4967
rect 8353 4213 8367 4227
rect 8413 4653 8427 4667
rect 8453 4653 8467 4667
rect 8433 4633 8447 4647
rect 8513 5153 8527 5167
rect 8493 5133 8507 5147
rect 8473 4613 8487 4627
rect 8473 4513 8487 4527
rect 8433 4493 8447 4507
rect 8453 4473 8467 4487
rect 8413 4353 8427 4367
rect 8433 4193 8447 4207
rect 8513 4933 8527 4947
rect 8573 6413 8587 6427
rect 8833 7893 8847 7907
rect 8793 7833 8807 7847
rect 8773 7813 8787 7827
rect 8793 7793 8807 7807
rect 8853 7853 8867 7867
rect 8773 7053 8787 7067
rect 8753 6953 8767 6967
rect 8753 6913 8767 6927
rect 8673 6833 8687 6847
rect 8673 6733 8687 6747
rect 8713 6733 8727 6747
rect 8693 6593 8707 6607
rect 8633 6413 8647 6427
rect 8733 6593 8747 6607
rect 8753 6593 8767 6607
rect 8713 6553 8727 6567
rect 8653 6373 8667 6387
rect 8693 6373 8707 6387
rect 8613 6273 8627 6287
rect 8693 6193 8707 6207
rect 8613 6173 8627 6187
rect 8673 6113 8687 6127
rect 8653 6093 8667 6107
rect 8693 6073 8707 6087
rect 8633 6033 8647 6047
rect 8593 6013 8607 6027
rect 8653 5933 8667 5947
rect 8613 5913 8627 5927
rect 8633 5893 8647 5907
rect 8573 5553 8587 5567
rect 8713 5813 8727 5827
rect 8733 5693 8747 5707
rect 8633 5533 8647 5547
rect 8553 5353 8567 5367
rect 8553 5153 8567 5167
rect 8753 5653 8767 5667
rect 8733 5533 8747 5547
rect 8693 5513 8707 5527
rect 8653 5433 8667 5447
rect 8713 5173 8727 5187
rect 8673 5133 8687 5147
rect 8593 5093 8607 5107
rect 8573 5033 8587 5047
rect 8533 4673 8547 4687
rect 8513 4653 8527 4667
rect 8513 4433 8527 4447
rect 8653 5013 8667 5027
rect 8693 5113 8707 5127
rect 8673 4953 8687 4967
rect 8633 4933 8647 4947
rect 8673 4933 8687 4947
rect 8753 4933 8767 4947
rect 8593 4753 8607 4767
rect 8573 4493 8587 4507
rect 8553 4273 8567 4287
rect 8573 4273 8587 4287
rect 8393 4153 8407 4167
rect 8413 4153 8427 4167
rect 8493 4153 8507 4167
rect 8333 4093 8347 4107
rect 8333 4013 8347 4027
rect 8253 3693 8267 3707
rect 8293 3693 8307 3707
rect 8273 3673 8287 3687
rect 8253 3633 8267 3647
rect 8213 3553 8227 3567
rect 8213 3493 8227 3507
rect 8233 3473 8247 3487
rect 8193 3393 8207 3407
rect 8193 3373 8207 3387
rect 8093 3293 8107 3307
rect 8093 3233 8107 3247
rect 8133 3233 8147 3247
rect 8073 2773 8087 2787
rect 8013 2733 8027 2747
rect 8013 2713 8027 2727
rect 7973 2573 7987 2587
rect 7973 2553 7987 2567
rect 7953 2533 7967 2547
rect 7993 2533 8007 2547
rect 7933 2173 7947 2187
rect 7933 2133 7947 2147
rect 8073 2613 8087 2627
rect 8153 3213 8167 3227
rect 8173 3193 8187 3207
rect 8113 3153 8127 3167
rect 8113 2773 8127 2787
rect 8093 2333 8107 2347
rect 8053 2253 8067 2267
rect 8033 2113 8047 2127
rect 8033 2073 8047 2087
rect 7893 1833 7907 1847
rect 8013 1853 8027 1867
rect 7993 1813 8007 1827
rect 7913 1793 7927 1807
rect 7873 1773 7887 1787
rect 7833 1753 7847 1767
rect 7773 1373 7787 1387
rect 7793 1333 7807 1347
rect 7833 1333 7847 1347
rect 7813 1313 7827 1327
rect 7593 1133 7607 1147
rect 7633 1133 7647 1147
rect 7653 1133 7667 1147
rect 7753 1133 7767 1147
rect 7773 1133 7787 1147
rect 7753 993 7767 1007
rect 7913 1613 7927 1627
rect 7893 1593 7907 1607
rect 7953 1553 7967 1567
rect 7893 1373 7907 1387
rect 7573 833 7587 847
rect 7593 813 7607 827
rect 7713 753 7727 767
rect 7733 693 7747 707
rect 7513 633 7527 647
rect 7533 633 7547 647
rect 7353 373 7367 387
rect 6733 333 6747 347
rect 6853 333 6867 347
rect 6893 333 6907 347
rect 6993 333 7007 347
rect 7113 333 7127 347
rect 6513 213 6527 227
rect 6493 173 6507 187
rect 6733 253 6747 267
rect 6593 193 6607 207
rect 6753 153 6767 167
rect 6553 113 6567 127
rect 6713 113 6727 127
rect 6773 133 6787 147
rect 6993 273 7007 287
rect 7153 293 7167 307
rect 7133 153 7147 167
rect 7193 153 7207 167
rect 6973 133 6987 147
rect 7413 313 7427 327
rect 7713 613 7727 627
rect 7933 1333 7947 1347
rect 7913 1073 7927 1087
rect 7993 1073 8007 1087
rect 7893 913 7907 927
rect 7933 913 7947 927
rect 7893 713 7907 727
rect 7873 573 7887 587
rect 7633 393 7647 407
rect 7873 373 7887 387
rect 7913 373 7927 387
rect 7673 333 7687 347
rect 7973 913 7987 927
rect 7993 813 8007 827
rect 8093 2193 8107 2207
rect 8093 2053 8107 2067
rect 8293 3153 8307 3167
rect 8273 3053 8287 3067
rect 8333 3713 8347 3727
rect 8313 3053 8327 3067
rect 8253 3033 8267 3047
rect 8293 3033 8307 3047
rect 8253 2853 8267 2867
rect 8193 2833 8207 2847
rect 8153 2693 8167 2707
rect 8293 2733 8307 2747
rect 8273 2693 8287 2707
rect 8273 2613 8287 2627
rect 8233 2593 8247 2607
rect 8253 2593 8267 2607
rect 8213 2553 8227 2567
rect 8233 2533 8247 2547
rect 8173 2513 8187 2527
rect 8233 2513 8247 2527
rect 8213 2473 8227 2487
rect 8213 2173 8227 2187
rect 8153 2113 8167 2127
rect 8133 2073 8147 2087
rect 8193 2073 8207 2087
rect 8133 2053 8147 2067
rect 8173 2053 8187 2067
rect 8213 2053 8227 2067
rect 8113 1853 8127 1867
rect 8093 1813 8107 1827
rect 8133 1813 8147 1827
rect 8113 1793 8127 1807
rect 8153 1793 8167 1807
rect 8073 1753 8087 1767
rect 8113 1593 8127 1607
rect 8173 1593 8187 1607
rect 8193 1593 8207 1607
rect 8113 1573 8127 1587
rect 8153 1573 8167 1587
rect 8133 1553 8147 1567
rect 8113 1533 8127 1547
rect 8313 2533 8327 2547
rect 8253 2273 8267 2287
rect 8413 4013 8427 4027
rect 8553 4013 8567 4027
rect 8393 3913 8407 3927
rect 8373 3693 8387 3707
rect 8453 3993 8467 4007
rect 8573 3993 8587 4007
rect 8573 3953 8587 3967
rect 8513 3853 8527 3867
rect 8513 3793 8527 3807
rect 8453 3633 8467 3647
rect 8533 3713 8547 3727
rect 8513 3693 8527 3707
rect 8553 3693 8567 3707
rect 8533 3673 8547 3687
rect 8553 3633 8567 3647
rect 8453 3613 8467 3627
rect 8493 3613 8507 3627
rect 8433 3573 8447 3587
rect 8413 3533 8427 3547
rect 8353 3493 8367 3507
rect 8453 3513 8467 3527
rect 8473 3473 8487 3487
rect 8433 3353 8447 3367
rect 8393 3213 8407 3227
rect 8373 3173 8387 3187
rect 8353 2253 8367 2267
rect 8253 2113 8267 2127
rect 8253 1793 8267 1807
rect 8353 2073 8367 2087
rect 8393 2133 8407 2147
rect 8453 3193 8467 3207
rect 8553 3393 8567 3407
rect 8633 4693 8647 4707
rect 8653 4673 8667 4687
rect 8733 4613 8747 4627
rect 8693 4593 8707 4607
rect 8613 4493 8627 4507
rect 8673 4493 8687 4507
rect 8693 4473 8707 4487
rect 8813 7693 8827 7707
rect 8953 9333 8967 9347
rect 8933 8493 8947 8507
rect 8913 8313 8927 8327
rect 8933 8253 8947 8267
rect 8933 7833 8947 7847
rect 8893 7813 8907 7827
rect 8913 7613 8927 7627
rect 8873 7473 8887 7487
rect 8873 7413 8887 7427
rect 8853 7333 8867 7347
rect 8853 7073 8867 7087
rect 9253 9993 9267 10007
rect 9233 9953 9247 9967
rect 9233 9773 9247 9787
rect 9193 9733 9207 9747
rect 9233 9733 9247 9747
rect 9213 9713 9227 9727
rect 9153 9653 9167 9667
rect 9173 9613 9187 9627
rect 9093 9473 9107 9487
rect 9053 9453 9067 9467
rect 9133 9273 9147 9287
rect 9073 9253 9087 9267
rect 9053 9233 9067 9247
rect 9013 9173 9027 9187
rect 9113 9233 9127 9247
rect 9073 8993 9087 9007
rect 9153 8993 9167 9007
rect 9093 8973 9107 8987
rect 8973 8893 8987 8907
rect 9133 8813 9147 8827
rect 9093 8793 9107 8807
rect 9073 8773 9087 8787
rect 9113 8773 9127 8787
rect 9333 10453 9347 10467
rect 9373 10453 9387 10467
rect 9413 10453 9427 10467
rect 9453 10453 9467 10467
rect 9473 10453 9487 10467
rect 9353 10433 9367 10447
rect 9393 10433 9407 10447
rect 9333 10373 9347 10387
rect 9313 10033 9327 10047
rect 9393 10193 9407 10207
rect 9413 10153 9427 10167
rect 9393 9973 9407 9987
rect 9313 9953 9327 9967
rect 9353 9953 9367 9967
rect 9373 9953 9387 9967
rect 9293 9933 9307 9947
rect 9293 9773 9307 9787
rect 9273 9713 9287 9727
rect 9313 9513 9327 9527
rect 9333 9513 9347 9527
rect 9353 9473 9367 9487
rect 9273 9453 9287 9467
rect 9333 9453 9347 9467
rect 9293 9433 9307 9447
rect 9373 9433 9387 9447
rect 9333 9313 9347 9327
rect 9293 9273 9307 9287
rect 9333 9273 9347 9287
rect 9233 9253 9247 9267
rect 9273 9253 9287 9267
rect 9193 8993 9207 9007
rect 9213 8793 9227 8807
rect 9193 8773 9207 8787
rect 9173 8753 9187 8767
rect 9033 8733 9047 8747
rect 9073 8733 9087 8747
rect 8993 8033 9007 8047
rect 9013 8013 9027 8027
rect 9013 7853 9027 7867
rect 9013 7833 9027 7847
rect 8973 7673 8987 7687
rect 8953 7613 8967 7627
rect 8933 7573 8947 7587
rect 8953 7553 8967 7567
rect 9013 7553 9027 7567
rect 8993 7493 9007 7507
rect 8993 7473 9007 7487
rect 8933 7433 8947 7447
rect 8913 7053 8927 7067
rect 8873 7033 8887 7047
rect 9013 7373 9027 7387
rect 8993 7313 9007 7327
rect 8933 6873 8947 6887
rect 9013 7033 9027 7047
rect 8993 6853 9007 6867
rect 8913 6713 8927 6727
rect 8953 6593 8967 6607
rect 8833 6533 8847 6547
rect 8913 6533 8927 6547
rect 8873 6393 8887 6407
rect 8973 6573 8987 6587
rect 8973 6413 8987 6427
rect 8813 6373 8827 6387
rect 8853 6373 8867 6387
rect 8893 6373 8907 6387
rect 8933 6373 8947 6387
rect 8793 6093 8807 6107
rect 8893 6113 8907 6127
rect 8913 6093 8927 6107
rect 8873 6053 8887 6067
rect 8913 6053 8927 6067
rect 8853 6033 8867 6047
rect 8893 6033 8907 6047
rect 8873 6013 8887 6027
rect 8793 5913 8807 5927
rect 8833 5913 8847 5927
rect 8773 4713 8787 4727
rect 8713 4453 8727 4467
rect 8753 4453 8767 4467
rect 8753 4413 8767 4427
rect 8853 5893 8867 5907
rect 8893 5893 8907 5907
rect 8813 5693 8827 5707
rect 8793 4393 8807 4407
rect 8613 4293 8627 4307
rect 8693 4273 8707 4287
rect 8733 4253 8747 4267
rect 8653 4173 8667 4187
rect 8713 4173 8727 4187
rect 8673 4153 8687 4167
rect 8613 4093 8627 4107
rect 8633 4093 8647 4107
rect 8613 4013 8627 4027
rect 8613 3793 8627 3807
rect 8593 3273 8607 3287
rect 8833 5653 8847 5667
rect 8873 5433 8887 5447
rect 8973 6113 8987 6127
rect 8933 6033 8947 6047
rect 8933 5973 8947 5987
rect 8933 5933 8947 5947
rect 8953 5933 8967 5947
rect 8973 5913 8987 5927
rect 8973 5613 8987 5627
rect 8933 5593 8947 5607
rect 9073 8513 9087 8527
rect 9113 8513 9127 8527
rect 9053 8493 9067 8507
rect 9093 8493 9107 8507
rect 9133 8473 9147 8487
rect 9133 8313 9147 8327
rect 9153 8313 9167 8327
rect 9173 8133 9187 8147
rect 9153 8073 9167 8087
rect 9213 8073 9227 8087
rect 9053 8033 9067 8047
rect 9133 7893 9147 7907
rect 9053 7833 9067 7847
rect 9093 7833 9107 7847
rect 9193 8053 9207 8067
rect 9353 9053 9367 9067
rect 9313 8953 9327 8967
rect 9253 8873 9267 8887
rect 9313 8773 9327 8787
rect 9293 8753 9307 8767
rect 9333 8753 9347 8767
rect 9253 8713 9267 8727
rect 9373 8973 9387 8987
rect 9373 8953 9387 8967
rect 9373 8753 9387 8767
rect 9353 8573 9367 8587
rect 9353 8533 9367 8547
rect 9293 8493 9307 8507
rect 9293 8373 9307 8387
rect 9253 8053 9267 8067
rect 9233 8033 9247 8047
rect 9153 7833 9167 7847
rect 9073 7813 9087 7827
rect 9113 7813 9127 7827
rect 9153 7813 9167 7827
rect 9193 7793 9207 7807
rect 9133 7573 9147 7587
rect 9073 7393 9087 7407
rect 9113 7373 9127 7387
rect 9233 7773 9247 7787
rect 9213 7473 9227 7487
rect 9173 7413 9187 7427
rect 9153 7353 9167 7367
rect 9053 7333 9067 7347
rect 9133 7333 9147 7347
rect 9093 7313 9107 7327
rect 9233 7273 9247 7287
rect 9273 8033 9287 8047
rect 9373 8493 9387 8507
rect 9333 8333 9347 8347
rect 9413 9773 9427 9787
rect 9433 9733 9447 9747
rect 9413 9413 9427 9427
rect 9393 8453 9407 8467
rect 9853 11113 9867 11127
rect 9833 10933 9847 10947
rect 9893 10933 9907 10947
rect 9793 10913 9807 10927
rect 9853 10893 9867 10907
rect 9933 10913 9947 10927
rect 10233 11173 10247 11187
rect 10373 11173 10387 11187
rect 10413 11173 10427 11187
rect 10613 11173 10627 11187
rect 10733 11173 10747 11187
rect 10833 11173 10847 11187
rect 10873 11173 10887 11187
rect 11073 11173 11087 11187
rect 10093 11153 10107 11167
rect 10133 11153 10147 11167
rect 10113 11113 10127 11127
rect 9913 10893 9927 10907
rect 9893 10873 9907 10887
rect 9873 10813 9887 10827
rect 9673 10693 9687 10707
rect 10093 10893 10107 10907
rect 10133 10873 10147 10887
rect 10193 10873 10207 10887
rect 9953 10813 9967 10827
rect 10073 10813 10087 10827
rect 9933 10733 9947 10747
rect 10213 10733 10227 10747
rect 9993 10713 10007 10727
rect 9893 10653 9907 10667
rect 9933 10653 9947 10667
rect 9973 10653 9987 10667
rect 9733 10493 9747 10507
rect 9613 10433 9627 10447
rect 9593 10413 9607 10427
rect 9633 10413 9647 10427
rect 9573 10373 9587 10387
rect 9673 10373 9687 10387
rect 9473 10213 9487 10227
rect 9533 10213 9547 10227
rect 9513 10193 9527 10207
rect 9673 10233 9687 10247
rect 9913 10413 9927 10427
rect 9873 10393 9887 10407
rect 9893 10393 9907 10407
rect 9833 10373 9847 10387
rect 9793 10233 9807 10247
rect 9773 10213 9787 10227
rect 9813 10213 9827 10227
rect 9873 10193 9887 10207
rect 9733 10133 9747 10147
rect 9813 10133 9827 10147
rect 9813 9973 9827 9987
rect 9853 9973 9867 9987
rect 9473 9893 9487 9907
rect 9833 9773 9847 9787
rect 9653 9753 9667 9767
rect 9513 9733 9527 9747
rect 9633 9733 9647 9747
rect 9713 9693 9727 9707
rect 9893 9773 9907 9787
rect 9993 10413 10007 10427
rect 9973 10193 9987 10207
rect 9913 9733 9927 9747
rect 10153 10653 10167 10667
rect 10113 10433 10127 10447
rect 10013 10393 10027 10407
rect 10033 10393 10047 10407
rect 10093 10393 10107 10407
rect 10013 10293 10027 10307
rect 10353 11153 10367 11167
rect 10293 11133 10307 11147
rect 10333 10913 10347 10927
rect 10553 10893 10567 10907
rect 10593 10893 10607 10907
rect 10633 10933 10647 10947
rect 10633 10913 10647 10927
rect 10713 10893 10727 10907
rect 10553 10873 10567 10887
rect 10613 10873 10627 10887
rect 10573 10753 10587 10767
rect 10693 10753 10707 10767
rect 10253 10613 10267 10627
rect 10313 10613 10327 10627
rect 10313 10433 10327 10447
rect 10453 10733 10467 10747
rect 10653 10713 10667 10727
rect 10713 10713 10727 10727
rect 10473 10693 10487 10707
rect 10633 10693 10647 10707
rect 10673 10693 10687 10707
rect 10713 10693 10727 10707
rect 10273 10413 10287 10427
rect 10253 10393 10267 10407
rect 10233 10213 10247 10227
rect 10353 10413 10367 10427
rect 10393 10413 10407 10427
rect 10013 10193 10027 10207
rect 10053 10193 10067 10207
rect 10293 10193 10307 10207
rect 10253 10153 10267 10167
rect 10333 10393 10347 10407
rect 10633 10653 10647 10667
rect 10593 10453 10607 10467
rect 10593 10433 10607 10447
rect 10553 10333 10567 10347
rect 10513 10233 10527 10247
rect 10453 10213 10467 10227
rect 10493 10213 10507 10227
rect 10313 10153 10327 10167
rect 10333 10013 10347 10027
rect 10193 9973 10207 9987
rect 10273 9973 10287 9987
rect 10293 9973 10307 9987
rect 9993 9953 10007 9967
rect 10153 9953 10167 9967
rect 9973 9713 9987 9727
rect 10033 9913 10047 9927
rect 10013 9773 10027 9787
rect 9873 9693 9887 9707
rect 9993 9693 10007 9707
rect 9853 9673 9867 9687
rect 9973 9673 9987 9687
rect 9673 9633 9687 9647
rect 9833 9633 9847 9647
rect 9513 9473 9527 9487
rect 9793 9473 9807 9487
rect 9673 9433 9687 9447
rect 9453 9353 9467 9367
rect 9713 9313 9727 9327
rect 9493 9293 9507 9307
rect 9633 9293 9647 9307
rect 9473 9253 9487 9267
rect 9593 9253 9607 9267
rect 9693 9273 9707 9287
rect 9673 9253 9687 9267
rect 9693 9233 9707 9247
rect 9633 9073 9647 9087
rect 9573 8973 9587 8987
rect 9613 8973 9627 8987
rect 9533 8953 9547 8967
rect 9613 8833 9627 8847
rect 9533 8793 9547 8807
rect 9573 8793 9587 8807
rect 9553 8773 9567 8787
rect 9493 8573 9507 8587
rect 9433 8373 9447 8387
rect 9393 8313 9407 8327
rect 9413 8313 9427 8327
rect 9433 8293 9447 8307
rect 9453 8233 9467 8247
rect 9413 8073 9427 8087
rect 9293 7733 9307 7747
rect 9293 7573 9307 7587
rect 9273 7533 9287 7547
rect 9373 7733 9387 7747
rect 9393 7533 9407 7547
rect 9333 7513 9347 7527
rect 9293 7493 9307 7507
rect 9333 7473 9347 7487
rect 9393 7433 9407 7447
rect 9353 7353 9367 7367
rect 9313 7333 9327 7347
rect 9553 8553 9567 8567
rect 9533 8533 9547 8547
rect 9513 8493 9527 8507
rect 9493 8293 9507 8307
rect 9573 8493 9587 8507
rect 9613 8473 9627 8487
rect 9653 8473 9667 8487
rect 9533 8453 9547 8467
rect 9873 9473 9887 9487
rect 9933 9293 9947 9307
rect 9913 9233 9927 9247
rect 9853 9213 9867 9227
rect 9933 9213 9947 9227
rect 9893 9053 9907 9067
rect 9713 8993 9727 9007
rect 9853 8993 9867 9007
rect 9833 8973 9847 8987
rect 9873 8973 9887 8987
rect 9873 8853 9887 8867
rect 9913 8853 9927 8867
rect 9753 8793 9767 8807
rect 9753 8753 9767 8767
rect 9713 8693 9727 8707
rect 9833 8793 9847 8807
rect 9853 8773 9867 8787
rect 9813 8693 9827 8707
rect 9833 8673 9847 8687
rect 9773 8553 9787 8567
rect 9793 8533 9807 8547
rect 9813 8513 9827 8527
rect 9773 8493 9787 8507
rect 9853 8493 9867 8507
rect 9833 8433 9847 8447
rect 9833 8313 9847 8327
rect 9913 8313 9927 8327
rect 9633 8273 9647 8287
rect 9513 8233 9527 8247
rect 9473 8133 9487 8147
rect 9513 8133 9527 8147
rect 9433 8013 9447 8027
rect 9453 8013 9467 8027
rect 9493 8013 9507 8027
rect 9533 7833 9547 7847
rect 9573 7833 9587 7847
rect 9613 7833 9627 7847
rect 9513 7813 9527 7827
rect 9553 7813 9567 7827
rect 9593 7813 9607 7827
rect 9693 8273 9707 8287
rect 9873 8293 9887 8307
rect 9673 8213 9687 8227
rect 9693 8213 9707 8227
rect 9833 8133 9847 8147
rect 9893 8133 9907 8147
rect 9693 8073 9707 8087
rect 9753 8053 9767 8067
rect 9753 8013 9767 8027
rect 9713 7833 9727 7847
rect 9913 8073 9927 8087
rect 9913 8013 9927 8027
rect 9873 7833 9887 7847
rect 9473 7673 9487 7687
rect 9433 7513 9447 7527
rect 9313 7313 9327 7327
rect 9413 7313 9427 7327
rect 9433 7313 9447 7327
rect 9253 7113 9267 7127
rect 9053 7093 9067 7107
rect 9113 7093 9127 7107
rect 9033 6833 9047 6847
rect 9073 7073 9087 7087
rect 9293 7053 9307 7067
rect 9133 7033 9147 7047
rect 9093 7013 9107 7027
rect 9093 6973 9107 6987
rect 9053 6793 9067 6807
rect 9233 6953 9247 6967
rect 9113 6853 9127 6867
rect 9153 6853 9167 6867
rect 9093 6733 9107 6747
rect 9133 6833 9147 6847
rect 9113 6613 9127 6627
rect 9173 6733 9187 6747
rect 9153 6613 9167 6627
rect 9173 6573 9187 6587
rect 9173 6513 9187 6527
rect 9133 6433 9147 6447
rect 9113 6413 9127 6427
rect 9033 6393 9047 6407
rect 9073 6393 9087 6407
rect 9013 5593 9027 5607
rect 8993 5473 9007 5487
rect 8973 5133 8987 5147
rect 8913 5093 8927 5107
rect 8893 4953 8907 4967
rect 8953 5113 8967 5127
rect 8933 5053 8947 5067
rect 8993 5093 9007 5107
rect 8933 4893 8947 4907
rect 8933 4793 8947 4807
rect 8873 4673 8887 4687
rect 8873 4633 8887 4647
rect 8853 4553 8867 4567
rect 8833 4533 8847 4547
rect 8813 4233 8827 4247
rect 8813 4213 8827 4227
rect 8733 4053 8747 4067
rect 8773 4033 8787 4047
rect 8793 3953 8807 3967
rect 8753 3933 8767 3947
rect 8733 3733 8747 3747
rect 8653 3713 8667 3727
rect 8713 3713 8727 3727
rect 8653 3673 8667 3687
rect 8633 3653 8647 3667
rect 8793 3633 8807 3647
rect 8693 3533 8707 3547
rect 8753 3533 8767 3547
rect 8793 3513 8807 3527
rect 8613 3253 8627 3267
rect 8493 3133 8507 3147
rect 8493 3073 8507 3087
rect 8433 3053 8447 3067
rect 8533 3053 8547 3067
rect 8493 2953 8507 2967
rect 8433 2773 8447 2787
rect 8453 2653 8467 2667
rect 8473 2613 8487 2627
rect 8453 2573 8467 2587
rect 8473 2553 8487 2567
rect 8633 3193 8647 3207
rect 8553 2753 8567 2767
rect 8593 2753 8607 2767
rect 8533 2733 8547 2747
rect 8573 2713 8587 2727
rect 8693 3253 8707 3267
rect 8673 3033 8687 3047
rect 8653 2793 8667 2807
rect 8653 2753 8667 2767
rect 8633 2733 8647 2747
rect 8513 2653 8527 2667
rect 8513 2593 8527 2607
rect 8533 2293 8547 2307
rect 8573 2293 8587 2307
rect 8553 2253 8567 2267
rect 8513 2153 8527 2167
rect 8493 2133 8507 2147
rect 8413 2033 8427 2047
rect 8373 1833 8387 1847
rect 8373 1813 8387 1827
rect 8333 1773 8347 1787
rect 8373 1693 8387 1707
rect 8313 1633 8327 1647
rect 8293 1373 8307 1387
rect 8293 1353 8307 1367
rect 8053 1313 8067 1327
rect 8193 1173 8207 1187
rect 8073 1153 8087 1167
rect 8193 1133 8207 1147
rect 8173 1113 8187 1127
rect 8213 1093 8227 1107
rect 8233 1093 8247 1107
rect 8273 1093 8287 1107
rect 8213 1073 8227 1087
rect 8173 1053 8187 1067
rect 8033 953 8047 967
rect 8033 913 8047 927
rect 8033 893 8047 907
rect 7613 253 7627 267
rect 7953 333 7967 347
rect 8013 333 8027 347
rect 7613 233 7627 247
rect 7893 233 7907 247
rect 7613 193 7627 207
rect 7393 173 7407 187
rect 7533 173 7547 187
rect 7693 173 7707 187
rect 7653 133 7667 147
rect 6873 113 6887 127
rect 7173 113 7187 127
rect 7213 113 7227 127
rect 7373 113 7387 127
rect 7413 113 7427 127
rect 7633 113 7647 127
rect 7933 153 7947 167
rect 7993 153 8007 167
rect 7893 133 7907 147
rect 7953 133 7967 147
rect 8073 853 8087 867
rect 8213 853 8227 867
rect 8233 833 8247 847
rect 8193 773 8207 787
rect 8173 693 8187 707
rect 8093 653 8107 667
rect 8153 653 8167 667
rect 8133 613 8147 627
rect 8193 653 8207 667
rect 8113 573 8127 587
rect 8093 553 8107 567
rect 8073 453 8087 467
rect 8033 113 8047 127
rect 6433 13 6447 27
rect 8153 333 8167 347
rect 8233 373 8247 387
rect 8193 293 8207 307
rect 8133 233 8147 247
rect 8273 993 8287 1007
rect 8393 1653 8407 1667
rect 8393 1393 8407 1407
rect 8453 2073 8467 2087
rect 8473 2073 8487 2087
rect 8473 2033 8487 2047
rect 8653 2593 8667 2607
rect 8673 2593 8687 2607
rect 8613 2293 8627 2307
rect 8593 2173 8607 2187
rect 8553 1773 8567 1787
rect 8573 1613 8587 1627
rect 8473 1593 8487 1607
rect 8453 1333 8467 1347
rect 8433 1293 8447 1307
rect 8493 1333 8507 1347
rect 8473 1313 8487 1327
rect 8513 1313 8527 1327
rect 8533 1293 8547 1307
rect 8453 1153 8467 1167
rect 8493 1153 8507 1167
rect 8473 1133 8487 1147
rect 8533 1133 8547 1147
rect 8553 1133 8567 1147
rect 8533 1073 8547 1087
rect 8373 893 8387 907
rect 8493 893 8507 907
rect 8313 853 8327 867
rect 8453 853 8467 867
rect 8393 833 8407 847
rect 8433 833 8447 847
rect 8573 853 8587 867
rect 8773 3193 8787 3207
rect 8793 3193 8807 3207
rect 8713 3033 8727 3047
rect 8753 3033 8767 3047
rect 8733 3013 8747 3027
rect 8853 4153 8867 4167
rect 8853 4033 8867 4047
rect 8853 3893 8867 3907
rect 8853 3853 8867 3867
rect 8833 3633 8847 3647
rect 8973 4653 8987 4667
rect 9153 6093 9167 6107
rect 9213 6373 9227 6387
rect 9113 6053 9127 6067
rect 9133 6053 9147 6067
rect 9173 6053 9187 6067
rect 9113 5953 9127 5967
rect 9113 5913 9127 5927
rect 9153 5913 9167 5927
rect 9093 5873 9107 5887
rect 9133 5873 9147 5887
rect 9073 5853 9087 5867
rect 9053 5833 9067 5847
rect 9053 5433 9067 5447
rect 9113 5513 9127 5527
rect 9073 5413 9087 5427
rect 9053 5213 9067 5227
rect 9033 4633 9047 4647
rect 8993 4553 9007 4567
rect 8953 4513 8967 4527
rect 9013 4473 9027 4487
rect 8893 4453 8907 4467
rect 8933 4453 8947 4467
rect 8973 4413 8987 4427
rect 8893 4373 8907 4387
rect 9033 4453 9047 4467
rect 8973 4193 8987 4207
rect 9013 4193 9027 4207
rect 8893 4173 8907 4187
rect 8913 4173 8927 4187
rect 8893 4153 8907 4167
rect 8873 3813 8887 3827
rect 8913 3973 8927 3987
rect 8993 4133 9007 4147
rect 8973 3953 8987 3967
rect 8933 3893 8947 3907
rect 8933 3793 8947 3807
rect 8913 3693 8927 3707
rect 8973 3673 8987 3687
rect 8893 3573 8907 3587
rect 8953 3573 8967 3587
rect 8933 3553 8947 3567
rect 8853 3513 8867 3527
rect 8893 3513 8907 3527
rect 8833 3233 8847 3247
rect 8813 3053 8827 3067
rect 8813 3033 8827 3047
rect 8753 2753 8767 2767
rect 8733 2733 8747 2747
rect 8733 2473 8747 2487
rect 8753 2353 8767 2367
rect 8693 2133 8707 2147
rect 8673 2113 8687 2127
rect 8613 2093 8627 2107
rect 8653 2093 8667 2107
rect 8653 2073 8667 2087
rect 8633 2053 8647 2067
rect 8813 2613 8827 2627
rect 8773 2313 8787 2327
rect 8773 2273 8787 2287
rect 9173 5633 9187 5647
rect 9213 5633 9227 5647
rect 9153 5613 9167 5627
rect 9213 5613 9227 5627
rect 9193 5593 9207 5607
rect 9153 5573 9167 5587
rect 9133 5213 9147 5227
rect 9153 5153 9167 5167
rect 9193 5153 9207 5167
rect 9133 5133 9147 5147
rect 9173 5113 9187 5127
rect 9133 5073 9147 5087
rect 9133 5053 9147 5067
rect 9113 4913 9127 4927
rect 9153 4893 9167 4907
rect 9193 4753 9207 4767
rect 9253 6873 9267 6887
rect 9413 7113 9427 7127
rect 9353 6953 9367 6967
rect 9333 6873 9347 6887
rect 9373 6893 9387 6907
rect 9413 6873 9427 6887
rect 9453 6813 9467 6827
rect 9393 6773 9407 6787
rect 9433 6753 9447 6767
rect 9373 6573 9387 6587
rect 9333 6533 9347 6547
rect 9333 6413 9347 6427
rect 9253 6113 9267 6127
rect 9253 5893 9267 5907
rect 9233 5593 9247 5607
rect 9213 4733 9227 4747
rect 9093 4653 9107 4667
rect 9133 4653 9147 4667
rect 9153 4633 9167 4647
rect 9213 4553 9227 4567
rect 9233 4513 9247 4527
rect 9193 4453 9207 4467
rect 9173 4433 9187 4447
rect 9153 4233 9167 4247
rect 9173 4213 9187 4227
rect 9113 4193 9127 4207
rect 9053 4153 9067 4167
rect 9093 4153 9107 4167
rect 9153 4173 9167 4187
rect 9193 4193 9207 4207
rect 9173 4153 9187 4167
rect 9153 4133 9167 4147
rect 9133 4113 9147 4127
rect 9073 4053 9087 4067
rect 9053 4033 9067 4047
rect 9013 3993 9027 4007
rect 9073 4013 9087 4027
rect 9093 4013 9107 4027
rect 9073 3993 9087 4007
rect 9013 3953 9027 3967
rect 9033 3913 9047 3927
rect 9013 3653 9027 3667
rect 8993 3513 9007 3527
rect 8993 3453 9007 3467
rect 8973 3433 8987 3447
rect 8893 3233 8907 3247
rect 8913 3213 8927 3227
rect 9013 3213 9027 3227
rect 8933 3193 8947 3207
rect 8993 3193 9007 3207
rect 8973 3073 8987 3087
rect 8873 3053 8887 3067
rect 8853 2653 8867 2667
rect 8833 2473 8847 2487
rect 8793 2253 8807 2267
rect 8813 2093 8827 2107
rect 8753 2073 8767 2087
rect 8693 2053 8707 2067
rect 8653 1813 8667 1827
rect 8713 1813 8727 1827
rect 8693 1793 8707 1807
rect 8613 1773 8627 1787
rect 8633 1633 8647 1647
rect 8613 1613 8627 1627
rect 8633 1593 8647 1607
rect 8693 1573 8707 1587
rect 8653 1553 8667 1567
rect 8733 1773 8747 1787
rect 8713 1553 8727 1567
rect 8693 1293 8707 1307
rect 8853 2073 8867 2087
rect 8893 3033 8907 3047
rect 9013 3033 9027 3047
rect 9053 3853 9067 3867
rect 9073 3773 9087 3787
rect 9053 3493 9067 3507
rect 9093 3553 9107 3567
rect 9073 3253 9087 3267
rect 9153 4033 9167 4047
rect 9413 6393 9427 6407
rect 9393 6153 9407 6167
rect 9353 6113 9367 6127
rect 9393 6073 9407 6087
rect 9373 6053 9387 6067
rect 9293 6033 9307 6047
rect 9313 5933 9327 5947
rect 9333 5933 9347 5947
rect 9353 5913 9367 5927
rect 9293 5633 9307 5647
rect 9293 5493 9307 5507
rect 9333 5473 9347 5487
rect 9313 5453 9327 5467
rect 9533 7573 9547 7587
rect 9613 7573 9627 7587
rect 9773 7633 9787 7647
rect 9673 7573 9687 7587
rect 9633 7553 9647 7567
rect 9573 7333 9587 7347
rect 9553 7313 9567 7327
rect 9593 7273 9607 7287
rect 9633 7273 9647 7287
rect 9573 7113 9587 7127
rect 9853 7793 9867 7807
rect 9833 7573 9847 7587
rect 9793 7553 9807 7567
rect 9853 7533 9867 7547
rect 9813 7373 9827 7387
rect 9833 7353 9847 7367
rect 9993 9233 10007 9247
rect 9973 8953 9987 8967
rect 9993 8793 10007 8807
rect 9953 8673 9967 8687
rect 10153 9773 10167 9787
rect 10053 9753 10067 9767
rect 10233 9953 10247 9967
rect 10293 9933 10307 9947
rect 10253 9913 10267 9927
rect 10173 9733 10187 9747
rect 10133 9713 10147 9727
rect 10053 9673 10067 9687
rect 10173 9653 10187 9667
rect 10133 9533 10147 9547
rect 10073 9473 10087 9487
rect 10093 9453 10107 9467
rect 10373 9973 10387 9987
rect 10493 9973 10507 9987
rect 10333 9513 10347 9527
rect 10053 9433 10067 9447
rect 10093 9433 10107 9447
rect 10173 9433 10187 9447
rect 10033 9413 10047 9427
rect 10073 9253 10087 9267
rect 10193 9413 10207 9427
rect 10153 9273 10167 9287
rect 10213 9293 10227 9307
rect 10173 9253 10187 9267
rect 10153 9053 10167 9067
rect 10193 9013 10207 9027
rect 10073 8973 10087 8987
rect 10133 8973 10147 8987
rect 10173 8953 10187 8967
rect 10113 8833 10127 8847
rect 10033 8793 10047 8807
rect 10073 8793 10087 8807
rect 10313 9453 10327 9467
rect 10353 9433 10367 9447
rect 10433 9953 10447 9967
rect 10533 9953 10547 9967
rect 10513 9933 10527 9947
rect 10473 9753 10487 9767
rect 10413 9733 10427 9747
rect 10453 9733 10467 9747
rect 10493 9733 10507 9747
rect 10453 9613 10467 9627
rect 10613 10413 10627 10427
rect 10933 11153 10947 11167
rect 11053 11153 11067 11167
rect 10813 11113 10827 11127
rect 10793 10933 10807 10947
rect 10893 10933 10907 10947
rect 10813 10893 10827 10907
rect 10753 10873 10767 10887
rect 11093 11133 11107 11147
rect 11193 11133 11207 11147
rect 11093 11113 11107 11127
rect 11033 10913 11047 10927
rect 11073 10913 11087 10927
rect 10933 10753 10947 10767
rect 10753 10693 10767 10707
rect 10873 10693 10887 10707
rect 10913 10693 10927 10707
rect 10813 10673 10827 10687
rect 10733 10433 10747 10447
rect 10833 10413 10847 10427
rect 10753 10333 10767 10347
rect 10733 10253 10747 10267
rect 10673 10213 10687 10227
rect 10773 10173 10787 10187
rect 10753 9993 10767 10007
rect 10813 9993 10827 10007
rect 10813 9933 10827 9947
rect 10773 9913 10787 9927
rect 10913 10453 10927 10467
rect 10653 9733 10667 9747
rect 10673 9733 10687 9747
rect 10613 9533 10627 9547
rect 10513 9473 10527 9487
rect 10533 9453 10547 9467
rect 10593 9453 10607 9467
rect 10633 9473 10647 9487
rect 10453 9273 10467 9287
rect 10513 9273 10527 9287
rect 10613 9273 10627 9287
rect 10713 9733 10727 9747
rect 10693 9533 10707 9547
rect 10693 9493 10707 9507
rect 10353 9253 10367 9267
rect 10373 9253 10387 9267
rect 10413 9253 10427 9267
rect 10313 9053 10327 9067
rect 10393 9233 10407 9247
rect 10353 9013 10367 9027
rect 10393 8993 10407 9007
rect 10373 8973 10387 8987
rect 10293 8873 10307 8887
rect 10313 8873 10327 8887
rect 10273 8793 10287 8807
rect 10053 8773 10067 8787
rect 10013 8733 10027 8747
rect 10193 8773 10207 8787
rect 10113 8753 10127 8767
rect 10353 8813 10367 8827
rect 10633 9233 10647 9247
rect 10693 9233 10707 9247
rect 10613 8993 10627 9007
rect 10553 8953 10567 8967
rect 10593 8953 10607 8967
rect 10053 8573 10067 8587
rect 10033 8533 10047 8547
rect 10253 8533 10267 8547
rect 9993 8513 10007 8527
rect 10013 8493 10027 8507
rect 10053 8493 10067 8507
rect 10033 8453 10047 8467
rect 10073 8453 10087 8467
rect 9993 8053 10007 8067
rect 9953 8033 9967 8047
rect 10053 8333 10067 8347
rect 10073 8313 10087 8327
rect 10113 8313 10127 8327
rect 10053 8293 10067 8307
rect 10093 8293 10107 8307
rect 10133 8293 10147 8307
rect 10293 8513 10307 8527
rect 10273 8493 10287 8507
rect 10313 8493 10327 8507
rect 10393 8513 10407 8527
rect 10353 8493 10367 8507
rect 10333 8473 10347 8487
rect 10373 8473 10387 8487
rect 10373 8353 10387 8367
rect 10293 8313 10307 8327
rect 10333 8293 10347 8307
rect 10353 8273 10367 8287
rect 10253 8253 10267 8267
rect 10153 8053 10167 8067
rect 10253 8053 10267 8067
rect 10033 8033 10047 8047
rect 10013 8013 10027 8027
rect 10133 7893 10147 7907
rect 10093 7853 10107 7867
rect 9973 7833 9987 7847
rect 10053 7833 10067 7847
rect 10073 7813 10087 7827
rect 10213 8033 10227 8047
rect 10573 8793 10587 8807
rect 10573 8773 10587 8787
rect 10693 8973 10707 8987
rect 10653 8793 10667 8807
rect 10533 8753 10547 8767
rect 10633 8753 10647 8767
rect 10533 8533 10547 8547
rect 10593 8533 10607 8547
rect 10493 8473 10507 8487
rect 10573 8493 10587 8507
rect 10613 8473 10627 8487
rect 10553 8433 10567 8447
rect 10493 8353 10507 8367
rect 10393 8333 10407 8347
rect 10453 8293 10467 8307
rect 10553 8333 10567 8347
rect 10553 8313 10567 8327
rect 10593 8313 10607 8327
rect 10693 8313 10707 8327
rect 10573 8293 10587 8307
rect 10573 8273 10587 8287
rect 10653 8293 10667 8307
rect 10593 8253 10607 8267
rect 10633 8253 10647 8267
rect 10493 8053 10507 8067
rect 10573 8053 10587 8067
rect 10373 8033 10387 8047
rect 10153 7853 10167 7867
rect 10093 7613 10107 7627
rect 9953 7533 9967 7547
rect 9913 7353 9927 7367
rect 9693 7173 9707 7187
rect 9673 6973 9687 6987
rect 10073 7533 10087 7547
rect 10113 7513 10127 7527
rect 10053 7413 10067 7427
rect 10053 7353 10067 7367
rect 10093 7353 10107 7367
rect 10033 7333 10047 7347
rect 10073 7333 10087 7347
rect 9953 7273 9967 7287
rect 10033 7273 10047 7287
rect 9553 6953 9567 6967
rect 9713 6953 9727 6967
rect 9793 6953 9807 6967
rect 9613 6893 9627 6907
rect 9893 6893 9907 6907
rect 9493 6773 9507 6787
rect 10053 6893 10067 6907
rect 10033 6813 10047 6827
rect 9653 6733 9667 6747
rect 9493 6573 9507 6587
rect 9633 6573 9647 6587
rect 9593 6433 9607 6447
rect 9953 6613 9967 6627
rect 9893 6573 9907 6587
rect 10113 6593 10127 6607
rect 9673 6433 9687 6447
rect 9693 6433 9707 6447
rect 9613 6413 9627 6427
rect 9653 6413 9667 6427
rect 9653 6393 9667 6407
rect 9553 6373 9567 6387
rect 9473 6353 9487 6367
rect 9593 6093 9607 6107
rect 9553 5933 9567 5947
rect 9633 6053 9647 6067
rect 9613 6033 9627 6047
rect 9453 5873 9467 5887
rect 9433 5633 9447 5647
rect 9473 5633 9487 5647
rect 9573 5633 9587 5647
rect 9453 5593 9467 5607
rect 9413 5573 9427 5587
rect 9433 5573 9447 5587
rect 9493 5573 9507 5587
rect 9393 5353 9407 5367
rect 9493 5413 9507 5427
rect 9533 5413 9547 5427
rect 9453 5393 9467 5407
rect 9513 5393 9527 5407
rect 9433 5193 9447 5207
rect 9373 5153 9387 5167
rect 9413 4993 9427 5007
rect 9353 4913 9367 4927
rect 9393 4913 9407 4927
rect 9313 4893 9327 4907
rect 9433 4933 9447 4947
rect 9273 4833 9287 4847
rect 9273 4753 9287 4767
rect 9293 4653 9307 4667
rect 9293 4453 9307 4467
rect 9273 4133 9287 4147
rect 9373 4653 9387 4667
rect 9333 4633 9347 4647
rect 9333 4553 9347 4567
rect 9313 4373 9327 4387
rect 9313 4313 9327 4327
rect 9313 4233 9327 4247
rect 9293 4013 9307 4027
rect 9313 4013 9327 4027
rect 9293 3993 9307 4007
rect 9193 3953 9207 3967
rect 9153 3933 9167 3947
rect 9253 3953 9267 3967
rect 9213 3853 9227 3867
rect 9233 3773 9247 3787
rect 9173 3653 9187 3667
rect 9113 3513 9127 3527
rect 9193 3513 9207 3527
rect 9133 3193 9147 3207
rect 9153 3173 9167 3187
rect 9093 3093 9107 3107
rect 9093 3073 9107 3087
rect 8973 2713 8987 2727
rect 8893 2593 8907 2607
rect 8933 2533 8947 2547
rect 8953 2513 8967 2527
rect 8913 2313 8927 2327
rect 8913 2233 8927 2247
rect 8893 2113 8907 2127
rect 8953 2113 8967 2127
rect 8873 1873 8887 1887
rect 8913 1833 8927 1847
rect 8833 1793 8847 1807
rect 8873 1793 8887 1807
rect 8813 1773 8827 1787
rect 8833 1773 8847 1787
rect 8933 1773 8947 1787
rect 8813 1653 8827 1667
rect 8873 1613 8887 1627
rect 8993 2553 9007 2567
rect 8993 2333 9007 2347
rect 9053 2653 9067 2667
rect 9193 3153 9207 3167
rect 9213 3053 9227 3067
rect 9193 3033 9207 3047
rect 9273 3913 9287 3927
rect 9373 4493 9387 4507
rect 9513 5353 9527 5367
rect 9493 5173 9507 5187
rect 9493 5113 9507 5127
rect 9493 5073 9507 5087
rect 9473 4813 9487 4827
rect 9453 4633 9467 4647
rect 9473 4533 9487 4547
rect 9433 4493 9447 4507
rect 9453 4493 9467 4507
rect 9413 4473 9427 4487
rect 9433 4433 9447 4447
rect 9393 4413 9407 4427
rect 9433 4413 9447 4427
rect 9373 4293 9387 4307
rect 9413 4193 9427 4207
rect 9393 4173 9407 4187
rect 9393 4153 9407 4167
rect 9333 3993 9347 4007
rect 9353 3753 9367 3767
rect 9373 3693 9387 3707
rect 9253 3013 9267 3027
rect 9293 3633 9307 3647
rect 9333 3553 9347 3567
rect 9293 2973 9307 2987
rect 9253 2733 9267 2747
rect 9293 2733 9307 2747
rect 9173 2613 9187 2627
rect 9233 2613 9247 2627
rect 9193 2553 9207 2567
rect 9213 2553 9227 2567
rect 8973 1813 8987 1827
rect 8893 1573 8907 1587
rect 8953 1573 8967 1587
rect 9033 2313 9047 2327
rect 9073 2293 9087 2307
rect 9013 2273 9027 2287
rect 9053 2273 9067 2287
rect 9093 2113 9107 2127
rect 9173 2473 9187 2487
rect 9173 2293 9187 2307
rect 9113 2073 9127 2087
rect 9193 2073 9207 2087
rect 9153 2053 9167 2067
rect 9153 1953 9167 1967
rect 9153 1773 9167 1787
rect 9193 1773 9207 1787
rect 9113 1713 9127 1727
rect 9093 1673 9107 1687
rect 9113 1613 9127 1627
rect 9193 1613 9207 1627
rect 9153 1593 9167 1607
rect 9093 1573 9107 1587
rect 8853 1553 8867 1567
rect 8993 1553 9007 1567
rect 9133 1553 9147 1567
rect 8933 1393 8947 1407
rect 8913 1353 8927 1367
rect 8813 1313 8827 1327
rect 8773 1293 8787 1307
rect 8773 1153 8787 1167
rect 8713 1113 8727 1127
rect 8673 1093 8687 1107
rect 9173 1373 9187 1387
rect 8933 1333 8947 1347
rect 8973 1333 8987 1347
rect 8993 1313 9007 1327
rect 9033 1293 9047 1307
rect 8953 1273 8967 1287
rect 9013 1253 9027 1267
rect 8953 1173 8967 1187
rect 8933 1133 8947 1147
rect 8933 1113 8947 1127
rect 8913 1093 8927 1107
rect 8693 1073 8707 1087
rect 8693 813 8707 827
rect 8373 773 8387 787
rect 8273 713 8287 727
rect 8493 773 8507 787
rect 8393 653 8407 667
rect 8373 633 8387 647
rect 8293 613 8307 627
rect 8373 453 8387 467
rect 8473 273 8487 287
rect 8473 213 8487 227
rect 8253 153 8267 167
rect 8273 153 8287 167
rect 8673 753 8687 767
rect 8673 693 8687 707
rect 8593 653 8607 667
rect 8573 613 8587 627
rect 8613 613 8627 627
rect 8633 613 8647 627
rect 8973 1093 8987 1107
rect 9173 1093 9187 1107
rect 9293 2253 9307 2267
rect 9273 2233 9287 2247
rect 9233 1793 9247 1807
rect 9533 5193 9547 5207
rect 9513 4433 9527 4447
rect 9493 4253 9507 4267
rect 9513 4093 9527 4107
rect 9553 5173 9567 5187
rect 9553 5153 9567 5167
rect 9553 4893 9567 4907
rect 9553 4653 9567 4667
rect 9553 4633 9567 4647
rect 9553 4153 9567 4167
rect 9533 4013 9547 4027
rect 10073 6573 10087 6587
rect 10133 6553 10147 6567
rect 9953 6453 9967 6467
rect 10093 6453 10107 6467
rect 9933 6413 9947 6427
rect 9873 6393 9887 6407
rect 9913 6393 9927 6407
rect 9793 6373 9807 6387
rect 9833 6373 9847 6387
rect 9813 6353 9827 6367
rect 9853 6353 9867 6367
rect 9813 6133 9827 6147
rect 9793 6093 9807 6107
rect 9833 6093 9847 6107
rect 9813 6033 9827 6047
rect 9873 6033 9887 6047
rect 9793 5953 9807 5967
rect 9673 5933 9687 5947
rect 9833 5913 9847 5927
rect 9773 5693 9787 5707
rect 9673 5653 9687 5667
rect 9713 5653 9727 5667
rect 9693 5613 9707 5627
rect 9673 5573 9687 5587
rect 9713 5573 9727 5587
rect 9693 5233 9707 5247
rect 9653 5193 9667 5207
rect 9633 5153 9647 5167
rect 9673 5153 9687 5167
rect 9593 5133 9607 5147
rect 9613 5113 9627 5127
rect 9633 4973 9647 4987
rect 9633 4913 9647 4927
rect 9613 4893 9627 4907
rect 9593 4873 9607 4887
rect 9593 4493 9607 4507
rect 9513 3973 9527 3987
rect 9533 3953 9547 3967
rect 9453 3913 9467 3927
rect 9433 3853 9447 3867
rect 9453 3833 9467 3847
rect 9513 3833 9527 3847
rect 9433 3713 9447 3727
rect 9473 3713 9487 3727
rect 9413 3693 9427 3707
rect 9393 3673 9407 3687
rect 9473 3673 9487 3687
rect 9453 3633 9467 3647
rect 9353 3513 9367 3527
rect 9393 3513 9407 3527
rect 9373 3493 9387 3507
rect 9373 3453 9387 3467
rect 9413 3453 9427 3467
rect 9433 3333 9447 3347
rect 9373 3173 9387 3187
rect 9453 3013 9467 3027
rect 9353 2713 9367 2727
rect 9513 3593 9527 3607
rect 9493 3533 9507 3547
rect 9513 3513 9527 3527
rect 9553 3873 9567 3887
rect 9553 3853 9567 3867
rect 9533 3213 9547 3227
rect 9513 3173 9527 3187
rect 9493 3133 9507 3147
rect 9473 2693 9487 2707
rect 9353 2573 9367 2587
rect 9413 2573 9427 2587
rect 9333 2333 9347 2347
rect 9393 2533 9407 2547
rect 9433 2533 9447 2547
rect 9533 2733 9547 2747
rect 9533 2693 9547 2707
rect 9513 2673 9527 2687
rect 9493 2533 9507 2547
rect 9473 2513 9487 2527
rect 9453 2473 9467 2487
rect 9353 2253 9367 2267
rect 9313 2233 9327 2247
rect 9433 2233 9447 2247
rect 9393 2113 9407 2127
rect 9353 2093 9367 2107
rect 9353 2073 9367 2087
rect 9413 2073 9427 2087
rect 9373 2053 9387 2067
rect 9353 1793 9367 1807
rect 9373 1773 9387 1787
rect 9333 1713 9347 1727
rect 9293 1613 9307 1627
rect 9213 1593 9227 1607
rect 9413 1653 9427 1667
rect 9413 1593 9427 1607
rect 9333 1573 9347 1587
rect 9353 1573 9367 1587
rect 9393 1573 9407 1587
rect 9273 1333 9287 1347
rect 9213 1293 9227 1307
rect 9293 1293 9307 1307
rect 9253 1253 9267 1267
rect 9273 1253 9287 1267
rect 9273 1153 9287 1167
rect 9233 1133 9247 1147
rect 9233 1113 9247 1127
rect 9253 1093 9267 1107
rect 8753 1053 8767 1067
rect 8733 653 8747 667
rect 8693 613 8707 627
rect 8713 613 8727 627
rect 8573 553 8587 567
rect 8553 373 8567 387
rect 8573 353 8587 367
rect 8613 333 8627 347
rect 8433 133 8447 147
rect 8633 133 8647 147
rect 8673 133 8687 147
rect 8713 133 8727 147
rect 8793 993 8807 1007
rect 8773 953 8787 967
rect 9253 933 9267 947
rect 9133 853 9147 867
rect 9173 853 9187 867
rect 8793 833 8807 847
rect 8893 813 8907 827
rect 9153 813 9167 827
rect 8933 793 8947 807
rect 8913 733 8927 747
rect 8893 713 8907 727
rect 8833 673 8847 687
rect 9153 673 9167 687
rect 9033 633 9047 647
rect 9113 633 9127 647
rect 8813 333 8827 347
rect 9013 333 9027 347
rect 8853 313 8867 327
rect 8833 293 8847 307
rect 8993 173 9007 187
rect 8813 153 8827 167
rect 8773 133 8787 147
rect 9133 613 9147 627
rect 9033 293 9047 307
rect 9413 893 9427 907
rect 9313 873 9327 887
rect 9393 873 9407 887
rect 9353 853 9367 867
rect 9373 833 9387 847
rect 9413 833 9427 847
rect 9353 813 9367 827
rect 9333 753 9347 767
rect 9353 673 9367 687
rect 9393 673 9407 687
rect 9333 653 9347 667
rect 9313 633 9327 647
rect 9373 633 9387 647
rect 9293 473 9307 487
rect 9113 333 9127 347
rect 9393 573 9407 587
rect 9473 2253 9487 2267
rect 9513 2213 9527 2227
rect 9493 2053 9507 2067
rect 9513 1773 9527 1787
rect 9493 1753 9507 1767
rect 9453 1633 9467 1647
rect 9453 1573 9467 1587
rect 9453 1333 9467 1347
rect 9493 1333 9507 1347
rect 9473 1233 9487 1247
rect 9473 1133 9487 1147
rect 9513 1093 9527 1107
rect 9453 713 9467 727
rect 9673 4793 9687 4807
rect 9653 4773 9667 4787
rect 9653 4693 9667 4707
rect 9733 5493 9747 5507
rect 9733 5433 9747 5447
rect 9733 5413 9747 5427
rect 9793 5413 9807 5427
rect 9713 4793 9727 4807
rect 9713 4673 9727 4687
rect 9693 4653 9707 4667
rect 9673 4533 9687 4547
rect 9713 4473 9727 4487
rect 9693 4453 9707 4467
rect 9673 4433 9687 4447
rect 9653 4413 9667 4427
rect 9713 4413 9727 4427
rect 9633 4213 9647 4227
rect 9653 4193 9667 4207
rect 9613 4173 9627 4187
rect 9613 4153 9627 4167
rect 9633 4133 9647 4147
rect 9613 3633 9627 3647
rect 9593 3593 9607 3607
rect 9593 3573 9607 3587
rect 9573 3513 9587 3527
rect 9613 3513 9627 3527
rect 9693 4393 9707 4407
rect 9673 4153 9687 4167
rect 9713 4173 9727 4187
rect 9693 4133 9707 4147
rect 9813 5113 9827 5127
rect 9853 5333 9867 5347
rect 9933 5673 9947 5687
rect 10073 6433 10087 6447
rect 10113 6393 10127 6407
rect 10073 6133 10087 6147
rect 10093 6113 10107 6127
rect 10173 7833 10187 7847
rect 10273 7893 10287 7907
rect 10373 7893 10387 7907
rect 10233 7813 10247 7827
rect 10173 7633 10187 7647
rect 10173 7513 10187 7527
rect 10173 7493 10187 7507
rect 10273 7433 10287 7447
rect 10233 7113 10247 7127
rect 10253 7113 10267 7127
rect 10333 7793 10347 7807
rect 10353 7633 10367 7647
rect 10533 7813 10547 7827
rect 10593 7853 10607 7867
rect 10553 7793 10567 7807
rect 10633 7833 10647 7847
rect 10613 7813 10627 7827
rect 10533 7573 10547 7587
rect 10473 7553 10487 7567
rect 10313 7533 10327 7547
rect 10333 7513 10347 7527
rect 10373 7413 10387 7427
rect 10313 7353 10327 7367
rect 10553 7553 10567 7567
rect 10593 7553 10607 7567
rect 10533 7513 10547 7527
rect 10573 7513 10587 7527
rect 10533 7373 10547 7387
rect 10553 7373 10567 7387
rect 10573 7373 10587 7387
rect 10473 7333 10487 7347
rect 10473 7113 10487 7127
rect 10253 6873 10267 6887
rect 10233 6853 10247 6867
rect 10153 6113 10167 6127
rect 10053 6093 10067 6107
rect 10133 6093 10147 6107
rect 10013 5913 10027 5927
rect 10533 7133 10547 7147
rect 10673 8073 10687 8087
rect 10653 7813 10667 7827
rect 10813 9493 10827 9507
rect 10773 9473 10787 9487
rect 10753 9453 10767 9467
rect 10753 9273 10767 9287
rect 10713 8073 10727 8087
rect 10733 8053 10747 8067
rect 10693 7933 10707 7947
rect 10733 7913 10747 7927
rect 10713 7893 10727 7907
rect 10693 7653 10707 7667
rect 10673 7553 10687 7567
rect 10733 7553 10747 7567
rect 10693 7513 10707 7527
rect 10633 7373 10647 7387
rect 10713 7373 10727 7387
rect 10613 7113 10627 7127
rect 10513 7093 10527 7107
rect 10633 7093 10647 7107
rect 10473 7073 10487 7087
rect 10513 7073 10527 7087
rect 10553 7073 10567 7087
rect 10313 7053 10327 7067
rect 10493 7053 10507 7067
rect 10393 6933 10407 6947
rect 10513 6933 10527 6947
rect 10293 6873 10307 6887
rect 10333 6873 10347 6887
rect 10313 6853 10327 6867
rect 10333 6573 10347 6587
rect 10273 6433 10287 6447
rect 10373 6433 10387 6447
rect 10313 6393 10327 6407
rect 10293 6373 10307 6387
rect 10353 6393 10367 6407
rect 10293 6353 10307 6367
rect 10313 6353 10327 6367
rect 10253 6053 10267 6067
rect 10093 5933 10107 5947
rect 10173 5933 10187 5947
rect 10573 7053 10587 7067
rect 10573 6873 10587 6887
rect 10553 6853 10567 6867
rect 10653 6813 10667 6827
rect 10533 6733 10547 6747
rect 10573 6733 10587 6747
rect 10533 6593 10547 6607
rect 10473 6573 10487 6587
rect 10493 6573 10507 6587
rect 10473 6373 10487 6387
rect 10413 6133 10427 6147
rect 10333 5993 10347 6007
rect 10113 5913 10127 5927
rect 10073 5873 10087 5887
rect 10033 5733 10047 5747
rect 10013 5633 10027 5647
rect 10133 5873 10147 5887
rect 9953 5613 9967 5627
rect 9993 5613 10007 5627
rect 9893 5173 9907 5187
rect 9913 5173 9927 5187
rect 9833 5073 9847 5087
rect 9873 5113 9887 5127
rect 9773 4953 9787 4967
rect 9793 4933 9807 4947
rect 9773 4913 9787 4927
rect 9873 4993 9887 5007
rect 10113 5613 10127 5627
rect 9973 5593 9987 5607
rect 10053 5453 10067 5467
rect 9993 5413 10007 5427
rect 10033 5393 10047 5407
rect 10053 5373 10067 5387
rect 10113 5373 10127 5387
rect 9973 4973 9987 4987
rect 9873 4933 9887 4947
rect 9913 4933 9927 4947
rect 9953 4933 9967 4947
rect 9893 4913 9907 4927
rect 9933 4913 9947 4927
rect 9853 4893 9867 4907
rect 9833 4793 9847 4807
rect 9793 4753 9807 4767
rect 9773 4673 9787 4687
rect 9813 4673 9827 4687
rect 9793 4653 9807 4667
rect 9753 4593 9767 4607
rect 9753 4473 9767 4487
rect 9753 4393 9767 4407
rect 9753 4353 9767 4367
rect 9753 4213 9767 4227
rect 9733 4153 9747 4167
rect 9733 4133 9747 4147
rect 9713 4033 9727 4047
rect 9673 3993 9687 4007
rect 9713 3993 9727 4007
rect 9753 3993 9767 4007
rect 9653 3673 9667 3687
rect 9793 4393 9807 4407
rect 9933 4693 9947 4707
rect 9853 4673 9867 4687
rect 9933 4653 9947 4667
rect 9953 4653 9967 4667
rect 9893 4613 9907 4627
rect 9873 4473 9887 4487
rect 9873 4433 9887 4447
rect 9933 4513 9947 4527
rect 9953 4433 9967 4447
rect 9873 4273 9887 4287
rect 9833 4213 9847 4227
rect 9913 4213 9927 4227
rect 9933 4213 9947 4227
rect 9873 4193 9887 4207
rect 9813 4173 9827 4187
rect 9793 3953 9807 3967
rect 9773 3793 9787 3807
rect 9713 3773 9727 3787
rect 9733 3773 9747 3787
rect 9733 3733 9747 3747
rect 9693 3693 9707 3707
rect 9713 3673 9727 3687
rect 9693 3593 9707 3607
rect 9673 3453 9687 3467
rect 9653 3333 9667 3347
rect 9593 3273 9607 3287
rect 9633 3273 9647 3287
rect 9573 2753 9587 2767
rect 9553 2213 9567 2227
rect 9573 1873 9587 1887
rect 9553 1793 9567 1807
rect 9553 1333 9567 1347
rect 9613 3253 9627 3267
rect 9613 3213 9627 3227
rect 9633 3193 9647 3207
rect 9633 3093 9647 3107
rect 9673 3033 9687 3047
rect 9693 2773 9707 2787
rect 9673 2753 9687 2767
rect 9653 2553 9667 2567
rect 9653 2313 9667 2327
rect 9653 2273 9667 2287
rect 9613 2233 9627 2247
rect 9613 2153 9627 2167
rect 9733 3593 9747 3607
rect 9613 2093 9627 2107
rect 9633 2073 9647 2087
rect 9673 2073 9687 2087
rect 9653 2053 9667 2067
rect 9753 3573 9767 3587
rect 9833 4153 9847 4167
rect 9853 4153 9867 4167
rect 9893 4133 9907 4147
rect 9893 4093 9907 4107
rect 9873 3993 9887 4007
rect 9833 3693 9847 3707
rect 9753 3493 9767 3507
rect 9733 2333 9747 2347
rect 9853 3513 9867 3527
rect 9873 3513 9887 3527
rect 9873 3493 9887 3507
rect 9833 3433 9847 3447
rect 9853 3433 9867 3447
rect 9793 3233 9807 3247
rect 9833 3033 9847 3047
rect 9773 2733 9787 2747
rect 9833 2733 9847 2747
rect 9793 2713 9807 2727
rect 9813 2713 9827 2727
rect 9813 2553 9827 2567
rect 9813 2353 9827 2367
rect 9813 2333 9827 2347
rect 9793 2313 9807 2327
rect 9753 2293 9767 2307
rect 9733 2273 9747 2287
rect 9713 2153 9727 2167
rect 9593 1793 9607 1807
rect 9613 1793 9627 1807
rect 9653 1773 9667 1787
rect 9593 1753 9607 1767
rect 9593 1613 9607 1627
rect 9613 1613 9627 1627
rect 9633 1593 9647 1607
rect 9613 1573 9627 1587
rect 9653 1553 9667 1567
rect 9653 1373 9667 1387
rect 9633 1273 9647 1287
rect 9593 1013 9607 1027
rect 9573 853 9587 867
rect 9633 913 9647 927
rect 9613 773 9627 787
rect 9613 733 9627 747
rect 9573 613 9587 627
rect 9633 573 9647 587
rect 9373 553 9387 567
rect 9433 553 9447 567
rect 9273 333 9287 347
rect 9333 333 9347 347
rect 9073 273 9087 287
rect 9053 233 9067 247
rect 9313 313 9327 327
rect 9293 293 9307 307
rect 9493 453 9507 467
rect 9533 373 9547 387
rect 9753 2153 9767 2167
rect 9753 2133 9767 2147
rect 9753 2053 9767 2067
rect 9933 4173 9947 4187
rect 9933 4133 9947 4147
rect 10153 5813 10167 5827
rect 10153 5613 10167 5627
rect 10133 5333 10147 5347
rect 10153 5173 10167 5187
rect 10113 5153 10127 5167
rect 10133 5153 10147 5167
rect 10093 5033 10107 5047
rect 10113 4973 10127 4987
rect 10153 4953 10167 4967
rect 10053 4933 10067 4947
rect 10093 4933 10107 4947
rect 10133 4933 10147 4947
rect 10313 5913 10327 5927
rect 10253 5893 10267 5907
rect 10233 5713 10247 5727
rect 10193 5673 10207 5687
rect 10333 5693 10347 5707
rect 10313 5653 10327 5667
rect 10273 5633 10287 5647
rect 10313 5633 10327 5647
rect 10333 5633 10347 5647
rect 10253 5613 10267 5627
rect 10293 5593 10307 5607
rect 10213 5513 10227 5527
rect 10253 5493 10267 5507
rect 10233 5473 10247 5487
rect 10273 5433 10287 5447
rect 10293 5393 10307 5407
rect 10253 5333 10267 5347
rect 10193 4933 10207 4947
rect 10133 4913 10147 4927
rect 10173 4913 10187 4927
rect 10053 4813 10067 4827
rect 10053 4773 10067 4787
rect 10013 4673 10027 4687
rect 9973 4093 9987 4107
rect 9973 4053 9987 4067
rect 9913 3973 9927 3987
rect 9953 3973 9967 3987
rect 9993 3973 10007 3987
rect 9913 3713 9927 3727
rect 10033 4653 10047 4667
rect 10113 4653 10127 4667
rect 10073 4433 10087 4447
rect 10073 4393 10087 4407
rect 10053 4293 10067 4307
rect 10033 3973 10047 3987
rect 10013 3933 10027 3947
rect 9973 3713 9987 3727
rect 9973 3653 9987 3667
rect 9953 3553 9967 3567
rect 9933 3433 9947 3447
rect 9873 3293 9887 3307
rect 9893 3293 9907 3307
rect 9913 3253 9927 3267
rect 9953 3193 9967 3207
rect 9893 3053 9907 3067
rect 9933 3053 9947 3067
rect 9873 3033 9887 3047
rect 9913 3033 9927 3047
rect 9873 2993 9887 3007
rect 9933 3013 9947 3027
rect 9853 2713 9867 2727
rect 9853 2593 9867 2607
rect 9893 2973 9907 2987
rect 9873 2553 9887 2567
rect 9913 2693 9927 2707
rect 9933 2533 9947 2547
rect 9913 2513 9927 2527
rect 9853 2353 9867 2367
rect 9913 2293 9927 2307
rect 9853 2273 9867 2287
rect 9833 2253 9847 2267
rect 9833 2073 9847 2087
rect 9833 2053 9847 2067
rect 9873 2053 9887 2067
rect 9813 1853 9827 1867
rect 9893 2033 9907 2047
rect 9873 1853 9887 1867
rect 9833 1813 9847 1827
rect 9813 1793 9827 1807
rect 9853 1793 9867 1807
rect 9833 1733 9847 1747
rect 9773 1713 9787 1727
rect 9793 1713 9807 1727
rect 9813 1613 9827 1627
rect 9733 1593 9747 1607
rect 9793 1593 9807 1607
rect 9693 1293 9707 1307
rect 9773 1293 9787 1307
rect 9353 133 9367 147
rect 9153 113 9167 127
rect 9653 473 9667 487
rect 9673 393 9687 407
rect 9733 1273 9747 1287
rect 9873 1273 9887 1287
rect 9733 1193 9747 1207
rect 9913 1133 9927 1147
rect 9773 1093 9787 1107
rect 9753 1073 9767 1087
rect 9713 973 9727 987
rect 9773 973 9787 987
rect 9733 373 9747 387
rect 9713 333 9727 347
rect 9753 313 9767 327
rect 9793 293 9807 307
rect 9693 233 9707 247
rect 9833 793 9847 807
rect 9993 3513 10007 3527
rect 9993 3193 10007 3207
rect 9973 2793 9987 2807
rect 10093 4153 10107 4167
rect 10073 3973 10087 3987
rect 10093 3913 10107 3927
rect 10073 3853 10087 3867
rect 10073 3753 10087 3767
rect 10073 3513 10087 3527
rect 10193 4673 10207 4687
rect 10173 4493 10187 4507
rect 10193 4433 10207 4447
rect 10153 4393 10167 4407
rect 10173 4133 10187 4147
rect 10113 3813 10127 3827
rect 10273 5133 10287 5147
rect 10353 5453 10367 5467
rect 10533 6433 10547 6447
rect 10593 6553 10607 6567
rect 10633 6493 10647 6507
rect 10593 6453 10607 6467
rect 10553 6413 10567 6427
rect 10573 6393 10587 6407
rect 10553 6373 10567 6387
rect 10693 6593 10707 6607
rect 10673 6353 10687 6367
rect 10833 9413 10847 9427
rect 10893 9733 10907 9747
rect 10893 9293 10907 9307
rect 10933 9913 10947 9927
rect 10933 9413 10947 9427
rect 10913 9273 10927 9287
rect 10873 9233 10887 9247
rect 10853 9213 10867 9227
rect 10893 9213 10907 9227
rect 10793 9013 10807 9027
rect 10833 8993 10847 9007
rect 10853 8973 10867 8987
rect 10873 8873 10887 8887
rect 10773 8813 10787 8827
rect 10813 8813 10827 8827
rect 10813 8793 10827 8807
rect 10853 8793 10867 8807
rect 10793 8773 10807 8787
rect 10833 8753 10847 8767
rect 10813 8513 10827 8527
rect 10773 8493 10787 8507
rect 10813 8333 10827 8347
rect 10833 8073 10847 8087
rect 10773 8053 10787 8067
rect 10773 7913 10787 7927
rect 10813 7833 10827 7847
rect 10853 7833 10867 7847
rect 10833 7813 10847 7827
rect 10773 7573 10787 7587
rect 10773 7513 10787 7527
rect 10753 7373 10767 7387
rect 10833 7553 10847 7567
rect 10813 7513 10827 7527
rect 10833 7413 10847 7427
rect 10853 7373 10867 7387
rect 10733 7333 10747 7347
rect 10813 7333 10827 7347
rect 10773 7313 10787 7327
rect 10853 7313 10867 7327
rect 10753 7133 10767 7147
rect 10793 7093 10807 7107
rect 10773 7073 10787 7087
rect 10733 6913 10747 6927
rect 10773 6873 10787 6887
rect 10813 6873 10827 6887
rect 10753 6853 10767 6867
rect 10793 6853 10807 6867
rect 10913 8533 10927 8547
rect 11053 10893 11067 10907
rect 11093 10893 11107 10907
rect 11233 10933 11247 10947
rect 11193 10873 11207 10887
rect 11073 10753 11087 10767
rect 11013 10733 11027 10747
rect 11013 10693 11027 10707
rect 11113 10733 11127 10747
rect 11153 10713 11167 10727
rect 11133 10693 11147 10707
rect 11073 10453 11087 10467
rect 10993 10273 11007 10287
rect 11093 10293 11107 10307
rect 11053 10253 11067 10267
rect 11033 10233 11047 10247
rect 11073 10233 11087 10247
rect 11013 10213 11027 10227
rect 11053 10213 11067 10227
rect 10993 10193 11007 10207
rect 10973 9933 10987 9947
rect 10973 9773 10987 9787
rect 10913 8073 10927 8087
rect 10953 8073 10967 8087
rect 10953 8053 10967 8067
rect 10933 7833 10947 7847
rect 11013 9973 11027 9987
rect 11053 9973 11067 9987
rect 11033 9933 11047 9947
rect 11213 10453 11227 10467
rect 11193 9933 11207 9947
rect 11213 9893 11227 9907
rect 11093 9773 11107 9787
rect 11053 9733 11067 9747
rect 11113 9733 11127 9747
rect 10993 9513 11007 9527
rect 11033 9473 11047 9487
rect 11293 10933 11307 10947
rect 11293 10913 11307 10927
rect 11273 10873 11287 10887
rect 11293 10713 11307 10727
rect 11253 10653 11267 10667
rect 11333 10453 11347 10467
rect 11313 10273 11327 10287
rect 11253 10213 11267 10227
rect 11273 10173 11287 10187
rect 11333 9993 11347 10007
rect 11293 9953 11307 9967
rect 11273 9933 11287 9947
rect 11253 9913 11267 9927
rect 11333 9893 11347 9907
rect 11053 9433 11067 9447
rect 11113 9433 11127 9447
rect 11053 9273 11067 9287
rect 11253 9433 11267 9447
rect 11213 9413 11227 9427
rect 11173 9293 11187 9307
rect 11273 9293 11287 9307
rect 11153 9273 11167 9287
rect 10993 9253 11007 9267
rect 10993 9013 11007 9027
rect 10973 7613 10987 7627
rect 11033 8813 11047 8827
rect 11133 9253 11147 9267
rect 11133 9013 11147 9027
rect 11093 8873 11107 8887
rect 11153 8973 11167 8987
rect 11173 8973 11187 8987
rect 11273 8973 11287 8987
rect 11113 8813 11127 8827
rect 11053 8793 11067 8807
rect 11093 8773 11107 8787
rect 11113 8753 11127 8767
rect 11013 8533 11027 8547
rect 11033 8353 11047 8367
rect 11093 8273 11107 8287
rect 11013 8193 11027 8207
rect 11113 8073 11127 8087
rect 11033 7853 11047 7867
rect 10993 7513 11007 7527
rect 10993 7493 11007 7507
rect 10973 7433 10987 7447
rect 11033 7453 11047 7467
rect 11013 7433 11027 7447
rect 10953 7333 10967 7347
rect 10953 7073 10967 7087
rect 11033 7413 11047 7427
rect 11093 7573 11107 7587
rect 11053 7373 11067 7387
rect 11053 7333 11067 7347
rect 11053 7073 11067 7087
rect 11053 6913 11067 6927
rect 11033 6873 11047 6887
rect 11013 6853 11027 6867
rect 11093 6893 11107 6907
rect 10893 6813 10907 6827
rect 11013 6813 11027 6827
rect 10993 6633 11007 6647
rect 10993 6573 11007 6587
rect 10833 6493 10847 6507
rect 10813 6433 10827 6447
rect 10793 6413 10807 6427
rect 10853 6473 10867 6487
rect 10813 6353 10827 6367
rect 10673 6213 10687 6227
rect 10713 6213 10727 6227
rect 10513 6173 10527 6187
rect 10433 6093 10447 6107
rect 10413 5433 10427 5447
rect 10393 5133 10407 5147
rect 10333 4993 10347 5007
rect 10373 4993 10387 5007
rect 10313 4933 10327 4947
rect 10353 4973 10367 4987
rect 10313 4693 10327 4707
rect 10333 4673 10347 4687
rect 10413 4673 10427 4687
rect 10293 4653 10307 4667
rect 10313 4653 10327 4667
rect 10293 4593 10307 4607
rect 10253 4273 10267 4287
rect 10213 4073 10227 4087
rect 10193 3993 10207 4007
rect 10273 3993 10287 4007
rect 10233 3973 10247 3987
rect 10153 3673 10167 3687
rect 10133 3653 10147 3667
rect 10073 3453 10087 3467
rect 10113 3453 10127 3467
rect 10053 3253 10067 3267
rect 10033 3133 10047 3147
rect 10033 3033 10047 3047
rect 10053 3033 10067 3047
rect 10033 2813 10047 2827
rect 10053 2733 10067 2747
rect 10033 2713 10047 2727
rect 10013 2693 10027 2707
rect 10013 2493 10027 2507
rect 9973 2473 9987 2487
rect 10013 2313 10027 2327
rect 9973 2293 9987 2307
rect 9993 2213 10007 2227
rect 9973 2113 9987 2127
rect 10013 2093 10027 2107
rect 10173 3653 10187 3667
rect 10153 3273 10167 3287
rect 10113 3233 10127 3247
rect 10153 3233 10167 3247
rect 10133 3213 10147 3227
rect 10113 3053 10127 3067
rect 10193 3533 10207 3547
rect 10193 3473 10207 3487
rect 10193 3273 10207 3287
rect 10173 3173 10187 3187
rect 10173 3053 10187 3067
rect 10133 3033 10147 3047
rect 10233 3813 10247 3827
rect 10253 3333 10267 3347
rect 10213 3213 10227 3227
rect 10213 3153 10227 3167
rect 10193 3013 10207 3027
rect 10113 2853 10127 2867
rect 10113 2793 10127 2807
rect 10153 2793 10167 2807
rect 10093 2713 10107 2727
rect 10093 2513 10107 2527
rect 10133 2513 10147 2527
rect 10073 2493 10087 2507
rect 10073 2333 10087 2347
rect 10033 2033 10047 2047
rect 10113 2493 10127 2507
rect 10093 2293 10107 2307
rect 10093 2233 10107 2247
rect 10093 2033 10107 2047
rect 10133 2033 10147 2047
rect 10173 2253 10187 2267
rect 10073 1813 10087 1827
rect 10073 1793 10087 1807
rect 10113 1793 10127 1807
rect 10013 1753 10027 1767
rect 10033 1653 10047 1667
rect 10053 1653 10067 1667
rect 10013 1613 10027 1627
rect 10073 1633 10087 1647
rect 10053 1613 10067 1627
rect 9973 1373 9987 1387
rect 10013 1373 10027 1387
rect 9953 1353 9967 1367
rect 9973 1333 9987 1347
rect 10033 1333 10047 1347
rect 9953 1293 9967 1307
rect 10013 1273 10027 1287
rect 9993 1153 10007 1167
rect 10113 1353 10127 1367
rect 10093 1273 10107 1287
rect 10093 1253 10107 1267
rect 9973 1033 9987 1047
rect 10053 933 10067 947
rect 10073 833 10087 847
rect 9933 753 9947 767
rect 9833 693 9847 707
rect 9833 393 9847 407
rect 9893 393 9907 407
rect 9853 373 9867 387
rect 9833 233 9847 247
rect 9813 193 9827 207
rect 9813 173 9827 187
rect 10153 1813 10167 1827
rect 10133 473 10147 487
rect 9993 353 10007 367
rect 9873 333 9887 347
rect 9893 333 9907 347
rect 9993 313 10007 327
rect 10293 3713 10307 3727
rect 10373 4473 10387 4487
rect 10653 6053 10667 6067
rect 10513 5933 10527 5947
rect 10573 5873 10587 5887
rect 10473 5773 10487 5787
rect 10653 5673 10667 5687
rect 10513 5653 10527 5667
rect 10493 5633 10507 5647
rect 10653 5593 10667 5607
rect 10453 5513 10467 5527
rect 10573 5473 10587 5487
rect 10453 5173 10467 5187
rect 10433 4653 10447 4667
rect 10753 6193 10767 6207
rect 10693 5933 10707 5947
rect 10533 5193 10547 5207
rect 10633 5193 10647 5207
rect 10673 5193 10687 5207
rect 10493 5153 10507 5167
rect 10473 5133 10487 5147
rect 10453 4473 10467 4487
rect 10433 4453 10447 4467
rect 10393 4433 10407 4447
rect 10393 4353 10407 4367
rect 10333 4293 10347 4307
rect 10373 4213 10387 4227
rect 10453 4033 10467 4047
rect 10773 6113 10787 6127
rect 10773 5893 10787 5907
rect 10813 5893 10827 5907
rect 10793 5873 10807 5887
rect 10773 5713 10787 5727
rect 10733 5653 10747 5667
rect 10713 5633 10727 5647
rect 10753 5633 10767 5647
rect 10813 5633 10827 5647
rect 10813 5613 10827 5627
rect 10773 5493 10787 5507
rect 10833 5473 10847 5487
rect 10713 5193 10727 5207
rect 10533 5013 10547 5027
rect 10613 4993 10627 5007
rect 10533 4633 10547 4647
rect 10493 4533 10507 4547
rect 10493 4513 10507 4527
rect 10413 3993 10427 4007
rect 10473 3993 10487 4007
rect 10333 3973 10347 3987
rect 10393 3953 10407 3967
rect 10333 3833 10347 3847
rect 10453 3973 10467 3987
rect 10433 3953 10447 3967
rect 10473 3913 10487 3927
rect 10433 3833 10447 3847
rect 10313 3673 10327 3687
rect 10413 3733 10427 3747
rect 10413 3713 10427 3727
rect 10373 3613 10387 3627
rect 10373 3553 10387 3567
rect 10333 3533 10347 3547
rect 10333 3493 10347 3507
rect 10273 3313 10287 3327
rect 10253 3073 10267 3087
rect 10233 3033 10247 3047
rect 10233 2933 10247 2947
rect 10213 2713 10227 2727
rect 10213 2353 10227 2367
rect 10293 3233 10307 3247
rect 10353 3453 10367 3467
rect 10353 3213 10367 3227
rect 10313 3053 10327 3067
rect 10333 3053 10347 3067
rect 10393 3193 10407 3207
rect 10393 3173 10407 3187
rect 10373 3053 10387 3067
rect 10353 3013 10367 3027
rect 10373 2993 10387 3007
rect 10333 2973 10347 2987
rect 10353 2953 10367 2967
rect 10273 2753 10287 2767
rect 10333 2753 10347 2767
rect 10293 2733 10307 2747
rect 10273 2713 10287 2727
rect 10313 2713 10327 2727
rect 10253 2633 10267 2647
rect 10293 2553 10307 2567
rect 10253 2493 10267 2507
rect 10233 2333 10247 2347
rect 10273 2253 10287 2267
rect 10253 2233 10267 2247
rect 10233 2213 10247 2227
rect 10353 2693 10367 2707
rect 10333 2553 10347 2567
rect 10313 2513 10327 2527
rect 10333 2513 10347 2527
rect 10333 2493 10347 2507
rect 10313 2293 10327 2307
rect 10313 2253 10327 2267
rect 10353 2333 10367 2347
rect 10373 2313 10387 2327
rect 10353 2213 10367 2227
rect 10373 2193 10387 2207
rect 10433 3493 10447 3507
rect 10433 3073 10447 3087
rect 10433 2993 10447 3007
rect 10513 4453 10527 4467
rect 10693 5113 10707 5127
rect 10673 4913 10687 4927
rect 10593 4893 10607 4907
rect 10553 4553 10567 4567
rect 10533 4213 10547 4227
rect 10673 4573 10687 4587
rect 10573 4493 10587 4507
rect 10593 4453 10607 4467
rect 10653 4453 10667 4467
rect 10673 4413 10687 4427
rect 10633 4393 10647 4407
rect 10653 4213 10667 4227
rect 10573 4153 10587 4167
rect 10573 4133 10587 4147
rect 10573 4113 10587 4127
rect 10553 4033 10567 4047
rect 10533 3953 10547 3967
rect 10533 3873 10547 3887
rect 10513 3733 10527 3747
rect 10473 2933 10487 2947
rect 10413 2873 10427 2887
rect 10393 2153 10407 2167
rect 10313 2033 10327 2047
rect 10373 2033 10387 2047
rect 10353 2013 10367 2027
rect 10333 1853 10347 1867
rect 10373 1793 10387 1807
rect 10313 1753 10327 1767
rect 10253 1613 10267 1627
rect 10293 1613 10307 1627
rect 10293 1593 10307 1607
rect 10253 1553 10267 1567
rect 10213 1333 10227 1347
rect 10293 1333 10307 1347
rect 10253 1253 10267 1267
rect 10233 1233 10247 1247
rect 10213 1133 10227 1147
rect 10193 1113 10207 1127
rect 10233 1113 10247 1127
rect 10273 1073 10287 1087
rect 10213 893 10227 907
rect 10193 753 10207 767
rect 10173 393 10187 407
rect 10173 353 10187 367
rect 10053 253 10067 267
rect 10153 253 10167 267
rect 9853 213 9867 227
rect 9853 193 9867 207
rect 10193 313 10207 327
rect 10173 153 10187 167
rect 10333 1293 10347 1307
rect 10313 1113 10327 1127
rect 10333 1093 10347 1107
rect 10373 1593 10387 1607
rect 10493 2773 10507 2787
rect 10473 2753 10487 2767
rect 10493 2733 10507 2747
rect 10433 2713 10447 2727
rect 10473 2333 10487 2347
rect 10433 2293 10447 2307
rect 10453 2273 10467 2287
rect 10453 2233 10467 2247
rect 10473 2093 10487 2107
rect 10453 1813 10467 1827
rect 10413 1573 10427 1587
rect 10453 1293 10467 1307
rect 10433 1273 10447 1287
rect 10453 1213 10467 1227
rect 10533 3693 10547 3707
rect 10593 3973 10607 3987
rect 10633 3993 10647 4007
rect 10613 3893 10627 3907
rect 10593 3853 10607 3867
rect 10573 3833 10587 3847
rect 10633 3753 10647 3767
rect 10593 3733 10607 3747
rect 10633 3733 10647 3747
rect 10613 3713 10627 3727
rect 10573 3513 10587 3527
rect 10633 3553 10647 3567
rect 10613 3493 10627 3507
rect 10573 3253 10587 3267
rect 10553 3213 10567 3227
rect 10593 3133 10607 3147
rect 10633 3053 10647 3067
rect 10573 3033 10587 3047
rect 10593 2993 10607 3007
rect 10553 2973 10567 2987
rect 10573 2973 10587 2987
rect 10533 2953 10547 2967
rect 10533 2933 10547 2947
rect 10553 2753 10567 2767
rect 10533 2733 10547 2747
rect 10533 2573 10547 2587
rect 10513 2113 10527 2127
rect 10593 2713 10607 2727
rect 10573 2593 10587 2607
rect 10633 2993 10647 3007
rect 10693 4113 10707 4127
rect 10673 4053 10687 4067
rect 10873 6353 10887 6367
rect 11073 6613 11087 6627
rect 11033 6513 11047 6527
rect 11093 6513 11107 6527
rect 11153 7993 11167 8007
rect 11113 6473 11127 6487
rect 11253 8773 11267 8787
rect 11293 8753 11307 8767
rect 11293 8533 11307 8547
rect 11213 8313 11227 8327
rect 11233 8173 11247 8187
rect 11293 8353 11307 8367
rect 11273 7933 11287 7947
rect 11233 7873 11247 7887
rect 11293 7793 11307 7807
rect 11233 7593 11247 7607
rect 11293 7533 11307 7547
rect 11193 7513 11207 7527
rect 11173 6313 11187 6327
rect 10873 6113 10887 6127
rect 10973 6053 10987 6067
rect 10913 5913 10927 5927
rect 10893 5713 10907 5727
rect 10893 5593 10907 5607
rect 11053 6093 11067 6107
rect 11013 6053 11027 6067
rect 11033 6033 11047 6047
rect 11033 5933 11047 5947
rect 10993 5913 11007 5927
rect 11093 5893 11107 5907
rect 11013 5673 11027 5687
rect 10973 5633 10987 5647
rect 10993 5593 11007 5607
rect 10953 5473 10967 5487
rect 10993 5453 11007 5467
rect 10933 5413 10947 5427
rect 10913 5253 10927 5267
rect 10853 5193 10867 5207
rect 10873 5153 10887 5167
rect 10793 5133 10807 5147
rect 10893 5133 10907 5147
rect 10853 5093 10867 5107
rect 10813 4973 10827 4987
rect 10733 4933 10747 4947
rect 10813 4693 10827 4707
rect 10773 4673 10787 4687
rect 10793 4653 10807 4667
rect 10733 4593 10747 4607
rect 10753 4593 10767 4607
rect 10773 4553 10787 4567
rect 10773 4473 10787 4487
rect 10733 4393 10747 4407
rect 10733 4193 10747 4207
rect 10793 4413 10807 4427
rect 10813 4213 10827 4227
rect 11033 5433 11047 5447
rect 11073 5413 11087 5427
rect 11053 5393 11067 5407
rect 11073 5373 11087 5387
rect 10953 5193 10967 5207
rect 10933 5053 10947 5067
rect 10913 4893 10927 4907
rect 10913 4673 10927 4687
rect 10873 4613 10887 4627
rect 10893 4573 10907 4587
rect 10913 4513 10927 4527
rect 10913 4473 10927 4487
rect 10773 4173 10787 4187
rect 10833 4193 10847 4207
rect 10813 4173 10827 4187
rect 10853 4153 10867 4167
rect 10713 4013 10727 4027
rect 10713 3993 10727 4007
rect 10733 3973 10747 3987
rect 10713 3953 10727 3967
rect 10693 3913 10707 3927
rect 10673 3733 10687 3747
rect 10673 3593 10687 3607
rect 10693 3533 10707 3547
rect 10673 3513 10687 3527
rect 10653 2793 10667 2807
rect 10653 2773 10667 2787
rect 10613 2573 10627 2587
rect 10633 2533 10647 2547
rect 10693 3493 10707 3507
rect 10733 3933 10747 3947
rect 10793 4113 10807 4127
rect 10813 4053 10827 4067
rect 10793 4033 10807 4047
rect 10773 4013 10787 4027
rect 10753 3513 10767 3527
rect 10753 3213 10767 3227
rect 10733 3153 10747 3167
rect 10753 3033 10767 3047
rect 10713 2973 10727 2987
rect 10693 2773 10707 2787
rect 10733 2773 10747 2787
rect 10673 2753 10687 2767
rect 10713 2753 10727 2767
rect 10693 2553 10707 2567
rect 10653 2513 10667 2527
rect 10633 2273 10647 2287
rect 10553 2233 10567 2247
rect 10553 2173 10567 2187
rect 10533 2093 10547 2107
rect 10513 2073 10527 2087
rect 10513 2053 10527 2067
rect 10713 2293 10727 2307
rect 10753 2273 10767 2287
rect 10673 2233 10687 2247
rect 10693 2233 10707 2247
rect 10653 2093 10667 2107
rect 10573 2033 10587 2047
rect 10513 1813 10527 1827
rect 10553 1813 10567 1827
rect 10733 2193 10747 2207
rect 10573 1793 10587 1807
rect 10693 1793 10707 1807
rect 10513 1753 10527 1767
rect 10533 1753 10547 1767
rect 10573 1753 10587 1767
rect 10613 1613 10627 1627
rect 10693 1593 10707 1607
rect 10593 1573 10607 1587
rect 10533 1553 10547 1567
rect 10833 4013 10847 4027
rect 10813 3773 10827 3787
rect 10933 4193 10947 4207
rect 10913 4153 10927 4167
rect 10933 4153 10947 4167
rect 10873 3933 10887 3947
rect 10833 3713 10847 3727
rect 10853 3693 10867 3707
rect 10973 5153 10987 5167
rect 11133 5653 11147 5667
rect 11153 5653 11167 5667
rect 11113 5633 11127 5647
rect 11093 5113 11107 5127
rect 11133 5173 11147 5187
rect 11153 5153 11167 5167
rect 11153 5093 11167 5107
rect 11113 4953 11127 4967
rect 11053 4933 11067 4947
rect 11073 4913 11087 4927
rect 11013 4673 11027 4687
rect 11033 4653 11047 4667
rect 10993 4633 11007 4647
rect 11053 4573 11067 4587
rect 10993 4553 11007 4567
rect 10973 4053 10987 4067
rect 10953 4033 10967 4047
rect 10953 4013 10967 4027
rect 10933 3993 10947 4007
rect 11053 4273 11067 4287
rect 11013 4033 11027 4047
rect 10953 3973 10967 3987
rect 10933 3793 10947 3807
rect 10873 3673 10887 3687
rect 10813 3653 10827 3667
rect 10833 3533 10847 3547
rect 10853 3533 10867 3547
rect 10813 3513 10827 3527
rect 10913 3513 10927 3527
rect 10813 3213 10827 3227
rect 10853 3213 10867 3227
rect 10913 3213 10927 3227
rect 10833 3073 10847 3087
rect 10813 3053 10827 3067
rect 10793 3033 10807 3047
rect 10833 3033 10847 3047
rect 10873 3033 10887 3047
rect 10853 2993 10867 3007
rect 10793 2953 10807 2967
rect 10813 2773 10827 2787
rect 10833 2773 10847 2787
rect 10833 2593 10847 2607
rect 10793 2553 10807 2567
rect 10853 2533 10867 2547
rect 10833 2513 10847 2527
rect 10793 2153 10807 2167
rect 10533 1353 10547 1367
rect 10713 1353 10727 1367
rect 10513 1193 10527 1207
rect 10493 1173 10507 1187
rect 10433 1133 10447 1147
rect 10473 1133 10487 1147
rect 10393 1113 10407 1127
rect 10413 1113 10427 1127
rect 10373 1053 10387 1067
rect 10353 913 10367 927
rect 10293 873 10307 887
rect 10273 853 10287 867
rect 10333 853 10347 867
rect 10373 853 10387 867
rect 10233 833 10247 847
rect 10293 813 10307 827
rect 10293 793 10307 807
rect 10313 713 10327 727
rect 10253 633 10267 647
rect 10313 613 10327 627
rect 10313 593 10327 607
rect 10273 533 10287 547
rect 10313 493 10327 507
rect 10253 393 10267 407
rect 10273 393 10287 407
rect 10413 833 10427 847
rect 10393 793 10407 807
rect 10453 1113 10467 1127
rect 10513 1113 10527 1127
rect 10473 1093 10487 1107
rect 10813 2033 10827 2047
rect 10773 2013 10787 2027
rect 10793 2013 10807 2027
rect 10753 1813 10767 1827
rect 10753 1733 10767 1747
rect 10893 3013 10907 3027
rect 10873 2513 10887 2527
rect 10853 2293 10867 2307
rect 10873 2293 10887 2307
rect 10853 2093 10867 2107
rect 10833 2013 10847 2027
rect 10813 1813 10827 1827
rect 10833 1773 10847 1787
rect 10853 1773 10867 1787
rect 10793 1753 10807 1767
rect 10833 1753 10847 1767
rect 10793 1733 10807 1747
rect 10773 1713 10787 1727
rect 10773 1593 10787 1607
rect 10813 1593 10827 1607
rect 10753 1553 10767 1567
rect 10733 1333 10747 1347
rect 10593 1313 10607 1327
rect 10673 1313 10687 1327
rect 10713 1313 10727 1327
rect 10793 1413 10807 1427
rect 10593 1273 10607 1287
rect 10733 1273 10747 1287
rect 10713 1253 10727 1267
rect 10653 1233 10667 1247
rect 10693 1233 10707 1247
rect 10693 1173 10707 1187
rect 10653 1113 10667 1127
rect 10533 893 10547 907
rect 10533 733 10547 747
rect 10553 713 10567 727
rect 10513 633 10527 647
rect 10533 633 10547 647
rect 10593 633 10607 647
rect 10613 633 10627 647
rect 10513 593 10527 607
rect 10573 573 10587 587
rect 10613 573 10627 587
rect 10493 493 10507 507
rect 10333 333 10347 347
rect 10353 333 10367 347
rect 10293 133 10307 147
rect 9673 113 9687 127
rect 10073 113 10087 127
rect 10213 113 10227 127
rect 10633 433 10647 447
rect 10473 273 10487 287
rect 10533 153 10547 167
rect 10653 353 10667 367
rect 10753 1213 10767 1227
rect 10713 1113 10727 1127
rect 10813 1333 10827 1347
rect 10773 653 10787 667
rect 10753 593 10767 607
rect 10793 593 10807 607
rect 10733 433 10747 447
rect 10713 353 10727 367
rect 10693 293 10707 307
rect 10733 293 10747 307
rect 10713 193 10727 207
rect 10753 153 10767 167
rect 10833 153 10847 167
rect 10873 1273 10887 1287
rect 10993 3753 11007 3767
rect 10973 3693 10987 3707
rect 10953 3673 10967 3687
rect 10933 3193 10947 3207
rect 10973 3533 10987 3547
rect 10973 2973 10987 2987
rect 10913 2793 10927 2807
rect 10953 2793 10967 2807
rect 10913 2773 10927 2787
rect 10953 2773 10967 2787
rect 10933 2753 10947 2767
rect 10933 2593 10947 2607
rect 10953 2573 10967 2587
rect 10933 2273 10947 2287
rect 10913 2233 10927 2247
rect 10933 2213 10947 2227
rect 10993 2773 11007 2787
rect 10973 2133 10987 2147
rect 10973 2113 10987 2127
rect 10953 1853 10967 1867
rect 11033 3993 11047 4007
rect 11093 4653 11107 4667
rect 11113 4633 11127 4647
rect 11133 4553 11147 4567
rect 11153 4513 11167 4527
rect 11133 4493 11147 4507
rect 11093 4213 11107 4227
rect 11133 4213 11147 4227
rect 11113 4193 11127 4207
rect 11093 4013 11107 4027
rect 11053 3673 11067 3687
rect 11073 3653 11087 3667
rect 11053 3513 11067 3527
rect 11093 3513 11107 3527
rect 11093 3213 11107 3227
rect 11073 3193 11087 3207
rect 11053 3173 11067 3187
rect 11033 3033 11047 3047
rect 11053 3013 11067 3027
rect 11053 2973 11067 2987
rect 11033 2773 11047 2787
rect 11013 2713 11027 2727
rect 11073 2953 11087 2967
rect 11073 2813 11087 2827
rect 11073 2733 11087 2747
rect 11053 2533 11067 2547
rect 11093 2533 11107 2547
rect 11073 2513 11087 2527
rect 11033 2493 11047 2507
rect 11073 2493 11087 2507
rect 11053 2333 11067 2347
rect 11013 2313 11027 2327
rect 11013 2253 11027 2267
rect 11073 2293 11087 2307
rect 11033 2093 11047 2107
rect 10993 1813 11007 1827
rect 10973 1773 10987 1787
rect 10933 1753 10947 1767
rect 11033 1753 11047 1767
rect 10913 1573 10927 1587
rect 11013 1573 11027 1587
rect 10933 1413 10947 1427
rect 10913 1353 10927 1367
rect 10913 1313 10927 1327
rect 10973 1333 10987 1347
rect 10953 1313 10967 1327
rect 11033 1553 11047 1567
rect 11013 1373 11027 1387
rect 11033 1333 11047 1347
rect 11013 1313 11027 1327
rect 10993 1253 11007 1267
rect 10933 1233 10947 1247
rect 10973 1153 10987 1167
rect 10993 1133 11007 1147
rect 10953 1113 10967 1127
rect 10913 853 10927 867
rect 10893 413 10907 427
rect 10893 333 10907 347
rect 11053 1153 11067 1167
rect 11093 1853 11107 1867
rect 11073 853 11087 867
rect 11053 793 11067 807
rect 10973 673 10987 687
rect 11013 673 11027 687
rect 10993 653 11007 667
rect 11013 653 11027 667
rect 11033 633 11047 647
rect 10973 413 10987 427
rect 11013 413 11027 427
rect 11033 413 11047 427
rect 10933 373 10947 387
rect 10973 373 10987 387
rect 11013 373 11027 387
rect 10953 353 10967 367
rect 11033 353 11047 367
rect 10993 333 11007 347
rect 10953 313 10967 327
rect 10873 173 10887 187
rect 10913 173 10927 187
rect 11133 3753 11147 3767
rect 11133 3733 11147 3747
rect 11253 7393 11267 7407
rect 11313 7313 11327 7327
rect 11293 7053 11307 7067
rect 11253 7013 11267 7027
rect 11213 6913 11227 6927
rect 11313 6913 11327 6927
rect 11253 6893 11267 6907
rect 11233 6853 11247 6867
rect 11293 6633 11307 6647
rect 11213 6573 11227 6587
rect 11293 6593 11307 6607
rect 11253 6493 11267 6507
rect 11253 6373 11267 6387
rect 11293 6373 11307 6387
rect 11213 6313 11227 6327
rect 11313 6293 11327 6307
rect 11253 6073 11267 6087
rect 11273 6053 11287 6067
rect 11293 5973 11307 5987
rect 11233 5893 11247 5907
rect 11273 5893 11287 5907
rect 11213 5873 11227 5887
rect 11253 5873 11267 5887
rect 11273 5853 11287 5867
rect 11213 5793 11227 5807
rect 11273 5673 11287 5687
rect 11213 5653 11227 5667
rect 11253 5653 11267 5667
rect 11233 5633 11247 5647
rect 11213 5153 11227 5167
rect 11193 4613 11207 4627
rect 11213 4033 11227 4047
rect 11213 4013 11227 4027
rect 11173 3993 11187 4007
rect 11193 3973 11207 3987
rect 11153 3673 11167 3687
rect 11153 3513 11167 3527
rect 11173 3293 11187 3307
rect 11153 3213 11167 3227
rect 11173 3193 11187 3207
rect 11253 5453 11267 5467
rect 11273 5413 11287 5427
rect 11313 5393 11327 5407
rect 11353 8533 11367 8547
rect 11253 5373 11267 5387
rect 11333 5373 11347 5387
rect 11273 4973 11287 4987
rect 11293 4693 11307 4707
rect 11273 4573 11287 4587
rect 11273 4373 11287 4387
rect 11253 3953 11267 3967
rect 11333 4593 11347 4607
rect 11333 4493 11347 4507
rect 11293 3733 11307 3747
rect 11353 3973 11367 3987
rect 11293 3693 11307 3707
rect 11333 3673 11347 3687
rect 11313 3553 11327 3567
rect 11293 3513 11307 3527
rect 11233 3213 11247 3227
rect 11273 3213 11287 3227
rect 11193 3153 11207 3167
rect 11213 2793 11227 2807
rect 11133 2773 11147 2787
rect 11193 2773 11207 2787
rect 11133 2733 11147 2747
rect 11173 2713 11187 2727
rect 11153 2353 11167 2367
rect 11193 2333 11207 2347
rect 11193 2313 11207 2327
rect 11153 2293 11167 2307
rect 11133 2273 11147 2287
rect 11173 2273 11187 2287
rect 11153 2133 11167 2147
rect 11133 1133 11147 1147
rect 11133 833 11147 847
rect 11133 793 11147 807
rect 11173 1813 11187 1827
rect 11173 1593 11187 1607
rect 11293 3193 11307 3207
rect 11293 2993 11307 3007
rect 11333 3173 11347 3187
rect 11333 3153 11347 3167
rect 11253 2953 11267 2967
rect 11293 2533 11307 2547
rect 11273 2513 11287 2527
rect 11253 2493 11267 2507
rect 11253 2213 11267 2227
rect 11313 2493 11327 2507
rect 11313 2313 11327 2327
rect 11273 2113 11287 2127
rect 11293 2113 11307 2127
rect 11273 2093 11287 2107
rect 11293 1833 11307 1847
rect 11253 1813 11267 1827
rect 11233 1773 11247 1787
rect 11193 1553 11207 1567
rect 11173 1273 11187 1287
rect 11213 1133 11227 1147
rect 11293 1753 11307 1767
rect 11253 1713 11267 1727
rect 11193 633 11207 647
rect 11173 433 11187 447
rect 11153 393 11167 407
rect 11193 393 11207 407
rect 11113 373 11127 387
rect 11153 373 11167 387
rect 11173 353 11187 367
rect 10973 173 10987 187
rect 11093 173 11107 187
rect 11193 173 11207 187
rect 10933 153 10947 167
rect 11233 873 11247 887
rect 11273 833 11287 847
rect 11233 653 11247 667
rect 11253 413 11267 427
rect 11353 2573 11367 2587
rect 11353 2533 11367 2547
rect 11333 353 11347 367
rect 11353 193 11367 207
rect 10853 133 10867 147
rect 11173 133 11187 147
rect 11213 133 11227 147
rect 10513 113 10527 127
rect 10813 113 10827 127
rect 10033 93 10047 107
rect 10453 93 10467 107
rect 9013 73 9027 87
<< metal3 >>
rect 4147 11296 4173 11304
rect 4347 11296 4373 11304
rect 7027 11296 7173 11304
rect 8167 11296 8193 11304
rect 2747 11236 3484 11244
rect 627 11216 793 11224
rect 947 11216 973 11224
rect 987 11216 1353 11224
rect 1627 11216 1793 11224
rect 1907 11216 2033 11224
rect 2047 11216 2713 11224
rect 3387 11216 3453 11224
rect 3476 11224 3484 11236
rect 4667 11236 6113 11244
rect 6147 11236 6773 11244
rect 3476 11216 4704 11224
rect 1027 11196 1784 11204
rect 1776 11187 1784 11196
rect 1827 11196 2673 11204
rect 2687 11196 2773 11204
rect 2787 11196 3413 11204
rect 3507 11196 3753 11204
rect 4187 11196 4593 11204
rect 4607 11196 4673 11204
rect 4696 11204 4704 11216
rect 4867 11216 5393 11224
rect 5407 11216 5553 11224
rect 6127 11216 6493 11224
rect 6516 11216 7273 11224
rect 6516 11204 6524 11216
rect 7687 11216 8153 11224
rect 8967 11216 9173 11224
rect 4696 11196 6524 11204
rect 6747 11196 6764 11204
rect 587 11176 633 11184
rect 787 11176 933 11184
rect 1007 11176 1193 11184
rect 1247 11176 1473 11184
rect 1547 11176 1733 11184
rect 1927 11176 2193 11184
rect 2307 11176 2453 11184
rect 2507 11176 2693 11184
rect 3416 11184 3424 11193
rect 3416 11176 4113 11184
rect 4307 11176 4373 11184
rect 5127 11176 5293 11184
rect 5347 11176 5533 11184
rect 5587 11176 6133 11184
rect 6527 11176 6733 11184
rect 6756 11167 6764 11196
rect 6987 11196 7004 11204
rect 6787 11176 6973 11184
rect 6996 11167 7004 11196
rect 7447 11196 7464 11204
rect 7227 11176 7253 11184
rect 7287 11176 7433 11184
rect 7456 11167 7464 11196
rect 8127 11196 8373 11204
rect 8436 11196 8673 11204
rect 8187 11176 8213 11184
rect 567 11156 953 11164
rect 1887 11156 2793 11164
rect 3447 11156 3713 11164
rect 4407 11156 4613 11164
rect 5707 11156 5913 11164
rect 6287 11156 6333 11164
rect 7147 11156 7193 11164
rect 7247 11156 7413 11164
rect 8167 11156 8193 11164
rect 8416 11164 8424 11193
rect 8436 11187 8444 11196
rect 8727 11196 8973 11204
rect 8987 11196 9153 11204
rect 9627 11196 10113 11204
rect 8667 11176 8933 11184
rect 8947 11176 8993 11184
rect 9407 11176 9613 11184
rect 9667 11176 9684 11184
rect 8416 11156 8453 11164
rect 8707 11156 9213 11164
rect 9676 11147 9684 11176
rect 9707 11176 9873 11184
rect 10247 11176 10373 11184
rect 10427 11176 10613 11184
rect 10747 11176 10833 11184
rect 10887 11176 11073 11184
rect 10147 11156 10353 11164
rect 10947 11156 11053 11164
rect 347 11136 573 11144
rect 2247 11136 3113 11144
rect 3127 11136 3553 11144
rect 6447 11136 6713 11144
rect 6727 11136 6953 11144
rect 6967 11136 7233 11144
rect 8487 11136 8853 11144
rect 8907 11136 8953 11144
rect 9147 11136 9413 11144
rect 10096 11144 10104 11153
rect 10096 11136 10293 11144
rect 11107 11136 11193 11144
rect 3167 11116 3473 11124
rect 5807 11116 6473 11124
rect 8147 11116 8633 11124
rect 9407 11116 9853 11124
rect 9867 11116 10113 11124
rect 10827 11116 11093 11124
rect 7947 11096 8573 11104
rect 4967 11076 5013 11084
rect 747 10956 1733 10964
rect 1747 10956 1873 10964
rect 8207 10956 8373 10964
rect 707 10936 753 10944
rect 2847 10936 2913 10944
rect 4707 10936 5273 10944
rect 5287 10936 5333 10944
rect 5347 10936 5653 10944
rect 6027 10936 6053 10944
rect 6287 10936 6393 10944
rect 8127 10936 8193 10944
rect 8247 10936 8333 10944
rect 8347 10936 8413 10944
rect 9847 10936 9893 10944
rect 10647 10936 10793 10944
rect 10807 10936 10893 10944
rect 11247 10936 11293 10944
rect 207 10916 373 10924
rect 387 10916 1053 10924
rect 1427 10916 1453 10924
rect 1687 10916 1713 10924
rect 1767 10916 1893 10924
rect 2127 10916 2153 10924
rect 2427 10916 2453 10924
rect 2807 10916 2873 10924
rect 3107 10916 3133 10924
rect 3156 10907 3164 10933
rect 3207 10916 3273 10924
rect 3887 10916 3913 10924
rect 4047 10916 4073 10924
rect 4367 10916 4553 10924
rect 4947 10916 4953 10924
rect 4967 10916 5673 10924
rect 5747 10916 5973 10924
rect 5987 10916 6473 10924
rect 6767 10916 6953 10924
rect 7007 10916 7213 10924
rect 7267 10916 7433 10924
rect 7487 10916 7693 10924
rect 8227 10916 8393 10924
rect 8827 10916 9093 10924
rect 9147 10916 9173 10924
rect 9347 10916 9433 10924
rect 9447 10916 9793 10924
rect 9807 10916 9933 10924
rect 10347 10916 10633 10924
rect 10596 10907 10604 10916
rect 10996 10916 11033 10924
rect 87 10896 533 10904
rect 1167 10896 1433 10904
rect 1447 10896 1533 10904
rect 1567 10896 1773 10904
rect 2536 10896 2773 10904
rect 207 10876 673 10884
rect 947 10876 993 10884
rect 1007 10876 1173 10884
rect 1727 10876 2053 10884
rect 2227 10876 2373 10884
rect 2536 10884 2544 10896
rect 2787 10896 2853 10904
rect 2907 10896 2953 10904
rect 3176 10896 4733 10904
rect 2387 10876 2544 10884
rect 2667 10876 2833 10884
rect 3176 10884 3184 10896
rect 6067 10896 6253 10904
rect 6687 10896 7393 10904
rect 7427 10896 7493 10904
rect 7507 10896 7933 10904
rect 7947 10896 8113 10904
rect 9127 10896 9393 10904
rect 9427 10896 9613 10904
rect 9867 10896 9913 10904
rect 10107 10896 10553 10904
rect 10727 10896 10813 10904
rect 10996 10904 11004 10916
rect 11087 10916 11293 10924
rect 10827 10896 11004 10904
rect 11067 10896 11093 10904
rect 3107 10876 3184 10884
rect 3207 10876 4093 10884
rect 4587 10876 4833 10884
rect 6227 10876 6373 10884
rect 6487 10876 6973 10884
rect 7167 10876 7413 10884
rect 9147 10876 9173 10884
rect 9667 10876 9893 10884
rect 10147 10876 10193 10884
rect 10567 10876 10613 10884
rect 10627 10876 10753 10884
rect 11207 10876 11273 10884
rect 487 10856 873 10864
rect 1667 10856 1893 10864
rect 2607 10856 2633 10864
rect 2647 10856 2733 10864
rect 2867 10856 3173 10864
rect 3227 10856 3893 10864
rect 3947 10856 4173 10864
rect 4347 10856 5113 10864
rect 5787 10856 7173 10864
rect 9247 10856 9353 10864
rect 1067 10836 2073 10844
rect 2087 10836 2093 10844
rect 2107 10836 2233 10844
rect 2947 10836 3193 10844
rect 3947 10836 4333 10844
rect 4747 10836 5313 10844
rect 6047 10836 6273 10844
rect 8587 10836 8613 10844
rect 607 10816 893 10824
rect 907 10816 1333 10824
rect 1347 10816 1913 10824
rect 4067 10816 4113 10824
rect 4767 10816 4893 10824
rect 6007 10816 6493 10824
rect 9887 10816 9953 10824
rect 9967 10816 10073 10824
rect 1407 10796 1733 10804
rect 4047 10796 4073 10804
rect 4107 10796 5493 10804
rect 967 10776 1173 10784
rect 1187 10776 1433 10784
rect 1447 10776 3533 10784
rect 4827 10776 5273 10784
rect 1667 10756 1693 10764
rect 1707 10756 2213 10764
rect 2767 10756 3113 10764
rect 3847 10756 4033 10764
rect 4407 10756 4733 10764
rect 4747 10756 5293 10764
rect 5307 10756 5353 10764
rect 5367 10756 5473 10764
rect 5487 10756 5953 10764
rect 5967 10756 6233 10764
rect 6447 10756 7213 10764
rect 8367 10756 9393 10764
rect 10587 10756 10693 10764
rect 10947 10756 11073 10764
rect 247 10736 313 10744
rect 467 10736 533 10744
rect 1207 10736 1453 10744
rect 1467 10736 2153 10744
rect 2467 10736 2713 10744
rect 2727 10736 3093 10744
rect 3807 10736 3993 10744
rect 4047 10736 4513 10744
rect 4807 10736 4833 10744
rect 5567 10736 5793 10744
rect 5807 10736 6073 10744
rect 6087 10736 6253 10744
rect 6267 10736 6493 10744
rect 6516 10736 6713 10744
rect -24 10716 413 10724
rect 527 10716 633 10724
rect 927 10716 1213 10724
rect 1227 10716 1393 10724
rect 1647 10716 1693 10724
rect 1747 10716 1844 10724
rect 707 10696 913 10704
rect 1427 10696 1493 10704
rect 1836 10704 1844 10716
rect 1867 10716 1893 10724
rect 2067 10716 2133 10724
rect 2927 10716 3413 10724
rect 3816 10716 4013 10724
rect 1836 10696 2473 10704
rect 2687 10696 2813 10704
rect 2827 10696 2953 10704
rect 3416 10696 3773 10704
rect -24 10676 173 10684
rect 667 10676 713 10684
rect 1207 10676 1373 10684
rect 1676 10684 1684 10693
rect 1387 10676 1684 10684
rect 2447 10676 2533 10684
rect 2547 10676 2913 10684
rect 2927 10676 2933 10684
rect 3416 10684 3424 10696
rect 3816 10704 3824 10716
rect 4207 10716 4313 10724
rect 4327 10716 4484 10724
rect 3787 10696 3824 10704
rect 4007 10696 4233 10704
rect 4267 10696 4333 10704
rect 4476 10704 4484 10716
rect 4587 10716 4773 10724
rect 5487 10716 5553 10724
rect 5647 10716 5753 10724
rect 6047 10716 6293 10724
rect 6516 10724 6524 10736
rect 6727 10736 6793 10744
rect 7227 10736 7453 10744
rect 7507 10736 7673 10744
rect 8147 10736 8513 10744
rect 8787 10736 9073 10744
rect 9947 10736 10213 10744
rect 10467 10736 11013 10744
rect 11027 10736 11113 10744
rect 6307 10716 6524 10724
rect 6587 10716 6973 10724
rect 7847 10716 7953 10724
rect 4476 10696 4753 10704
rect 4807 10696 4833 10704
rect 4907 10696 5033 10704
rect 5236 10704 5244 10713
rect 5047 10696 5244 10704
rect 5407 10696 5513 10704
rect 5827 10696 6033 10704
rect 6327 10696 6513 10704
rect 6967 10696 7013 10704
rect 7047 10696 7093 10704
rect 7407 10696 7673 10704
rect 7856 10704 7864 10716
rect 7967 10716 8353 10724
rect 8567 10716 8733 10724
rect 8796 10716 8993 10724
rect 8796 10707 8804 10716
rect 9047 10716 9993 10724
rect 10727 10716 11144 10724
rect 7687 10696 7864 10704
rect 7887 10696 8313 10704
rect 8467 10696 8533 10704
rect 8947 10696 8973 10704
rect 8987 10696 9153 10704
rect 9267 10696 9413 10704
rect 9687 10696 10473 10704
rect 10487 10696 10633 10704
rect 2987 10676 3424 10684
rect 4247 10676 4993 10684
rect 5227 10676 5373 10684
rect 5467 10676 5533 10684
rect 5547 10676 5773 10684
rect 5787 10676 6053 10684
rect 6367 10676 7053 10684
rect 8707 10676 9013 10684
rect 9327 10676 9413 10684
rect 10656 10684 10664 10713
rect 11136 10707 11144 10716
rect 11167 10716 11293 10724
rect 10687 10696 10713 10704
rect 10767 10696 10873 10704
rect 10927 10696 11013 10704
rect 10656 10676 10813 10684
rect 527 10656 933 10664
rect 1527 10656 1713 10664
rect 3507 10656 4553 10664
rect 5267 10656 5313 10664
rect 5327 10656 6013 10664
rect 9907 10656 9933 10664
rect 9947 10656 9973 10664
rect 9987 10656 10153 10664
rect 10647 10656 11253 10664
rect 3467 10636 4473 10644
rect 4487 10636 5493 10644
rect 3887 10616 4293 10624
rect 10267 10616 10313 10624
rect 2007 10596 3233 10604
rect 3247 10596 6573 10604
rect 3207 10576 4093 10584
rect 3127 10556 3373 10564
rect 387 10536 1153 10544
rect 707 10516 2413 10524
rect 3447 10516 3573 10524
rect 3587 10516 4273 10524
rect 67 10496 733 10504
rect 1167 10496 2613 10504
rect 4127 10496 4773 10504
rect 8307 10496 8893 10504
rect 8907 10496 9733 10504
rect 1616 10476 1633 10484
rect 1616 10467 1624 10476
rect 1727 10476 1793 10484
rect 1807 10476 4853 10484
rect 6296 10476 6393 10484
rect 6296 10467 6304 10476
rect 6407 10476 6733 10484
rect 7067 10476 7513 10484
rect 7527 10476 7833 10484
rect 467 10456 673 10464
rect 1247 10456 1573 10464
rect 1887 10456 1933 10464
rect 2307 10456 2513 10464
rect 2627 10456 3313 10464
rect 3367 10456 3793 10464
rect 3867 10456 4213 10464
rect 4647 10456 4693 10464
rect 4707 10456 4713 10464
rect 5367 10456 5513 10464
rect 5567 10456 5973 10464
rect 427 10436 513 10444
rect 667 10436 693 10444
rect 716 10436 1373 10444
rect 716 10424 724 10436
rect 1467 10436 1593 10444
rect 1867 10436 1893 10444
rect 2267 10436 2333 10444
rect 2567 10436 3033 10444
rect 3127 10436 3153 10444
rect 3627 10436 3653 10444
rect 4067 10436 4584 10444
rect 627 10416 724 10424
rect 767 10416 1833 10424
rect 1887 10416 1913 10424
rect 1927 10416 1953 10424
rect 2327 10416 2393 10424
rect 2927 10416 3053 10424
rect 3076 10424 3084 10433
rect 3076 10416 3333 10424
rect 3387 10416 3593 10424
rect 4576 10424 4584 10436
rect 4607 10436 4733 10444
rect 5347 10436 5593 10444
rect 4576 10416 4873 10424
rect 5616 10424 5624 10456
rect 6347 10456 6453 10464
rect 7827 10456 8173 10464
rect 8327 10456 8373 10464
rect 9096 10456 9133 10464
rect 6107 10436 6533 10444
rect 6827 10436 7413 10444
rect 7807 10436 7873 10444
rect 7896 10436 8033 10444
rect 5507 10416 5624 10424
rect 5707 10416 6013 10424
rect 6027 10416 6353 10424
rect 6367 10416 6673 10424
rect 6907 10416 7073 10424
rect 7087 10416 7193 10424
rect 7896 10424 7904 10436
rect 8047 10436 8213 10444
rect 8367 10436 8553 10444
rect 8867 10436 8953 10444
rect 7507 10416 7904 10424
rect 8407 10416 8493 10424
rect 9096 10424 9104 10456
rect 9347 10456 9373 10464
rect 9427 10456 9453 10464
rect 9487 10456 10593 10464
rect 10927 10456 11073 10464
rect 11227 10456 11333 10464
rect 9127 10436 9213 10444
rect 9227 10436 9353 10444
rect 9407 10436 9613 10444
rect 10127 10436 10313 10444
rect 10607 10436 10733 10444
rect 9096 10416 9133 10424
rect 9607 10416 9633 10424
rect 9927 10416 9993 10424
rect 10287 10416 10353 10424
rect 10367 10416 10393 10424
rect 10627 10416 10833 10424
rect 187 10396 393 10404
rect 1407 10396 1493 10404
rect 1867 10396 1893 10404
rect 2587 10396 2673 10404
rect 3027 10396 3093 10404
rect 3147 10396 4313 10404
rect 4487 10396 4573 10404
rect 4907 10396 5113 10404
rect 5587 10396 5833 10404
rect 5987 10396 6553 10404
rect 6847 10396 7113 10404
rect 9107 10396 9173 10404
rect 9187 10396 9873 10404
rect 9907 10396 10013 10404
rect 10047 10396 10093 10404
rect 10267 10396 10333 10404
rect 907 10376 2273 10384
rect 3167 10376 3833 10384
rect 4687 10376 7313 10384
rect 7327 10376 7893 10384
rect 7907 10376 8913 10384
rect 9127 10376 9153 10384
rect 9347 10376 9573 10384
rect 9587 10376 9673 10384
rect 9687 10376 9833 10384
rect -24 10356 153 10364
rect 2087 10356 2113 10364
rect 2127 10356 2273 10364
rect 3567 10356 4093 10364
rect 5107 10356 5533 10364
rect 227 10336 633 10344
rect 647 10336 973 10344
rect 2787 10336 2993 10344
rect 3007 10336 3913 10344
rect 5907 10336 6013 10344
rect 7687 10336 7713 10344
rect 8647 10336 8733 10344
rect 10567 10336 10753 10344
rect -24 10316 733 10324
rect 2847 10316 5013 10324
rect 8587 10316 8693 10324
rect 2847 10296 3713 10304
rect 4927 10296 7093 10304
rect 10027 10296 11093 10304
rect -24 10276 193 10284
rect 407 10276 1173 10284
rect 1887 10276 2193 10284
rect 2207 10276 2733 10284
rect 3607 10276 3653 10284
rect 3667 10276 3833 10284
rect 4307 10276 4353 10284
rect 6387 10276 6513 10284
rect 6527 10276 7253 10284
rect 7887 10276 7973 10284
rect 11007 10276 11313 10284
rect 887 10256 1653 10264
rect 1667 10256 1773 10264
rect 2307 10256 2333 10264
rect 2347 10256 2533 10264
rect 2547 10256 2573 10264
rect 2587 10256 3093 10264
rect 3107 10256 3273 10264
rect 3307 10256 3373 10264
rect 3407 10256 3513 10264
rect 3587 10256 3653 10264
rect 3667 10256 3773 10264
rect 3827 10256 3873 10264
rect 4167 10256 4293 10264
rect 5587 10256 5733 10264
rect 6087 10256 6473 10264
rect 6747 10256 6893 10264
rect 7007 10256 7453 10264
rect 7707 10256 7753 10264
rect 7967 10256 8193 10264
rect 8887 10256 9093 10264
rect 10747 10256 11053 10264
rect -24 10236 13 10244
rect 287 10236 473 10244
rect 527 10236 593 10244
rect 627 10236 2333 10244
rect 2387 10236 2793 10244
rect 3327 10236 3813 10244
rect 3867 10236 4193 10244
rect 4207 10236 4213 10244
rect 4267 10236 4333 10244
rect 4347 10236 4553 10244
rect 4567 10236 4813 10244
rect 4827 10236 5593 10244
rect 5767 10236 5853 10244
rect 5867 10236 6504 10244
rect 427 10216 453 10224
rect 476 10216 764 10224
rect -24 10184 -16 10204
rect 476 10204 484 10216
rect 27 10196 484 10204
rect 547 10196 733 10204
rect 756 10204 764 10216
rect 1647 10216 1813 10224
rect 2367 10216 2553 10224
rect 2927 10216 3033 10224
rect 3316 10224 3324 10233
rect 6496 10227 6504 10236
rect 6787 10236 6953 10244
rect 7247 10236 7293 10244
rect 8027 10236 8153 10244
rect 8587 10236 8673 10244
rect 8687 10236 8853 10244
rect 8907 10236 9273 10244
rect 9687 10236 9793 10244
rect 10527 10236 11024 10244
rect 3087 10216 3324 10224
rect 3387 10216 3533 10224
rect 3587 10216 3633 10224
rect 4067 10216 4273 10224
rect 4527 10216 4753 10224
rect 4807 10216 5273 10224
rect 5747 10216 5813 10224
rect 7016 10224 7024 10233
rect 6767 10216 7073 10224
rect 7267 10216 7353 10224
rect 7367 10216 7413 10224
rect 7687 10216 7893 10224
rect 7916 10207 7924 10233
rect 11016 10227 11024 10236
rect 8187 10216 8333 10224
rect 8387 10216 8613 10224
rect 8667 10216 9473 10224
rect 9547 10216 9773 10224
rect 9827 10216 10233 10224
rect 10247 10216 10453 10224
rect 10507 10216 10673 10224
rect 756 10196 2053 10204
rect 2327 10196 2813 10204
rect 3727 10196 3833 10204
rect 3847 10196 4033 10204
rect 5047 10196 5253 10204
rect 5487 10196 5553 10204
rect 5627 10196 6673 10204
rect 8407 10196 8433 10204
rect 8447 10196 8573 10204
rect 9127 10196 9213 10204
rect 9407 10196 9513 10204
rect 9887 10196 9973 10204
rect 9987 10196 10013 10204
rect 10067 10196 10293 10204
rect 11036 10204 11044 10233
rect 11056 10227 11064 10253
rect 11076 10224 11084 10233
rect 11076 10216 11253 10224
rect 11007 10196 11044 10204
rect -24 10176 1393 10184
rect 3807 10176 4073 10184
rect 4087 10176 4253 10184
rect 4927 10176 5033 10184
rect 5107 10176 5293 10184
rect 5467 10176 5513 10184
rect 7947 10176 8353 10184
rect 8367 10176 8453 10184
rect 10787 10176 11273 10184
rect 247 10156 253 10164
rect 267 10156 613 10164
rect 2747 10156 3073 10164
rect 3927 10156 4493 10164
rect 4627 10156 5773 10164
rect 6467 10156 6873 10164
rect 7127 10156 7213 10164
rect 7227 10156 7973 10164
rect 9427 10156 10253 10164
rect 10267 10156 10313 10164
rect 6007 10136 6233 10144
rect 9027 10136 9093 10144
rect 9747 10136 9813 10144
rect 507 10116 633 10124
rect 5987 10116 6753 10124
rect 7747 10116 7853 10124
rect 1487 10056 2073 10064
rect 2087 10056 2373 10064
rect 607 10036 1173 10044
rect 1187 10036 6933 10044
rect 8907 10036 9313 10044
rect 2107 10016 2293 10024
rect 3547 10016 4873 10024
rect 4887 10016 5313 10024
rect 8827 10016 10333 10024
rect 1267 9996 1873 10004
rect 1887 9996 2313 10004
rect 3267 9996 4713 10004
rect 5667 9996 5993 10004
rect 6687 9996 7273 10004
rect 9267 9996 10753 10004
rect 10767 9996 10813 10004
rect 10827 9996 11333 10004
rect 67 9976 253 9984
rect 1027 9976 1213 9984
rect 2127 9976 2353 9984
rect 3467 9976 3993 9984
rect 4067 9976 4973 9984
rect 5327 9976 5413 9984
rect 5447 9976 5713 9984
rect 5787 9976 5933 9984
rect 6607 9976 6853 9984
rect 7347 9976 7433 9984
rect 7587 9976 7833 9984
rect 7856 9976 8113 9984
rect 607 9956 1073 9964
rect 1167 9956 1193 9964
rect 2107 9956 2313 9964
rect 2367 9956 2393 9964
rect 2747 9956 2793 9964
rect 2827 9956 2973 9964
rect 2987 9956 3033 9964
rect 3087 9956 3273 9964
rect 3427 9956 3493 9964
rect 3607 9956 3793 9964
rect 4167 9956 4253 9964
rect 4307 9956 4573 9964
rect 4687 9956 4733 9964
rect 5027 9956 5153 9964
rect 5167 9956 5193 9964
rect 5607 9956 5653 9964
rect 5707 9956 5813 9964
rect 5887 9956 6033 9964
rect 6147 9956 6593 9964
rect 6647 9956 6673 9964
rect 6907 9956 6993 9964
rect 7007 9956 7373 9964
rect 7487 9956 7613 9964
rect 7667 9956 7773 9964
rect 7856 9964 7864 9976
rect 8447 9976 9393 9984
rect 9827 9976 9853 9984
rect 10207 9976 10273 9984
rect 10387 9976 10493 9984
rect 11027 9976 11053 9984
rect 7787 9956 7864 9964
rect 8567 9956 8773 9964
rect 9007 9956 9033 9964
rect 9247 9956 9313 9964
rect 9367 9956 9373 9964
rect 9387 9956 9993 9964
rect 10167 9956 10233 9964
rect 647 9936 873 9944
rect 1476 9936 1613 9944
rect 287 9916 413 9924
rect 907 9916 933 9924
rect 1476 9924 1484 9936
rect 1667 9936 1713 9944
rect 1807 9936 1893 9944
rect 1907 9936 2033 9944
rect 2147 9936 3053 9944
rect 3067 9936 3453 9944
rect 3527 9936 3544 9944
rect 3536 9927 3544 9936
rect 3567 9936 3633 9944
rect 3667 9936 3773 9944
rect 3796 9944 3804 9953
rect 3796 9936 3993 9944
rect 4027 9936 4933 9944
rect 5476 9944 5484 9953
rect 5476 9936 5673 9944
rect 5927 9936 6313 9944
rect 6407 9936 6533 9944
rect 6667 9936 6713 9944
rect 6927 9936 6953 9944
rect 7447 9936 7593 9944
rect 7727 9936 7853 9944
rect 7876 9927 7884 9953
rect 10296 9947 10304 9973
rect 10447 9956 10533 9964
rect 11176 9956 11293 9964
rect 8607 9936 8833 9944
rect 8947 9936 9053 9944
rect 9107 9936 9293 9944
rect 10527 9936 10813 9944
rect 10827 9936 10973 9944
rect 11176 9944 11184 9956
rect 11047 9936 11184 9944
rect 11207 9936 11273 9944
rect 1387 9916 1484 9924
rect 1507 9916 1633 9924
rect 1887 9916 1913 9924
rect 3007 9916 3393 9924
rect 3487 9916 3513 9924
rect 4567 9916 4953 9924
rect 6627 9916 6873 9924
rect 7807 9916 7833 9924
rect 9047 9916 9073 9924
rect 9087 9916 9153 9924
rect 10047 9916 10253 9924
rect 10787 9916 10933 9924
rect 10947 9916 11253 9924
rect 927 9896 1393 9904
rect 1407 9896 3593 9904
rect 7427 9896 7813 9904
rect 7827 9896 7953 9904
rect 8427 9896 9473 9904
rect 11227 9896 11333 9904
rect 227 9876 553 9884
rect 567 9876 1853 9884
rect 3907 9876 4673 9884
rect 7787 9876 7873 9884
rect 327 9856 353 9864
rect 1627 9856 1833 9864
rect 2387 9856 2633 9864
rect 2827 9856 3833 9864
rect 7887 9856 7973 9864
rect 7987 9856 8093 9864
rect 687 9836 693 9844
rect 707 9836 1233 9844
rect 1987 9836 2813 9844
rect 2827 9836 2853 9844
rect 2867 9836 3633 9844
rect 5027 9836 5293 9844
rect 6127 9836 8013 9844
rect 8267 9836 9013 9844
rect 3867 9816 4213 9824
rect 4567 9816 5253 9824
rect 6167 9816 6313 9824
rect 6687 9816 7573 9824
rect 1087 9796 1113 9804
rect 1127 9796 1353 9804
rect 1407 9796 3193 9804
rect 3207 9796 3593 9804
rect 3847 9796 4493 9804
rect 5467 9796 5513 9804
rect 6587 9796 7053 9804
rect 1107 9776 1353 9784
rect 1667 9776 1753 9784
rect 2127 9776 2333 9784
rect 3287 9776 3533 9784
rect 3567 9776 3693 9784
rect 3747 9776 3793 9784
rect 4847 9776 4893 9784
rect 5267 9776 5373 9784
rect 5587 9776 5833 9784
rect 6067 9776 6353 9784
rect 6927 9776 7013 9784
rect 8607 9776 8793 9784
rect 9247 9776 9293 9784
rect 9307 9776 9413 9784
rect 9847 9776 9893 9784
rect 10027 9776 10153 9784
rect 10987 9776 11093 9784
rect 727 9756 913 9764
rect 927 9756 1113 9764
rect 1167 9756 1813 9764
rect 1927 9756 1993 9764
rect 2667 9756 2853 9764
rect 2907 9756 3013 9764
rect 4027 9756 4073 9764
rect 4227 9756 4513 9764
rect 4687 9756 4753 9764
rect 4807 9756 4993 9764
rect 5087 9756 5293 9764
rect 5827 9756 5944 9764
rect 167 9736 193 9744
rect 887 9736 904 9744
rect 436 9707 444 9733
rect 467 9716 553 9724
rect 896 9707 904 9736
rect 1147 9736 1253 9744
rect 1427 9736 1433 9744
rect 1447 9736 1673 9744
rect 1687 9736 1973 9744
rect 2387 9736 3033 9744
rect 3047 9736 3053 9744
rect 3547 9736 3733 9744
rect 4267 9736 4293 9744
rect 4507 9736 4653 9744
rect 4827 9736 5173 9744
rect 5367 9736 5513 9744
rect 5936 9744 5944 9756
rect 5967 9756 5993 9764
rect 6047 9756 6273 9764
rect 6667 9756 6753 9764
rect 6807 9756 7084 9764
rect 7076 9747 7084 9756
rect 7547 9756 7633 9764
rect 7647 9756 7753 9764
rect 8307 9756 8353 9764
rect 9667 9756 9924 9764
rect 9916 9747 9924 9756
rect 10067 9756 10473 9764
rect 10487 9756 10664 9764
rect 10656 9747 10664 9756
rect 5936 9736 6293 9744
rect 6347 9736 6553 9744
rect 7127 9736 7293 9744
rect 7307 9736 7513 9744
rect 7907 9736 7993 9744
rect 8227 9736 8413 9744
rect 8827 9736 8973 9744
rect 8987 9736 9193 9744
rect 9247 9736 9433 9744
rect 9527 9736 9633 9744
rect 9647 9736 9804 9744
rect 1387 9716 1473 9724
rect 1707 9716 1893 9724
rect 2627 9716 2653 9724
rect 2807 9716 2873 9724
rect 3627 9716 3773 9724
rect 4207 9716 4233 9724
rect 4287 9716 4313 9724
rect 5007 9716 5033 9724
rect 5287 9716 5653 9724
rect 5707 9716 5713 9724
rect 5727 9716 5793 9724
rect 5807 9716 5953 9724
rect 7047 9716 7133 9724
rect 9227 9716 9273 9724
rect 9796 9724 9804 9736
rect 10187 9736 10413 9744
rect 10467 9736 10493 9744
rect 10687 9736 10713 9744
rect 10727 9736 10893 9744
rect 11067 9736 11113 9744
rect 9796 9716 9973 9724
rect 9987 9716 10133 9724
rect 3687 9696 4013 9704
rect 6327 9696 8333 9704
rect 8347 9696 8453 9704
rect 9727 9696 9873 9704
rect 9887 9696 9993 9704
rect 5147 9676 5953 9684
rect 5967 9676 6453 9684
rect 7527 9676 7733 9684
rect 7747 9676 7853 9684
rect 8767 9676 9853 9684
rect 9987 9676 10053 9684
rect 2987 9656 3033 9664
rect 3267 9656 3293 9664
rect 3636 9656 4053 9664
rect 187 9636 233 9644
rect 247 9636 413 9644
rect 427 9636 473 9644
rect 487 9636 853 9644
rect 867 9636 953 9644
rect 967 9636 2393 9644
rect 2407 9636 3093 9644
rect 3636 9644 3644 9656
rect 4447 9656 4533 9664
rect 4547 9656 5273 9664
rect 5787 9656 6013 9664
rect 6027 9656 6453 9664
rect 8207 9656 8873 9664
rect 9167 9656 10173 9664
rect 3107 9636 3644 9644
rect 3887 9636 4533 9644
rect 7967 9636 8233 9644
rect 8647 9636 9673 9644
rect 9687 9636 9833 9644
rect 3647 9616 3773 9624
rect 9187 9616 10453 9624
rect 2847 9596 4213 9604
rect 7147 9596 7553 9604
rect 7327 9576 7353 9584
rect 1647 9556 2673 9564
rect 2647 9536 3073 9544
rect 10147 9536 10613 9544
rect 10627 9536 10693 9544
rect 1467 9516 2253 9524
rect 3067 9516 4333 9524
rect 5607 9516 6713 9524
rect 6727 9516 6773 9524
rect 8087 9516 8933 9524
rect 8947 9516 9313 9524
rect 9327 9516 9333 9524
rect 10347 9516 10993 9524
rect 1387 9496 1593 9504
rect 1887 9496 2153 9504
rect 2167 9496 2413 9504
rect 2807 9496 3233 9504
rect 3247 9496 3413 9504
rect 3447 9496 3473 9504
rect 3707 9496 3733 9504
rect 3756 9496 4573 9504
rect 167 9476 193 9484
rect 527 9476 693 9484
rect 707 9476 853 9484
rect 976 9476 1173 9484
rect 976 9467 984 9476
rect 1187 9476 1333 9484
rect 1427 9476 1453 9484
rect 1607 9476 1633 9484
rect 1656 9467 1664 9493
rect 1927 9476 1973 9484
rect 2207 9476 2233 9484
rect 2407 9476 2433 9484
rect 2487 9476 2513 9484
rect 2527 9476 3413 9484
rect 3756 9484 3764 9496
rect 4587 9496 4813 9504
rect 5647 9496 6213 9504
rect 6227 9496 6413 9504
rect 6507 9496 6573 9504
rect 7067 9496 7453 9504
rect 7467 9496 7513 9504
rect 8287 9496 8813 9504
rect 10707 9496 10813 9504
rect 3467 9476 3764 9484
rect 4067 9476 4113 9484
rect 4387 9476 4413 9484
rect 4567 9476 4613 9484
rect 4787 9476 4833 9484
rect 5007 9476 5073 9484
rect 5116 9476 5433 9484
rect 267 9456 673 9464
rect 1407 9456 1473 9464
rect 1687 9456 1893 9464
rect 2087 9456 2133 9464
rect 2187 9456 2253 9464
rect 2467 9456 2573 9464
rect 2727 9456 3173 9464
rect 3347 9456 3433 9464
rect 3587 9456 3673 9464
rect 4147 9456 4193 9464
rect 4307 9456 4393 9464
rect 4647 9456 4913 9464
rect 5116 9464 5124 9476
rect 5867 9476 6013 9484
rect 6067 9476 6093 9484
rect 6107 9476 6133 9484
rect 6767 9476 6953 9484
rect 6967 9476 7033 9484
rect 7427 9476 7493 9484
rect 7507 9476 7553 9484
rect 7947 9476 8013 9484
rect 8167 9476 8364 9484
rect 5067 9456 5124 9464
rect 5147 9456 5293 9464
rect 5516 9464 5524 9473
rect 8356 9467 8364 9476
rect 9007 9476 9093 9484
rect 9367 9476 9513 9484
rect 9807 9476 9873 9484
rect 10087 9476 10513 9484
rect 10647 9476 10773 9484
rect 10787 9476 11033 9484
rect 5307 9456 5524 9464
rect 5567 9456 5684 9464
rect 867 9436 1313 9444
rect 1327 9436 1613 9444
rect 1647 9436 1833 9444
rect 1947 9436 2213 9444
rect 2227 9436 2793 9444
rect 2967 9436 3153 9444
rect 3967 9436 4093 9444
rect 4367 9436 4593 9444
rect 5327 9436 5593 9444
rect 5676 9444 5684 9456
rect 5827 9456 5993 9464
rect 6427 9456 6653 9464
rect 6667 9456 6693 9464
rect 6747 9456 6913 9464
rect 7127 9456 7573 9464
rect 7587 9456 7853 9464
rect 7867 9456 8213 9464
rect 8627 9456 8673 9464
rect 8847 9456 9053 9464
rect 9287 9456 9333 9464
rect 10107 9456 10313 9464
rect 10547 9456 10593 9464
rect 10607 9456 10753 9464
rect 5676 9436 6033 9444
rect 6047 9436 6233 9444
rect 6247 9436 6613 9444
rect 8607 9436 8773 9444
rect 8807 9436 8933 9444
rect 9307 9436 9373 9444
rect 9687 9436 10053 9444
rect 10107 9436 10173 9444
rect 10367 9436 11053 9444
rect 11067 9436 11113 9444
rect 11127 9436 11253 9444
rect 1207 9416 2073 9424
rect 2427 9416 2493 9424
rect 2507 9416 3393 9424
rect 4427 9416 4733 9424
rect 4867 9416 6453 9424
rect 6647 9416 6673 9424
rect 8407 9416 8793 9424
rect 9427 9416 10033 9424
rect 10207 9416 10833 9424
rect 10847 9416 10933 9424
rect 10947 9416 11213 9424
rect 2667 9396 2913 9404
rect 3167 9396 3913 9404
rect 3927 9396 4053 9404
rect 5527 9396 5613 9404
rect 6527 9396 6733 9404
rect 8807 9396 8893 9404
rect 2967 9376 3013 9384
rect 3407 9376 3493 9384
rect 3507 9376 4893 9384
rect 5807 9376 5973 9384
rect 6487 9376 6513 9384
rect 6687 9376 6833 9384
rect 7807 9376 7833 9384
rect 887 9356 933 9364
rect 4227 9356 4333 9364
rect 4347 9356 6433 9364
rect 6467 9356 7553 9364
rect 7567 9356 9453 9364
rect 707 9336 713 9344
rect 727 9336 1813 9344
rect 1827 9336 1853 9344
rect 3207 9336 3213 9344
rect 3227 9336 4853 9344
rect 7007 9336 7033 9344
rect 7767 9336 7913 9344
rect 8547 9336 8833 9344
rect 8927 9336 8953 9344
rect 487 9316 633 9324
rect 647 9316 2393 9324
rect 3147 9316 3833 9324
rect 4107 9316 4473 9324
rect 9347 9316 9713 9324
rect 667 9296 853 9304
rect 1387 9296 1613 9304
rect 1667 9296 1873 9304
rect 2587 9296 2613 9304
rect 2627 9296 2853 9304
rect 3407 9296 3873 9304
rect 3887 9296 4113 9304
rect 4487 9296 4793 9304
rect 4807 9296 4953 9304
rect 5547 9296 5733 9304
rect 6747 9296 6993 9304
rect 7007 9296 7193 9304
rect 7227 9296 7373 9304
rect 8227 9296 8453 9304
rect 9507 9296 9633 9304
rect 9947 9296 10213 9304
rect 10907 9296 11173 9304
rect 11187 9296 11273 9304
rect 687 9276 2353 9284
rect 2427 9276 2533 9284
rect 3027 9276 3113 9284
rect 3167 9276 3373 9284
rect 3687 9276 3893 9284
rect 3907 9276 4184 9284
rect 387 9256 593 9264
rect 1147 9256 1193 9264
rect 1407 9256 1733 9264
rect 1907 9256 2113 9264
rect 2127 9256 2193 9264
rect 2387 9256 2573 9264
rect 2607 9256 2673 9264
rect 2827 9256 2893 9264
rect 3067 9256 3133 9264
rect 3636 9264 3644 9273
rect 3636 9256 3793 9264
rect 3847 9256 4153 9264
rect 4176 9264 4184 9276
rect 4207 9276 4233 9284
rect 4267 9276 4373 9284
rect 4407 9276 4453 9284
rect 4467 9276 4793 9284
rect 5507 9276 5613 9284
rect 5936 9276 6213 9284
rect 4176 9256 4213 9264
rect 4527 9256 5173 9264
rect 5227 9256 5253 9264
rect 5487 9256 5573 9264
rect 5916 9264 5924 9273
rect 5936 9267 5944 9276
rect 6507 9276 6713 9284
rect 7187 9276 7453 9284
rect 7507 9276 7713 9284
rect 8427 9276 8473 9284
rect 8527 9276 8784 9284
rect 8776 9267 8784 9276
rect 8847 9276 9133 9284
rect 9147 9276 9293 9284
rect 9307 9276 9333 9284
rect 9707 9276 10153 9284
rect 10467 9276 10513 9284
rect 10527 9276 10613 9284
rect 10767 9276 10913 9284
rect 11067 9276 11153 9284
rect 5727 9256 5924 9264
rect 6247 9256 6333 9264
rect 6927 9256 6953 9264
rect 7387 9256 7473 9264
rect 8307 9256 8393 9264
rect 9087 9256 9233 9264
rect 9287 9256 9473 9264
rect 9607 9256 9673 9264
rect 10087 9256 10173 9264
rect 10367 9256 10373 9264
rect 10387 9256 10413 9264
rect 11007 9256 11133 9264
rect 2687 9236 2913 9244
rect 3427 9236 3613 9244
rect 3807 9236 4233 9244
rect 4507 9236 4553 9244
rect 4707 9236 5133 9244
rect 5147 9236 5193 9244
rect 5247 9236 5333 9244
rect 5767 9236 6293 9244
rect 6307 9236 6393 9244
rect 6827 9236 6973 9244
rect 7027 9236 7733 9244
rect 7747 9236 7873 9244
rect 8387 9236 8493 9244
rect 8587 9236 9053 9244
rect 9067 9236 9113 9244
rect 9127 9236 9693 9244
rect 9707 9236 9913 9244
rect 10007 9236 10393 9244
rect 10407 9236 10633 9244
rect 10707 9236 10873 9244
rect 1327 9216 1353 9224
rect 2887 9216 2993 9224
rect 3347 9216 3633 9224
rect 4767 9216 5253 9224
rect 5587 9216 6173 9224
rect 6187 9216 6753 9224
rect 6767 9216 7133 9224
rect 7407 9216 7693 9224
rect 9867 9216 9933 9224
rect 10867 9216 10893 9224
rect 2307 9196 2933 9204
rect 2947 9196 4613 9204
rect 4967 9196 5553 9204
rect 5567 9196 5633 9204
rect 5787 9196 5973 9204
rect 47 9176 53 9184
rect 67 9176 273 9184
rect 287 9176 713 9184
rect 2447 9176 4393 9184
rect 4947 9176 6473 9184
rect 6847 9176 7433 9184
rect 8427 9176 9013 9184
rect 4907 9156 5933 9164
rect 6007 9156 6433 9164
rect 6447 9156 7713 9164
rect 8787 9156 8813 9164
rect 4127 9136 6533 9144
rect 1807 9116 1833 9124
rect 1867 9116 1913 9124
rect 1927 9116 3873 9124
rect 3887 9116 4973 9124
rect 4987 9116 5173 9124
rect 5287 9116 5293 9124
rect 5307 9116 5393 9124
rect 5407 9116 5993 9124
rect 6427 9116 6913 9124
rect 587 9096 773 9104
rect 1827 9096 1853 9104
rect 2927 9096 3173 9104
rect 3187 9096 4073 9104
rect 4087 9096 7693 9104
rect 8487 9096 8573 9104
rect 4547 9076 6093 9084
rect 6107 9076 6273 9084
rect 6527 9076 7013 9084
rect 7027 9076 7253 9084
rect 7887 9076 8233 9084
rect 8547 9076 9633 9084
rect 3727 9056 5953 9064
rect 6227 9056 9353 9064
rect 9367 9056 9893 9064
rect 9907 9056 10153 9064
rect 10167 9056 10313 9064
rect 2827 9036 2844 9044
rect 2836 9027 2844 9036
rect 3467 9036 3493 9044
rect 3707 9036 3813 9044
rect 3927 9036 4033 9044
rect 4047 9036 5753 9044
rect 5867 9036 6033 9044
rect 6407 9036 6613 9044
rect 6687 9036 6973 9044
rect 7167 9036 7653 9044
rect 7667 9036 7933 9044
rect 7947 9036 8073 9044
rect 8187 9036 8273 9044
rect 8287 9036 8633 9044
rect 967 9016 1113 9024
rect 1907 9016 2133 9024
rect 2147 9016 2353 9024
rect 2367 9016 2493 9024
rect 3007 9016 3053 9024
rect 3167 9016 3213 9024
rect 3227 9016 3293 9024
rect 4767 9016 4824 9024
rect -24 8984 -16 9004
rect 167 8996 313 9004
rect 927 8996 1073 9004
rect 1287 8996 1393 9004
rect 1447 8996 1493 9004
rect 1667 8996 1693 9004
rect 2167 8996 2233 9004
rect 2387 8996 2573 9004
rect 2667 8996 2853 9004
rect 3207 8996 3613 9004
rect 3847 8996 4053 9004
rect 4727 8996 4793 9004
rect 4816 9004 4824 9016
rect 5047 9016 5113 9024
rect 5387 9016 5733 9024
rect 5747 9016 5873 9024
rect 5947 9016 7993 9024
rect 8347 9016 8513 9024
rect 10207 9016 10353 9024
rect 10807 9016 10993 9024
rect 11007 9016 11133 9024
rect 4816 8996 4833 9004
rect 5087 8996 5133 9004
rect 5607 8996 5613 9004
rect 5627 8996 5813 9004
rect 5967 8996 7113 9004
rect 7147 8996 7353 9004
rect 8096 9004 8104 9013
rect 7867 8996 8104 9004
rect 8127 8996 8193 9004
rect 8567 8996 8593 9004
rect 8887 8996 9073 9004
rect 9167 8996 9193 9004
rect 9727 8996 9853 9004
rect 10356 8996 10393 9004
rect -24 8976 193 8984
rect 436 8967 444 8993
rect 627 8976 1033 8984
rect 1167 8976 1373 8984
rect 1547 8976 1633 8984
rect 1747 8976 2093 8984
rect 2627 8976 2813 8984
rect 4327 8976 4433 8984
rect 4527 8976 4693 8984
rect 4707 8976 4773 8984
rect 4827 8976 4953 8984
rect 5316 8984 5324 8993
rect 5067 8976 5324 8984
rect 5487 8976 5533 8984
rect 5667 8976 5853 8984
rect 6167 8976 6373 8984
rect 6387 8976 6393 8984
rect 6447 8976 6513 8984
rect 6627 8976 6813 8984
rect 6827 8976 6853 8984
rect 6947 8976 7093 8984
rect 7396 8984 7404 8993
rect 7267 8976 7404 8984
rect 7827 8976 7893 8984
rect 8127 8976 8253 8984
rect 8287 8976 8393 8984
rect 8527 8976 8573 8984
rect 8627 8976 8733 8984
rect 8927 8976 9093 8984
rect 9387 8976 9573 8984
rect 9627 8976 9833 8984
rect 9887 8976 10073 8984
rect 10356 8984 10364 8996
rect 10627 8996 10833 9004
rect 10147 8976 10364 8984
rect 10387 8976 10693 8984
rect 10867 8976 11153 8984
rect 11167 8976 11173 8984
rect 11187 8976 11273 8984
rect 1487 8956 1933 8964
rect 3307 8956 3733 8964
rect 3747 8956 4293 8964
rect 4307 8956 4553 8964
rect 4807 8956 5013 8964
rect 5327 8956 5413 8964
rect 6207 8956 6813 8964
rect 7027 8956 7073 8964
rect 7427 8956 8033 8964
rect 8367 8956 9313 8964
rect 9327 8956 9373 8964
rect 9547 8956 9973 8964
rect 9987 8956 10173 8964
rect 10567 8956 10593 8964
rect 1167 8936 1673 8944
rect 2207 8936 2444 8944
rect 1227 8916 2373 8924
rect 2436 8924 2444 8936
rect 3647 8936 3853 8944
rect 3867 8936 4513 8944
rect 4587 8936 5573 8944
rect 6887 8936 7333 8944
rect 7607 8936 8353 8944
rect 8387 8936 8413 8944
rect 8427 8936 8513 8944
rect 8567 8936 8893 8944
rect 2436 8916 6333 8924
rect 7027 8916 8433 8924
rect 747 8896 893 8904
rect 907 8896 2773 8904
rect 3827 8896 3853 8904
rect 5947 8896 6133 8904
rect 6527 8896 6653 8904
rect 6907 8896 8973 8904
rect 1427 8876 3733 8884
rect 4387 8876 7773 8884
rect 8367 8876 8813 8884
rect 9267 8876 10293 8884
rect 10327 8876 10873 8884
rect 10887 8876 11093 8884
rect 247 8856 2553 8864
rect 2607 8856 4073 8864
rect 4287 8856 4433 8864
rect 4447 8856 5093 8864
rect 5227 8856 5773 8864
rect 6827 8856 7193 8864
rect 8167 8856 8393 8864
rect 8607 8856 8633 8864
rect 8667 8856 9873 8864
rect 9887 8856 9913 8864
rect 2147 8836 2153 8844
rect 2167 8836 2253 8844
rect 2267 8836 2913 8844
rect 3167 8836 3313 8844
rect 3647 8836 3933 8844
rect 4127 8836 4253 8844
rect 4267 8836 5373 8844
rect 6167 8836 6453 8844
rect 6467 8836 6593 8844
rect 6747 8836 7173 8844
rect 9627 8836 10113 8844
rect 267 8816 333 8824
rect 347 8816 1133 8824
rect 1907 8816 3313 8824
rect 3427 8816 3553 8824
rect 3567 8816 3673 8824
rect 4767 8816 4813 8824
rect 5987 8816 6273 8824
rect 6447 8816 6493 8824
rect 6607 8816 6833 8824
rect 6847 8816 7093 8824
rect 7127 8816 7213 8824
rect 8587 8816 9133 8824
rect 10367 8816 10773 8824
rect 10787 8816 10813 8824
rect 11047 8816 11113 8824
rect 727 8796 913 8804
rect 1387 8796 1613 8804
rect 1667 8796 1873 8804
rect 1896 8796 2113 8804
rect 176 8776 213 8784
rect 176 8747 184 8776
rect 707 8776 733 8784
rect 947 8776 1253 8784
rect 1327 8776 1353 8784
rect 1896 8784 1904 8796
rect 2427 8796 2473 8804
rect 2827 8796 2873 8804
rect 4487 8796 4573 8804
rect 4927 8796 5253 8804
rect 5427 8796 5433 8804
rect 5447 8796 5713 8804
rect 5907 8796 5993 8804
rect 6947 8796 7033 8804
rect 7207 8796 7253 8804
rect 1407 8776 1904 8784
rect 1987 8776 2173 8784
rect 2367 8776 2453 8784
rect 2567 8776 2993 8784
rect 3087 8776 3133 8784
rect 3196 8784 3204 8793
rect 8356 8787 8364 8813
rect 8467 8796 8753 8804
rect 8767 8796 8793 8804
rect 8867 8796 9093 8804
rect 9227 8796 9533 8804
rect 9587 8796 9753 8804
rect 9847 8796 9993 8804
rect 10087 8796 10273 8804
rect 10287 8796 10573 8804
rect 10667 8796 10813 8804
rect 10867 8796 11053 8804
rect 3196 8776 3273 8784
rect 3287 8776 3393 8784
rect 3727 8776 4053 8784
rect 4067 8776 4333 8784
rect 4567 8776 4833 8784
rect 4987 8776 5193 8784
rect 5247 8776 5593 8784
rect 5607 8776 5613 8784
rect 5627 8776 5693 8784
rect 5767 8776 5913 8784
rect 6567 8776 7033 8784
rect 7047 8776 7573 8784
rect 7647 8776 8133 8784
rect 8147 8776 8333 8784
rect 8387 8776 8473 8784
rect 8627 8776 8813 8784
rect 8907 8776 9073 8784
rect 9127 8776 9193 8784
rect 9207 8776 9313 8784
rect 9567 8776 9853 8784
rect 10036 8784 10044 8793
rect 9867 8776 10044 8784
rect 10067 8776 10193 8784
rect 10587 8776 10793 8784
rect 11107 8776 11253 8784
rect 907 8756 953 8764
rect 1147 8756 1313 8764
rect 1327 8756 1753 8764
rect 1867 8756 1913 8764
rect 2587 8756 2633 8764
rect 3467 8756 3613 8764
rect 1936 8736 2393 8744
rect 1936 8724 1944 8736
rect 2407 8736 3293 8744
rect 3636 8744 3644 8773
rect 3667 8756 3673 8764
rect 3687 8756 3873 8764
rect 4107 8756 4313 8764
rect 4516 8764 4524 8773
rect 4516 8756 4553 8764
rect 4607 8756 4733 8764
rect 5107 8756 6493 8764
rect 6767 8756 6893 8764
rect 6907 8756 7053 8764
rect 7067 8756 7233 8764
rect 7887 8756 8073 8764
rect 8187 8756 8553 8764
rect 8607 8756 9173 8764
rect 9187 8756 9293 8764
rect 9347 8756 9373 8764
rect 9767 8756 10113 8764
rect 10547 8756 10633 8764
rect 10847 8756 11113 8764
rect 11127 8756 11293 8764
rect 3627 8736 3644 8744
rect 3847 8736 4353 8744
rect 4847 8736 5693 8744
rect 6427 8736 6593 8744
rect 6756 8736 7133 8744
rect 1707 8716 1944 8724
rect 2287 8716 2573 8724
rect 3907 8716 4673 8724
rect 4767 8716 6313 8724
rect 6756 8724 6764 8736
rect 8707 8736 9033 8744
rect 9087 8736 10013 8744
rect 6416 8716 6764 8724
rect 6416 8704 6424 8716
rect 8047 8716 9253 8724
rect 6207 8696 6424 8704
rect 6447 8696 8593 8704
rect 8907 8696 9713 8704
rect 9727 8696 9813 8704
rect 3127 8676 3173 8684
rect 3187 8676 3633 8684
rect 3747 8676 5753 8684
rect 6327 8676 7533 8684
rect 7587 8676 9833 8684
rect 9847 8676 9953 8684
rect 2187 8656 2273 8664
rect 3147 8656 3153 8664
rect 5187 8656 8493 8664
rect 8607 8656 8653 8664
rect 1367 8636 2393 8644
rect 2407 8636 4333 8644
rect 4567 8636 5053 8644
rect 5867 8636 8233 8644
rect 5507 8616 7273 8624
rect 7527 8616 7673 8624
rect 7967 8616 8453 8624
rect 1687 8596 2953 8604
rect 2967 8596 4113 8604
rect 4307 8596 4513 8604
rect 4687 8596 5353 8604
rect 7667 8596 8033 8604
rect 2087 8576 2433 8584
rect 2447 8576 3013 8584
rect 3027 8576 3833 8584
rect 4347 8576 5113 8584
rect 5587 8576 7233 8584
rect 8107 8576 8173 8584
rect 8487 8576 9353 8584
rect 9507 8576 10053 8584
rect 207 8556 233 8564
rect 247 8556 673 8564
rect 687 8556 953 8564
rect 2627 8556 4773 8564
rect 4827 8556 5213 8564
rect 5647 8556 5713 8564
rect 5767 8556 6113 8564
rect 6307 8556 9553 8564
rect 1167 8536 1593 8544
rect 1607 8536 1753 8544
rect 1847 8536 1933 8544
rect 2767 8536 3453 8544
rect 3587 8536 3813 8544
rect 3827 8536 3973 8544
rect 4807 8536 4873 8544
rect 4987 8536 5493 8544
rect 5687 8536 5853 8544
rect 5867 8536 5973 8544
rect 6087 8536 6173 8544
rect 6187 8536 6213 8544
rect 6227 8536 7173 8544
rect 7327 8536 7613 8544
rect 7627 8536 7873 8544
rect 8176 8536 8533 8544
rect 707 8516 913 8524
rect 1176 8516 1273 8524
rect 1176 8507 1184 8516
rect 1447 8516 1573 8524
rect 3047 8516 3093 8524
rect 3107 8516 3133 8524
rect 3327 8516 4033 8524
rect 4087 8516 4193 8524
rect 4307 8516 4553 8524
rect 4787 8516 4813 8524
rect 4867 8516 4953 8524
rect 5407 8516 5433 8524
rect 5647 8516 5824 8524
rect 287 8496 453 8504
rect 1207 8496 1413 8504
rect 1667 8496 1913 8504
rect 1956 8496 2813 8504
rect 1956 8484 1964 8496
rect 3007 8496 3073 8504
rect 3127 8496 3753 8504
rect 3867 8496 4304 8504
rect 507 8476 1964 8484
rect 1987 8476 2173 8484
rect 3067 8476 3093 8484
rect 3327 8476 3793 8484
rect 4296 8484 4304 8496
rect 4367 8496 4413 8504
rect 4587 8496 4933 8504
rect 5027 8496 5093 8504
rect 5147 8496 5233 8504
rect 5627 8496 5793 8504
rect 5816 8504 5824 8516
rect 5907 8516 6013 8524
rect 6127 8516 6193 8524
rect 6407 8516 6573 8524
rect 6587 8516 6653 8524
rect 6727 8516 6893 8524
rect 7007 8516 7324 8524
rect 5816 8496 5833 8504
rect 6107 8496 6293 8504
rect 6327 8496 6373 8504
rect 6427 8496 6453 8504
rect 6567 8496 6673 8504
rect 6687 8496 6793 8504
rect 6827 8496 7013 8504
rect 7107 8496 7193 8504
rect 7316 8504 7324 8516
rect 7347 8516 7433 8524
rect 7547 8516 7653 8524
rect 7867 8516 7913 8524
rect 8176 8507 8184 8536
rect 8667 8536 8773 8544
rect 8787 8536 9124 8544
rect 9116 8527 9124 8536
rect 9367 8536 9533 8544
rect 8207 8516 8253 8524
rect 8407 8516 8644 8524
rect 7316 8496 7393 8504
rect 7427 8496 7573 8504
rect 7687 8496 8153 8504
rect 8227 8496 8373 8504
rect 8427 8496 8513 8504
rect 8636 8504 8644 8516
rect 8867 8516 9073 8524
rect 9776 8524 9784 8553
rect 9807 8536 10033 8544
rect 10267 8536 10533 8544
rect 10547 8536 10593 8544
rect 10927 8536 11013 8544
rect 11307 8536 11353 8544
rect 9776 8516 9813 8524
rect 10007 8516 10293 8524
rect 10407 8516 10813 8524
rect 8636 8496 8873 8504
rect 8947 8496 9053 8504
rect 9107 8496 9293 8504
rect 9387 8496 9513 8504
rect 9587 8496 9773 8504
rect 9867 8496 10013 8504
rect 10067 8496 10273 8504
rect 10327 8496 10353 8504
rect 10587 8496 10773 8504
rect 4296 8476 4693 8484
rect 4847 8476 5273 8484
rect 5367 8476 5513 8484
rect 5567 8476 5593 8484
rect 5647 8476 5873 8484
rect 5887 8476 5953 8484
rect 5987 8476 6453 8484
rect 6507 8476 6873 8484
rect 6927 8476 6993 8484
rect 7027 8476 7113 8484
rect 7167 8476 8273 8484
rect 9147 8476 9613 8484
rect 9667 8476 10333 8484
rect 10387 8476 10493 8484
rect 10507 8476 10613 8484
rect 1687 8456 1733 8464
rect 1787 8456 2813 8464
rect 2867 8456 3193 8464
rect 3847 8456 4293 8464
rect 4327 8456 4673 8464
rect 4847 8456 5853 8464
rect 5927 8456 5993 8464
rect 6107 8456 6433 8464
rect 6647 8456 7264 8464
rect 1587 8436 2193 8444
rect 2207 8436 2593 8444
rect 4067 8436 4993 8444
rect 5127 8436 6733 8444
rect 6807 8436 6913 8444
rect 7256 8444 7264 8456
rect 7287 8456 7633 8464
rect 7647 8456 7733 8464
rect 8447 8456 9393 8464
rect 9547 8456 10033 8464
rect 10047 8456 10073 8464
rect 7256 8436 7853 8444
rect 9847 8436 10553 8444
rect 267 8416 673 8424
rect 687 8416 1133 8424
rect 1147 8416 1553 8424
rect 3627 8416 6793 8424
rect 6887 8416 7093 8424
rect 7607 8416 7633 8424
rect 887 8396 933 8404
rect 987 8396 1373 8404
rect 1387 8396 1653 8404
rect 1767 8396 2353 8404
rect 2647 8396 3924 8404
rect 1607 8376 2293 8384
rect 2607 8376 3733 8384
rect 3916 8384 3924 8396
rect 4347 8396 4933 8404
rect 5027 8396 5573 8404
rect 6336 8396 6553 8404
rect 3916 8376 4053 8384
rect 4307 8376 5473 8384
rect 5487 8376 5633 8384
rect 6336 8384 6344 8396
rect 6607 8396 7073 8404
rect 7127 8396 7573 8404
rect 7627 8396 8633 8404
rect 6047 8376 6344 8384
rect 6367 8376 7593 8384
rect 7607 8376 8213 8384
rect 8227 8376 8833 8384
rect 9307 8376 9433 8384
rect 2167 8356 2433 8364
rect 2447 8356 2893 8364
rect 2907 8356 4313 8364
rect 4327 8356 4493 8364
rect 4527 8356 4873 8364
rect 4887 8356 4913 8364
rect 5087 8356 5573 8364
rect 5836 8356 6053 8364
rect 487 8336 633 8344
rect 647 8336 1093 8344
rect 1167 8336 1333 8344
rect 1347 8336 1773 8344
rect 1807 8336 2073 8344
rect 2367 8336 3253 8344
rect 3767 8336 4113 8344
rect 4127 8336 5173 8344
rect 5836 8344 5844 8356
rect 6147 8356 6293 8364
rect 6307 8356 6913 8364
rect 6927 8356 6933 8364
rect 7107 8356 7293 8364
rect 8207 8356 8593 8364
rect 8727 8356 10373 8364
rect 10507 8356 11033 8364
rect 11307 8356 11404 8364
rect 5187 8336 5844 8344
rect 5867 8336 6553 8344
rect 6647 8336 6673 8344
rect 6767 8336 6813 8344
rect 6827 8336 6833 8344
rect 6887 8336 7353 8344
rect 7387 8336 7613 8344
rect 7687 8336 8113 8344
rect 8407 8336 9333 8344
rect 10067 8336 10393 8344
rect 10567 8336 10813 8344
rect 387 8316 593 8324
rect 607 8316 1053 8324
rect 1467 8316 1873 8324
rect 1887 8316 1933 8324
rect 2127 8316 2493 8324
rect 2847 8316 3033 8324
rect 3127 8316 3313 8324
rect 3587 8316 3833 8324
rect 3887 8316 3913 8324
rect 3927 8316 4013 8324
rect 4087 8316 4233 8324
rect 4267 8316 4373 8324
rect 4507 8316 5033 8324
rect 5087 8316 5513 8324
rect 5547 8316 6033 8324
rect 6056 8316 6313 8324
rect 647 8296 753 8304
rect 1067 8296 1193 8304
rect 1787 8296 2093 8304
rect 2147 8296 2253 8304
rect 2347 8296 2513 8304
rect 2627 8296 2853 8304
rect 3267 8296 3293 8304
rect 3347 8296 3413 8304
rect 3827 8296 3953 8304
rect 3987 8296 4353 8304
rect 4367 8296 4533 8304
rect 4647 8296 4813 8304
rect 4947 8296 5313 8304
rect 6056 8304 6064 8316
rect 6407 8316 6513 8324
rect 6547 8316 6713 8324
rect 6856 8324 6864 8333
rect 6816 8316 7313 8324
rect 6816 8307 6824 8316
rect 7567 8316 7893 8324
rect 7907 8316 7953 8324
rect 8167 8316 8424 8324
rect 8416 8307 8424 8316
rect 8696 8316 8913 8324
rect 8696 8307 8704 8316
rect 8927 8316 9133 8324
rect 9167 8316 9393 8324
rect 9427 8316 9833 8324
rect 9927 8316 10073 8324
rect 10127 8316 10293 8324
rect 10307 8316 10553 8324
rect 10607 8316 10693 8324
rect 11227 8316 11404 8324
rect 5527 8296 6064 8304
rect 6087 8296 6193 8304
rect 6207 8296 6333 8304
rect 6667 8296 6813 8304
rect 7027 8296 7093 8304
rect 7907 8296 8073 8304
rect 8107 8296 8133 8304
rect 8187 8296 8213 8304
rect 8467 8296 8553 8304
rect 8567 8296 8573 8304
rect 9447 8296 9493 8304
rect 9887 8296 10044 8304
rect 1107 8276 1813 8284
rect 1867 8276 2133 8284
rect 2667 8276 2893 8284
rect 3067 8276 3553 8284
rect 3607 8276 3653 8284
rect 3847 8276 4473 8284
rect 4627 8276 4653 8284
rect 4747 8276 5133 8284
rect 5387 8276 5453 8284
rect 5627 8276 5673 8284
rect 5847 8276 6093 8284
rect 6127 8276 6173 8284
rect 6187 8276 6373 8284
rect 6747 8276 6853 8284
rect 8367 8276 8433 8284
rect 9647 8276 9693 8284
rect 10036 8284 10044 8296
rect 10067 8296 10093 8304
rect 10347 8296 10453 8304
rect 10587 8296 10653 8304
rect 10136 8284 10144 8293
rect 10036 8276 10344 8284
rect 3527 8256 3553 8264
rect 3747 8256 4633 8264
rect 4687 8256 4713 8264
rect 4867 8256 5353 8264
rect 5807 8256 6613 8264
rect 6727 8256 7973 8264
rect 7987 8256 7993 8264
rect 8947 8256 10253 8264
rect 10336 8264 10344 8276
rect 10367 8276 10573 8284
rect 11107 8276 11404 8284
rect 10336 8256 10593 8264
rect 10607 8256 10633 8264
rect 2247 8236 3153 8244
rect 5047 8236 5673 8244
rect 6567 8236 7013 8244
rect 7927 8236 8573 8244
rect 8587 8236 8753 8244
rect 9467 8236 9513 8244
rect 4107 8216 4193 8224
rect 4207 8216 4953 8224
rect 4967 8216 5093 8224
rect 5107 8216 6573 8224
rect 6687 8216 7753 8224
rect 7947 8216 9673 8224
rect 9687 8216 9693 8224
rect 1247 8196 2813 8204
rect 5007 8196 6533 8204
rect 6556 8196 7133 8204
rect 3147 8176 4553 8184
rect 5267 8176 5553 8184
rect 6556 8184 6564 8196
rect 7147 8196 7333 8204
rect 7587 8196 11013 8204
rect 5587 8176 6564 8184
rect 6587 8176 7113 8184
rect 7887 8176 8313 8184
rect 8647 8176 11233 8184
rect 2487 8156 3053 8164
rect 3067 8156 4273 8164
rect 4867 8156 4893 8164
rect 5287 8156 7353 8164
rect 7407 8156 7453 8164
rect 4247 8136 5793 8144
rect 5827 8136 5873 8144
rect 6087 8136 6133 8144
rect 6187 8136 9173 8144
rect 9187 8136 9473 8144
rect 9487 8136 9513 8144
rect 9847 8136 9893 8144
rect 3047 8116 5273 8124
rect 5527 8116 5613 8124
rect 5647 8116 8133 8124
rect 687 8096 773 8104
rect 787 8096 833 8104
rect 2807 8096 3853 8104
rect 3967 8096 4373 8104
rect 4407 8096 5533 8104
rect 5787 8096 6153 8104
rect 6227 8096 6713 8104
rect 7087 8096 8273 8104
rect 47 8076 53 8084
rect 67 8076 713 8084
rect 727 8076 873 8084
rect 887 8076 1013 8084
rect 2867 8076 3013 8084
rect 3027 8076 3213 8084
rect 3227 8076 3513 8084
rect 3527 8076 3873 8084
rect 4307 8076 4573 8084
rect 4647 8076 7613 8084
rect 7627 8076 8093 8084
rect 8607 8076 8793 8084
rect 8807 8076 9153 8084
rect 9227 8076 9413 8084
rect 9707 8076 9913 8084
rect 10687 8076 10713 8084
rect 10847 8076 10913 8084
rect 10967 8076 11113 8084
rect 407 8056 813 8064
rect 1827 8056 2313 8064
rect 4367 8056 4433 8064
rect 4456 8056 5833 8064
rect 647 8036 913 8044
rect 1307 8036 1473 8044
rect 1547 8036 1573 8044
rect 1867 8036 2013 8044
rect 2727 8036 2753 8044
rect 2787 8036 3253 8044
rect 3587 8036 3713 8044
rect 3887 8036 3953 8044
rect 4007 8036 4033 8044
rect 4456 8044 4464 8056
rect 5927 8056 6593 8064
rect 6807 8056 7084 8064
rect 7076 8047 7084 8056
rect 7187 8056 7493 8064
rect 9207 8056 9253 8064
rect 9767 8056 9993 8064
rect 10167 8056 10253 8064
rect 10507 8056 10573 8064
rect 10747 8056 10773 8064
rect 10787 8056 10953 8064
rect 4287 8036 4464 8044
rect 4847 8036 5053 8044
rect 5107 8036 5193 8044
rect 5287 8036 5313 8044
rect 5367 8036 5533 8044
rect 5567 8036 5793 8044
rect 5847 8036 6053 8044
rect 6067 8036 6313 8044
rect 6747 8036 6853 8044
rect 7127 8036 7253 8044
rect 7327 8036 7393 8044
rect 7847 8036 8053 8044
rect 8227 8036 8333 8044
rect 8747 8036 8993 8044
rect 9007 8036 9053 8044
rect 9247 8036 9273 8044
rect 9967 8036 10033 8044
rect 10227 8036 10373 8044
rect 367 8016 493 8024
rect 507 8016 633 8024
rect 1267 8016 1553 8024
rect 1667 8016 1733 8024
rect 1747 8016 2213 8024
rect 2267 8016 2293 8024
rect 2327 8016 2733 8024
rect 2827 8016 2973 8024
rect 3007 8016 3913 8024
rect 4007 8016 4153 8024
rect 5127 8016 5424 8024
rect 1587 7996 1773 8004
rect 2807 7996 2893 8004
rect 2907 7996 3033 8004
rect 3047 7996 3193 8004
rect 4207 7996 4313 8004
rect 4447 7996 4513 8004
rect 4647 7996 4693 8004
rect 5367 7996 5393 8004
rect 5416 8004 5424 8016
rect 5447 8016 5493 8024
rect 5667 8016 5793 8024
rect 5827 8016 5913 8024
rect 5947 8016 6033 8024
rect 6316 8024 6324 8033
rect 6316 8016 6353 8024
rect 6627 8016 6813 8024
rect 7147 8016 7213 8024
rect 7387 8016 7573 8024
rect 7607 8016 7933 8024
rect 8127 8016 8193 8024
rect 8296 8016 9004 8024
rect 5416 7996 5933 8004
rect 5967 7996 6073 8004
rect 6227 7996 6593 8004
rect 6847 7996 7704 8004
rect 687 7976 713 7984
rect 1227 7976 1773 7984
rect 2187 7976 2773 7984
rect 2787 7976 3193 7984
rect 4247 7976 4413 7984
rect 4427 7976 5013 7984
rect 5107 7976 5713 7984
rect 5747 7976 5813 7984
rect 6007 7976 7613 7984
rect 7696 7984 7704 7996
rect 7727 7996 7833 8004
rect 8296 8004 8304 8016
rect 8087 7996 8304 8004
rect 8327 7996 8533 8004
rect 8996 8004 9004 8016
rect 9027 8016 9433 8024
rect 9447 8016 9453 8024
rect 9507 8016 9753 8024
rect 9927 8016 10013 8024
rect 8996 7996 11153 8004
rect 7696 7976 7813 7984
rect 8247 7976 8753 7984
rect 3507 7956 5673 7964
rect 5707 7956 7753 7964
rect 1047 7936 1133 7944
rect 3247 7936 5253 7944
rect 5327 7936 5453 7944
rect 6047 7936 6413 7944
rect 7267 7936 7373 7944
rect 10707 7936 11273 7944
rect 3727 7916 5573 7924
rect 5727 7916 6613 7924
rect 6767 7916 6973 7924
rect 7447 7916 7633 7924
rect 7647 7916 7933 7924
rect 7947 7916 8353 7924
rect 10747 7916 10773 7924
rect 3607 7896 3693 7904
rect 3927 7896 5384 7904
rect 2087 7876 2273 7884
rect 2287 7876 2773 7884
rect 3487 7876 3533 7884
rect 3547 7876 3753 7884
rect 3767 7876 3933 7884
rect 4167 7876 4253 7884
rect 5376 7884 5384 7896
rect 5407 7896 5633 7904
rect 5687 7896 6373 7904
rect 6667 7896 8833 7904
rect 8847 7896 9133 7904
rect 9147 7896 10133 7904
rect 10147 7896 10273 7904
rect 10387 7896 10713 7904
rect 5376 7876 5633 7884
rect 5867 7876 6253 7884
rect 6447 7876 6573 7884
rect 6587 7876 6813 7884
rect 8167 7876 11233 7884
rect 1327 7856 1353 7864
rect 1447 7856 1653 7864
rect 1847 7856 1873 7864
rect 2247 7856 2573 7864
rect 2587 7856 2713 7864
rect 2727 7856 2993 7864
rect 3247 7856 3293 7864
rect 3707 7856 3893 7864
rect 3987 7856 4033 7864
rect 4067 7856 4973 7864
rect 5207 7856 5733 7864
rect 5847 7856 5873 7864
rect 5887 7856 6113 7864
rect 6267 7856 6493 7864
rect 6507 7856 6673 7864
rect 6687 7856 6833 7864
rect 7227 7856 7433 7864
rect 7627 7856 7853 7864
rect 7867 7856 7873 7864
rect 7907 7856 8413 7864
rect 8867 7856 9013 7864
rect 9076 7856 9604 7864
rect 247 7836 413 7844
rect 1347 7836 1393 7844
rect 1467 7836 1673 7844
rect 1687 7836 1893 7844
rect 1907 7836 2144 7844
rect 187 7816 453 7824
rect 927 7816 1153 7824
rect 1427 7816 2113 7824
rect 2136 7824 2144 7836
rect 2327 7836 2833 7844
rect 2847 7836 2933 7844
rect 2947 7836 3433 7844
rect 3987 7836 4113 7844
rect 4247 7836 5053 7844
rect 5347 7836 5373 7844
rect 5427 7836 5453 7844
rect 5667 7836 5724 7844
rect 2136 7816 2213 7824
rect 2227 7816 2333 7824
rect 3007 7816 3053 7824
rect 3747 7816 3873 7824
rect 3887 7816 3953 7824
rect 4107 7816 4253 7824
rect 4467 7816 4704 7824
rect 4696 7807 4704 7816
rect 5136 7824 5144 7833
rect 5716 7827 5724 7836
rect 5907 7836 5973 7844
rect 6136 7844 6144 7853
rect 6136 7836 6524 7844
rect 6176 7827 6184 7836
rect 4947 7816 5144 7824
rect 5747 7816 5913 7824
rect 6347 7816 6413 7824
rect 6467 7816 6493 7824
rect 6516 7824 6524 7836
rect 6867 7836 6913 7844
rect 7107 7836 7644 7844
rect 7636 7827 7644 7836
rect 7667 7836 7873 7844
rect 8207 7836 8273 7844
rect 8807 7836 8933 7844
rect 9027 7836 9053 7844
rect 9076 7827 9084 7856
rect 9167 7836 9533 7844
rect 6516 7816 6673 7824
rect 6947 7816 7133 7824
rect 7187 7816 7253 7824
rect 7407 7816 7593 7824
rect 8107 7816 8173 7824
rect 8187 7816 8253 7824
rect 8407 7816 8433 7824
rect 8587 7816 8613 7824
rect 8787 7816 8893 7824
rect 8907 7816 9073 7824
rect 447 7796 893 7804
rect 907 7796 1073 7804
rect 1387 7796 1453 7804
rect 1627 7796 1753 7804
rect 2047 7796 2473 7804
rect 3027 7796 4193 7804
rect 4367 7796 4433 7804
rect 4987 7796 5513 7804
rect 5547 7796 5853 7804
rect 5887 7796 6113 7804
rect 6147 7796 6293 7804
rect 6307 7796 6613 7804
rect 6827 7796 6913 7804
rect 7027 7796 7153 7804
rect 7407 7796 7513 7804
rect 7927 7796 8113 7804
rect 8587 7796 8653 7804
rect 8747 7796 8793 7804
rect 9096 7804 9104 7833
rect 9127 7816 9153 7824
rect 9527 7816 9553 7824
rect 9096 7796 9193 7804
rect 9576 7804 9584 7833
rect 9596 7827 9604 7856
rect 10107 7856 10153 7864
rect 10607 7856 11033 7864
rect 9627 7836 9713 7844
rect 9887 7836 9973 7844
rect 10067 7836 10173 7844
rect 10647 7836 10813 7844
rect 10867 7836 10933 7844
rect 10087 7816 10233 7824
rect 10547 7816 10613 7824
rect 10667 7816 10833 7824
rect 9576 7796 9853 7804
rect 10347 7796 10553 7804
rect 11307 7796 11404 7804
rect 1087 7776 1113 7784
rect 1947 7776 2453 7784
rect 2467 7776 3273 7784
rect 3287 7776 4253 7784
rect 4267 7776 5293 7784
rect 5307 7776 6073 7784
rect 6087 7776 6533 7784
rect 6547 7776 7333 7784
rect 7347 7776 9233 7784
rect 227 7756 1333 7764
rect 2927 7756 3953 7764
rect 3967 7756 4313 7764
rect 4327 7756 5804 7764
rect 947 7736 1473 7744
rect 4147 7736 5133 7744
rect 5147 7736 5773 7744
rect 5796 7744 5804 7756
rect 6107 7756 6293 7764
rect 6887 7756 7513 7764
rect 5796 7736 5893 7744
rect 6447 7736 6513 7744
rect 7047 7736 7153 7744
rect 7247 7736 7573 7744
rect 7747 7736 9293 7744
rect 9307 7736 9373 7744
rect 4047 7716 6573 7724
rect 4747 7696 4993 7704
rect 5067 7696 6284 7704
rect 2307 7676 4613 7684
rect 4627 7676 4733 7684
rect 5187 7676 5613 7684
rect 5907 7676 6253 7684
rect 6276 7684 6284 7696
rect 6307 7696 6733 7704
rect 6976 7696 7673 7704
rect 6976 7684 6984 7696
rect 7707 7696 8813 7704
rect 6276 7676 6984 7684
rect 7007 7676 7193 7684
rect 8987 7676 9473 7684
rect 967 7656 5253 7664
rect 5267 7656 5553 7664
rect 5587 7656 7013 7664
rect 8047 7656 8133 7664
rect 8687 7656 10693 7664
rect 3647 7636 4353 7644
rect 4447 7636 4933 7644
rect 5207 7636 5273 7644
rect 5287 7636 6113 7644
rect 6167 7636 6773 7644
rect 6787 7636 6793 7644
rect 3167 7616 4053 7624
rect 4147 7616 4293 7624
rect 4707 7616 5833 7624
rect 6087 7616 6753 7624
rect 6847 7616 6933 7624
rect 7056 7624 7064 7653
rect 8447 7636 9773 7644
rect 10187 7636 10353 7644
rect 7056 7616 7093 7624
rect 7307 7616 8253 7624
rect 8267 7616 8413 7624
rect 8927 7616 8953 7624
rect 10107 7616 10973 7624
rect 4627 7596 4753 7604
rect 4807 7596 4873 7604
rect 5427 7596 5493 7604
rect 5527 7596 5653 7604
rect 5727 7596 6713 7604
rect 6767 7596 6773 7604
rect 6787 7596 7253 7604
rect 7347 7596 7453 7604
rect 7647 7596 11233 7604
rect 647 7576 673 7584
rect 687 7576 1633 7584
rect 1647 7576 1793 7584
rect 3307 7576 3353 7584
rect 3407 7576 3693 7584
rect 4047 7576 4153 7584
rect 4567 7576 4573 7584
rect 4587 7576 4973 7584
rect 5087 7576 5293 7584
rect 5407 7576 5553 7584
rect 5807 7576 5993 7584
rect 6256 7576 6373 7584
rect 6256 7567 6264 7576
rect 6487 7576 6633 7584
rect 7167 7576 8313 7584
rect 8467 7576 8513 7584
rect 8947 7576 9133 7584
rect 9307 7576 9533 7584
rect 9547 7576 9613 7584
rect 9687 7576 9833 7584
rect 10547 7576 10773 7584
rect 11107 7576 11404 7584
rect 507 7556 653 7564
rect 887 7556 933 7564
rect 1487 7556 1613 7564
rect 1667 7556 1733 7564
rect 1847 7556 1893 7564
rect 1947 7556 1973 7564
rect 2396 7556 2633 7564
rect 2396 7547 2404 7556
rect 2647 7556 2753 7564
rect 2907 7556 3233 7564
rect 3607 7556 3793 7564
rect 3847 7556 3993 7564
rect 4327 7556 4473 7564
rect 4487 7556 4773 7564
rect 5047 7556 5064 7564
rect 567 7536 693 7544
rect 707 7536 1653 7544
rect 2107 7536 2133 7544
rect 2487 7536 2873 7544
rect 3387 7536 3473 7544
rect 3627 7536 4393 7544
rect 4467 7536 4533 7544
rect 4796 7544 4804 7553
rect 4567 7536 4804 7544
rect 5056 7544 5064 7556
rect 5087 7556 5673 7564
rect 5687 7556 5733 7564
rect 5767 7556 5933 7564
rect 6507 7556 6553 7564
rect 6747 7556 6824 7564
rect 5056 7536 5173 7544
rect 5467 7536 5533 7544
rect 5627 7536 5793 7544
rect 6027 7536 6153 7544
rect 6687 7536 6793 7544
rect 6816 7544 6824 7556
rect 7367 7556 7593 7564
rect 7607 7556 7653 7564
rect 7747 7556 7953 7564
rect 8227 7556 8293 7564
rect 8447 7556 8713 7564
rect 8967 7556 9013 7564
rect 9647 7556 9793 7564
rect 10487 7556 10553 7564
rect 10607 7556 10673 7564
rect 10747 7556 10833 7564
rect 6816 7536 7133 7544
rect 7216 7544 7224 7553
rect 7167 7536 7224 7544
rect 7447 7536 7633 7544
rect 7727 7536 7913 7544
rect 7947 7536 8153 7544
rect 8247 7536 8273 7544
rect 9287 7536 9393 7544
rect 9867 7536 9953 7544
rect 10087 7536 10313 7544
rect 11307 7536 11404 7544
rect 207 7516 673 7524
rect 1987 7516 2153 7524
rect 2187 7516 2413 7524
rect 3127 7516 3333 7524
rect 4607 7516 4693 7524
rect 4947 7516 5053 7524
rect 5347 7516 5453 7524
rect 5667 7516 5753 7524
rect 5867 7516 6213 7524
rect 6287 7516 6513 7524
rect 6747 7516 6813 7524
rect 6967 7516 7173 7524
rect 7267 7516 7673 7524
rect 7687 7516 7813 7524
rect 7987 7516 8353 7524
rect 8527 7516 8653 7524
rect 8667 7516 9333 7524
rect 9347 7516 9433 7524
rect 10127 7516 10173 7524
rect 10347 7516 10533 7524
rect 10587 7516 10693 7524
rect 10787 7516 10813 7524
rect 11007 7516 11193 7524
rect 1767 7496 1953 7504
rect 1967 7496 2373 7504
rect 2787 7496 3093 7504
rect 3107 7496 4433 7504
rect 4787 7496 4793 7504
rect 4807 7496 5273 7504
rect 5987 7496 6293 7504
rect 6667 7496 6833 7504
rect 7287 7496 7413 7504
rect 7487 7496 7493 7504
rect 7507 7496 7953 7504
rect 8167 7496 8993 7504
rect 9007 7496 9293 7504
rect 10187 7496 10993 7504
rect 4207 7476 4673 7484
rect 5327 7476 5553 7484
rect 5707 7476 6353 7484
rect 6707 7476 6733 7484
rect 6927 7476 7133 7484
rect 7887 7476 8173 7484
rect 8487 7476 8693 7484
rect 8887 7476 8993 7484
rect 9227 7476 9333 7484
rect 2127 7456 2393 7464
rect 2407 7456 2613 7464
rect 2627 7456 2853 7464
rect 2867 7456 3093 7464
rect 3867 7456 4673 7464
rect 4687 7456 5373 7464
rect 5447 7456 6413 7464
rect 6567 7456 7053 7464
rect 7087 7456 7373 7464
rect 8207 7456 11033 7464
rect 3787 7436 4593 7444
rect 4987 7436 5193 7444
rect 5527 7436 6193 7444
rect 6367 7436 8933 7444
rect 9407 7436 10273 7444
rect 10987 7436 11013 7444
rect 3467 7416 3553 7424
rect 3567 7416 3813 7424
rect 3827 7416 5533 7424
rect 5556 7416 5853 7424
rect 3507 7396 3773 7404
rect 5556 7404 5564 7416
rect 5907 7416 6953 7424
rect 7067 7416 7873 7424
rect 7896 7416 8873 7424
rect 4867 7396 5564 7404
rect 5587 7396 5773 7404
rect 5787 7396 6033 7404
rect 6247 7396 6273 7404
rect 6507 7396 6553 7404
rect 6587 7396 6773 7404
rect 7896 7404 7904 7416
rect 9187 7416 10053 7424
rect 10067 7416 10373 7424
rect 10387 7416 10833 7424
rect 10847 7416 11033 7424
rect 6887 7396 7904 7404
rect 7927 7396 8633 7404
rect 9087 7396 11253 7404
rect 1327 7376 1433 7384
rect 1447 7376 1453 7384
rect 2587 7376 2793 7384
rect 2847 7376 2973 7384
rect 2987 7376 3233 7384
rect 3267 7376 3433 7384
rect 3727 7376 3753 7384
rect 3867 7376 3953 7384
rect 3987 7376 4013 7384
rect 4027 7376 4073 7384
rect 4707 7376 5073 7384
rect 5167 7376 5313 7384
rect 5707 7376 5953 7384
rect 6247 7376 6333 7384
rect 6447 7376 6833 7384
rect 7287 7376 7493 7384
rect 8147 7376 8173 7384
rect 8247 7376 9013 7384
rect 9027 7376 9113 7384
rect 9827 7376 10533 7384
rect 10547 7376 10553 7384
rect 10587 7376 10633 7384
rect 10727 7376 10753 7384
rect 10867 7376 11053 7384
rect 107 7356 213 7364
rect 307 7356 713 7364
rect 727 7356 973 7364
rect 1136 7364 1144 7373
rect 1136 7356 1393 7364
rect 1407 7356 1493 7364
rect 1827 7356 1873 7364
rect 2087 7356 2193 7364
rect 2927 7356 3213 7364
rect 3227 7356 3293 7364
rect 3527 7356 4193 7364
rect 4307 7356 4393 7364
rect 4847 7356 4913 7364
rect 4967 7356 5093 7364
rect 5227 7356 5253 7364
rect 5476 7347 5484 7373
rect 5507 7356 5793 7364
rect 6467 7356 6693 7364
rect 6747 7356 6893 7364
rect 7007 7356 7293 7364
rect 7327 7356 7453 7364
rect 7967 7356 8233 7364
rect 8707 7356 9153 7364
rect 9367 7356 9833 7364
rect 9927 7356 10053 7364
rect 10107 7356 10313 7364
rect 10327 7356 10744 7364
rect 10736 7347 10744 7356
rect 207 7336 453 7344
rect 587 7336 653 7344
rect 1087 7336 1113 7344
rect 1167 7336 1373 7344
rect 1647 7336 1853 7344
rect 2007 7336 2273 7344
rect 2287 7336 2333 7344
rect 2767 7336 2813 7344
rect 3047 7336 3113 7344
rect 4107 7336 4213 7344
rect 4947 7336 4973 7344
rect 5007 7336 5393 7344
rect 5627 7336 5753 7344
rect 6347 7336 6513 7344
rect 6736 7336 6873 7344
rect 247 7316 293 7324
rect 947 7316 1613 7324
rect 1907 7316 2293 7324
rect 2367 7316 2373 7324
rect 2387 7316 2553 7324
rect 2687 7316 2813 7324
rect 2987 7316 3013 7324
rect 4896 7324 4904 7333
rect 4896 7316 4933 7324
rect 5087 7316 5193 7324
rect 5207 7316 5333 7324
rect 5447 7316 5533 7324
rect 5547 7316 6073 7324
rect 6736 7324 6744 7336
rect 6927 7336 6973 7344
rect 7147 7336 7473 7344
rect 7747 7336 7933 7344
rect 8227 7336 8253 7344
rect 8867 7336 9053 7344
rect 9147 7336 9313 7344
rect 9587 7336 10033 7344
rect 10087 7336 10473 7344
rect 10827 7336 10953 7344
rect 10967 7336 11053 7344
rect 6727 7316 6744 7324
rect 7016 7324 7024 7333
rect 7007 7316 7024 7324
rect 7307 7316 7653 7324
rect 7947 7316 8093 7324
rect 9007 7316 9093 7324
rect 9327 7316 9413 7324
rect 9447 7316 9553 7324
rect 10787 7316 10853 7324
rect 11327 7316 11404 7324
rect 287 7296 413 7304
rect 427 7296 433 7304
rect 447 7296 533 7304
rect 707 7296 1193 7304
rect 1367 7296 1393 7304
rect 1527 7296 2113 7304
rect 2527 7296 4733 7304
rect 4747 7296 4913 7304
rect 5167 7296 5613 7304
rect 6756 7304 6764 7313
rect 6567 7296 6764 7304
rect 6787 7296 7024 7304
rect 4907 7276 4933 7284
rect 5167 7276 5233 7284
rect 5287 7276 5413 7284
rect 5527 7276 5833 7284
rect 6687 7276 6993 7284
rect 7016 7284 7024 7296
rect 7016 7276 8073 7284
rect 9247 7276 9593 7284
rect 9607 7276 9633 7284
rect 9967 7276 10033 7284
rect 3267 7256 3793 7264
rect 3807 7256 5393 7264
rect 6227 7256 7313 7264
rect 5487 7236 6053 7244
rect 6487 7236 6773 7244
rect 6987 7236 7253 7244
rect 7527 7236 8253 7244
rect 8547 7236 8633 7244
rect 3767 7216 4193 7224
rect 5267 7216 5513 7224
rect 5967 7216 6273 7224
rect 6307 7216 6533 7224
rect 7127 7216 8293 7224
rect 8567 7216 8613 7224
rect 5027 7196 5073 7204
rect 5607 7196 5933 7204
rect 6027 7196 7153 7204
rect 7167 7196 7253 7204
rect 7867 7196 8333 7204
rect 8347 7196 8413 7204
rect 1067 7182 1133 7190
rect 1287 7176 1333 7184
rect 1507 7176 1633 7184
rect 2127 7176 5193 7184
rect 5347 7176 5693 7184
rect 5707 7176 5713 7184
rect 5947 7176 6313 7184
rect 6527 7176 7213 7184
rect 8327 7176 9693 7184
rect 4127 7156 8513 7164
rect 1927 7136 3033 7144
rect 3067 7136 3193 7144
rect 3207 7136 5053 7144
rect 5067 7136 5353 7144
rect 5367 7136 6793 7144
rect 6827 7136 7633 7144
rect 8147 7136 8173 7144
rect 10547 7136 10753 7144
rect 507 7116 553 7124
rect 1847 7116 1913 7124
rect 4067 7116 4813 7124
rect 4947 7116 5984 7124
rect 67 7096 513 7104
rect 527 7096 813 7104
rect 827 7096 1253 7104
rect 1807 7096 1873 7104
rect 3167 7096 3193 7104
rect 3527 7096 3573 7104
rect 3627 7096 3733 7104
rect 4527 7096 5133 7104
rect 5147 7096 5273 7104
rect 5667 7096 5773 7104
rect 5976 7104 5984 7116
rect 6007 7116 6213 7124
rect 6507 7116 6573 7124
rect 6967 7116 7293 7124
rect 7427 7116 7893 7124
rect 7907 7116 8153 7124
rect 9267 7116 9413 7124
rect 9427 7116 9573 7124
rect 9587 7116 10233 7124
rect 10247 7116 10253 7124
rect 10487 7116 10613 7124
rect 5976 7096 6104 7104
rect 87 7076 173 7084
rect 407 7076 853 7084
rect 907 7076 933 7084
rect 947 7076 953 7084
rect 1207 7076 1233 7084
rect 1747 7076 1893 7084
rect 2287 7076 2413 7084
rect 2627 7076 2653 7084
rect 2747 7076 2893 7084
rect 3407 7076 3473 7084
rect 3647 7076 3813 7084
rect 4527 7076 4684 7084
rect 1227 7056 1273 7064
rect 2156 7064 2164 7073
rect 2156 7056 2633 7064
rect 4327 7056 4393 7064
rect 4407 7056 4633 7064
rect 4676 7064 4684 7076
rect 4707 7076 4733 7084
rect 4787 7076 4813 7084
rect 4827 7076 4993 7084
rect 5247 7076 5733 7084
rect 5747 7076 5853 7084
rect 6047 7076 6073 7084
rect 6096 7084 6104 7096
rect 6127 7096 6713 7104
rect 6727 7096 6793 7104
rect 6927 7096 7013 7104
rect 7476 7096 8373 7104
rect 6096 7076 6453 7084
rect 6676 7076 6753 7084
rect 4676 7056 4713 7064
rect 4907 7056 5033 7064
rect 5087 7056 5253 7064
rect 5307 7056 5353 7064
rect 5656 7056 5713 7064
rect 107 7036 193 7044
rect 1147 7036 1293 7044
rect 2147 7036 2213 7044
rect 2407 7036 2713 7044
rect 2887 7036 3133 7044
rect 3347 7036 3593 7044
rect 4147 7036 4293 7044
rect 4747 7036 4853 7044
rect 5656 7044 5664 7056
rect 5767 7056 5953 7064
rect 6027 7056 6233 7064
rect 6676 7064 6684 7076
rect 7476 7084 7484 7096
rect 8527 7096 8613 7104
rect 9067 7096 9113 7104
rect 10527 7096 10544 7104
rect 6936 7076 7484 7084
rect 6307 7056 6684 7064
rect 6936 7064 6944 7076
rect 8167 7076 8273 7084
rect 8407 7076 8593 7084
rect 8867 7076 9073 7084
rect 10487 7076 10513 7084
rect 6707 7056 6944 7064
rect 6967 7056 6993 7064
rect 7047 7056 7173 7064
rect 7496 7047 7504 7073
rect 8227 7056 8633 7064
rect 8787 7056 8913 7064
rect 8927 7056 9293 7064
rect 10327 7056 10493 7064
rect 10536 7064 10544 7096
rect 10647 7096 10793 7104
rect 10567 7076 10773 7084
rect 10967 7076 11053 7084
rect 10536 7056 10573 7064
rect 11396 7064 11404 7084
rect 11307 7056 11404 7064
rect 4887 7036 5664 7044
rect 5687 7036 5973 7044
rect 5987 7036 6153 7044
rect 6467 7036 6973 7044
rect 7067 7036 7273 7044
rect 7687 7036 7713 7044
rect 7867 7036 8133 7044
rect 8687 7036 8873 7044
rect 9027 7036 9133 7044
rect 687 7016 1173 7024
rect 2687 7016 2733 7024
rect 3367 7016 3873 7024
rect 3887 7016 4033 7024
rect 4287 7016 4753 7024
rect 4987 7016 5073 7024
rect 5127 7016 5713 7024
rect 7547 7016 7693 7024
rect 7787 7016 8413 7024
rect 9107 7016 11253 7024
rect 987 6996 1093 7004
rect 1107 6996 2173 7004
rect 4267 6996 4453 7004
rect 4467 6996 4493 7004
rect 4507 6996 4933 7004
rect 5716 6996 6493 7004
rect 587 6976 693 6984
rect 947 6976 1153 6984
rect 5716 6984 5724 6996
rect 6527 6996 6913 7004
rect 7227 6996 8133 7004
rect 1747 6976 5724 6984
rect 5747 6976 6473 6984
rect 6507 6976 7764 6984
rect 867 6956 1393 6964
rect 1407 6956 1593 6964
rect 1727 6956 3213 6964
rect 4447 6956 5333 6964
rect 5407 6956 6073 6964
rect 6387 6956 6993 6964
rect 7756 6964 7764 6976
rect 9107 6976 9673 6984
rect 7756 6956 7913 6964
rect 8767 6956 9233 6964
rect 9367 6956 9553 6964
rect 9727 6956 9793 6964
rect 1207 6936 1653 6944
rect 3847 6936 4053 6944
rect 4067 6936 4493 6944
rect 5307 6936 5593 6944
rect 5627 6936 6133 6944
rect 6427 6936 7613 6944
rect 7827 6936 10393 6944
rect 10407 6936 10513 6944
rect 1127 6916 1513 6924
rect 3627 6916 3853 6924
rect 4087 6916 4253 6924
rect 4347 6916 5113 6924
rect 5127 6916 5673 6924
rect 5727 6916 8753 6924
rect 10747 6916 11053 6924
rect 11067 6916 11213 6924
rect 11227 6916 11313 6924
rect 267 6896 473 6904
rect 487 6896 673 6904
rect 1667 6896 1693 6904
rect 2167 6896 2433 6904
rect 3547 6896 3853 6904
rect 3867 6896 4073 6904
rect 4367 6896 4433 6904
rect 5427 6896 6553 6904
rect 6567 6896 6813 6904
rect 6827 6896 7433 6904
rect 7447 6896 7553 6904
rect 7947 6896 8093 6904
rect 9387 6896 9613 6904
rect 9907 6896 10053 6904
rect 11107 6896 11253 6904
rect 447 6876 493 6884
rect 747 6876 893 6884
rect 907 6876 1113 6884
rect 1187 6876 1413 6884
rect 1487 6876 1533 6884
rect 1587 6876 1693 6884
rect 1867 6876 2293 6884
rect 3767 6876 3813 6884
rect 4107 6876 4353 6884
rect 4367 6876 4513 6884
rect 4527 6876 4613 6884
rect 4847 6876 5193 6884
rect 5267 6876 5293 6884
rect 5387 6876 5753 6884
rect 5767 6876 5793 6884
rect 5807 6876 5993 6884
rect 6047 6876 7024 6884
rect 227 6856 613 6864
rect 727 6856 913 6864
rect 927 6856 1153 6864
rect 1247 6856 1453 6864
rect 1687 6856 1933 6864
rect 2187 6856 2193 6864
rect 2207 6856 2353 6864
rect 2407 6856 2573 6864
rect 2667 6856 2713 6864
rect 2887 6856 2933 6864
rect 2947 6856 3053 6864
rect 3347 6856 3393 6864
rect 3416 6856 3573 6864
rect 467 6836 653 6844
rect 887 6836 913 6844
rect 2307 6836 2373 6844
rect 2616 6844 2624 6853
rect 2616 6836 2833 6844
rect 3087 6836 3293 6844
rect 3416 6844 3424 6856
rect 3647 6856 3833 6864
rect 4307 6856 4413 6864
rect 4507 6856 4553 6864
rect 4727 6856 4773 6864
rect 4827 6856 4853 6864
rect 5007 6856 5053 6864
rect 5327 6856 5593 6864
rect 5707 6856 5813 6864
rect 6027 6856 6113 6864
rect 6407 6856 6493 6864
rect 6767 6856 6973 6864
rect 7016 6864 7024 6876
rect 7047 6876 7473 6884
rect 7487 6876 7513 6884
rect 7767 6876 7973 6884
rect 8947 6876 9253 6884
rect 9347 6876 9413 6884
rect 10267 6876 10293 6884
rect 10347 6876 10573 6884
rect 10787 6876 10813 6884
rect 11047 6876 11164 6884
rect 7016 6856 7204 6864
rect 3367 6836 3424 6844
rect 4667 6836 5273 6844
rect 5607 6836 5853 6844
rect 5867 6836 6053 6844
rect 6747 6836 6953 6844
rect 6967 6836 7013 6844
rect 7196 6844 7204 6856
rect 7227 6856 7333 6864
rect 7467 6856 7533 6864
rect 8007 6856 8073 6864
rect 8147 6856 8193 6864
rect 8487 6856 8993 6864
rect 9127 6856 9153 6864
rect 10247 6856 10313 6864
rect 10567 6856 10753 6864
rect 10807 6856 11013 6864
rect 11156 6864 11164 6876
rect 11156 6856 11233 6864
rect 7196 6836 7713 6844
rect 8147 6836 8233 6844
rect 8567 6836 8573 6844
rect 8587 6836 8673 6844
rect 9047 6836 9133 6844
rect 2847 6816 3173 6824
rect 3207 6816 3353 6824
rect 3447 6816 4033 6824
rect 4047 6816 4333 6824
rect 4347 6816 4613 6824
rect 4667 6816 5573 6824
rect 5827 6816 6493 6824
rect 6967 6816 7953 6824
rect 7967 6816 8373 6824
rect 8547 6816 9453 6824
rect 9467 6816 10033 6824
rect 10047 6816 10653 6824
rect 10907 6816 11013 6824
rect 3327 6796 4113 6804
rect 4547 6796 4573 6804
rect 4607 6796 6033 6804
rect 6127 6796 6773 6804
rect 6987 6796 7253 6804
rect 8127 6796 8233 6804
rect 8247 6796 9053 6804
rect 4187 6776 4873 6784
rect 4967 6776 5233 6784
rect 5287 6776 6013 6784
rect 6087 6776 7413 6784
rect 7427 6776 8433 6784
rect 9407 6776 9493 6784
rect 2427 6756 2653 6764
rect 3667 6756 5973 6764
rect 6187 6756 6313 6764
rect 6907 6756 7053 6764
rect 8027 6756 9433 6764
rect 207 6736 1613 6744
rect 1627 6736 1953 6744
rect 1967 6736 2093 6744
rect 4347 6736 5473 6744
rect 7847 6736 8673 6744
rect 8727 6736 9093 6744
rect 9187 6736 9653 6744
rect 10547 6736 10573 6744
rect 4487 6716 5093 6724
rect 5107 6716 5413 6724
rect 5847 6716 6113 6724
rect 6347 6716 6513 6724
rect 6947 6716 7193 6724
rect 8207 6716 8253 6724
rect 8267 6716 8913 6724
rect 3127 6696 4533 6704
rect 4627 6696 4693 6704
rect 4927 6696 5373 6704
rect 5547 6696 6173 6704
rect 1467 6676 2313 6684
rect 4727 6676 7673 6684
rect 727 6656 4713 6664
rect 5427 6656 6213 6664
rect 6867 6656 7453 6664
rect 1827 6636 1913 6644
rect 1927 6636 2213 6644
rect 4616 6636 4673 6644
rect 627 6616 673 6624
rect 1387 6616 1453 6624
rect 1467 6616 1713 6624
rect 1787 6616 1824 6624
rect 427 6596 653 6604
rect 1207 6596 1253 6604
rect 1267 6596 1413 6604
rect 1767 6596 1793 6604
rect 1816 6604 1824 6616
rect 2247 6616 2713 6624
rect 2727 6616 2873 6624
rect 3427 6616 3593 6624
rect 3827 6616 3873 6624
rect 4616 6624 4624 6636
rect 5107 6636 5153 6644
rect 5167 6636 5353 6644
rect 5367 6636 5533 6644
rect 5567 6636 5673 6644
rect 6047 6636 6353 6644
rect 7527 6636 7833 6644
rect 4487 6616 4624 6624
rect 5327 6616 5573 6624
rect 5847 6616 5993 6624
rect 6047 6616 6193 6624
rect 6396 6616 6713 6624
rect 1816 6596 1893 6604
rect 1907 6596 2373 6604
rect 2687 6596 2833 6604
rect 3047 6596 3133 6604
rect 3187 6596 3893 6604
rect 4527 6596 4644 6604
rect 4636 6587 4644 6596
rect 5367 6596 5553 6604
rect 6396 6604 6404 6616
rect 6727 6616 7493 6624
rect 7507 6616 7973 6624
rect 9127 6616 9153 6624
rect 10996 6624 11004 6633
rect 9967 6616 11073 6624
rect 11296 6607 11304 6633
rect 6027 6596 6404 6604
rect 6427 6596 6453 6604
rect 6687 6596 6793 6604
rect 6807 6596 6973 6604
rect 7047 6596 7233 6604
rect 7787 6596 7813 6604
rect 8307 6596 8453 6604
rect 8507 6596 8693 6604
rect 8747 6596 8753 6604
rect 8767 6596 8953 6604
rect 10127 6596 10344 6604
rect 647 6576 813 6584
rect 1327 6576 1473 6584
rect 1747 6576 1833 6584
rect 3767 6576 4033 6584
rect 4047 6576 4133 6584
rect 4367 6576 4473 6584
rect 4507 6576 4573 6584
rect 5027 6576 5213 6584
rect 5247 6576 5293 6584
rect 7276 6584 7284 6593
rect 10336 6587 10344 6596
rect 10547 6596 10693 6604
rect 6487 6576 7284 6584
rect 7307 6576 7533 6584
rect 7907 6576 7953 6584
rect 8987 6576 9173 6584
rect 9187 6576 9373 6584
rect 9507 6576 9633 6584
rect 9647 6576 9893 6584
rect 9907 6576 10073 6584
rect 10347 6576 10473 6584
rect 10507 6576 10993 6584
rect 11007 6576 11213 6584
rect 387 6556 1113 6564
rect 1407 6556 1773 6564
rect 1787 6556 1813 6564
rect 2947 6556 3153 6564
rect 3467 6556 3653 6564
rect 3667 6556 3853 6564
rect 3887 6556 4113 6564
rect 4567 6556 4713 6564
rect 4847 6556 5333 6564
rect 5447 6556 6433 6564
rect 6787 6556 6813 6564
rect 7567 6556 7693 6564
rect 7707 6556 7753 6564
rect 7767 6556 7953 6564
rect 8027 6556 8153 6564
rect 8487 6556 8713 6564
rect 10147 6556 10593 6564
rect 1447 6536 1573 6544
rect 4727 6536 5433 6544
rect 5807 6536 5833 6544
rect 5867 6536 6673 6544
rect 6707 6536 6793 6544
rect 6987 6536 7093 6544
rect 7207 6536 7253 6544
rect 8847 6536 8913 6544
rect 8927 6536 9333 6544
rect 947 6516 1473 6524
rect 3067 6516 4313 6524
rect 5927 6516 6233 6524
rect 6247 6516 6553 6524
rect 6747 6516 7013 6524
rect 7227 6516 7393 6524
rect 7827 6516 9173 6524
rect 11047 6516 11093 6524
rect 927 6496 973 6504
rect 1047 6496 1153 6504
rect 1167 6496 2053 6504
rect 2087 6496 2493 6504
rect 2567 6496 2753 6504
rect 3687 6496 4553 6504
rect 4607 6496 4673 6504
rect 5447 6496 5933 6504
rect 6287 6496 6513 6504
rect 6536 6496 7813 6504
rect 1527 6476 2533 6484
rect 2547 6476 4593 6484
rect 5147 6476 5273 6484
rect 5987 6476 6013 6484
rect 6536 6484 6544 6496
rect 10647 6496 10833 6504
rect 10847 6496 11253 6504
rect 6027 6476 6544 6484
rect 6676 6476 6913 6484
rect 1707 6456 1753 6464
rect 1767 6456 2013 6464
rect 3787 6456 4753 6464
rect 4787 6456 4993 6464
rect 5047 6456 5333 6464
rect 6676 6464 6684 6476
rect 10867 6476 11113 6484
rect 5407 6456 6684 6464
rect 6787 6456 7413 6464
rect 8527 6456 9953 6464
rect 10107 6456 10593 6464
rect 1727 6436 1953 6444
rect 4147 6436 4793 6444
rect 4907 6436 5193 6444
rect 5207 6436 5473 6444
rect 5967 6436 7373 6444
rect 9147 6436 9593 6444
rect 9607 6436 9673 6444
rect 9707 6436 10073 6444
rect 10087 6436 10273 6444
rect 10387 6436 10533 6444
rect 10547 6436 10813 6444
rect 247 6416 273 6424
rect 296 6416 453 6424
rect 296 6404 304 6416
rect 487 6416 673 6424
rect 767 6416 1013 6424
rect 1027 6416 1393 6424
rect 1747 6416 1913 6424
rect 3587 6416 3613 6424
rect 3927 6416 4073 6424
rect 4087 6416 4093 6424
rect 4307 6416 4353 6424
rect 4827 6416 5313 6424
rect 5347 6416 5513 6424
rect 5827 6416 5973 6424
rect 6067 6416 6133 6424
rect 6147 6416 6413 6424
rect 7007 6416 7093 6424
rect 7107 6416 8093 6424
rect 8587 6416 8633 6424
rect 8987 6416 9113 6424
rect 9127 6416 9333 6424
rect 9627 6416 9653 6424
rect 9667 6416 9933 6424
rect 10567 6416 10793 6424
rect 216 6396 304 6404
rect 216 6387 224 6396
rect 507 6396 933 6404
rect 1147 6396 1193 6404
rect 1247 6396 1453 6404
rect 1647 6396 1713 6404
rect 2007 6396 2073 6404
rect 2247 6396 2473 6404
rect 2647 6396 2653 6404
rect 2667 6396 2713 6404
rect 3407 6396 3593 6404
rect 3767 6396 3813 6404
rect 3867 6396 4104 6404
rect 4096 6387 4104 6396
rect 5227 6396 5333 6404
rect 5747 6396 5813 6404
rect 6167 6396 6193 6404
rect 6367 6396 6453 6404
rect 7507 6396 7653 6404
rect 7936 6396 7993 6404
rect 267 6376 1093 6384
rect 1927 6376 1973 6384
rect 2067 6376 2253 6384
rect 2327 6376 2513 6384
rect 2587 6376 2773 6384
rect 3347 6376 3433 6384
rect 3487 6376 3833 6384
rect 3847 6376 3913 6384
rect 4547 6376 5033 6384
rect 5547 6376 5753 6384
rect 6596 6384 6604 6393
rect 7936 6387 7944 6396
rect 8227 6396 8413 6404
rect 8467 6396 8873 6404
rect 9047 6396 9073 6404
rect 9427 6396 9653 6404
rect 9667 6396 9873 6404
rect 9927 6396 10113 6404
rect 10127 6396 10304 6404
rect 10296 6387 10304 6396
rect 10367 6396 10573 6404
rect 6527 6376 6993 6384
rect 7167 6376 7393 6384
rect 7527 6376 7673 6384
rect 7987 6376 8193 6384
rect 8667 6376 8693 6384
rect 8827 6376 8853 6384
rect 8907 6376 8933 6384
rect 9227 6376 9553 6384
rect 9807 6376 9833 6384
rect 10316 6367 10324 6393
rect 10487 6376 10553 6384
rect 11267 6376 11293 6384
rect 707 6356 953 6364
rect 967 6356 1013 6364
rect 1027 6356 1373 6364
rect 1867 6356 1973 6364
rect 2567 6356 2733 6364
rect 2747 6356 2893 6364
rect 3907 6356 3993 6364
rect 4007 6356 4573 6364
rect 5507 6356 5593 6364
rect 5607 6356 5773 6364
rect 5967 6356 6053 6364
rect 6267 6356 6444 6364
rect 1547 6336 1933 6344
rect 1947 6336 2553 6344
rect 5307 6336 5733 6344
rect 6436 6344 6444 6356
rect 6647 6356 6773 6364
rect 7007 6356 7133 6364
rect 7447 6356 7813 6364
rect 7827 6356 7893 6364
rect 8387 6356 8433 6364
rect 9487 6356 9813 6364
rect 9867 6356 10293 6364
rect 10687 6356 10813 6364
rect 10827 6356 10873 6364
rect 6436 6336 6953 6344
rect 7547 6336 7713 6344
rect 7727 6336 7853 6344
rect 8427 6336 8533 6344
rect 6456 6316 7093 6324
rect 3907 6296 4473 6304
rect 4487 6296 4873 6304
rect 5567 6296 5673 6304
rect 5687 6296 5953 6304
rect 6456 6304 6464 6316
rect 7327 6316 7713 6324
rect 11187 6316 11213 6324
rect 6167 6296 6464 6304
rect 6547 6296 6693 6304
rect 6927 6296 11313 6304
rect 807 6276 6673 6284
rect 6696 6276 8613 6284
rect 847 6256 3113 6264
rect 4387 6256 5093 6264
rect 6696 6264 6704 6276
rect 6487 6256 6704 6264
rect 6767 6256 7053 6264
rect 87 6236 393 6244
rect 1187 6236 1213 6244
rect 3407 6236 4373 6244
rect 4387 6236 6013 6244
rect 6327 6236 6373 6244
rect 6387 6236 6573 6244
rect 6687 6236 7973 6244
rect 8007 6236 8133 6244
rect 2267 6216 3373 6224
rect 4647 6216 5524 6224
rect 5247 6196 5493 6204
rect 5516 6204 5524 6216
rect 6567 6216 7113 6224
rect 7127 6216 7153 6224
rect 7647 6216 8193 6224
rect 10687 6216 10713 6224
rect 5516 6196 7053 6204
rect 8707 6196 10753 6204
rect 247 6176 1273 6184
rect 2107 6176 2473 6184
rect 2487 6176 3133 6184
rect 4027 6176 5533 6184
rect 6127 6176 8433 6184
rect 8627 6176 10513 6184
rect 1007 6156 1233 6164
rect 1247 6156 1533 6164
rect 2527 6156 2793 6164
rect 3767 6156 4173 6164
rect 4587 6156 5833 6164
rect 6187 6156 6273 6164
rect 6567 6156 7033 6164
rect 7047 6156 7173 6164
rect 7187 6156 7193 6164
rect 7207 6156 7473 6164
rect 7647 6156 8033 6164
rect 8047 6156 9393 6164
rect 547 6136 693 6144
rect 707 6136 1173 6144
rect 1187 6136 1273 6144
rect 1367 6136 1953 6144
rect 1967 6136 2433 6144
rect 2447 6136 2493 6144
rect 3187 6136 3473 6144
rect 4647 6136 5744 6144
rect 5736 6127 5744 6136
rect 6047 6136 6213 6144
rect 6227 6136 6553 6144
rect 6707 6136 6933 6144
rect 7627 6136 7684 6144
rect 7676 6127 7684 6136
rect 8187 6136 8213 6144
rect 9827 6136 10073 6144
rect 10087 6136 10413 6144
rect 207 6116 253 6124
rect 696 6116 913 6124
rect 696 6104 704 6116
rect 967 6116 1433 6124
rect 1447 6116 1493 6124
rect 1507 6116 1513 6124
rect 1807 6116 2053 6124
rect 2407 6116 2453 6124
rect 2467 6116 2533 6124
rect 2847 6116 2973 6124
rect 3427 6116 3473 6124
rect 3747 6116 3833 6124
rect 3867 6116 3973 6124
rect 4167 6116 4613 6124
rect 4627 6116 5473 6124
rect 5487 6116 5624 6124
rect 687 6096 704 6104
rect 727 6096 1153 6104
rect 1207 6096 1473 6104
rect 2007 6096 2093 6104
rect 2107 6096 2373 6104
rect 2387 6096 2833 6104
rect 2987 6096 3553 6104
rect 4827 6096 4873 6104
rect 5616 6104 5624 6116
rect 5647 6116 5693 6124
rect 6007 6116 6193 6124
rect 6667 6116 6733 6124
rect 6967 6116 6993 6124
rect 7187 6116 7393 6124
rect 7447 6116 7493 6124
rect 7867 6116 7913 6124
rect 8107 6116 8113 6124
rect 8347 6116 8373 6124
rect 8547 6116 8673 6124
rect 8907 6116 8973 6124
rect 9267 6116 9353 6124
rect 10107 6116 10153 6124
rect 10787 6116 10873 6124
rect 5616 6096 5673 6104
rect 5787 6096 5933 6104
rect 5947 6096 6033 6104
rect 6187 6096 6353 6104
rect 6367 6096 6373 6104
rect 6387 6096 6653 6104
rect 6867 6096 6893 6104
rect 7067 6096 7653 6104
rect 7907 6096 8073 6104
rect 8116 6104 8124 6113
rect 8116 6096 8653 6104
rect 8807 6096 8913 6104
rect 9167 6096 9593 6104
rect 9807 6096 9833 6104
rect 10067 6096 10133 6104
rect 10447 6096 11053 6104
rect 267 6076 453 6084
rect 587 6076 653 6084
rect 667 6076 733 6084
rect 1467 6076 1793 6084
rect 2087 6076 2273 6084
rect 2467 6076 2633 6084
rect 3347 6076 3733 6084
rect 4167 6076 4293 6084
rect 4367 6076 4633 6084
rect 4647 6076 4773 6084
rect 5327 6076 5453 6084
rect 5467 6076 6113 6084
rect 7587 6076 7653 6084
rect 7967 6076 8053 6084
rect 8187 6076 8213 6084
rect 8707 6076 9393 6084
rect 9407 6076 11253 6084
rect 227 6056 273 6064
rect 287 6056 433 6064
rect 4307 6056 4613 6064
rect 4627 6056 4833 6064
rect 6067 6056 7853 6064
rect 7947 6056 8293 6064
rect 8327 6056 8873 6064
rect 8927 6056 9113 6064
rect 9147 6056 9173 6064
rect 9387 6056 9633 6064
rect 10267 6056 10653 6064
rect 10987 6056 11013 6064
rect 11027 6056 11273 6064
rect 787 6036 933 6044
rect 967 6036 4093 6044
rect 4207 6036 4873 6044
rect 5987 6036 6533 6044
rect 6947 6036 7873 6044
rect 8147 6036 8393 6044
rect 8647 6036 8853 6044
rect 8907 6036 8933 6044
rect 9307 6036 9613 6044
rect 9627 6036 9813 6044
rect 9887 6036 11033 6044
rect 1647 6016 1673 6024
rect 1767 6016 1813 6024
rect 2627 6016 2653 6024
rect 2747 6016 2813 6024
rect 3307 6016 3713 6024
rect 5387 6016 6853 6024
rect 7207 6016 7353 6024
rect 8287 6016 8393 6024
rect 8607 6016 8873 6024
rect 1907 5996 1933 6004
rect 1956 5996 3293 6004
rect 1587 5976 1833 5984
rect 1956 5984 1964 5996
rect 3307 5996 4113 6004
rect 4136 5996 4733 6004
rect 1847 5976 1964 5984
rect 3207 5976 3893 5984
rect 4136 5984 4144 5996
rect 4747 5996 5273 6004
rect 6347 5996 6373 6004
rect 6587 5996 7493 6004
rect 7567 5996 10333 6004
rect 3907 5976 4144 5984
rect 4767 5976 5733 5984
rect 5747 5976 5813 5984
rect 6107 5976 6453 5984
rect 6667 5976 7173 5984
rect 7367 5976 7413 5984
rect 7587 5976 7613 5984
rect 8947 5976 11293 5984
rect 1567 5956 1993 5964
rect 2067 5956 2373 5964
rect 2387 5956 2893 5964
rect 3387 5956 4273 5964
rect 4387 5956 4533 5964
rect 4707 5956 5273 5964
rect 6707 5956 7013 5964
rect 7707 5956 8353 5964
rect 9127 5956 9793 5964
rect -24 5936 953 5944
rect 1387 5936 1873 5944
rect 2167 5936 2293 5944
rect 2307 5936 2313 5944
rect 2327 5936 2853 5944
rect 2867 5936 3353 5944
rect 4107 5936 4573 5944
rect 5127 5936 5453 5944
rect 5727 5936 6353 5944
rect 6787 5936 6793 5944
rect 6807 5936 6873 5944
rect 6907 5936 7033 5944
rect 7627 5936 7713 5944
rect 7847 5936 8133 5944
rect 8287 5936 8653 5944
rect 8667 5936 8933 5944
rect 8967 5936 9313 5944
rect 9347 5936 9553 5944
rect 9687 5936 10093 5944
rect 10187 5936 10513 5944
rect 10707 5936 11033 5944
rect 387 5916 393 5924
rect 407 5916 593 5924
rect 1107 5916 1173 5924
rect 1907 5916 2113 5924
rect 2367 5916 2633 5924
rect 3027 5916 3233 5924
rect 3527 5916 3633 5924
rect 3707 5916 3853 5924
rect 3887 5916 4793 5924
rect 4887 5916 5793 5924
rect 6547 5916 6993 5924
rect 7747 5916 7833 5924
rect 8027 5916 8173 5924
rect 8487 5916 8613 5924
rect 8807 5916 8833 5924
rect 8856 5916 8973 5924
rect 8856 5907 8864 5916
rect 8987 5916 9113 5924
rect 9167 5916 9353 5924
rect 9847 5916 10013 5924
rect 10127 5916 10313 5924
rect 10927 5916 10993 5924
rect 527 5896 573 5904
rect 787 5896 893 5904
rect 1287 5896 2133 5904
rect 2147 5896 2333 5904
rect 2807 5896 3313 5904
rect 3367 5896 3393 5904
rect 4567 5896 4593 5904
rect 4687 5896 4773 5904
rect 4827 5896 4853 5904
rect 5827 5896 5973 5904
rect 6007 5896 6173 5904
rect 6367 5896 6733 5904
rect 6787 5896 7613 5904
rect 8427 5896 8433 5904
rect 8447 5896 8633 5904
rect 8907 5896 9124 5904
rect 47 5876 933 5884
rect 947 5876 1193 5884
rect 1207 5876 1213 5884
rect 1227 5876 1353 5884
rect 3667 5876 3833 5884
rect 3847 5876 3993 5884
rect 4867 5876 5113 5884
rect 5127 5876 5253 5884
rect 5787 5876 5833 5884
rect 5847 5876 7693 5884
rect 7847 5876 8373 5884
rect 9116 5884 9124 5896
rect 9267 5896 10253 5904
rect 10787 5896 10813 5904
rect 11107 5896 11233 5904
rect 9116 5876 9133 5884
rect 9467 5876 10073 5884
rect 10087 5876 10133 5884
rect 10587 5876 10793 5884
rect 11227 5876 11253 5884
rect 1527 5856 1553 5864
rect 1567 5856 1853 5864
rect 1867 5856 2593 5864
rect 4407 5856 4693 5864
rect 4707 5856 6013 5864
rect 6067 5856 7013 5864
rect 7047 5856 7053 5864
rect 7067 5856 7213 5864
rect 7227 5856 7933 5864
rect 9096 5864 9104 5873
rect 11276 5867 11284 5893
rect 9087 5856 9104 5864
rect 4447 5836 7053 5844
rect 7947 5836 9053 5844
rect 5207 5816 6224 5824
rect 1647 5796 1813 5804
rect 1827 5796 2073 5804
rect 3547 5796 5793 5804
rect 6216 5804 6224 5816
rect 6807 5816 7913 5824
rect 8727 5816 10153 5824
rect 6216 5796 7033 5804
rect 7207 5796 7313 5804
rect 7747 5796 7753 5804
rect 7767 5796 11213 5804
rect 3367 5776 5233 5784
rect 5247 5776 5513 5784
rect 6047 5776 6713 5784
rect 6747 5776 6953 5784
rect 6987 5776 7013 5784
rect 7087 5776 7353 5784
rect 8507 5776 10473 5784
rect 2627 5756 5853 5764
rect 5987 5756 6473 5764
rect 6527 5756 6673 5764
rect 6687 5756 6973 5764
rect 6987 5756 7513 5764
rect 5607 5736 5753 5744
rect 6507 5736 6693 5744
rect 6727 5736 7673 5744
rect 7807 5736 10033 5744
rect 2507 5716 3593 5724
rect 3967 5716 4053 5724
rect 5007 5716 5293 5724
rect 5587 5716 6353 5724
rect 7507 5716 7853 5724
rect 8087 5716 8353 5724
rect 8447 5716 10233 5724
rect 10247 5716 10773 5724
rect 10787 5716 10893 5724
rect 2367 5696 2873 5704
rect 2887 5696 3733 5704
rect 4247 5696 4333 5704
rect 4807 5696 6033 5704
rect 8047 5696 8153 5704
rect 8747 5696 8813 5704
rect 9787 5696 10333 5704
rect 2576 5676 3153 5684
rect 2576 5667 2584 5676
rect 3747 5676 3913 5684
rect 4407 5676 4553 5684
rect 4567 5676 5073 5684
rect 5087 5676 5933 5684
rect 6027 5676 7773 5684
rect 7787 5676 8073 5684
rect 8107 5676 8433 5684
rect 9947 5676 10193 5684
rect 10667 5676 11013 5684
rect 467 5656 473 5664
rect 487 5656 633 5664
rect 687 5656 1013 5664
rect 1027 5656 1653 5664
rect 3127 5656 3473 5664
rect 3807 5656 5193 5664
rect 5487 5656 5573 5664
rect 5627 5656 5953 5664
rect 5967 5656 6233 5664
rect 6567 5656 6613 5664
rect 6627 5656 6913 5664
rect 7336 5656 7453 5664
rect 7336 5647 7344 5656
rect 7467 5656 7904 5664
rect 947 5636 1233 5644
rect 1547 5636 1593 5644
rect 1667 5636 1853 5644
rect 1947 5636 2033 5644
rect 2787 5636 2813 5644
rect 2867 5636 2933 5644
rect 3027 5636 3113 5644
rect 3127 5636 3613 5644
rect 3627 5636 3853 5644
rect 3867 5636 4353 5644
rect 4967 5636 5693 5644
rect 5727 5636 5753 5644
rect 5887 5636 5913 5644
rect 5947 5636 6793 5644
rect 7447 5636 7593 5644
rect 7607 5636 7633 5644
rect 7896 5644 7904 5656
rect 7927 5656 8013 5664
rect 8027 5656 8753 5664
rect 8767 5656 8833 5664
rect 9687 5656 9713 5664
rect 10327 5656 10513 5664
rect 10747 5656 11133 5664
rect 11167 5656 11213 5664
rect 11276 5664 11284 5673
rect 11267 5656 11284 5664
rect 7896 5636 8493 5644
rect 9227 5636 9293 5644
rect 9487 5636 9573 5644
rect 9976 5636 10013 5644
rect 367 5616 853 5624
rect 1847 5616 2593 5624
rect 2847 5616 3053 5624
rect 3307 5616 3593 5624
rect 3647 5616 3793 5624
rect 3927 5616 3953 5624
rect 4047 5616 4333 5624
rect 5207 5616 5733 5624
rect 6627 5616 6653 5624
rect 6767 5616 6773 5624
rect 6787 5616 7033 5624
rect 7667 5616 7853 5624
rect 7876 5624 7884 5633
rect 7876 5616 7953 5624
rect 8987 5616 9153 5624
rect 9176 5624 9184 5633
rect 9176 5616 9213 5624
rect 9436 5624 9444 5633
rect 9436 5616 9693 5624
rect 9976 5624 9984 5636
rect 10287 5636 10313 5644
rect 10347 5636 10493 5644
rect 10507 5636 10713 5644
rect 10767 5636 10813 5644
rect 10987 5636 11113 5644
rect 9967 5616 9984 5624
rect 10007 5616 10113 5624
rect 10167 5616 10253 5624
rect 11236 5624 11244 5633
rect 10827 5616 11244 5624
rect 2027 5596 2553 5604
rect 2707 5596 2973 5604
rect 2987 5596 3133 5604
rect 3447 5596 3813 5604
rect 5067 5596 5213 5604
rect 5607 5596 5673 5604
rect 6187 5596 6533 5604
rect 6727 5596 6933 5604
rect 7407 5596 7613 5604
rect 7707 5596 8113 5604
rect 8387 5596 8933 5604
rect 9027 5596 9193 5604
rect 9247 5596 9453 5604
rect 9987 5596 10293 5604
rect 10307 5596 10653 5604
rect 10907 5596 10993 5604
rect 1107 5576 1153 5584
rect 1167 5576 1333 5584
rect 1347 5576 2833 5584
rect 2847 5576 2913 5584
rect 3247 5576 3253 5584
rect 3267 5576 3293 5584
rect 3307 5576 3593 5584
rect 3767 5576 5933 5584
rect 6107 5576 6193 5584
rect 6207 5576 7433 5584
rect 9167 5576 9413 5584
rect 9447 5576 9493 5584
rect 9507 5576 9673 5584
rect 9687 5576 9713 5584
rect 1767 5556 1793 5564
rect 2207 5556 2413 5564
rect 2787 5556 3033 5564
rect 3067 5556 3313 5564
rect 4167 5556 4573 5564
rect 4827 5556 5244 5564
rect 1367 5536 1413 5544
rect 3187 5536 3573 5544
rect 3947 5536 4313 5544
rect 5236 5544 5244 5556
rect 5687 5556 5813 5564
rect 6307 5556 6813 5564
rect 6967 5556 7013 5564
rect 7127 5556 7293 5564
rect 7307 5556 7373 5564
rect 7387 5556 8573 5564
rect 5236 5536 6333 5544
rect 6427 5536 7993 5544
rect 8647 5536 8733 5544
rect 927 5516 1013 5524
rect 2807 5516 3213 5524
rect 3227 5516 3393 5524
rect 3407 5516 3893 5524
rect 4467 5516 4573 5524
rect 5207 5516 6113 5524
rect 6407 5516 6573 5524
rect 6627 5516 6833 5524
rect 7447 5516 7533 5524
rect 7907 5516 8153 5524
rect 8167 5516 8493 5524
rect 8507 5516 8693 5524
rect 9127 5516 10213 5524
rect 10227 5516 10453 5524
rect 2787 5496 2933 5504
rect 3267 5496 3513 5504
rect 4767 5496 6073 5504
rect 6647 5496 6693 5504
rect 7847 5496 7893 5504
rect 9307 5496 9733 5504
rect 10267 5496 10773 5504
rect 227 5476 433 5484
rect 447 5476 1453 5484
rect 2767 5476 3153 5484
rect 4147 5476 4413 5484
rect 4847 5476 4893 5484
rect 4927 5476 5153 5484
rect 5167 5476 5733 5484
rect 5747 5476 6133 5484
rect 6907 5476 7593 5484
rect 7607 5476 7933 5484
rect 9007 5476 9333 5484
rect 10036 5476 10233 5484
rect 287 5456 453 5464
rect 567 5456 593 5464
rect 607 5456 913 5464
rect 927 5456 1213 5464
rect 1467 5456 1613 5464
rect 1647 5456 1693 5464
rect 2927 5456 3313 5464
rect 3327 5456 3373 5464
rect 3647 5456 3833 5464
rect 5387 5456 5553 5464
rect 5887 5456 6213 5464
rect 7027 5456 7073 5464
rect 7287 5456 7533 5464
rect 7547 5456 7873 5464
rect 7887 5456 8273 5464
rect 8307 5456 8373 5464
rect 10036 5464 10044 5476
rect 10587 5476 10833 5484
rect 10847 5476 10953 5484
rect 9327 5456 10044 5464
rect 10067 5456 10353 5464
rect 11007 5456 11253 5464
rect 907 5436 953 5444
rect 1627 5436 1673 5444
rect 1727 5436 1873 5444
rect 2387 5436 2453 5444
rect 2587 5436 2653 5444
rect 2907 5436 2973 5444
rect 3607 5436 3993 5444
rect 4127 5436 4173 5444
rect 4227 5436 4253 5444
rect 4267 5436 4313 5444
rect 4647 5436 5184 5444
rect 5176 5427 5184 5436
rect 6067 5436 7153 5444
rect 7327 5436 7573 5444
rect 7847 5436 7993 5444
rect 8007 5436 8473 5444
rect 8667 5436 8873 5444
rect 8887 5436 9053 5444
rect 9747 5436 10273 5444
rect 10427 5436 11033 5444
rect 207 5416 273 5424
rect 987 5416 1173 5424
rect 1447 5416 1633 5424
rect 1867 5416 1933 5424
rect 1947 5416 1973 5424
rect 2167 5416 2393 5424
rect 2447 5416 2493 5424
rect 2687 5416 2773 5424
rect 2867 5416 2953 5424
rect 3047 5416 3193 5424
rect 3207 5416 3413 5424
rect 3467 5416 3513 5424
rect 3807 5416 3953 5424
rect 4007 5416 4273 5424
rect 4287 5416 4593 5424
rect 4687 5416 4853 5424
rect 4887 5416 4913 5424
rect 5047 5416 5133 5424
rect 5227 5416 5833 5424
rect 6167 5416 6453 5424
rect 7887 5416 7973 5424
rect 8107 5416 8153 5424
rect 8407 5416 9073 5424
rect 9087 5416 9493 5424
rect 9547 5416 9733 5424
rect 9807 5416 9993 5424
rect 10947 5416 11073 5424
rect 11087 5416 11273 5424
rect 696 5364 704 5413
rect 727 5396 793 5404
rect 947 5396 1473 5404
rect 1487 5396 1573 5404
rect 1847 5396 1913 5404
rect 1967 5396 2013 5404
rect 2047 5396 2133 5404
rect 2287 5396 2713 5404
rect 2727 5396 2893 5404
rect 3747 5396 4253 5404
rect 4967 5396 5073 5404
rect 6036 5404 6044 5413
rect 6036 5396 6053 5404
rect 6347 5396 6493 5404
rect 6787 5396 6953 5404
rect 6967 5396 7033 5404
rect 7527 5396 7693 5404
rect 7707 5396 7713 5404
rect 7767 5396 8013 5404
rect 9467 5396 9513 5404
rect 10047 5396 10293 5404
rect 11327 5396 11404 5404
rect 1227 5376 2173 5384
rect 2187 5376 2373 5384
rect 3427 5376 3913 5384
rect 4207 5376 4613 5384
rect 4747 5376 5433 5384
rect 5667 5376 6373 5384
rect 6387 5376 6733 5384
rect 6807 5376 6973 5384
rect 6996 5376 7893 5384
rect 687 5356 704 5364
rect 967 5356 1153 5364
rect 1167 5356 1873 5364
rect 4867 5356 5053 5364
rect 5887 5356 5973 5364
rect 5987 5356 6153 5364
rect 6996 5364 7004 5376
rect 8027 5376 8053 5384
rect 10067 5376 10113 5384
rect 11056 5384 11064 5393
rect 11056 5376 11073 5384
rect 11267 5376 11333 5384
rect 6327 5356 7004 5364
rect 7267 5356 7453 5364
rect 7627 5356 8553 5364
rect 9407 5356 9513 5364
rect 4887 5336 4933 5344
rect 5527 5336 6813 5344
rect 6927 5336 6993 5344
rect 7007 5336 9853 5344
rect 10147 5336 10253 5344
rect 4227 5316 8333 5324
rect 4907 5296 5613 5304
rect 5927 5296 7273 5304
rect 547 5276 1013 5284
rect 5107 5276 5173 5284
rect 5636 5276 5753 5284
rect 1007 5256 1113 5264
rect 5636 5264 5644 5276
rect 5767 5276 6013 5284
rect 6267 5276 6533 5284
rect 7487 5276 8453 5284
rect 3487 5256 5644 5264
rect 7556 5256 10913 5264
rect 227 5156 393 5164
rect 487 5156 513 5164
rect 187 5136 453 5144
rect 427 5116 573 5124
rect 636 5087 644 5253
rect 4167 5236 4813 5244
rect 7556 5244 7564 5256
rect 4987 5236 7564 5244
rect 7587 5236 8373 5244
rect 8387 5236 9693 5244
rect 2227 5216 7433 5224
rect 7647 5216 8113 5224
rect 9067 5216 9133 5224
rect 3687 5196 3753 5204
rect 4627 5196 5353 5204
rect 6387 5196 6473 5204
rect 6707 5196 6833 5204
rect 7207 5196 9433 5204
rect 9547 5196 9653 5204
rect 10547 5196 10633 5204
rect 10687 5196 10713 5204
rect 10867 5196 10953 5204
rect 1947 5176 2133 5184
rect 2907 5176 3453 5184
rect 3467 5176 3593 5184
rect 3607 5176 3633 5184
rect 5116 5176 5213 5184
rect 887 5156 1353 5164
rect 1547 5156 1673 5164
rect 1727 5156 1793 5164
rect 2007 5156 2113 5164
rect 2727 5156 2804 5164
rect 1467 5136 1653 5144
rect 1707 5136 2193 5144
rect 2467 5136 2653 5144
rect 2796 5144 2804 5156
rect 2907 5156 2933 5164
rect 3347 5156 3393 5164
rect 3627 5156 3773 5164
rect 4396 5156 4613 5164
rect 4396 5147 4404 5156
rect 4627 5156 4733 5164
rect 4896 5147 4904 5173
rect 5116 5167 5124 5176
rect 5247 5176 5413 5184
rect 5427 5176 5613 5184
rect 5627 5176 5873 5184
rect 5987 5176 6093 5184
rect 6267 5176 7553 5184
rect 7667 5176 7853 5184
rect 7936 5176 8213 5184
rect 5167 5156 5213 5164
rect 6027 5156 6073 5164
rect 6447 5156 6473 5164
rect 6827 5156 6953 5164
rect 7007 5156 7033 5164
rect 7247 5156 7353 5164
rect 7367 5156 7413 5164
rect 7936 5164 7944 5176
rect 8727 5176 9493 5184
rect 9567 5176 9684 5184
rect 9676 5167 9684 5176
rect 9927 5176 10153 5184
rect 10467 5176 11133 5184
rect 7467 5156 7944 5164
rect 7967 5156 8053 5164
rect 8447 5156 8513 5164
rect 8567 5156 9153 5164
rect 9207 5156 9373 5164
rect 9567 5156 9633 5164
rect 9896 5164 9904 5173
rect 9876 5156 10113 5164
rect 2796 5136 2913 5144
rect 2927 5136 2973 5144
rect 2987 5136 3013 5144
rect 3087 5136 3293 5144
rect 3447 5136 3513 5144
rect 4307 5136 4353 5144
rect 4847 5136 4873 5144
rect 4916 5144 4924 5153
rect 4916 5136 5433 5144
rect 6007 5136 6053 5144
rect 6107 5136 6273 5144
rect 6307 5136 6713 5144
rect 7027 5136 7173 5144
rect 7287 5136 7933 5144
rect 8467 5136 8493 5144
rect 8507 5136 8673 5144
rect 8987 5136 9133 5144
rect 9876 5144 9884 5156
rect 10147 5156 10493 5164
rect 10887 5156 10973 5164
rect 11167 5156 11213 5164
rect 9607 5136 9884 5144
rect 10287 5136 10393 5144
rect 10487 5136 10793 5144
rect 10807 5136 10893 5144
rect 707 5116 893 5124
rect 1187 5116 1493 5124
rect 2347 5116 2693 5124
rect 3307 5116 3893 5124
rect 4387 5116 4413 5124
rect 5727 5116 6053 5124
rect 6467 5116 6893 5124
rect 7147 5116 7173 5124
rect 7227 5116 7433 5124
rect 8167 5116 8693 5124
rect 8967 5116 9173 5124
rect 9507 5116 9613 5124
rect 9827 5116 9873 5124
rect 10707 5116 11093 5124
rect 1367 5096 2053 5104
rect 2067 5096 2373 5104
rect 3047 5096 3153 5104
rect 4467 5096 4973 5104
rect 5967 5096 6493 5104
rect 6527 5096 6973 5104
rect 7867 5096 7913 5104
rect 7927 5096 8413 5104
rect 8427 5096 8593 5104
rect 8927 5096 8993 5104
rect 10867 5096 11153 5104
rect 1327 5076 1853 5084
rect 1867 5076 1933 5084
rect 3827 5076 4053 5084
rect 4487 5076 4593 5084
rect 5227 5076 5613 5084
rect 5627 5076 5813 5084
rect 8207 5076 8273 5084
rect 8407 5076 9133 5084
rect 9507 5076 9833 5084
rect 507 5056 533 5064
rect 547 5056 993 5064
rect 1267 5056 4113 5064
rect 5507 5056 5973 5064
rect 5987 5056 6213 5064
rect 7387 5056 7673 5064
rect 8247 5056 8933 5064
rect 9147 5056 10933 5064
rect 247 5036 413 5044
rect 427 5036 1253 5044
rect 3187 5036 3373 5044
rect 3567 5036 4153 5044
rect 4167 5036 4213 5044
rect 4327 5036 4493 5044
rect 4527 5036 5013 5044
rect 5067 5036 5133 5044
rect 5787 5036 5813 5044
rect 7447 5036 8353 5044
rect 8587 5036 10093 5044
rect 27 5016 1773 5024
rect 1967 5016 3693 5024
rect 4327 5016 4593 5024
rect 5547 5016 7093 5024
rect 7667 5016 8653 5024
rect 8667 5016 10533 5024
rect 3027 4996 3653 5004
rect 4147 4996 4333 5004
rect 5347 4996 5513 5004
rect 5607 4996 6453 5004
rect 7047 4996 9413 5004
rect 9887 4996 10333 5004
rect 10387 4996 10613 5004
rect 647 4976 664 4984
rect -24 4956 13 4964
rect 447 4956 473 4964
rect 487 4956 633 4964
rect 656 4924 664 4976
rect 967 4976 1193 4984
rect 1427 4976 1453 4984
rect 1527 4976 1693 4984
rect 2907 4976 3453 4984
rect 3467 4976 3553 4984
rect 4087 4976 4253 4984
rect 4587 4976 5833 4984
rect 6467 4976 6493 4984
rect 6547 4976 8393 4984
rect 9647 4976 9973 4984
rect 10127 4976 10353 4984
rect 10827 4976 11273 4984
rect 11116 4967 11124 4976
rect 727 4956 833 4964
rect 1147 4956 1213 4964
rect 1427 4956 1613 4964
rect 1627 4956 1713 4964
rect 1787 4956 2433 4964
rect 2447 4956 2713 4964
rect 2727 4956 2793 4964
rect 2807 4956 2893 4964
rect 3007 4956 3113 4964
rect 3187 4956 3413 4964
rect 3607 4956 3693 4964
rect 3707 4956 3993 4964
rect 4127 4956 4573 4964
rect 4647 4956 6213 4964
rect 6267 4956 6473 4964
rect 7147 4956 7393 4964
rect 7407 4956 7753 4964
rect 8187 4956 8413 4964
rect 8687 4956 8893 4964
rect 9787 4956 10153 4964
rect 707 4936 773 4944
rect 787 4936 933 4944
rect 1487 4936 1513 4944
rect 1707 4936 1833 4944
rect 1847 4936 1973 4944
rect 2667 4936 2873 4944
rect 2987 4936 3133 4944
rect 3687 4936 3873 4944
rect 3927 4936 4093 4944
rect 4107 4936 4193 4944
rect 5207 4936 5533 4944
rect 5547 4936 5893 4944
rect 5907 4936 5933 4944
rect 6067 4936 6233 4944
rect 6287 4936 6593 4944
rect 6747 4936 6953 4944
rect 7687 4936 7733 4944
rect 8527 4936 8633 4944
rect 8687 4936 8753 4944
rect 8767 4936 9433 4944
rect 9807 4936 9873 4944
rect 9927 4936 9953 4944
rect 10067 4936 10093 4944
rect 10147 4936 10193 4944
rect 10207 4936 10313 4944
rect 10747 4936 11053 4944
rect 656 4916 673 4924
rect 827 4916 973 4924
rect 987 4916 1033 4924
rect 1447 4916 1973 4924
rect 2047 4916 2133 4924
rect 2147 4916 2473 4924
rect 3707 4916 3793 4924
rect 3887 4916 4613 4924
rect 5527 4916 5573 4924
rect 5907 4916 5993 4924
rect 6987 4916 7073 4924
rect 7207 4916 7533 4924
rect 7867 4916 7893 4924
rect 7947 4916 8053 4924
rect 9127 4916 9353 4924
rect 9407 4916 9633 4924
rect 9647 4916 9773 4924
rect 9907 4916 9933 4924
rect 10147 4916 10173 4924
rect 10687 4916 11073 4924
rect 867 4896 2373 4904
rect 4427 4896 4713 4904
rect 5647 4896 6533 4904
rect 6947 4896 8933 4904
rect 9167 4896 9313 4904
rect 9567 4896 9613 4904
rect 9867 4896 10593 4904
rect 10607 4896 10913 4904
rect 2467 4876 2693 4884
rect 2707 4876 2953 4884
rect 2967 4876 3193 4884
rect 3207 4876 3433 4884
rect 3447 4876 3593 4884
rect 3607 4876 4133 4884
rect 4147 4876 4433 4884
rect 5807 4876 7193 4884
rect 7767 4876 9593 4884
rect 667 4856 1733 4864
rect 1767 4856 4753 4864
rect 4907 4856 4953 4864
rect 4967 4856 5413 4864
rect 7647 4856 8113 4864
rect 4607 4836 9273 4844
rect 947 4816 1053 4824
rect 4307 4816 5953 4824
rect 9487 4816 10053 4824
rect 227 4796 413 4804
rect 2387 4796 4233 4804
rect 4247 4796 4953 4804
rect 4967 4796 5693 4804
rect 5727 4796 8313 4804
rect 8947 4796 9673 4804
rect 9727 4796 9833 4804
rect 4327 4776 4833 4784
rect 9667 4776 10053 4784
rect 2116 4756 2173 4764
rect 2116 4747 2124 4756
rect 3147 4756 3873 4764
rect 5027 4756 7793 4764
rect 8607 4756 9193 4764
rect 9287 4756 9793 4764
rect 2747 4736 3133 4744
rect 3147 4736 4653 4744
rect 5427 4736 5773 4744
rect 5787 4736 6253 4744
rect 6267 4736 6793 4744
rect 7807 4736 9213 4744
rect 487 4716 553 4724
rect 767 4716 853 4724
rect 1587 4716 1933 4724
rect 3347 4716 3393 4724
rect 3447 4716 4773 4724
rect 5707 4716 5733 4724
rect 5787 4716 6193 4724
rect 6667 4716 6733 4724
rect 7947 4716 7973 4724
rect 8067 4716 8773 4724
rect 407 4696 1553 4704
rect 1567 4696 1933 4704
rect 2027 4696 2653 4704
rect 2667 4696 3053 4704
rect 3187 4696 3333 4704
rect 3767 4696 3933 4704
rect 3947 4696 4633 4704
rect 4787 4696 5053 4704
rect 5067 4696 5553 4704
rect 5847 4696 6693 4704
rect 6987 4696 7033 4704
rect 7407 4696 7813 4704
rect 7827 4696 7873 4704
rect 7927 4696 8013 4704
rect 8047 4696 8073 4704
rect 8127 4696 8213 4704
rect 8647 4696 9653 4704
rect 9947 4696 10313 4704
rect 10827 4696 11293 4704
rect 187 4676 453 4684
rect 527 4676 1633 4684
rect 1687 4676 1793 4684
rect 1807 4676 1993 4684
rect 2107 4676 2613 4684
rect 2907 4676 3093 4684
rect 3987 4676 4073 4684
rect 5547 4676 5733 4684
rect 5887 4676 5913 4684
rect 6507 4676 6713 4684
rect 7416 4676 7573 4684
rect 7416 4667 7424 4676
rect 7767 4676 7953 4684
rect 8047 4676 8193 4684
rect 8247 4676 8533 4684
rect 8547 4676 8653 4684
rect 8887 4676 9364 4684
rect 247 4656 413 4664
rect 427 4656 593 4664
rect 1347 4656 1393 4664
rect 1447 4656 1613 4664
rect 1667 4656 1893 4664
rect 1967 4656 1973 4664
rect 1987 4656 2493 4664
rect 2507 4656 2673 4664
rect 3627 4656 3833 4664
rect 3907 4656 4413 4664
rect 4987 4656 5213 4664
rect 5056 4647 5064 4656
rect 5547 4656 5673 4664
rect 6327 4656 6513 4664
rect 6747 4656 6873 4664
rect 7007 4656 7013 4664
rect 7027 4656 7193 4664
rect 7207 4656 7393 4664
rect 7467 4656 7793 4664
rect 8167 4656 8413 4664
rect 8467 4656 8513 4664
rect 8987 4656 9093 4664
rect 9147 4656 9293 4664
rect 9356 4664 9364 4676
rect 9727 4676 9773 4684
rect 9827 4676 9853 4684
rect 10027 4676 10193 4684
rect 10347 4676 10413 4684
rect 10927 4676 11013 4684
rect 9356 4656 9373 4664
rect 9567 4656 9693 4664
rect 9807 4656 9933 4664
rect 9967 4656 10033 4664
rect 10127 4656 10293 4664
rect 10327 4656 10433 4664
rect 10776 4664 10784 4673
rect 10776 4656 10793 4664
rect 11047 4656 11093 4664
rect 367 4636 853 4644
rect 867 4636 873 4644
rect 1047 4636 1133 4644
rect 1927 4636 2253 4644
rect 3847 4636 4253 4644
rect 4267 4636 4273 4644
rect 4387 4636 4553 4644
rect 5287 4636 5493 4644
rect 5587 4636 5793 4644
rect 6107 4636 6473 4644
rect 7447 4636 7633 4644
rect 7687 4636 7733 4644
rect 8027 4636 8253 4644
rect 8287 4636 8433 4644
rect 8887 4636 9033 4644
rect 9167 4636 9333 4644
rect 9467 4636 9553 4644
rect 10547 4636 10993 4644
rect 11007 4636 11113 4644
rect 1227 4616 2393 4624
rect 2407 4616 2613 4624
rect 3967 4616 4093 4624
rect 5047 4616 5093 4624
rect 5107 4616 5293 4624
rect 6387 4616 6453 4624
rect 6547 4616 7693 4624
rect 7907 4616 8473 4624
rect 8487 4616 8733 4624
rect 8747 4616 9893 4624
rect 9907 4616 10873 4624
rect 10887 4616 11193 4624
rect 727 4596 853 4604
rect 4047 4596 4693 4604
rect 5047 4596 5253 4604
rect 6167 4596 6333 4604
rect 6447 4596 6653 4604
rect 6867 4596 7493 4604
rect 8327 4596 8693 4604
rect 8707 4596 9753 4604
rect 10307 4596 10733 4604
rect 10767 4596 11333 4604
rect 2847 4576 4893 4584
rect 5467 4576 5513 4584
rect 5567 4576 10673 4584
rect 10907 4576 11053 4584
rect 11067 4576 11273 4584
rect 2167 4556 2373 4564
rect 2687 4556 3113 4564
rect 3187 4556 3313 4564
rect 3327 4556 4153 4564
rect 4247 4556 4913 4564
rect 4927 4556 5953 4564
rect 6027 4556 6873 4564
rect 6887 4556 7573 4564
rect 8867 4556 8993 4564
rect 9227 4556 9333 4564
rect 10567 4556 10773 4564
rect 11007 4556 11133 4564
rect 1927 4536 4613 4544
rect 5467 4536 5853 4544
rect 8847 4536 9473 4544
rect 9687 4536 10493 4544
rect 2827 4516 3353 4524
rect 4387 4516 4413 4524
rect 5807 4516 6073 4524
rect 6087 4516 6313 4524
rect 7187 4516 7753 4524
rect 7947 4516 7973 4524
rect 8227 4516 8473 4524
rect 8487 4516 8953 4524
rect 9247 4516 9933 4524
rect 10507 4516 10913 4524
rect 10927 4516 11153 4524
rect 1067 4496 1213 4504
rect 1387 4496 1433 4504
rect 1447 4496 1793 4504
rect 1807 4496 2053 4504
rect 2087 4496 2253 4504
rect 2447 4496 2633 4504
rect 2727 4496 2873 4504
rect 2887 4496 2933 4504
rect 2947 4496 3093 4504
rect 3107 4496 3153 4504
rect 3347 4496 3833 4504
rect 4647 4496 4853 4504
rect 5087 4496 5233 4504
rect 5667 4496 5893 4504
rect 6247 4496 6573 4504
rect 6647 4496 7073 4504
rect 7527 4496 7704 4504
rect 507 4476 513 4484
rect 527 4476 673 4484
rect 707 4476 913 4484
rect 927 4476 1313 4484
rect 1407 4476 1593 4484
rect 1627 4476 1833 4484
rect 2647 4476 2833 4484
rect 2947 4476 3053 4484
rect 3807 4476 3853 4484
rect 4007 4476 4093 4484
rect 4107 4476 4124 4484
rect 467 4456 553 4464
rect 567 4456 733 4464
rect 1147 4456 1233 4464
rect 1247 4456 1573 4464
rect 1587 4456 2013 4464
rect 2127 4456 2173 4464
rect 2867 4456 2993 4464
rect 3127 4456 3673 4464
rect 4116 4464 4124 4476
rect 4147 4476 4173 4484
rect 4207 4476 4413 4484
rect 4667 4476 4693 4484
rect 5367 4476 5773 4484
rect 5927 4476 6113 4484
rect 6207 4476 6353 4484
rect 7067 4476 7193 4484
rect 7567 4476 7653 4484
rect 7667 4476 7673 4484
rect 7696 4484 7704 4496
rect 7747 4496 8433 4504
rect 8447 4496 8573 4504
rect 8627 4496 8673 4504
rect 8687 4496 9373 4504
rect 9447 4496 9453 4504
rect 9607 4496 10173 4504
rect 10187 4496 10573 4504
rect 11147 4496 11333 4504
rect 7696 4476 8013 4484
rect 8167 4476 8193 4484
rect 8467 4476 8693 4484
rect 9027 4476 9413 4484
rect 9727 4476 9753 4484
rect 9887 4476 10373 4484
rect 10387 4476 10453 4484
rect 10787 4476 10913 4484
rect 4116 4456 4353 4464
rect 4487 4456 4533 4464
rect 4547 4456 4973 4464
rect 5267 4456 5353 4464
rect 5947 4456 6093 4464
rect 6147 4456 6353 4464
rect 6587 4456 7373 4464
rect 7547 4456 7753 4464
rect 7767 4456 7953 4464
rect 7987 4456 8233 4464
rect 8727 4456 8753 4464
rect 8907 4456 8933 4464
rect 9047 4456 9193 4464
rect 9307 4456 9693 4464
rect 10447 4456 10513 4464
rect 10607 4456 10653 4464
rect 47 4436 53 4444
rect 67 4436 713 4444
rect 907 4436 953 4444
rect 967 4436 1113 4444
rect 1127 4436 1353 4444
rect 2787 4436 3053 4444
rect 3087 4436 3193 4444
rect 3207 4436 3493 4444
rect 3927 4436 4113 4444
rect 6387 4436 6413 4444
rect 6987 4436 7053 4444
rect 7067 4436 7133 4444
rect 7147 4436 7273 4444
rect 7347 4436 7733 4444
rect 7787 4436 7973 4444
rect 8027 4436 8173 4444
rect 8527 4436 9173 4444
rect 9376 4436 9433 4444
rect 427 4416 933 4424
rect 4707 4416 4913 4424
rect 4927 4416 5093 4424
rect 6187 4416 6613 4424
rect 7047 4416 7073 4424
rect 7667 4416 7853 4424
rect 7967 4416 8153 4424
rect 8767 4416 8973 4424
rect 9376 4424 9384 4436
rect 9527 4436 9673 4444
rect 9687 4436 9873 4444
rect 9967 4436 10073 4444
rect 10207 4436 10393 4444
rect 8987 4416 9384 4424
rect 9407 4416 9433 4424
rect 9667 4416 9713 4424
rect 9727 4416 10673 4424
rect 10687 4416 10793 4424
rect 847 4396 1153 4404
rect 1167 4396 1633 4404
rect 1647 4396 2033 4404
rect 4887 4396 7644 4404
rect 827 4376 1813 4384
rect 1827 4376 2073 4384
rect 2087 4376 2113 4384
rect 2607 4376 5513 4384
rect 5987 4376 7613 4384
rect 7636 4384 7644 4396
rect 7787 4396 7813 4404
rect 8187 4396 8793 4404
rect 9707 4396 9753 4404
rect 9807 4396 10073 4404
rect 10087 4396 10153 4404
rect 10167 4396 10633 4404
rect 10647 4396 10733 4404
rect 7636 4376 8064 4384
rect 6787 4356 8033 4364
rect 8056 4364 8064 4376
rect 8147 4376 8893 4384
rect 9327 4376 11273 4384
rect 8056 4356 8413 4364
rect 9767 4356 10393 4364
rect 5187 4336 5633 4344
rect 2387 4316 7713 4324
rect 8007 4316 8193 4324
rect 8207 4316 9313 4324
rect 2627 4296 3073 4304
rect 3087 4296 3473 4304
rect 4687 4296 5073 4304
rect 5227 4296 5433 4304
rect 7407 4296 8233 4304
rect 8247 4296 8613 4304
rect 9387 4296 10053 4304
rect 10067 4296 10333 4304
rect 2367 4276 2453 4284
rect 2547 4276 3733 4284
rect 4447 4276 5633 4284
rect 6527 4276 6553 4284
rect 6627 4276 7433 4284
rect 7707 4276 7753 4284
rect 8567 4276 8573 4284
rect 8587 4276 8693 4284
rect 8707 4276 9873 4284
rect 10267 4276 11053 4284
rect 2467 4256 2573 4264
rect 2927 4256 3313 4264
rect 3887 4256 4593 4264
rect 5827 4256 5873 4264
rect 6087 4256 6293 4264
rect 6307 4256 6793 4264
rect 7247 4256 7633 4264
rect 7647 4256 8313 4264
rect 8747 4256 9493 4264
rect 667 4236 913 4244
rect 947 4236 1133 4244
rect 2107 4236 2653 4244
rect 3567 4236 4453 4244
rect 5807 4236 7253 4244
rect 7707 4236 8813 4244
rect 9167 4236 9313 4244
rect 727 4216 993 4224
rect 1007 4216 1053 4224
rect 1427 4216 1593 4224
rect 1607 4216 1873 4224
rect 2556 4216 2933 4224
rect 2556 4207 2564 4216
rect 3247 4216 3513 4224
rect 4147 4216 4253 4224
rect 4287 4216 4393 4224
rect 4407 4216 4693 4224
rect 4707 4216 5093 4224
rect 5327 4216 5373 4224
rect 6296 4216 6333 4224
rect 247 4196 393 4204
rect 407 4196 933 4204
rect 2307 4196 2533 4204
rect 2667 4196 2713 4204
rect 2747 4196 2913 4204
rect 2947 4196 3273 4204
rect 3307 4196 3773 4204
rect 3867 4196 4433 4204
rect 4487 4196 4713 4204
rect 5847 4196 5933 4204
rect 5967 4196 6033 4204
rect 6296 4204 6304 4216
rect 6347 4216 6473 4224
rect 6487 4216 6593 4224
rect 6607 4216 6673 4224
rect 7287 4216 7413 4224
rect 7447 4216 7473 4224
rect 8367 4216 8813 4224
rect 9187 4216 9633 4224
rect 9647 4216 9753 4224
rect 9847 4216 9913 4224
rect 9947 4216 10373 4224
rect 10387 4216 10533 4224
rect 10667 4216 10813 4224
rect 11107 4216 11133 4224
rect 6047 4196 6304 4204
rect 6327 4196 6513 4204
rect 7267 4196 7693 4204
rect 7747 4196 7813 4204
rect 7827 4196 7933 4204
rect 7987 4196 8133 4204
rect 8327 4196 8433 4204
rect 8987 4196 9013 4204
rect 9127 4196 9193 4204
rect 9427 4196 9653 4204
rect 9887 4196 10733 4204
rect 10747 4196 10833 4204
rect 10947 4196 11113 4204
rect 207 4176 473 4184
rect 887 4176 1033 4184
rect 2087 4176 2253 4184
rect 2267 4176 2273 4184
rect 2296 4167 2304 4193
rect 3047 4176 3333 4184
rect 3727 4176 3873 4184
rect 3947 4176 3973 4184
rect 4467 4176 4793 4184
rect 5596 4184 5604 4193
rect 5387 4176 5613 4184
rect 5647 4176 6053 4184
rect 6107 4176 6613 4184
rect 7727 4176 8204 4184
rect 707 4156 813 4164
rect 1167 4156 1393 4164
rect 2327 4156 2913 4164
rect 3547 4156 3613 4164
rect 3627 4156 3913 4164
rect 3987 4156 5333 4164
rect 5867 4156 6373 4164
rect 6787 4156 6993 4164
rect 7027 4156 7073 4164
rect 7507 4156 7533 4164
rect 7556 4156 7893 4164
rect 367 4136 1333 4144
rect 2367 4136 3273 4144
rect 4367 4136 4893 4144
rect 4907 4136 5593 4144
rect 7556 4144 7564 4156
rect 7967 4156 8113 4164
rect 8196 4164 8204 4176
rect 8227 4176 8653 4184
rect 8727 4176 8893 4184
rect 8907 4176 8913 4184
rect 9167 4176 9393 4184
rect 9627 4176 9713 4184
rect 9827 4176 9933 4184
rect 10787 4176 10813 4184
rect 8196 4156 8393 4164
rect 8427 4156 8493 4164
rect 8687 4156 8853 4164
rect 8907 4156 9053 4164
rect 9107 4156 9173 4164
rect 9407 4156 9553 4164
rect 9627 4156 9673 4164
rect 9747 4156 9833 4164
rect 9867 4156 10093 4164
rect 10587 4156 10853 4164
rect 10867 4156 10913 4164
rect 10927 4156 10933 4164
rect 6347 4136 7564 4144
rect 7587 4136 8993 4144
rect 9167 4136 9273 4144
rect 9647 4136 9693 4144
rect 9707 4136 9733 4144
rect 9907 4136 9933 4144
rect 9947 4136 10173 4144
rect 10187 4136 10573 4144
rect 267 4116 393 4124
rect 1847 4116 2753 4124
rect 3707 4116 4713 4124
rect 6067 4116 6433 4124
rect 7047 4116 9133 4124
rect 10587 4116 10693 4124
rect 10707 4116 10793 4124
rect 1187 4096 1513 4104
rect 1887 4096 2993 4104
rect 6467 4096 7313 4104
rect 7527 4096 8333 4104
rect 8347 4096 8613 4104
rect 8647 4096 9513 4104
rect 9907 4096 9973 4104
rect 1247 4076 1433 4084
rect 1987 4076 2253 4084
rect 2267 4076 7733 4084
rect 8007 4076 10213 4084
rect 867 4056 1453 4064
rect 1467 4056 1693 4064
rect 2847 4056 3013 4064
rect 5827 4056 8733 4064
rect 9087 4056 9973 4064
rect 10687 4056 10813 4064
rect 10827 4056 10973 4064
rect 667 4036 993 4044
rect 2927 4036 3253 4044
rect 3267 4036 4164 4044
rect 627 4016 1953 4024
rect 2247 4016 2573 4024
rect 2627 4016 2713 4024
rect 2727 4016 2953 4024
rect 3727 4016 3953 4024
rect 4156 4024 4164 4036
rect 4187 4036 4913 4044
rect 5067 4036 6413 4044
rect 6427 4036 7593 4044
rect 7887 4036 8773 4044
rect 8867 4036 9053 4044
rect 9167 4036 9713 4044
rect 10467 4036 10553 4044
rect 10807 4036 10953 4044
rect 11027 4036 11213 4044
rect 4156 4016 4973 4024
rect 5267 4016 5273 4024
rect 5287 4016 5673 4024
rect 6647 4016 6673 4024
rect 6827 4016 6933 4024
rect 7007 4016 7133 4024
rect 7167 4016 7353 4024
rect 7367 4016 7473 4024
rect 7527 4016 8133 4024
rect 8167 4016 8333 4024
rect 8427 4016 8553 4024
rect 8627 4016 9073 4024
rect 9107 4016 9293 4024
rect 9327 4016 9533 4024
rect 10727 4016 10773 4024
rect 10847 4016 10953 4024
rect 11107 4016 11213 4024
rect 507 3996 913 4004
rect 967 3996 1004 4004
rect 467 3976 473 3984
rect 487 3976 973 3984
rect 996 3984 1004 3996
rect 1027 3996 1233 4004
rect 1267 3996 1313 4004
rect 1327 3996 1473 4004
rect 1667 3996 1713 4004
rect 2487 3996 2753 4004
rect 2787 3996 3033 4004
rect 3107 3996 3273 4004
rect 3647 3996 3733 4004
rect 4487 3996 4633 4004
rect 4867 3996 5173 4004
rect 5347 3996 5473 4004
rect 5707 3996 5913 4004
rect 6667 3996 6693 4004
rect 6947 3996 6953 4004
rect 6967 3996 7313 4004
rect 7327 3996 7533 4004
rect 7707 3996 7833 4004
rect 7907 3996 7953 4004
rect 8047 3996 8073 4004
rect 8107 3996 8144 4004
rect 996 3976 1413 3984
rect 1596 3976 1673 3984
rect 647 3956 673 3964
rect 727 3956 853 3964
rect 1227 3956 1353 3964
rect 1436 3947 1444 3973
rect 1596 3964 1604 3976
rect 1936 3984 1944 3993
rect 1936 3976 2273 3984
rect 2287 3976 2373 3984
rect 2527 3976 2813 3984
rect 3027 3976 3193 3984
rect 3207 3976 3233 3984
rect 3247 3976 3253 3984
rect 3507 3976 3653 3984
rect 3667 3976 4293 3984
rect 4447 3976 4693 3984
rect 5087 3976 5193 3984
rect 5207 3976 5393 3984
rect 5447 3976 5553 3984
rect 5627 3976 5993 3984
rect 6547 3976 6713 3984
rect 7167 3976 7373 3984
rect 7487 3976 7633 3984
rect 7867 3976 7913 3984
rect 8087 3976 8113 3984
rect 1507 3956 1604 3964
rect 1627 3956 1693 3964
rect 2547 3956 2633 3964
rect 2747 3956 2933 3964
rect 2967 3956 2973 3964
rect 2987 3956 3213 3964
rect 3547 3956 4213 3964
rect 4427 3956 4533 3964
rect 4667 3956 4933 3964
rect 5007 3956 5193 3964
rect 5207 3956 6233 3964
rect 6547 3956 7513 3964
rect 7587 3956 7653 3964
rect 7747 3956 7833 3964
rect 8136 3964 8144 3996
rect 8467 3996 8573 4004
rect 9027 3996 9073 4004
rect 9347 3996 9673 4004
rect 9687 3996 9713 4004
rect 9767 3996 9873 4004
rect 10207 3996 10273 4004
rect 10427 3996 10473 4004
rect 10647 3996 10713 4004
rect 11047 3996 11173 4004
rect 9296 3984 9304 3993
rect 8927 3976 9513 3984
rect 9927 3976 9953 3984
rect 10007 3976 10033 3984
rect 10087 3976 10233 3984
rect 10347 3976 10453 3984
rect 10607 3976 10733 3984
rect 10936 3984 10944 3993
rect 10936 3976 10953 3984
rect 11207 3976 11353 3984
rect 8107 3956 8144 3964
rect 8267 3956 8573 3964
rect 8807 3956 8973 3964
rect 8987 3956 9013 3964
rect 9207 3956 9253 3964
rect 9547 3956 9793 3964
rect 10407 3956 10433 3964
rect 10447 3956 10533 3964
rect 10727 3956 11253 3964
rect 2507 3936 2593 3944
rect 2607 3936 3173 3944
rect 3267 3936 3473 3944
rect 3487 3936 3793 3944
rect 5247 3936 5493 3944
rect 6927 3936 7453 3944
rect 7807 3936 8753 3944
rect 8767 3936 9153 3944
rect 10027 3936 10124 3944
rect 1427 3916 1653 3924
rect 2587 3916 3313 3924
rect 3607 3916 3693 3924
rect 5547 3916 5953 3924
rect 7387 3916 7773 3924
rect 8407 3916 9033 3924
rect 9047 3916 9273 3924
rect 9467 3916 10093 3924
rect 10116 3924 10124 3936
rect 10747 3936 10873 3944
rect 10116 3916 10473 3924
rect 10487 3916 10693 3924
rect 947 3896 973 3904
rect 987 3896 1153 3904
rect 2527 3896 4853 3904
rect 7847 3896 8853 3904
rect 8947 3896 10613 3904
rect 4507 3876 5253 3884
rect 5707 3876 7993 3884
rect 9567 3876 10533 3884
rect 3847 3856 4413 3864
rect 6527 3856 7113 3864
rect 7527 3856 8073 3864
rect 8527 3856 8853 3864
rect 9067 3856 9213 3864
rect 9447 3856 9553 3864
rect 10087 3856 10593 3864
rect 4087 3836 4313 3844
rect 4947 3836 6853 3844
rect 6867 3836 9453 3844
rect 9527 3836 10333 3844
rect 10447 3836 10573 3844
rect 2507 3816 3633 3824
rect 4047 3816 8873 3824
rect 10127 3816 10233 3824
rect 2207 3796 2433 3804
rect 2447 3796 5673 3804
rect 6387 3796 7453 3804
rect 7547 3796 8513 3804
rect 8627 3796 8933 3804
rect 9787 3796 10933 3804
rect 247 3776 393 3784
rect 407 3776 1173 3784
rect 2387 3776 2393 3784
rect 2407 3776 4273 3784
rect 4867 3776 5553 3784
rect 7087 3776 7913 3784
rect 8016 3776 9073 3784
rect 607 3756 733 3764
rect 1187 3756 1533 3764
rect 2167 3756 2693 3764
rect 2827 3756 3853 3764
rect 3867 3756 3893 3764
rect 4127 3756 4333 3764
rect 4567 3756 5053 3764
rect 5507 3756 5933 3764
rect 6667 3756 6893 3764
rect 6907 3756 7133 3764
rect 7207 3756 7753 3764
rect 8016 3764 8024 3776
rect 9247 3776 9713 3784
rect 9747 3776 10813 3784
rect 7767 3756 8024 3764
rect 8047 3756 8073 3764
rect 9367 3756 10073 3764
rect 10596 3756 10633 3764
rect 10596 3747 10604 3756
rect 11007 3756 11133 3764
rect 707 3736 793 3744
rect 1147 3736 1413 3744
rect 1707 3736 1753 3744
rect 1767 3736 2213 3744
rect 2876 3736 3093 3744
rect 2876 3727 2884 3736
rect 3187 3736 3293 3744
rect 3307 3736 4233 3744
rect 4327 3736 4893 3744
rect 5067 3736 5373 3744
rect 5607 3736 5893 3744
rect 5987 3736 6153 3744
rect 6627 3736 6673 3744
rect 6687 3736 7073 3744
rect 7127 3736 7233 3744
rect 7867 3736 8053 3744
rect 8127 3736 8733 3744
rect 8747 3736 9733 3744
rect 10427 3736 10513 3744
rect 10647 3736 10673 3744
rect 11147 3736 11293 3744
rect 207 3716 253 3724
rect 547 3716 913 3724
rect 927 3716 1113 3724
rect 1227 3716 1433 3724
rect 1547 3716 1913 3724
rect 2667 3716 2733 3724
rect 3127 3716 3193 3724
rect 3227 3716 3373 3724
rect 3387 3716 3593 3724
rect 3616 3716 4373 3724
rect 427 3696 493 3704
rect 687 3696 713 3704
rect 947 3696 1253 3704
rect 2187 3696 2513 3704
rect 2547 3696 2673 3704
rect 3616 3704 3624 3716
rect 4507 3716 4613 3724
rect 4707 3716 5013 3724
rect 5147 3716 5353 3724
rect 5427 3716 5673 3724
rect 5947 3716 6433 3724
rect 6647 3716 7133 3724
rect 7336 3716 7533 3724
rect 7336 3707 7344 3716
rect 8047 3716 8093 3724
rect 8347 3716 8533 3724
rect 8547 3716 8653 3724
rect 8727 3716 9433 3724
rect 9927 3716 9973 3724
rect 10307 3716 10413 3724
rect 10627 3716 10833 3724
rect 2707 3696 3624 3704
rect 3667 3696 3873 3704
rect 4147 3696 4173 3704
rect 4467 3696 4593 3704
rect 5187 3696 5513 3704
rect 6167 3696 6553 3704
rect 6607 3696 6653 3704
rect 6887 3696 6953 3704
rect 7107 3696 7293 3704
rect 7747 3696 7993 3704
rect 8027 3696 8253 3704
rect 8307 3696 8373 3704
rect 8387 3696 8513 3704
rect 8567 3696 8913 3704
rect 9387 3696 9413 3704
rect 9476 3704 9484 3713
rect 9476 3696 9693 3704
rect 9707 3696 9833 3704
rect 10547 3696 10853 3704
rect 10987 3696 11293 3704
rect 267 3676 433 3684
rect 467 3676 1013 3684
rect 1127 3676 1673 3684
rect 1907 3676 2133 3684
rect 3147 3676 3353 3684
rect 4167 3676 4373 3684
rect 4427 3676 4833 3684
rect 4887 3676 5393 3684
rect 5447 3676 5613 3684
rect 5647 3676 6133 3684
rect 6707 3676 6853 3684
rect 7327 3676 7513 3684
rect 7567 3676 7733 3684
rect 7787 3676 7813 3684
rect 7827 3676 8113 3684
rect 8287 3676 8533 3684
rect 8667 3676 8973 3684
rect 9407 3676 9473 3684
rect 9667 3676 9713 3684
rect 10167 3676 10313 3684
rect 10887 3676 10953 3684
rect 10967 3676 11053 3684
rect 11167 3676 11333 3684
rect 227 3656 453 3664
rect 667 3656 713 3664
rect 967 3656 1013 3664
rect 1027 3656 1633 3664
rect 4107 3656 4153 3664
rect 4587 3656 4633 3664
rect 5027 3656 5113 3664
rect 6247 3656 6913 3664
rect 7247 3656 7753 3664
rect 8067 3656 8633 3664
rect 9027 3656 9173 3664
rect 9187 3656 9973 3664
rect 10147 3656 10173 3664
rect 10827 3656 11073 3664
rect 1627 3636 5033 3644
rect 5187 3636 5573 3644
rect 5607 3636 5813 3644
rect 6767 3636 7253 3644
rect 8267 3636 8453 3644
rect 8567 3636 8793 3644
rect 8807 3636 8833 3644
rect 8847 3636 9293 3644
rect 9467 3636 9613 3644
rect 5567 3616 5813 3624
rect 5927 3616 5953 3624
rect 6867 3616 7713 3624
rect 8107 3616 8453 3624
rect 8507 3616 10373 3624
rect 1347 3596 1413 3604
rect 1427 3596 2133 3604
rect 3067 3596 3433 3604
rect 3467 3596 3793 3604
rect 5167 3596 5633 3604
rect 5647 3596 6273 3604
rect 6787 3596 6833 3604
rect 7227 3596 7313 3604
rect 7687 3596 7713 3604
rect 7747 3596 9513 3604
rect 9607 3596 9693 3604
rect 9747 3596 10673 3604
rect 1207 3576 1233 3584
rect 1447 3576 1893 3584
rect 2767 3576 2893 3584
rect 3207 3576 3813 3584
rect 3827 3576 4593 3584
rect 5787 3576 6113 3584
rect 6287 3576 6433 3584
rect 6447 3576 7113 3584
rect 7147 3576 7173 3584
rect 7187 3576 7513 3584
rect 8447 3576 8893 3584
rect 8907 3576 8953 3584
rect 9607 3576 9753 3584
rect 1967 3556 2433 3564
rect 2527 3556 2893 3564
rect 2927 3556 3373 3564
rect 3687 3556 4513 3564
rect 5627 3556 5793 3564
rect 6107 3556 6153 3564
rect 6167 3556 7193 3564
rect 7267 3556 7293 3564
rect 7307 3556 7733 3564
rect 7927 3556 8213 3564
rect 8947 3556 9093 3564
rect 9347 3556 9953 3564
rect 10387 3556 10633 3564
rect 10647 3556 11313 3564
rect 2427 3536 2444 3544
rect 787 3516 933 3524
rect 2436 3524 2444 3536
rect 2467 3536 2533 3544
rect 2887 3536 3193 3544
rect 3407 3536 3613 3544
rect 3867 3536 3913 3544
rect 3927 3536 4093 3544
rect 4127 3536 4564 3544
rect 2436 3516 2453 3524
rect 2727 3516 2813 3524
rect 2827 3516 3133 3524
rect 3207 3516 3233 3524
rect 4147 3516 4213 3524
rect 427 3496 453 3504
rect 747 3496 793 3504
rect 807 3496 953 3504
rect 1067 3496 1773 3504
rect 2687 3496 3093 3504
rect 2207 3476 2353 3484
rect 2607 3476 2653 3484
rect 2707 3476 2733 3484
rect 3156 3484 3164 3513
rect 3187 3496 3373 3504
rect 3887 3496 4413 3504
rect 3156 3476 3173 3484
rect 4107 3476 4153 3484
rect 387 3456 893 3464
rect 1727 3456 1733 3464
rect 1747 3456 3633 3464
rect 3987 3456 4193 3464
rect 4536 3464 4544 3493
rect 4556 3487 4564 3536
rect 5227 3536 5273 3544
rect 5327 3536 5353 3544
rect 5587 3536 5793 3544
rect 5807 3536 6573 3544
rect 6807 3536 7033 3544
rect 7047 3536 7733 3544
rect 7747 3536 8413 3544
rect 8707 3536 8753 3544
rect 8767 3536 9493 3544
rect 10207 3536 10333 3544
rect 10347 3536 10693 3544
rect 10707 3536 10833 3544
rect 10867 3536 10973 3544
rect 4827 3516 4973 3524
rect 5107 3516 5493 3524
rect 6507 3516 6533 3524
rect 7027 3516 7093 3524
rect 7127 3516 7213 3524
rect 7227 3516 7373 3524
rect 7787 3516 7833 3524
rect 7947 3516 7973 3524
rect 8467 3516 8793 3524
rect 8867 3516 8893 3524
rect 9007 3516 9113 3524
rect 9127 3516 9193 3524
rect 9527 3516 9573 3524
rect 9596 3516 9613 3524
rect 4767 3496 5033 3504
rect 5187 3496 5233 3504
rect 5527 3496 5593 3504
rect 5927 3496 6033 3504
rect 6327 3496 6793 3504
rect 6976 3504 6984 3513
rect 6976 3496 7073 3504
rect 7767 3496 7973 3504
rect 8227 3496 8353 3504
rect 8367 3496 9053 3504
rect 9356 3504 9364 3513
rect 9356 3496 9373 3504
rect 9396 3504 9404 3513
rect 9596 3504 9604 3516
rect 9627 3516 9853 3524
rect 9887 3516 9993 3524
rect 10087 3516 10573 3524
rect 10687 3516 10753 3524
rect 10827 3516 10913 3524
rect 10927 3516 11053 3524
rect 11107 3516 11153 3524
rect 11167 3516 11293 3524
rect 9396 3496 9604 3504
rect 9767 3496 9873 3504
rect 9887 3496 10333 3504
rect 10347 3496 10433 3504
rect 10627 3496 10693 3504
rect 5147 3476 5273 3484
rect 5887 3476 6073 3484
rect 6307 3476 6353 3484
rect 6387 3476 7233 3484
rect 7247 3476 7304 3484
rect 4536 3456 4773 3464
rect 4787 3456 4813 3464
rect 5007 3456 5313 3464
rect 6147 3456 6333 3464
rect 7107 3456 7273 3464
rect 7296 3464 7304 3476
rect 7467 3476 7533 3484
rect 7547 3476 7933 3484
rect 8007 3476 8233 3484
rect 8247 3476 8473 3484
rect 8487 3476 10193 3484
rect 7296 3456 8993 3464
rect 9387 3456 9413 3464
rect 9687 3456 10073 3464
rect 10127 3456 10353 3464
rect 987 3436 2333 3444
rect 4347 3436 4433 3444
rect 4447 3436 4513 3444
rect 4527 3436 5553 3444
rect 8987 3436 9833 3444
rect 9847 3436 9853 3444
rect 9867 3436 9933 3444
rect 2447 3416 5713 3424
rect 6487 3416 6573 3424
rect 4607 3396 7553 3404
rect 7707 3396 7773 3404
rect 8207 3396 8553 3404
rect 327 3376 353 3384
rect 3247 3376 5073 3384
rect 7707 3376 8193 3384
rect 5667 3356 6013 3364
rect 7427 3356 7693 3364
rect 7716 3356 8433 3364
rect 7716 3344 7724 3356
rect 7567 3336 7724 3344
rect 9447 3336 9653 3344
rect 9667 3336 10253 3344
rect 787 3316 1673 3324
rect 2267 3316 2633 3324
rect 4747 3316 10273 3324
rect 187 3296 1653 3304
rect 1667 3296 3793 3304
rect 6047 3296 6853 3304
rect 7107 3296 7973 3304
rect 7987 3296 8093 3304
rect 9887 3296 9893 3304
rect 9907 3296 11173 3304
rect 1687 3276 2373 3284
rect 3007 3276 3073 3284
rect 5307 3276 5453 3284
rect 5467 3276 5733 3284
rect 5767 3276 5813 3284
rect 6727 3276 6913 3284
rect 7967 3276 8593 3284
rect 9607 3276 9633 3284
rect 10167 3276 10193 3284
rect -24 3256 173 3264
rect 747 3256 1113 3264
rect 2147 3256 2313 3264
rect 2387 3256 2593 3264
rect 2647 3256 2653 3264
rect 2667 3256 2833 3264
rect 4127 3256 4673 3264
rect 5547 3256 5773 3264
rect 6227 3256 6293 3264
rect 6567 3256 6733 3264
rect 7447 3256 7473 3264
rect 7667 3256 7753 3264
rect 7827 3256 8613 3264
rect 8707 3256 9073 3264
rect 9627 3256 9913 3264
rect 9927 3256 10053 3264
rect 10067 3256 10573 3264
rect 227 3236 413 3244
rect 427 3236 533 3244
rect 587 3236 653 3244
rect 667 3236 773 3244
rect 1087 3236 1313 3244
rect 1367 3236 1513 3244
rect 1707 3236 2673 3244
rect 3387 3236 3573 3244
rect 3587 3236 3613 3244
rect 3727 3236 3933 3244
rect 4647 3236 4713 3244
rect 4807 3236 4853 3244
rect 5287 3236 5713 3244
rect 6207 3236 6233 3244
rect 6367 3236 6453 3244
rect 6487 3236 6533 3244
rect 6547 3236 6724 3244
rect 6716 3227 6724 3236
rect 6907 3236 6933 3244
rect 6987 3236 7013 3244
rect 7027 3236 7353 3244
rect 7387 3236 7673 3244
rect 8107 3236 8133 3244
rect 8847 3236 8893 3244
rect 9807 3236 10113 3244
rect 10167 3236 10293 3244
rect 407 3216 513 3224
rect 567 3216 633 3224
rect 707 3216 953 3224
rect 967 3216 1053 3224
rect 1487 3216 1753 3224
rect 2467 3216 2733 3224
rect 3047 3216 3593 3224
rect 3647 3216 4613 3224
rect 4667 3216 4673 3224
rect 4687 3216 6253 3224
rect 6267 3216 6493 3224
rect 7247 3216 7313 3224
rect 7327 3216 7813 3224
rect 7927 3216 7953 3224
rect 8167 3216 8393 3224
rect 8927 3216 9013 3224
rect 9547 3216 9613 3224
rect 10147 3216 10213 3224
rect 10367 3216 10553 3224
rect 10767 3216 10813 3224
rect 10867 3216 10913 3224
rect 11107 3216 11153 3224
rect 11247 3216 11273 3224
rect 727 3196 793 3204
rect 1107 3196 1133 3204
rect 1367 3196 2033 3204
rect 2047 3196 2053 3204
rect 2067 3196 2404 3204
rect 487 3176 993 3184
rect 1887 3176 2113 3184
rect 2396 3184 2404 3196
rect 2427 3196 2653 3204
rect 2867 3196 3353 3204
rect 4267 3196 5793 3204
rect 6747 3196 6953 3204
rect 7887 3196 8173 3204
rect 8187 3196 8453 3204
rect 8467 3196 8633 3204
rect 8647 3196 8773 3204
rect 8807 3196 8933 3204
rect 9007 3196 9133 3204
rect 9147 3196 9633 3204
rect 9967 3196 9993 3204
rect 10007 3196 10393 3204
rect 10947 3196 11073 3204
rect 11187 3196 11293 3204
rect 2396 3176 3013 3184
rect 3027 3176 3033 3184
rect 3147 3176 3553 3184
rect 3627 3176 5233 3184
rect 5247 3176 5493 3184
rect 6067 3176 6213 3184
rect 6227 3176 7193 3184
rect 7587 3176 8373 3184
rect 9167 3176 9373 3184
rect 9387 3176 9513 3184
rect 10187 3176 10393 3184
rect 11067 3176 11333 3184
rect 967 3156 1333 3164
rect 1347 3156 4153 3164
rect 4187 3156 4713 3164
rect 4727 3156 6013 3164
rect 6127 3156 7533 3164
rect 8127 3156 8293 3164
rect 9207 3156 10213 3164
rect 10227 3156 10733 3164
rect 11207 3156 11333 3164
rect 3307 3136 3393 3144
rect 6007 3136 6133 3144
rect 6147 3136 8493 3144
rect 9507 3136 10033 3144
rect 10047 3136 10593 3144
rect 2647 3116 3053 3124
rect 3147 3116 4293 3124
rect 4387 3116 5033 3124
rect 6807 3116 7293 3124
rect 2227 3096 2613 3104
rect 3067 3096 3333 3104
rect 6087 3096 6153 3104
rect 6947 3096 7053 3104
rect 7587 3096 7913 3104
rect 9107 3096 9633 3104
rect 3367 3076 4033 3084
rect 4347 3076 4973 3084
rect 6827 3076 6993 3084
rect 7007 3076 7053 3084
rect 7067 3076 7373 3084
rect 7387 3076 7993 3084
rect 8007 3076 8493 3084
rect 8987 3076 9093 3084
rect 10267 3076 10433 3084
rect 10447 3076 10833 3084
rect 447 3056 613 3064
rect 1167 3056 1373 3064
rect 1887 3056 2553 3064
rect 2867 3056 3273 3064
rect 3327 3056 3533 3064
rect 3827 3056 3993 3064
rect 4407 3056 4533 3064
rect 4547 3056 4733 3064
rect 6387 3056 6413 3064
rect 6467 3056 6833 3064
rect 6887 3056 7073 3064
rect 7667 3056 7713 3064
rect 7727 3056 8013 3064
rect 8287 3056 8313 3064
rect 8447 3056 8533 3064
rect 8827 3056 8873 3064
rect 8887 3056 9213 3064
rect 9907 3056 9933 3064
rect 10127 3056 10173 3064
rect 10327 3056 10333 3064
rect 10347 3056 10373 3064
rect 10647 3056 10813 3064
rect 647 3036 713 3044
rect 1467 3036 1633 3044
rect 1687 3036 1733 3044
rect 2087 3036 2193 3044
rect 3996 3036 4253 3044
rect 3996 3027 4004 3036
rect 4647 3036 4713 3044
rect 4727 3036 5173 3044
rect 5327 3036 5453 3044
rect 6227 3036 6393 3044
rect 6627 3036 6653 3044
rect 7107 3036 7133 3044
rect 7347 3036 7553 3044
rect 7627 3036 7873 3044
rect 7967 3036 8033 3044
rect 8067 3036 8253 3044
rect 8307 3036 8673 3044
rect 8687 3036 8713 3044
rect 8767 3036 8813 3044
rect 8907 3036 9013 3044
rect 9027 3036 9193 3044
rect 9687 3036 9833 3044
rect 9847 3036 9873 3044
rect 9927 3036 10033 3044
rect 10067 3036 10133 3044
rect 10247 3036 10573 3044
rect 10767 3036 10793 3044
rect 10847 3036 10873 3044
rect 10887 3036 11033 3044
rect 287 3016 393 3024
rect 427 3016 653 3024
rect 1427 3016 1613 3024
rect 2187 3016 2333 3024
rect 2347 3016 2433 3024
rect 2847 3016 3233 3024
rect 3267 3016 3353 3024
rect 4247 3016 4773 3024
rect 5127 3016 5233 3024
rect 5387 3016 5433 3024
rect 5487 3016 5693 3024
rect 6647 3016 7204 3024
rect 247 2996 413 3004
rect 927 2996 953 3004
rect 967 2996 1653 3004
rect 1907 2996 2253 3004
rect 2287 2996 2533 3004
rect 2547 2996 3033 3004
rect 3087 2996 3093 3004
rect 3107 2996 3393 3004
rect 5407 2996 5673 3004
rect 5727 2996 5853 3004
rect 5947 2996 6033 3004
rect 6047 2996 6173 3004
rect 6607 2996 7173 3004
rect 7196 3004 7204 3016
rect 7547 3016 7593 3024
rect 7767 3016 7813 3024
rect 8747 3016 9253 3024
rect 9267 3016 9453 3024
rect 9876 3016 9933 3024
rect 9876 3007 9884 3016
rect 10207 3016 10353 3024
rect 10907 3016 11053 3024
rect 7196 2996 7793 3004
rect 10387 2996 10433 3004
rect 10607 2996 10633 3004
rect 10867 2996 11293 3004
rect 707 2976 753 2984
rect 2307 2976 2533 2984
rect 2547 2976 2613 2984
rect 3307 2976 3413 2984
rect 7807 2976 7833 2984
rect 9307 2976 9893 2984
rect 9907 2976 10333 2984
rect 10347 2976 10553 2984
rect 10587 2976 10713 2984
rect 10987 2976 11053 2984
rect 467 2956 793 2964
rect 1527 2956 2573 2964
rect 7027 2956 7353 2964
rect 7367 2956 8493 2964
rect 10367 2956 10533 2964
rect 10807 2956 11073 2964
rect 11087 2956 11253 2964
rect 767 2936 993 2944
rect 1007 2936 1693 2944
rect 1707 2936 1713 2944
rect 5967 2936 10233 2944
rect 10487 2936 10533 2944
rect 4527 2916 5333 2924
rect 1587 2896 1853 2904
rect 5067 2896 5133 2904
rect 1607 2876 10413 2884
rect 4887 2856 5173 2864
rect 5247 2856 5353 2864
rect 7647 2856 8253 2864
rect 8267 2856 10113 2864
rect 3327 2836 8193 2844
rect 10047 2816 11073 2824
rect 1147 2796 2993 2804
rect 3007 2796 3053 2804
rect 4027 2796 4213 2804
rect 5127 2796 5193 2804
rect 6627 2796 6653 2804
rect 6667 2796 6773 2804
rect 6987 2796 8653 2804
rect 9987 2796 10113 2804
rect 10167 2796 10653 2804
rect 10927 2796 10944 2804
rect 247 2776 413 2784
rect 427 2776 653 2784
rect 667 2776 873 2784
rect 1087 2776 1353 2784
rect 1667 2776 2313 2784
rect 2596 2776 2793 2784
rect 207 2756 433 2764
rect 447 2756 613 2764
rect 627 2756 673 2764
rect 807 2736 893 2744
rect 967 2736 1124 2744
rect 1116 2727 1124 2736
rect 1287 2736 1333 2744
rect 227 2716 593 2724
rect 927 2716 973 2724
rect 1356 2724 1364 2753
rect 1376 2747 1384 2773
rect 1407 2756 1453 2764
rect 2147 2756 2573 2764
rect 2596 2764 2604 2776
rect 3387 2776 3593 2784
rect 4947 2776 5253 2784
rect 5767 2776 6653 2784
rect 6667 2776 6993 2784
rect 8087 2776 8113 2784
rect 8447 2776 9693 2784
rect 10507 2776 10653 2784
rect 10667 2776 10693 2784
rect 10747 2776 10813 2784
rect 10847 2776 10913 2784
rect 10936 2767 10944 2796
rect 10967 2796 11213 2804
rect 10967 2776 10993 2784
rect 11007 2776 11033 2784
rect 11147 2776 11193 2784
rect 2587 2756 2604 2764
rect 2627 2756 3104 2764
rect 1687 2736 1733 2744
rect 1747 2736 2633 2744
rect 2807 2736 3033 2744
rect 3047 2736 3073 2744
rect 3096 2744 3104 2756
rect 3447 2756 3633 2764
rect 3747 2756 3933 2764
rect 4107 2756 4233 2764
rect 5127 2756 5153 2764
rect 5207 2756 5273 2764
rect 5687 2756 5713 2764
rect 6387 2756 6753 2764
rect 6847 2756 7084 2764
rect 7076 2747 7084 2756
rect 7127 2756 7273 2764
rect 7507 2756 7553 2764
rect 7607 2756 7733 2764
rect 8567 2756 8593 2764
rect 8667 2756 8753 2764
rect 9587 2756 9673 2764
rect 10287 2756 10333 2764
rect 10487 2756 10553 2764
rect 10687 2756 10713 2764
rect 3096 2736 3493 2744
rect 3507 2736 4273 2744
rect 4287 2736 4453 2744
rect 4467 2736 4573 2744
rect 4707 2736 4813 2744
rect 5147 2736 5293 2744
rect 6067 2736 6093 2744
rect 6347 2736 6593 2744
rect 7007 2736 7033 2744
rect 7187 2736 7293 2744
rect 7747 2736 7873 2744
rect 7887 2736 8013 2744
rect 8307 2736 8533 2744
rect 8647 2736 8733 2744
rect 8747 2736 9253 2744
rect 9307 2736 9533 2744
rect 9787 2736 9833 2744
rect 9847 2736 10053 2744
rect 10067 2736 10293 2744
rect 10507 2736 10533 2744
rect 11087 2736 11133 2744
rect 1347 2716 1513 2724
rect 1787 2716 2593 2724
rect 2616 2716 3213 2724
rect 2616 2704 2624 2716
rect 3347 2716 3533 2724
rect 4667 2716 4953 2724
rect 5327 2716 5413 2724
rect 6427 2716 6633 2724
rect 6647 2716 6813 2724
rect 7167 2716 7353 2724
rect 8027 2716 8573 2724
rect 8987 2716 9353 2724
rect 9367 2716 9793 2724
rect 9827 2716 9853 2724
rect 10047 2716 10093 2724
rect 10227 2716 10273 2724
rect 10327 2716 10433 2724
rect 10447 2716 10593 2724
rect 11027 2716 11173 2724
rect 2327 2696 2624 2704
rect 2647 2696 3313 2704
rect 5787 2696 5893 2704
rect 8167 2696 8273 2704
rect 9487 2696 9533 2704
rect 9927 2696 10013 2704
rect 10027 2696 10353 2704
rect 1827 2676 1873 2684
rect 2387 2676 3953 2684
rect 3967 2676 4413 2684
rect 5367 2676 5393 2684
rect 7067 2676 9513 2684
rect 1887 2656 2093 2664
rect 2567 2656 2713 2664
rect 5567 2656 8453 2664
rect 8527 2656 8853 2664
rect 8867 2656 9053 2664
rect 1607 2636 1733 2644
rect 1747 2636 2273 2644
rect 2667 2636 2833 2644
rect 3327 2636 4293 2644
rect 4827 2636 5193 2644
rect 5647 2636 5873 2644
rect 5887 2636 6333 2644
rect 6347 2636 7693 2644
rect 7847 2636 7953 2644
rect 7967 2636 10253 2644
rect 1207 2616 1633 2624
rect 2107 2616 2153 2624
rect 2767 2616 2813 2624
rect 3347 2616 3513 2624
rect 3527 2616 3713 2624
rect 4427 2616 5553 2624
rect 7227 2616 8073 2624
rect 8087 2616 8273 2624
rect 8287 2616 8473 2624
rect 8827 2616 9173 2624
rect 9187 2616 9233 2624
rect 607 2596 613 2604
rect 627 2596 1073 2604
rect 1567 2596 1633 2604
rect 1647 2596 2413 2604
rect 2427 2596 2513 2604
rect 2607 2596 2833 2604
rect 3567 2596 4053 2604
rect 4567 2596 5913 2604
rect 7967 2596 8233 2604
rect 8247 2596 8253 2604
rect 8267 2596 8513 2604
rect 8667 2596 8673 2604
rect 8687 2596 8893 2604
rect 8956 2596 9853 2604
rect 227 2576 393 2584
rect 427 2576 693 2584
rect 1307 2576 1373 2584
rect 1407 2576 1573 2584
rect 1867 2576 2033 2584
rect 2047 2576 2113 2584
rect 2127 2576 2653 2584
rect 3467 2576 4073 2584
rect 4267 2576 4633 2584
rect 4647 2576 4813 2584
rect 4847 2576 5053 2584
rect 5127 2576 5313 2584
rect 5627 2576 5753 2584
rect 5847 2576 6393 2584
rect 6507 2576 6753 2584
rect 7987 2576 8004 2584
rect 667 2556 733 2564
rect 2067 2556 2193 2564
rect 2207 2556 2553 2564
rect 3287 2556 3973 2564
rect 4607 2556 4733 2564
rect 4787 2556 4853 2564
rect 5607 2556 5713 2564
rect 5807 2556 6013 2564
rect 6187 2556 6293 2564
rect 6367 2556 6513 2564
rect 6747 2556 6893 2564
rect 7027 2556 7053 2564
rect 7187 2556 7253 2564
rect 207 2536 273 2544
rect 307 2536 573 2544
rect 587 2536 773 2544
rect 1167 2536 1433 2544
rect 2047 2536 2073 2544
rect 2207 2536 2273 2544
rect 2447 2536 2573 2544
rect 2627 2536 2653 2544
rect 3027 2536 3233 2544
rect 3247 2536 3733 2544
rect 3887 2536 4033 2544
rect 4087 2536 4353 2544
rect 4367 2536 4393 2544
rect 4467 2536 4573 2544
rect 4627 2536 4773 2544
rect 4807 2536 5073 2544
rect 5187 2536 5333 2544
rect 6267 2536 6293 2544
rect 6727 2536 6793 2544
rect 6927 2536 6993 2544
rect 7007 2536 7073 2544
rect 7147 2536 7233 2544
rect 7907 2536 7953 2544
rect 47 2516 173 2524
rect 187 2516 253 2524
rect 267 2516 733 2524
rect 747 2516 753 2524
rect 1787 2516 2293 2524
rect 2347 2516 2493 2524
rect 3827 2516 4253 2524
rect 5927 2516 5953 2524
rect 5967 2516 6213 2524
rect 6227 2516 6233 2524
rect 6287 2516 6353 2524
rect 6407 2516 6513 2524
rect 6527 2516 6673 2524
rect 6707 2516 6953 2524
rect 6967 2516 7113 2524
rect 7527 2516 7633 2524
rect 7647 2516 7653 2524
rect 7976 2524 7984 2553
rect 7996 2547 8004 2576
rect 8956 2584 8964 2596
rect 10587 2596 10833 2604
rect 10847 2596 10933 2604
rect 8467 2576 8964 2584
rect 9367 2576 9413 2584
rect 10547 2576 10613 2584
rect 10967 2576 11353 2584
rect 8487 2556 8993 2564
rect 9207 2556 9213 2564
rect 9227 2556 9653 2564
rect 9827 2556 9873 2564
rect 10307 2556 10333 2564
rect 10707 2556 10793 2564
rect 7976 2516 8173 2524
rect 8216 2524 8224 2553
rect 8247 2536 8313 2544
rect 8947 2536 9393 2544
rect 9447 2536 9493 2544
rect 10647 2536 10853 2544
rect 11067 2536 11093 2544
rect 11307 2536 11353 2544
rect 8216 2516 8233 2524
rect 8967 2516 9473 2524
rect 9936 2524 9944 2533
rect 9936 2516 10093 2524
rect 10147 2516 10313 2524
rect 10347 2516 10653 2524
rect 10847 2516 10873 2524
rect 11087 2516 11273 2524
rect 687 2496 1613 2504
rect 2167 2496 4313 2504
rect 5847 2496 6153 2504
rect 6167 2496 6473 2504
rect 7487 2496 7613 2504
rect 9916 2504 9924 2513
rect 9916 2496 10013 2504
rect 10087 2496 10113 2504
rect 10267 2496 10333 2504
rect 11047 2496 11073 2504
rect 11267 2496 11313 2504
rect 687 2476 713 2484
rect 1727 2476 2353 2484
rect 2367 2476 3293 2484
rect 5307 2476 5693 2484
rect 6147 2476 8213 2484
rect 8747 2476 8833 2484
rect 8847 2476 9173 2484
rect 9187 2476 9453 2484
rect 9467 2476 9973 2484
rect 3307 2456 4433 2464
rect 4447 2456 5213 2464
rect 567 2436 793 2444
rect 1767 2416 1833 2424
rect 4847 2396 4913 2404
rect 5987 2396 6273 2404
rect 4607 2376 5013 2384
rect 5987 2376 6593 2384
rect 287 2356 353 2364
rect 3987 2356 4473 2364
rect 6207 2356 7393 2364
rect 7727 2356 8753 2364
rect 9827 2356 9853 2364
rect 10227 2356 11153 2364
rect 2667 2336 2673 2344
rect 2687 2336 3393 2344
rect 3407 2336 3773 2344
rect 3787 2336 3793 2344
rect 3807 2336 4073 2344
rect 6507 2336 6873 2344
rect 7147 2336 8093 2344
rect 8107 2336 8993 2344
rect 9007 2336 9333 2344
rect 9747 2336 9813 2344
rect 10087 2336 10233 2344
rect 10367 2336 10473 2344
rect 11067 2336 11193 2344
rect 3907 2316 4713 2324
rect 6607 2316 7413 2324
rect 8536 2316 8773 2324
rect 8536 2307 8544 2316
rect 8927 2316 9033 2324
rect 9667 2316 9793 2324
rect 10027 2316 10373 2324
rect 11027 2316 11193 2324
rect 11207 2316 11313 2324
rect 607 2296 673 2304
rect 1376 2296 1393 2304
rect 1376 2287 1384 2296
rect 2187 2296 2333 2304
rect 2347 2296 2533 2304
rect 2547 2296 2593 2304
rect 2647 2296 3293 2304
rect 3327 2296 3353 2304
rect 3367 2296 3913 2304
rect 4087 2296 5193 2304
rect 5207 2296 5253 2304
rect 5727 2296 5913 2304
rect 5927 2296 5993 2304
rect 6127 2296 6553 2304
rect 6567 2296 6833 2304
rect 7727 2296 7853 2304
rect 8587 2296 8613 2304
rect 9087 2296 9173 2304
rect 9767 2296 9913 2304
rect 9987 2296 10093 2304
rect 10327 2296 10433 2304
rect 10727 2296 10853 2304
rect 10867 2296 10873 2304
rect 11087 2296 11153 2304
rect 467 2276 653 2284
rect 667 2276 793 2284
rect 1427 2276 1473 2284
rect 1747 2276 1793 2284
rect 1847 2276 1893 2284
rect 2327 2276 2553 2284
rect 3247 2276 3433 2284
rect 3747 2276 3813 2284
rect 3947 2276 3973 2284
rect 3996 2284 4004 2293
rect 3996 2276 4013 2284
rect 4047 2276 4113 2284
rect 4507 2276 4673 2284
rect 5687 2276 5813 2284
rect 5827 2276 5873 2284
rect 6107 2276 6213 2284
rect 6247 2276 6553 2284
rect 6567 2276 6693 2284
rect 6856 2276 7093 2284
rect 387 2256 613 2264
rect 707 2256 1133 2264
rect 1156 2264 1164 2273
rect 1156 2256 1393 2264
rect 1447 2256 1773 2264
rect 2347 2256 2393 2264
rect 2467 2256 2533 2264
rect 3767 2256 3993 2264
rect 6067 2256 6153 2264
rect 6307 2256 6633 2264
rect 6687 2256 6813 2264
rect 6856 2264 6864 2276
rect 7107 2276 7293 2284
rect 7307 2276 7353 2284
rect 7367 2276 7473 2284
rect 7487 2276 7664 2284
rect 7656 2267 7664 2276
rect 7816 2276 8253 2284
rect 7816 2267 7824 2276
rect 8787 2276 9013 2284
rect 9067 2276 9653 2284
rect 9747 2276 9853 2284
rect 10467 2276 10633 2284
rect 10767 2276 10933 2284
rect 11147 2276 11173 2284
rect 6827 2256 6864 2264
rect 6887 2256 7113 2264
rect 7167 2256 7193 2264
rect 7387 2256 7593 2264
rect 7676 2256 7813 2264
rect 107 2236 193 2244
rect 1127 2236 1193 2244
rect 2107 2236 2273 2244
rect 2287 2236 2373 2244
rect 2587 2236 2813 2244
rect 3107 2236 3273 2244
rect 3947 2236 3993 2244
rect 4447 2236 5413 2244
rect 6047 2236 6133 2244
rect 6407 2236 6433 2244
rect 7676 2244 7684 2256
rect 8067 2256 8353 2264
rect 8567 2256 8793 2264
rect 9307 2256 9353 2264
rect 9487 2256 9833 2264
rect 10187 2256 10273 2264
rect 10287 2256 10313 2264
rect 10327 2256 11013 2264
rect 7427 2236 7684 2244
rect 7807 2236 7833 2244
rect 7847 2236 8913 2244
rect 9287 2236 9313 2244
rect 9447 2236 9613 2244
rect 10107 2236 10253 2244
rect 10467 2236 10553 2244
rect 10687 2236 10693 2244
rect 10707 2236 10913 2244
rect 87 2216 713 2224
rect 887 2216 1193 2224
rect 3107 2216 3613 2224
rect 3867 2216 4233 2224
rect 4807 2216 5033 2224
rect 7867 2216 9513 2224
rect 9527 2216 9553 2224
rect 9567 2216 9993 2224
rect 10247 2216 10353 2224
rect 10367 2216 10933 2224
rect 10947 2216 11253 2224
rect 1187 2196 1413 2204
rect 3627 2196 3873 2204
rect 7687 2196 7893 2204
rect 7907 2196 8093 2204
rect 10387 2196 10733 2204
rect 4287 2176 4413 2184
rect 4427 2176 4853 2184
rect 4867 2176 4933 2184
rect 4947 2176 5213 2184
rect 5227 2176 5593 2184
rect 6827 2176 7933 2184
rect 8227 2176 8593 2184
rect 8607 2176 10553 2184
rect 747 2156 913 2164
rect 5167 2156 5193 2164
rect 7627 2156 7753 2164
rect 7767 2156 8513 2164
rect 9627 2156 9713 2164
rect 9767 2156 10393 2164
rect 10407 2156 10793 2164
rect 2147 2136 3393 2144
rect 5207 2136 5293 2144
rect 6767 2136 6993 2144
rect 7007 2136 7313 2144
rect 7947 2136 8393 2144
rect 8507 2136 8693 2144
rect 8707 2136 9753 2144
rect 10987 2136 11153 2144
rect 1707 2116 2153 2124
rect 2527 2116 2553 2124
rect 2567 2116 2673 2124
rect 3027 2116 3133 2124
rect 3307 2116 3813 2124
rect 6187 2116 6253 2124
rect 6947 2116 7013 2124
rect 7187 2116 7213 2124
rect 7267 2116 8033 2124
rect 8167 2116 8253 2124
rect 8687 2116 8893 2124
rect 8907 2116 8953 2124
rect 9107 2116 9393 2124
rect 9987 2116 10513 2124
rect 10987 2116 11273 2124
rect 11287 2116 11293 2124
rect 947 2096 1073 2104
rect 1467 2096 2573 2104
rect 2587 2096 2773 2104
rect 2907 2096 3313 2104
rect 3447 2096 4273 2104
rect 4387 2096 4553 2104
rect 5327 2096 5473 2104
rect 6207 2096 6224 2104
rect 87 2076 493 2084
rect 607 2076 664 2084
rect 427 2056 453 2064
rect 527 2056 633 2064
rect 656 2044 664 2076
rect 776 2067 784 2093
rect 907 2076 973 2084
rect 987 2076 1224 2084
rect 1216 2067 1224 2076
rect 1247 2076 1533 2084
rect 1827 2076 2113 2084
rect 2307 2076 2353 2084
rect 2767 2076 2813 2084
rect 2867 2076 3073 2084
rect 3347 2076 3844 2084
rect 1127 2056 1173 2064
rect 1667 2056 1753 2064
rect 1767 2056 1873 2064
rect 2396 2064 2404 2073
rect 3836 2067 3844 2076
rect 3967 2076 4673 2084
rect 4687 2076 4753 2084
rect 5967 2076 6153 2084
rect 1967 2056 2404 2064
rect 2787 2056 2833 2064
rect 3927 2056 3973 2064
rect 4747 2056 4813 2064
rect 4927 2056 5193 2064
rect 5507 2056 5773 2064
rect 627 2036 664 2044
rect 1147 2036 1193 2044
rect 1767 2036 1913 2044
rect 1927 2036 2293 2044
rect 2627 2036 2873 2044
rect 2887 2036 3153 2044
rect 3367 2036 3413 2044
rect 3587 2036 3633 2044
rect 3807 2036 3933 2044
rect 4627 2036 4833 2044
rect 4847 2036 4873 2044
rect 4887 2036 5313 2044
rect 6196 2044 6204 2073
rect 6216 2067 6224 2096
rect 6427 2096 6593 2104
rect 6747 2096 6933 2104
rect 6987 2096 7613 2104
rect 8196 2096 8613 2104
rect 8196 2087 8204 2096
rect 8627 2096 8653 2104
rect 8667 2096 8813 2104
rect 9367 2096 9613 2104
rect 9627 2096 10013 2104
rect 10487 2096 10533 2104
rect 10667 2096 10853 2104
rect 10867 2096 11033 2104
rect 11056 2096 11273 2104
rect 6447 2076 6533 2084
rect 6627 2076 6713 2084
rect 7187 2076 7353 2084
rect 7407 2076 7453 2084
rect 8047 2076 8133 2084
rect 8367 2076 8453 2084
rect 8487 2076 8653 2084
rect 8767 2076 8853 2084
rect 9207 2076 9353 2084
rect 9427 2076 9633 2084
rect 9687 2076 9833 2084
rect 11056 2084 11064 2096
rect 10527 2076 11064 2084
rect 6907 2056 7193 2064
rect 7447 2056 7593 2064
rect 8107 2056 8133 2064
rect 8187 2056 8213 2064
rect 8647 2056 8693 2064
rect 9116 2064 9124 2073
rect 9116 2056 9153 2064
rect 9387 2056 9493 2064
rect 9667 2056 9753 2064
rect 9847 2056 9873 2064
rect 10096 2056 10513 2064
rect 10096 2047 10104 2056
rect 6196 2036 6393 2044
rect 6947 2036 7453 2044
rect 8427 2036 8473 2044
rect 9907 2036 10033 2044
rect 10147 2036 10313 2044
rect 10327 2036 10373 2044
rect 10587 2036 10813 2044
rect 5667 2016 6173 2024
rect 10367 2016 10773 2024
rect 10807 2016 10833 2024
rect 6167 1996 6493 2004
rect 6227 1976 6413 1984
rect 1667 1956 1693 1964
rect 5987 1956 9153 1964
rect 2407 1916 2653 1924
rect 2667 1916 2693 1924
rect 4307 1916 5893 1924
rect 5107 1896 5493 1904
rect 1307 1876 3133 1884
rect 3147 1876 3593 1884
rect 3667 1876 4513 1884
rect 7347 1876 8873 1884
rect 8887 1876 9573 1884
rect 4067 1856 4453 1864
rect 4467 1856 4573 1864
rect 5287 1856 7133 1864
rect 8027 1856 8113 1864
rect 9827 1856 9873 1864
rect 10347 1856 10953 1864
rect 10967 1856 11093 1864
rect 947 1836 2593 1844
rect 3287 1836 4513 1844
rect 4527 1836 4773 1844
rect 5247 1836 5333 1844
rect 7907 1836 8124 1844
rect 1787 1816 1833 1824
rect 2496 1816 2513 1824
rect 2496 1807 2504 1816
rect 4027 1816 4393 1824
rect 4407 1816 4553 1824
rect 4567 1816 4753 1824
rect 5087 1816 5313 1824
rect 6127 1816 6453 1824
rect 6487 1816 6673 1824
rect 7567 1816 7653 1824
rect 8007 1816 8093 1824
rect 8116 1824 8124 1836
rect 8387 1836 8913 1844
rect 8927 1836 11293 1844
rect 8116 1816 8133 1824
rect 8147 1816 8373 1824
rect 8667 1816 8713 1824
rect 8727 1816 8973 1824
rect 9847 1816 9864 1824
rect 9856 1807 9864 1816
rect 10087 1816 10124 1824
rect 10116 1807 10124 1816
rect 10167 1816 10453 1824
rect 10527 1816 10553 1824
rect 10767 1816 10813 1824
rect 11007 1816 11173 1824
rect 11187 1816 11253 1824
rect 87 1796 493 1804
rect 1107 1796 1153 1804
rect 1167 1796 1273 1804
rect 1587 1796 1933 1804
rect 2547 1796 2753 1804
rect 2767 1796 2893 1804
rect 2947 1796 2973 1804
rect 3027 1796 3053 1804
rect 3507 1796 3873 1804
rect 3947 1796 3973 1804
rect 4207 1796 4233 1804
rect 4607 1796 5253 1804
rect 5747 1796 5933 1804
rect 5947 1796 6093 1804
rect 6467 1796 6533 1804
rect 7927 1796 8113 1804
rect 8167 1796 8253 1804
rect 8707 1796 8833 1804
rect 8847 1796 8873 1804
rect 9247 1796 9353 1804
rect 9567 1796 9593 1804
rect 9627 1796 9813 1804
rect 10387 1796 10573 1804
rect 10707 1796 11204 1804
rect 727 1776 853 1784
rect 867 1776 953 1784
rect 1827 1776 1853 1784
rect 2107 1776 2173 1784
rect 2447 1776 2513 1784
rect 2747 1776 2764 1784
rect 947 1756 1293 1764
rect 1367 1756 1393 1764
rect 1807 1756 2113 1764
rect 2287 1756 2553 1764
rect 2756 1747 2764 1776
rect 3187 1776 3233 1784
rect 3367 1776 3473 1784
rect 3727 1776 3953 1784
rect 4007 1776 4073 1784
rect 4267 1776 4433 1784
rect 5207 1776 5353 1784
rect 5667 1776 5713 1784
rect 5727 1776 5753 1784
rect 5847 1776 5993 1784
rect 6007 1776 6193 1784
rect 6207 1776 6213 1784
rect 6247 1776 6333 1784
rect 6487 1776 6493 1784
rect 6507 1776 6753 1784
rect 6767 1776 6933 1784
rect 6947 1776 7113 1784
rect 7127 1776 7293 1784
rect 7587 1776 7873 1784
rect 8347 1776 8553 1784
rect 8627 1776 8733 1784
rect 8827 1776 8833 1784
rect 8847 1776 8933 1784
rect 9167 1776 9193 1784
rect 9387 1776 9513 1784
rect 10076 1784 10084 1793
rect 9667 1776 10833 1784
rect 10867 1776 10973 1784
rect 11196 1784 11204 1796
rect 11196 1776 11233 1784
rect 3207 1756 3393 1764
rect 4367 1756 4653 1764
rect 5067 1756 5233 1764
rect 5807 1756 6633 1764
rect 7087 1756 7373 1764
rect 7407 1756 7553 1764
rect 7847 1756 8073 1764
rect 9507 1756 9593 1764
rect 10027 1756 10313 1764
rect 10327 1756 10513 1764
rect 10547 1756 10573 1764
rect 10807 1756 10833 1764
rect 10947 1756 11033 1764
rect 11047 1756 11293 1764
rect 927 1736 1013 1744
rect 1147 1736 1393 1744
rect 3127 1736 3193 1744
rect 3967 1736 4493 1744
rect 4547 1736 4773 1744
rect 7427 1736 9833 1744
rect 10767 1736 10793 1744
rect 167 1716 193 1724
rect 2567 1716 3553 1724
rect 6027 1716 6893 1724
rect 6907 1716 7693 1724
rect 7707 1716 9113 1724
rect 9347 1716 9773 1724
rect 9787 1716 9793 1724
rect 10787 1716 11253 1724
rect 107 1696 213 1704
rect 547 1696 673 1704
rect 687 1696 2053 1704
rect 2747 1696 2853 1704
rect 2947 1696 4193 1704
rect 4507 1696 4973 1704
rect 5287 1696 5473 1704
rect 6627 1696 8373 1704
rect 687 1676 773 1684
rect 2067 1676 4713 1684
rect 6967 1676 7153 1684
rect 7287 1676 9093 1684
rect 1627 1656 1973 1664
rect 1987 1656 2333 1664
rect 2587 1656 3033 1664
rect 3047 1656 3853 1664
rect 3867 1656 3993 1664
rect 4287 1656 4673 1664
rect 4687 1656 5233 1664
rect 8407 1656 8813 1664
rect 9427 1656 10033 1664
rect 10047 1656 10053 1664
rect 1087 1636 2573 1644
rect 3587 1636 3753 1644
rect 4367 1636 4473 1644
rect 4487 1636 4533 1644
rect 5467 1636 5753 1644
rect 6787 1636 6993 1644
rect 7727 1636 8313 1644
rect 8327 1636 8633 1644
rect 9467 1636 10073 1644
rect 627 1616 713 1624
rect 827 1616 1593 1624
rect 1607 1616 1953 1624
rect 1967 1616 2093 1624
rect 2147 1616 2153 1624
rect 2167 1616 2193 1624
rect 2207 1616 2353 1624
rect 2887 1616 3093 1624
rect 3247 1616 3553 1624
rect 3687 1616 4053 1624
rect 4087 1616 4473 1624
rect 4527 1616 5213 1624
rect 5307 1616 5953 1624
rect 6987 1616 7153 1624
rect 7207 1616 7473 1624
rect 7927 1616 8573 1624
rect 8627 1616 8873 1624
rect 9127 1616 9193 1624
rect 9307 1616 9593 1624
rect 9827 1616 10013 1624
rect 10067 1616 10253 1624
rect 10307 1616 10613 1624
rect 807 1596 873 1604
rect 1747 1596 1893 1604
rect 2107 1596 2433 1604
rect 2627 1596 2813 1604
rect 2827 1596 3044 1604
rect 427 1576 553 1584
rect 707 1576 853 1584
rect 867 1576 893 1584
rect 147 1556 193 1564
rect 916 1564 924 1593
rect 1387 1576 1433 1584
rect 1947 1576 2493 1584
rect 3036 1584 3044 1596
rect 3367 1596 3493 1604
rect 3507 1596 3593 1604
rect 3827 1596 3873 1604
rect 3887 1596 4093 1604
rect 4107 1596 4213 1604
rect 4387 1596 4493 1604
rect 4687 1596 4713 1604
rect 4767 1596 5044 1604
rect 5036 1587 5044 1596
rect 5067 1596 5093 1604
rect 5587 1596 5833 1604
rect 5987 1596 6033 1604
rect 6107 1596 6713 1604
rect 6787 1596 7253 1604
rect 7507 1596 7573 1604
rect 7647 1596 7893 1604
rect 8127 1596 8173 1604
rect 8207 1596 8473 1604
rect 8487 1596 8633 1604
rect 9167 1596 9213 1604
rect 9227 1596 9413 1604
rect 3036 1576 3073 1584
rect 5227 1576 5453 1584
rect 5467 1576 5513 1584
rect 247 1556 924 1564
rect 1707 1556 1873 1564
rect 1927 1556 1973 1564
rect 1987 1556 2073 1564
rect 2407 1556 2953 1564
rect 3027 1556 3333 1564
rect 4487 1556 5473 1564
rect 5536 1564 5544 1593
rect 5567 1576 5633 1584
rect 5827 1576 5853 1584
rect 7456 1584 7464 1593
rect 9616 1587 9624 1613
rect 9647 1596 9733 1604
rect 9747 1596 9793 1604
rect 10387 1596 10693 1604
rect 10707 1596 10773 1604
rect 10827 1596 11173 1604
rect 6507 1576 7444 1584
rect 7456 1576 7693 1584
rect 5536 1556 6053 1564
rect 6067 1556 6513 1564
rect 6647 1556 6733 1564
rect 7247 1556 7273 1564
rect 7436 1564 7444 1576
rect 8127 1576 8153 1584
rect 8707 1576 8893 1584
rect 8967 1576 9093 1584
rect 9107 1576 9333 1584
rect 9347 1576 9353 1584
rect 9407 1576 9453 1584
rect 10296 1584 10304 1593
rect 10296 1576 10413 1584
rect 10427 1576 10593 1584
rect 10927 1576 11013 1584
rect 7436 1556 7673 1564
rect 7967 1556 8133 1564
rect 8667 1556 8713 1564
rect 8867 1556 8993 1564
rect 9007 1556 9133 1564
rect 9147 1556 9653 1564
rect 10267 1556 10533 1564
rect 10547 1556 10753 1564
rect 11047 1556 11193 1564
rect 2967 1536 4253 1544
rect 4267 1536 4433 1544
rect 5007 1536 5253 1544
rect 6447 1536 6473 1544
rect 7167 1536 8113 1544
rect 2627 1496 2833 1504
rect 3127 1436 3153 1444
rect 3527 1436 3613 1444
rect 4307 1436 4513 1444
rect 4527 1436 5773 1444
rect 5787 1436 6013 1444
rect 10807 1416 10933 1424
rect 7067 1396 7493 1404
rect 8407 1396 8933 1404
rect 2107 1376 2153 1384
rect 6867 1376 7553 1384
rect 7787 1376 7893 1384
rect 8307 1376 9173 1384
rect 9667 1376 9973 1384
rect 10027 1376 11013 1384
rect 267 1356 413 1364
rect 1027 1356 1193 1364
rect 1207 1356 1493 1364
rect 1507 1356 3213 1364
rect 5487 1356 5733 1364
rect 7367 1356 8293 1364
rect 8307 1356 8913 1364
rect 9967 1356 10113 1364
rect 10547 1356 10713 1364
rect 207 1336 393 1344
rect 1167 1336 1184 1344
rect 176 1304 184 1333
rect 247 1316 433 1324
rect 627 1316 633 1324
rect 647 1316 673 1324
rect 727 1316 1093 1324
rect 1107 1316 1153 1324
rect 1176 1307 1184 1336
rect 1347 1336 1673 1344
rect 1687 1336 1933 1344
rect 2427 1336 3093 1344
rect 3107 1336 3173 1344
rect 3207 1336 3313 1344
rect 3527 1336 3773 1344
rect 5227 1336 5273 1344
rect 5347 1336 5533 1344
rect 6036 1336 6833 1344
rect 1327 1316 1433 1324
rect 1456 1316 1893 1324
rect 1456 1307 1464 1316
rect 1907 1316 2013 1324
rect 2047 1316 2593 1324
rect 2607 1316 2833 1324
rect 2847 1316 3633 1324
rect 3807 1316 3933 1324
rect 4207 1316 4273 1324
rect 4527 1316 4553 1324
rect 4607 1316 4693 1324
rect 4747 1316 4933 1324
rect 5047 1316 5233 1324
rect 5267 1316 5293 1324
rect 6036 1324 6044 1336
rect 7007 1336 7053 1344
rect 7567 1336 7793 1344
rect 7847 1336 7933 1344
rect 8467 1336 8493 1344
rect 8947 1336 8973 1344
rect 9287 1336 9453 1344
rect 9507 1336 9553 1344
rect 9987 1336 10033 1344
rect 10047 1336 10213 1344
rect 10227 1336 10293 1344
rect 10747 1336 10813 1344
rect 10916 1327 10924 1353
rect 10987 1336 11033 1344
rect 5527 1316 6044 1324
rect 6067 1316 6113 1324
rect 7127 1316 7173 1324
rect 7187 1316 7313 1324
rect 7827 1316 8053 1324
rect 8487 1316 8513 1324
rect 8827 1316 8993 1324
rect 10607 1316 10673 1324
rect 10967 1316 11013 1324
rect 176 1296 213 1304
rect 487 1296 693 1304
rect 747 1296 1133 1304
rect 1247 1296 1413 1304
rect 1607 1296 2313 1304
rect 2327 1296 2333 1304
rect 2387 1296 2493 1304
rect 3307 1296 3333 1304
rect 3507 1296 3573 1304
rect 4227 1296 4253 1304
rect 4547 1296 5793 1304
rect 5807 1296 5993 1304
rect 6087 1296 6193 1304
rect 6207 1296 6413 1304
rect 6467 1296 6573 1304
rect 6587 1296 6753 1304
rect 8447 1296 8533 1304
rect 8707 1296 8773 1304
rect 9047 1296 9213 1304
rect 9307 1296 9693 1304
rect 9787 1296 9953 1304
rect 10347 1296 10453 1304
rect 187 1276 353 1284
rect 667 1276 713 1284
rect 1147 1276 1313 1284
rect 1927 1276 2253 1284
rect 2267 1276 2593 1284
rect 3287 1276 3333 1284
rect 4327 1276 4573 1284
rect 6347 1276 6533 1284
rect 8967 1276 9633 1284
rect 9747 1276 9873 1284
rect 10027 1276 10093 1284
rect 10447 1276 10593 1284
rect 10716 1284 10724 1313
rect 10716 1276 10733 1284
rect 10887 1276 11173 1284
rect 167 1256 213 1264
rect 687 1256 733 1264
rect 967 1256 993 1264
rect 1007 1256 2113 1264
rect 2167 1256 2353 1264
rect 2447 1256 2993 1264
rect 3007 1256 3533 1264
rect 4307 1256 4913 1264
rect 5767 1256 7073 1264
rect 7107 1256 7404 1264
rect 1127 1236 1153 1244
rect 1747 1236 2533 1244
rect 2547 1236 2553 1244
rect 2567 1236 2793 1244
rect 2807 1236 3013 1244
rect 4067 1236 4413 1244
rect 4427 1236 4693 1244
rect 4707 1236 5593 1244
rect 5927 1236 7373 1244
rect 7396 1244 7404 1256
rect 9027 1256 9253 1264
rect 9287 1256 10093 1264
rect 10107 1256 10253 1264
rect 10267 1256 10713 1264
rect 10727 1256 10993 1264
rect 7396 1236 9473 1244
rect 10247 1236 10653 1244
rect 10707 1236 10933 1244
rect 1027 1216 2093 1224
rect 2107 1216 2573 1224
rect 2587 1216 3233 1224
rect 3247 1216 3513 1224
rect 3567 1216 5393 1224
rect 5407 1216 5473 1224
rect 6707 1216 7333 1224
rect 10467 1216 10753 1224
rect 3187 1196 3993 1204
rect 5987 1196 7113 1204
rect 9747 1196 10513 1204
rect 2907 1176 3553 1184
rect 3587 1176 4933 1184
rect 6607 1176 6713 1184
rect 8207 1176 8953 1184
rect 10507 1176 10693 1184
rect 487 1156 693 1164
rect 707 1156 1173 1164
rect 1427 1156 1453 1164
rect 1467 1156 1733 1164
rect 2327 1156 3493 1164
rect 3507 1156 3673 1164
rect 4247 1156 4733 1164
rect 4747 1156 4893 1164
rect 6067 1156 6133 1164
rect 6367 1156 6433 1164
rect 6667 1156 6693 1164
rect 6827 1156 7053 1164
rect 8087 1156 8453 1164
rect 8467 1156 8493 1164
rect 8787 1156 9273 1164
rect 10007 1156 10973 1164
rect 10987 1156 11053 1164
rect 627 1136 913 1144
rect 927 1136 1393 1144
rect 1407 1136 1433 1144
rect 1507 1136 1653 1144
rect 1667 1136 1793 1144
rect 1907 1136 2313 1144
rect 2327 1136 2613 1144
rect 3067 1136 3293 1144
rect 4047 1136 4233 1144
rect 4727 1136 4873 1144
rect 4927 1136 5053 1144
rect 5467 1136 5653 1144
rect 5667 1136 6193 1144
rect 6427 1136 6673 1144
rect 6687 1136 6933 1144
rect 7147 1136 7173 1144
rect 7607 1136 7633 1144
rect 7667 1136 7753 1144
rect 7787 1136 8193 1144
rect 8487 1136 8533 1144
rect 8567 1136 8933 1144
rect 9247 1136 9473 1144
rect 9927 1136 10213 1144
rect 10447 1136 10473 1144
rect 11007 1136 11133 1144
rect 11147 1136 11213 1144
rect 747 1116 773 1124
rect 1247 1116 1373 1124
rect 1387 1116 1593 1124
rect 1627 1116 2053 1124
rect 2087 1116 2104 1124
rect 247 1096 393 1104
rect 407 1096 413 1104
rect 427 1096 453 1104
rect 516 1104 524 1113
rect 516 1096 753 1104
rect 767 1096 953 1104
rect 1136 1104 1144 1113
rect 1136 1096 1253 1104
rect 1647 1096 1853 1104
rect 2096 1104 2104 1116
rect 2127 1116 2293 1124
rect 2307 1116 2373 1124
rect 2587 1116 2973 1124
rect 3087 1116 3573 1124
rect 3807 1116 4393 1124
rect 4487 1116 4693 1124
rect 4827 1116 5433 1124
rect 5707 1116 5873 1124
rect 6107 1116 6364 1124
rect 2096 1096 2553 1104
rect 2847 1096 3033 1104
rect 3087 1096 3133 1104
rect 3247 1096 3273 1104
rect 3407 1096 3553 1104
rect 3627 1096 4253 1104
rect 3816 1087 3824 1096
rect 4267 1096 5213 1104
rect 5427 1096 5453 1104
rect 6127 1096 6293 1104
rect 6356 1104 6364 1116
rect 6387 1116 6573 1124
rect 6596 1116 6633 1124
rect 6356 1096 6533 1104
rect 6596 1104 6604 1116
rect 6827 1116 6853 1124
rect 6907 1116 8164 1124
rect 6567 1096 6604 1104
rect 6667 1096 6693 1104
rect 6927 1096 7013 1104
rect 7427 1096 7453 1104
rect 8156 1104 8164 1116
rect 8187 1116 8713 1124
rect 8947 1116 9233 1124
rect 10207 1116 10233 1124
rect 10247 1116 10313 1124
rect 10407 1116 10413 1124
rect 10427 1116 10453 1124
rect 10527 1116 10653 1124
rect 10727 1116 10953 1124
rect 8156 1096 8213 1104
rect 8247 1096 8273 1104
rect 8516 1096 8673 1104
rect 507 1076 673 1084
rect 987 1076 1013 1084
rect 1447 1076 1873 1084
rect 2287 1076 2393 1084
rect 2407 1076 2813 1084
rect 2827 1076 2873 1084
rect 3147 1076 3513 1084
rect 3527 1076 3533 1084
rect 3867 1076 4533 1084
rect 6407 1076 7033 1084
rect 7367 1076 7393 1084
rect 7927 1076 7993 1084
rect 8516 1084 8524 1096
rect 8927 1096 8973 1104
rect 9187 1096 9253 1104
rect 9527 1096 9773 1104
rect 10347 1096 10473 1104
rect 8227 1076 8524 1084
rect 8547 1076 8693 1084
rect 9767 1076 10273 1084
rect 1847 1056 1893 1064
rect 3027 1056 3833 1064
rect 3847 1056 5333 1064
rect 5347 1056 5373 1064
rect 6587 1056 7153 1064
rect 7167 1056 8173 1064
rect 8767 1056 10373 1064
rect 2067 1036 3313 1044
rect 6207 1036 6813 1044
rect 7467 1036 9973 1044
rect 3567 1016 4473 1024
rect 4487 1016 4493 1024
rect 5447 1016 6353 1024
rect 6567 1016 9593 1024
rect 1707 996 2853 1004
rect 2867 996 3733 1004
rect 5287 996 7353 1004
rect 7767 996 8273 1004
rect 8287 996 8793 1004
rect 6367 976 6613 984
rect 6627 976 6873 984
rect 9727 976 9773 984
rect 1947 956 2133 964
rect 2147 956 2813 964
rect 2827 956 3393 964
rect 8047 956 8773 964
rect 2367 936 3793 944
rect 4427 936 7373 944
rect 9267 936 10053 944
rect 2567 916 2793 924
rect 3227 916 4053 924
rect 6047 916 7353 924
rect 7447 916 7533 924
rect 7907 916 7933 924
rect 7987 916 8033 924
rect 9647 916 10353 924
rect 287 896 693 904
rect 707 896 1113 904
rect 1127 896 1353 904
rect 1367 896 2153 904
rect 2627 896 4913 904
rect 6287 896 6353 904
rect 7127 896 7553 904
rect 7567 896 8033 904
rect 8387 896 8464 904
rect 947 876 993 884
rect 1887 876 3093 884
rect 3107 876 3773 884
rect 4967 876 5193 884
rect 5207 876 5433 884
rect 5527 876 7393 884
rect 7476 876 8424 884
rect 216 856 413 864
rect 216 844 224 856
rect 747 856 1753 864
rect 2027 856 2053 864
rect 2767 856 2853 864
rect 3767 856 4724 864
rect 207 836 224 844
rect 247 836 564 844
rect 147 816 213 824
rect 487 816 533 824
rect 556 824 564 836
rect 907 836 944 844
rect 556 816 673 824
rect 787 816 913 824
rect 936 824 944 836
rect 1207 836 1433 844
rect 1447 836 1993 844
rect 2007 836 2093 844
rect 2167 836 2573 844
rect 2587 836 2933 844
rect 3187 836 3273 844
rect 3327 836 3833 844
rect 4227 836 4253 844
rect 4307 836 4453 844
rect 4467 836 4513 844
rect 4716 844 4724 856
rect 4747 856 4993 864
rect 5047 856 6253 864
rect 7007 856 7033 864
rect 7147 856 7224 864
rect 7216 847 7224 856
rect 7367 856 7453 864
rect 7476 864 7484 876
rect 7467 856 7484 864
rect 7507 856 8073 864
rect 8227 856 8313 864
rect 8416 864 8424 876
rect 8456 867 8464 896
rect 8507 896 9413 904
rect 10227 896 10533 904
rect 9327 876 9393 884
rect 10307 876 11233 884
rect 8416 856 8444 864
rect 8436 847 8444 856
rect 8587 856 9133 864
rect 9187 856 9353 864
rect 9587 856 10273 864
rect 10347 856 10373 864
rect 10927 856 11073 864
rect 4716 836 4753 844
rect 4887 836 5253 844
rect 5587 836 6013 844
rect 6027 836 6093 844
rect 7116 836 7153 844
rect 936 816 1173 824
rect 1767 816 1853 824
rect 1987 816 2333 824
rect 2387 816 2473 824
rect 2847 816 3033 824
rect 3087 816 3113 824
rect 3207 816 3293 824
rect 3547 816 4053 824
rect 4287 816 4413 824
rect 4547 816 4713 824
rect 5027 816 5053 824
rect 5067 816 5413 824
rect 5427 816 5473 824
rect 5607 816 5993 824
rect 7116 824 7124 836
rect 7387 836 7433 844
rect 7487 836 7573 844
rect 8247 836 8393 844
rect 8807 836 9373 844
rect 9427 836 10073 844
rect 10247 836 10413 844
rect 11147 836 11273 844
rect 6047 816 7124 824
rect 7136 816 7173 824
rect 967 796 1013 804
rect 1187 796 1233 804
rect 1487 796 1633 804
rect 1887 796 1993 804
rect 2027 796 2073 804
rect 2087 796 3013 804
rect 3027 796 3033 804
rect 3067 796 3173 804
rect 3267 796 3513 804
rect 3847 796 5173 804
rect 5187 796 5233 804
rect 5247 796 5493 804
rect 5807 796 6073 804
rect 6087 796 6333 804
rect 6507 796 6733 804
rect 7136 804 7144 816
rect 7427 816 7593 824
rect 8007 816 8693 824
rect 8907 816 9153 824
rect 9367 816 10293 824
rect 6767 796 7144 804
rect 7167 796 8933 804
rect 8947 796 9833 804
rect 10307 796 10393 804
rect 11067 796 11133 804
rect 707 776 753 784
rect 767 776 853 784
rect 1227 776 2033 784
rect 3167 776 3333 784
rect 3347 776 3573 784
rect 4047 776 4073 784
rect 4087 776 4213 784
rect 4807 776 5733 784
rect 6307 776 6673 784
rect 6687 776 6773 784
rect 6787 776 6953 784
rect 7407 776 8193 784
rect 8207 776 8373 784
rect 8507 776 9613 784
rect 667 756 1573 764
rect 2127 756 2344 764
rect 187 736 433 744
rect 1167 736 1293 744
rect 1307 736 1633 744
rect 1667 736 2213 744
rect 2336 744 2344 756
rect 2367 756 2393 764
rect 4507 756 4673 764
rect 4687 756 5113 764
rect 5267 756 5933 764
rect 6007 756 6633 764
rect 6647 756 6833 764
rect 7267 756 7713 764
rect 8687 756 9333 764
rect 9947 756 10193 764
rect 2336 736 5573 744
rect 5727 736 6113 744
rect 7207 736 8913 744
rect 9627 736 10533 744
rect 447 716 1724 724
rect 1007 696 1693 704
rect 1716 704 1724 716
rect 2587 716 5693 724
rect 5707 716 5733 724
rect 6127 716 7893 724
rect 7907 716 8273 724
rect 8907 716 9453 724
rect 10327 716 10553 724
rect 1716 696 3013 704
rect 3027 696 5193 704
rect 5207 696 6153 704
rect 7267 696 7313 704
rect 7347 696 7733 704
rect 7747 696 8173 704
rect 8687 696 9833 704
rect 1847 676 1893 684
rect 2127 676 2373 684
rect 2387 676 3973 684
rect 4027 676 4193 684
rect 4407 676 5253 684
rect 5767 676 6653 684
rect 6667 676 6993 684
rect 7007 676 8833 684
rect 9167 676 9353 684
rect 9367 676 9393 684
rect 10987 676 11013 684
rect 507 656 553 664
rect 567 656 673 664
rect 687 656 1413 664
rect 1867 656 2093 664
rect 2167 656 3273 664
rect 3347 656 3533 664
rect 3787 656 4213 664
rect 4227 656 4273 664
rect 5227 656 5313 664
rect 5676 656 5933 664
rect 247 636 453 644
rect 547 636 953 644
rect 1387 636 1413 644
rect 1467 636 1613 644
rect 1667 636 1853 644
rect 1967 636 2493 644
rect 2507 636 3073 644
rect 3087 636 3213 644
rect 3327 636 3473 644
rect 3536 636 3553 644
rect 3536 627 3544 636
rect 3567 636 3773 644
rect 3976 636 4673 644
rect 227 616 253 624
rect 487 616 553 624
rect 667 616 733 624
rect 1407 616 1773 624
rect 1787 616 2153 624
rect 2316 616 2813 624
rect 2316 607 2324 616
rect 2827 616 2953 624
rect 3647 616 3953 624
rect 3976 624 3984 636
rect 5676 644 5684 656
rect 7067 656 7273 664
rect 7287 656 7473 664
rect 7507 656 8093 664
rect 8167 656 8193 664
rect 8407 656 8593 664
rect 8747 656 9333 664
rect 10787 656 10993 664
rect 11027 656 11233 664
rect 4967 636 5684 644
rect 5707 636 5753 644
rect 7047 636 7233 644
rect 7547 636 8373 644
rect 9047 636 9113 644
rect 9327 636 9373 644
rect 10267 636 10513 644
rect 10527 636 10533 644
rect 10627 636 11033 644
rect 11047 636 11193 644
rect 3967 616 3984 624
rect 4007 616 4073 624
rect 4727 616 4933 624
rect 5467 616 5673 624
rect 7516 624 7524 633
rect 7516 616 7713 624
rect 8147 616 8293 624
rect 8587 616 8613 624
rect 8647 616 8693 624
rect 8727 616 9133 624
rect 9147 616 9573 624
rect 10596 624 10604 633
rect 10327 616 10804 624
rect 10796 607 10804 616
rect 1447 596 1953 604
rect 2467 596 2593 604
rect 2887 596 3293 604
rect 4547 596 4733 604
rect 4747 596 4973 604
rect 5027 596 10313 604
rect 10527 596 10753 604
rect 927 576 1673 584
rect 1687 576 2553 584
rect 5107 576 5773 584
rect 5787 576 7113 584
rect 7887 576 8113 584
rect 9407 576 9633 584
rect 10587 576 10613 584
rect 987 556 1193 564
rect 1207 556 1933 564
rect 2987 556 5713 564
rect 8107 556 8573 564
rect 9387 556 9433 564
rect 6207 536 10273 544
rect 10327 496 10493 504
rect 6027 476 9293 484
rect 9667 476 10133 484
rect 8087 456 8373 464
rect 8387 456 9493 464
rect 4747 436 4873 444
rect 10647 436 10733 444
rect 10747 436 11173 444
rect 507 416 513 424
rect 527 416 2293 424
rect 3187 416 4693 424
rect 4707 416 4753 424
rect 4987 416 5393 424
rect 5487 416 10893 424
rect 10987 416 11013 424
rect 11047 416 11253 424
rect 1387 396 1453 404
rect 2487 396 2573 404
rect 3067 396 3953 404
rect 3967 396 4373 404
rect 4387 396 4413 404
rect 4507 396 4933 404
rect 5007 396 6133 404
rect 6987 396 7633 404
rect 9687 396 9833 404
rect 9847 396 9893 404
rect 10187 396 10253 404
rect 10267 396 10273 404
rect 11167 396 11193 404
rect 1267 376 1373 384
rect 1427 376 1613 384
rect 1667 376 1933 384
rect 2067 376 2233 384
rect 2247 376 2533 384
rect 2547 376 2793 384
rect 2947 376 3133 384
rect 3147 376 3253 384
rect 3487 376 3753 384
rect 3807 376 3993 384
rect 4007 376 4353 384
rect 4947 376 5433 384
rect 5447 376 5613 384
rect 6107 376 6173 384
rect 6767 376 7353 384
rect 7887 376 7913 384
rect 8247 376 8553 384
rect 9547 376 9733 384
rect 9867 376 10933 384
rect 10987 376 11013 384
rect 11127 376 11153 384
rect 216 347 224 373
rect 247 356 533 364
rect 616 356 713 364
rect 616 344 624 356
rect 767 356 913 364
rect 927 356 933 364
rect 1167 356 1324 364
rect 487 336 624 344
rect 647 336 693 344
rect 1316 344 1324 356
rect 1347 356 1393 364
rect 1607 356 1873 364
rect 1887 356 1973 364
rect 2116 356 2313 364
rect 2116 347 2124 356
rect 3027 356 3213 364
rect 4067 356 4213 364
rect 4367 356 4453 364
rect 4507 356 4533 364
rect 4867 356 5953 364
rect 6667 356 8573 364
rect 10007 356 10173 364
rect 10187 356 10653 364
rect 10667 356 10713 364
rect 10967 356 11033 364
rect 11187 356 11333 364
rect 1316 336 1633 344
rect 1687 336 1824 344
rect 407 316 513 324
rect 527 316 1793 324
rect 1816 324 1824 336
rect 2787 336 3193 344
rect 3247 336 3964 344
rect 1816 316 1893 324
rect 1907 316 2053 324
rect 2107 316 2153 324
rect 2307 316 2313 324
rect 2327 316 2473 324
rect 3507 316 3833 324
rect 3956 324 3964 336
rect 3987 336 4033 344
rect 4047 336 4193 344
rect 4247 336 4953 344
rect 5327 336 5693 344
rect 5767 336 5913 344
rect 6247 336 6413 344
rect 6747 336 6853 344
rect 6907 336 6993 344
rect 7007 336 7113 344
rect 7687 336 7953 344
rect 8027 336 8153 344
rect 8627 336 8813 344
rect 9027 336 9113 344
rect 9287 336 9333 344
rect 9727 336 9873 344
rect 9907 336 10333 344
rect 10347 336 10353 344
rect 10907 336 10993 344
rect 3956 316 5013 324
rect 5027 316 5453 324
rect 5707 316 5893 324
rect 7427 316 8853 324
rect 8867 316 9313 324
rect 9767 316 9993 324
rect 10207 316 10953 324
rect 187 296 453 304
rect 1567 296 1913 304
rect 1927 296 2033 304
rect 2047 296 3273 304
rect 3287 296 3973 304
rect 7167 296 8193 304
rect 8847 296 9033 304
rect 9307 296 9793 304
rect 10707 296 10733 304
rect 7007 276 8473 284
rect 9087 276 10473 284
rect 6747 256 7613 264
rect 10067 256 10153 264
rect 747 236 873 244
rect 3907 236 4473 244
rect 6047 236 7613 244
rect 7907 236 8133 244
rect 8456 236 9053 244
rect 2967 216 3853 224
rect 4147 216 4713 224
rect 5347 216 5753 224
rect 8456 224 8464 236
rect 9707 236 9833 244
rect 6527 216 8464 224
rect 8487 216 9853 224
rect 927 196 2213 204
rect 2287 196 2933 204
rect 3747 196 5093 204
rect 5107 196 5493 204
rect 5507 196 6593 204
rect 7627 196 9813 204
rect 9867 196 10713 204
rect 10727 196 11353 204
rect 227 176 413 184
rect 1147 176 1293 184
rect 1387 176 1573 184
rect 1847 176 2013 184
rect 2507 176 2713 184
rect 2727 176 2973 184
rect 2987 176 3153 184
rect 3427 176 3453 184
rect 3887 176 4033 184
rect 4327 176 4553 184
rect 4596 176 4813 184
rect 447 156 653 164
rect 967 156 1013 164
rect 1027 156 1993 164
rect 2007 156 2553 164
rect 2567 156 3113 164
rect 3127 156 3193 164
rect 3207 156 3473 164
rect 4087 156 4313 164
rect 4596 164 4604 176
rect 4847 176 5073 184
rect 5527 176 5713 184
rect 5807 176 6253 184
rect 6267 176 6493 184
rect 7407 176 7533 184
rect 7707 176 8993 184
rect 9827 176 10873 184
rect 10927 176 10973 184
rect 11107 176 11193 184
rect 4367 156 4604 164
rect 4627 156 5533 164
rect 5767 156 6153 164
rect 6767 156 7133 164
rect 7207 156 7933 164
rect 8007 156 8253 164
rect 8287 156 8813 164
rect 8827 156 10173 164
rect 10547 156 10753 164
rect 10767 156 10833 164
rect 10847 156 10933 164
rect 907 136 1113 144
rect 2487 136 2593 144
rect 5127 136 5313 144
rect 5536 136 6053 144
rect 687 116 813 124
rect 1987 116 2253 124
rect 4047 116 4093 124
rect 4387 116 4593 124
rect 4607 116 4793 124
rect 5536 124 5544 136
rect 6787 136 6973 144
rect 7667 136 7893 144
rect 7967 136 8433 144
rect 8447 136 8633 144
rect 8687 136 8713 144
rect 8787 136 9353 144
rect 10307 136 10853 144
rect 11187 136 11213 144
rect 5067 116 5544 124
rect 5567 116 5773 124
rect 6567 116 6713 124
rect 6887 116 7173 124
rect 7227 116 7373 124
rect 7387 116 7413 124
rect 8047 116 9153 124
rect 9167 116 9673 124
rect 10087 116 10213 124
rect 10527 116 10813 124
rect 2227 96 2693 104
rect 2707 96 3053 104
rect 7636 104 7644 113
rect 6287 96 7644 104
rect 10047 96 10453 104
rect 6087 76 9013 84
rect 6367 16 6433 24
use INVX1  _1744_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304789
transform -1 0 4590 0 1 10810
box -12 -8 72 252
use NAND2X1  _1745_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304996
transform 1 0 4350 0 -1 11290
box -12 -8 92 252
use OAI21X1  _1746_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305162
transform -1 0 4390 0 1 10810
box -12 -8 112 252
use INVX1  _1747_
timestamp 1728304789
transform -1 0 5830 0 -1 11290
box -12 -8 72 252
use NAND2X1  _1748_
timestamp 1728304996
transform 1 0 6710 0 -1 11290
box -12 -8 92 252
use OAI21X1  _1749_
timestamp 1728305162
transform 1 0 6450 0 -1 11290
box -12 -8 112 252
use INVX1  _1750_
timestamp 1728304789
transform 1 0 5310 0 -1 11290
box -12 -8 72 252
use NAND2X1  _1751_
timestamp 1728304996
transform 1 0 6950 0 -1 11290
box -12 -8 92 252
use OAI21X1  _1752_
timestamp 1728305162
transform 1 0 5510 0 -1 11290
box -12 -8 112 252
use INVX1  _1753_
timestamp 1728304789
transform 1 0 7670 0 1 10810
box -12 -8 72 252
use NAND2X1  _1754_
timestamp 1728304996
transform -1 0 7250 0 -1 11290
box -12 -8 92 252
use OAI21X1  _1755_
timestamp 1728305162
transform -1 0 7510 0 1 10810
box -12 -8 112 252
use INVX8  _1756_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304916
transform -1 0 6610 0 1 1210
box -12 -8 133 252
use OR2X2  _1757_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305284
transform 1 0 7150 0 1 10810
box -12 -8 112 252
use OAI21X1  _1758_
timestamp 1728305162
transform 1 0 6930 0 -1 10810
box -12 -8 112 252
use INVX1  _1759_
timestamp 1728304789
transform -1 0 3230 0 -1 10810
box -12 -8 72 252
use INVX1  _1760_
timestamp 1728304789
transform 1 0 2470 0 -1 11290
box -12 -8 72 252
use NAND2X1  _1761_
timestamp 1728304996
transform 1 0 7410 0 -1 11290
box -12 -8 92 252
use OAI21X1  _1762_
timestamp 1728305162
transform 1 0 2670 0 -1 11290
box -12 -8 112 252
use INVX1  _1763_
timestamp 1728304789
transform -1 0 8370 0 1 9850
box -12 -8 72 252
use NAND2X1  _1764_
timestamp 1728304996
transform -1 0 8210 0 1 10810
box -12 -8 92 252
use OAI21X1  _1765_
timestamp 1728305162
transform -1 0 8210 0 -1 10330
box -12 -8 112 252
use MUX2X1  _1766_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304958
transform -1 0 8050 0 -1 9370
box -12 -8 131 252
use INVX1  _1767_
timestamp 1728304789
transform -1 0 7970 0 -1 6010
box -12 -8 72 252
use INVX1  _1768_
timestamp 1728304789
transform -1 0 5870 0 1 4090
box -12 -8 72 252
use INVX1  _1769_
timestamp 1728304789
transform 1 0 3270 0 1 2170
box -12 -8 72 252
use INVX1  _1770_
timestamp 1728304789
transform 1 0 10910 0 1 2170
box -12 -8 72 252
use INVX1  _1771_
timestamp 1728304789
transform 1 0 11170 0 1 1210
box -12 -8 72 252
use NAND2X1  _1772_
timestamp 1728304996
transform 1 0 10910 0 1 2650
box -12 -8 92 252
use NAND2X1  _1773_
timestamp 1728304996
transform 1 0 10430 0 1 2170
box -12 -8 92 252
use NOR2X1  _1774_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305106
transform 1 0 10810 0 1 3130
box -12 -8 92 252
use INVX2  _1775_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304826
transform -1 0 9650 0 1 4090
box -12 -8 72 252
use NAND2X1  _1776_
timestamp 1728304996
transform 1 0 9670 0 -1 4570
box -12 -8 92 252
use INVX4  _1777_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304878
transform -1 0 8910 0 -1 5530
box -12 -8 92 252
use NAND2X1  _1778_
timestamp 1728304996
transform -1 0 11090 0 -1 3130
box -12 -8 92 252
use INVX1  _1779_
timestamp 1728304789
transform 1 0 10270 0 -1 250
box -12 -8 72 252
use INVX1  _1780_
timestamp 1728304789
transform 1 0 11030 0 1 1690
box -12 -8 72 252
use NAND2X1  _1781_
timestamp 1728304996
transform -1 0 11090 0 -1 2650
box -12 -8 92 252
use NOR2X1  _1782_
timestamp 1728305106
transform -1 0 11350 0 1 3610
box -12 -8 92 252
use OAI21X1  _1783_
timestamp 1728305162
transform -1 0 10150 0 -1 3610
box -12 -8 112 252
use AND2X2  _1784_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304163
transform 1 0 10670 0 1 2170
box -12 -8 112 252
use NOR2X1  _1785_
timestamp 1728305106
transform 1 0 11010 0 -1 2170
box -12 -8 92 252
use NAND2X1  _1786_
timestamp 1728304996
transform -1 0 10390 0 -1 2650
box -12 -8 92 252
use INVX2  _1787_
timestamp 1728304826
transform 1 0 9350 0 -1 250
box -12 -8 72 252
use NAND2X1  _1788_
timestamp 1728304996
transform 1 0 10630 0 -1 4570
box -12 -8 92 252
use OAI21X1  _1789_
timestamp 1728305162
transform -1 0 9550 0 -1 4090
box -12 -8 112 252
use NOR2X1  _1790_
timestamp 1728305106
transform -1 0 10910 0 1 3610
box -12 -8 92 252
use INVX1  _1791_
timestamp 1728304789
transform 1 0 11050 0 1 3610
box -12 -8 72 252
use NOR2X1  _1792_
timestamp 1728305106
transform 1 0 5770 0 -1 3610
box -12 -8 92 252
use AOI22X1  _1793_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304278
transform 1 0 5490 0 -1 3610
box -14 -8 132 252
use INVX1  _1794_
timestamp 1728304789
transform -1 0 5090 0 1 3130
box -12 -8 72 252
use INVX1  _1795_
timestamp 1728304789
transform 1 0 3850 0 -1 3610
box -12 -8 72 252
use NAND2X1  _1796_
timestamp 1728304996
transform 1 0 4290 0 -1 3610
box -12 -8 92 252
use OAI22X1  _1797_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305200
transform -1 0 4930 0 1 3610
box -12 -8 132 252
use NAND2X1  _1798_
timestamp 1728304996
transform -1 0 11210 0 1 2170
box -12 -8 92 252
use NOR3X1  _1799_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728303224
transform -1 0 11190 0 1 4090
box -12 -8 192 252
use NOR2X1  _1800_
timestamp 1728305106
transform -1 0 10630 0 -1 2650
box -12 -8 92 252
use NOR2X1  _1801_
timestamp 1728305106
transform -1 0 10290 0 1 2170
box -12 -8 92 252
use NAND2X1  _1802_
timestamp 1728304996
transform 1 0 10090 0 -1 2650
box -12 -8 92 252
use NOR2X1  _1803_
timestamp 1728305106
transform 1 0 10350 0 1 3130
box -12 -8 92 252
use NAND2X1  _1804_
timestamp 1728304996
transform 1 0 10330 0 -1 3130
box -12 -8 92 252
use NAND2X1  _1805_
timestamp 1728304996
transform -1 0 10210 0 -1 4570
box -12 -8 92 252
use OAI21X1  _1806_
timestamp 1728305162
transform 1 0 10090 0 1 3130
box -12 -8 112 252
use OAI21X1  _1807_
timestamp 1728305162
transform -1 0 10270 0 -1 4090
box -12 -8 112 252
use NAND2X1  _1808_
timestamp 1728304996
transform -1 0 10570 0 -1 250
box -12 -8 92 252
use NOR2X1  _1809_
timestamp 1728305106
transform -1 0 11230 0 -1 4090
box -12 -8 92 252
use NAND2X1  _1810_
timestamp 1728304996
transform -1 0 6390 0 1 3610
box -12 -8 92 252
use AND2X2  _1811_
timestamp 1728304163
transform -1 0 11330 0 -1 1690
box -12 -8 112 252
use NAND2X1  _1812_
timestamp 1728304996
transform -1 0 10370 0 -1 2170
box -12 -8 92 252
use INVX1  _1813_
timestamp 1728304789
transform -1 0 7850 0 1 2650
box -12 -8 72 252
use NAND2X1  _1814_
timestamp 1728304996
transform -1 0 7710 0 1 3130
box -12 -8 92 252
use NOR2X1  _1815_
timestamp 1728305106
transform -1 0 11110 0 -1 3610
box -12 -8 92 252
use INVX2  _1816_
timestamp 1728304826
transform -1 0 7750 0 1 4090
box -12 -8 72 252
use NOR2X1  _1817_
timestamp 1728305106
transform 1 0 6810 0 -1 3130
box -12 -8 92 252
use INVX1  _1818_
timestamp 1728304789
transform 1 0 6770 0 -1 3610
box -12 -8 72 252
use NAND3X1  _1819_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305047
transform 1 0 6270 0 -1 3610
box -12 -8 112 252
use NAND2X1  _1820_
timestamp 1728304996
transform 1 0 10450 0 1 2650
box -12 -8 92 252
use NOR2X1  _1821_
timestamp 1728305106
transform -1 0 6890 0 1 3610
box -12 -8 92 252
use NOR2X1  _1822_
timestamp 1728305106
transform 1 0 11250 0 -1 2170
box -12 -8 92 252
use NAND2X1  _1823_
timestamp 1728304996
transform -1 0 10150 0 -1 2170
box -12 -8 92 252
use NOR2X1  _1824_
timestamp 1728305106
transform 1 0 7410 0 1 4570
box -12 -8 92 252
use NOR2X1  _1825_
timestamp 1728305106
transform 1 0 6610 0 -1 4090
box -12 -8 92 252
use NOR2X1  _1826_
timestamp 1728305106
transform 1 0 11050 0 1 3130
box -12 -8 92 252
use NAND2X1  _1827_
timestamp 1728304996
transform -1 0 7550 0 -1 3610
box -12 -8 92 252
use NAND3X1  _1828_
timestamp 1728305047
transform 1 0 11230 0 1 1690
box -12 -8 112 252
use INVX1  _1829_
timestamp 1728304789
transform -1 0 7550 0 -1 5530
box -12 -8 72 252
use NAND2X1  _1830_
timestamp 1728304996
transform 1 0 7650 0 1 5050
box -12 -8 92 252
use NOR2X1  _1831_
timestamp 1728305106
transform 1 0 10770 0 -1 1690
box -12 -8 92 252
use NAND2X1  _1832_
timestamp 1728304996
transform 1 0 10770 0 -1 2170
box -12 -8 92 252
use OAI21X1  _1833_
timestamp 1728305162
transform 1 0 7310 0 -1 4090
box -12 -8 112 252
use INVX1  _1834_
timestamp 1728304789
transform -1 0 7170 0 -1 4090
box -12 -8 72 252
use NAND3X1  _1835_
timestamp 1728305047
transform -1 0 6650 0 1 3610
box -12 -8 112 252
use NOR2X1  _1836_
timestamp 1728305106
transform -1 0 6170 0 1 3610
box -12 -8 92 252
use NAND2X1  _1837_
timestamp 1728304996
transform -1 0 5710 0 1 3610
box -12 -8 92 252
use AOI21X1  _1838_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304211
transform 1 0 5370 0 1 3610
box -12 -8 112 252
use OAI21X1  _1839_
timestamp 1728305162
transform 1 0 5930 0 -1 4090
box -12 -8 112 252
use INVX1  _1840_
timestamp 1728304789
transform -1 0 8190 0 -1 7450
box -12 -8 72 252
use INVX2  _1841_
timestamp 1728304826
transform -1 0 5110 0 1 6010
box -12 -8 72 252
use NOR2X1  _1842_
timestamp 1728305106
transform -1 0 7010 0 1 4570
box -12 -8 92 252
use INVX2  _1843_
timestamp 1728304826
transform 1 0 7270 0 -1 4570
box -12 -8 72 252
use INVX4  _1844_
timestamp 1728304878
transform -1 0 10390 0 1 4090
box -12 -8 92 252
use NAND2X1  _1845_
timestamp 1728304996
transform 1 0 11250 0 -1 3130
box -12 -8 92 252
use NOR2X1  _1846_
timestamp 1728305106
transform 1 0 11250 0 -1 3610
box -12 -8 92 252
use NAND2X1  _1847_
timestamp 1728304996
transform -1 0 8250 0 1 4090
box -12 -8 92 252
use NOR2X1  _1848_
timestamp 1728305106
transform 1 0 10790 0 -1 2650
box -12 -8 92 252
use NAND2X1  _1849_
timestamp 1728304996
transform -1 0 10750 0 1 2650
box -12 -8 92 252
use OAI21X1  _1850_
timestamp 1728305162
transform -1 0 8730 0 1 4090
box -12 -8 112 252
use NAND2X1  _1851_
timestamp 1728304996
transform -1 0 11330 0 -1 2650
box -12 -8 92 252
use NOR2X1  _1852_
timestamp 1728305106
transform 1 0 9810 0 -1 250
box -12 -8 92 252
use NAND2X1  _1853_
timestamp 1728304996
transform 1 0 9350 0 -1 5050
box -12 -8 92 252
use OAI21X1  _1854_
timestamp 1728305162
transform 1 0 9130 0 1 5050
box -12 -8 112 252
use NOR2X1  _1855_
timestamp 1728305106
transform 1 0 8910 0 1 5050
box -12 -8 92 252
use INVX1  _1856_
timestamp 1728304789
transform 1 0 9430 0 -1 3130
box -12 -8 72 252
use NOR2X1  _1857_
timestamp 1728305106
transform 1 0 9190 0 -1 3130
box -12 -8 92 252
use NOR2X1  _1858_
timestamp 1728305106
transform 1 0 7390 0 -1 5050
box -12 -8 92 252
use NAND2X1  _1859_
timestamp 1728304996
transform -1 0 10870 0 1 1690
box -12 -8 92 252
use OAI21X1  _1860_
timestamp 1728305162
transform 1 0 7170 0 1 5050
box -12 -8 112 252
use INVX1  _1861_
timestamp 1728304789
transform 1 0 7430 0 1 5050
box -12 -8 72 252
use NAND2X1  _1862_
timestamp 1728304996
transform -1 0 9970 0 -1 4570
box -12 -8 92 252
use NOR2X1  _1863_
timestamp 1728305106
transform 1 0 8670 0 -1 2650
box -12 -8 92 252
use NAND2X1  _1864_
timestamp 1728304996
transform 1 0 9970 0 1 2170
box -12 -8 92 252
use NOR2X1  _1865_
timestamp 1728305106
transform 1 0 7810 0 1 2170
box -12 -8 92 252
use NOR2X1  _1866_
timestamp 1728305106
transform -1 0 9070 0 -1 4090
box -12 -8 92 252
use INVX1  _1867_
timestamp 1728304789
transform 1 0 9390 0 1 5050
box -12 -8 72 252
use NOR2X1  _1868_
timestamp 1728305106
transform 1 0 10930 0 -1 250
box -12 -8 92 252
use OAI21X1  _1869_
timestamp 1728305162
transform 1 0 9410 0 -1 4570
box -12 -8 112 252
use NAND3X1  _1870_
timestamp 1728305047
transform -1 0 9250 0 -1 4570
box -12 -8 112 252
use NAND2X1  _1871_
timestamp 1728304996
transform 1 0 8630 0 1 4570
box -12 -8 92 252
use OAI21X1  _1872_
timestamp 1728305162
transform 1 0 7910 0 1 4090
box -12 -8 112 252
use INVX1  _1873_
timestamp 1728304789
transform 1 0 6450 0 1 3130
box -12 -8 72 252
use OAI21X1  _1874_
timestamp 1728305162
transform -1 0 7010 0 1 3130
box -12 -8 112 252
use OR2X2  _1875_
timestamp 1728305284
transform -1 0 6750 0 1 3130
box -12 -8 112 252
use INVX1  _1876_
timestamp 1728304789
transform 1 0 6750 0 1 4090
box -12 -8 72 252
use NAND3X1  _1877_
timestamp 1728305047
transform -1 0 8250 0 1 4570
box -12 -8 112 252
use NOR2X1  _1878_
timestamp 1728305106
transform -1 0 8470 0 1 4570
box -12 -8 92 252
use NAND3X1  _1879_
timestamp 1728305047
transform -1 0 8250 0 1 5050
box -12 -8 112 252
use OAI22X1  _1880_
timestamp 1728305200
transform -1 0 7210 0 -1 8890
box -12 -8 132 252
use INVX1  _1881_
timestamp 1728304789
transform -1 0 6450 0 -1 8890
box -12 -8 72 252
use INVX2  _1882_
timestamp 1728304826
transform 1 0 3590 0 1 7450
box -12 -8 72 252
use OAI22X1  _1883_
timestamp 1728305200
transform -1 0 7210 0 1 8410
box -12 -8 132 252
use INVX2  _1884_
timestamp 1728304826
transform -1 0 6690 0 1 8890
box -12 -8 72 252
use INVX1  _1885_
timestamp 1728304789
transform 1 0 5930 0 1 5530
box -12 -8 72 252
use OAI22X1  _1886_
timestamp 1728305200
transform -1 0 6410 0 -1 8410
box -12 -8 132 252
use INVX2  _1887_
timestamp 1728304826
transform 1 0 6950 0 1 9370
box -12 -8 72 252
use INVX2  _1888_
timestamp 1728304826
transform 1 0 3710 0 1 7930
box -12 -8 72 252
use OAI22X1  _1889_
timestamp 1728305200
transform -1 0 6150 0 -1 8410
box -12 -8 132 252
use INVX1  _1890_
timestamp 1728304789
transform 1 0 6530 0 -1 9850
box -12 -8 72 252
use OAI22X1  _1891_
timestamp 1728305200
transform -1 0 6250 0 -1 8890
box -12 -8 132 252
use INVX2  _1892_
timestamp 1728304826
transform 1 0 5730 0 -1 10330
box -12 -8 72 252
use INVX2  _1893_
timestamp 1728304826
transform 1 0 1130 0 -1 8890
box -12 -8 72 252
use OAI22X1  _1894_
timestamp 1728305200
transform 1 0 6050 0 1 8410
box -12 -8 132 252
use INVX2  _1895_
timestamp 1728304826
transform 1 0 6950 0 1 10810
box -12 -8 72 252
use INVX2  _1896_
timestamp 1728304826
transform 1 0 5250 0 1 6010
box -12 -8 72 252
use OAI22X1  _1897_
timestamp 1728305200
transform 1 0 6110 0 -1 7930
box -12 -8 132 252
use INVX2  _1898_
timestamp 1728304826
transform 1 0 6530 0 1 10330
box -12 -8 72 252
use OAI22X1  _1899_
timestamp 1728305200
transform 1 0 6610 0 -1 7930
box -12 -8 132 252
use INVX1  _1900_
timestamp 1728304789
transform 1 0 650 0 1 2170
box -12 -8 72 252
use NAND2X1  _1901_
timestamp 1728304996
transform 1 0 8090 0 1 5530
box -12 -8 92 252
use OAI21X1  _1902_
timestamp 1728305162
transform 1 0 8610 0 -1 5050
box -12 -8 112 252
use NOR2X1  _1903_
timestamp 1728305106
transform 1 0 7990 0 -1 3130
box -12 -8 92 252
use NOR2X1  _1904_
timestamp 1728305106
transform -1 0 10190 0 1 3610
box -12 -8 92 252
use NOR2X1  _1905_
timestamp 1728305106
transform 1 0 7650 0 1 4570
box -12 -8 92 252
use NAND3X1  _1906_
timestamp 1728305047
transform 1 0 7630 0 -1 5050
box -12 -8 112 252
use NAND2X1  _1907_
timestamp 1728304996
transform 1 0 8750 0 -1 4090
box -12 -8 92 252
use NAND3X1  _1908_
timestamp 1728305047
transform -1 0 7910 0 -1 4090
box -12 -8 112 252
use NOR2X1  _1909_
timestamp 1728305106
transform 1 0 1930 0 -1 4090
box -12 -8 92 252
use NAND3X1  _1910_
timestamp 1728305047
transform -1 0 9950 0 -1 2650
box -12 -8 112 252
use NAND2X1  _1911_
timestamp 1728304996
transform 1 0 9610 0 1 3130
box -12 -8 92 252
use OAI21X1  _1912_
timestamp 1728305162
transform 1 0 6210 0 1 3130
box -12 -8 112 252
use NOR2X1  _1913_
timestamp 1728305106
transform 1 0 10750 0 1 4570
box -12 -8 92 252
use NOR2X1  _1914_
timestamp 1728305106
transform 1 0 10810 0 -1 3610
box -12 -8 92 252
use NAND2X1  _1915_
timestamp 1728304996
transform -1 0 10410 0 1 3610
box -12 -8 92 252
use OAI21X1  _1916_
timestamp 1728305162
transform -1 0 6070 0 1 3130
box -12 -8 112 252
use NOR2X1  _1917_
timestamp 1728305106
transform 1 0 4130 0 1 3130
box -12 -8 92 252
use AND2X2  _1918_
timestamp 1728304163
transform -1 0 970 0 -1 3130
box -12 -8 112 252
use NAND2X1  _1919_
timestamp 1728304996
transform -1 0 250 0 -1 3130
box -12 -8 92 252
use INVX1  _1920_
timestamp 1728304789
transform 1 0 1110 0 1 2650
box -12 -8 72 252
use INVX1  _1921_
timestamp 1728304789
transform -1 0 1350 0 1 3130
box -12 -8 72 252
use AOI21X1  _1922_
timestamp 1728304211
transform -1 0 1130 0 1 3130
box -12 -8 112 252
use OAI21X1  _1923_
timestamp 1728305162
transform 1 0 630 0 -1 3130
box -12 -8 112 252
use OAI21X1  _1924_
timestamp 1728305162
transform -1 0 4670 0 1 3130
box -12 -8 112 252
use INVX1  _1925_
timestamp 1728304789
transform -1 0 450 0 -1 1690
box -12 -8 72 252
use NOR2X1  _1926_
timestamp 1728305106
transform 1 0 890 0 1 2650
box -12 -8 92 252
use NOR3X1  _1927_
timestamp 1728303224
transform -1 0 2350 0 -1 4090
box -12 -8 192 252
use AND2X2  _1928_
timestamp 1728304163
transform -1 0 1770 0 -1 3610
box -12 -8 112 252
use NAND3X1  _1929_
timestamp 1728305047
transform 1 0 390 0 1 2650
box -12 -8 112 252
use AOI21X1  _1930_
timestamp 1728304211
transform 1 0 770 0 1 3130
box -12 -8 112 252
use NAND3X1  _1931_
timestamp 1728305047
transform 1 0 630 0 1 2650
box -12 -8 112 252
use AOI22X1  _1932_
timestamp 1728304278
transform -1 0 770 0 -1 3610
box -14 -8 132 252
use AOI22X1  _1933_
timestamp 1728304278
transform 1 0 630 0 -1 5050
box -14 -8 132 252
use AND2X2  _1934_
timestamp 1728304163
transform -1 0 750 0 1 3610
box -12 -8 112 252
use NAND3X1  _1935_
timestamp 1728305047
transform -1 0 1730 0 1 3610
box -12 -8 112 252
use OAI21X1  _1936_
timestamp 1728305162
transform 1 0 890 0 1 3610
box -12 -8 112 252
use NAND3X1  _1937_
timestamp 1728305047
transform -1 0 750 0 1 4570
box -12 -8 112 252
use INVX1  _1938_
timestamp 1728304789
transform -1 0 230 0 -1 2650
box -12 -8 72 252
use NAND3X1  _1939_
timestamp 1728305047
transform 1 0 390 0 -1 3130
box -12 -8 112 252
use AOI22X1  _1940_
timestamp 1728304278
transform 1 0 930 0 -1 3610
box -14 -8 132 252
use NAND2X1  _1941_
timestamp 1728304996
transform 1 0 630 0 1 5530
box -12 -8 92 252
use NAND3X1  _1942_
timestamp 1728305047
transform 1 0 650 0 -1 5530
box -12 -8 112 252
use INVX1  _1943_
timestamp 1728304789
transform 1 0 8210 0 1 6490
box -12 -8 72 252
use AOI21X1  _1944_
timestamp 1728304211
transform -1 0 7810 0 1 3610
box -12 -8 112 252
use INVX1  _1945_
timestamp 1728304789
transform -1 0 7570 0 1 3610
box -12 -8 72 252
use NOR2X1  _1946_
timestamp 1728305106
transform 1 0 8530 0 -1 4090
box -12 -8 92 252
use NOR2X1  _1947_
timestamp 1728305106
transform -1 0 7790 0 -1 3610
box -12 -8 92 252
use NAND2X1  _1948_
timestamp 1728304996
transform -1 0 7130 0 1 3610
box -12 -8 92 252
use NOR2X1  _1949_
timestamp 1728305106
transform -1 0 7350 0 1 3610
box -12 -8 92 252
use OAI21X1  _1950_
timestamp 1728305162
transform 1 0 8410 0 1 5050
box -12 -8 112 252
use INVX1  _1951_
timestamp 1728304789
transform 1 0 8410 0 1 4090
box -12 -8 72 252
use INVX2  _1952_
timestamp 1728304826
transform 1 0 9910 0 1 3610
box -12 -8 72 252
use OAI21X1  _1953_
timestamp 1728305162
transform -1 0 8570 0 1 3610
box -12 -8 112 252
use NOR2X1  _1954_
timestamp 1728305106
transform 1 0 8310 0 -1 4090
box -12 -8 92 252
use NOR2X1  _1955_
timestamp 1728305106
transform 1 0 6530 0 -1 3610
box -12 -8 92 252
use NAND3X1  _1956_
timestamp 1728305047
transform -1 0 8170 0 -1 4090
box -12 -8 112 252
use INVX2  _1957_
timestamp 1728304826
transform 1 0 8150 0 -1 5530
box -12 -8 72 252
use NAND2X1  _1958_
timestamp 1728304996
transform 1 0 10530 0 -1 2170
box -12 -8 92 252
use OAI21X1  _1959_
timestamp 1728305162
transform 1 0 7890 0 1 4570
box -12 -8 112 252
use INVX1  _1960_
timestamp 1728304789
transform 1 0 7950 0 -1 4570
box -12 -8 72 252
use NOR2X1  _1961_
timestamp 1728305106
transform 1 0 10790 0 -1 3130
box -12 -8 92 252
use NAND2X1  _1962_
timestamp 1728304996
transform 1 0 10570 0 1 3130
box -12 -8 92 252
use OAI21X1  _1963_
timestamp 1728305162
transform 1 0 9930 0 -1 4090
box -12 -8 112 252
use NOR2X1  _1964_
timestamp 1728305106
transform -1 0 7530 0 1 4090
box -12 -8 92 252
use NAND3X1  _1965_
timestamp 1728305047
transform -1 0 7810 0 -1 4570
box -12 -8 112 252
use NAND2X1  _1966_
timestamp 1728304996
transform -1 0 3670 0 -1 8890
box -12 -8 92 252
use OAI21X1  _1967_
timestamp 1728305162
transform -1 0 7150 0 1 7930
box -12 -8 112 252
use AOI21X1  _1968_
timestamp 1728304211
transform 1 0 7590 0 -1 7930
box -12 -8 112 252
use OAI21X1  _1969_
timestamp 1728305162
transform -1 0 7950 0 -1 7930
box -12 -8 112 252
use NAND2X1  _1970_
timestamp 1728304996
transform 1 0 1590 0 1 4090
box -12 -8 92 252
use AOI22X1  _1971_
timestamp 1728304278
transform -1 0 1010 0 -1 4090
box -14 -8 132 252
use NAND3X1  _1972_
timestamp 1728305047
transform 1 0 1430 0 -1 4090
box -12 -8 112 252
use NAND3X1  _1973_
timestamp 1728305047
transform 1 0 1670 0 -1 4090
box -12 -8 112 252
use INVX1  _1974_
timestamp 1728304789
transform 1 0 8450 0 -1 6970
box -12 -8 72 252
use INVX1  _1975_
timestamp 1728304789
transform 1 0 3050 0 -1 9850
box -12 -8 72 252
use NAND2X1  _1976_
timestamp 1728304996
transform -1 0 7290 0 1 4090
box -12 -8 92 252
use NOR2X1  _1977_
timestamp 1728305106
transform -1 0 2990 0 1 9370
box -12 -8 92 252
use INVX1  _1978_
timestamp 1728304789
transform -1 0 3930 0 1 9370
box -12 -8 72 252
use OAI21X1  _1979_
timestamp 1728305162
transform -1 0 6690 0 1 8410
box -12 -8 112 252
use AOI21X1  _1980_
timestamp 1728304211
transform 1 0 7870 0 1 8410
box -12 -8 112 252
use OAI21X1  _1981_
timestamp 1728305162
transform 1 0 8370 0 1 8410
box -12 -8 112 252
use NAND2X1  _1982_
timestamp 1728304996
transform -1 0 3190 0 1 6010
box -12 -8 92 252
use AOI22X1  _1983_
timestamp 1728304278
transform 1 0 1790 0 1 5530
box -14 -8 132 252
use NAND3X1  _1984_
timestamp 1728305047
transform 1 0 1890 0 -1 5530
box -12 -8 112 252
use NAND3X1  _1985_
timestamp 1728305047
transform 1 0 2550 0 1 5530
box -12 -8 112 252
use INVX1  _1986_
timestamp 1728304789
transform -1 0 7250 0 -1 6970
box -12 -8 72 252
use INVX1  _1987_
timestamp 1728304789
transform 1 0 5170 0 1 9850
box -12 -8 72 252
use OAI22X1  _1988_
timestamp 1728305200
transform -1 0 5170 0 -1 8410
box -12 -8 132 252
use AOI21X1  _1989_
timestamp 1728304211
transform 1 0 6810 0 -1 8410
box -12 -8 112 252
use OAI21X1  _1990_
timestamp 1728305162
transform -1 0 7430 0 -1 8410
box -12 -8 112 252
use NAND2X1  _1991_
timestamp 1728304996
transform -1 0 2190 0 -1 5050
box -12 -8 92 252
use AOI22X1  _1992_
timestamp 1728304278
transform -1 0 1750 0 1 5050
box -14 -8 132 252
use NAND3X1  _1993_
timestamp 1728305047
transform -1 0 2010 0 1 5050
box -12 -8 112 252
use NAND3X1  _1994_
timestamp 1728305047
transform 1 0 2150 0 1 5050
box -12 -8 112 252
use INVX1  _1995_
timestamp 1728304789
transform 1 0 8130 0 1 6970
box -12 -8 72 252
use NAND2X1  _1996_
timestamp 1728304996
transform -1 0 2410 0 1 8890
box -12 -8 92 252
use OAI21X1  _1997_
timestamp 1728305162
transform -1 0 4130 0 -1 8410
box -12 -8 112 252
use AOI21X1  _1998_
timestamp 1728304211
transform -1 0 6670 0 -1 8410
box -12 -8 112 252
use OAI21X1  _1999_
timestamp 1728305162
transform -1 0 8370 0 1 7930
box -12 -8 112 252
use NAND2X1  _2000_
timestamp 1728304996
transform 1 0 1910 0 -1 6970
box -12 -8 92 252
use AOI22X1  _2001_
timestamp 1728304278
transform 1 0 1390 0 1 6490
box -14 -8 132 252
use NAND3X1  _2002_
timestamp 1728305047
transform 1 0 1610 0 1 7450
box -12 -8 112 252
use NAND3X1  _2003_
timestamp 1728305047
transform 1 0 1650 0 -1 6970
box -12 -8 112 252
use INVX1  _2004_
timestamp 1728304789
transform 1 0 7910 0 1 6970
box -12 -8 72 252
use NAND2X1  _2005_
timestamp 1728304996
transform 1 0 2090 0 -1 9370
box -12 -8 92 252
use OAI21X1  _2006_
timestamp 1728305162
transform -1 0 6430 0 1 8410
box -12 -8 112 252
use AOI21X1  _2007_
timestamp 1728304211
transform 1 0 7610 0 1 8410
box -12 -8 112 252
use OAI21X1  _2008_
timestamp 1728305162
transform -1 0 8230 0 1 8410
box -12 -8 112 252
use NAND2X1  _2009_
timestamp 1728304996
transform 1 0 890 0 -1 7450
box -12 -8 92 252
use AOI22X1  _2010_
timestamp 1728304278
transform -1 0 1030 0 -1 6490
box -14 -8 132 252
use NAND3X1  _2011_
timestamp 1728305047
transform 1 0 650 0 1 7450
box -12 -8 112 252
use NAND3X1  _2012_
timestamp 1728305047
transform 1 0 890 0 1 7450
box -12 -8 112 252
use INVX1  _2013_
timestamp 1728304789
transform 1 0 5550 0 1 7930
box -12 -8 72 252
use NAND2X1  _2014_
timestamp 1728304996
transform 1 0 1850 0 1 8890
box -12 -8 92 252
use OAI21X1  _2015_
timestamp 1728305162
transform -1 0 4110 0 1 8410
box -12 -8 112 252
use AOI21X1  _2016_
timestamp 1728304211
transform 1 0 6850 0 1 8410
box -12 -8 112 252
use OAI21X1  _2017_
timestamp 1728305162
transform -1 0 7470 0 1 8410
box -12 -8 112 252
use NAND2X1  _2018_
timestamp 1728304996
transform -1 0 1670 0 -1 7450
box -12 -8 92 252
use AOI22X1  _2019_
timestamp 1728304278
transform -1 0 1790 0 1 6490
box -14 -8 132 252
use NAND3X1  _2020_
timestamp 1728305047
transform 1 0 1850 0 1 6970
box -12 -8 112 252
use NAND3X1  _2021_
timestamp 1728305047
transform 1 0 1830 0 -1 7450
box -12 -8 112 252
use INVX1  _2022_
timestamp 1728304789
transform 1 0 4610 0 1 7930
box -12 -8 72 252
use INVX1  _2023_
timestamp 1728304789
transform 1 0 630 0 -1 8410
box -12 -8 72 252
use NOR2X1  _2024_
timestamp 1728305106
transform 1 0 1550 0 -1 8410
box -12 -8 92 252
use INVX1  _2025_
timestamp 1728304789
transform 1 0 2590 0 1 8410
box -12 -8 72 252
use OAI21X1  _2026_
timestamp 1728305162
transform -1 0 4890 0 1 8410
box -12 -8 112 252
use AOI21X1  _2027_
timestamp 1728304211
transform 1 0 7310 0 1 7930
box -12 -8 112 252
use OAI21X1  _2028_
timestamp 1728305162
transform -1 0 7650 0 1 7930
box -12 -8 112 252
use NAND2X1  _2029_
timestamp 1728304996
transform -1 0 250 0 -1 6970
box -12 -8 92 252
use AOI22X1  _2030_
timestamp 1728304278
transform -1 0 770 0 -1 6490
box -14 -8 132 252
use NAND3X1  _2031_
timestamp 1728305047
transform -1 0 490 0 -1 6970
box -12 -8 112 252
use NAND3X1  _2032_
timestamp 1728305047
transform 1 0 650 0 1 6490
box -12 -8 112 252
use INVX1  _2033_
timestamp 1728304789
transform 1 0 7710 0 1 6970
box -12 -8 72 252
use INVX1  _2034_
timestamp 1728304789
transform 1 0 1330 0 -1 8410
box -12 -8 72 252
use NOR2X1  _2035_
timestamp 1728305106
transform 1 0 2210 0 1 7930
box -12 -8 92 252
use INVX1  _2036_
timestamp 1728304789
transform 1 0 2990 0 -1 7930
box -12 -8 72 252
use OAI21X1  _2037_
timestamp 1728305162
transform -1 0 4290 0 -1 7930
box -12 -8 112 252
use AOI21X1  _2038_
timestamp 1728304211
transform 1 0 7650 0 1 7450
box -12 -8 112 252
use OAI21X1  _2039_
timestamp 1728305162
transform -1 0 7990 0 1 7450
box -12 -8 112 252
use NAND2X1  _2040_
timestamp 1728304996
transform -1 0 3110 0 1 2650
box -12 -8 92 252
use INVX8  _2041_
timestamp 1728304916
transform -1 0 750 0 1 1690
box -12 -8 133 252
use INVX1  _2042_
timestamp 1728304789
transform 1 0 1830 0 1 4090
box -12 -8 72 252
use INVX1  _2043_
timestamp 1728304789
transform -1 0 3970 0 -1 11290
box -12 -8 72 252
use INVX1  _2044_
timestamp 1728304789
transform 1 0 5450 0 1 6010
box -12 -8 72 252
use OAI21X1  _2045_
timestamp 1728305162
transform -1 0 4250 0 -1 7450
box -12 -8 112 252
use AOI21X1  _2046_
timestamp 1728304211
transform 1 0 2970 0 -1 4090
box -12 -8 112 252
use OAI21X1  _2047_
timestamp 1728305162
transform 1 0 2710 0 -1 4090
box -12 -8 112 252
use INVX1  _2048_
timestamp 1728304789
transform -1 0 3710 0 -1 4570
box -12 -8 72 252
use AOI21X1  _2049_
timestamp 1728304211
transform -1 0 3130 0 -1 4570
box -12 -8 112 252
use OAI21X1  _2050_
timestamp 1728305162
transform -1 0 2630 0 1 4090
box -12 -8 112 252
use NAND2X1  _2051_
timestamp 1728304996
transform -1 0 2590 0 1 250
box -12 -8 92 252
use INVX1  _2052_
timestamp 1728304789
transform -1 0 970 0 1 250
box -12 -8 72 252
use INVX1  _2053_
timestamp 1728304789
transform -1 0 3550 0 1 4090
box -12 -8 72 252
use AOI21X1  _2054_
timestamp 1728304211
transform 1 0 3210 0 -1 4090
box -12 -8 112 252
use OAI21X1  _2055_
timestamp 1728305162
transform -1 0 2950 0 1 3610
box -12 -8 112 252
use INVX1  _2056_
timestamp 1728304789
transform 1 0 4490 0 1 6970
box -12 -8 72 252
use NAND2X1  _2057_
timestamp 1728304996
transform -1 0 4090 0 1 7450
box -12 -8 92 252
use OAI21X1  _2058_
timestamp 1728305162
transform 1 0 4710 0 1 6970
box -12 -8 112 252
use INVX2  _2059_
timestamp 1728304826
transform -1 0 2110 0 1 4090
box -12 -8 72 252
use INVX1  _2060_
timestamp 1728304789
transform -1 0 3910 0 -1 5050
box -12 -8 72 252
use NAND2X1  _2061_
timestamp 1728304996
transform 1 0 3630 0 1 5050
box -12 -8 92 252
use OAI21X1  _2062_
timestamp 1728305162
transform -1 0 3710 0 -1 5050
box -12 -8 112 252
use NAND2X1  _2063_
timestamp 1728304996
transform 1 0 2590 0 1 3130
box -12 -8 92 252
use NAND2X1  _2064_
timestamp 1728304996
transform -1 0 2750 0 -1 250
box -12 -8 92 252
use INVX1  _2065_
timestamp 1728304789
transform -1 0 2510 0 -1 250
box -12 -8 72 252
use NAND2X1  _2066_
timestamp 1728304996
transform 1 0 2550 0 -1 730
box -12 -8 92 252
use NAND2X1  _2067_
timestamp 1728304996
transform -1 0 2930 0 1 4570
box -12 -8 92 252
use OAI21X1  _2068_
timestamp 1728305162
transform -1 0 3170 0 1 4570
box -12 -8 112 252
use NAND2X1  _2069_
timestamp 1728304996
transform 1 0 2650 0 -1 3610
box -12 -8 92 252
use INVX2  _2070_
timestamp 1728304826
transform -1 0 1210 0 -1 730
box -12 -8 72 252
use OAI21X1  _2071_
timestamp 1728305162
transform -1 0 2990 0 -1 5530
box -12 -8 112 252
use AOI21X1  _2072_
timestamp 1728304211
transform -1 0 2730 0 -1 5530
box -12 -8 112 252
use NOR2X1  _2073_
timestamp 1728305106
transform -1 0 1430 0 -1 1210
box -12 -8 92 252
use NAND2X1  _2074_
timestamp 1728304996
transform 1 0 3330 0 1 4570
box -12 -8 92 252
use OAI21X1  _2075_
timestamp 1728305162
transform -1 0 2890 0 -1 4570
box -12 -8 112 252
use NAND2X1  _2076_
timestamp 1728304996
transform 1 0 2490 0 -1 4090
box -12 -8 92 252
use MUX2X1  _2077_
timestamp 1728304958
transform -1 0 3470 0 1 5050
box -12 -8 131 252
use NOR2X1  _2078_
timestamp 1728305106
transform 1 0 2870 0 -1 3610
box -12 -8 92 252
use NAND2X1  _2079_
timestamp 1728304996
transform -1 0 4070 0 -1 1210
box -12 -8 92 252
use INVX1  _2080_
timestamp 1728304789
transform 1 0 4230 0 -1 1210
box -12 -8 72 252
use NAND2X1  _2081_
timestamp 1728304996
transform -1 0 3830 0 -1 1210
box -12 -8 92 252
use NOR2X1  _2082_
timestamp 1728305106
transform 1 0 5870 0 -1 1210
box -12 -8 92 252
use AOI22X1  _2083_
timestamp 1728304278
transform -1 0 6690 0 -1 1210
box -14 -8 132 252
use NOR2X1  _2084_
timestamp 1728305106
transform 1 0 10030 0 -1 1690
box -12 -8 92 252
use OAI21X1  _2085_
timestamp 1728305162
transform -1 0 10630 0 -1 1690
box -12 -8 112 252
use NAND2X1  _2086_
timestamp 1728304996
transform 1 0 10550 0 1 1690
box -12 -8 92 252
use NOR2X1  _2087_
timestamp 1728305106
transform 1 0 11110 0 -1 4570
box -12 -8 92 252
use OAI21X1  _2088_
timestamp 1728305162
transform 1 0 10310 0 1 1690
box -12 -8 112 252
use NAND2X1  _2089_
timestamp 1728304996
transform -1 0 9650 0 1 730
box -12 -8 92 252
use NOR2X1  _2090_
timestamp 1728305106
transform 1 0 10790 0 -1 5050
box -12 -8 92 252
use INVX1  _2091_
timestamp 1728304789
transform 1 0 11270 0 -1 5050
box -12 -8 72 252
use NOR2X1  _2092_
timestamp 1728305106
transform -1 0 10310 0 1 2650
box -12 -8 92 252
use NAND2X1  _2093_
timestamp 1728304996
transform 1 0 10310 0 -1 3610
box -12 -8 92 252
use OAI21X1  _2094_
timestamp 1728305162
transform -1 0 10870 0 1 4090
box -12 -8 112 252
use NOR2X1  _2095_
timestamp 1728305106
transform 1 0 10870 0 -1 4570
box -12 -8 92 252
use OAI21X1  _2096_
timestamp 1728305162
transform -1 0 11350 0 1 4570
box -12 -8 112 252
use INVX1  _2097_
timestamp 1728304789
transform -1 0 11230 0 -1 1210
box -12 -8 72 252
use INVX1  _2098_
timestamp 1728304789
transform 1 0 10290 0 -1 730
box -12 -8 72 252
use NAND2X1  _2099_
timestamp 1728304996
transform 1 0 10750 0 -1 730
box -12 -8 92 252
use NOR2X1  _2100_
timestamp 1728305106
transform 1 0 10990 0 -1 730
box -12 -8 92 252
use INVX1  _2101_
timestamp 1728304789
transform 1 0 11230 0 -1 730
box -12 -8 72 252
use OAI21X1  _2102_
timestamp 1728305162
transform 1 0 4090 0 -1 4570
box -12 -8 112 252
use AOI21X1  _2103_
timestamp 1728304211
transform 1 0 4350 0 -1 4570
box -12 -8 112 252
use NAND2X1  _2104_
timestamp 1728304996
transform 1 0 3950 0 1 250
box -12 -8 92 252
use INVX1  _2105_
timestamp 1728304789
transform -1 0 1910 0 1 250
box -12 -8 72 252
use NAND2X1  _2106_
timestamp 1728304996
transform -1 0 2310 0 -1 250
box -12 -8 92 252
use NAND2X1  _2107_
timestamp 1728304996
transform -1 0 2810 0 1 250
box -12 -8 92 252
use INVX2  _2108_
timestamp 1728304826
transform 1 0 1570 0 1 1690
box -12 -8 72 252
use NAND2X1  _2109_
timestamp 1728304996
transform -1 0 3050 0 1 250
box -12 -8 92 252
use OAI22X1  _2110_
timestamp 1728305200
transform 1 0 3190 0 1 250
box -12 -8 132 252
use NAND3X1  _2111_
timestamp 1728305047
transform 1 0 5410 0 1 250
box -12 -8 112 252
use NOR2X1  _2112_
timestamp 1728305106
transform 1 0 11270 0 1 3130
box -12 -8 92 252
use NAND2X1  _2113_
timestamp 1728304996
transform -1 0 9930 0 1 3130
box -12 -8 92 252
use OAI21X1  _2114_
timestamp 1728305162
transform 1 0 9870 0 -1 3130
box -12 -8 112 252
use INVX1  _2115_
timestamp 1728304789
transform -1 0 11210 0 -1 250
box -12 -8 72 252
use INVX1  _2116_
timestamp 1728304789
transform -1 0 11170 0 1 5050
box -12 -8 72 252
use NAND2X1  _2117_
timestamp 1728304996
transform -1 0 10790 0 1 5530
box -12 -8 92 252
use NAND2X1  _2118_
timestamp 1728304996
transform 1 0 9110 0 -1 5050
box -12 -8 92 252
use NAND3X1  _2119_
timestamp 1728305047
transform -1 0 11290 0 1 5530
box -12 -8 112 252
use NOR2X1  _2120_
timestamp 1728305106
transform 1 0 11130 0 1 2650
box -12 -8 92 252
use INVX1  _2121_
timestamp 1728304789
transform 1 0 11250 0 1 730
box -12 -8 72 252
use NOR2X1  _2122_
timestamp 1728305106
transform 1 0 10950 0 -1 1210
box -12 -8 92 252
use NAND2X1  _2123_
timestamp 1728304996
transform 1 0 10990 0 -1 1690
box -12 -8 92 252
use NOR2X1  _2124_
timestamp 1728305106
transform 1 0 9470 0 1 2170
box -12 -8 92 252
use INVX1  _2125_
timestamp 1728304789
transform 1 0 9590 0 1 1690
box -12 -8 72 252
use NOR2X1  _2126_
timestamp 1728305106
transform -1 0 10070 0 1 2650
box -12 -8 92 252
use NAND2X1  _2127_
timestamp 1728304996
transform 1 0 9850 0 -1 2170
box -12 -8 92 252
use OAI21X1  _2128_
timestamp 1728305162
transform 1 0 9790 0 1 1690
box -12 -8 112 252
use NAND2X1  _2129_
timestamp 1728304996
transform -1 0 9090 0 1 2170
box -12 -8 92 252
use OAI21X1  _2130_
timestamp 1728305162
transform 1 0 9710 0 1 2170
box -12 -8 112 252
use NOR2X1  _2131_
timestamp 1728305106
transform 1 0 9790 0 -1 1690
box -12 -8 92 252
use OR2X2  _2132_
timestamp 1728305284
transform 1 0 10270 0 -1 1690
box -12 -8 112 252
use NOR2X1  _2133_
timestamp 1728305106
transform 1 0 10410 0 1 1210
box -12 -8 92 252
use NOR2X1  _2134_
timestamp 1728305106
transform -1 0 10270 0 1 1210
box -12 -8 92 252
use NOR2X1  _2135_
timestamp 1728305106
transform 1 0 10710 0 -1 1210
box -12 -8 92 252
use AOI22X1  _2136_
timestamp 1728304278
transform -1 0 10750 0 1 1210
box -14 -8 132 252
use NAND3X1  _2137_
timestamp 1728305047
transform 1 0 10910 0 1 1210
box -12 -8 112 252
use AOI21X1  _2138_
timestamp 1728304211
transform -1 0 11090 0 1 730
box -12 -8 112 252
use NAND3X1  _2139_
timestamp 1728305047
transform -1 0 11010 0 1 250
box -12 -8 112 252
use OR2X2  _2140_
timestamp 1728305284
transform -1 0 8510 0 -1 250
box -12 -8 112 252
use INVX1  _2141_
timestamp 1728304789
transform 1 0 8650 0 -1 250
box -12 -8 72 252
use NOR2X1  _2142_
timestamp 1728305106
transform 1 0 1990 0 -1 250
box -12 -8 92 252
use NAND3X1  _2143_
timestamp 1728305047
transform -1 0 3110 0 -1 730
box -12 -8 112 252
use INVX1  _2144_
timestamp 1728304789
transform -1 0 6150 0 -1 1210
box -12 -8 72 252
use AOI22X1  _2145_
timestamp 1728304278
transform -1 0 6430 0 -1 1210
box -14 -8 132 252
use NOR2X1  _2146_
timestamp 1728305106
transform 1 0 5630 0 -1 1210
box -12 -8 92 252
use AOI22X1  _2147_
timestamp 1728304278
transform -1 0 6950 0 -1 1210
box -14 -8 132 252
use NOR2X1  _2148_
timestamp 1728305106
transform 1 0 9770 0 1 2650
box -12 -8 92 252
use OAI21X1  _2149_
timestamp 1728305162
transform 1 0 8830 0 -1 1690
box -12 -8 112 252
use OAI21X1  _2150_
timestamp 1728305162
transform -1 0 8690 0 -1 1690
box -12 -8 112 252
use NOR2X1  _2151_
timestamp 1728305106
transform 1 0 8270 0 1 2170
box -12 -8 92 252
use OAI21X1  _2152_
timestamp 1728305162
transform -1 0 9170 0 -1 1690
box -12 -8 112 252
use OAI21X1  _2153_
timestamp 1728305162
transform -1 0 9290 0 -1 1210
box -12 -8 112 252
use NOR2X1  _2154_
timestamp 1728305106
transform 1 0 8930 0 1 3610
box -12 -8 92 252
use OAI21X1  _2155_
timestamp 1728305162
transform 1 0 8110 0 1 3130
box -12 -8 112 252
use OAI21X1  _2156_
timestamp 1728305162
transform -1 0 8470 0 1 3130
box -12 -8 112 252
use NAND3X1  _2157_
timestamp 1728305047
transform -1 0 8570 0 1 1210
box -12 -8 112 252
use NAND2X1  _2158_
timestamp 1728304996
transform 1 0 10430 0 -1 4090
box -12 -8 92 252
use INVX1  _2159_
timestamp 1728304789
transform 1 0 6130 0 -1 3130
box -12 -8 72 252
use NAND2X1  _2160_
timestamp 1728304996
transform -1 0 6530 0 -1 2650
box -12 -8 92 252
use OAI21X1  _2161_
timestamp 1728305162
transform 1 0 6690 0 -1 2650
box -12 -8 112 252
use OAI21X1  _2162_
timestamp 1728305162
transform -1 0 8090 0 1 2650
box -12 -8 112 252
use INVX2  _2163_
timestamp 1728304826
transform -1 0 8490 0 -1 3610
box -12 -8 72 252
use OAI21X1  _2164_
timestamp 1728305162
transform 1 0 7210 0 -1 2650
box -12 -8 112 252
use AOI21X1  _2165_
timestamp 1728304211
transform -1 0 7250 0 -1 2170
box -12 -8 112 252
use NOR2X1  _2166_
timestamp 1728305106
transform -1 0 8310 0 -1 3130
box -12 -8 92 252
use OAI21X1  _2167_
timestamp 1728305162
transform -1 0 8030 0 -1 2650
box -12 -8 112 252
use OAI21X1  _2168_
timestamp 1728305162
transform -1 0 8270 0 -1 2650
box -12 -8 112 252
use NAND2X1  _2169_
timestamp 1728304996
transform 1 0 8250 0 1 1210
box -12 -8 92 252
use NOR2X1  _2170_
timestamp 1728305106
transform -1 0 8510 0 -1 1210
box -12 -8 92 252
use NAND3X1  _2171_
timestamp 1728305047
transform 1 0 8670 0 -1 1210
box -12 -8 112 252
use OAI21X1  _2172_
timestamp 1728305162
transform -1 0 10610 0 -1 730
box -12 -8 112 252
use OAI21X1  _2173_
timestamp 1728305162
transform 1 0 10250 0 1 730
box -12 -8 112 252
use NOR2X1  _2174_
timestamp 1728305106
transform 1 0 4490 0 -1 1690
box -12 -8 92 252
use NOR2X1  _2175_
timestamp 1728305106
transform -1 0 4110 0 -1 1690
box -12 -8 92 252
use AOI22X1  _2176_
timestamp 1728304278
transform -1 0 5590 0 -1 1690
box -14 -8 132 252
use OAI21X1  _2177_
timestamp 1728305162
transform -1 0 6250 0 -1 2170
box -12 -8 112 252
use OAI21X1  _2178_
timestamp 1728305162
transform -1 0 6490 0 1 1690
box -12 -8 112 252
use NAND2X1  _2179_
timestamp 1728304996
transform 1 0 6470 0 -1 1690
box -12 -8 92 252
use MUX2X1  _2180_
timestamp 1728304958
transform 1 0 7270 0 1 2650
box -12 -8 131 252
use NAND2X1  _2181_
timestamp 1728304996
transform 1 0 7390 0 1 3130
box -12 -8 92 252
use NOR2X1  _2182_
timestamp 1728305106
transform -1 0 7330 0 -1 5530
box -12 -8 92 252
use NAND2X1  _2183_
timestamp 1728304996
transform 1 0 6230 0 -1 2650
box -12 -8 92 252
use OAI21X1  _2184_
timestamp 1728305162
transform 1 0 6570 0 1 2170
box -12 -8 112 252
use NOR2X1  _2185_
timestamp 1728305106
transform -1 0 6770 0 -1 2170
box -12 -8 92 252
use NAND2X1  _2186_
timestamp 1728304996
transform -1 0 9190 0 -1 6970
box -12 -8 92 252
use OR2X2  _2187_
timestamp 1728305284
transform -1 0 9630 0 -1 6490
box -12 -8 112 252
use NAND2X1  _2188_
timestamp 1728304996
transform 1 0 9150 0 1 6490
box -12 -8 92 252
use OAI21X1  _2189_
timestamp 1728305162
transform -1 0 8990 0 1 6490
box -12 -8 112 252
use NOR2X1  _2190_
timestamp 1728305106
transform 1 0 8610 0 -1 6010
box -12 -8 92 252
use OAI21X1  _2191_
timestamp 1728305162
transform 1 0 8830 0 -1 6490
box -12 -8 112 252
use NAND2X1  _2192_
timestamp 1728304996
transform 1 0 7410 0 -1 2170
box -12 -8 92 252
use NOR2X1  _2193_
timestamp 1728305106
transform 1 0 7630 0 -1 1210
box -12 -8 92 252
use NAND2X1  _2194_
timestamp 1728304996
transform -1 0 8790 0 1 3610
box -12 -8 92 252
use INVX1  _2195_
timestamp 1728304789
transform -1 0 8710 0 -1 3610
box -12 -8 72 252
use OAI21X1  _2196_
timestamp 1728305162
transform 1 0 8710 0 -1 3130
box -12 -8 112 252
use OAI21X1  _2197_
timestamp 1728305162
transform 1 0 8730 0 1 2650
box -12 -8 112 252
use OAI21X1  _2198_
timestamp 1728305162
transform -1 0 7430 0 1 2170
box -12 -8 112 252
use OAI21X1  _2199_
timestamp 1728305162
transform -1 0 7670 0 1 2170
box -12 -8 112 252
use INVX1  _2200_
timestamp 1728304789
transform 1 0 9130 0 1 3130
box -12 -8 72 252
use OAI21X1  _2201_
timestamp 1728305162
transform 1 0 8990 0 1 2650
box -12 -8 112 252
use OAI21X1  _2202_
timestamp 1728305162
transform -1 0 8850 0 1 2170
box -12 -8 112 252
use NAND3X1  _2203_
timestamp 1728305047
transform 1 0 8510 0 1 2170
box -12 -8 112 252
use OAI21X1  _2204_
timestamp 1728305162
transform -1 0 8590 0 1 2650
box -12 -8 112 252
use OAI21X1  _2205_
timestamp 1728305162
transform 1 0 8230 0 1 2650
box -12 -8 112 252
use OAI21X1  _2206_
timestamp 1728305162
transform -1 0 8210 0 -1 2170
box -12 -8 112 252
use OAI21X1  _2207_
timestamp 1728305162
transform 1 0 8610 0 -1 2170
box -12 -8 112 252
use AND2X2  _2208_
timestamp 1728304163
transform -1 0 8470 0 -1 2170
box -12 -8 112 252
use INVX1  _2209_
timestamp 1728304789
transform -1 0 7950 0 -1 2170
box -12 -8 72 252
use INVX4  _2210_
timestamp 1728304878
transform 1 0 2830 0 -1 6970
box -12 -8 92 252
use OAI21X1  _2211_
timestamp 1728305162
transform -1 0 7390 0 -1 3130
box -12 -8 112 252
use OAI21X1  _2212_
timestamp 1728305162
transform -1 0 7630 0 -1 3130
box -12 -8 112 252
use NAND3X1  _2213_
timestamp 1728305047
transform -1 0 8170 0 1 1690
box -12 -8 112 252
use NOR2X1  _2214_
timestamp 1728305106
transform 1 0 8650 0 1 730
box -12 -8 92 252
use NAND3X1  _2215_
timestamp 1728305047
transform 1 0 9330 0 1 730
box -12 -8 112 252
use NOR2X1  _2216_
timestamp 1728305106
transform 1 0 9330 0 -1 730
box -12 -8 92 252
use NAND2X1  _2217_
timestamp 1728304996
transform -1 0 9650 0 -1 730
box -12 -8 92 252
use NOR2X1  _2218_
timestamp 1728305106
transform 1 0 4010 0 1 730
box -12 -8 92 252
use AND2X2  _2219_
timestamp 1728304163
transform -1 0 2430 0 1 3130
box -12 -8 112 252
use NAND2X1  _2220_
timestamp 1728304996
transform -1 0 3810 0 -1 730
box -12 -8 92 252
use INVX1  _2221_
timestamp 1728304789
transform 1 0 4210 0 -1 730
box -12 -8 72 252
use NOR2X1  _2222_
timestamp 1728305106
transform 1 0 4430 0 -1 730
box -12 -8 92 252
use OAI21X1  _2223_
timestamp 1728305162
transform 1 0 4230 0 1 730
box -12 -8 112 252
use NOR2X1  _2224_
timestamp 1728305106
transform -1 0 2990 0 -1 250
box -12 -8 92 252
use AOI22X1  _2225_
timestamp 1728304278
transform -1 0 6090 0 1 1210
box -14 -8 132 252
use NOR2X1  _2226_
timestamp 1728305106
transform 1 0 6090 0 1 2650
box -12 -8 92 252
use OAI21X1  _2227_
timestamp 1728305162
transform -1 0 7170 0 1 2170
box -12 -8 112 252
use OAI21X1  _2228_
timestamp 1728305162
transform 1 0 6810 0 1 2170
box -12 -8 112 252
use NAND2X1  _2229_
timestamp 1728304996
transform 1 0 7890 0 -1 5050
box -12 -8 92 252
use NAND2X1  _2230_
timestamp 1728304996
transform -1 0 6350 0 1 4090
box -12 -8 92 252
use OAI21X1  _2231_
timestamp 1728305162
transform -1 0 6590 0 1 4090
box -12 -8 112 252
use AOI21X1  _2232_
timestamp 1728304211
transform 1 0 6950 0 -1 2650
box -12 -8 112 252
use AND2X2  _2233_
timestamp 1728304163
transform 1 0 7510 0 1 1210
box -12 -8 112 252
use NAND3X1  _2234_
timestamp 1728305047
transform 1 0 7430 0 1 730
box -12 -8 112 252
use INVX1  _2235_
timestamp 1728304789
transform 1 0 9510 0 1 250
box -12 -8 72 252
use NAND2X1  _2236_
timestamp 1728304996
transform 1 0 10550 0 -1 3130
box -12 -8 92 252
use OAI21X1  _2237_
timestamp 1728305162
transform 1 0 10050 0 1 1690
box -12 -8 112 252
use NAND3X1  _2238_
timestamp 1728305047
transform -1 0 10050 0 -1 1210
box -12 -8 112 252
use OR2X2  _2239_
timestamp 1728305284
transform -1 0 5990 0 -1 2170
box -12 -8 112 252
use INVX1  _2240_
timestamp 1728304789
transform 1 0 2790 0 -1 730
box -12 -8 72 252
use NAND2X1  _2241_
timestamp 1728304996
transform -1 0 4510 0 -1 1210
box -12 -8 92 252
use NOR2X1  _2242_
timestamp 1728305106
transform -1 0 4750 0 -1 1210
box -12 -8 92 252
use NOR2X1  _2243_
timestamp 1728305106
transform 1 0 3470 0 1 250
box -12 -8 92 252
use NAND3X1  _2244_
timestamp 1728305047
transform 1 0 5210 0 1 730
box -12 -8 112 252
use NAND3X1  _2245_
timestamp 1728305047
transform 1 0 7370 0 -1 1210
box -12 -8 112 252
use INVX1  _2246_
timestamp 1728304789
transform 1 0 7390 0 -1 250
box -12 -8 72 252
use NAND2X1  _2247_
timestamp 1728304996
transform -1 0 3390 0 -1 1690
box -12 -8 92 252
use NOR2X1  _2248_
timestamp 1728305106
transform 1 0 3530 0 1 1210
box -12 -8 92 252
use NAND2X1  _2249_
timestamp 1728304996
transform 1 0 5490 0 1 1210
box -12 -8 92 252
use OAI22X1  _2250_
timestamp 1728305200
transform 1 0 6770 0 1 1210
box -12 -8 132 252
use NAND2X1  _2251_
timestamp 1728304996
transform 1 0 7290 0 1 1210
box -12 -8 92 252
use NOR2X1  _2252_
timestamp 1728305106
transform -1 0 9770 0 -1 4090
box -12 -8 92 252
use NAND2X1  _2253_
timestamp 1728304996
transform 1 0 9450 0 1 1210
box -12 -8 92 252
use NAND2X1  _2254_
timestamp 1728304996
transform 1 0 5730 0 1 1210
box -12 -8 92 252
use NAND3X1  _2255_
timestamp 1728305047
transform -1 0 7130 0 1 1210
box -12 -8 112 252
use NOR2X1  _2256_
timestamp 1728305106
transform 1 0 7230 0 -1 730
box -12 -8 92 252
use NOR2X1  _2257_
timestamp 1728305106
transform -1 0 3210 0 -1 250
box -12 -8 92 252
use OAI21X1  _2258_
timestamp 1728305162
transform -1 0 3210 0 -1 3610
box -12 -8 112 252
use NOR2X1  _2259_
timestamp 1728305106
transform 1 0 3550 0 -1 1690
box -12 -8 92 252
use NAND3X1  _2260_
timestamp 1728305047
transform 1 0 4710 0 1 730
box -12 -8 112 252
use OAI21X1  _2261_
timestamp 1728305162
transform -1 0 5810 0 1 730
box -12 -8 112 252
use NOR2X1  _2262_
timestamp 1728305106
transform 1 0 4890 0 -1 1210
box -12 -8 92 252
use NAND3X1  _2263_
timestamp 1728305047
transform 1 0 4970 0 1 730
box -12 -8 112 252
use OAI21X1  _2264_
timestamp 1728305162
transform -1 0 6350 0 1 730
box -12 -8 112 252
use INVX1  _2265_
timestamp 1728304789
transform 1 0 3550 0 1 3130
box -12 -8 72 252
use INVX1  _2266_
timestamp 1728304789
transform 1 0 7610 0 1 5530
box -12 -8 72 252
use NAND2X1  _2267_
timestamp 1728304996
transform -1 0 5570 0 1 4570
box -12 -8 92 252
use OAI21X1  _2268_
timestamp 1728305162
transform -1 0 5810 0 1 4570
box -12 -8 112 252
use INVX1  _2269_
timestamp 1728304789
transform 1 0 5510 0 -1 5050
box -12 -8 72 252
use NAND2X1  _2270_
timestamp 1728304996
transform -1 0 6390 0 -1 4570
box -12 -8 92 252
use OAI21X1  _2271_
timestamp 1728305162
transform 1 0 6070 0 -1 4570
box -12 -8 112 252
use MUX2X1  _2272_
timestamp 1728304958
transform 1 0 5670 0 -1 4090
box -12 -8 131 252
use OR2X2  _2273_
timestamp 1728305284
transform 1 0 5470 0 1 3130
box -12 -8 112 252
use NAND2X1  _2274_
timestamp 1728304996
transform 1 0 5250 0 1 3130
box -12 -8 92 252
use NAND2X1  _2275_
timestamp 1728304996
transform 1 0 5730 0 1 3130
box -12 -8 92 252
use NOR2X1  _2276_
timestamp 1728305106
transform -1 0 6410 0 -1 3130
box -12 -8 92 252
use NOR2X1  _2277_
timestamp 1728305106
transform 1 0 7870 0 1 3130
box -12 -8 92 252
use INVX1  _2278_
timestamp 1728304789
transform -1 0 7830 0 -1 3130
box -12 -8 72 252
use OAI21X1  _2279_
timestamp 1728305162
transform 1 0 6570 0 -1 3130
box -12 -8 112 252
use AOI21X1  _2280_
timestamp 1728304211
transform -1 0 6670 0 1 2650
box -12 -8 112 252
use OAI21X1  _2281_
timestamp 1728305162
transform -1 0 6410 0 1 2650
box -12 -8 112 252
use NOR3X1  _2282_
timestamp 1728303224
transform 1 0 6630 0 -1 730
box -12 -8 192 252
use NAND3X1  _2283_
timestamp 1728305047
transform 1 0 7330 0 1 250
box -12 -8 112 252
use NOR2X1  _2284_
timestamp 1728305106
transform 1 0 9270 0 1 250
box -12 -8 92 252
use NAND2X1  _2285_
timestamp 1728304996
transform 1 0 9730 0 1 250
box -12 -8 92 252
use OAI21X1  _2286_
timestamp 1728305162
transform -1 0 2690 0 1 3610
box -12 -8 112 252
use INVX1  _2287_
timestamp 1728304789
transform -1 0 1930 0 1 1210
box -12 -8 72 252
use NOR2X1  _2288_
timestamp 1728305106
transform -1 0 2390 0 1 730
box -12 -8 92 252
use INVX1  _2289_
timestamp 1728304789
transform 1 0 2270 0 1 1690
box -12 -8 72 252
use NOR2X1  _2290_
timestamp 1728305106
transform -1 0 1910 0 1 730
box -12 -8 92 252
use AOI21X1  _2291_
timestamp 1728304211
transform 1 0 2050 0 1 730
box -12 -8 112 252
use OAI21X1  _2292_
timestamp 1728305162
transform 1 0 4190 0 1 250
box -12 -8 112 252
use MUX2X1  _2293_
timestamp 1728304958
transform 1 0 4930 0 1 250
box -12 -8 131 252
use NAND2X1  _2294_
timestamp 1728304996
transform 1 0 6130 0 1 250
box -12 -8 92 252
use NOR2X1  _2295_
timestamp 1728305106
transform -1 0 2390 0 1 1210
box -12 -8 92 252
use OAI21X1  _2296_
timestamp 1728305162
transform 1 0 3770 0 1 730
box -12 -8 112 252
use INVX1  _2297_
timestamp 1728304789
transform 1 0 2290 0 1 250
box -12 -8 72 252
use NOR2X1  _2298_
timestamp 1728305106
transform 1 0 2070 0 1 250
box -12 -8 92 252
use NOR2X1  _2299_
timestamp 1728305106
transform 1 0 3510 0 -1 730
box -12 -8 92 252
use OAI21X1  _2300_
timestamp 1728305162
transform 1 0 3270 0 -1 730
box -12 -8 112 252
use AND2X2  _2301_
timestamp 1728304163
transform -1 0 3810 0 1 250
box -12 -8 112 252
use INVX1  _2302_
timestamp 1728304789
transform 1 0 5190 0 1 250
box -12 -8 72 252
use OAI21X1  _2303_
timestamp 1728305162
transform -1 0 5270 0 -1 730
box -12 -8 112 252
use NAND2X1  _2304_
timestamp 1728304996
transform 1 0 5430 0 -1 730
box -12 -8 92 252
use INVX2  _2305_
timestamp 1728304826
transform -1 0 1650 0 1 2170
box -12 -8 72 252
use OAI21X1  _2306_
timestamp 1728305162
transform 1 0 2530 0 -1 1210
box -12 -8 112 252
use OAI21X1  _2307_
timestamp 1728305162
transform -1 0 5750 0 -1 730
box -12 -8 112 252
use NOR2X1  _2308_
timestamp 1728305106
transform -1 0 5750 0 1 250
box -12 -8 92 252
use NAND2X1  _2309_
timestamp 1728304996
transform 1 0 4690 0 1 250
box -12 -8 92 252
use OAI21X1  _2310_
timestamp 1728305162
transform 1 0 4430 0 1 250
box -12 -8 112 252
use NOR2X1  _2311_
timestamp 1728305106
transform -1 0 3910 0 -1 250
box -12 -8 92 252
use AND2X2  _2312_
timestamp 1728304163
transform -1 0 4150 0 -1 250
box -12 -8 112 252
use AOI21X1  _2313_
timestamp 1728304211
transform 1 0 5370 0 -1 1210
box -12 -8 112 252
use AND2X2  _2314_
timestamp 1728304163
transform 1 0 4550 0 -1 250
box -12 -8 112 252
use NAND3X1  _2315_
timestamp 1728305047
transform 1 0 5490 0 -1 250
box -12 -8 112 252
use AND2X2  _2316_
timestamp 1728304163
transform -1 0 10030 0 1 1210
box -12 -8 112 252
use NOR2X1  _2317_
timestamp 1728305106
transform 1 0 11250 0 1 6010
box -12 -8 92 252
use NOR2X1  _2318_
timestamp 1728305106
transform -1 0 10990 0 -1 4090
box -12 -8 92 252
use OAI21X1  _2319_
timestamp 1728305162
transform -1 0 10650 0 -1 3610
box -12 -8 112 252
use NOR2X1  _2320_
timestamp 1728305106
transform 1 0 10710 0 -1 250
box -12 -8 92 252
use OAI21X1  _2321_
timestamp 1728305162
transform 1 0 10670 0 -1 4090
box -12 -8 112 252
use NAND3X1  _2322_
timestamp 1728305047
transform 1 0 10570 0 1 3610
box -12 -8 112 252
use INVX1  _2323_
timestamp 1728304789
transform 1 0 6810 0 1 2650
box -12 -8 72 252
use NOR2X1  _2324_
timestamp 1728305106
transform 1 0 7030 0 1 2650
box -12 -8 92 252
use NAND2X1  _2325_
timestamp 1728304996
transform 1 0 9390 0 1 6490
box -12 -8 92 252
use NAND2X1  _2326_
timestamp 1728304996
transform -1 0 8970 0 -1 2650
box -12 -8 92 252
use OAI21X1  _2327_
timestamp 1728305162
transform -1 0 9470 0 -1 2650
box -12 -8 112 252
use OAI21X1  _2328_
timestamp 1728305162
transform -1 0 9690 0 -1 2170
box -12 -8 112 252
use OAI21X1  _2329_
timestamp 1728305162
transform 1 0 9350 0 -1 2170
box -12 -8 112 252
use OAI21X1  _2330_
timestamp 1728305162
transform -1 0 9190 0 -1 2170
box -12 -8 112 252
use NOR2X1  _2331_
timestamp 1728305106
transform -1 0 9310 0 1 2170
box -12 -8 92 252
use OAI21X1  _2332_
timestamp 1728305162
transform 1 0 9250 0 1 2650
box -12 -8 112 252
use OR2X2  _2333_
timestamp 1728305284
transform 1 0 9510 0 1 2650
box -12 -8 112 252
use AOI21X1  _2334_
timestamp 1728304211
transform -1 0 9770 0 1 1210
box -12 -8 112 252
use OAI21X1  _2335_
timestamp 1728305162
transform 1 0 5750 0 -1 250
box -12 -8 112 252
use INVX1  _2336_
timestamp 1728304789
transform 1 0 6250 0 -1 250
box -12 -8 72 252
use INVX1  _2337_
timestamp 1728304789
transform -1 0 6090 0 -1 2650
box -12 -8 72 252
use OAI22X1  _2338_
timestamp 1728305200
transform -1 0 6090 0 1 730
box -12 -8 132 252
use OAI21X1  _2339_
timestamp 1728305162
transform 1 0 10450 0 -1 1210
box -12 -8 112 252
use OAI21X1  _2340_
timestamp 1728305162
transform -1 0 9430 0 -1 1690
box -12 -8 112 252
use OAI21X1  _2341_
timestamp 1728305162
transform 1 0 9330 0 1 1690
box -12 -8 112 252
use OR2X2  _2342_
timestamp 1728305284
transform 1 0 10210 0 -1 1210
box -12 -8 112 252
use NAND3X1  _2343_
timestamp 1728305047
transform -1 0 9790 0 -1 1210
box -12 -8 112 252
use NOR2X1  _2344_
timestamp 1728305106
transform 1 0 9790 0 1 730
box -12 -8 92 252
use OR2X2  _2345_
timestamp 1728305284
transform -1 0 7070 0 -1 730
box -12 -8 112 252
use NOR2X1  _2346_
timestamp 1728305106
transform 1 0 6850 0 1 250
box -12 -8 92 252
use NAND2X1  _2347_
timestamp 1728304996
transform -1 0 7230 0 -1 250
box -12 -8 92 252
use NAND3X1  _2348_
timestamp 1728305047
transform 1 0 8190 0 -1 1210
box -12 -8 112 252
use NOR3X1  _2349_
timestamp 1728303224
transform -1 0 8030 0 -1 250
box -12 -8 192 252
use NAND3X1  _2350_
timestamp 1728305047
transform 1 0 7610 0 -1 250
box -12 -8 112 252
use INVX1  _2351_
timestamp 1728304789
transform -1 0 5350 0 -1 250
box -12 -8 72 252
use OR2X2  _2352_
timestamp 1728305284
transform 1 0 5890 0 1 250
box -12 -8 112 252
use NAND2X1  _2353_
timestamp 1728304996
transform -1 0 4390 0 -1 250
box -12 -8 92 252
use NOR2X1  _2354_
timestamp 1728305106
transform 1 0 4810 0 -1 250
box -12 -8 92 252
use NAND3X1  _2355_
timestamp 1728305047
transform -1 0 5130 0 -1 250
box -12 -8 112 252
use NAND3X1  _2356_
timestamp 1728305047
transform 1 0 6010 0 -1 250
box -12 -8 112 252
use AOI22X1  _2357_
timestamp 1728304278
transform -1 0 5850 0 -1 1690
box -14 -8 132 252
use NOR2X1  _2358_
timestamp 1728305106
transform 1 0 7050 0 -1 3130
box -12 -8 92 252
use MUX2X1  _2359_
timestamp 1728304958
transform 1 0 6410 0 -1 2170
box -12 -8 131 252
use AND2X2  _2360_
timestamp 1728304163
transform 1 0 6630 0 1 1690
box -12 -8 112 252
use NAND2X1  _2361_
timestamp 1728304996
transform 1 0 7950 0 -1 3610
box -12 -8 92 252
use NAND2X1  _2362_
timestamp 1728304996
transform 1 0 7470 0 -1 2650
box -12 -8 92 252
use OAI21X1  _2363_
timestamp 1728305162
transform -1 0 7630 0 1 2650
box -12 -8 112 252
use NAND2X1  _2364_
timestamp 1728304996
transform 1 0 8190 0 -1 3610
box -12 -8 92 252
use NOR2X1  _2365_
timestamp 1728305106
transform -1 0 8110 0 1 2170
box -12 -8 92 252
use NOR2X1  _2366_
timestamp 1728305106
transform 1 0 7830 0 1 1690
box -12 -8 92 252
use NAND2X1  _2367_
timestamp 1728304996
transform 1 0 8110 0 -1 730
box -12 -8 92 252
use NOR2X1  _2368_
timestamp 1728305106
transform 1 0 8310 0 1 250
box -12 -8 92 252
use NAND2X1  _2369_
timestamp 1728304996
transform -1 0 10110 0 1 730
box -12 -8 92 252
use NAND3X1  _2370_
timestamp 1728305047
transform 1 0 5450 0 1 730
box -12 -8 112 252
use OAI21X1  _2371_
timestamp 1728305162
transform -1 0 8950 0 1 1690
box -12 -8 112 252
use OAI21X1  _2372_
timestamp 1728305162
transform -1 0 8690 0 1 1690
box -12 -8 112 252
use NAND3X1  _2373_
timestamp 1728305047
transform -1 0 8250 0 1 730
box -12 -8 112 252
use INVX1  _2374_
timestamp 1728304789
transform 1 0 8190 0 -1 250
box -12 -8 72 252
use OR2X2  _2375_
timestamp 1728305284
transform 1 0 6590 0 1 250
box -12 -8 112 252
use NAND3X1  _2376_
timestamp 1728305047
transform 1 0 8530 0 1 250
box -12 -8 112 252
use NOR2X1  _2377_
timestamp 1728305106
transform -1 0 8870 0 1 250
box -12 -8 92 252
use NAND3X1  _2378_
timestamp 1728305047
transform -1 0 9170 0 -1 730
box -12 -8 112 252
use INVX1  _2379_
timestamp 1728304789
transform -1 0 7010 0 -1 250
box -12 -8 72 252
use NOR2X1  _2380_
timestamp 1728305106
transform -1 0 7170 0 1 250
box -12 -8 92 252
use NOR2X1  _2381_
timestamp 1728305106
transform -1 0 7010 0 1 730
box -12 -8 92 252
use INVX1  _2382_
timestamp 1728304789
transform -1 0 8090 0 1 1210
box -12 -8 72 252
use NAND3X1  _2383_
timestamp 1728305047
transform 1 0 7770 0 1 1210
box -12 -8 112 252
use NOR3X1  _2384_
timestamp 1728303224
transform 1 0 7850 0 -1 1210
box -12 -8 192 252
use AND2X2  _2385_
timestamp 1728304163
transform -1 0 7690 0 1 250
box -12 -8 112 252
use NAND3X1  _2386_
timestamp 1728305047
transform -1 0 6790 0 -1 250
box -12 -8 112 252
use NOR2X1  _2387_
timestamp 1728305106
transform -1 0 6550 0 -1 250
box -12 -8 92 252
use OAI21X1  _2388_
timestamp 1728305162
transform -1 0 9130 0 1 250
box -12 -8 112 252
use NAND3X1  _2389_
timestamp 1728305047
transform -1 0 8490 0 1 730
box -12 -8 112 252
use NOR2X1  _2390_
timestamp 1728305106
transform -1 0 8430 0 -1 730
box -12 -8 92 252
use NOR2X1  _2391_
timestamp 1728305106
transform -1 0 9650 0 -1 1690
box -12 -8 92 252
use INVX1  _2392_
timestamp 1728304789
transform 1 0 8370 0 -1 1690
box -12 -8 72 252
use AND2X2  _2393_
timestamp 1728304163
transform 1 0 8330 0 1 1690
box -12 -8 112 252
use NAND3X1  _2394_
timestamp 1728305047
transform 1 0 8950 0 1 1210
box -12 -8 112 252
use NAND3X1  _2395_
timestamp 1728305047
transform 1 0 8930 0 -1 1210
box -12 -8 112 252
use NOR2X1  _2396_
timestamp 1728305106
transform 1 0 9210 0 1 1210
box -12 -8 92 252
use NAND3X1  _2397_
timestamp 1728305047
transform -1 0 9530 0 -1 1210
box -12 -8 112 252
use NOR2X1  _2398_
timestamp 1728305106
transform 1 0 8850 0 -1 730
box -12 -8 92 252
use INVX1  _2399_
timestamp 1728304789
transform -1 0 7750 0 -1 730
box -12 -8 72 252
use NOR2X1  _2400_
timestamp 1728305106
transform 1 0 7470 0 -1 730
box -12 -8 92 252
use NAND3X1  _2401_
timestamp 1728305047
transform 1 0 8590 0 -1 730
box -12 -8 112 252
use INVX1  _2402_
timestamp 1728304789
transform -1 0 6550 0 1 730
box -12 -8 72 252
use NOR2X1  _2403_
timestamp 1728305106
transform -1 0 6790 0 1 730
box -12 -8 92 252
use INVX1  _2404_
timestamp 1728304789
transform -1 0 7730 0 -1 1690
box -12 -8 72 252
use NOR2X1  _2405_
timestamp 1728305106
transform -1 0 7510 0 -1 1690
box -12 -8 92 252
use AND2X2  _2406_
timestamp 1728304163
transform 1 0 7190 0 -1 1690
box -12 -8 112 252
use AND2X2  _2407_
timestamp 1728304163
transform -1 0 6790 0 -1 1690
box -12 -8 112 252
use AND2X2  _2408_
timestamp 1728304163
transform -1 0 6110 0 -1 1690
box -12 -8 112 252
use AND2X2  _2409_
timestamp 1728304163
transform 1 0 7110 0 -1 1210
box -12 -8 112 252
use NOR2X1  _2410_
timestamp 1728305106
transform -1 0 7430 0 1 1690
box -12 -8 92 252
use NOR2X1  _2411_
timestamp 1728305106
transform -1 0 7010 0 -1 2170
box -12 -8 92 252
use NAND2X1  _2412_
timestamp 1728304996
transform -1 0 7670 0 1 1690
box -12 -8 92 252
use OAI21X1  _2413_
timestamp 1728305162
transform 1 0 7110 0 1 1690
box -12 -8 112 252
use NOR2X1  _2414_
timestamp 1728305106
transform 1 0 6950 0 -1 1690
box -12 -8 92 252
use NAND3X1  _2415_
timestamp 1728305047
transform -1 0 8210 0 -1 1690
box -12 -8 112 252
use NOR2X1  _2416_
timestamp 1728305106
transform 1 0 7890 0 -1 1690
box -12 -8 92 252
use NAND2X1  _2417_
timestamp 1728304996
transform -1 0 9190 0 1 730
box -12 -8 92 252
use NOR2X1  _2418_
timestamp 1728305106
transform -1 0 8950 0 1 730
box -12 -8 92 252
use NAND3X1  _2419_
timestamp 1728305047
transform 1 0 7170 0 1 730
box -12 -8 112 252
use INVX1  _2420_
timestamp 1728304789
transform 1 0 2310 0 -1 3130
box -12 -8 72 252
use INVX2  _2421_
timestamp 1728304826
transform -1 0 9830 0 -1 6010
box -12 -8 72 252
use INVX1  _2422_
timestamp 1728304789
transform 1 0 8370 0 -1 5530
box -12 -8 72 252
use NAND3X1  _2423_
timestamp 1728305047
transform 1 0 9070 0 -1 6010
box -12 -8 112 252
use OAI21X1  _2424_
timestamp 1728305162
transform 1 0 8870 0 1 6010
box -12 -8 112 252
use INVX1  _2425_
timestamp 1728304789
transform 1 0 3270 0 1 2650
box -12 -8 72 252
use OAI21X1  _2426_
timestamp 1728305162
transform 1 0 8830 0 -1 6010
box -12 -8 112 252
use INVX1  _2427_
timestamp 1728304789
transform 1 0 8930 0 1 5530
box -12 -8 72 252
use NOR2X1  _2428_
timestamp 1728305106
transform 1 0 9310 0 -1 6010
box -12 -8 92 252
use INVX1  _2429_
timestamp 1728304789
transform 1 0 9550 0 -1 6010
box -12 -8 72 252
use INVX2  _2430_
timestamp 1728304826
transform 1 0 8910 0 -1 6970
box -12 -8 72 252
use OAI21X1  _2431_
timestamp 1728305162
transform -1 0 9430 0 1 6010
box -12 -8 112 252
use NOR2X1  _2432_
timestamp 1728305106
transform 1 0 9590 0 1 6010
box -12 -8 92 252
use AOI22X1  _2433_
timestamp 1728304278
transform -1 0 10110 0 -1 6010
box -14 -8 132 252
use NAND2X1  _2434_
timestamp 1728304996
transform -1 0 10130 0 1 6010
box -12 -8 92 252
use INVX1  _2435_
timestamp 1728304789
transform 1 0 4550 0 1 4570
box -12 -8 72 252
use NOR2X1  _2436_
timestamp 1728305106
transform 1 0 9290 0 -1 6490
box -12 -8 92 252
use OAI21X1  _2437_
timestamp 1728305162
transform 1 0 10990 0 1 4570
box -12 -8 112 252
use OAI21X1  _2438_
timestamp 1728305162
transform -1 0 11130 0 -1 5050
box -12 -8 112 252
use NAND3X1  _2439_
timestamp 1728305047
transform -1 0 11090 0 -1 5530
box -12 -8 112 252
use OAI21X1  _2440_
timestamp 1728305162
transform 1 0 9150 0 1 5530
box -12 -8 112 252
use OAI21X1  _2441_
timestamp 1728305162
transform -1 0 6350 0 -1 5530
box -12 -8 112 252
use NAND2X1  _2442_
timestamp 1728304996
transform -1 0 8430 0 1 6970
box -12 -8 92 252
use OAI21X1  _2443_
timestamp 1728305162
transform 1 0 3930 0 -1 7930
box -12 -8 112 252
use INVX1  _2444_
timestamp 1728304789
transform -1 0 4830 0 1 5530
box -12 -8 72 252
use NAND2X1  _2445_
timestamp 1728304996
transform -1 0 8770 0 1 5530
box -12 -8 92 252
use OAI21X1  _2446_
timestamp 1728305162
transform 1 0 8350 0 -1 6010
box -12 -8 112 252
use AOI22X1  _2447_
timestamp 1728304278
transform 1 0 8170 0 -1 6970
box -14 -8 132 252
use NAND3X1  _2448_
timestamp 1728305047
transform 1 0 8590 0 1 6970
box -12 -8 112 252
use INVX1  _2449_
timestamp 1728304789
transform -1 0 8890 0 1 6970
box -12 -8 72 252
use OAI21X1  _2450_
timestamp 1728305162
transform -1 0 9150 0 1 6970
box -12 -8 112 252
use OAI21X1  _2451_
timestamp 1728305162
transform 1 0 3930 0 1 7930
box -12 -8 112 252
use NOR2X1  _2452_
timestamp 1728305106
transform 1 0 7690 0 -1 6010
box -12 -8 92 252
use OAI21X1  _2453_
timestamp 1728305162
transform -1 0 6810 0 -1 6010
box -12 -8 112 252
use AOI22X1  _2454_
timestamp 1728304278
transform -1 0 6550 0 -1 7450
box -14 -8 132 252
use NAND3X1  _2455_
timestamp 1728305047
transform -1 0 6790 0 -1 7450
box -12 -8 112 252
use INVX1  _2456_
timestamp 1728304789
transform -1 0 8890 0 -1 7450
box -12 -8 72 252
use OAI21X1  _2457_
timestamp 1728305162
transform -1 0 9130 0 -1 7450
box -12 -8 112 252
use NAND2X1  _2458_
timestamp 1728304996
transform -1 0 6970 0 -1 7930
box -12 -8 92 252
use OAI21X1  _2459_
timestamp 1728305162
transform -1 0 3770 0 -1 7930
box -12 -8 112 252
use AOI22X1  _2460_
timestamp 1728304278
transform 1 0 7190 0 -1 7450
box -14 -8 132 252
use NAND3X1  _2461_
timestamp 1728305047
transform 1 0 7130 0 -1 7930
box -12 -8 112 252
use INVX1  _2462_
timestamp 1728304789
transform -1 0 7450 0 -1 7930
box -12 -8 72 252
use OAI21X1  _2463_
timestamp 1728305162
transform -1 0 7490 0 1 7450
box -12 -8 112 252
use INVX1  _2464_
timestamp 1728304789
transform 1 0 4590 0 1 5050
box -12 -8 72 252
use INVX1  _2465_
timestamp 1728304789
transform -1 0 7510 0 -1 7450
box -12 -8 72 252
use OAI21X1  _2466_
timestamp 1728305162
transform -1 0 3550 0 1 7930
box -12 -8 112 252
use OAI21X1  _2467_
timestamp 1728305162
transform 1 0 6290 0 1 7930
box -12 -8 112 252
use AOI21X1  _2468_
timestamp 1728304211
transform -1 0 6470 0 -1 7930
box -12 -8 112 252
use OAI21X1  _2469_
timestamp 1728305162
transform -1 0 6330 0 1 7450
box -12 -8 112 252
use INVX1  _2470_
timestamp 1728304789
transform -1 0 6530 0 1 7450
box -12 -8 72 252
use OAI21X1  _2471_
timestamp 1728305162
transform -1 0 8250 0 1 7450
box -12 -8 112 252
use AOI21X1  _2472_
timestamp 1728304211
transform -1 0 6270 0 -1 7450
box -12 -8 112 252
use OAI21X1  _2473_
timestamp 1728305162
transform -1 0 5590 0 1 7450
box -12 -8 112 252
use INVX1  _2474_
timestamp 1728304789
transform -1 0 5490 0 -1 8890
box -12 -8 72 252
use OAI21X1  _2475_
timestamp 1728305162
transform -1 0 7990 0 1 5050
box -12 -8 112 252
use OAI21X1  _2476_
timestamp 1728305162
transform -1 0 2890 0 -1 8410
box -12 -8 112 252
use OAI21X1  _2477_
timestamp 1728305162
transform -1 0 5390 0 1 7930
box -12 -8 112 252
use NOR2X1  _2478_
timestamp 1728305106
transform 1 0 5370 0 -1 7930
box -12 -8 92 252
use OAI21X1  _2479_
timestamp 1728305162
transform -1 0 8210 0 -1 7930
box -12 -8 112 252
use OAI21X1  _2480_
timestamp 1728305162
transform 1 0 6030 0 1 7930
box -12 -8 112 252
use INVX1  _2481_
timestamp 1728304789
transform 1 0 4270 0 -1 8890
box -12 -8 72 252
use OAI21X1  _2482_
timestamp 1728305162
transform -1 0 2650 0 -1 8410
box -12 -8 112 252
use OAI21X1  _2483_
timestamp 1728305162
transform -1 0 4890 0 -1 8410
box -12 -8 112 252
use NOR2X1  _2484_
timestamp 1728305106
transform -1 0 5890 0 -1 8410
box -12 -8 92 252
use OAI21X1  _2485_
timestamp 1728305162
transform -1 0 7170 0 -1 8410
box -12 -8 112 252
use OAI21X1  _2486_
timestamp 1728305162
transform 1 0 3190 0 1 7930
box -12 -8 112 252
use OAI21X1  _2487_
timestamp 1728305162
transform -1 0 5870 0 1 7930
box -12 -8 112 252
use AOI21X1  _2488_
timestamp 1728304211
transform 1 0 6550 0 1 7930
box -12 -8 112 252
use OAI21X1  _2489_
timestamp 1728305162
transform -1 0 6890 0 1 7930
box -12 -8 112 252
use INVX1  _2490_
timestamp 1728304789
transform 1 0 7810 0 1 7930
box -12 -8 72 252
use OAI21X1  _2491_
timestamp 1728305162
transform -1 0 8130 0 1 7930
box -12 -8 112 252
use OAI21X1  _2492_
timestamp 1728305162
transform -1 0 3050 0 1 7930
box -12 -8 112 252
use OAI21X1  _2493_
timestamp 1728305162
transform -1 0 5710 0 -1 7930
box -12 -8 112 252
use AOI21X1  _2494_
timestamp 1728304211
transform -1 0 6770 0 1 7450
box -12 -8 112 252
use OAI21X1  _2495_
timestamp 1728305162
transform 1 0 6950 0 -1 7450
box -12 -8 112 252
use INVX1  _2496_
timestamp 1728304789
transform 1 0 7670 0 -1 7450
box -12 -8 72 252
use OAI21X1  _2497_
timestamp 1728305162
transform -1 0 7970 0 -1 7450
box -12 -8 112 252
use OAI21X1  _2498_
timestamp 1728305162
transform -1 0 8970 0 -1 5050
box -12 -8 112 252
use NOR2X1  _2499_
timestamp 1728305106
transform 1 0 9110 0 1 6010
box -12 -8 92 252
use INVX2  _2500_
timestamp 1728304826
transform -1 0 7790 0 1 6490
box -12 -8 72 252
use OAI21X1  _2501_
timestamp 1728305162
transform -1 0 6950 0 -1 4090
box -12 -8 112 252
use NAND2X1  _2502_
timestamp 1728304996
transform -1 0 7770 0 -1 5530
box -12 -8 92 252
use NAND3X1  _2503_
timestamp 1728305047
transform 1 0 11230 0 -1 6010
box -12 -8 112 252
use NOR2X1  _2504_
timestamp 1728305106
transform -1 0 4730 0 -1 7450
box -12 -8 92 252
use INVX2  _2505_
timestamp 1728304826
transform -1 0 5830 0 -1 6970
box -12 -8 72 252
use NOR2X1  _2506_
timestamp 1728305106
transform -1 0 6890 0 -1 4570
box -12 -8 92 252
use NAND2X1  _2507_
timestamp 1728304996
transform 1 0 5950 0 -1 6490
box -12 -8 92 252
use NOR2X1  _2508_
timestamp 1728305106
transform 1 0 5770 0 1 6490
box -12 -8 92 252
use OAI21X1  _2509_
timestamp 1728305162
transform -1 0 9010 0 -1 4570
box -12 -8 112 252
use NAND3X1  _2510_
timestamp 1728305047
transform -1 0 8250 0 -1 4570
box -12 -8 112 252
use NOR2X1  _2511_
timestamp 1728305106
transform -1 0 7570 0 -1 4570
box -12 -8 92 252
use NAND3X1  _2512_
timestamp 1728305047
transform 1 0 7210 0 -1 3610
box -12 -8 112 252
use NOR2X1  _2513_
timestamp 1728305106
transform 1 0 6970 0 -1 3610
box -12 -8 92 252
use NAND2X1  _2514_
timestamp 1728304996
transform 1 0 7150 0 -1 5050
box -12 -8 92 252
use NAND2X1  _2515_
timestamp 1728304996
transform 1 0 10470 0 1 5530
box -12 -8 92 252
use INVX1  _2516_
timestamp 1728304789
transform 1 0 8630 0 -1 6490
box -12 -8 72 252
use NAND3X1  _2517_
timestamp 1728305047
transform 1 0 10730 0 -1 6010
box -12 -8 112 252
use OAI22X1  _2518_
timestamp 1728305200
transform -1 0 9910 0 1 4090
box -12 -8 132 252
use OR2X2  _2519_
timestamp 1728305284
transform 1 0 10070 0 1 4090
box -12 -8 112 252
use NOR2X1  _2520_
timestamp 1728305106
transform -1 0 10570 0 -1 6010
box -12 -8 92 252
use OAI21X1  _2521_
timestamp 1728305162
transform -1 0 8710 0 1 6010
box -12 -8 112 252
use NOR2X1  _2522_
timestamp 1728305106
transform 1 0 6190 0 -1 6490
box -12 -8 92 252
use NAND2X1  _2523_
timestamp 1728304996
transform 1 0 5990 0 1 6490
box -12 -8 92 252
use NAND2X1  _2524_
timestamp 1728304996
transform 1 0 8390 0 -1 6490
box -12 -8 92 252
use OAI21X1  _2525_
timestamp 1728305162
transform 1 0 6890 0 1 6010
box -12 -8 112 252
use OAI21X1  _2526_
timestamp 1728305162
transform -1 0 7950 0 1 6010
box -12 -8 112 252
use AOI21X1  _2527_
timestamp 1728304211
transform 1 0 8110 0 1 6010
box -12 -8 112 252
use AND2X2  _2528_
timestamp 1728304163
transform -1 0 8230 0 -1 6490
box -12 -8 112 252
use OAI21X1  _2529_
timestamp 1728305162
transform 1 0 7950 0 1 6490
box -12 -8 112 252
use AOI21X1  _2530_
timestamp 1728304211
transform -1 0 7990 0 -1 6490
box -12 -8 112 252
use INVX1  _2531_
timestamp 1728304789
transform -1 0 7950 0 -1 730
box -12 -8 72 252
use OAI21X1  _2532_
timestamp 1728305162
transform 1 0 7930 0 -1 6970
box -12 -8 112 252
use INVX1  _2533_
timestamp 1728304789
transform -1 0 5630 0 -1 6970
box -12 -8 72 252
use AOI22X1  _2534_
timestamp 1728304278
transform -1 0 6090 0 -1 6970
box -14 -8 132 252
use AND2X2  _2535_
timestamp 1728304163
transform -1 0 7770 0 -1 6970
box -12 -8 112 252
use OAI21X1  _2536_
timestamp 1728305162
transform 1 0 7470 0 1 6970
box -12 -8 112 252
use AOI21X1  _2537_
timestamp 1728304211
transform 1 0 7410 0 -1 6970
box -12 -8 112 252
use INVX1  _2538_
timestamp 1728304789
transform 1 0 8130 0 -1 6010
box -12 -8 72 252
use OAI21X1  _2539_
timestamp 1728305162
transform 1 0 5970 0 1 6970
box -12 -8 112 252
use AOI22X1  _2540_
timestamp 1728304278
transform 1 0 5710 0 1 6970
box -14 -8 132 252
use AND2X2  _2541_
timestamp 1728304163
transform 1 0 6230 0 1 6970
box -12 -8 112 252
use OAI21X1  _2542_
timestamp 1728305162
transform -1 0 6830 0 1 6970
box -12 -8 112 252
use AOI21X1  _2543_
timestamp 1728304211
transform -1 0 6810 0 1 6490
box -12 -8 112 252
use INVX1  _2544_
timestamp 1728304789
transform 1 0 6250 0 -1 1690
box -12 -8 72 252
use OR2X2  _2545_
timestamp 1728305284
transform 1 0 6970 0 1 6490
box -12 -8 112 252
use INVX1  _2546_
timestamp 1728304789
transform 1 0 6230 0 1 6490
box -12 -8 72 252
use OAI22X1  _2547_
timestamp 1728305200
transform 1 0 6430 0 1 6490
box -12 -8 132 252
use AOI21X1  _2548_
timestamp 1728304211
transform 1 0 7230 0 1 6490
box -12 -8 112 252
use OAI21X1  _2549_
timestamp 1728305162
transform 1 0 7470 0 1 6490
box -12 -8 112 252
use AOI21X1  _2550_
timestamp 1728304211
transform -1 0 7730 0 -1 6490
box -12 -8 112 252
use INVX1  _2551_
timestamp 1728304789
transform -1 0 6410 0 1 2170
box -12 -8 72 252
use NAND2X1  _2552_
timestamp 1728304996
transform -1 0 4970 0 -1 7930
box -12 -8 92 252
use INVX1  _2553_
timestamp 1728304789
transform -1 0 6010 0 -1 7450
box -12 -8 72 252
use OAI22X1  _2554_
timestamp 1728305200
transform -1 0 5790 0 -1 7450
box -12 -8 132 252
use AOI21X1  _2555_
timestamp 1728304211
transform 1 0 5730 0 1 7450
box -12 -8 112 252
use AND2X2  _2556_
timestamp 1728304163
transform 1 0 5130 0 -1 7930
box -12 -8 112 252
use OAI21X1  _2557_
timestamp 1728305162
transform 1 0 5850 0 -1 7930
box -12 -8 112 252
use AOI21X1  _2558_
timestamp 1728304211
transform -1 0 6590 0 1 6970
box -12 -8 112 252
use INVX1  _2559_
timestamp 1728304789
transform 1 0 6190 0 -1 4090
box -12 -8 72 252
use NAND2X1  _2560_
timestamp 1728304996
transform 1 0 4430 0 -1 7930
box -12 -8 92 252
use INVX1  _2561_
timestamp 1728304789
transform -1 0 5550 0 1 6970
box -12 -8 72 252
use OAI22X1  _2562_
timestamp 1728305200
transform 1 0 5130 0 -1 7450
box -12 -8 132 252
use AOI21X1  _2563_
timestamp 1728304211
transform -1 0 5090 0 1 7450
box -12 -8 112 252
use NAND2X1  _2564_
timestamp 1728304996
transform -1 0 4750 0 -1 7930
box -12 -8 92 252
use INVX1  _2565_
timestamp 1728304789
transform 1 0 4810 0 1 7930
box -12 -8 72 252
use OAI21X1  _2566_
timestamp 1728305162
transform -1 0 5130 0 1 7930
box -12 -8 112 252
use AOI21X1  _2567_
timestamp 1728304211
transform 1 0 5250 0 1 7450
box -12 -8 112 252
use INVX1  _2568_
timestamp 1728304789
transform 1 0 5370 0 -1 5530
box -12 -8 72 252
use OAI21X1  _2569_
timestamp 1728305162
transform -1 0 4350 0 1 7450
box -12 -8 112 252
use AOI22X1  _2570_
timestamp 1728304278
transform 1 0 5290 0 -1 6970
box -14 -8 132 252
use AND2X2  _2571_
timestamp 1728304163
transform 1 0 4390 0 -1 7450
box -12 -8 112 252
use OAI21X1  _2572_
timestamp 1728305162
transform -1 0 4610 0 1 7450
box -12 -8 112 252
use AOI21X1  _2573_
timestamp 1728304211
transform 1 0 4750 0 1 7450
box -12 -8 112 252
use INVX1  _2574_
timestamp 1728304789
transform 1 0 5490 0 -1 6010
box -12 -8 72 252
use OAI21X1  _2575_
timestamp 1728305162
transform -1 0 5130 0 -1 6970
box -12 -8 112 252
use AOI22X1  _2576_
timestamp 1728304278
transform 1 0 5210 0 1 6970
box -14 -8 132 252
use AND2X2  _2577_
timestamp 1728304163
transform 1 0 4970 0 1 6970
box -12 -8 112 252
use OAI21X1  _2578_
timestamp 1728305162
transform -1 0 4970 0 -1 7450
box -12 -8 112 252
use AOI21X1  _2579_
timestamp 1728304211
transform 1 0 4770 0 -1 6970
box -12 -8 112 252
use INVX1  _2580_
timestamp 1728304789
transform 1 0 4810 0 -1 5050
box -12 -8 72 252
use INVX2  _2581_
timestamp 1728304826
transform -1 0 4270 0 1 9850
box -12 -8 72 252
use INVX1  _2582_
timestamp 1728304789
transform -1 0 3430 0 -1 8890
box -12 -8 72 252
use INVX2  _2583_
timestamp 1728304826
transform 1 0 2330 0 -1 8410
box -12 -8 72 252
use OAI21X1  _2584_
timestamp 1728305162
transform 1 0 3270 0 -1 8410
box -12 -8 112 252
use INVX2  _2585_
timestamp 1728304826
transform -1 0 6490 0 -1 6490
box -12 -8 72 252
use AOI22X1  _2586_
timestamp 1728304278
transform -1 0 3890 0 -1 8410
box -14 -8 132 252
use NAND3X1  _2587_
timestamp 1728305047
transform -1 0 3630 0 -1 8410
box -12 -8 112 252
use NOR2X1  _2588_
timestamp 1728305106
transform -1 0 3130 0 -1 8410
box -12 -8 92 252
use OAI21X1  _2589_
timestamp 1728305162
transform -1 0 3130 0 1 8410
box -12 -8 112 252
use INVX1  _2590_
timestamp 1728304789
transform 1 0 3690 0 -1 11290
box -12 -8 72 252
use AOI21X1  _2591_
timestamp 1728304211
transform -1 0 3250 0 1 9370
box -12 -8 112 252
use OAI21X1  _2592_
timestamp 1728305162
transform 1 0 2650 0 1 9370
box -12 -8 112 252
use AOI21X1  _2593_
timestamp 1728304211
transform -1 0 2850 0 1 9850
box -12 -8 112 252
use OAI21X1  _2594_
timestamp 1728305162
transform -1 0 2850 0 -1 10330
box -12 -8 112 252
use INVX1  _2595_
timestamp 1728304789
transform -1 0 3910 0 1 10810
box -12 -8 72 252
use AOI22X1  _2596_
timestamp 1728304278
transform 1 0 3470 0 1 9850
box -14 -8 132 252
use OAI21X1  _2597_
timestamp 1728305162
transform 1 0 3390 0 1 9370
box -12 -8 112 252
use NAND2X1  _2598_
timestamp 1728304996
transform -1 0 3350 0 -1 9850
box -12 -8 92 252
use INVX1  _2599_
timestamp 1728304789
transform -1 0 3310 0 1 9850
box -12 -8 72 252
use OAI21X1  _2600_
timestamp 1728305162
transform 1 0 3010 0 1 9850
box -12 -8 112 252
use INVX2  _2601_
timestamp 1728304826
transform -1 0 2610 0 -1 10330
box -12 -8 72 252
use AOI22X1  _2602_
timestamp 1728304278
transform -1 0 2910 0 -1 9850
box -14 -8 132 252
use OAI21X1  _2603_
timestamp 1728305162
transform -1 0 2510 0 1 9370
box -12 -8 112 252
use NAND2X1  _2604_
timestamp 1728304996
transform 1 0 2570 0 -1 9850
box -12 -8 92 252
use INVX1  _2605_
timestamp 1728304789
transform -1 0 2590 0 1 9850
box -12 -8 72 252
use OAI21X1  _2606_
timestamp 1728305162
transform 1 0 2290 0 -1 10330
box -12 -8 112 252
use INVX1  _2607_
timestamp 1728304789
transform -1 0 1670 0 -1 10330
box -12 -8 72 252
use INVX1  _2608_
timestamp 1728304789
transform -1 0 1210 0 1 9370
box -12 -8 72 252
use AOI22X1  _2609_
timestamp 1728304278
transform 1 0 2130 0 1 9370
box -14 -8 132 252
use OAI21X1  _2610_
timestamp 1728305162
transform 1 0 1350 0 1 9370
box -12 -8 112 252
use AOI21X1  _2611_
timestamp 1728304211
transform -1 0 1430 0 -1 9850
box -12 -8 112 252
use OAI21X1  _2612_
timestamp 1728305162
transform -1 0 1170 0 -1 9850
box -12 -8 112 252
use INVX1  _2613_
timestamp 1728304789
transform -1 0 2090 0 1 10330
box -12 -8 72 252
use INVX1  _2614_
timestamp 1728304789
transform -1 0 730 0 1 9370
box -12 -8 72 252
use AOI22X1  _2615_
timestamp 1728304278
transform 1 0 1850 0 1 9370
box -14 -8 132 252
use OAI21X1  _2616_
timestamp 1728305162
transform 1 0 1610 0 1 9370
box -12 -8 112 252
use AOI21X1  _2617_
timestamp 1728304211
transform -1 0 1690 0 -1 9850
box -12 -8 112 252
use OAI21X1  _2618_
timestamp 1728305162
transform -1 0 1910 0 1 9850
box -12 -8 112 252
use INVX1  _2619_
timestamp 1728304789
transform 1 0 890 0 1 8890
box -12 -8 72 252
use AOI21X1  _2620_
timestamp 1728304211
transform -1 0 1490 0 1 8410
box -12 -8 112 252
use OAI21X1  _2621_
timestamp 1728305162
transform 1 0 1130 0 1 8410
box -12 -8 112 252
use AOI21X1  _2622_
timestamp 1728304211
transform -1 0 1450 0 1 8890
box -12 -8 112 252
use OAI21X1  _2623_
timestamp 1728305162
transform 1 0 1090 0 1 8890
box -12 -8 112 252
use INVX1  _2624_
timestamp 1728304789
transform -1 0 690 0 -1 9850
box -12 -8 72 252
use AOI21X1  _2625_
timestamp 1728304211
transform -1 0 2810 0 1 7930
box -12 -8 112 252
use OAI21X1  _2626_
timestamp 1728305162
transform 1 0 1730 0 1 7930
box -12 -8 112 252
use AOI21X1  _2627_
timestamp 1728304211
transform 1 0 1490 0 1 7930
box -12 -8 112 252
use OAI21X1  _2628_
timestamp 1728305162
transform 1 0 870 0 -1 8890
box -12 -8 112 252
use INVX1  _2629_
timestamp 1728304789
transform -1 0 3530 0 -1 4090
box -12 -8 72 252
use NOR2X1  _2630_
timestamp 1728305106
transform 1 0 4350 0 1 5050
box -12 -8 92 252
use INVX1  _2631_
timestamp 1728304789
transform -1 0 5030 0 1 5530
box -12 -8 72 252
use NOR2X1  _2632_
timestamp 1728305106
transform 1 0 10990 0 -1 6010
box -12 -8 92 252
use INVX1  _2633_
timestamp 1728304789
transform 1 0 3990 0 -1 3130
box -12 -8 72 252
use NOR2X1  _2634_
timestamp 1728305106
transform 1 0 9070 0 -1 6490
box -12 -8 92 252
use INVX8  _2635_
timestamp 1728304916
transform -1 0 2470 0 -1 5050
box -12 -8 133 252
use OAI21X1  _2636_
timestamp 1728305162
transform -1 0 9310 0 -1 4090
box -12 -8 112 252
use NOR2X1  _2637_
timestamp 1728305106
transform 1 0 4450 0 -1 9370
box -12 -8 92 252
use INVX1  _2638_
timestamp 1728304789
transform 1 0 4950 0 -1 9370
box -12 -8 72 252
use OAI21X1  _2639_
timestamp 1728305162
transform -1 0 10090 0 1 4570
box -12 -8 112 252
use OAI21X1  _2640_
timestamp 1728305162
transform -1 0 10050 0 1 5530
box -12 -8 112 252
use NOR2X1  _2641_
timestamp 1728305106
transform 1 0 10270 0 -1 6010
box -12 -8 92 252
use AOI21X1  _2642_
timestamp 1728304211
transform -1 0 9670 0 -1 5050
box -12 -8 112 252
use NOR2X1  _2643_
timestamp 1728305106
transform 1 0 11010 0 1 6010
box -12 -8 92 252
use AND2X2  _2644_
timestamp 1728304163
transform -1 0 9910 0 1 6010
box -12 -8 112 252
use NAND3X1  _2645_
timestamp 1728305047
transform -1 0 9890 0 -1 6490
box -12 -8 112 252
use OAI22X1  _2646_
timestamp 1728305200
transform 1 0 10210 0 1 5530
box -12 -8 132 252
use NAND3X1  _2647_
timestamp 1728305047
transform -1 0 8750 0 1 6490
box -12 -8 112 252
use NOR2X1  _2648_
timestamp 1728305106
transform -1 0 4330 0 1 6970
box -12 -8 92 252
use AOI22X1  _2649_
timestamp 1728304278
transform -1 0 5990 0 -1 8890
box -14 -8 132 252
use AOI22X1  _2650_
timestamp 1728304278
transform 1 0 9410 0 1 5530
box -14 -8 132 252
use NOR3X1  _2651_
timestamp 1728303224
transform -1 0 5950 0 1 8890
box -12 -8 192 252
use OAI21X1  _2652_
timestamp 1728305162
transform -1 0 8010 0 -1 5530
box -12 -8 112 252
use AOI21X1  _2653_
timestamp 1728304211
transform -1 0 7930 0 1 5530
box -12 -8 112 252
use OAI21X1  _2654_
timestamp 1728305162
transform 1 0 4770 0 1 8890
box -12 -8 112 252
use AOI21X1  _2655_
timestamp 1728304211
transform -1 0 5610 0 1 8890
box -12 -8 112 252
use OAI21X1  _2656_
timestamp 1728305162
transform -1 0 6210 0 1 8890
box -12 -8 112 252
use NOR2X1  _2657_
timestamp 1728305106
transform -1 0 6910 0 1 8890
box -12 -8 92 252
use AND2X2  _2658_
timestamp 1728304163
transform 1 0 6370 0 1 8890
box -12 -8 112 252
use OR2X2  _2659_
timestamp 1728305284
transform 1 0 7070 0 1 8890
box -12 -8 112 252
use OAI22X1  _2660_
timestamp 1728305200
transform -1 0 7430 0 1 8890
box -12 -8 132 252
use NAND2X1  _2661_
timestamp 1728304996
transform -1 0 4630 0 -1 8410
box -12 -8 92 252
use OAI21X1  _2662_
timestamp 1728305162
transform 1 0 4530 0 1 8410
box -12 -8 112 252
use AOI21X1  _2663_
timestamp 1728304211
transform 1 0 6430 0 -1 9370
box -12 -8 112 252
use OAI21X1  _2664_
timestamp 1728305162
transform -1 0 6790 0 -1 9370
box -12 -8 112 252
use NOR2X1  _2665_
timestamp 1728305106
transform 1 0 7190 0 -1 9370
box -12 -8 92 252
use NAND3X1  _2666_
timestamp 1728305047
transform 1 0 6950 0 -1 9370
box -12 -8 112 252
use NAND2X1  _2667_
timestamp 1728304996
transform 1 0 7690 0 -1 9370
box -12 -8 92 252
use OAI22X1  _2668_
timestamp 1728305200
transform 1 0 7410 0 -1 9370
box -12 -8 132 252
use INVX1  _2669_
timestamp 1728304789
transform 1 0 8090 0 1 9850
box -12 -8 72 252
use OAI21X1  _2670_
timestamp 1728305162
transform -1 0 4390 0 -1 8410
box -12 -8 112 252
use AOI22X1  _2671_
timestamp 1728304278
transform -1 0 5510 0 -1 7450
box -14 -8 132 252
use NAND2X1  _2672_
timestamp 1728304996
transform 1 0 5330 0 -1 8410
box -12 -8 92 252
use INVX1  _2673_
timestamp 1728304789
transform 1 0 7270 0 -1 9850
box -12 -8 72 252
use OAI21X1  _2674_
timestamp 1728305162
transform -1 0 7590 0 -1 9850
box -12 -8 112 252
use NOR2X1  _2675_
timestamp 1728305106
transform 1 0 7750 0 -1 9850
box -12 -8 92 252
use INVX1  _2676_
timestamp 1728304789
transform -1 0 7710 0 -1 10330
box -12 -8 72 252
use OAI21X1  _2677_
timestamp 1728305162
transform 1 0 7870 0 -1 10330
box -12 -8 112 252
use OAI22X1  _2678_
timestamp 1728305200
transform 1 0 7810 0 1 9850
box -12 -8 132 252
use NOR2X1  _2679_
timestamp 1728305106
transform 1 0 4270 0 1 8890
box -12 -8 92 252
use NAND3X1  _2680_
timestamp 1728305047
transform -1 0 4610 0 1 8890
box -12 -8 112 252
use INVX2  _2681_
timestamp 1728304826
transform 1 0 6210 0 1 9370
box -12 -8 72 252
use AOI21X1  _2682_
timestamp 1728304211
transform 1 0 6850 0 1 9850
box -12 -8 112 252
use INVX1  _2683_
timestamp 1728304789
transform 1 0 4190 0 1 7930
box -12 -8 72 252
use AOI21X1  _2684_
timestamp 1728304211
transform -1 0 5910 0 1 8410
box -12 -8 112 252
use OAI21X1  _2685_
timestamp 1728305162
transform 1 0 5570 0 1 8410
box -12 -8 112 252
use NOR2X1  _2686_
timestamp 1728305106
transform -1 0 7030 0 -1 10330
box -12 -8 92 252
use INVX1  _2687_
timestamp 1728304789
transform 1 0 7450 0 -1 10330
box -12 -8 72 252
use AOI21X1  _2688_
timestamp 1728304211
transform -1 0 7670 0 1 9850
box -12 -8 112 252
use AOI21X1  _2689_
timestamp 1728304211
transform 1 0 6590 0 1 9850
box -12 -8 112 252
use OAI22X1  _2690_
timestamp 1728305200
transform 1 0 6690 0 -1 10330
box -12 -8 132 252
use OAI21X1  _2691_
timestamp 1728305162
transform 1 0 7190 0 -1 10330
box -12 -8 112 252
use OAI22X1  _2692_
timestamp 1728305200
transform -1 0 7410 0 1 9850
box -12 -8 132 252
use NAND3X1  _2693_
timestamp 1728305047
transform 1 0 5170 0 -1 9370
box -12 -8 112 252
use NOR2X1  _2694_
timestamp 1728305106
transform -1 0 5350 0 1 9370
box -12 -8 92 252
use OAI21X1  _2695_
timestamp 1728305162
transform 1 0 6750 0 -1 9850
box -12 -8 112 252
use OAI21X1  _2696_
timestamp 1728305162
transform 1 0 6690 0 1 9370
box -12 -8 112 252
use INVX1  _2697_
timestamp 1728304789
transform 1 0 7090 0 1 9850
box -12 -8 72 252
use AOI22X1  _2698_
timestamp 1728304278
transform 1 0 7010 0 -1 9850
box -14 -8 132 252
use NAND3X1  _2699_
timestamp 1728305047
transform -1 0 6530 0 1 9370
box -12 -8 112 252
use OAI21X1  _2700_
timestamp 1728305162
transform 1 0 5490 0 1 9370
box -12 -8 112 252
use AOI21X1  _2701_
timestamp 1728304211
transform -1 0 5670 0 -1 8410
box -12 -8 112 252
use OAI21X1  _2702_
timestamp 1728305162
transform -1 0 5730 0 -1 8890
box -12 -8 112 252
use AOI21X1  _2703_
timestamp 1728304211
transform -1 0 5770 0 -1 9370
box -12 -8 112 252
use AND2X2  _2704_
timestamp 1728304163
transform 1 0 5750 0 -1 9850
box -12 -8 112 252
use OAI21X1  _2705_
timestamp 1728305162
transform 1 0 5990 0 -1 9850
box -12 -8 112 252
use OAI22X1  _2706_
timestamp 1728305200
transform -1 0 6370 0 -1 9850
box -12 -8 132 252
use AOI21X1  _2707_
timestamp 1728304211
transform -1 0 6070 0 1 9370
box -12 -8 112 252
use INVX2  _2708_
timestamp 1728304826
transform -1 0 2450 0 1 8410
box -12 -8 72 252
use OAI21X1  _2709_
timestamp 1728305162
transform -1 0 5150 0 1 8410
box -12 -8 112 252
use INVX1  _2710_
timestamp 1728304789
transform -1 0 5010 0 -1 8890
box -12 -8 72 252
use OAI21X1  _2711_
timestamp 1728305162
transform -1 0 5270 0 -1 8890
box -12 -8 112 252
use NOR2X1  _2712_
timestamp 1728305106
transform -1 0 5830 0 1 9370
box -12 -8 92 252
use OAI21X1  _2713_
timestamp 1728305162
transform -1 0 5970 0 1 9850
box -12 -8 112 252
use AOI21X1  _2714_
timestamp 1728304211
transform -1 0 6290 0 -1 9370
box -12 -8 112 252
use OAI22X1  _2715_
timestamp 1728305200
transform 1 0 5910 0 -1 9370
box -12 -8 132 252
use NOR3X1  _2716_
timestamp 1728303224
transform -1 0 6930 0 1 10330
box -12 -8 192 252
use INVX1  _2717_
timestamp 1728304789
transform 1 0 6710 0 -1 10810
box -12 -8 72 252
use NAND3X1  _2718_
timestamp 1728305047
transform 1 0 6270 0 1 10330
box -12 -8 112 252
use OAI21X1  _2719_
timestamp 1728305162
transform -1 0 6530 0 -1 10330
box -12 -8 112 252
use INVX1  _2720_
timestamp 1728304789
transform 1 0 4750 0 -1 8890
box -12 -8 72 252
use OAI21X1  _2721_
timestamp 1728305162
transform 1 0 5010 0 1 8890
box -12 -8 112 252
use AOI21X1  _2722_
timestamp 1728304211
transform 1 0 5270 0 1 8890
box -12 -8 112 252
use OAI21X1  _2723_
timestamp 1728305162
transform -1 0 5590 0 -1 9850
box -12 -8 112 252
use NOR2X1  _2724_
timestamp 1728305106
transform 1 0 6250 0 -1 10810
box -12 -8 92 252
use INVX1  _2725_
timestamp 1728304789
transform 1 0 6490 0 -1 10810
box -12 -8 72 252
use OAI21X1  _2726_
timestamp 1728305162
transform -1 0 6310 0 1 10810
box -12 -8 112 252
use OAI22X1  _2727_
timestamp 1728305200
transform 1 0 5950 0 1 10810
box -12 -8 132 252
use INVX1  _2728_
timestamp 1728304789
transform -1 0 4450 0 1 7930
box -12 -8 72 252
use OAI21X1  _2729_
timestamp 1728305162
transform -1 0 4370 0 1 8410
box -12 -8 112 252
use AOI21X1  _2730_
timestamp 1728304211
transform -1 0 5410 0 1 8410
box -12 -8 112 252
use OAI21X1  _2731_
timestamp 1728305162
transform -1 0 5510 0 -1 9370
box -12 -8 112 252
use AOI21X1  _2732_
timestamp 1728304211
transform -1 0 5830 0 -1 10810
box -12 -8 112 252
use NAND3X1  _2733_
timestamp 1728305047
transform -1 0 6090 0 -1 10810
box -12 -8 112 252
use NAND2X1  _2734_
timestamp 1728304996
transform -1 0 5370 0 1 10330
box -12 -8 92 252
use OAI22X1  _2735_
timestamp 1728305200
transform 1 0 5530 0 1 10330
box -12 -8 132 252
use AOI21X1  _2736_
timestamp 1728304211
transform -1 0 8510 0 1 6490
box -12 -8 112 252
use OAI21X1  _2737_
timestamp 1728305162
transform 1 0 3850 0 -1 9370
box -12 -8 112 252
use NAND2X1  _2738_
timestamp 1728304996
transform 1 0 4030 0 1 8890
box -12 -8 92 252
use NAND2X1  _2739_
timestamp 1728304996
transform -1 0 3890 0 -1 8890
box -12 -8 92 252
use NAND3X1  _2740_
timestamp 1728305047
transform -1 0 3870 0 1 8890
box -12 -8 112 252
use NOR3X1  _2741_
timestamp 1728303224
transform -1 0 4290 0 -1 9370
box -12 -8 192 252
use OAI21X1  _2742_
timestamp 1728305162
transform -1 0 4330 0 -1 10810
box -12 -8 112 252
use INVX1  _2743_
timestamp 1728304789
transform 1 0 5010 0 -1 10810
box -12 -8 72 252
use AND2X2  _2744_
timestamp 1728304163
transform 1 0 4730 0 1 10810
box -12 -8 112 252
use OAI21X1  _2745_
timestamp 1728305162
transform 1 0 5230 0 -1 10810
box -12 -8 112 252
use OAI22X1  _2746_
timestamp 1728305200
transform 1 0 4730 0 -1 10810
box -12 -8 132 252
use OAI21X1  _2747_
timestamp 1728305162
transform 1 0 5630 0 1 9850
box -12 -8 112 252
use AOI21X1  _2748_
timestamp 1728304211
transform -1 0 5130 0 1 9370
box -12 -8 112 252
use AOI21X1  _2749_
timestamp 1728304211
transform -1 0 5490 0 1 9850
box -12 -8 112 252
use NAND3X1  _2750_
timestamp 1728305047
transform -1 0 5570 0 -1 10810
box -12 -8 112 252
use NOR2X1  _2751_
timestamp 1728305106
transform 1 0 4490 0 -1 10810
box -12 -8 92 252
use NOR2X1  _2752_
timestamp 1728305106
transform 1 0 3970 0 -1 9850
box -12 -8 92 252
use INVX1  _2753_
timestamp 1728304789
transform -1 0 3570 0 -1 9850
box -12 -8 72 252
use AOI22X1  _2754_
timestamp 1728304278
transform -1 0 3210 0 -1 9370
box -14 -8 132 252
use NAND3X1  _2755_
timestamp 1728305047
transform 1 0 3350 0 -1 9370
box -12 -8 112 252
use AOI21X1  _2756_
timestamp 1728304211
transform -1 0 3830 0 -1 9850
box -12 -8 112 252
use OAI21X1  _2757_
timestamp 1728305162
transform -1 0 3830 0 1 9850
box -12 -8 112 252
use AOI21X1  _2758_
timestamp 1728304211
transform -1 0 3830 0 -1 10810
box -12 -8 112 252
use NOR2X1  _2759_
timestamp 1728305106
transform -1 0 3690 0 -1 9370
box -12 -8 92 252
use OAI21X1  _2760_
timestamp 1728305162
transform -1 0 3730 0 1 9370
box -12 -8 112 252
use NOR2X1  _2761_
timestamp 1728305106
transform -1 0 3870 0 -1 10330
box -12 -8 92 252
use OAI21X1  _2762_
timestamp 1728305162
transform -1 0 3650 0 1 10330
box -12 -8 112 252
use OAI21X1  _2763_
timestamp 1728305162
transform 1 0 3110 0 1 10810
box -12 -8 112 252
use OAI22X1  _2764_
timestamp 1728305200
transform 1 0 3410 0 -1 11290
box -12 -8 132 252
use NOR2X1  _2765_
timestamp 1728305106
transform -1 0 2770 0 -1 10810
box -12 -8 92 252
use INVX1  _2766_
timestamp 1728304789
transform 1 0 3810 0 1 7450
box -12 -8 72 252
use OAI21X1  _2767_
timestamp 1728305162
transform -1 0 4590 0 -1 8890
box -12 -8 112 252
use AOI21X1  _2768_
timestamp 1728304211
transform 1 0 4570 0 1 9370
box -12 -8 112 252
use OAI21X1  _2769_
timestamp 1728305162
transform 1 0 5250 0 -1 9850
box -12 -8 112 252
use AOI22X1  _2770_
timestamp 1728304278
transform -1 0 4850 0 -1 9850
box -14 -8 132 252
use AND2X2  _2771_
timestamp 1728304163
transform -1 0 5090 0 -1 9850
box -12 -8 112 252
use AND2X2  _2772_
timestamp 1728304163
transform -1 0 5090 0 -1 10330
box -12 -8 112 252
use MUX2X1  _2773_
timestamp 1728304958
transform 1 0 2750 0 1 10330
box -12 -8 131 252
use NOR2X1  _2774_
timestamp 1728305106
transform -1 0 2690 0 1 10810
box -12 -8 92 252
use NAND3X1  _2775_
timestamp 1728305047
transform 1 0 3990 0 -1 10810
box -12 -8 112 252
use NAND2X1  _2776_
timestamp 1728304996
transform 1 0 4490 0 -1 10330
box -12 -8 92 252
use NAND2X1  _2777_
timestamp 1728304996
transform 1 0 5250 0 -1 10330
box -12 -8 92 252
use OAI21X1  _2778_
timestamp 1728305162
transform -1 0 4830 0 -1 10330
box -12 -8 112 252
use OAI21X1  _2779_
timestamp 1728305162
transform 1 0 4050 0 1 10810
box -12 -8 112 252
use OAI22X1  _2780_
timestamp 1728305200
transform 1 0 2850 0 1 10810
box -12 -8 132 252
use OAI21X1  _2781_
timestamp 1728305162
transform -1 0 4130 0 -1 8890
box -12 -8 112 252
use AOI21X1  _2782_
timestamp 1728304211
transform -1 0 2950 0 -1 8890
box -12 -8 112 252
use NAND3X1  _2783_
timestamp 1728305047
transform 1 0 2570 0 1 8890
box -12 -8 112 252
use INVX1  _2784_
timestamp 1728304789
transform 1 0 630 0 -1 9370
box -12 -8 72 252
use MUX2X1  _2785_
timestamp 1728304958
transform -1 0 2450 0 -1 9370
box -12 -8 131 252
use AOI21X1  _2786_
timestamp 1728304211
transform 1 0 2590 0 -1 9370
box -12 -8 112 252
use OAI21X1  _2787_
timestamp 1728305162
transform -1 0 3110 0 -1 10330
box -12 -8 112 252
use AOI21X1  _2788_
timestamp 1728304211
transform -1 0 2610 0 1 10330
box -12 -8 112 252
use NAND2X1  _2789_
timestamp 1728304996
transform -1 0 3870 0 1 10330
box -12 -8 92 252
use NAND2X1  _2790_
timestamp 1728304996
transform 1 0 3310 0 1 10330
box -12 -8 92 252
use AOI22X1  _2791_
timestamp 1728304278
transform -1 0 3150 0 1 10330
box -14 -8 132 252
use NAND3X1  _2792_
timestamp 1728305047
transform -1 0 3010 0 -1 10810
box -12 -8 112 252
use OAI21X1  _2793_
timestamp 1728305162
transform -1 0 2450 0 1 10810
box -12 -8 112 252
use OAI22X1  _2794_
timestamp 1728305200
transform 1 0 2230 0 1 10330
box -12 -8 132 252
use NAND2X1  _2795_
timestamp 1728304996
transform 1 0 890 0 -1 10810
box -12 -8 92 252
use OAI21X1  _2796_
timestamp 1728305162
transform 1 0 1830 0 -1 9370
box -12 -8 112 252
use AOI21X1  _2797_
timestamp 1728304211
transform -1 0 2170 0 1 8890
box -12 -8 112 252
use OAI21X1  _2798_
timestamp 1728305162
transform 1 0 1330 0 -1 9370
box -12 -8 112 252
use NOR2X1  _2799_
timestamp 1728305106
transform -1 0 1670 0 -1 9370
box -12 -8 92 252
use OAI21X1  _2800_
timestamp 1728305162
transform -1 0 1930 0 -1 9850
box -12 -8 112 252
use NOR2X1  _2801_
timestamp 1728305106
transform 1 0 1830 0 -1 10330
box -12 -8 92 252
use NOR2X1  _2802_
timestamp 1728305106
transform 1 0 1890 0 -1 10810
box -12 -8 92 252
use NOR3X1  _2803_
timestamp 1728303224
transform 1 0 3390 0 -1 10810
box -12 -8 192 252
use NAND2X1  _2804_
timestamp 1728304996
transform -1 0 610 0 -1 11290
box -12 -8 92 252
use NOR2X1  _2805_
timestamp 1728305106
transform 1 0 7070 0 1 10330
box -12 -8 92 252
use NAND2X1  _2806_
timestamp 1728304996
transform -1 0 5570 0 -1 10330
box -12 -8 92 252
use NOR2X1  _2807_
timestamp 1728305106
transform -1 0 5150 0 1 10330
box -12 -8 92 252
use NAND2X1  _2808_
timestamp 1728304996
transform 1 0 4030 0 -1 10330
box -12 -8 92 252
use OAI21X1  _2809_
timestamp 1728305162
transform -1 0 4570 0 -1 9850
box -12 -8 112 252
use INVX1  _2810_
timestamp 1728304789
transform -1 0 4870 0 1 9370
box -12 -8 72 252
use OAI21X1  _2811_
timestamp 1728305162
transform -1 0 4790 0 -1 9370
box -12 -8 112 252
use AOI21X1  _2812_
timestamp 1728304211
transform 1 0 4330 0 1 9370
box -12 -8 112 252
use AOI21X1  _2813_
timestamp 1728304211
transform 1 0 4070 0 1 9370
box -12 -8 112 252
use NAND3X1  _2814_
timestamp 1728305047
transform 1 0 4210 0 -1 9850
box -12 -8 112 252
use OAI21X1  _2815_
timestamp 1728305162
transform -1 0 4350 0 -1 10330
box -12 -8 112 252
use AND2X2  _2816_
timestamp 1728304163
transform 1 0 2590 0 -1 8890
box -12 -8 112 252
use NAND2X1  _2817_
timestamp 1728304996
transform -1 0 2930 0 -1 9370
box -12 -8 92 252
use NAND3X1  _2818_
timestamp 1728305047
transform 1 0 2810 0 1 8890
box -12 -8 112 252
use NOR2X1  _2819_
timestamp 1728305106
transform 1 0 3270 0 -1 10330
box -12 -8 92 252
use OAI22X1  _2820_
timestamp 1728305200
transform 1 0 3510 0 -1 10330
box -12 -8 132 252
use NOR3X1  _2821_
timestamp 1728303224
transform -1 0 4190 0 1 10330
box -12 -8 192 252
use NAND3X1  _2822_
timestamp 1728305047
transform -1 0 4930 0 1 10330
box -12 -8 112 252
use OAI21X1  _2823_
timestamp 1728305162
transform -1 0 1890 0 1 10330
box -12 -8 112 252
use AND2X2  _2824_
timestamp 1728304163
transform 1 0 650 0 1 10810
box -12 -8 112 252
use OAI21X1  _2825_
timestamp 1728305162
transform 1 0 630 0 -1 10810
box -12 -8 112 252
use INVX1  _2826_
timestamp 1728304789
transform -1 0 810 0 -1 11290
box -12 -8 72 252
use OAI21X1  _2827_
timestamp 1728305162
transform 1 0 1830 0 -1 8890
box -12 -8 112 252
use AOI21X1  _2828_
timestamp 1728304211
transform -1 0 2190 0 -1 8890
box -12 -8 112 252
use OAI21X1  _2829_
timestamp 1728305162
transform 1 0 1330 0 -1 8890
box -12 -8 112 252
use NOR2X1  _2830_
timestamp 1728305106
transform -1 0 1670 0 -1 8890
box -12 -8 92 252
use OAI21X1  _2831_
timestamp 1728305162
transform -1 0 1690 0 1 8890
box -12 -8 112 252
use NOR2X1  _2832_
timestamp 1728305106
transform 1 0 2130 0 -1 10810
box -12 -8 92 252
use NOR2X1  _2833_
timestamp 1728305106
transform -1 0 1210 0 1 10810
box -12 -8 92 252
use AOI21X1  _2834_
timestamp 1728304211
transform 1 0 950 0 -1 11290
box -12 -8 112 252
use INVX1  _2835_
timestamp 1728304789
transform 1 0 1210 0 -1 11290
box -12 -8 72 252
use NOR3X1  _2836_
timestamp 1728303224
transform 1 0 1410 0 -1 11290
box -12 -8 192 252
use OAI21X1  _2837_
timestamp 1728305162
transform 1 0 1750 0 -1 11290
box -12 -8 112 252
use OAI21X1  _2838_
timestamp 1728305162
transform -1 0 1710 0 1 10810
box -12 -8 112 252
use NOR2X1  _2839_
timestamp 1728305106
transform 1 0 890 0 1 10810
box -12 -8 92 252
use NOR2X1  _2840_
timestamp 1728305106
transform 1 0 1350 0 1 9850
box -12 -8 92 252
use NOR2X1  _2841_
timestamp 1728305106
transform 1 0 2150 0 1 8410
box -12 -8 92 252
use AOI22X1  _2842_
timestamp 1728304278
transform -1 0 1890 0 -1 8410
box -14 -8 132 252
use AND2X2  _2843_
timestamp 1728304163
transform -1 0 1990 0 1 8410
box -12 -8 112 252
use OAI21X1  _2844_
timestamp 1728305162
transform -1 0 1730 0 1 8410
box -12 -8 112 252
use NOR2X1  _2845_
timestamp 1728305106
transform -1 0 1670 0 1 9850
box -12 -8 92 252
use NAND3X1  _2846_
timestamp 1728305047
transform 1 0 1390 0 -1 10810
box -12 -8 112 252
use OAI21X1  _2847_
timestamp 1728305162
transform -1 0 1450 0 1 10810
box -12 -8 112 252
use INVX1  _2848_
timestamp 1728304789
transform -1 0 1410 0 1 10330
box -12 -8 72 252
use OAI21X1  _2849_
timestamp 1728305162
transform -1 0 1750 0 -1 10810
box -12 -8 112 252
use NAND3X1  _2850_
timestamp 1728305047
transform -1 0 1650 0 1 10330
box -12 -8 112 252
use NAND2X1  _2851_
timestamp 1728304996
transform -1 0 1190 0 1 9850
box -12 -8 92 252
use AND2X2  _2852_
timestamp 1728304163
transform -1 0 1250 0 -1 10330
box -12 -8 112 252
use NOR3X1  _2853_
timestamp 1728303224
transform -1 0 2550 0 -1 10810
box -12 -8 192 252
use NOR2X1  _2854_
timestamp 1728305106
transform 1 0 870 0 1 9850
box -12 -8 92 252
use NOR2X1  _2855_
timestamp 1728305106
transform 1 0 2530 0 -1 7930
box -12 -8 92 252
use AOI22X1  _2856_
timestamp 1728304278
transform -1 0 2170 0 -1 8410
box -14 -8 132 252
use AND2X2  _2857_
timestamp 1728304163
transform -1 0 2550 0 1 7930
box -12 -8 112 252
use OAI21X1  _2858_
timestamp 1728305162
transform -1 0 2430 0 -1 8890
box -12 -8 112 252
use NOR2X1  _2859_
timestamp 1728305106
transform -1 0 1010 0 -1 10330
box -12 -8 92 252
use NAND3X1  _2860_
timestamp 1728305047
transform 1 0 610 0 1 10330
box -12 -8 112 252
use INVX1  _2861_
timestamp 1728304789
transform -1 0 230 0 1 10330
box -12 -8 72 252
use NAND3X1  _2862_
timestamp 1728305047
transform -1 0 1230 0 -1 10810
box -12 -8 112 252
use AOI21X1  _2863_
timestamp 1728304211
transform 1 0 370 0 1 10330
box -12 -8 112 252
use AOI22X1  _2864_
timestamp 1728304278
transform -1 0 530 0 -1 10330
box -14 -8 132 252
use INVX1  _2865_
timestamp 1728304789
transform 1 0 4530 0 -1 6010
box -12 -8 72 252
use NAND3X1  _2866_
timestamp 1728305047
transform 1 0 4570 0 1 6010
box -12 -8 112 252
use OAI21X1  _2867_
timestamp 1728305162
transform 1 0 5670 0 1 6010
box -12 -8 112 252
use NAND2X1  _2868_
timestamp 1728304996
transform -1 0 3090 0 -1 3130
box -12 -8 92 252
use OAI21X1  _2869_
timestamp 1728305162
transform -1 0 3410 0 1 3130
box -12 -8 112 252
use NAND2X1  _2870_
timestamp 1728304996
transform -1 0 2450 0 1 3610
box -12 -8 92 252
use OAI21X1  _2871_
timestamp 1728305162
transform 1 0 2390 0 -1 3610
box -12 -8 112 252
use NAND2X1  _2872_
timestamp 1728304996
transform -1 0 4750 0 1 4090
box -12 -8 92 252
use OAI21X1  _2873_
timestamp 1728305162
transform 1 0 4410 0 1 4090
box -12 -8 112 252
use INVX1  _2874_
timestamp 1728304789
transform -1 0 4270 0 1 2650
box -12 -8 72 252
use INVX2  _2875_
timestamp 1728304826
transform -1 0 1830 0 -1 250
box -12 -8 72 252
use NOR2X1  _2876_
timestamp 1728305106
transform -1 0 970 0 1 1690
box -12 -8 92 252
use NAND2X1  _2877_
timestamp 1728304996
transform -1 0 3650 0 -1 2170
box -12 -8 92 252
use OAI21X1  _2878_
timestamp 1728305162
transform -1 0 4110 0 -1 2650
box -12 -8 112 252
use INVX1  _2879_
timestamp 1728304789
transform -1 0 1390 0 -1 2650
box -12 -8 72 252
use NOR2X1  _2880_
timestamp 1728305106
transform 1 0 1550 0 -1 2650
box -12 -8 92 252
use NAND2X1  _2881_
timestamp 1728304996
transform -1 0 1910 0 -1 3130
box -12 -8 92 252
use OAI22X1  _2882_
timestamp 1728305200
transform -1 0 2650 0 -1 3130
box -12 -8 132 252
use OAI21X1  _2883_
timestamp 1728305162
transform 1 0 4550 0 -1 2650
box -12 -8 112 252
use NAND2X1  _2884_
timestamp 1728304996
transform 1 0 4250 0 -1 1690
box -12 -8 92 252
use OR2X2  _2885_
timestamp 1728305284
transform 1 0 3210 0 1 1690
box -12 -8 112 252
use OAI21X1  _2886_
timestamp 1728305162
transform 1 0 4750 0 -1 2170
box -12 -8 112 252
use INVX1  _2887_
timestamp 1728304789
transform 1 0 5230 0 1 1690
box -12 -8 72 252
use NOR2X1  _2888_
timestamp 1728305106
transform 1 0 3490 0 1 2650
box -12 -8 92 252
use NAND2X1  _2889_
timestamp 1728304996
transform 1 0 3690 0 1 1690
box -12 -8 92 252
use OAI22X1  _2890_
timestamp 1728305200
transform -1 0 4590 0 1 1690
box -12 -8 132 252
use OAI21X1  _2891_
timestamp 1728305162
transform -1 0 4310 0 -1 3130
box -12 -8 112 252
use NOR2X1  _2892_
timestamp 1728305106
transform -1 0 2130 0 -1 1210
box -12 -8 92 252
use NAND2X1  _2893_
timestamp 1728304996
transform 1 0 3770 0 1 1210
box -12 -8 92 252
use OAI21X1  _2894_
timestamp 1728305162
transform 1 0 3950 0 1 2170
box -12 -8 112 252
use INVX1  _2895_
timestamp 1728304789
transform 1 0 4550 0 -1 2170
box -12 -8 72 252
use OAI22X1  _2896_
timestamp 1728305200
transform -1 0 4050 0 1 1690
box -12 -8 132 252
use OAI21X1  _2897_
timestamp 1728305162
transform -1 0 6010 0 1 1690
box -12 -8 112 252
use NAND2X1  _2898_
timestamp 1728304996
transform 1 0 5270 0 1 1210
box -12 -8 92 252
use OAI21X1  _2899_
timestamp 1728305162
transform 1 0 5230 0 -1 1690
box -12 -8 112 252
use INVX1  _2900_
timestamp 1728304789
transform 1 0 5470 0 -1 2170
box -12 -8 72 252
use OAI22X1  _2901_
timestamp 1728305200
transform -1 0 5070 0 -1 1690
box -12 -8 132 252
use OAI21X1  _2902_
timestamp 1728305162
transform -1 0 1690 0 -1 3130
box -12 -8 112 252
use NOR2X1  _2903_
timestamp 1728305106
transform 1 0 2290 0 -1 1210
box -12 -8 92 252
use NAND2X1  _2904_
timestamp 1728304996
transform 1 0 2550 0 1 730
box -12 -8 92 252
use NOR2X1  _2905_
timestamp 1728305106
transform 1 0 1330 0 1 1690
box -12 -8 92 252
use INVX1  _2906_
timestamp 1728304789
transform 1 0 1130 0 1 1690
box -12 -8 72 252
use OAI21X1  _2907_
timestamp 1728305162
transform 1 0 1330 0 1 2650
box -12 -8 112 252
use NAND3X1  _2908_
timestamp 1728305047
transform -1 0 1710 0 1 1210
box -12 -8 112 252
use NAND3X1  _2909_
timestamp 1728305047
transform -1 0 1950 0 -1 1690
box -12 -8 112 252
use NOR2X1  _2910_
timestamp 1728305106
transform -1 0 1690 0 -1 1690
box -12 -8 92 252
use INVX1  _2911_
timestamp 1728304789
transform -1 0 1690 0 -1 2170
box -12 -8 72 252
use OAI21X1  _2912_
timestamp 1728305162
transform -1 0 2650 0 1 2650
box -12 -8 112 252
use OAI21X1  _2913_
timestamp 1728305162
transform -1 0 1870 0 -1 2650
box -12 -8 112 252
use NOR2X1  _2914_
timestamp 1728305106
transform 1 0 2330 0 -1 1690
box -12 -8 92 252
use NOR2X1  _2915_
timestamp 1728305106
transform 1 0 2090 0 -1 1690
box -12 -8 92 252
use AND2X2  _2916_
timestamp 1728304163
transform 1 0 1790 0 1 1690
box -12 -8 112 252
use OAI21X1  _2917_
timestamp 1728305162
transform -1 0 1950 0 -1 2170
box -12 -8 112 252
use AOI21X1  _2918_
timestamp 1728304211
transform 1 0 1790 0 1 2170
box -12 -8 112 252
use NOR2X1  _2919_
timestamp 1728305106
transform -1 0 2410 0 -1 2170
box -12 -8 92 252
use INVX1  _2920_
timestamp 1728304789
transform -1 0 2110 0 1 2170
box -12 -8 72 252
use NOR2X1  _2921_
timestamp 1728305106
transform -1 0 2170 0 -1 2170
box -12 -8 92 252
use AOI21X1  _2922_
timestamp 1728304211
transform -1 0 2130 0 -1 2650
box -12 -8 112 252
use AOI22X1  _2923_
timestamp 1728304278
transform -1 0 2170 0 -1 3130
box -14 -8 132 252
use NAND2X1  _2924_
timestamp 1728304996
transform -1 0 3110 0 1 1210
box -12 -8 92 252
use NOR2X1  _2925_
timestamp 1728305106
transform 1 0 3530 0 -1 1210
box -12 -8 92 252
use OAI21X1  _2926_
timestamp 1728305162
transform -1 0 2570 0 1 1690
box -12 -8 112 252
use AOI22X1  _2927_
timestamp 1728304278
transform -1 0 2650 0 -1 2650
box -14 -8 132 252
use INVX1  _2928_
timestamp 1728304789
transform 1 0 4690 0 1 2170
box -12 -8 72 252
use AND2X2  _2929_
timestamp 1728304163
transform 1 0 3510 0 1 730
box -12 -8 112 252
use NAND2X1  _2930_
timestamp 1728304996
transform -1 0 2870 0 1 730
box -12 -8 92 252
use NOR2X1  _2931_
timestamp 1728305106
transform -1 0 3090 0 1 730
box -12 -8 92 252
use AOI22X1  _2932_
timestamp 1728304278
transform 1 0 3250 0 1 730
box -14 -8 132 252
use NAND2X1  _2933_
timestamp 1728304996
transform -1 0 2870 0 -1 1210
box -12 -8 92 252
use OAI21X1  _2934_
timestamp 1728305162
transform 1 0 3010 0 -1 1210
box -12 -8 112 252
use INVX2  _2935_
timestamp 1728304826
transform -1 0 1450 0 1 730
box -12 -8 72 252
use NAND2X1  _2936_
timestamp 1728304996
transform -1 0 990 0 -1 1210
box -12 -8 92 252
use OR2X2  _2937_
timestamp 1728305284
transform 1 0 670 0 -1 730
box -12 -8 112 252
use NAND2X1  _2938_
timestamp 1728304996
transform 1 0 1830 0 -1 1210
box -12 -8 92 252
use OAI21X1  _2939_
timestamp 1728305162
transform -1 0 1670 0 -1 1210
box -12 -8 112 252
use AOI21X1  _2940_
timestamp 1728304211
transform 1 0 3270 0 -1 1210
box -12 -8 112 252
use AND2X2  _2941_
timestamp 1728304163
transform 1 0 3270 0 1 1210
box -12 -8 112 252
use AOI21X1  _2942_
timestamp 1728304211
transform -1 0 3550 0 1 1690
box -12 -8 112 252
use AND2X2  _2943_
timestamp 1728304163
transform -1 0 3410 0 -1 2170
box -12 -8 112 252
use AOI22X1  _2944_
timestamp 1728304278
transform -1 0 3910 0 -1 2170
box -14 -8 132 252
use INVX1  _2945_
timestamp 1728304789
transform 1 0 3270 0 1 4090
box -12 -8 72 252
use OAI21X1  _2946_
timestamp 1728305162
transform 1 0 3710 0 1 4090
box -12 -8 112 252
use OAI21X1  _2947_
timestamp 1728305162
transform 1 0 3270 0 -1 2650
box -12 -8 112 252
use OAI22X1  _2948_
timestamp 1728305200
transform -1 0 4390 0 -1 2650
box -12 -8 132 252
use AOI21X1  _2949_
timestamp 1728304211
transform 1 0 3250 0 -1 3130
box -12 -8 112 252
use NOR2X1  _2950_
timestamp 1728305106
transform 1 0 2550 0 -1 2170
box -12 -8 92 252
use AOI22X1  _2951_
timestamp 1728304278
transform -1 0 2910 0 -1 2170
box -14 -8 132 252
use OAI21X1  _2952_
timestamp 1728305162
transform -1 0 3150 0 -1 2170
box -12 -8 112 252
use NAND2X1  _2953_
timestamp 1728304996
transform -1 0 2350 0 1 2170
box -12 -8 92 252
use OAI22X1  _2954_
timestamp 1728305200
transform -1 0 2630 0 1 2170
box -12 -8 132 252
use OAI21X1  _2955_
timestamp 1728305162
transform 1 0 3090 0 1 3610
box -12 -8 112 252
use INVX1  _2956_
timestamp 1728304789
transform 1 0 3350 0 1 3610
box -12 -8 72 252
use NAND2X1  _2957_
timestamp 1728304996
transform 1 0 3850 0 1 3610
box -12 -8 92 252
use NAND3X1  _2958_
timestamp 1728305047
transform 1 0 2270 0 -1 2650
box -12 -8 112 252
use OAI22X1  _2959_
timestamp 1728305200
transform 1 0 3570 0 1 3610
box -12 -8 132 252
use OAI21X1  _2960_
timestamp 1728305162
transform 1 0 3670 0 -1 4090
box -12 -8 112 252
use INVX1  _2961_
timestamp 1728304789
transform 1 0 2810 0 1 1210
box -12 -8 72 252
use NAND3X1  _2962_
timestamp 1728305047
transform 1 0 2550 0 1 1210
box -12 -8 112 252
use AOI22X1  _2963_
timestamp 1728304278
transform 1 0 3050 0 -1 1690
box -14 -8 132 252
use OAI21X1  _2964_
timestamp 1728305162
transform 1 0 2810 0 -1 1690
box -12 -8 112 252
use OAI21X1  _2965_
timestamp 1728305162
transform -1 0 5950 0 1 2170
box -12 -8 112 252
use OAI21X1  _2966_
timestamp 1728305162
transform 1 0 4210 0 1 1690
box -12 -8 112 252
use NAND2X1  _2967_
timestamp 1728304996
transform -1 0 4750 0 -1 730
box -12 -8 92 252
use OAI22X1  _2968_
timestamp 1728305200
transform -1 0 5010 0 -1 730
box -12 -8 132 252
use INVX1  _2969_
timestamp 1728304789
transform -1 0 1470 0 -1 2170
box -12 -8 72 252
use OAI21X1  _2970_
timestamp 1728305162
transform -1 0 1690 0 1 2650
box -12 -8 112 252
use NOR2X1  _2971_
timestamp 1728305106
transform -1 0 1670 0 1 730
box -12 -8 92 252
use OAI21X1  _2972_
timestamp 1728305162
transform -1 0 1450 0 1 2170
box -12 -8 112 252
use OAI21X1  _2973_
timestamp 1728305162
transform -1 0 1190 0 1 2170
box -12 -8 112 252
use INVX1  _2974_
timestamp 1728304789
transform -1 0 1910 0 -1 730
box -12 -8 72 252
use NOR2X1  _2975_
timestamp 1728305106
transform -1 0 2150 0 -1 730
box -12 -8 92 252
use AOI21X1  _2976_
timestamp 1728304211
transform 1 0 3950 0 -1 730
box -12 -8 112 252
use AOI22X1  _2977_
timestamp 1728304278
transform -1 0 4630 0 1 1210
box -14 -8 132 252
use OAI21X1  _2978_
timestamp 1728305162
transform 1 0 4250 0 1 1210
box -12 -8 112 252
use NOR2X1  _2979_
timestamp 1728305106
transform 1 0 1610 0 -1 730
box -12 -8 92 252
use INVX1  _2980_
timestamp 1728304789
transform -1 0 1150 0 -1 250
box -12 -8 72 252
use OAI21X1  _2981_
timestamp 1728305162
transform -1 0 930 0 -1 250
box -12 -8 112 252
use NAND2X1  _2982_
timestamp 1728304996
transform 1 0 2310 0 -1 730
box -12 -8 92 252
use NAND2X1  _2983_
timestamp 1728304996
transform -1 0 690 0 -1 250
box -12 -8 92 252
use NOR2X1  _2984_
timestamp 1728305106
transform -1 0 450 0 -1 250
box -12 -8 92 252
use INVX1  _2985_
timestamp 1728304789
transform -1 0 230 0 -1 250
box -12 -8 72 252
use OAI21X1  _2986_
timestamp 1728305162
transform -1 0 530 0 1 250
box -12 -8 112 252
use AOI21X1  _2987_
timestamp 1728304211
transform -1 0 770 0 1 250
box -12 -8 112 252
use OAI21X1  _2988_
timestamp 1728305162
transform -1 0 750 0 1 1210
box -12 -8 112 252
use NAND2X1  _2989_
timestamp 1728304996
transform 1 0 410 0 1 1210
box -12 -8 92 252
use OAI21X1  _2990_
timestamp 1728305162
transform 1 0 170 0 1 1210
box -12 -8 112 252
use OAI21X1  _2991_
timestamp 1728305162
transform -1 0 530 0 -1 1210
box -12 -8 112 252
use NAND2X1  _2992_
timestamp 1728304996
transform -1 0 2150 0 1 1210
box -12 -8 92 252
use OAI21X1  _2993_
timestamp 1728305162
transform -1 0 1230 0 1 730
box -12 -8 112 252
use OAI21X1  _2994_
timestamp 1728305162
transform -1 0 970 0 1 730
box -12 -8 112 252
use NOR2X1  _2995_
timestamp 1728305106
transform 1 0 690 0 -1 1210
box -12 -8 92 252
use AOI22X1  _2996_
timestamp 1728304278
transform -1 0 730 0 -1 1690
box -14 -8 132 252
use OAI21X1  _2997_
timestamp 1728305162
transform -1 0 1010 0 -1 730
box -12 -8 112 252
use OAI21X1  _2998_
timestamp 1728305162
transform -1 0 270 0 1 250
box -12 -8 112 252
use OAI21X1  _2999_
timestamp 1728305162
transform -1 0 510 0 -1 730
box -12 -8 112 252
use OAI21X1  _3000_
timestamp 1728305162
transform -1 0 250 0 -1 730
box -12 -8 112 252
use OAI21X1  _3001_
timestamp 1728305162
transform -1 0 270 0 -1 1210
box -12 -8 112 252
use OAI21X1  _3002_
timestamp 1728305162
transform -1 0 730 0 1 730
box -12 -8 112 252
use OAI21X1  _3003_
timestamp 1728305162
transform -1 0 270 0 1 730
box -12 -8 112 252
use INVX1  _3004_
timestamp 1728304789
transform -1 0 970 0 1 1210
box -12 -8 72 252
use AOI22X1  _3005_
timestamp 1728304278
transform 1 0 870 0 -1 1690
box -14 -8 132 252
use NAND2X1  _3006_
timestamp 1728304996
transform -1 0 250 0 -1 1690
box -12 -8 92 252
use INVX1  _3007_
timestamp 1728304789
transform 1 0 1890 0 1 3610
box -12 -8 72 252
use OAI22X1  _3008_
timestamp 1728305200
transform -1 0 1230 0 1 1210
box -12 -8 132 252
use NAND2X1  _3009_
timestamp 1728304996
transform -1 0 1470 0 -1 1690
box -12 -8 92 252
use OAI21X1  _3010_
timestamp 1728305162
transform -1 0 1470 0 1 1210
box -12 -8 112 252
use NOR2X1  _3011_
timestamp 1728305106
transform -1 0 1230 0 -1 1690
box -12 -8 92 252
use NOR2X1  _3012_
timestamp 1728305106
transform -1 0 1610 0 -1 250
box -12 -8 92 252
use NAND2X1  _3013_
timestamp 1728304996
transform -1 0 1370 0 -1 250
box -12 -8 92 252
use INVX1  _3014_
timestamp 1728304789
transform 1 0 1130 0 1 250
box -12 -8 72 252
use NAND3X1  _3015_
timestamp 1728305047
transform -1 0 1690 0 1 250
box -12 -8 112 252
use OAI21X1  _3016_
timestamp 1728305162
transform -1 0 1470 0 -1 730
box -12 -8 112 252
use NAND3X1  _3017_
timestamp 1728305047
transform -1 0 1450 0 1 250
box -12 -8 112 252
use NOR2X1  _3018_
timestamp 1728305106
transform 1 0 1130 0 -1 1210
box -12 -8 92 252
use AOI22X1  _3019_
timestamp 1728304278
transform -1 0 1250 0 -1 2170
box -14 -8 132 252
use AND2X2  _3020_
timestamp 1728304163
transform -1 0 3870 0 1 8410
box -12 -8 112 252
use OAI21X1  _3021_
timestamp 1728305162
transform -1 0 6110 0 1 4090
box -12 -8 112 252
use NOR2X1  _3022_
timestamp 1728305106
transform 1 0 2890 0 -1 5050
box -12 -8 92 252
use INVX2  _3023_
timestamp 1728304826
transform 1 0 2890 0 1 5050
box -12 -8 72 252
use OAI21X1  _3024_
timestamp 1728305162
transform 1 0 3890 0 -1 5530
box -12 -8 112 252
use OAI21X1  _3025_
timestamp 1728305162
transform -1 0 4390 0 1 5530
box -12 -8 112 252
use OAI21X1  _3026_
timestamp 1728305162
transform -1 0 3230 0 -1 5530
box -12 -8 112 252
use OAI21X1  _3027_
timestamp 1728305162
transform -1 0 3650 0 1 5530
box -12 -8 112 252
use OAI21X1  _3028_
timestamp 1728305162
transform -1 0 4170 0 -1 5050
box -12 -8 112 252
use OAI21X1  _3029_
timestamp 1728305162
transform -1 0 4650 0 -1 5050
box -12 -8 112 252
use OAI21X1  _3030_
timestamp 1728305162
transform 1 0 3570 0 1 4570
box -12 -8 112 252
use OAI21X1  _3031_
timestamp 1728305162
transform -1 0 3910 0 1 4570
box -12 -8 112 252
use OAI21X1  _3032_
timestamp 1728305162
transform -1 0 2730 0 -1 5050
box -12 -8 112 252
use OAI21X1  _3033_
timestamp 1728305162
transform -1 0 2750 0 1 5050
box -12 -8 112 252
use OAI21X1  _3034_
timestamp 1728305162
transform 1 0 2790 0 1 5530
box -12 -8 112 252
use OAI21X1  _3035_
timestamp 1728305162
transform -1 0 3150 0 1 5530
box -12 -8 112 252
use OAI21X1  _3036_
timestamp 1728305162
transform 1 0 3390 0 -1 5530
box -12 -8 112 252
use OAI21X1  _3037_
timestamp 1728305162
transform -1 0 3890 0 1 5530
box -12 -8 112 252
use OAI21X1  _3038_
timestamp 1728305162
transform -1 0 3470 0 -1 5050
box -12 -8 112 252
use OAI21X1  _3039_
timestamp 1728305162
transform 1 0 3110 0 -1 5050
box -12 -8 112 252
use OAI21X1  _3040_
timestamp 1728305162
transform 1 0 2270 0 1 4090
box -12 -8 112 252
use INVX1  _3041_
timestamp 1728304789
transform 1 0 2810 0 -1 3130
box -12 -8 72 252
use OAI21X1  _3042_
timestamp 1728305162
transform 1 0 7550 0 -1 4090
box -12 -8 112 252
use INVX1  _3043_
timestamp 1728304789
transform 1 0 6410 0 -1 4090
box -12 -8 72 252
use OAI21X1  _3044_
timestamp 1728305162
transform 1 0 5410 0 -1 4090
box -12 -8 112 252
use INVX1  _3045_
timestamp 1728304789
transform 1 0 5850 0 -1 4570
box -12 -8 72 252
use NOR2X1  _3046_
timestamp 1728305106
transform 1 0 5570 0 1 4090
box -12 -8 92 252
use INVX1  _3047_
timestamp 1728304789
transform 1 0 4890 0 1 4090
box -12 -8 72 252
use NOR2X1  _3048_
timestamp 1728305106
transform 1 0 5250 0 1 4570
box -12 -8 92 252
use AOI21X1  _3049_
timestamp 1728304211
transform 1 0 5950 0 -1 5050
box -12 -8 112 252
use OAI21X1  _3050_
timestamp 1728305162
transform -1 0 7030 0 1 5050
box -12 -8 112 252
use NAND2X1  _3051_
timestamp 1728304996
transform -1 0 6490 0 1 5530
box -12 -8 92 252
use OAI21X1  _3052_
timestamp 1728305162
transform 1 0 6450 0 1 5050
box -12 -8 112 252
use AND2X2  _3053_
timestamp 1728304163
transform 1 0 6210 0 1 5050
box -12 -8 112 252
use OAI21X1  _3054_
timestamp 1728305162
transform 1 0 5950 0 1 5050
box -12 -8 112 252
use OAI21X1  _3055_
timestamp 1728305162
transform -1 0 6110 0 -1 5530
box -12 -8 112 252
use NOR2X1  _3056_
timestamp 1728305106
transform 1 0 4710 0 -1 3130
box -12 -8 92 252
use NAND2X1  _3057_
timestamp 1728304996
transform 1 0 4470 0 -1 3130
box -12 -8 92 252
use OAI21X1  _3058_
timestamp 1728305162
transform -1 0 4650 0 1 3610
box -12 -8 112 252
use NAND2X1  _3059_
timestamp 1728304996
transform 1 0 4410 0 -1 4090
box -12 -8 92 252
use INVX1  _3060_
timestamp 1728304789
transform -1 0 4410 0 1 3130
box -12 -8 72 252
use OAI21X1  _3061_
timestamp 1728305162
transform 1 0 4090 0 1 3610
box -12 -8 112 252
use MUX2X1  _3062_
timestamp 1728304958
transform -1 0 5010 0 -1 4090
box -12 -8 131 252
use OAI21X1  _3063_
timestamp 1728305162
transform 1 0 4630 0 -1 4090
box -12 -8 112 252
use NOR2X1  _3064_
timestamp 1728305106
transform 1 0 6110 0 1 2170
box -12 -8 92 252
use NAND2X1  _3065_
timestamp 1728304996
transform 1 0 5890 0 -1 3130
box -12 -8 92 252
use AOI21X1  _3066_
timestamp 1728304211
transform -1 0 5950 0 1 3610
box -12 -8 112 252
use OAI21X1  _3067_
timestamp 1728305162
transform -1 0 6110 0 -1 3610
box -12 -8 112 252
use NOR2X1  _3068_
timestamp 1728305106
transform -1 0 7110 0 -1 4570
box -12 -8 92 252
use OAI21X1  _3069_
timestamp 1728305162
transform -1 0 6650 0 -1 4570
box -12 -8 112 252
use OAI21X1  _3070_
timestamp 1728305162
transform 1 0 6210 0 -1 5050
box -12 -8 112 252
use NOR2X1  _3071_
timestamp 1728305106
transform -1 0 6530 0 -1 5050
box -12 -8 92 252
use NAND2X1  _3072_
timestamp 1728304996
transform 1 0 6690 0 1 4570
box -12 -8 92 252
use OAI21X1  _3073_
timestamp 1728305162
transform 1 0 6430 0 1 4570
box -12 -8 112 252
use OAI21X1  _3074_
timestamp 1728305162
transform 1 0 510 0 1 3130
box -12 -8 112 252
use NAND2X1  _3075_
timestamp 1728304996
transform -1 0 730 0 -1 4090
box -12 -8 92 252
use NAND2X1  _3076_
timestamp 1728304996
transform -1 0 4410 0 1 3610
box -12 -8 92 252
use AOI21X1  _3077_
timestamp 1728304211
transform 1 0 2110 0 1 3610
box -12 -8 112 252
use AOI21X1  _3078_
timestamp 1728304211
transform -1 0 5690 0 -1 4570
box -12 -8 112 252
use AOI21X1  _3079_
timestamp 1728304211
transform 1 0 5130 0 -1 5530
box -12 -8 112 252
use INVX1  _3080_
timestamp 1728304789
transform 1 0 4350 0 1 6010
box -12 -8 72 252
use AOI21X1  _3081_
timestamp 1728304211
transform 1 0 5970 0 -1 6010
box -12 -8 112 252
use AOI21X1  _3082_
timestamp 1728304211
transform -1 0 7070 0 -1 6010
box -12 -8 112 252
use AOI21X1  _3083_
timestamp 1728304211
transform 1 0 6150 0 1 5530
box -12 -8 112 252
use NAND2X1  _3084_
timestamp 1728304996
transform -1 0 5870 0 -1 5530
box -12 -8 92 252
use OAI21X1  _3085_
timestamp 1728305162
transform -1 0 5190 0 1 5050
box -12 -8 112 252
use INVX1  _3086_
timestamp 1728304789
transform 1 0 5590 0 -1 5530
box -12 -8 72 252
use AOI22X1  _3087_
timestamp 1728304278
transform -1 0 5270 0 -1 4090
box -14 -8 132 252
use MUX2X1  _3088_
timestamp 1728304958
transform -1 0 5830 0 -1 6010
box -12 -8 131 252
use MUX2X1  _3089_
timestamp 1728304958
transform -1 0 5770 0 1 5530
box -12 -8 131 252
use MUX2X1  _3090_
timestamp 1728304958
transform 1 0 4870 0 -1 5530
box -12 -8 131 252
use MUX2X1  _3091_
timestamp 1728304958
transform -1 0 4930 0 1 5050
box -12 -8 131 252
use NOR2X1  _3092_
timestamp 1728305106
transform 1 0 5670 0 -1 2170
box -12 -8 92 252
use NOR2X1  _3093_
timestamp 1728305106
transform -1 0 4150 0 -1 3610
box -12 -8 92 252
use NAND2X1  _3094_
timestamp 1728304996
transform 1 0 4510 0 -1 3610
box -12 -8 92 252
use INVX1  _3095_
timestamp 1728304789
transform 1 0 4830 0 1 3130
box -12 -8 72 252
use NOR2X1  _3096_
timestamp 1728305106
transform 1 0 4810 0 -1 2650
box -12 -8 92 252
use NAND3X1  _3097_
timestamp 1728305047
transform 1 0 5030 0 -1 2650
box -12 -8 112 252
use OAI21X1  _3098_
timestamp 1728305162
transform -1 0 5230 0 1 2650
box -12 -8 112 252
use AOI21X1  _3099_
timestamp 1728304211
transform 1 0 5290 0 -1 2650
box -12 -8 112 252
use NAND2X1  _3100_
timestamp 1728304996
transform -1 0 5730 0 -1 3130
box -12 -8 92 252
use AOI21X1  _3101_
timestamp 1728304211
transform 1 0 5230 0 -1 3610
box -12 -8 112 252
use NAND2X1  _3102_
timestamp 1728304996
transform 1 0 4730 0 -1 3610
box -12 -8 92 252
use OAI21X1  _3103_
timestamp 1728305162
transform 1 0 4970 0 -1 3610
box -12 -8 112 252
use MUX2X1  _3104_
timestamp 1728304958
transform -1 0 5210 0 1 3610
box -12 -8 131 252
use OAI21X1  _3105_
timestamp 1728305162
transform 1 0 5410 0 -1 3130
box -12 -8 112 252
use INVX1  _3106_
timestamp 1728304789
transform 1 0 8610 0 1 10810
box -12 -8 72 252
use NAND2X1  _3107_
timestamp 1728304996
transform 1 0 8370 0 1 10810
box -12 -8 92 252
use OAI21X1  _3108_
timestamp 1728305162
transform 1 0 8110 0 -1 11290
box -12 -8 112 252
use OAI21X1  _3109_
timestamp 1728305162
transform -1 0 8750 0 -1 4570
box -12 -8 112 252
use NAND3X1  _3110_
timestamp 1728305047
transform -1 0 8490 0 -1 4570
box -12 -8 112 252
use NOR2X1  _3111_
timestamp 1728305106
transform 1 0 4610 0 -1 4570
box -12 -8 92 252
use OAI21X1  _3112_
timestamp 1728305162
transform 1 0 4850 0 -1 4570
box -12 -8 112 252
use INVX1  _3113_
timestamp 1728304789
transform -1 0 1390 0 -1 4570
box -12 -8 72 252
use NAND3X1  _3114_
timestamp 1728305047
transform 1 0 870 0 -1 4570
box -12 -8 112 252
use NAND2X1  _3115_
timestamp 1728304996
transform 1 0 4550 0 1 5530
box -12 -8 92 252
use OAI21X1  _3116_
timestamp 1728305162
transform -1 0 4230 0 -1 5530
box -12 -8 112 252
use NAND2X1  _3117_
timestamp 1728304996
transform -1 0 490 0 1 4570
box -12 -8 92 252
use OAI21X1  _3118_
timestamp 1728305162
transform -1 0 250 0 1 4570
box -12 -8 112 252
use AND2X2  _3119_
timestamp 1728304163
transform -1 0 5110 0 -1 6010
box -12 -8 112 252
use NAND2X1  _3120_
timestamp 1728304996
transform 1 0 4530 0 -1 6970
box -12 -8 92 252
use NAND2X1  _3121_
timestamp 1728304996
transform 1 0 5250 0 -1 6010
box -12 -8 92 252
use OAI21X1  _3122_
timestamp 1728305162
transform -1 0 4650 0 1 6490
box -12 -8 112 252
use INVX1  _3123_
timestamp 1728304789
transform -1 0 3850 0 1 6970
box -12 -8 72 252
use NOR2X1  _3124_
timestamp 1728305106
transform -1 0 4110 0 -1 6970
box -12 -8 92 252
use OAI21X1  _3125_
timestamp 1728305162
transform -1 0 3870 0 -1 6970
box -12 -8 112 252
use INVX1  _3126_
timestamp 1728304789
transform 1 0 4790 0 -1 6490
box -12 -8 72 252
use NOR2X1  _3127_
timestamp 1728305106
transform 1 0 4830 0 1 6010
box -12 -8 92 252
use OAI21X1  _3128_
timestamp 1728305162
transform 1 0 4750 0 -1 6010
box -12 -8 112 252
use OAI21X1  _3129_
timestamp 1728305162
transform 1 0 3810 0 -1 6010
box -12 -8 112 252
use INVX1  _3130_
timestamp 1728304789
transform -1 0 1970 0 -1 5050
box -12 -8 72 252
use NAND2X1  _3131_
timestamp 1728304996
transform -1 0 1470 0 1 3610
box -12 -8 92 252
use OAI21X1  _3132_
timestamp 1728305162
transform 1 0 1150 0 1 3610
box -12 -8 112 252
use NOR2X1  _3133_
timestamp 1728305106
transform 1 0 4010 0 1 6970
box -12 -8 92 252
use NOR2X1  _3134_
timestamp 1728305106
transform 1 0 3570 0 1 6970
box -12 -8 92 252
use OR2X2  _3135_
timestamp 1728305284
transform 1 0 3330 0 1 6970
box -12 -8 112 252
use OAI21X1  _3136_
timestamp 1728305162
transform 1 0 3810 0 -1 6490
box -12 -8 112 252
use AOI21X1  _3137_
timestamp 1728304211
transform 1 0 4050 0 -1 6490
box -12 -8 112 252
use AOI21X1  _3138_
timestamp 1728304211
transform -1 0 4190 0 1 6010
box -12 -8 112 252
use NAND2X1  _3139_
timestamp 1728304996
transform 1 0 1150 0 -1 5530
box -12 -8 92 252
use OAI21X1  _3140_
timestamp 1728305162
transform 1 0 910 0 -1 5530
box -12 -8 112 252
use NOR2X1  _3141_
timestamp 1728305106
transform -1 0 4150 0 1 6490
box -12 -8 92 252
use NOR2X1  _3142_
timestamp 1728305106
transform 1 0 3830 0 1 6490
box -12 -8 92 252
use OAI21X1  _3143_
timestamp 1728305162
transform -1 0 4370 0 -1 6970
box -12 -8 112 252
use NAND2X1  _3144_
timestamp 1728304996
transform -1 0 3610 0 -1 6970
box -12 -8 92 252
use NAND2X1  _3145_
timestamp 1728304996
transform 1 0 3310 0 -1 6970
box -12 -8 92 252
use AND2X2  _3146_
timestamp 1728304163
transform -1 0 3470 0 1 6490
box -12 -8 112 252
use NOR2X1  _3147_
timestamp 1728305106
transform 1 0 3610 0 1 6490
box -12 -8 92 252
use NOR2X1  _3148_
timestamp 1728305106
transform -1 0 3650 0 -1 6490
box -12 -8 92 252
use MUX2X1  _3149_
timestamp 1728304958
transform -1 0 3670 0 -1 6010
box -12 -8 131 252
use NAND2X1  _3150_
timestamp 1728304996
transform 1 0 2130 0 -1 5530
box -12 -8 92 252
use OAI21X1  _3151_
timestamp 1728305162
transform -1 0 2470 0 -1 5530
box -12 -8 112 252
use OAI21X1  _3152_
timestamp 1728305162
transform 1 0 7610 0 1 6010
box -12 -8 112 252
use OAI21X1  _3153_
timestamp 1728305162
transform 1 0 4550 0 -1 6490
box -12 -8 112 252
use NAND2X1  _3154_
timestamp 1728304996
transform -1 0 950 0 -1 7930
box -12 -8 92 252
use OAI21X1  _3155_
timestamp 1728305162
transform 1 0 1090 0 -1 7930
box -12 -8 112 252
use NAND2X1  _3156_
timestamp 1728304996
transform 1 0 3070 0 -1 6970
box -12 -8 92 252
use OAI21X1  _3157_
timestamp 1728305162
transform -1 0 2930 0 1 7450
box -12 -8 112 252
use OR2X2  _3158_
timestamp 1728305284
transform 1 0 2050 0 -1 7930
box -12 -8 112 252
use INVX1  _3159_
timestamp 1728304789
transform 1 0 2610 0 1 7450
box -12 -8 72 252
use NOR2X1  _3160_
timestamp 1728305106
transform 1 0 3210 0 -1 7450
box -12 -8 92 252
use OAI21X1  _3161_
timestamp 1728305162
transform -1 0 2850 0 -1 7450
box -12 -8 112 252
use INVX1  _3162_
timestamp 1728304789
transform -1 0 2590 0 -1 7450
box -12 -8 72 252
use NOR2X1  _3163_
timestamp 1728305106
transform -1 0 1690 0 -1 7930
box -12 -8 92 252
use AOI22X1  _3164_
timestamp 1728304278
transform 1 0 1350 0 -1 7930
box -14 -8 132 252
use NAND2X1  _3165_
timestamp 1728304996
transform -1 0 490 0 -1 7930
box -12 -8 92 252
use OAI21X1  _3166_
timestamp 1728305162
transform -1 0 250 0 -1 7930
box -12 -8 112 252
use INVX1  _3167_
timestamp 1728304789
transform 1 0 2150 0 -1 6970
box -12 -8 72 252
use NOR2X1  _3168_
timestamp 1728305106
transform 1 0 2070 0 -1 7450
box -12 -8 92 252
use NOR2X1  _3169_
timestamp 1728305106
transform -1 0 2450 0 1 7450
box -12 -8 92 252
use NOR2X1  _3170_
timestamp 1728305106
transform 1 0 2130 0 1 7450
box -12 -8 92 252
use NAND2X1  _3171_
timestamp 1728304996
transform -1 0 2370 0 -1 7450
box -12 -8 92 252
use INVX1  _3172_
timestamp 1728304789
transform 1 0 1990 0 1 7930
box -12 -8 72 252
use NOR2X1  _3173_
timestamp 1728305106
transform -1 0 1910 0 -1 7930
box -12 -8 92 252
use OAI21X1  _3174_
timestamp 1728305162
transform -1 0 1970 0 1 7450
box -12 -8 112 252
use OAI21X1  _3175_
timestamp 1728305162
transform -1 0 3210 0 1 6490
box -12 -8 112 252
use INVX1  _3176_
timestamp 1728304789
transform -1 0 2950 0 1 6490
box -12 -8 72 252
use NAND2X1  _3177_
timestamp 1728304996
transform 1 0 2370 0 -1 6970
box -12 -8 92 252
use OAI21X1  _3178_
timestamp 1728305162
transform 1 0 2710 0 -1 6490
box -12 -8 112 252
use OAI21X1  _3179_
timestamp 1728305162
transform 1 0 2350 0 1 6970
box -12 -8 112 252
use OAI21X1  _3180_
timestamp 1728305162
transform 1 0 3310 0 -1 6490
box -12 -8 112 252
use NAND2X1  _3181_
timestamp 1728304996
transform -1 0 3070 0 -1 7450
box -12 -8 92 252
use NAND2X1  _3182_
timestamp 1728304996
transform -1 0 3170 0 1 6970
box -12 -8 92 252
use INVX1  _3183_
timestamp 1728304789
transform 1 0 2870 0 1 6970
box -12 -8 72 252
use OAI21X1  _3184_
timestamp 1728305162
transform -1 0 2690 0 -1 6970
box -12 -8 112 252
use AOI21X1  _3185_
timestamp 1728304211
transform -1 0 2710 0 1 6970
box -12 -8 112 252
use AOI21X1  _3186_
timestamp 1728304211
transform 1 0 2110 0 1 6970
box -12 -8 112 252
use NAND2X1  _3187_
timestamp 1728304996
transform -1 0 490 0 -1 7450
box -12 -8 92 252
use OAI21X1  _3188_
timestamp 1728305162
transform -1 0 270 0 -1 7450
box -12 -8 112 252
use NAND2X1  _3189_
timestamp 1728304996
transform 1 0 1110 0 -1 4570
box -12 -8 92 252
use OAI21X1  _3190_
timestamp 1728305162
transform -1 0 1010 0 -1 5050
box -12 -8 112 252
use OAI21X1  _3191_
timestamp 1728305162
transform -1 0 1270 0 -1 5050
box -12 -8 112 252
use OAI21X1  _3192_
timestamp 1728305162
transform 1 0 1790 0 -1 4570
box -12 -8 112 252
use OAI21X1  _3193_
timestamp 1728305162
transform 1 0 1550 0 -1 4570
box -12 -8 112 252
use OAI21X1  _3194_
timestamp 1728305162
transform 1 0 3350 0 1 6010
box -12 -8 112 252
use OAI21X1  _3195_
timestamp 1728305162
transform 1 0 3290 0 -1 6010
box -12 -8 112 252
use OAI21X1  _3196_
timestamp 1728305162
transform 1 0 2050 0 -1 4570
box -12 -8 112 252
use OAI21X1  _3197_
timestamp 1728305162
transform -1 0 2690 0 1 4570
box -12 -8 112 252
use OAI21X1  _3198_
timestamp 1728305162
transform -1 0 2290 0 -1 6490
box -12 -8 112 252
use OAI21X1  _3199_
timestamp 1728305162
transform -1 0 2550 0 -1 6490
box -12 -8 112 252
use OAI21X1  _3200_
timestamp 1728305162
transform 1 0 890 0 -1 6970
box -12 -8 112 252
use OAI21X1  _3201_
timestamp 1728305162
transform -1 0 1230 0 1 6970
box -12 -8 112 252
use OAI21X1  _3202_
timestamp 1728305162
transform 1 0 1130 0 -1 6970
box -12 -8 112 252
use OAI21X1  _3203_
timestamp 1728305162
transform -1 0 1490 0 -1 6970
box -12 -8 112 252
use OAI21X1  _3204_
timestamp 1728305162
transform -1 0 750 0 -1 6970
box -12 -8 112 252
use OAI21X1  _3205_
timestamp 1728305162
transform -1 0 730 0 -1 7450
box -12 -8 112 252
use AND2X2  _3206_
timestamp 1728304163
transform 1 0 1170 0 -1 4090
box -12 -8 112 252
use NOR2X1  _3207_
timestamp 1728305106
transform -1 0 490 0 -1 5530
box -12 -8 92 252
use AOI21X1  _3208_
timestamp 1728304211
transform -1 0 250 0 -1 5530
box -12 -8 112 252
use NOR2X1  _3209_
timestamp 1728305106
transform 1 0 410 0 1 3610
box -12 -8 92 252
use AOI21X1  _3210_
timestamp 1728304211
transform -1 0 250 0 1 3610
box -12 -8 112 252
use NOR2X1  _3211_
timestamp 1728305106
transform -1 0 1730 0 -1 5530
box -12 -8 92 252
use AOI21X1  _3212_
timestamp 1728304211
transform -1 0 1490 0 -1 5530
box -12 -8 112 252
use NOR2X1  _3213_
timestamp 1728305106
transform 1 0 1670 0 -1 5050
box -12 -8 92 252
use AOI21X1  _3214_
timestamp 1728304211
transform 1 0 1430 0 -1 5050
box -12 -8 112 252
use NOR2X1  _3215_
timestamp 1728305106
transform -1 0 1450 0 -1 7450
box -12 -8 92 252
use AOI21X1  _3216_
timestamp 1728304211
transform 1 0 1110 0 -1 7450
box -12 -8 112 252
use NOR2X1  _3217_
timestamp 1728305106
transform -1 0 490 0 1 6010
box -12 -8 92 252
use AOI21X1  _3218_
timestamp 1728304211
transform -1 0 250 0 1 6010
box -12 -8 112 252
use NOR2X1  _3219_
timestamp 1728305106
transform -1 0 1770 0 -1 6490
box -12 -8 92 252
use AOI21X1  _3220_
timestamp 1728304211
transform 1 0 1930 0 -1 6490
box -12 -8 112 252
use NOR2X1  _3221_
timestamp 1728305106
transform -1 0 490 0 -1 6490
box -12 -8 92 252
use AOI21X1  _3222_
timestamp 1728304211
transform -1 0 270 0 -1 6490
box -12 -8 112 252
use NAND2X1  _3223_
timestamp 1728304996
transform -1 0 970 0 1 4090
box -12 -8 92 252
use INVX2  _3224_
timestamp 1728304826
transform 1 0 650 0 -1 4570
box -12 -8 72 252
use OAI21X1  _3225_
timestamp 1728305162
transform -1 0 510 0 1 5050
box -12 -8 112 252
use OAI21X1  _3226_
timestamp 1728305162
transform -1 0 250 0 1 5050
box -12 -8 112 252
use OAI21X1  _3227_
timestamp 1728305162
transform -1 0 530 0 1 4090
box -12 -8 112 252
use OAI21X1  _3228_
timestamp 1728305162
transform -1 0 270 0 1 4090
box -12 -8 112 252
use OAI21X1  _3229_
timestamp 1728305162
transform -1 0 2170 0 -1 6010
box -12 -8 112 252
use OAI21X1  _3230_
timestamp 1728305162
transform 1 0 1830 0 -1 6010
box -12 -8 112 252
use OAI21X1  _3231_
timestamp 1728305162
transform 1 0 1610 0 1 4570
box -12 -8 112 252
use OAI21X1  _3232_
timestamp 1728305162
transform -1 0 1970 0 1 4570
box -12 -8 112 252
use OAI21X1  _3233_
timestamp 1728305162
transform 1 0 1190 0 -1 6490
box -12 -8 112 252
use OAI21X1  _3234_
timestamp 1728305162
transform -1 0 1530 0 -1 6490
box -12 -8 112 252
use OAI21X1  _3235_
timestamp 1728305162
transform 1 0 1150 0 1 6010
box -12 -8 112 252
use OAI21X1  _3236_
timestamp 1728305162
transform 1 0 1410 0 1 6010
box -12 -8 112 252
use OAI21X1  _3237_
timestamp 1728305162
transform 1 0 2310 0 -1 6010
box -12 -8 112 252
use OAI21X1  _3238_
timestamp 1728305162
transform 1 0 2570 0 -1 6010
box -12 -8 112 252
use OAI21X1  _3239_
timestamp 1728305162
transform -1 0 730 0 1 6010
box -12 -8 112 252
use OAI21X1  _3240_
timestamp 1728305162
transform -1 0 990 0 1 6010
box -12 -8 112 252
use OAI21X1  _3241_
timestamp 1728305162
transform 1 0 9810 0 -1 3610
box -12 -8 112 252
use OAI21X1  _3242_
timestamp 1728305162
transform -1 0 9210 0 -1 2650
box -12 -8 112 252
use NOR2X1  _3243_
timestamp 1728305106
transform 1 0 9570 0 -1 3610
box -12 -8 92 252
use OAI21X1  _3244_
timestamp 1728305162
transform 1 0 8870 0 1 3130
box -12 -8 112 252
use AOI21X1  _3245_
timestamp 1728304211
transform 1 0 9150 0 1 3610
box -12 -8 112 252
use AND2X2  _3246_
timestamp 1728304163
transform -1 0 9770 0 1 3610
box -12 -8 112 252
use INVX1  _3247_
timestamp 1728304789
transform 1 0 10570 0 -1 5050
box -12 -8 72 252
use OAI21X1  _3248_
timestamp 1728305162
transform 1 0 10850 0 1 5050
box -12 -8 112 252
use AND2X2  _3249_
timestamp 1728304163
transform -1 0 9670 0 -1 250
box -12 -8 112 252
use NAND3X1  _3250_
timestamp 1728305047
transform 1 0 9490 0 -1 5530
box -12 -8 112 252
use OR2X2  _3251_
timestamp 1728305284
transform 1 0 9350 0 1 3130
box -12 -8 112 252
use NOR2X1  _3252_
timestamp 1728305106
transform -1 0 9410 0 -1 3610
box -12 -8 92 252
use OAI21X1  _3253_
timestamp 1728305162
transform -1 0 8070 0 1 3610
box -12 -8 112 252
use NOR2X1  _3254_
timestamp 1728305106
transform -1 0 8310 0 1 3610
box -12 -8 92 252
use AOI22X1  _3255_
timestamp 1728304278
transform -1 0 9510 0 1 3610
box -14 -8 132 252
use OAI21X1  _3256_
timestamp 1728305162
transform 1 0 8370 0 -1 5050
box -12 -8 112 252
use NOR2X1  _3257_
timestamp 1728305106
transform 1 0 8130 0 -1 5050
box -12 -8 92 252
use NAND3X1  _3258_
timestamp 1728305047
transform 1 0 8650 0 1 5050
box -12 -8 112 252
use OAI21X1  _3259_
timestamp 1728305162
transform 1 0 9610 0 1 5050
box -12 -8 112 252
use AOI21X1  _3260_
timestamp 1728304211
transform -1 0 11030 0 1 5530
box -12 -8 112 252
use AND2X2  _3261_
timestamp 1728304163
transform -1 0 10590 0 -1 5530
box -12 -8 112 252
use NAND3X1  _3262_
timestamp 1728305047
transform 1 0 10090 0 1 5050
box -12 -8 112 252
use OAI21X1  _3263_
timestamp 1728305162
transform 1 0 9750 0 1 4570
box -12 -8 112 252
use NOR2X1  _3264_
timestamp 1728305106
transform 1 0 9110 0 -1 3610
box -12 -8 92 252
use NAND3X1  _3265_
timestamp 1728305047
transform -1 0 9930 0 -1 5050
box -12 -8 112 252
use NOR2X1  _3266_
timestamp 1728305106
transform 1 0 9850 0 1 5050
box -12 -8 92 252
use NAND2X1  _3267_
timestamp 1728304996
transform -1 0 9830 0 -1 5530
box -12 -8 92 252
use OAI21X1  _3268_
timestamp 1728305162
transform -1 0 10170 0 -1 5050
box -12 -8 112 252
use AND2X2  _3269_
timestamp 1728304163
transform -1 0 10690 0 1 5050
box -12 -8 112 252
use NAND3X1  _3270_
timestamp 1728305047
transform 1 0 10330 0 -1 5050
box -12 -8 112 252
use NOR2X1  _3271_
timestamp 1728305106
transform -1 0 10190 0 -1 3130
box -12 -8 92 252
use OAI21X1  _3272_
timestamp 1728305162
transform 1 0 10370 0 -1 4570
box -12 -8 112 252
use NAND3X1  _3273_
timestamp 1728305047
transform -1 0 10350 0 1 4570
box -12 -8 112 252
use OR2X2  _3274_
timestamp 1728305284
transform -1 0 10430 0 1 5050
box -12 -8 112 252
use OAI21X1  _3275_
timestamp 1728305162
transform 1 0 9690 0 1 5530
box -12 -8 112 252
use NOR2X1  _3276_
timestamp 1728305106
transform -1 0 9350 0 -1 5530
box -12 -8 92 252
use AND2X2  _3277_
timestamp 1728304163
transform -1 0 10850 0 -1 5530
box -12 -8 112 252
use NAND3X1  _3278_
timestamp 1728305047
transform 1 0 10230 0 -1 5530
box -12 -8 112 252
use OAI21X1  _3279_
timestamp 1728305162
transform -1 0 10070 0 -1 5530
box -12 -8 112 252
use OAI21X1  _3280_
timestamp 1728305162
transform 1 0 9350 0 1 4090
box -12 -8 112 252
use OAI21X1  _3281_
timestamp 1728305162
transform 1 0 9090 0 1 4090
box -12 -8 112 252
use NOR2X1  _3282_
timestamp 1728305106
transform -1 0 7050 0 1 4090
box -12 -8 92 252
use NAND2X1  _3283_
timestamp 1728304996
transform -1 0 6990 0 -1 5050
box -12 -8 92 252
use NAND2X1  _3284_
timestamp 1728304996
transform 1 0 6670 0 -1 5050
box -12 -8 92 252
use NAND2X1  _3285_
timestamp 1728304996
transform 1 0 7130 0 -1 6490
box -12 -8 92 252
use OAI21X1  _3286_
timestamp 1728305162
transform -1 0 7470 0 -1 6490
box -12 -8 112 252
use NAND2X1  _3287_
timestamp 1728304996
transform -1 0 6790 0 -1 6970
box -12 -8 92 252
use OAI21X1  _3288_
timestamp 1728305162
transform -1 0 7050 0 -1 6970
box -12 -8 112 252
use NAND2X1  _3289_
timestamp 1728304996
transform -1 0 6970 0 1 5530
box -12 -8 92 252
use OAI21X1  _3290_
timestamp 1728305162
transform 1 0 6650 0 1 5530
box -12 -8 112 252
use NAND2X1  _3291_
timestamp 1728304996
transform 1 0 7150 0 1 6010
box -12 -8 92 252
use OAI21X1  _3292_
timestamp 1728305162
transform -1 0 7470 0 1 6010
box -12 -8 112 252
use NAND2X1  _3293_
timestamp 1728304996
transform 1 0 7250 0 1 6970
box -12 -8 92 252
use OAI21X1  _3294_
timestamp 1728305162
transform 1 0 6990 0 1 6970
box -12 -8 112 252
use NAND2X1  _3295_
timestamp 1728304996
transform 1 0 6170 0 1 6010
box -12 -8 92 252
use OAI21X1  _3296_
timestamp 1728305162
transform 1 0 5930 0 1 6010
box -12 -8 112 252
use NAND2X1  _3297_
timestamp 1728304996
transform 1 0 5530 0 1 6490
box -12 -8 92 252
use OAI21X1  _3298_
timestamp 1728305162
transform 1 0 5290 0 1 6490
box -12 -8 112 252
use NAND2X1  _3299_
timestamp 1728304996
transform 1 0 5730 0 -1 6490
box -12 -8 92 252
use OAI21X1  _3300_
timestamp 1728305162
transform 1 0 5470 0 -1 6490
box -12 -8 112 252
use AOI21X1  _3301_
timestamp 1728304211
transform 1 0 6990 0 -1 5530
box -12 -8 112 252
use NAND2X1  _3302_
timestamp 1728304996
transform 1 0 3050 0 1 8890
box -12 -8 92 252
use OAI21X1  _3303_
timestamp 1728305162
transform -1 0 3210 0 -1 8890
box -12 -8 112 252
use NAND2X1  _3304_
timestamp 1728304996
transform 1 0 2070 0 1 9850
box -12 -8 92 252
use OAI21X1  _3305_
timestamp 1728305162
transform -1 0 2390 0 1 9850
box -12 -8 112 252
use NAND2X1  _3306_
timestamp 1728304996
transform 1 0 3990 0 1 9850
box -12 -8 92 252
use OAI21X1  _3307_
timestamp 1728305162
transform -1 0 5010 0 1 9850
box -12 -8 112 252
use NAND2X1  _3308_
timestamp 1728304996
transform -1 0 230 0 -1 9850
box -12 -8 92 252
use OAI21X1  _3309_
timestamp 1728305162
transform -1 0 270 0 1 9370
box -12 -8 112 252
use NAND2X1  _3310_
timestamp 1728304996
transform -1 0 910 0 -1 9850
box -12 -8 92 252
use OAI21X1  _3311_
timestamp 1728305162
transform -1 0 990 0 1 9370
box -12 -8 112 252
use NAND2X1  _3312_
timestamp 1728304996
transform -1 0 470 0 -1 9850
box -12 -8 92 252
use OAI21X1  _3313_
timestamp 1728305162
transform -1 0 510 0 1 9370
box -12 -8 112 252
use NAND2X1  _3314_
timestamp 1728304996
transform -1 0 250 0 -1 8890
box -12 -8 92 252
use OAI21X1  _3315_
timestamp 1728305162
transform -1 0 270 0 1 8410
box -12 -8 112 252
use NAND2X1  _3316_
timestamp 1728304996
transform -1 0 730 0 1 8410
box -12 -8 92 252
use OAI21X1  _3317_
timestamp 1728305162
transform -1 0 990 0 1 8410
box -12 -8 112 252
use DFFSR  _3318_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728387359
transform 1 0 10350 0 1 730
box -12 -8 492 252
use DFFSR  _3319_
timestamp 1728387359
transform 1 0 9810 0 1 250
box -12 -8 492 252
use DFFSR  _3320_
timestamp 1728387359
transform -1 0 9190 0 -1 250
box -12 -8 492 252
use DFFSR  _3321_
timestamp 1728387359
transform 1 0 10290 0 1 250
box -12 -8 492 252
use DFFSR  _3322_
timestamp 1728387359
transform 1 0 9650 0 -1 730
box -12 -8 492 252
use DFFSR  _3323_
timestamp 1728387359
transform 1 0 7530 0 1 730
box -12 -8 492 252
use DFFSR  _3324_
timestamp 1728387359
transform 1 0 7210 0 -1 8890
box -12 -8 492 252
use DFFSR  _3325_
timestamp 1728387359
transform -1 0 6930 0 -1 8890
box -12 -8 492 252
use DFFSR  _3326_
timestamp 1728387359
transform -1 0 7870 0 1 10330
box -12 -8 492 252
use DFFSR  _3327_
timestamp 1728387359
transform -1 0 7490 0 1 9370
box -12 -8 492 252
use DFFSR  _3328_
timestamp 1728387359
transform 1 0 5970 0 1 9850
box -12 -8 492 252
use DFFSR  _3329_
timestamp 1728387359
transform -1 0 6270 0 -1 10330
box -12 -8 492 252
use DFFSR  _3330_
timestamp 1728387359
transform 1 0 6310 0 1 10810
box -12 -8 492 252
use DFFSR  _3331_
timestamp 1728387359
transform 1 0 5650 0 1 10330
box -12 -8 492 252
use DFFSR  _3332_
timestamp 1728387359
transform -1 0 4670 0 1 10330
box -12 -8 492 252
use DFFSR  _3333_
timestamp 1728387359
transform 1 0 3210 0 1 10810
box -12 -8 492 252
use DFFSR  _3334_
timestamp 1728387359
transform 1 0 2770 0 -1 11290
box -12 -8 492 252
use DFFSR  _3335_
timestamp 1728387359
transform 1 0 710 0 1 10330
box -12 -8 492 252
use DFFSR  _3336_
timestamp 1728387359
transform 1 0 10 0 1 10810
box -12 -8 492 252
use DFFSR  _3337_
timestamp 1728387359
transform 1 0 1710 0 1 10810
box -12 -8 492 252
use DFFSR  _3338_
timestamp 1728387359
transform 1 0 250 0 -1 8890
box -12 -8 492 252
use DFFSR  _3339_
timestamp 1728387359
transform 1 0 230 0 1 9850
box -12 -8 492 252
use DFFSR  _3340_
timestamp 1728387359
transform 1 0 3910 0 -1 6010
box -12 -8 492 252
use DFFSR  _3341_
timestamp 1728387359
transform -1 0 6550 0 -1 6010
box -12 -8 492 252
use DFFSR  _3342_
timestamp 1728387359
transform 1 0 2670 0 1 3130
box -12 -8 492 252
use DFFSR  _3343_
timestamp 1728387359
transform 1 0 1770 0 -1 3610
box -12 -8 492 252
use DFFSR  _3344_
timestamp 1728387359
transform 1 0 4610 0 1 4570
box -12 -8 492 252
use DFFSR  _3345_
timestamp 1728387359
transform 1 0 3370 0 -1 2650
box -12 -8 492 252
use DFFSR  _3346_
timestamp 1728387359
transform 1 0 3710 0 1 5050
box -12 -8 492 252
use DFFSR  _3347_
timestamp 1728387359
transform -1 0 5230 0 1 2170
box -12 -8 492 252
use DFFSR  _3348_
timestamp 1728387359
transform 1 0 4590 0 1 1690
box -12 -8 492 252
use DFFSR  _3349_
timestamp 1728387359
transform 1 0 3570 0 1 2650
box -12 -8 492 252
use DFFSR  _3350_
timestamp 1728387359
transform 1 0 3910 0 -1 2170
box -12 -8 492 252
use DFFSR  _3351_
timestamp 1728387359
transform 1 0 5290 0 1 1690
box -12 -8 492 252
use DFFSR  _3352_
timestamp 1728387359
transform 1 0 4850 0 -1 2170
box -12 -8 492 252
use DFFSR  _3353_
timestamp 1728387359
transform 1 0 970 0 -1 3130
box -12 -8 492 252
use DFFSR  _3354_
timestamp 1728387359
transform 1 0 1690 0 1 2650
box -12 -8 492 252
use DFFSR  _3355_
timestamp 1728387359
transform 1 0 1690 0 1 3130
box -12 -8 492 252
use DFFSR  _3356_
timestamp 1728387359
transform 1 0 2650 0 -1 2650
box -12 -8 492 252
use DFFSR  _3357_
timestamp 1728387359
transform 1 0 4050 0 1 2170
box -12 -8 492 252
use DFFSR  _3358_
timestamp 1728387359
transform 1 0 3910 0 1 4570
box -12 -8 492 252
use DFFSR  _3359_
timestamp 1728387359
transform 1 0 4790 0 -1 3130
box -12 -8 492 252
use DFFSR  _3360_
timestamp 1728387359
transform 1 0 3350 0 -1 3130
box -12 -8 492 252
use DFFSR  _3361_
timestamp 1728387359
transform -1 0 3810 0 1 2170
box -12 -8 492 252
use DFFSR  _3362_
timestamp 1728387359
transform 1 0 2630 0 1 2170
box -12 -8 492 252
use DFFSR  _3363_
timestamp 1728387359
transform 1 0 3210 0 -1 3610
box -12 -8 492 252
use DFFSR  _3364_
timestamp 1728387359
transform 1 0 3770 0 -1 4090
box -12 -8 492 252
use DFFSR  _3365_
timestamp 1728387359
transform 1 0 2570 0 1 1690
box -12 -8 492 252
use DFFSR  _3366_
timestamp 1728387359
transform 1 0 5230 0 1 2170
box -12 -8 492 252
use DFFSR  _3367_
timestamp 1728387359
transform 1 0 5750 0 -1 730
box -12 -8 492 252
use DFFSR  _3368_
timestamp 1728387359
transform 1 0 230 0 -1 2650
box -12 -8 492 252
use DFFSR  _3369_
timestamp 1728387359
transform -1 0 5110 0 1 1210
box -12 -8 492 252
use DFFSR  _3370_
timestamp 1728387359
transform 1 0 10 0 -1 2170
box -12 -8 492 252
use DFFSR  _3371_
timestamp 1728387359
transform -1 0 970 0 -1 2170
box -12 -8 492 252
use DFFSR  _3372_
timestamp 1728387359
transform 1 0 10 0 1 1690
box -12 -8 492 252
use DFFSR  _3373_
timestamp 1728387359
transform 1 0 10 0 1 2170
box -12 -8 492 252
use DFFSR  _3374_
timestamp 1728387359
transform 1 0 710 0 -1 2650
box -12 -8 492 252
use DFFSR  _3375_
timestamp 1728387359
transform -1 0 5310 0 1 10810
box -12 -8 492 252
use DFFSR  _3376_
timestamp 1728387359
transform -1 0 6310 0 -1 11290
box -12 -8 492 252
use DFFSR  _3377_
timestamp 1728387359
transform 1 0 4670 0 -1 11290
box -12 -8 492 252
use DFFSR  _3378_
timestamp 1728387359
transform 1 0 7030 0 -1 10810
box -12 -8 492 252
use DFFSR  _3379_
timestamp 1728387359
transform 1 0 5310 0 1 10810
box -12 -8 492 252
use DFFSR  _3380_
timestamp 1728387359
transform 1 0 1850 0 -1 11290
box -12 -8 492 252
use DFFSR  _3381_
timestamp 1728387359
transform 1 0 7830 0 -1 9850
box -12 -8 492 252
use DFFSR  _3382_
timestamp 1728387359
transform 1 0 7490 0 1 9370
box -12 -8 492 252
use DFFSR  _3383_
timestamp 1728387359
transform 1 0 3130 0 1 8410
box -12 -8 492 252
use DFFPOSX1  _3384_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728340458
transform -1 0 4130 0 1 5530
box -13 -8 253 252
use DFFPOSX1  _3385_
timestamp 1728340458
transform -1 0 3390 0 1 5530
box -13 -8 253 252
use DFFPOSX1  _3386_
timestamp 1728340458
transform -1 0 4410 0 -1 5050
box -13 -8 253 252
use DFFPOSX1  _3387_
timestamp 1728340458
transform 1 0 3710 0 -1 4570
box -13 -8 253 252
use DFFPOSX1  _3388_
timestamp 1728340458
transform 1 0 2250 0 1 5050
box -13 -8 253 252
use DFFPOSX1  _3389_
timestamp 1728340458
transform -1 0 3150 0 -1 6010
box -13 -8 253 252
use DFFPOSX1  _3390_
timestamp 1728340458
transform -1 0 3730 0 -1 5530
box -13 -8 253 252
use DFFPOSX1  _3391_
timestamp 1728340458
transform 1 0 2950 0 1 5050
box -13 -8 253 252
use DFFSR  _3392_
timestamp 1728387359
transform -1 0 3110 0 1 4090
box -12 -8 492 252
use DFFSR  _3393_
timestamp 1728387359
transform 1 0 6970 0 1 5530
box -12 -8 492 252
use DFFSR  _3394_
timestamp 1728387359
transform -1 0 5430 0 -1 4570
box -12 -8 492 252
use DFFSR  _3395_
timestamp 1728387359
transform -1 0 6290 0 1 4570
box -12 -8 492 252
use DFFSR  _3396_
timestamp 1728387359
transform 1 0 4870 0 -1 5050
box -12 -8 492 252
use DFFSR  _3397_
timestamp 1728387359
transform 1 0 5030 0 1 5530
box -12 -8 492 252
use DFFSR  _3398_
timestamp 1728387359
transform 1 0 5230 0 1 2650
box -12 -8 492 252
use DFFSR  _3399_
timestamp 1728387359
transform 1 0 7490 0 -1 11290
box -12 -8 492 252
use DFFSR  _3400_
timestamp 1728387359
transform 1 0 10 0 -1 4570
box -12 -8 492 252
use DFFSR  _3401_
timestamp 1728387359
transform 1 0 1050 0 -1 3610
box -12 -8 492 252
use DFFSR  _3402_
timestamp 1728387359
transform 1 0 510 0 1 5050
box -12 -8 492 252
use DFFSR  _3403_
timestamp 1728387359
transform -1 0 2390 0 1 5530
box -12 -8 492 252
use DFFSR  _3404_
timestamp 1728387359
transform 1 0 850 0 1 7930
box -12 -8 492 252
use DFFSR  _3405_
timestamp 1728387359
transform 1 0 10 0 1 7930
box -12 -8 492 252
use DFFSR  _3406_
timestamp 1728387359
transform -1 0 2750 0 1 6490
box -12 -8 492 252
use DFFSR  _3407_
timestamp 1728387359
transform 1 0 10 0 1 6970
box -12 -8 492 252
use DFFSR  _3408_
timestamp 1728387359
transform -1 0 1230 0 1 4570
box -12 -8 492 252
use DFFSR  _3409_
timestamp 1728387359
transform 1 0 970 0 1 4090
box -12 -8 492 252
use DFFSR  _3410_
timestamp 1728387359
transform -1 0 3930 0 1 6010
box -12 -8 492 252
use DFFSR  _3411_
timestamp 1728387359
transform -1 0 2630 0 -1 4570
box -12 -8 492 252
use DFFSR  _3412_
timestamp 1728387359
transform -1 0 2270 0 1 6490
box -12 -8 492 252
use DFFSR  _3413_
timestamp 1728387359
transform 1 0 490 0 1 6970
box -12 -8 492 252
use DFFSR  _3414_
timestamp 1728387359
transform 1 0 1230 0 1 6970
box -12 -8 492 252
use DFFSR  _3415_
timestamp 1728387359
transform 1 0 10 0 1 7450
box -12 -8 492 252
use DFFSR  _3416_
timestamp 1728387359
transform 1 0 10 0 1 5530
box -12 -8 492 252
use DFFSR  _3417_
timestamp 1728387359
transform 1 0 10 0 -1 3610
box -12 -8 492 252
use DFFSR  _3418_
timestamp 1728387359
transform 1 0 1170 0 1 5530
box -12 -8 492 252
use DFFSR  _3419_
timestamp 1728387359
transform 1 0 990 0 1 5050
box -12 -8 492 252
use DFFSR  _3420_
timestamp 1728387359
transform 1 0 990 0 1 7450
box -12 -8 492 252
use DFFSR  _3421_
timestamp 1728387359
transform 1 0 10 0 -1 6010
box -12 -8 492 252
use DFFSR  _3422_
timestamp 1728387359
transform -1 0 2470 0 1 6010
box -12 -8 492 252
use DFFSR  _3423_
timestamp 1728387359
transform 1 0 10 0 1 6490
box -12 -8 492 252
use DFFSR  _3424_
timestamp 1728387359
transform 1 0 4230 0 -1 5530
box -12 -8 492 252
use DFFSR  _3425_
timestamp 1728387359
transform 1 0 10 0 -1 5050
box -12 -8 492 252
use DFFSR  _3426_
timestamp 1728387359
transform 1 0 10 0 -1 4090
box -12 -8 492 252
use DFFSR  _3427_
timestamp 1728387359
transform 1 0 1190 0 -1 6010
box -12 -8 492 252
use DFFSR  _3428_
timestamp 1728387359
transform -1 0 2450 0 1 4570
box -12 -8 492 252
use DFFSR  _3429_
timestamp 1728387359
transform 1 0 750 0 1 6490
box -12 -8 492 252
use DFFSR  _3430_
timestamp 1728387359
transform -1 0 1990 0 1 6010
box -12 -8 492 252
use DFFSR  _3431_
timestamp 1728387359
transform 1 0 2470 0 1 6010
box -12 -8 492 252
use DFFSR  _3432_
timestamp 1728387359
transform -1 0 970 0 -1 6010
box -12 -8 492 252
use DFFSR  _3433_
timestamp 1728387359
transform -1 0 6970 0 -1 6490
box -12 -8 492 252
use DFFSR  _3434_
timestamp 1728387359
transform -1 0 6570 0 -1 6970
box -12 -8 492 252
use DFFSR  _3435_
timestamp 1728387359
transform -1 0 6830 0 -1 5530
box -12 -8 492 252
use DFFSR  _3436_
timestamp 1728387359
transform -1 0 7550 0 -1 6010
box -12 -8 492 252
use DFFSR  _3437_
timestamp 1728387359
transform 1 0 6770 0 1 7450
box -12 -8 492 252
use DFFSR  _3438_
timestamp 1728387359
transform -1 0 6730 0 1 6010
box -12 -8 492 252
use DFFSR  _3439_
timestamp 1728387359
transform 1 0 4650 0 1 6490
box -12 -8 492 252
use DFFSR  _3440_
timestamp 1728387359
transform 1 0 4850 0 -1 6490
box -12 -8 492 252
use DFFSR  _3441_
timestamp 1728387359
transform 1 0 3130 0 1 8890
box -12 -8 492 252
use DFFSR  _3442_
timestamp 1728387359
transform 1 0 1930 0 -1 9850
box -12 -8 492 252
use DFFSR  _3443_
timestamp 1728387359
transform -1 0 4750 0 1 9850
box -12 -8 492 252
use DFFSR  _3444_
timestamp 1728387359
transform 1 0 10 0 -1 9370
box -12 -8 492 252
use DFFSR  _3445_
timestamp 1728387359
transform 1 0 690 0 -1 9370
box -12 -8 492 252
use DFFSR  _3446_
timestamp 1728387359
transform 1 0 250 0 1 8890
box -12 -8 492 252
use DFFSR  _3447_
timestamp 1728387359
transform 1 0 10 0 -1 8410
box -12 -8 492 252
use DFFSR  _3448_
timestamp 1728387359
transform 1 0 690 0 -1 8410
box -12 -8 492 252
use OR2X2  _3449_
timestamp 1728305284
transform -1 0 3990 0 -1 7450
box -12 -8 112 252
use NOR2X1  _3450_
timestamp 1728305106
transform 1 0 3090 0 1 7450
box -12 -8 92 252
use NOR2X1  _3451_
timestamp 1728305106
transform 1 0 3210 0 -1 7930
box -12 -8 92 252
use NOR2X1  _3452_
timestamp 1728305106
transform -1 0 3510 0 -1 7450
box -12 -8 92 252
use NAND3X1  _3453_
timestamp 1728305047
transform 1 0 3330 0 1 7450
box -12 -8 112 252
use NOR2X1  _3454_
timestamp 1728305106
transform -1 0 3750 0 -1 7450
box -12 -8 92 252
use INVX1  _3455_
timestamp 1728304789
transform 1 0 10050 0 -1 6970
box -12 -8 72 252
use AND2X2  _3456_
timestamp 1728304163
transform 1 0 9630 0 1 6490
box -12 -8 112 252
use NOR2X1  _3457_
timestamp 1728305106
transform -1 0 9950 0 1 6490
box -12 -8 92 252
use NOR2X1  _3458_
timestamp 1728305106
transform -1 0 10130 0 -1 6490
box -12 -8 92 252
use INVX1  _3459_
timestamp 1728304789
transform 1 0 10510 0 -1 6970
box -12 -8 72 252
use NOR2X1  _3460_
timestamp 1728305106
transform -1 0 10850 0 -1 6490
box -12 -8 92 252
use NAND2X1  _3461_
timestamp 1728304996
transform -1 0 10630 0 1 6490
box -12 -8 92 252
use INVX1  _3462_
timestamp 1728304789
transform -1 0 10150 0 1 6490
box -12 -8 72 252
use OAI21X1  _3463_
timestamp 1728305162
transform 1 0 10530 0 -1 6490
box -12 -8 112 252
use NOR2X1  _3464_
timestamp 1728305106
transform -1 0 10390 0 1 6490
box -12 -8 92 252
use OAI21X1  _3465_
timestamp 1728305162
transform 1 0 10270 0 -1 6490
box -12 -8 112 252
use NAND2X1  _3466_
timestamp 1728304996
transform -1 0 10370 0 1 6010
box -12 -8 92 252
use INVX4  _3467_
timestamp 1728304878
transform 1 0 8370 0 1 6010
box -12 -8 92 252
use INVX4  _3468_
timestamp 1728304878
transform 1 0 9190 0 1 7930
box -12 -8 92 252
use NAND2X1  _3469_
timestamp 1728304996
transform 1 0 8670 0 -1 6970
box -12 -8 92 252
use INVX2  _3470_
timestamp 1728304826
transform -1 0 8630 0 -1 7930
box -12 -8 72 252
use NAND2X1  _3471_
timestamp 1728304996
transform 1 0 8750 0 1 7930
box -12 -8 92 252
use INVX2  _3472_
timestamp 1728304826
transform 1 0 8990 0 1 7930
box -12 -8 72 252
use AND2X2  _3473_
timestamp 1728304163
transform -1 0 8870 0 -1 7930
box -12 -8 112 252
use NAND2X1  _3474_
timestamp 1728304996
transform -1 0 8990 0 1 7450
box -12 -8 92 252
use AOI22X1  _3475_
timestamp 1728304278
transform -1 0 9150 0 -1 7930
box -14 -8 132 252
use INVX2  _3476_
timestamp 1728304826
transform 1 0 9830 0 1 7450
box -12 -8 72 252
use OAI21X1  _3477_
timestamp 1728305162
transform 1 0 9290 0 -1 7450
box -12 -8 112 252
use OAI21X1  _3478_
timestamp 1728305162
transform -1 0 9230 0 1 7450
box -12 -8 112 252
use INVX4  _3479_
timestamp 1728304878
transform 1 0 10650 0 -1 9850
box -12 -8 92 252
use OAI21X1  _3480_
timestamp 1728305162
transform -1 0 10290 0 1 7930
box -12 -8 112 252
use AOI21X1  _3481_
timestamp 1728304211
transform -1 0 10130 0 -1 7930
box -12 -8 112 252
use NOR2X1  _3482_
timestamp 1728305106
transform -1 0 9930 0 1 10330
box -12 -8 92 252
use OR2X2  _3483_
timestamp 1728305284
transform 1 0 10990 0 -1 7450
box -12 -8 112 252
use OAI21X1  _3484_
timestamp 1728305162
transform 1 0 10990 0 1 6970
box -12 -8 112 252
use NAND2X1  _3485_
timestamp 1728304996
transform 1 0 11270 0 1 6490
box -12 -8 92 252
use OAI21X1  _3486_
timestamp 1728305162
transform 1 0 11210 0 -1 6970
box -12 -8 112 252
use NAND2X1  _3487_
timestamp 1728304996
transform 1 0 10990 0 -1 6970
box -12 -8 92 252
use NAND2X1  _3488_
timestamp 1728304996
transform 1 0 9630 0 -1 8410
box -12 -8 92 252
use AND2X2  _3489_
timestamp 1728304163
transform 1 0 9510 0 1 8410
box -12 -8 112 252
use NAND2X1  _3490_
timestamp 1728304996
transform -1 0 9850 0 1 8410
box -12 -8 92 252
use AOI22X1  _3491_
timestamp 1728304278
transform -1 0 9890 0 -1 8890
box -14 -8 132 252
use OAI21X1  _3492_
timestamp 1728305162
transform 1 0 10010 0 1 8410
box -12 -8 112 252
use OAI21X1  _3493_
timestamp 1728305162
transform 1 0 10270 0 1 8410
box -12 -8 112 252
use NAND2X1  _3494_
timestamp 1728304996
transform 1 0 10390 0 -1 9370
box -12 -8 92 252
use INVX2  _3495_
timestamp 1728304826
transform -1 0 8950 0 -1 8410
box -12 -8 72 252
use OAI21X1  _3496_
timestamp 1728305162
transform 1 0 9530 0 -1 8890
box -12 -8 112 252
use OAI21X1  _3497_
timestamp 1728305162
transform 1 0 10030 0 -1 8890
box -12 -8 112 252
use NAND2X1  _3498_
timestamp 1728304996
transform 1 0 9910 0 -1 9370
box -12 -8 92 252
use AND2X2  _3499_
timestamp 1728304163
transform 1 0 9310 0 1 8890
box -12 -8 112 252
use NAND2X1  _3500_
timestamp 1728304996
transform -1 0 9650 0 1 8890
box -12 -8 92 252
use AOI22X1  _3501_
timestamp 1728304278
transform -1 0 9930 0 1 8890
box -14 -8 132 252
use OAI21X1  _3502_
timestamp 1728305162
transform 1 0 9650 0 -1 9370
box -12 -8 112 252
use OAI21X1  _3503_
timestamp 1728305162
transform 1 0 10150 0 -1 9370
box -12 -8 112 252
use OAI21X1  _3504_
timestamp 1728305162
transform -1 0 10190 0 1 8890
box -12 -8 112 252
use OAI21X1  _3505_
timestamp 1728305162
transform 1 0 10330 0 1 8890
box -12 -8 112 252
use NAND2X1  _3506_
timestamp 1728304996
transform 1 0 10870 0 -1 9370
box -12 -8 92 252
use INVX1  _3507_
timestamp 1728304789
transform -1 0 9510 0 -1 9370
box -12 -8 72 252
use INVX1  _3508_
timestamp 1728304789
transform -1 0 8650 0 -1 8890
box -12 -8 72 252
use INVX1  _3509_
timestamp 1728304789
transform 1 0 8530 0 1 7930
box -12 -8 72 252
use NAND2X1  _3510_
timestamp 1728304996
transform 1 0 9290 0 -1 8890
box -12 -8 92 252
use OAI21X1  _3511_
timestamp 1728305162
transform -1 0 9150 0 -1 8890
box -12 -8 112 252
use OAI21X1  _3512_
timestamp 1728305162
transform 1 0 8790 0 -1 8890
box -12 -8 112 252
use AOI21X1  _3513_
timestamp 1728304211
transform -1 0 9170 0 1 8890
box -12 -8 112 252
use NAND2X1  _3514_
timestamp 1728304996
transform -1 0 8910 0 1 8890
box -12 -8 92 252
use OAI21X1  _3515_
timestamp 1728305162
transform -1 0 9310 0 -1 9370
box -12 -8 112 252
use INVX1  _3516_
timestamp 1728304789
transform 1 0 11090 0 -1 9850
box -12 -8 72 252
use OAI21X1  _3517_
timestamp 1728305162
transform -1 0 10490 0 -1 9850
box -12 -8 112 252
use OAI21X1  _3518_
timestamp 1728305162
transform 1 0 10470 0 1 9850
box -12 -8 112 252
use AND2X2  _3519_
timestamp 1728304163
transform 1 0 10970 0 1 9850
box -12 -8 112 252
use OR2X2  _3520_
timestamp 1728305284
transform -1 0 11330 0 -1 10330
box -12 -8 112 252
use NAND3X1  _3521_
timestamp 1728305047
transform 1 0 7590 0 -1 8410
box -12 -8 112 252
use AOI22X1  _3522_
timestamp 1728304278
transform -1 0 8210 0 -1 8410
box -14 -8 132 252
use INVX1  _3523_
timestamp 1728304789
transform 1 0 8830 0 1 8410
box -12 -8 72 252
use INVX1  _3524_
timestamp 1728304789
transform 1 0 8630 0 1 8410
box -12 -8 72 252
use OAI21X1  _3525_
timestamp 1728305162
transform 1 0 9050 0 1 8410
box -12 -8 112 252
use NAND2X1  _3526_
timestamp 1728304996
transform -1 0 9370 0 1 8410
box -12 -8 92 252
use OAI22X1  _3527_
timestamp 1728305200
transform -1 0 8490 0 -1 8410
box -12 -8 132 252
use NOR2X1  _3528_
timestamp 1728305106
transform -1 0 10070 0 1 9850
box -12 -8 92 252
use AOI21X1  _3529_
timestamp 1728304211
transform 1 0 10130 0 -1 9850
box -12 -8 112 252
use AOI21X1  _3530_
timestamp 1728304211
transform 1 0 10230 0 1 9850
box -12 -8 112 252
use NAND2X1  _3531_
timestamp 1728304996
transform -1 0 10310 0 -1 10330
box -12 -8 92 252
use INVX1  _3532_
timestamp 1728304789
transform 1 0 10410 0 -1 10810
box -12 -8 72 252
use NAND3X1  _3533_
timestamp 1728305047
transform -1 0 8410 0 1 8890
box -12 -8 112 252
use AOI22X1  _3534_
timestamp 1728304278
transform -1 0 8670 0 1 8890
box -14 -8 132 252
use INVX1  _3535_
timestamp 1728304789
transform -1 0 8190 0 1 9370
box -12 -8 72 252
use NOR2X1  _3536_
timestamp 1728305106
transform -1 0 8410 0 1 9370
box -12 -8 92 252
use OAI21X1  _3537_
timestamp 1728305162
transform 1 0 8470 0 -1 9370
box -12 -8 112 252
use OAI22X1  _3538_
timestamp 1728305200
transform -1 0 8850 0 -1 9370
box -12 -8 132 252
use OAI21X1  _3539_
timestamp 1728305162
transform -1 0 9710 0 -1 9850
box -12 -8 112 252
use AOI21X1  _3540_
timestamp 1728304211
transform 1 0 9870 0 -1 9850
box -12 -8 112 252
use OAI21X1  _3541_
timestamp 1728305162
transform -1 0 10010 0 -1 10810
box -12 -8 112 252
use NAND2X1  _3542_
timestamp 1728304996
transform -1 0 7670 0 1 8890
box -12 -8 92 252
use NAND2X1  _3543_
timestamp 1728304996
transform -1 0 7930 0 -1 8410
box -12 -8 92 252
use AOI22X1  _3544_
timestamp 1728304278
transform 1 0 8070 0 -1 8890
box -14 -8 132 252
use INVX1  _3545_
timestamp 1728304789
transform 1 0 8950 0 -1 9850
box -12 -8 72 252
use INVX1  _3546_
timestamp 1728304789
transform -1 0 8430 0 -1 7930
box -12 -8 72 252
use OAI21X1  _3547_
timestamp 1728305162
transform 1 0 8790 0 1 9370
box -12 -8 112 252
use NAND2X1  _3548_
timestamp 1728304996
transform -1 0 9130 0 1 9370
box -12 -8 92 252
use NAND2X1  _3549_
timestamp 1728304996
transform -1 0 9070 0 -1 9370
box -12 -8 92 252
use OAI21X1  _3550_
timestamp 1728305162
transform 1 0 9010 0 1 9850
box -12 -8 112 252
use OAI21X1  _3551_
timestamp 1728305162
transform 1 0 9290 0 1 9370
box -12 -8 112 252
use INVX1  _3552_
timestamp 1728304789
transform 1 0 9410 0 -1 9850
box -12 -8 72 252
use OAI21X1  _3553_
timestamp 1728305162
transform 1 0 9170 0 -1 9850
box -12 -8 112 252
use OAI21X1  _3554_
timestamp 1728305162
transform 1 0 9090 0 1 10330
box -12 -8 112 252
use OAI21X1  _3555_
timestamp 1728305162
transform -1 0 8730 0 -1 8410
box -12 -8 112 252
use NOR2X1  _3556_
timestamp 1728305106
transform 1 0 8570 0 1 9370
box -12 -8 92 252
use MUX2X1  _3557_
timestamp 1728304958
transform -1 0 8310 0 -1 9370
box -12 -8 131 252
use NAND2X1  _3558_
timestamp 1728304996
transform -1 0 7930 0 -1 8890
box -12 -8 92 252
use NAND2X1  _3559_
timestamp 1728304996
transform 1 0 7830 0 1 8890
box -12 -8 92 252
use AOI21X1  _3560_
timestamp 1728304211
transform 1 0 8330 0 -1 8890
box -12 -8 112 252
use NAND2X1  _3561_
timestamp 1728304996
transform -1 0 8150 0 1 8890
box -12 -8 92 252
use NAND3X1  _3562_
timestamp 1728305047
transform -1 0 9150 0 -1 10330
box -12 -8 112 252
use AOI22X1  _3563_
timestamp 1728304278
transform -1 0 9170 0 1 10810
box -14 -8 132 252
use NOR2X1  _3564_
timestamp 1728305106
transform 1 0 10170 0 -1 10810
box -12 -8 92 252
use OAI21X1  _3565_
timestamp 1728305162
transform -1 0 10150 0 1 10810
box -12 -8 112 252
use NAND2X1  _3566_
timestamp 1728304996
transform 1 0 10010 0 -1 10330
box -12 -8 92 252
use INVX1  _3567_
timestamp 1728304789
transform 1 0 10090 0 1 10330
box -12 -8 72 252
use OAI21X1  _3568_
timestamp 1728305162
transform 1 0 10290 0 1 10330
box -12 -8 112 252
use INVX1  _3569_
timestamp 1728304789
transform 1 0 10310 0 1 10810
box -12 -8 72 252
use AND2X2  _3570_
timestamp 1728304163
transform 1 0 10750 0 1 10810
box -12 -8 112 252
use NAND2X1  _3571_
timestamp 1728304996
transform -1 0 10810 0 1 9850
box -12 -8 92 252
use OAI21X1  _3572_
timestamp 1728305162
transform -1 0 11330 0 1 9850
box -12 -8 112 252
use OAI21X1  _3573_
timestamp 1728305162
transform 1 0 11110 0 -1 10810
box -12 -8 112 252
use AOI21X1  _3574_
timestamp 1728304211
transform 1 0 10870 0 -1 10810
box -12 -8 112 252
use INVX1  _3575_
timestamp 1728304789
transform 1 0 11270 0 1 10810
box -12 -8 72 252
use NAND2X1  _3576_
timestamp 1728304996
transform 1 0 10030 0 -1 250
box -12 -8 92 252
use NAND2X1  _3577_
timestamp 1728304996
transform -1 0 11350 0 1 10330
box -12 -8 92 252
use INVX1  _3578_
timestamp 1728304789
transform 1 0 10870 0 -1 9850
box -12 -8 72 252
use NAND2X1  _3579_
timestamp 1728304996
transform -1 0 10650 0 -1 11290
box -12 -8 92 252
use AOI21X1  _3580_
timestamp 1728304211
transform -1 0 9370 0 1 9850
box -12 -8 112 252
use OAI21X1  _3581_
timestamp 1728305162
transform -1 0 9050 0 -1 10810
box -12 -8 112 252
use INVX1  _3582_
timestamp 1728304789
transform 1 0 8830 0 1 10810
box -12 -8 72 252
use NOR2X1  _3583_
timestamp 1728305106
transform -1 0 9210 0 -1 11290
box -12 -8 92 252
use OAI21X1  _3584_
timestamp 1728305162
transform 1 0 8870 0 -1 11290
box -12 -8 112 252
use INVX1  _3585_
timestamp 1728304789
transform -1 0 9670 0 1 10810
box -12 -8 72 252
use OAI21X1  _3586_
timestamp 1728305162
transform 1 0 9190 0 -1 10810
box -12 -8 112 252
use MUX2X1  _3587_
timestamp 1728304958
transform -1 0 9450 0 1 10810
box -12 -8 131 252
use NAND2X1  _3588_
timestamp 1728304996
transform 1 0 9370 0 -1 11290
box -12 -8 92 252
use NAND3X1  _3589_
timestamp 1728305047
transform 1 0 10070 0 -1 11290
box -12 -8 112 252
use NAND2X1  _3590_
timestamp 1728304996
transform -1 0 10410 0 -1 11290
box -12 -8 92 252
use OAI21X1  _3591_
timestamp 1728305162
transform 1 0 9810 0 1 10810
box -12 -8 112 252
use NAND2X1  _3592_
timestamp 1728304996
transform 1 0 9850 0 -1 11290
box -12 -8 92 252
use NAND2X1  _3593_
timestamp 1728304996
transform -1 0 9690 0 -1 11290
box -12 -8 92 252
use AOI21X1  _3594_
timestamp 1728304211
transform 1 0 10450 0 -1 10330
box -12 -8 112 252
use NAND2X1  _3595_
timestamp 1728304996
transform 1 0 11030 0 1 10330
box -12 -8 92 252
use AOI22X1  _3596_
timestamp 1728304278
transform -1 0 11090 0 -1 10330
box -14 -8 132 252
use OAI21X1  _3597_
timestamp 1728305162
transform 1 0 10610 0 -1 9370
box -12 -8 112 252
use INVX1  _3598_
timestamp 1728304789
transform 1 0 11270 0 -1 11290
box -12 -8 72 252
use OAI21X1  _3599_
timestamp 1728305162
transform 1 0 11210 0 1 9370
box -12 -8 112 252
use OAI21X1  _3600_
timestamp 1728305162
transform 1 0 11110 0 -1 9370
box -12 -8 112 252
use NAND2X1  _3601_
timestamp 1728304996
transform 1 0 10290 0 -1 8890
box -12 -8 92 252
use OAI21X1  _3602_
timestamp 1728305162
transform 1 0 10510 0 -1 8890
box -12 -8 112 252
use INVX1  _3603_
timestamp 1728304789
transform 1 0 10590 0 1 8890
box -12 -8 72 252
use OAI21X1  _3604_
timestamp 1728305162
transform 1 0 10810 0 1 8890
box -12 -8 112 252
use INVX1  _3605_
timestamp 1728304789
transform 1 0 11270 0 -1 8890
box -12 -8 72 252
use AOI22X1  _3606_
timestamp 1728304278
transform 1 0 10770 0 -1 8890
box -14 -8 132 252
use OAI21X1  _3607_
timestamp 1728305162
transform -1 0 10130 0 1 7450
box -12 -8 112 252
use OAI21X1  _3608_
timestamp 1728305162
transform -1 0 10390 0 1 7450
box -12 -8 112 252
use INVX1  _3609_
timestamp 1728304789
transform 1 0 10810 0 1 7450
box -12 -8 72 252
use NAND2X1  _3610_
timestamp 1728304996
transform 1 0 9610 0 1 7450
box -12 -8 92 252
use AND2X2  _3611_
timestamp 1728304163
transform 1 0 9430 0 1 7930
box -12 -8 112 252
use NAND2X1  _3612_
timestamp 1728304996
transform 1 0 9690 0 1 7930
box -12 -8 92 252
use AOI22X1  _3613_
timestamp 1728304278
transform 1 0 9530 0 -1 7930
box -14 -8 132 252
use OAI21X1  _3614_
timestamp 1728305162
transform -1 0 10030 0 1 7930
box -12 -8 112 252
use OAI21X1  _3615_
timestamp 1728305162
transform -1 0 9890 0 -1 7930
box -12 -8 112 252
use OAI21X1  _3616_
timestamp 1728305162
transform -1 0 9210 0 -1 8410
box -12 -8 112 252
use OAI21X1  _3617_
timestamp 1728305162
transform -1 0 9470 0 -1 8410
box -12 -8 112 252
use NAND2X1  _3618_
timestamp 1728304996
transform 1 0 9850 0 -1 8410
box -12 -8 92 252
use INVX1  _3619_
timestamp 1728304789
transform 1 0 11030 0 -1 7930
box -12 -8 72 252
use AOI22X1  _3620_
timestamp 1728304278
transform -1 0 10850 0 -1 7450
box -14 -8 132 252
use OAI21X1  _3621_
timestamp 1728305162
transform -1 0 10630 0 1 8410
box -12 -8 112 252
use INVX1  _3622_
timestamp 1728304789
transform 1 0 10790 0 1 8410
box -12 -8 72 252
use OAI21X1  _3623_
timestamp 1728305162
transform 1 0 10070 0 -1 8410
box -12 -8 112 252
use INVX1  _3624_
timestamp 1728304789
transform 1 0 10810 0 -1 8410
box -12 -8 72 252
use NAND2X1  _3625_
timestamp 1728304996
transform 1 0 10910 0 1 7930
box -12 -8 92 252
use OAI21X1  _3626_
timestamp 1728305162
transform -1 0 10870 0 -1 7930
box -12 -8 112 252
use NOR2X1  _3627_
timestamp 1728305106
transform -1 0 9850 0 -1 7450
box -12 -8 92 252
use OR2X2  _3628_
timestamp 1728305284
transform -1 0 10590 0 -1 7450
box -12 -8 112 252
use NAND2X1  _3629_
timestamp 1728304996
transform 1 0 10750 0 1 6970
box -12 -8 92 252
use OAI21X1  _3630_
timestamp 1728305162
transform 1 0 10550 0 -1 8410
box -12 -8 112 252
use NAND2X1  _3631_
timestamp 1728304996
transform -1 0 10750 0 1 7930
box -12 -8 92 252
use NAND2X1  _3632_
timestamp 1728304996
transform -1 0 11110 0 -1 11290
box -12 -8 92 252
use OAI21X1  _3633_
timestamp 1728305162
transform 1 0 11010 0 1 10810
box -12 -8 112 252
use NAND2X1  _3634_
timestamp 1728304996
transform -1 0 10870 0 -1 11290
box -12 -8 92 252
use NOR2X1  _3635_
timestamp 1728305106
transform -1 0 10610 0 1 10810
box -12 -8 92 252
use OAI21X1  _3636_
timestamp 1728305162
transform -1 0 10710 0 -1 10810
box -12 -8 112 252
use NAND2X1  _3637_
timestamp 1728304996
transform -1 0 10870 0 1 10330
box -12 -8 92 252
use OAI21X1  _3638_
timestamp 1728305162
transform -1 0 10810 0 -1 10330
box -12 -8 112 252
use OAI21X1  _3639_
timestamp 1728305162
transform -1 0 10630 0 1 10330
box -12 -8 112 252
use INVX1  _3640_
timestamp 1728304789
transform -1 0 11070 0 1 9370
box -12 -8 72 252
use AOI22X1  _3641_
timestamp 1728304278
transform -1 0 10850 0 1 9370
box -14 -8 132 252
use OAI21X1  _3642_
timestamp 1728305162
transform -1 0 11170 0 1 8890
box -12 -8 112 252
use NAND2X1  _3643_
timestamp 1728304996
transform 1 0 11010 0 1 8410
box -12 -8 92 252
use NAND3X1  _3644_
timestamp 1728305047
transform -1 0 10630 0 -1 7930
box -12 -8 112 252
use AND2X2  _3645_
timestamp 1728304163
transform -1 0 10390 0 -1 7930
box -12 -8 112 252
use NAND2X1  _3646_
timestamp 1728304996
transform -1 0 11130 0 -1 8890
box -12 -8 92 252
use NAND2X1  _3647_
timestamp 1728304996
transform 1 0 11150 0 1 250
box -12 -8 92 252
use NAND2X1  _3648_
timestamp 1728304996
transform 1 0 11250 0 1 8410
box -12 -8 92 252
use NAND2X1  _3649_
timestamp 1728304996
transform 1 0 10310 0 -1 8410
box -12 -8 92 252
use NAND2X1  _3650_
timestamp 1728304996
transform 1 0 10450 0 1 7930
box -12 -8 92 252
use AOI21X1  _3651_
timestamp 1728304211
transform 1 0 10550 0 1 7450
box -12 -8 112 252
use AOI22X1  _3652_
timestamp 1728304278
transform -1 0 10590 0 1 6970
box -14 -8 132 252
use OAI21X1  _3653_
timestamp 1728305162
transform 1 0 10730 0 -1 6970
box -12 -8 112 252
use NAND2X1  _3654_
timestamp 1728304996
transform 1 0 8530 0 1 9850
box -12 -8 92 252
use OAI21X1  _3655_
timestamp 1728305162
transform -1 0 8850 0 1 9850
box -12 -8 112 252
use NAND2X1  _3656_
timestamp 1728304996
transform 1 0 8370 0 1 10330
box -12 -8 92 252
use AOI21X1  _3657_
timestamp 1728304211
transform -1 0 8810 0 -1 10810
box -12 -8 112 252
use OAI21X1  _3658_
timestamp 1728305162
transform -1 0 8730 0 -1 11290
box -12 -8 112 252
use OAI21X1  _3659_
timestamp 1728305162
transform -1 0 8470 0 -1 11290
box -12 -8 112 252
use OAI21X1  _3660_
timestamp 1728305162
transform -1 0 8570 0 -1 10810
box -12 -8 112 252
use NAND2X1  _3661_
timestamp 1728304996
transform -1 0 9430 0 1 10330
box -12 -8 92 252
use OAI21X1  _3662_
timestamp 1728305162
transform -1 0 9690 0 1 10330
box -12 -8 112 252
use NAND2X1  _3663_
timestamp 1728304996
transform 1 0 9510 0 -1 10330
box -12 -8 92 252
use OAI21X1  _3664_
timestamp 1728305162
transform -1 0 9850 0 -1 10330
box -12 -8 112 252
use NAND2X1  _3665_
timestamp 1728304996
transform 1 0 8350 0 -1 10330
box -12 -8 92 252
use OAI21X1  _3666_
timestamp 1728305162
transform -1 0 8690 0 -1 10330
box -12 -8 112 252
use NAND2X1  _3667_
timestamp 1728304996
transform -1 0 9390 0 -1 7930
box -12 -8 92 252
use NOR2X1  _3668_
timestamp 1728305106
transform -1 0 10590 0 1 9370
box -12 -8 92 252
use OAI21X1  _3669_
timestamp 1728305162
transform -1 0 10370 0 1 9370
box -12 -8 112 252
use OAI21X1  _3670_
timestamp 1728305162
transform -1 0 10110 0 1 9370
box -12 -8 112 252
use NAND2X1  _3671_
timestamp 1728304996
transform 1 0 8410 0 1 7450
box -12 -8 92 252
use OAI21X1  _3672_
timestamp 1728305162
transform 1 0 8650 0 1 7450
box -12 -8 112 252
use NAND2X1  _3673_
timestamp 1728304996
transform -1 0 9610 0 -1 7450
box -12 -8 92 252
use OAI21X1  _3674_
timestamp 1728305162
transform -1 0 10110 0 -1 7450
box -12 -8 112 252
use NAND2X1  _3675_
timestamp 1728304996
transform 1 0 10250 0 1 6970
box -12 -8 92 252
use OAI21X1  _3676_
timestamp 1728305162
transform -1 0 10350 0 -1 6970
box -12 -8 112 252
use NAND2X1  _3677_
timestamp 1728304996
transform 1 0 9530 0 1 6970
box -12 -8 92 252
use OAI21X1  _3678_
timestamp 1728305162
transform -1 0 9430 0 -1 6970
box -12 -8 112 252
use DFFSR  _3679_
timestamp 1728387359
transform 1 0 10850 0 -1 6490
box -12 -8 492 252
use DFFSR  _3680_
timestamp 1728387359
transform 1 0 10630 0 1 6490
box -12 -8 492 252
use DFFSR  _3681_
timestamp 1728387359
transform -1 0 8790 0 -1 9850
box -12 -8 492 252
use DFFSR  _3682_
timestamp 1728387359
transform -1 0 8330 0 -1 10810
box -12 -8 492 252
use DFFSR  _3683_
timestamp 1728387359
transform -1 0 9770 0 -1 10810
box -12 -8 492 252
use DFFSR  _3684_
timestamp 1728387359
transform -1 0 9850 0 1 9850
box -12 -8 492 252
use DFFSR  _3685_
timestamp 1728387359
transform -1 0 8930 0 1 10330
box -12 -8 492 252
use DFFSR  _3686_
timestamp 1728387359
transform -1 0 9870 0 1 9370
box -12 -8 492 252
use DFFSR  _3687_
timestamp 1728387359
transform -1 0 8670 0 -1 7450
box -12 -8 492 252
use DFFSR  _3688_
timestamp 1728387359
transform -1 0 10090 0 1 6970
box -12 -8 492 252
use DFFSR  _3689_
timestamp 1728387359
transform -1 0 10850 0 1 6010
box -12 -8 492 252
use DFFSR  _3690_
timestamp 1728387359
transform 1 0 9430 0 -1 6970
box -12 -8 492 252
use BUFX2  _3691_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304320
transform 1 0 7850 0 1 250
box -12 -8 92 252
use BUFX2  _3692_
timestamp 1728304320
transform -1 0 8170 0 1 250
box -12 -8 92 252
use BUFX2  _3693_
timestamp 1728304320
transform -1 0 2130 0 -1 10330
box -12 -8 92 252
use BUFX2  _3694_
timestamp 1728304320
transform -1 0 250 0 -1 10330
box -12 -8 92 252
use BUFX2  _3695_
timestamp 1728304320
transform 1 0 690 0 -1 10330
box -12 -8 92 252
use BUFX2  _3696_
timestamp 1728304320
transform -1 0 230 0 1 9850
box -12 -8 92 252
use BUFX2  _3697_
timestamp 1728304320
transform -1 0 250 0 -1 10810
box -12 -8 92 252
use BUFX2  _3698_
timestamp 1728304320
transform -1 0 470 0 -1 10810
box -12 -8 92 252
use BUFX2  _3699_
timestamp 1728304320
transform 1 0 6250 0 1 1210
box -12 -8 92 252
use BUFX2  _3700_
timestamp 1728304320
transform -1 0 6470 0 -1 730
box -12 -8 92 252
use BUFX2  _3701_
timestamp 1728304320
transform -1 0 6430 0 1 250
box -12 -8 92 252
use BUFX2  _3702_
timestamp 1728304320
transform -1 0 5430 0 1 5050
box -12 -8 92 252
use BUFX2  _3703_
timestamp 1728304320
transform -1 0 3670 0 -1 250
box -12 -8 92 252
use BUFX2  _3704_
timestamp 1728304320
transform -1 0 3430 0 -1 250
box -12 -8 92 252
use BUFX2  _3705_
timestamp 1728304320
transform -1 0 250 0 1 8890
box -12 -8 92 252
use BUFX2  _3706_
timestamp 1728304320
transform -1 0 1470 0 -1 10330
box -12 -8 92 252
use BUFX2  _3707_
timestamp 1728304320
transform 1 0 11250 0 1 6970
box -12 -8 92 252
use BUFX2  _3708_
timestamp 1728304320
transform 1 0 11250 0 -1 7450
box -12 -8 92 252
use BUFX2  _3709_
timestamp 1728304320
transform 1 0 11250 0 1 7450
box -12 -8 92 252
use BUFX2  _3710_
timestamp 1728304320
transform 1 0 11030 0 1 7450
box -12 -8 92 252
use BUFX2  _3711_
timestamp 1728304320
transform 1 0 11230 0 -1 7930
box -12 -8 92 252
use BUFX2  _3712_
timestamp 1728304320
transform 1 0 11030 0 -1 8410
box -12 -8 92 252
use BUFX2  _3713_
timestamp 1728304320
transform 1 0 11150 0 1 7930
box -12 -8 92 252
use BUFX2  _3714_
timestamp 1728304320
transform 1 0 11250 0 -1 8410
box -12 -8 92 252
use BUFX2  _3715_
timestamp 1728304320
transform 1 0 11250 0 -1 5530
box -12 -8 92 252
use BUFX2  BUFX2_insert0
timestamp 1728304320
transform 1 0 7890 0 1 10810
box -12 -8 92 252
use BUFX2  BUFX2_insert1
timestamp 1728304320
transform 1 0 9110 0 1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert2
timestamp 1728304320
transform 1 0 9290 0 1 6970
box -12 -8 92 252
use BUFX2  BUFX2_insert3
timestamp 1728304320
transform 1 0 5790 0 -1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert4
timestamp 1728304320
transform 1 0 6890 0 1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert5
timestamp 1728304320
transform -1 0 4190 0 -1 11290
box -12 -8 92 252
use BUFX2  BUFX2_insert6
timestamp 1728304320
transform 1 0 7310 0 1 10330
box -12 -8 92 252
use BUFX2  BUFX2_insert7
timestamp 1728304320
transform -1 0 4270 0 1 4090
box -12 -8 92 252
use BUFX2  BUFX2_insert8
timestamp 1728304320
transform -1 0 7730 0 -1 2170
box -12 -8 92 252
use BUFX2  BUFX2_insert9
timestamp 1728304320
transform 1 0 4590 0 -1 11290
box -12 -8 92 252
use BUFX2  BUFX2_insert10
timestamp 1728304320
transform -1 0 750 0 1 4090
box -12 -8 92 252
use BUFX2  BUFX2_insert11
timestamp 1728304320
transform -1 0 4970 0 1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert12
timestamp 1728304320
transform 1 0 850 0 1 5530
box -12 -8 92 252
use BUFX2  BUFX2_insert13
timestamp 1728304320
transform -1 0 6070 0 1 7450
box -12 -8 92 252
use BUFX2  BUFX2_insert14
timestamp 1728304320
transform 1 0 4650 0 1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert15
timestamp 1728304320
transform 1 0 5710 0 -1 5050
box -12 -8 92 252
use BUFX2  BUFX2_insert16
timestamp 1728304320
transform 1 0 2810 0 1 8410
box -12 -8 92 252
use BUFX2  BUFX2_insert17
timestamp 1728304320
transform 1 0 4310 0 1 6490
box -12 -8 92 252
use BUFX2  BUFX2_insert18
timestamp 1728304320
transform -1 0 230 0 1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert19
timestamp 1728304320
transform -1 0 510 0 1 8410
box -12 -8 92 252
use BUFX2  BUFX2_insert20
timestamp 1728304320
transform 1 0 630 0 -1 7930
box -12 -8 92 252
use BUFX2  BUFX2_insert21
timestamp 1728304320
transform -1 0 7250 0 1 4570
box -12 -8 92 252
use BUFX2  BUFX2_insert22
timestamp 1728304320
transform -1 0 10630 0 1 4090
box -12 -8 92 252
use BUFX2  BUFX2_insert23
timestamp 1728304320
transform -1 0 8950 0 1 4090
box -12 -8 92 252
use BUFX2  BUFX2_insert24
timestamp 1728304320
transform 1 0 8630 0 1 3130
box -12 -8 92 252
use BUFX2  BUFX2_insert25
timestamp 1728304320
transform -1 0 7250 0 1 3130
box -12 -8 92 252
use BUFX2  BUFX2_insert37
timestamp 1728304320
transform -1 0 1170 0 1 5530
box -12 -8 92 252
use BUFX2  BUFX2_insert38
timestamp 1728304320
transform 1 0 1390 0 1 4570
box -12 -8 92 252
use BUFX2  BUFX2_insert39
timestamp 1728304320
transform -1 0 1190 0 -1 6010
box -12 -8 92 252
use BUFX2  BUFX2_insert40
timestamp 1728304320
transform -1 0 2910 0 -1 6010
box -12 -8 92 252
use BUFX2  BUFX2_insert41
timestamp 1728304320
transform 1 0 9630 0 -1 3130
box -12 -8 92 252
use BUFX2  BUFX2_insert42
timestamp 1728304320
transform 1 0 8970 0 -1 3130
box -12 -8 92 252
use BUFX2  BUFX2_insert43
timestamp 1728304320
transform -1 0 8950 0 -1 3610
box -12 -8 92 252
use BUFX2  BUFX2_insert44
timestamp 1728304320
transform -1 0 9150 0 1 4570
box -12 -8 92 252
use BUFX2  BUFX2_insert45
timestamp 1728304320
transform 1 0 3970 0 1 4090
box -12 -8 92 252
use BUFX2  BUFX2_insert46
timestamp 1728304320
transform 1 0 5330 0 1 4090
box -12 -8 92 252
use BUFX2  BUFX2_insert47
timestamp 1728304320
transform 1 0 4410 0 1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert48
timestamp 1728304320
transform 1 0 5550 0 -1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert49
timestamp 1728304320
transform -1 0 2390 0 1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert50
timestamp 1728304320
transform 1 0 8430 0 -1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert51
timestamp 1728304320
transform -1 0 10590 0 1 4570
box -12 -8 92 252
use BUFX2  BUFX2_insert52
timestamp 1728304320
transform -1 0 9610 0 1 4570
box -12 -8 92 252
use BUFX2  BUFX2_insert53
timestamp 1728304320
transform -1 0 9710 0 -1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert54
timestamp 1728304320
transform -1 0 8550 0 -1 3130
box -12 -8 92 252
use BUFX2  BUFX2_insert55
timestamp 1728304320
transform -1 0 490 0 1 730
box -12 -8 92 252
use BUFX2  BUFX2_insert56
timestamp 1728304320
transform 1 0 5130 0 -1 1210
box -12 -8 92 252
use BUFX2  BUFX2_insert57
timestamp 1728304320
transform 1 0 4710 0 -1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert58
timestamp 1728304320
transform 1 0 2050 0 1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert59
timestamp 1728304320
transform 1 0 4490 0 1 730
box -12 -8 92 252
use BUFX2  BUFX2_insert60
timestamp 1728304320
transform -1 0 8910 0 -1 10330
box -12 -8 92 252
use BUFX2  BUFX2_insert61
timestamp 1728304320
transform 1 0 10270 0 -1 7450
box -12 -8 92 252
use BUFX2  BUFX2_insert62
timestamp 1728304320
transform 1 0 9290 0 -1 10330
box -12 -8 92 252
use BUFX2  BUFX2_insert63
timestamp 1728304320
transform 1 0 9390 0 1 7450
box -12 -8 92 252
use BUFX2  BUFX2_insert64
timestamp 1728304320
transform 1 0 8730 0 1 1210
box -12 -8 92 252
use BUFX2  BUFX2_insert65
timestamp 1728304320
transform -1 0 5170 0 1 4090
box -12 -8 92 252
use BUFX2  BUFX2_insert66
timestamp 1728304320
transform 1 0 5870 0 1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert67
timestamp 1728304320
transform 1 0 6710 0 1 5050
box -12 -8 92 252
use BUFX2  BUFX2_insert68
timestamp 1728304320
transform 1 0 7690 0 -1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert69
timestamp 1728304320
transform -1 0 6250 0 1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert70
timestamp 1728304320
transform 1 0 8850 0 -1 2170
box -12 -8 92 252
use BUFX2  BUFX2_insert71
timestamp 1728304320
transform 1 0 2570 0 -1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert72
timestamp 1728304320
transform 1 0 4010 0 1 1210
box -12 -8 92 252
use BUFX2  BUFX2_insert73
timestamp 1728304320
transform 1 0 2790 0 1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert74
timestamp 1728304320
transform -1 0 3870 0 -1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert75
timestamp 1728304320
transform -1 0 950 0 1 2170
box -12 -8 92 252
use BUFX2  BUFX2_insert76
timestamp 1728304320
transform 1 0 8850 0 1 4570
box -12 -8 92 252
use BUFX2  BUFX2_insert77
timestamp 1728304320
transform -1 0 8670 0 -1 5530
box -12 -8 92 252
use BUFX2  BUFX2_insert78
timestamp 1728304320
transform 1 0 9050 0 -1 5530
box -12 -8 92 252
use BUFX2  BUFX2_insert79
timestamp 1728304320
transform -1 0 9390 0 1 4570
box -12 -8 92 252
use BUFX2  BUFX2_insert80
timestamp 1728304320
transform 1 0 4310 0 -1 6490
box -12 -8 92 252
use BUFX2  BUFX2_insert81
timestamp 1728304320
transform 1 0 3430 0 -1 7930
box -12 -8 92 252
use BUFX2  BUFX2_insert82
timestamp 1728304320
transform 1 0 2310 0 -1 7930
box -12 -8 92 252
use BUFX2  BUFX2_insert83
timestamp 1728304320
transform -1 0 2850 0 -1 7930
box -12 -8 92 252
use CLKBUF1  CLKBUF1_insert26 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304421
transform -1 0 1690 0 1 3130
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert27
timestamp 1728304421
transform 1 0 3770 0 1 3130
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert28
timestamp 1728304421
transform 1 0 150 0 1 3130
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert29
timestamp 1728304421
transform 1 0 650 0 1 7930
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert30
timestamp 1728304421
transform 1 0 8330 0 1 5530
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert31
timestamp 1728304421
transform -1 0 7850 0 -1 10810
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert32
timestamp 1728304421
transform -1 0 3490 0 -1 4570
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert33
timestamp 1728304421
transform -1 0 8210 0 1 10330
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert34
timestamp 1728304421
transform -1 0 370 0 -1 11290
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert35
timestamp 1728304421
transform -1 0 5790 0 1 5050
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert36
timestamp 1728304421
transform -1 0 3150 0 -1 6490
box -12 -8 212 252
use FILL  FILL167250x144150 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728341909
transform -1 0 11170 0 -1 9850
box -12 -8 32 252
use FILL  FILL167550x75750
timestamp 1728341909
transform 1 0 11170 0 1 5050
box -12 -8 32 252
use FILL  FILL167550x133350
timestamp 1728341909
transform 1 0 11170 0 1 8890
box -12 -8 32 252
use FILL  FILL167550x144150
timestamp 1728341909
transform -1 0 11190 0 -1 9850
box -12 -8 32 252
use FILL  FILL167850x61350
timestamp 1728341909
transform 1 0 11190 0 1 4090
box -12 -8 32 252
use FILL  FILL167850x64950
timestamp 1728341909
transform -1 0 11210 0 -1 4570
box -12 -8 32 252
use FILL  FILL167850x75750
timestamp 1728341909
transform 1 0 11190 0 1 5050
box -12 -8 32 252
use FILL  FILL167850x133350
timestamp 1728341909
transform 1 0 11190 0 1 8890
box -12 -8 32 252
use FILL  FILL167850x144150
timestamp 1728341909
transform -1 0 11210 0 -1 9850
box -12 -8 32 252
use FILL  FILL168150x150
timestamp 1728341909
transform -1 0 11230 0 -1 250
box -12 -8 32 252
use FILL  FILL168150x32550
timestamp 1728341909
transform 1 0 11210 0 1 2170
box -12 -8 32 252
use FILL  FILL168150x39750
timestamp 1728341909
transform 1 0 11210 0 1 2650
box -12 -8 32 252
use FILL  FILL168150x61350
timestamp 1728341909
transform 1 0 11210 0 1 4090
box -12 -8 32 252
use FILL  FILL168150x64950
timestamp 1728341909
transform -1 0 11230 0 -1 4570
box -12 -8 32 252
use FILL  FILL168150x75750
timestamp 1728341909
transform 1 0 11210 0 1 5050
box -12 -8 32 252
use FILL  FILL168150x133350
timestamp 1728341909
transform 1 0 11210 0 1 8890
box -12 -8 32 252
use FILL  FILL168150x136950
timestamp 1728341909
transform -1 0 11230 0 -1 9370
box -12 -8 32 252
use FILL  FILL168150x144150
timestamp 1728341909
transform -1 0 11230 0 -1 9850
box -12 -8 32 252
use FILL  FILL168150x158550
timestamp 1728341909
transform -1 0 11230 0 -1 10810
box -12 -8 32 252
use FILL  FILL168450x150
timestamp 1728341909
transform -1 0 11250 0 -1 250
box -12 -8 32 252
use FILL  FILL168450x3750
timestamp 1728341909
transform 1 0 11230 0 1 250
box -12 -8 32 252
use FILL  FILL168450x14550
timestamp 1728341909
transform -1 0 11250 0 -1 1210
box -12 -8 32 252
use FILL  FILL168450x18150
timestamp 1728341909
transform 1 0 11230 0 1 1210
box -12 -8 32 252
use FILL  FILL168450x32550
timestamp 1728341909
transform 1 0 11230 0 1 2170
box -12 -8 32 252
use FILL  FILL168450x39750
timestamp 1728341909
transform 1 0 11230 0 1 2650
box -12 -8 32 252
use FILL  FILL168450x57750
timestamp 1728341909
transform -1 0 11250 0 -1 4090
box -12 -8 32 252
use FILL  FILL168450x61350
timestamp 1728341909
transform 1 0 11230 0 1 4090
box -12 -8 32 252
use FILL  FILL168450x64950
timestamp 1728341909
transform -1 0 11250 0 -1 4570
box -12 -8 32 252
use FILL  FILL168450x75750
timestamp 1728341909
transform 1 0 11230 0 1 5050
box -12 -8 32 252
use FILL  FILL168450x118950
timestamp 1728341909
transform 1 0 11230 0 1 7930
box -12 -8 32 252
use FILL  FILL168450x133350
timestamp 1728341909
transform 1 0 11230 0 1 8890
box -12 -8 32 252
use FILL  FILL168450x136950
timestamp 1728341909
transform -1 0 11250 0 -1 9370
box -12 -8 32 252
use FILL  FILL168450x144150
timestamp 1728341909
transform -1 0 11250 0 -1 9850
box -12 -8 32 252
use FILL  FILL168450x158550
timestamp 1728341909
transform -1 0 11250 0 -1 10810
box -12 -8 32 252
use FILL  FILL168750x150
timestamp 1728341909
transform -1 0 11270 0 -1 250
box -12 -8 32 252
use FILL  FILL168750x3750
timestamp 1728341909
transform 1 0 11250 0 1 250
box -12 -8 32 252
use FILL  FILL168750x14550
timestamp 1728341909
transform -1 0 11270 0 -1 1210
box -12 -8 32 252
use FILL  FILL168750x18150
timestamp 1728341909
transform 1 0 11250 0 1 1210
box -12 -8 32 252
use FILL  FILL168750x32550
timestamp 1728341909
transform 1 0 11250 0 1 2170
box -12 -8 32 252
use FILL  FILL168750x39750
timestamp 1728341909
transform 1 0 11250 0 1 2650
box -12 -8 32 252
use FILL  FILL168750x57750
timestamp 1728341909
transform -1 0 11270 0 -1 4090
box -12 -8 32 252
use FILL  FILL168750x61350
timestamp 1728341909
transform 1 0 11250 0 1 4090
box -12 -8 32 252
use FILL  FILL168750x64950
timestamp 1728341909
transform -1 0 11270 0 -1 4570
box -12 -8 32 252
use FILL  FILL168750x75750
timestamp 1728341909
transform 1 0 11250 0 1 5050
box -12 -8 32 252
use FILL  FILL168750x118950
timestamp 1728341909
transform 1 0 11250 0 1 7930
box -12 -8 32 252
use FILL  FILL168750x133350
timestamp 1728341909
transform 1 0 11250 0 1 8890
box -12 -8 32 252
use FILL  FILL168750x136950
timestamp 1728341909
transform -1 0 11270 0 -1 9370
box -12 -8 32 252
use FILL  FILL168750x144150
timestamp 1728341909
transform -1 0 11270 0 -1 9850
box -12 -8 32 252
use FILL  FILL168750x158550
timestamp 1728341909
transform -1 0 11270 0 -1 10810
box -12 -8 32 252
use FILL  FILL169050x150
timestamp 1728341909
transform -1 0 11290 0 -1 250
box -12 -8 32 252
use FILL  FILL169050x3750
timestamp 1728341909
transform 1 0 11270 0 1 250
box -12 -8 32 252
use FILL  FILL169050x14550
timestamp 1728341909
transform -1 0 11290 0 -1 1210
box -12 -8 32 252
use FILL  FILL169050x18150
timestamp 1728341909
transform 1 0 11270 0 1 1210
box -12 -8 32 252
use FILL  FILL169050x32550
timestamp 1728341909
transform 1 0 11270 0 1 2170
box -12 -8 32 252
use FILL  FILL169050x39750
timestamp 1728341909
transform 1 0 11270 0 1 2650
box -12 -8 32 252
use FILL  FILL169050x57750
timestamp 1728341909
transform -1 0 11290 0 -1 4090
box -12 -8 32 252
use FILL  FILL169050x61350
timestamp 1728341909
transform 1 0 11270 0 1 4090
box -12 -8 32 252
use FILL  FILL169050x64950
timestamp 1728341909
transform -1 0 11290 0 -1 4570
box -12 -8 32 252
use FILL  FILL169050x75750
timestamp 1728341909
transform 1 0 11270 0 1 5050
box -12 -8 32 252
use FILL  FILL169050x118950
timestamp 1728341909
transform 1 0 11270 0 1 7930
box -12 -8 32 252
use FILL  FILL169050x133350
timestamp 1728341909
transform 1 0 11270 0 1 8890
box -12 -8 32 252
use FILL  FILL169050x136950
timestamp 1728341909
transform -1 0 11290 0 -1 9370
box -12 -8 32 252
use FILL  FILL169050x144150
timestamp 1728341909
transform -1 0 11290 0 -1 9850
box -12 -8 32 252
use FILL  FILL169050x158550
timestamp 1728341909
transform -1 0 11290 0 -1 10810
box -12 -8 32 252
use FILL  FILL169350x150
timestamp 1728341909
transform -1 0 11310 0 -1 250
box -12 -8 32 252
use FILL  FILL169350x3750
timestamp 1728341909
transform 1 0 11290 0 1 250
box -12 -8 32 252
use FILL  FILL169350x7350
timestamp 1728341909
transform -1 0 11310 0 -1 730
box -12 -8 32 252
use FILL  FILL169350x14550
timestamp 1728341909
transform -1 0 11310 0 -1 1210
box -12 -8 32 252
use FILL  FILL169350x18150
timestamp 1728341909
transform 1 0 11290 0 1 1210
box -12 -8 32 252
use FILL  FILL169350x32550
timestamp 1728341909
transform 1 0 11290 0 1 2170
box -12 -8 32 252
use FILL  FILL169350x39750
timestamp 1728341909
transform 1 0 11290 0 1 2650
box -12 -8 32 252
use FILL  FILL169350x57750
timestamp 1728341909
transform -1 0 11310 0 -1 4090
box -12 -8 32 252
use FILL  FILL169350x61350
timestamp 1728341909
transform 1 0 11290 0 1 4090
box -12 -8 32 252
use FILL  FILL169350x64950
timestamp 1728341909
transform -1 0 11310 0 -1 4570
box -12 -8 32 252
use FILL  FILL169350x75750
timestamp 1728341909
transform 1 0 11290 0 1 5050
box -12 -8 32 252
use FILL  FILL169350x82950
timestamp 1728341909
transform 1 0 11290 0 1 5530
box -12 -8 32 252
use FILL  FILL169350x118950
timestamp 1728341909
transform 1 0 11290 0 1 7930
box -12 -8 32 252
use FILL  FILL169350x133350
timestamp 1728341909
transform 1 0 11290 0 1 8890
box -12 -8 32 252
use FILL  FILL169350x136950
timestamp 1728341909
transform -1 0 11310 0 -1 9370
box -12 -8 32 252
use FILL  FILL169350x144150
timestamp 1728341909
transform -1 0 11310 0 -1 9850
box -12 -8 32 252
use FILL  FILL169350x158550
timestamp 1728341909
transform -1 0 11310 0 -1 10810
box -12 -8 32 252
use FILL  FILL169650x150
timestamp 1728341909
transform -1 0 11330 0 -1 250
box -12 -8 32 252
use FILL  FILL169650x3750
timestamp 1728341909
transform 1 0 11310 0 1 250
box -12 -8 32 252
use FILL  FILL169650x7350
timestamp 1728341909
transform -1 0 11330 0 -1 730
box -12 -8 32 252
use FILL  FILL169650x10950
timestamp 1728341909
transform 1 0 11310 0 1 730
box -12 -8 32 252
use FILL  FILL169650x14550
timestamp 1728341909
transform -1 0 11330 0 -1 1210
box -12 -8 32 252
use FILL  FILL169650x18150
timestamp 1728341909
transform 1 0 11310 0 1 1210
box -12 -8 32 252
use FILL  FILL169650x32550
timestamp 1728341909
transform 1 0 11310 0 1 2170
box -12 -8 32 252
use FILL  FILL169650x39750
timestamp 1728341909
transform 1 0 11310 0 1 2650
box -12 -8 32 252
use FILL  FILL169650x57750
timestamp 1728341909
transform -1 0 11330 0 -1 4090
box -12 -8 32 252
use FILL  FILL169650x61350
timestamp 1728341909
transform 1 0 11310 0 1 4090
box -12 -8 32 252
use FILL  FILL169650x64950
timestamp 1728341909
transform -1 0 11330 0 -1 4570
box -12 -8 32 252
use FILL  FILL169650x75750
timestamp 1728341909
transform 1 0 11310 0 1 5050
box -12 -8 32 252
use FILL  FILL169650x82950
timestamp 1728341909
transform 1 0 11310 0 1 5530
box -12 -8 32 252
use FILL  FILL169650x100950
timestamp 1728341909
transform -1 0 11330 0 -1 6970
box -12 -8 32 252
use FILL  FILL169650x115350
timestamp 1728341909
transform -1 0 11330 0 -1 7930
box -12 -8 32 252
use FILL  FILL169650x118950
timestamp 1728341909
transform 1 0 11310 0 1 7930
box -12 -8 32 252
use FILL  FILL169650x133350
timestamp 1728341909
transform 1 0 11310 0 1 8890
box -12 -8 32 252
use FILL  FILL169650x136950
timestamp 1728341909
transform -1 0 11330 0 -1 9370
box -12 -8 32 252
use FILL  FILL169650x140550
timestamp 1728341909
transform 1 0 11310 0 1 9370
box -12 -8 32 252
use FILL  FILL169650x144150
timestamp 1728341909
transform -1 0 11330 0 -1 9850
box -12 -8 32 252
use FILL  FILL169650x158550
timestamp 1728341909
transform -1 0 11330 0 -1 10810
box -12 -8 32 252
use FILL  FILL169950x150
timestamp 1728341909
transform -1 0 11350 0 -1 250
box -12 -8 32 252
use FILL  FILL169950x3750
timestamp 1728341909
transform 1 0 11330 0 1 250
box -12 -8 32 252
use FILL  FILL169950x7350
timestamp 1728341909
transform -1 0 11350 0 -1 730
box -12 -8 32 252
use FILL  FILL169950x10950
timestamp 1728341909
transform 1 0 11330 0 1 730
box -12 -8 32 252
use FILL  FILL169950x14550
timestamp 1728341909
transform -1 0 11350 0 -1 1210
box -12 -8 32 252
use FILL  FILL169950x18150
timestamp 1728341909
transform 1 0 11330 0 1 1210
box -12 -8 32 252
use FILL  FILL169950x21750
timestamp 1728341909
transform -1 0 11350 0 -1 1690
box -12 -8 32 252
use FILL  FILL169950x25350
timestamp 1728341909
transform 1 0 11330 0 1 1690
box -12 -8 32 252
use FILL  FILL169950x28950
timestamp 1728341909
transform -1 0 11350 0 -1 2170
box -12 -8 32 252
use FILL  FILL169950x32550
timestamp 1728341909
transform 1 0 11330 0 1 2170
box -12 -8 32 252
use FILL  FILL169950x36150
timestamp 1728341909
transform -1 0 11350 0 -1 2650
box -12 -8 32 252
use FILL  FILL169950x39750
timestamp 1728341909
transform 1 0 11330 0 1 2650
box -12 -8 32 252
use FILL  FILL169950x43350
timestamp 1728341909
transform -1 0 11350 0 -1 3130
box -12 -8 32 252
use FILL  FILL169950x50550
timestamp 1728341909
transform -1 0 11350 0 -1 3610
box -12 -8 32 252
use FILL  FILL169950x57750
timestamp 1728341909
transform -1 0 11350 0 -1 4090
box -12 -8 32 252
use FILL  FILL169950x61350
timestamp 1728341909
transform 1 0 11330 0 1 4090
box -12 -8 32 252
use FILL  FILL169950x64950
timestamp 1728341909
transform -1 0 11350 0 -1 4570
box -12 -8 32 252
use FILL  FILL169950x72150
timestamp 1728341909
transform -1 0 11350 0 -1 5050
box -12 -8 32 252
use FILL  FILL169950x75750
timestamp 1728341909
transform 1 0 11330 0 1 5050
box -12 -8 32 252
use FILL  FILL169950x79350
timestamp 1728341909
transform -1 0 11350 0 -1 5530
box -12 -8 32 252
use FILL  FILL169950x82950
timestamp 1728341909
transform 1 0 11330 0 1 5530
box -12 -8 32 252
use FILL  FILL169950x86550
timestamp 1728341909
transform -1 0 11350 0 -1 6010
box -12 -8 32 252
use FILL  FILL169950x90150
timestamp 1728341909
transform 1 0 11330 0 1 6010
box -12 -8 32 252
use FILL  FILL169950x93750
timestamp 1728341909
transform -1 0 11350 0 -1 6490
box -12 -8 32 252
use FILL  FILL169950x100950
timestamp 1728341909
transform -1 0 11350 0 -1 6970
box -12 -8 32 252
use FILL  FILL169950x104550
timestamp 1728341909
transform 1 0 11330 0 1 6970
box -12 -8 32 252
use FILL  FILL169950x108150
timestamp 1728341909
transform -1 0 11350 0 -1 7450
box -12 -8 32 252
use FILL  FILL169950x111750
timestamp 1728341909
transform 1 0 11330 0 1 7450
box -12 -8 32 252
use FILL  FILL169950x115350
timestamp 1728341909
transform -1 0 11350 0 -1 7930
box -12 -8 32 252
use FILL  FILL169950x118950
timestamp 1728341909
transform 1 0 11330 0 1 7930
box -12 -8 32 252
use FILL  FILL169950x122550
timestamp 1728341909
transform -1 0 11350 0 -1 8410
box -12 -8 32 252
use FILL  FILL169950x126150
timestamp 1728341909
transform 1 0 11330 0 1 8410
box -12 -8 32 252
use FILL  FILL169950x129750
timestamp 1728341909
transform -1 0 11350 0 -1 8890
box -12 -8 32 252
use FILL  FILL169950x133350
timestamp 1728341909
transform 1 0 11330 0 1 8890
box -12 -8 32 252
use FILL  FILL169950x136950
timestamp 1728341909
transform -1 0 11350 0 -1 9370
box -12 -8 32 252
use FILL  FILL169950x140550
timestamp 1728341909
transform 1 0 11330 0 1 9370
box -12 -8 32 252
use FILL  FILL169950x144150
timestamp 1728341909
transform -1 0 11350 0 -1 9850
box -12 -8 32 252
use FILL  FILL169950x147750
timestamp 1728341909
transform 1 0 11330 0 1 9850
box -12 -8 32 252
use FILL  FILL169950x151350
timestamp 1728341909
transform -1 0 11350 0 -1 10330
box -12 -8 32 252
use FILL  FILL169950x158550
timestamp 1728341909
transform -1 0 11350 0 -1 10810
box -12 -8 32 252
use FILL  FILL169950x162150
timestamp 1728341909
transform 1 0 11330 0 1 10810
box -12 -8 32 252
use FILL  FILL169950x165750
timestamp 1728341909
transform -1 0 11350 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__1744_
timestamp 1728341909
transform -1 0 4410 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__1745_
timestamp 1728341909
transform 1 0 4190 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__1746_
timestamp 1728341909
transform -1 0 4170 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__1747_
timestamp 1728341909
transform -1 0 5630 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__1748_
timestamp 1728341909
transform 1 0 6550 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__1749_
timestamp 1728341909
transform 1 0 6310 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__1750_
timestamp 1728341909
transform 1 0 5150 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__1751_
timestamp 1728341909
transform 1 0 6790 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__1752_
timestamp 1728341909
transform 1 0 5370 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__1753_
timestamp 1728341909
transform 1 0 7510 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__1754_
timestamp 1728341909
transform -1 0 7050 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__1755_
timestamp 1728341909
transform -1 0 7270 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__1756_
timestamp 1728341909
transform -1 0 6350 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1757_
timestamp 1728341909
transform 1 0 7010 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__1758_
timestamp 1728341909
transform 1 0 6770 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__1759_
timestamp 1728341909
transform -1 0 3030 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__1760_
timestamp 1728341909
transform 1 0 2330 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__1761_
timestamp 1728341909
transform 1 0 7250 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__1762_
timestamp 1728341909
transform 1 0 2530 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__1763_
timestamp 1728341909
transform -1 0 8170 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__1764_
timestamp 1728341909
transform -1 0 7990 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__1765_
timestamp 1728341909
transform -1 0 7990 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__1766_
timestamp 1728341909
transform -1 0 7790 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__1767_
timestamp 1728341909
transform -1 0 7790 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__1768_
timestamp 1728341909
transform -1 0 5670 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1769_
timestamp 1728341909
transform 1 0 3110 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1770_
timestamp 1728341909
transform 1 0 10770 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1771_
timestamp 1728341909
transform 1 0 11010 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1772_
timestamp 1728341909
transform 1 0 10750 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1773_
timestamp 1728341909
transform 1 0 10290 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1774_
timestamp 1728341909
transform 1 0 10650 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1775_
timestamp 1728341909
transform -1 0 9470 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1776_
timestamp 1728341909
transform 1 0 9510 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1777_
timestamp 1728341909
transform -1 0 8690 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1778_
timestamp 1728341909
transform -1 0 10890 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1779_
timestamp 1728341909
transform 1 0 10110 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1780_
timestamp 1728341909
transform 1 0 10870 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1781_
timestamp 1728341909
transform -1 0 10890 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1782_
timestamp 1728341909
transform -1 0 11130 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1783_
timestamp 1728341909
transform -1 0 9930 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1784_
timestamp 1728341909
transform 1 0 10510 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1785_
timestamp 1728341909
transform 1 0 10850 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1786_
timestamp 1728341909
transform -1 0 10190 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1787_
timestamp 1728341909
transform 1 0 9190 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1788_
timestamp 1728341909
transform 1 0 10470 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1789_
timestamp 1728341909
transform -1 0 9330 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1790_
timestamp 1728341909
transform -1 0 10690 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1791_
timestamp 1728341909
transform 1 0 10910 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1792_
timestamp 1728341909
transform 1 0 5610 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1793_
timestamp 1728341909
transform 1 0 5330 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1794_
timestamp 1728341909
transform -1 0 4910 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1795_
timestamp 1728341909
transform 1 0 3690 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1796_
timestamp 1728341909
transform 1 0 4150 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1797_
timestamp 1728341909
transform -1 0 4670 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1798_
timestamp 1728341909
transform -1 0 10990 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1799_
timestamp 1728341909
transform -1 0 10890 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1800_
timestamp 1728341909
transform -1 0 10410 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1801_
timestamp 1728341909
transform -1 0 10070 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1802_
timestamp 1728341909
transform 1 0 9950 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1803_
timestamp 1728341909
transform 1 0 10190 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1804_
timestamp 1728341909
transform 1 0 10190 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1805_
timestamp 1728341909
transform -1 0 9990 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1806_
timestamp 1728341909
transform 1 0 9930 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1807_
timestamp 1728341909
transform -1 0 10050 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1808_
timestamp 1728341909
transform -1 0 10350 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1809_
timestamp 1728341909
transform -1 0 11010 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1810_
timestamp 1728341909
transform -1 0 6190 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1811_
timestamp 1728341909
transform -1 0 11090 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1812_
timestamp 1728341909
transform -1 0 10170 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1813_
timestamp 1728341909
transform -1 0 7650 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1814_
timestamp 1728341909
transform -1 0 7490 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1815_
timestamp 1728341909
transform -1 0 10910 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1816_
timestamp 1728341909
transform -1 0 7550 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1817_
timestamp 1728341909
transform 1 0 6670 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1818_
timestamp 1728341909
transform 1 0 6610 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1819_
timestamp 1728341909
transform 1 0 6110 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1820_
timestamp 1728341909
transform 1 0 10310 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1821_
timestamp 1728341909
transform -1 0 6670 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1822_
timestamp 1728341909
transform 1 0 11090 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1823_
timestamp 1728341909
transform -1 0 9950 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1824_
timestamp 1728341909
transform 1 0 7250 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1825_
timestamp 1728341909
transform 1 0 6470 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1826_
timestamp 1728341909
transform 1 0 10890 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1827_
timestamp 1728341909
transform -1 0 7330 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1828_
timestamp 1728341909
transform 1 0 11090 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1829_
timestamp 1728341909
transform -1 0 7350 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1830_
timestamp 1728341909
transform 1 0 7490 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1831_
timestamp 1728341909
transform 1 0 10630 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1832_
timestamp 1728341909
transform 1 0 10610 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1833_
timestamp 1728341909
transform 1 0 7170 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1834_
timestamp 1728341909
transform -1 0 6970 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1835_
timestamp 1728341909
transform -1 0 6410 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1836_
timestamp 1728341909
transform -1 0 5970 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1837_
timestamp 1728341909
transform -1 0 5490 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1838_
timestamp 1728341909
transform 1 0 5210 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1839_
timestamp 1728341909
transform 1 0 5790 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1840_
timestamp 1728341909
transform -1 0 7990 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__1841_
timestamp 1728341909
transform -1 0 4930 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__1842_
timestamp 1728341909
transform -1 0 6790 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1843_
timestamp 1728341909
transform 1 0 7110 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1844_
timestamp 1728341909
transform -1 0 10190 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1845_
timestamp 1728341909
transform 1 0 11090 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1846_
timestamp 1728341909
transform 1 0 11110 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1847_
timestamp 1728341909
transform -1 0 8030 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1848_
timestamp 1728341909
transform 1 0 10630 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1849_
timestamp 1728341909
transform -1 0 10550 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1850_
timestamp 1728341909
transform -1 0 8490 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1851_
timestamp 1728341909
transform -1 0 11110 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1852_
timestamp 1728341909
transform 1 0 9670 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1853_
timestamp 1728341909
transform 1 0 9190 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1854_
timestamp 1728341909
transform 1 0 8990 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1855_
timestamp 1728341909
transform 1 0 8750 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1856_
timestamp 1728341909
transform 1 0 9270 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1857_
timestamp 1728341909
transform 1 0 9050 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1858_
timestamp 1728341909
transform 1 0 7230 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1859_
timestamp 1728341909
transform -1 0 10650 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1860_
timestamp 1728341909
transform 1 0 7030 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1861_
timestamp 1728341909
transform 1 0 7270 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1862_
timestamp 1728341909
transform -1 0 9770 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1863_
timestamp 1728341909
transform 1 0 8510 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1864_
timestamp 1728341909
transform 1 0 9810 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1865_
timestamp 1728341909
transform 1 0 7670 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1866_
timestamp 1728341909
transform -1 0 8850 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1867_
timestamp 1728341909
transform 1 0 9230 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1868_
timestamp 1728341909
transform 1 0 10790 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1869_
timestamp 1728341909
transform 1 0 9250 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1870_
timestamp 1728341909
transform -1 0 9030 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1871_
timestamp 1728341909
transform 1 0 8470 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1872_
timestamp 1728341909
transform 1 0 7750 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1873_
timestamp 1728341909
transform 1 0 6310 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1874_
timestamp 1728341909
transform -1 0 6770 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1875_
timestamp 1728341909
transform -1 0 6530 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1876_
timestamp 1728341909
transform 1 0 6590 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1877_
timestamp 1728341909
transform -1 0 8010 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1878_
timestamp 1728341909
transform -1 0 8270 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1879_
timestamp 1728341909
transform -1 0 8010 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1880_
timestamp 1728341909
transform -1 0 6950 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__1881_
timestamp 1728341909
transform -1 0 6270 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__1882_
timestamp 1728341909
transform 1 0 3430 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__1883_
timestamp 1728341909
transform -1 0 6970 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__1884_
timestamp 1728341909
transform -1 0 6490 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__1885_
timestamp 1728341909
transform 1 0 5770 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1886_
timestamp 1728341909
transform -1 0 6170 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__1887_
timestamp 1728341909
transform 1 0 6790 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__1888_
timestamp 1728341909
transform 1 0 3550 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__1889_
timestamp 1728341909
transform -1 0 5910 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__1890_
timestamp 1728341909
transform 1 0 6370 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__1891_
timestamp 1728341909
transform -1 0 6010 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__1892_
timestamp 1728341909
transform 1 0 5570 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__1893_
timestamp 1728341909
transform 1 0 970 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__1894_
timestamp 1728341909
transform 1 0 5910 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__1895_
timestamp 1728341909
transform 1 0 6790 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__1896_
timestamp 1728341909
transform 1 0 5110 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__1897_
timestamp 1728341909
transform 1 0 5950 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__1898_
timestamp 1728341909
transform 1 0 6370 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__1899_
timestamp 1728341909
transform 1 0 6470 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__1900_
timestamp 1728341909
transform 1 0 490 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1901_
timestamp 1728341909
transform 1 0 7930 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1902_
timestamp 1728341909
transform 1 0 8470 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1903_
timestamp 1728341909
transform 1 0 7830 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1904_
timestamp 1728341909
transform -1 0 9990 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1905_
timestamp 1728341909
transform 1 0 7490 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1906_
timestamp 1728341909
transform 1 0 7470 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1907_
timestamp 1728341909
transform 1 0 8610 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1908_
timestamp 1728341909
transform -1 0 7670 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1909_
timestamp 1728341909
transform 1 0 1770 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1910_
timestamp 1728341909
transform -1 0 9730 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1911_
timestamp 1728341909
transform 1 0 9450 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1912_
timestamp 1728341909
transform 1 0 6070 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1913_
timestamp 1728341909
transform 1 0 10590 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1914_
timestamp 1728341909
transform 1 0 10650 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1915_
timestamp 1728341909
transform -1 0 10210 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1916_
timestamp 1728341909
transform -1 0 5830 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1917_
timestamp 1728341909
transform 1 0 3970 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1918_
timestamp 1728341909
transform -1 0 750 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1919_
timestamp 1728341909
transform -1 0 30 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1920_
timestamp 1728341909
transform 1 0 970 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1921_
timestamp 1728341909
transform -1 0 1150 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1922_
timestamp 1728341909
transform -1 0 890 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1923_
timestamp 1728341909
transform 1 0 490 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1924_
timestamp 1728341909
transform -1 0 4430 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1925_
timestamp 1728341909
transform -1 0 270 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1926_
timestamp 1728341909
transform 1 0 730 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1927_
timestamp 1728341909
transform -1 0 2030 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1928_
timestamp 1728341909
transform -1 0 1550 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1929_
timestamp 1728341909
transform 1 0 230 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1930_
timestamp 1728341909
transform 1 0 610 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1931_
timestamp 1728341909
transform 1 0 490 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1932_
timestamp 1728341909
transform -1 0 510 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1933_
timestamp 1728341909
transform 1 0 490 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1934_
timestamp 1728341909
transform -1 0 510 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1935_
timestamp 1728341909
transform -1 0 1490 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1936_
timestamp 1728341909
transform 1 0 750 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1937_
timestamp 1728341909
transform -1 0 510 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1938_
timestamp 1728341909
transform -1 0 30 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1939_
timestamp 1728341909
transform 1 0 250 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1940_
timestamp 1728341909
transform 1 0 770 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1941_
timestamp 1728341909
transform 1 0 490 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1942_
timestamp 1728341909
transform 1 0 490 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1943_
timestamp 1728341909
transform 1 0 8050 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__1944_
timestamp 1728341909
transform -1 0 7590 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1945_
timestamp 1728341909
transform -1 0 7370 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1946_
timestamp 1728341909
transform 1 0 8390 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1947_
timestamp 1728341909
transform -1 0 7570 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1948_
timestamp 1728341909
transform -1 0 6910 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1949_
timestamp 1728341909
transform -1 0 7150 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1950_
timestamp 1728341909
transform 1 0 8250 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1951_
timestamp 1728341909
transform 1 0 8250 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1952_
timestamp 1728341909
transform 1 0 9770 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1953_
timestamp 1728341909
transform -1 0 8330 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1954_
timestamp 1728341909
transform 1 0 8170 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1955_
timestamp 1728341909
transform 1 0 6370 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1956_
timestamp 1728341909
transform -1 0 7930 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1957_
timestamp 1728341909
transform 1 0 8010 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1958_
timestamp 1728341909
transform 1 0 10370 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1959_
timestamp 1728341909
transform 1 0 7730 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1960_
timestamp 1728341909
transform 1 0 7810 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1961_
timestamp 1728341909
transform 1 0 10630 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1962_
timestamp 1728341909
transform 1 0 10430 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1963_
timestamp 1728341909
transform 1 0 9770 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1964_
timestamp 1728341909
transform -1 0 7310 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1965_
timestamp 1728341909
transform -1 0 7590 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1966_
timestamp 1728341909
transform -1 0 3450 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__1967_
timestamp 1728341909
transform -1 0 6910 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__1968_
timestamp 1728341909
transform 1 0 7450 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__1969_
timestamp 1728341909
transform -1 0 7710 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__1970_
timestamp 1728341909
transform 1 0 1450 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1971_
timestamp 1728341909
transform -1 0 750 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1972_
timestamp 1728341909
transform 1 0 1270 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1973_
timestamp 1728341909
transform 1 0 1530 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1974_
timestamp 1728341909
transform 1 0 8290 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__1975_
timestamp 1728341909
transform 1 0 2910 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__1976_
timestamp 1728341909
transform -1 0 7070 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1977_
timestamp 1728341909
transform -1 0 2770 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__1978_
timestamp 1728341909
transform -1 0 3750 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__1979_
timestamp 1728341909
transform -1 0 6450 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__1980_
timestamp 1728341909
transform 1 0 7710 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__1981_
timestamp 1728341909
transform 1 0 8230 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__1982_
timestamp 1728341909
transform -1 0 2970 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__1983_
timestamp 1728341909
transform 1 0 1650 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1984_
timestamp 1728341909
transform 1 0 1730 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1985_
timestamp 1728341909
transform 1 0 2390 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1986_
timestamp 1728341909
transform -1 0 7070 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__1987_
timestamp 1728341909
transform 1 0 5010 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__1988_
timestamp 1728341909
transform -1 0 4910 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__1989_
timestamp 1728341909
transform 1 0 6670 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__1990_
timestamp 1728341909
transform -1 0 7190 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__1991_
timestamp 1728341909
transform -1 0 1990 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1992_
timestamp 1728341909
transform -1 0 1490 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1993_
timestamp 1728341909
transform -1 0 1770 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1994_
timestamp 1728341909
transform 1 0 2010 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1995_
timestamp 1728341909
transform 1 0 7970 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__1996_
timestamp 1728341909
transform -1 0 2190 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__1997_
timestamp 1728341909
transform -1 0 3910 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__1998_
timestamp 1728341909
transform -1 0 6430 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__1999_
timestamp 1728341909
transform -1 0 8150 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2000_
timestamp 1728341909
transform 1 0 1750 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2001_
timestamp 1728341909
transform 1 0 1230 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2002_
timestamp 1728341909
transform 1 0 1470 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2003_
timestamp 1728341909
transform 1 0 1490 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2004_
timestamp 1728341909
transform 1 0 7770 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2005_
timestamp 1728341909
transform 1 0 1930 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2006_
timestamp 1728341909
transform -1 0 6190 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2007_
timestamp 1728341909
transform 1 0 7470 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2008_
timestamp 1728341909
transform -1 0 7990 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2009_
timestamp 1728341909
transform 1 0 730 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2010_
timestamp 1728341909
transform -1 0 790 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2011_
timestamp 1728341909
transform 1 0 490 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2012_
timestamp 1728341909
transform 1 0 750 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2013_
timestamp 1728341909
transform 1 0 5390 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2014_
timestamp 1728341909
transform 1 0 1690 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2015_
timestamp 1728341909
transform -1 0 3890 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2016_
timestamp 1728341909
transform 1 0 6690 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2017_
timestamp 1728341909
transform -1 0 7230 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2018_
timestamp 1728341909
transform -1 0 1470 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2019_
timestamp 1728341909
transform -1 0 1530 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2020_
timestamp 1728341909
transform 1 0 1710 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2021_
timestamp 1728341909
transform 1 0 1670 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2022_
timestamp 1728341909
transform 1 0 4450 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2023_
timestamp 1728341909
transform 1 0 490 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2024_
timestamp 1728341909
transform 1 0 1390 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2025_
timestamp 1728341909
transform 1 0 2450 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2026_
timestamp 1728341909
transform -1 0 4650 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2027_
timestamp 1728341909
transform 1 0 7150 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2028_
timestamp 1728341909
transform -1 0 7430 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2029_
timestamp 1728341909
transform -1 0 30 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2030_
timestamp 1728341909
transform -1 0 510 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2031_
timestamp 1728341909
transform -1 0 270 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2032_
timestamp 1728341909
transform 1 0 490 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2033_
timestamp 1728341909
transform 1 0 7570 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2034_
timestamp 1728341909
transform 1 0 1170 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2035_
timestamp 1728341909
transform 1 0 2050 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2036_
timestamp 1728341909
transform 1 0 2850 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2037_
timestamp 1728341909
transform -1 0 4050 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2038_
timestamp 1728341909
transform 1 0 7490 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2039_
timestamp 1728341909
transform -1 0 7770 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2040_
timestamp 1728341909
transform -1 0 2890 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2041_
timestamp 1728341909
transform -1 0 510 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2042_
timestamp 1728341909
transform 1 0 1670 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2043_
timestamp 1728341909
transform -1 0 3770 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__2044_
timestamp 1728341909
transform 1 0 5310 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2045_
timestamp 1728341909
transform -1 0 4010 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2046_
timestamp 1728341909
transform 1 0 2810 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2047_
timestamp 1728341909
transform 1 0 2570 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2048_
timestamp 1728341909
transform -1 0 3510 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2049_
timestamp 1728341909
transform -1 0 2910 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2050_
timestamp 1728341909
transform -1 0 2390 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2051_
timestamp 1728341909
transform -1 0 2370 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2052_
timestamp 1728341909
transform -1 0 790 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2053_
timestamp 1728341909
transform -1 0 3350 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2054_
timestamp 1728341909
transform 1 0 3070 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2055_
timestamp 1728341909
transform -1 0 2710 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2056_
timestamp 1728341909
transform 1 0 4330 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2057_
timestamp 1728341909
transform -1 0 3890 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2058_
timestamp 1728341909
transform 1 0 4550 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2059_
timestamp 1728341909
transform -1 0 1910 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2060_
timestamp 1728341909
transform -1 0 3730 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2061_
timestamp 1728341909
transform 1 0 3470 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2062_
timestamp 1728341909
transform -1 0 3490 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2063_
timestamp 1728341909
transform 1 0 2430 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2064_
timestamp 1728341909
transform -1 0 2530 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2065_
timestamp 1728341909
transform -1 0 2330 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2066_
timestamp 1728341909
transform 1 0 2390 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2067_
timestamp 1728341909
transform -1 0 2710 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2068_
timestamp 1728341909
transform -1 0 2950 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2069_
timestamp 1728341909
transform 1 0 2490 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2070_
timestamp 1728341909
transform -1 0 1030 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2071_
timestamp 1728341909
transform -1 0 2750 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2072_
timestamp 1728341909
transform -1 0 2490 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2073_
timestamp 1728341909
transform -1 0 1230 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2074_
timestamp 1728341909
transform 1 0 3170 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2075_
timestamp 1728341909
transform -1 0 2650 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2076_
timestamp 1728341909
transform 1 0 2350 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2077_
timestamp 1728341909
transform -1 0 3210 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2078_
timestamp 1728341909
transform 1 0 2730 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2079_
timestamp 1728341909
transform -1 0 3850 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2080_
timestamp 1728341909
transform 1 0 4070 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2081_
timestamp 1728341909
transform -1 0 3630 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2082_
timestamp 1728341909
transform 1 0 5710 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2083_
timestamp 1728341909
transform -1 0 6450 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2084_
timestamp 1728341909
transform 1 0 9870 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2085_
timestamp 1728341909
transform -1 0 10390 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2086_
timestamp 1728341909
transform 1 0 10410 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2087_
timestamp 1728341909
transform 1 0 10950 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2088_
timestamp 1728341909
transform 1 0 10150 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2089_
timestamp 1728341909
transform -1 0 9450 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2090_
timestamp 1728341909
transform 1 0 10630 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2091_
timestamp 1728341909
transform 1 0 11130 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2092_
timestamp 1728341909
transform -1 0 10090 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2093_
timestamp 1728341909
transform 1 0 10150 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2094_
timestamp 1728341909
transform -1 0 10650 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2095_
timestamp 1728341909
transform 1 0 10710 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2096_
timestamp 1728341909
transform -1 0 11110 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2097_
timestamp 1728341909
transform -1 0 11050 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2098_
timestamp 1728341909
transform 1 0 10130 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2099_
timestamp 1728341909
transform 1 0 10610 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2100_
timestamp 1728341909
transform 1 0 10830 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2101_
timestamp 1728341909
transform 1 0 11070 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2102_
timestamp 1728341909
transform 1 0 3950 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2103_
timestamp 1728341909
transform 1 0 4190 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2104_
timestamp 1728341909
transform 1 0 3810 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2105_
timestamp 1728341909
transform -1 0 1710 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2106_
timestamp 1728341909
transform -1 0 2090 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2107_
timestamp 1728341909
transform -1 0 2610 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2108_
timestamp 1728341909
transform 1 0 1410 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2109_
timestamp 1728341909
transform -1 0 2830 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2110_
timestamp 1728341909
transform 1 0 3050 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2111_
timestamp 1728341909
transform 1 0 5250 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2112_
timestamp 1728341909
transform 1 0 11130 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2113_
timestamp 1728341909
transform -1 0 9710 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2114_
timestamp 1728341909
transform 1 0 9710 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2115_
timestamp 1728341909
transform -1 0 11030 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2116_
timestamp 1728341909
transform -1 0 10970 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2117_
timestamp 1728341909
transform -1 0 10570 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2118_
timestamp 1728341909
transform 1 0 8970 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2119_
timestamp 1728341909
transform -1 0 11050 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2120_
timestamp 1728341909
transform 1 0 10990 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2121_
timestamp 1728341909
transform 1 0 11090 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2122_
timestamp 1728341909
transform 1 0 10790 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2123_
timestamp 1728341909
transform 1 0 10850 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2124_
timestamp 1728341909
transform 1 0 9310 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2125_
timestamp 1728341909
transform 1 0 9430 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2126_
timestamp 1728341909
transform -1 0 9870 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2127_
timestamp 1728341909
transform 1 0 9690 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2128_
timestamp 1728341909
transform 1 0 9650 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2129_
timestamp 1728341909
transform -1 0 8870 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2130_
timestamp 1728341909
transform 1 0 9550 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2131_
timestamp 1728341909
transform 1 0 9650 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2132_
timestamp 1728341909
transform 1 0 10110 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2133_
timestamp 1728341909
transform 1 0 10270 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2134_
timestamp 1728341909
transform -1 0 10050 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2135_
timestamp 1728341909
transform 1 0 10550 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2136_
timestamp 1728341909
transform -1 0 10510 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2137_
timestamp 1728341909
transform 1 0 10750 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2138_
timestamp 1728341909
transform -1 0 10850 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2139_
timestamp 1728341909
transform -1 0 10790 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2140_
timestamp 1728341909
transform -1 0 8270 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2141_
timestamp 1728341909
transform 1 0 8510 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2142_
timestamp 1728341909
transform 1 0 1830 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2143_
timestamp 1728341909
transform -1 0 2870 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2144_
timestamp 1728341909
transform -1 0 5970 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2145_
timestamp 1728341909
transform -1 0 6170 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2146_
timestamp 1728341909
transform 1 0 5470 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2147_
timestamp 1728341909
transform -1 0 6710 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2148_
timestamp 1728341909
transform 1 0 9610 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2149_
timestamp 1728341909
transform 1 0 8690 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2150_
timestamp 1728341909
transform -1 0 8450 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2151_
timestamp 1728341909
transform 1 0 8110 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2152_
timestamp 1728341909
transform -1 0 8950 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2153_
timestamp 1728341909
transform -1 0 9050 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2154_
timestamp 1728341909
transform 1 0 8790 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2155_
timestamp 1728341909
transform 1 0 7950 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2156_
timestamp 1728341909
transform -1 0 8230 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2157_
timestamp 1728341909
transform -1 0 8350 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2158_
timestamp 1728341909
transform 1 0 10270 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2159_
timestamp 1728341909
transform 1 0 5970 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2160_
timestamp 1728341909
transform -1 0 6330 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2161_
timestamp 1728341909
transform 1 0 6530 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2162_
timestamp 1728341909
transform -1 0 7870 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2163_
timestamp 1728341909
transform -1 0 8290 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2164_
timestamp 1728341909
transform 1 0 7050 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2165_
timestamp 1728341909
transform -1 0 7030 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2166_
timestamp 1728341909
transform -1 0 8090 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2167_
timestamp 1728341909
transform -1 0 7790 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2168_
timestamp 1728341909
transform -1 0 8050 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2169_
timestamp 1728341909
transform 1 0 8090 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2170_
timestamp 1728341909
transform -1 0 8310 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2171_
timestamp 1728341909
transform 1 0 8510 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2172_
timestamp 1728341909
transform -1 0 10370 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2173_
timestamp 1728341909
transform 1 0 10110 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2174_
timestamp 1728341909
transform 1 0 4330 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2175_
timestamp 1728341909
transform -1 0 3890 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2176_
timestamp 1728341909
transform -1 0 5350 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2177_
timestamp 1728341909
transform -1 0 6010 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2178_
timestamp 1728341909
transform -1 0 6270 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2179_
timestamp 1728341909
transform 1 0 6310 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2180_
timestamp 1728341909
transform 1 0 7110 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2181_
timestamp 1728341909
transform 1 0 7250 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2182_
timestamp 1728341909
transform -1 0 7110 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2183_
timestamp 1728341909
transform 1 0 6090 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2184_
timestamp 1728341909
transform 1 0 6410 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2185_
timestamp 1728341909
transform -1 0 6550 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2186_
timestamp 1728341909
transform -1 0 8990 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2187_
timestamp 1728341909
transform -1 0 9390 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2188_
timestamp 1728341909
transform 1 0 8990 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2189_
timestamp 1728341909
transform -1 0 8770 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2190_
timestamp 1728341909
transform 1 0 8450 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2191_
timestamp 1728341909
transform 1 0 8690 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2192_
timestamp 1728341909
transform 1 0 7250 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2193_
timestamp 1728341909
transform 1 0 7470 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2194_
timestamp 1728341909
transform -1 0 8590 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2195_
timestamp 1728341909
transform -1 0 8510 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2196_
timestamp 1728341909
transform 1 0 8550 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2197_
timestamp 1728341909
transform 1 0 8590 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2198_
timestamp 1728341909
transform -1 0 7190 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2199_
timestamp 1728341909
transform -1 0 7450 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2200_
timestamp 1728341909
transform 1 0 8970 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2201_
timestamp 1728341909
transform 1 0 8830 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2202_
timestamp 1728341909
transform -1 0 8630 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2203_
timestamp 1728341909
transform 1 0 8350 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2204_
timestamp 1728341909
transform -1 0 8350 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2205_
timestamp 1728341909
transform 1 0 8090 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2206_
timestamp 1728341909
transform -1 0 7970 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2207_
timestamp 1728341909
transform 1 0 8470 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2208_
timestamp 1728341909
transform -1 0 8230 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2209_
timestamp 1728341909
transform -1 0 7750 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2210_
timestamp 1728341909
transform 1 0 2690 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2211_
timestamp 1728341909
transform -1 0 7150 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2212_
timestamp 1728341909
transform -1 0 7410 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2213_
timestamp 1728341909
transform -1 0 7930 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2214_
timestamp 1728341909
transform 1 0 8490 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2215_
timestamp 1728341909
transform 1 0 9190 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2216_
timestamp 1728341909
transform 1 0 9170 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2217_
timestamp 1728341909
transform -1 0 9430 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2218_
timestamp 1728341909
transform 1 0 3870 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2219_
timestamp 1728341909
transform -1 0 2190 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2220_
timestamp 1728341909
transform -1 0 3610 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2221_
timestamp 1728341909
transform 1 0 4050 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2222_
timestamp 1728341909
transform 1 0 4270 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2223_
timestamp 1728341909
transform 1 0 4090 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2224_
timestamp 1728341909
transform -1 0 2770 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2225_
timestamp 1728341909
transform -1 0 5830 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2226_
timestamp 1728341909
transform 1 0 5950 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2227_
timestamp 1728341909
transform -1 0 6930 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2228_
timestamp 1728341909
transform 1 0 6670 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2229_
timestamp 1728341909
transform 1 0 7730 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2230_
timestamp 1728341909
transform -1 0 6130 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2231_
timestamp 1728341909
transform -1 0 6370 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2232_
timestamp 1728341909
transform 1 0 6790 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2233_
timestamp 1728341909
transform 1 0 7370 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2234_
timestamp 1728341909
transform 1 0 7270 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2235_
timestamp 1728341909
transform 1 0 9350 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2236_
timestamp 1728341909
transform 1 0 10410 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2237_
timestamp 1728341909
transform 1 0 9890 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2238_
timestamp 1728341909
transform -1 0 9810 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2239_
timestamp 1728341909
transform -1 0 5770 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2240_
timestamp 1728341909
transform 1 0 2630 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2241_
timestamp 1728341909
transform -1 0 4310 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2242_
timestamp 1728341909
transform -1 0 4530 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2243_
timestamp 1728341909
transform 1 0 3310 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2244_
timestamp 1728341909
transform 1 0 5070 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2245_
timestamp 1728341909
transform 1 0 7210 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2246_
timestamp 1728341909
transform 1 0 7230 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2247_
timestamp 1728341909
transform -1 0 3190 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2248_
timestamp 1728341909
transform 1 0 3370 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2249_
timestamp 1728341909
transform 1 0 5350 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2250_
timestamp 1728341909
transform 1 0 6610 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2251_
timestamp 1728341909
transform 1 0 7130 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2252_
timestamp 1728341909
transform -1 0 9570 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2253_
timestamp 1728341909
transform 1 0 9290 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2254_
timestamp 1728341909
transform 1 0 5570 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2255_
timestamp 1728341909
transform -1 0 6910 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2256_
timestamp 1728341909
transform 1 0 7070 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2257_
timestamp 1728341909
transform -1 0 3010 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2258_
timestamp 1728341909
transform -1 0 2970 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2259_
timestamp 1728341909
transform 1 0 3390 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2260_
timestamp 1728341909
transform 1 0 4570 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2261_
timestamp 1728341909
transform -1 0 5570 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2262_
timestamp 1728341909
transform 1 0 4750 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2263_
timestamp 1728341909
transform 1 0 4810 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2264_
timestamp 1728341909
transform -1 0 6110 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2265_
timestamp 1728341909
transform 1 0 3410 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2266_
timestamp 1728341909
transform 1 0 7450 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2267_
timestamp 1728341909
transform -1 0 5350 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2268_
timestamp 1728341909
transform -1 0 5590 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2269_
timestamp 1728341909
transform 1 0 5350 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2270_
timestamp 1728341909
transform -1 0 6190 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2271_
timestamp 1728341909
transform 1 0 5910 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2272_
timestamp 1728341909
transform 1 0 5510 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2273_
timestamp 1728341909
transform 1 0 5330 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2274_
timestamp 1728341909
transform 1 0 5090 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2275_
timestamp 1728341909
transform 1 0 5570 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2276_
timestamp 1728341909
transform -1 0 6210 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2277_
timestamp 1728341909
transform 1 0 7710 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2278_
timestamp 1728341909
transform -1 0 7650 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2279_
timestamp 1728341909
transform 1 0 6410 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2280_
timestamp 1728341909
transform -1 0 6430 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2281_
timestamp 1728341909
transform -1 0 6190 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2282_
timestamp 1728341909
transform 1 0 6470 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2283_
timestamp 1728341909
transform 1 0 7170 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2284_
timestamp 1728341909
transform 1 0 9130 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2285_
timestamp 1728341909
transform 1 0 9570 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2286_
timestamp 1728341909
transform -1 0 2470 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2287_
timestamp 1728341909
transform -1 0 1730 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2288_
timestamp 1728341909
transform -1 0 2170 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2289_
timestamp 1728341909
transform 1 0 2130 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2290_
timestamp 1728341909
transform -1 0 1690 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2291_
timestamp 1728341909
transform 1 0 1910 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2292_
timestamp 1728341909
transform 1 0 4030 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2293_
timestamp 1728341909
transform 1 0 4770 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2294_
timestamp 1728341909
transform 1 0 5990 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2295_
timestamp 1728341909
transform -1 0 2170 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2296_
timestamp 1728341909
transform 1 0 3610 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2297_
timestamp 1728341909
transform 1 0 2150 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2298_
timestamp 1728341909
transform 1 0 1910 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2299_
timestamp 1728341909
transform 1 0 3370 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2300_
timestamp 1728341909
transform 1 0 3110 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2301_
timestamp 1728341909
transform -1 0 3570 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2302_
timestamp 1728341909
transform 1 0 5050 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2303_
timestamp 1728341909
transform -1 0 5030 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2304_
timestamp 1728341909
transform 1 0 5270 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2305_
timestamp 1728341909
transform -1 0 1470 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2306_
timestamp 1728341909
transform 1 0 2370 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2307_
timestamp 1728341909
transform -1 0 5530 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2308_
timestamp 1728341909
transform -1 0 5530 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2309_
timestamp 1728341909
transform 1 0 4530 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2310_
timestamp 1728341909
transform 1 0 4290 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2311_
timestamp 1728341909
transform -1 0 3690 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2312_
timestamp 1728341909
transform -1 0 3930 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2313_
timestamp 1728341909
transform 1 0 5210 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2314_
timestamp 1728341909
transform 1 0 4390 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2315_
timestamp 1728341909
transform 1 0 5350 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2316_
timestamp 1728341909
transform -1 0 9790 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2317_
timestamp 1728341909
transform 1 0 11090 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2318_
timestamp 1728341909
transform -1 0 10790 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2319_
timestamp 1728341909
transform -1 0 10410 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2320_
timestamp 1728341909
transform 1 0 10570 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2321_
timestamp 1728341909
transform 1 0 10510 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2322_
timestamp 1728341909
transform 1 0 10410 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2323_
timestamp 1728341909
transform 1 0 6670 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2324_
timestamp 1728341909
transform 1 0 6870 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2325_
timestamp 1728341909
transform 1 0 9230 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2326_
timestamp 1728341909
transform -1 0 8770 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2327_
timestamp 1728341909
transform -1 0 9230 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2328_
timestamp 1728341909
transform -1 0 9470 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2329_
timestamp 1728341909
transform 1 0 9190 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2330_
timestamp 1728341909
transform -1 0 8950 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2331_
timestamp 1728341909
transform -1 0 9110 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2332_
timestamp 1728341909
transform 1 0 9090 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2333_
timestamp 1728341909
transform 1 0 9350 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2334_
timestamp 1728341909
transform -1 0 9550 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2335_
timestamp 1728341909
transform 1 0 5590 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2336_
timestamp 1728341909
transform 1 0 6110 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2337_
timestamp 1728341909
transform -1 0 5890 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2338_
timestamp 1728341909
transform -1 0 5830 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2339_
timestamp 1728341909
transform 1 0 10310 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2340_
timestamp 1728341909
transform -1 0 9190 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2341_
timestamp 1728341909
transform 1 0 9190 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2342_
timestamp 1728341909
transform 1 0 10050 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2343_
timestamp 1728341909
transform -1 0 9550 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2344_
timestamp 1728341909
transform 1 0 9650 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2345_
timestamp 1728341909
transform -1 0 6830 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2346_
timestamp 1728341909
transform 1 0 6690 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2347_
timestamp 1728341909
transform -1 0 7030 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2348_
timestamp 1728341909
transform 1 0 8030 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2349_
timestamp 1728341909
transform -1 0 7730 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2350_
timestamp 1728341909
transform 1 0 7450 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2351_
timestamp 1728341909
transform -1 0 5150 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2352_
timestamp 1728341909
transform 1 0 5750 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2353_
timestamp 1728341909
transform -1 0 4170 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2354_
timestamp 1728341909
transform 1 0 4650 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2355_
timestamp 1728341909
transform -1 0 4910 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2356_
timestamp 1728341909
transform 1 0 5850 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2357_
timestamp 1728341909
transform -1 0 5610 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2358_
timestamp 1728341909
transform 1 0 6890 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2359_
timestamp 1728341909
transform 1 0 6250 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2360_
timestamp 1728341909
transform 1 0 6490 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2361_
timestamp 1728341909
transform 1 0 7790 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2362_
timestamp 1728341909
transform 1 0 7310 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2363_
timestamp 1728341909
transform -1 0 7410 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2364_
timestamp 1728341909
transform 1 0 8030 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2365_
timestamp 1728341909
transform -1 0 7910 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2366_
timestamp 1728341909
transform 1 0 7670 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2367_
timestamp 1728341909
transform 1 0 7950 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2368_
timestamp 1728341909
transform 1 0 8170 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2369_
timestamp 1728341909
transform -1 0 9890 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2370_
timestamp 1728341909
transform 1 0 5310 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2371_
timestamp 1728341909
transform -1 0 8710 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2372_
timestamp 1728341909
transform -1 0 8450 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2373_
timestamp 1728341909
transform -1 0 8030 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2374_
timestamp 1728341909
transform 1 0 8030 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2375_
timestamp 1728341909
transform 1 0 6430 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2376_
timestamp 1728341909
transform 1 0 8390 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2377_
timestamp 1728341909
transform -1 0 8650 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2378_
timestamp 1728341909
transform -1 0 8950 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2379_
timestamp 1728341909
transform -1 0 6810 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2380_
timestamp 1728341909
transform -1 0 6950 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2381_
timestamp 1728341909
transform -1 0 6810 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2382_
timestamp 1728341909
transform -1 0 7890 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2383_
timestamp 1728341909
transform 1 0 7610 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2384_
timestamp 1728341909
transform 1 0 7710 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2385_
timestamp 1728341909
transform -1 0 7450 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2386_
timestamp 1728341909
transform -1 0 6570 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2387_
timestamp 1728341909
transform -1 0 6330 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2388_
timestamp 1728341909
transform -1 0 8890 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2389_
timestamp 1728341909
transform -1 0 8270 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2390_
timestamp 1728341909
transform -1 0 8210 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2391_
timestamp 1728341909
transform -1 0 9450 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2392_
timestamp 1728341909
transform 1 0 8210 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2393_
timestamp 1728341909
transform 1 0 8170 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2394_
timestamp 1728341909
transform 1 0 8810 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2395_
timestamp 1728341909
transform 1 0 8770 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2396_
timestamp 1728341909
transform 1 0 9050 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2397_
timestamp 1728341909
transform -1 0 9310 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2398_
timestamp 1728341909
transform 1 0 8690 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2399_
timestamp 1728341909
transform -1 0 7570 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2400_
timestamp 1728341909
transform 1 0 7310 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2401_
timestamp 1728341909
transform 1 0 8430 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2402_
timestamp 1728341909
transform -1 0 6370 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2403_
timestamp 1728341909
transform -1 0 6570 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2404_
timestamp 1728341909
transform -1 0 7530 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2405_
timestamp 1728341909
transform -1 0 7310 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2406_
timestamp 1728341909
transform 1 0 7030 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2407_
timestamp 1728341909
transform -1 0 6570 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2408_
timestamp 1728341909
transform -1 0 5870 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2409_
timestamp 1728341909
transform 1 0 6950 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2410_
timestamp 1728341909
transform -1 0 7230 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2411_
timestamp 1728341909
transform -1 0 6790 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2412_
timestamp 1728341909
transform -1 0 7450 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2413_
timestamp 1728341909
transform 1 0 6970 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2414_
timestamp 1728341909
transform 1 0 6790 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2415_
timestamp 1728341909
transform -1 0 7990 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2416_
timestamp 1728341909
transform 1 0 7730 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2417_
timestamp 1728341909
transform -1 0 8970 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2418_
timestamp 1728341909
transform -1 0 8750 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2419_
timestamp 1728341909
transform 1 0 7010 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2420_
timestamp 1728341909
transform 1 0 2170 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2421_
timestamp 1728341909
transform -1 0 9630 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2422_
timestamp 1728341909
transform 1 0 8210 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2423_
timestamp 1728341909
transform 1 0 8930 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2424_
timestamp 1728341909
transform 1 0 8710 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2425_
timestamp 1728341909
transform 1 0 3110 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2426_
timestamp 1728341909
transform 1 0 8690 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2427_
timestamp 1728341909
transform 1 0 8770 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2428_
timestamp 1728341909
transform 1 0 9170 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2429_
timestamp 1728341909
transform 1 0 9390 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2430_
timestamp 1728341909
transform 1 0 8750 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2431_
timestamp 1728341909
transform -1 0 9210 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2432_
timestamp 1728341909
transform 1 0 9430 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2433_
timestamp 1728341909
transform -1 0 9850 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2434_
timestamp 1728341909
transform -1 0 9930 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2435_
timestamp 1728341909
transform 1 0 4390 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2436_
timestamp 1728341909
transform 1 0 9150 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2437_
timestamp 1728341909
transform 1 0 10830 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2438_
timestamp 1728341909
transform -1 0 10890 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2439_
timestamp 1728341909
transform -1 0 10870 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2440_
timestamp 1728341909
transform 1 0 8990 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2441_
timestamp 1728341909
transform -1 0 6130 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2442_
timestamp 1728341909
transform -1 0 8210 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2443_
timestamp 1728341909
transform 1 0 3770 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2444_
timestamp 1728341909
transform -1 0 4650 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2445_
timestamp 1728341909
transform -1 0 8550 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2446_
timestamp 1728341909
transform 1 0 8190 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2447_
timestamp 1728341909
transform 1 0 8030 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2448_
timestamp 1728341909
transform 1 0 8430 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2449_
timestamp 1728341909
transform -1 0 8710 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2450_
timestamp 1728341909
transform -1 0 8910 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2451_
timestamp 1728341909
transform 1 0 3770 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2452_
timestamp 1728341909
transform 1 0 7550 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2453_
timestamp 1728341909
transform -1 0 6570 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2454_
timestamp 1728341909
transform -1 0 6290 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2455_
timestamp 1728341909
transform -1 0 6570 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2456_
timestamp 1728341909
transform -1 0 8690 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2457_
timestamp 1728341909
transform -1 0 8910 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2458_
timestamp 1728341909
transform -1 0 6750 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2459_
timestamp 1728341909
transform -1 0 3530 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2460_
timestamp 1728341909
transform 1 0 7050 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2461_
timestamp 1728341909
transform 1 0 6970 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2462_
timestamp 1728341909
transform -1 0 7250 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2463_
timestamp 1728341909
transform -1 0 7270 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2464_
timestamp 1728341909
transform 1 0 4430 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2465_
timestamp 1728341909
transform -1 0 7330 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2466_
timestamp 1728341909
transform -1 0 3310 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2467_
timestamp 1728341909
transform 1 0 6130 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2468_
timestamp 1728341909
transform -1 0 6250 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2469_
timestamp 1728341909
transform -1 0 6090 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2470_
timestamp 1728341909
transform -1 0 6350 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2471_
timestamp 1728341909
transform -1 0 8010 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2472_
timestamp 1728341909
transform -1 0 6030 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2473_
timestamp 1728341909
transform -1 0 5370 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2474_
timestamp 1728341909
transform -1 0 5290 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2475_
timestamp 1728341909
transform -1 0 7750 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2476_
timestamp 1728341909
transform -1 0 2670 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2477_
timestamp 1728341909
transform -1 0 5150 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2478_
timestamp 1728341909
transform 1 0 5230 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2479_
timestamp 1728341909
transform -1 0 7970 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2480_
timestamp 1728341909
transform 1 0 5870 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2481_
timestamp 1728341909
transform 1 0 4130 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2482_
timestamp 1728341909
transform -1 0 2410 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2483_
timestamp 1728341909
transform -1 0 4650 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2484_
timestamp 1728341909
transform -1 0 5690 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2485_
timestamp 1728341909
transform -1 0 6930 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2486_
timestamp 1728341909
transform 1 0 3050 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2487_
timestamp 1728341909
transform -1 0 5630 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2488_
timestamp 1728341909
transform 1 0 6390 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2489_
timestamp 1728341909
transform -1 0 6670 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2490_
timestamp 1728341909
transform 1 0 7650 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2491_
timestamp 1728341909
transform -1 0 7890 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2492_
timestamp 1728341909
transform -1 0 2830 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2493_
timestamp 1728341909
transform -1 0 5470 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2494_
timestamp 1728341909
transform -1 0 6550 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2495_
timestamp 1728341909
transform 1 0 6790 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2496_
timestamp 1728341909
transform 1 0 7510 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2497_
timestamp 1728341909
transform -1 0 7750 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2498_
timestamp 1728341909
transform -1 0 8730 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2499_
timestamp 1728341909
transform 1 0 8970 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2500_
timestamp 1728341909
transform -1 0 7590 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2501_
timestamp 1728341909
transform -1 0 6710 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2502_
timestamp 1728341909
transform -1 0 7570 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2503_
timestamp 1728341909
transform 1 0 11070 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2504_
timestamp 1728341909
transform -1 0 4510 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2505_
timestamp 1728341909
transform -1 0 5650 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2506_
timestamp 1728341909
transform -1 0 6670 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2507_
timestamp 1728341909
transform 1 0 5810 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2508_
timestamp 1728341909
transform 1 0 5610 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2509_
timestamp 1728341909
transform -1 0 8770 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2510_
timestamp 1728341909
transform -1 0 8030 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2511_
timestamp 1728341909
transform -1 0 7350 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2512_
timestamp 1728341909
transform 1 0 7050 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2513_
timestamp 1728341909
transform 1 0 6830 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2514_
timestamp 1728341909
transform 1 0 6990 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2515_
timestamp 1728341909
transform 1 0 10330 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2516_
timestamp 1728341909
transform 1 0 8470 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2517_
timestamp 1728341909
transform 1 0 10570 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2518_
timestamp 1728341909
transform -1 0 9670 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2519_
timestamp 1728341909
transform 1 0 9910 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2520_
timestamp 1728341909
transform -1 0 10370 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2521_
timestamp 1728341909
transform -1 0 8470 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2522_
timestamp 1728341909
transform 1 0 6030 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2523_
timestamp 1728341909
transform 1 0 5850 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2524_
timestamp 1728341909
transform 1 0 8230 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2525_
timestamp 1728341909
transform 1 0 6730 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2526_
timestamp 1728341909
transform -1 0 7730 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2527_
timestamp 1728341909
transform 1 0 7950 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2528_
timestamp 1728341909
transform -1 0 8010 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2529_
timestamp 1728341909
transform 1 0 7790 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2530_
timestamp 1728341909
transform -1 0 7750 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2531_
timestamp 1728341909
transform -1 0 7770 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2532_
timestamp 1728341909
transform 1 0 7770 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2533_
timestamp 1728341909
transform -1 0 5430 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2534_
timestamp 1728341909
transform -1 0 5850 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2535_
timestamp 1728341909
transform -1 0 7530 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2536_
timestamp 1728341909
transform 1 0 7330 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2537_
timestamp 1728341909
transform 1 0 7250 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2538_
timestamp 1728341909
transform 1 0 7970 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2539_
timestamp 1728341909
transform 1 0 5830 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2540_
timestamp 1728341909
transform 1 0 5550 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2541_
timestamp 1728341909
transform 1 0 6070 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2542_
timestamp 1728341909
transform -1 0 6610 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2543_
timestamp 1728341909
transform -1 0 6570 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2544_
timestamp 1728341909
transform 1 0 6110 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2545_
timestamp 1728341909
transform 1 0 6810 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2546_
timestamp 1728341909
transform 1 0 6070 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2547_
timestamp 1728341909
transform 1 0 6290 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2548_
timestamp 1728341909
transform 1 0 7070 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2549_
timestamp 1728341909
transform 1 0 7330 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2550_
timestamp 1728341909
transform -1 0 7490 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2551_
timestamp 1728341909
transform -1 0 6210 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2552_
timestamp 1728341909
transform -1 0 4770 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2553_
timestamp 1728341909
transform -1 0 5810 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2554_
timestamp 1728341909
transform -1 0 5530 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2555_
timestamp 1728341909
transform 1 0 5590 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2556_
timestamp 1728341909
transform 1 0 4970 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2557_
timestamp 1728341909
transform 1 0 5710 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2558_
timestamp 1728341909
transform -1 0 6350 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2559_
timestamp 1728341909
transform 1 0 6030 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2560_
timestamp 1728341909
transform 1 0 4290 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2561_
timestamp 1728341909
transform -1 0 5350 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2562_
timestamp 1728341909
transform 1 0 4970 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2563_
timestamp 1728341909
transform -1 0 4870 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2564_
timestamp 1728341909
transform -1 0 4530 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2565_
timestamp 1728341909
transform 1 0 4670 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2566_
timestamp 1728341909
transform -1 0 4890 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2567_
timestamp 1728341909
transform 1 0 5090 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2568_
timestamp 1728341909
transform 1 0 5230 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2569_
timestamp 1728341909
transform -1 0 4110 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2570_
timestamp 1728341909
transform 1 0 5130 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2571_
timestamp 1728341909
transform 1 0 4250 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2572_
timestamp 1728341909
transform -1 0 4370 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2573_
timestamp 1728341909
transform 1 0 4610 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2574_
timestamp 1728341909
transform 1 0 5330 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2575_
timestamp 1728341909
transform -1 0 4890 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2576_
timestamp 1728341909
transform 1 0 5070 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2577_
timestamp 1728341909
transform 1 0 4810 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2578_
timestamp 1728341909
transform -1 0 4750 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2579_
timestamp 1728341909
transform 1 0 4610 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__2580_
timestamp 1728341909
transform 1 0 4650 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2581_
timestamp 1728341909
transform -1 0 4090 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2582_
timestamp 1728341909
transform -1 0 3230 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2583_
timestamp 1728341909
transform 1 0 2170 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2584_
timestamp 1728341909
transform 1 0 3130 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2585_
timestamp 1728341909
transform -1 0 6290 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2586_
timestamp 1728341909
transform -1 0 3650 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2587_
timestamp 1728341909
transform -1 0 3390 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2588_
timestamp 1728341909
transform -1 0 2910 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2589_
timestamp 1728341909
transform -1 0 2910 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2590_
timestamp 1728341909
transform 1 0 3530 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__2591_
timestamp 1728341909
transform -1 0 3010 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2592_
timestamp 1728341909
transform 1 0 2510 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2593_
timestamp 1728341909
transform -1 0 2610 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2594_
timestamp 1728341909
transform -1 0 2630 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2595_
timestamp 1728341909
transform -1 0 3710 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__2596_
timestamp 1728341909
transform 1 0 3310 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2597_
timestamp 1728341909
transform 1 0 3250 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2598_
timestamp 1728341909
transform -1 0 3130 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2599_
timestamp 1728341909
transform -1 0 3130 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2600_
timestamp 1728341909
transform 1 0 2850 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2601_
timestamp 1728341909
transform -1 0 2410 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2602_
timestamp 1728341909
transform -1 0 2670 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2603_
timestamp 1728341909
transform -1 0 2270 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2604_
timestamp 1728341909
transform 1 0 2410 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2605_
timestamp 1728341909
transform -1 0 2410 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2606_
timestamp 1728341909
transform 1 0 2130 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2607_
timestamp 1728341909
transform -1 0 1490 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2608_
timestamp 1728341909
transform -1 0 1010 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2609_
timestamp 1728341909
transform 1 0 1970 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2610_
timestamp 1728341909
transform 1 0 1210 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2611_
timestamp 1728341909
transform -1 0 1190 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2612_
timestamp 1728341909
transform -1 0 930 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2613_
timestamp 1728341909
transform -1 0 1910 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2614_
timestamp 1728341909
transform -1 0 530 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2615_
timestamp 1728341909
transform 1 0 1710 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2616_
timestamp 1728341909
transform 1 0 1450 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2617_
timestamp 1728341909
transform -1 0 1450 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2618_
timestamp 1728341909
transform -1 0 1690 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2619_
timestamp 1728341909
transform 1 0 730 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2620_
timestamp 1728341909
transform -1 0 1250 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2621_
timestamp 1728341909
transform 1 0 990 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2622_
timestamp 1728341909
transform -1 0 1210 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2623_
timestamp 1728341909
transform 1 0 950 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2624_
timestamp 1728341909
transform -1 0 490 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2625_
timestamp 1728341909
transform -1 0 2570 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2626_
timestamp 1728341909
transform 1 0 1590 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2627_
timestamp 1728341909
transform 1 0 1330 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2628_
timestamp 1728341909
transform 1 0 730 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2629_
timestamp 1728341909
transform -1 0 3330 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2630_
timestamp 1728341909
transform 1 0 4190 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2631_
timestamp 1728341909
transform -1 0 4850 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2632_
timestamp 1728341909
transform 1 0 10830 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2633_
timestamp 1728341909
transform 1 0 3830 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2634_
timestamp 1728341909
transform 1 0 8930 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2635_
timestamp 1728341909
transform -1 0 2210 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2636_
timestamp 1728341909
transform -1 0 9090 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2637_
timestamp 1728341909
transform 1 0 4290 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2638_
timestamp 1728341909
transform 1 0 4790 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2639_
timestamp 1728341909
transform -1 0 9870 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2640_
timestamp 1728341909
transform -1 0 9810 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2641_
timestamp 1728341909
transform 1 0 10110 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2642_
timestamp 1728341909
transform -1 0 9450 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2643_
timestamp 1728341909
transform 1 0 10850 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2644_
timestamp 1728341909
transform -1 0 9690 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2645_
timestamp 1728341909
transform -1 0 9650 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__2646_
timestamp 1728341909
transform 1 0 10050 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2647_
timestamp 1728341909
transform -1 0 8530 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2648_
timestamp 1728341909
transform -1 0 4110 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__2649_
timestamp 1728341909
transform -1 0 5750 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2650_
timestamp 1728341909
transform 1 0 9250 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2651_
timestamp 1728341909
transform -1 0 5630 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2652_
timestamp 1728341909
transform -1 0 7790 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2653_
timestamp 1728341909
transform -1 0 7690 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2654_
timestamp 1728341909
transform 1 0 4610 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2655_
timestamp 1728341909
transform -1 0 5390 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2656_
timestamp 1728341909
transform -1 0 5970 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2657_
timestamp 1728341909
transform -1 0 6710 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2658_
timestamp 1728341909
transform 1 0 6210 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2659_
timestamp 1728341909
transform 1 0 6910 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2660_
timestamp 1728341909
transform -1 0 7190 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2661_
timestamp 1728341909
transform -1 0 4410 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2662_
timestamp 1728341909
transform 1 0 4370 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2663_
timestamp 1728341909
transform 1 0 6290 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2664_
timestamp 1728341909
transform -1 0 6550 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2665_
timestamp 1728341909
transform 1 0 7050 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2666_
timestamp 1728341909
transform 1 0 6790 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2667_
timestamp 1728341909
transform 1 0 7530 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2668_
timestamp 1728341909
transform 1 0 7270 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2669_
timestamp 1728341909
transform 1 0 7930 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2670_
timestamp 1728341909
transform -1 0 4150 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2671_
timestamp 1728341909
transform -1 0 5270 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__2672_
timestamp 1728341909
transform 1 0 5170 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2673_
timestamp 1728341909
transform 1 0 7130 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2674_
timestamp 1728341909
transform -1 0 7350 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2675_
timestamp 1728341909
transform 1 0 7590 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2676_
timestamp 1728341909
transform -1 0 7530 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2677_
timestamp 1728341909
transform 1 0 7710 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2678_
timestamp 1728341909
transform 1 0 7670 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2679_
timestamp 1728341909
transform 1 0 4110 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2680_
timestamp 1728341909
transform -1 0 4370 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2681_
timestamp 1728341909
transform 1 0 6070 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2682_
timestamp 1728341909
transform 1 0 6690 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2683_
timestamp 1728341909
transform 1 0 4030 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2684_
timestamp 1728341909
transform -1 0 5690 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2685_
timestamp 1728341909
transform 1 0 5410 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2686_
timestamp 1728341909
transform -1 0 6830 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2687_
timestamp 1728341909
transform 1 0 7290 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2688_
timestamp 1728341909
transform -1 0 7430 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2689_
timestamp 1728341909
transform 1 0 6450 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2690_
timestamp 1728341909
transform 1 0 6530 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2691_
timestamp 1728341909
transform 1 0 7030 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2692_
timestamp 1728341909
transform -1 0 7170 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2693_
timestamp 1728341909
transform 1 0 5010 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2694_
timestamp 1728341909
transform -1 0 5150 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2695_
timestamp 1728341909
transform 1 0 6590 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2696_
timestamp 1728341909
transform 1 0 6530 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2697_
timestamp 1728341909
transform 1 0 6950 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2698_
timestamp 1728341909
transform 1 0 6850 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2699_
timestamp 1728341909
transform -1 0 6290 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2700_
timestamp 1728341909
transform 1 0 5350 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2701_
timestamp 1728341909
transform -1 0 5430 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2702_
timestamp 1728341909
transform -1 0 5510 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2703_
timestamp 1728341909
transform -1 0 5530 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2704_
timestamp 1728341909
transform 1 0 5590 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2705_
timestamp 1728341909
transform 1 0 5850 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2706_
timestamp 1728341909
transform -1 0 6110 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2707_
timestamp 1728341909
transform -1 0 5850 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2708_
timestamp 1728341909
transform -1 0 2250 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2709_
timestamp 1728341909
transform -1 0 4910 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2710_
timestamp 1728341909
transform -1 0 4830 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2711_
timestamp 1728341909
transform -1 0 5030 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2712_
timestamp 1728341909
transform -1 0 5610 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2713_
timestamp 1728341909
transform -1 0 5750 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2714_
timestamp 1728341909
transform -1 0 6050 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2715_
timestamp 1728341909
transform 1 0 5770 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2716_
timestamp 1728341909
transform -1 0 6610 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2717_
timestamp 1728341909
transform 1 0 6550 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2718_
timestamp 1728341909
transform 1 0 6130 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2719_
timestamp 1728341909
transform -1 0 6290 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2720_
timestamp 1728341909
transform 1 0 4590 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2721_
timestamp 1728341909
transform 1 0 4870 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2722_
timestamp 1728341909
transform 1 0 5110 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2723_
timestamp 1728341909
transform -1 0 5370 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2724_
timestamp 1728341909
transform 1 0 6090 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2725_
timestamp 1728341909
transform 1 0 6330 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2726_
timestamp 1728341909
transform -1 0 6090 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__2727_
timestamp 1728341909
transform 1 0 5790 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__2728_
timestamp 1728341909
transform -1 0 4270 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2729_
timestamp 1728341909
transform -1 0 4130 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2730_
timestamp 1728341909
transform -1 0 5170 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2731_
timestamp 1728341909
transform -1 0 5290 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2732_
timestamp 1728341909
transform -1 0 5590 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2733_
timestamp 1728341909
transform -1 0 5850 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2734_
timestamp 1728341909
transform -1 0 5170 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2735_
timestamp 1728341909
transform 1 0 5370 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2736_
timestamp 1728341909
transform -1 0 8290 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__2737_
timestamp 1728341909
transform 1 0 3690 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2738_
timestamp 1728341909
transform 1 0 3870 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2739_
timestamp 1728341909
transform -1 0 3690 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2740_
timestamp 1728341909
transform -1 0 3630 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2741_
timestamp 1728341909
transform -1 0 3970 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2742_
timestamp 1728341909
transform -1 0 4110 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2743_
timestamp 1728341909
transform 1 0 4850 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2744_
timestamp 1728341909
transform 1 0 4590 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__2745_
timestamp 1728341909
transform 1 0 5070 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2746_
timestamp 1728341909
transform 1 0 4570 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2747_
timestamp 1728341909
transform 1 0 5490 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2748_
timestamp 1728341909
transform -1 0 4890 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2749_
timestamp 1728341909
transform -1 0 5250 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2750_
timestamp 1728341909
transform -1 0 5350 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2751_
timestamp 1728341909
transform 1 0 4330 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2752_
timestamp 1728341909
transform 1 0 3830 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2753_
timestamp 1728341909
transform -1 0 3370 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2754_
timestamp 1728341909
transform -1 0 2950 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2755_
timestamp 1728341909
transform 1 0 3210 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2756_
timestamp 1728341909
transform -1 0 3590 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2757_
timestamp 1728341909
transform -1 0 3610 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2758_
timestamp 1728341909
transform -1 0 3590 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2759_
timestamp 1728341909
transform -1 0 3470 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2760_
timestamp 1728341909
transform -1 0 3510 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2761_
timestamp 1728341909
transform -1 0 3650 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2762_
timestamp 1728341909
transform -1 0 3410 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2763_
timestamp 1728341909
transform 1 0 2970 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__2764_
timestamp 1728341909
transform 1 0 3250 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__2765_
timestamp 1728341909
transform -1 0 2570 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2766_
timestamp 1728341909
transform 1 0 3650 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__2767_
timestamp 1728341909
transform -1 0 4350 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2768_
timestamp 1728341909
transform 1 0 4430 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2769_
timestamp 1728341909
transform 1 0 5090 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2770_
timestamp 1728341909
transform -1 0 4590 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2771_
timestamp 1728341909
transform -1 0 4870 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2772_
timestamp 1728341909
transform -1 0 4850 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2773_
timestamp 1728341909
transform 1 0 2610 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2774_
timestamp 1728341909
transform -1 0 2470 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__2775_
timestamp 1728341909
transform 1 0 3830 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2776_
timestamp 1728341909
transform 1 0 4350 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2777_
timestamp 1728341909
transform 1 0 5090 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2778_
timestamp 1728341909
transform -1 0 4590 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2779_
timestamp 1728341909
transform 1 0 3910 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__2780_
timestamp 1728341909
transform 1 0 2690 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__2781_
timestamp 1728341909
transform -1 0 3910 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2782_
timestamp 1728341909
transform -1 0 2710 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2783_
timestamp 1728341909
transform 1 0 2410 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2784_
timestamp 1728341909
transform 1 0 490 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2785_
timestamp 1728341909
transform -1 0 2190 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2786_
timestamp 1728341909
transform 1 0 2450 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2787_
timestamp 1728341909
transform -1 0 2870 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2788_
timestamp 1728341909
transform -1 0 2370 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2789_
timestamp 1728341909
transform -1 0 3670 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2790_
timestamp 1728341909
transform 1 0 3150 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2791_
timestamp 1728341909
transform -1 0 2890 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2792_
timestamp 1728341909
transform -1 0 2790 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2793_
timestamp 1728341909
transform -1 0 2210 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__2794_
timestamp 1728341909
transform 1 0 2090 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2795_
timestamp 1728341909
transform 1 0 730 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2796_
timestamp 1728341909
transform 1 0 1670 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2797_
timestamp 1728341909
transform -1 0 1950 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2798_
timestamp 1728341909
transform 1 0 1170 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2799_
timestamp 1728341909
transform -1 0 1450 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2800_
timestamp 1728341909
transform -1 0 1710 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2801_
timestamp 1728341909
transform 1 0 1670 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2802_
timestamp 1728341909
transform 1 0 1750 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2803_
timestamp 1728341909
transform 1 0 3230 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2804_
timestamp 1728341909
transform -1 0 390 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__2805_
timestamp 1728341909
transform 1 0 6930 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2806_
timestamp 1728341909
transform -1 0 5350 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2807_
timestamp 1728341909
transform -1 0 4950 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2808_
timestamp 1728341909
transform 1 0 3870 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2809_
timestamp 1728341909
transform -1 0 4330 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2810_
timestamp 1728341909
transform -1 0 4690 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2811_
timestamp 1728341909
transform -1 0 4550 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2812_
timestamp 1728341909
transform 1 0 4170 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2813_
timestamp 1728341909
transform 1 0 3930 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__2814_
timestamp 1728341909
transform 1 0 4050 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__2815_
timestamp 1728341909
transform -1 0 4130 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2816_
timestamp 1728341909
transform 1 0 2430 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2817_
timestamp 1728341909
transform -1 0 2710 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__2818_
timestamp 1728341909
transform 1 0 2670 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2819_
timestamp 1728341909
transform 1 0 3110 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2820_
timestamp 1728341909
transform 1 0 3350 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2821_
timestamp 1728341909
transform -1 0 3890 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2822_
timestamp 1728341909
transform -1 0 4690 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2823_
timestamp 1728341909
transform -1 0 1670 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2824_
timestamp 1728341909
transform 1 0 490 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__2825_
timestamp 1728341909
transform 1 0 470 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2826_
timestamp 1728341909
transform -1 0 630 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__2827_
timestamp 1728341909
transform 1 0 1670 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2828_
timestamp 1728341909
transform -1 0 1950 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2829_
timestamp 1728341909
transform 1 0 1190 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2830_
timestamp 1728341909
transform -1 0 1450 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2831_
timestamp 1728341909
transform -1 0 1470 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__2832_
timestamp 1728341909
transform 1 0 1970 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2833_
timestamp 1728341909
transform -1 0 990 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__2834_
timestamp 1728341909
transform 1 0 810 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__2835_
timestamp 1728341909
transform 1 0 1050 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__2836_
timestamp 1728341909
transform 1 0 1270 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__2837_
timestamp 1728341909
transform 1 0 1590 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__2838_
timestamp 1728341909
transform -1 0 1470 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__2839_
timestamp 1728341909
transform 1 0 750 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__2840_
timestamp 1728341909
transform 1 0 1190 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2841_
timestamp 1728341909
transform 1 0 1990 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2842_
timestamp 1728341909
transform -1 0 1650 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2843_
timestamp 1728341909
transform -1 0 1750 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2844_
timestamp 1728341909
transform -1 0 1510 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__2845_
timestamp 1728341909
transform -1 0 1450 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2846_
timestamp 1728341909
transform 1 0 1230 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2847_
timestamp 1728341909
transform -1 0 1230 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__2848_
timestamp 1728341909
transform -1 0 1210 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2849_
timestamp 1728341909
transform -1 0 1510 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2850_
timestamp 1728341909
transform -1 0 1430 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2851_
timestamp 1728341909
transform -1 0 970 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2852_
timestamp 1728341909
transform -1 0 1030 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2853_
timestamp 1728341909
transform -1 0 2230 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2854_
timestamp 1728341909
transform 1 0 710 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__2855_
timestamp 1728341909
transform 1 0 2390 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__2856_
timestamp 1728341909
transform -1 0 1910 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__2857_
timestamp 1728341909
transform -1 0 2310 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__2858_
timestamp 1728341909
transform -1 0 2210 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__2859_
timestamp 1728341909
transform -1 0 790 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2860_
timestamp 1728341909
transform 1 0 470 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2861_
timestamp 1728341909
transform -1 0 30 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2862_
timestamp 1728341909
transform -1 0 990 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__2863_
timestamp 1728341909
transform 1 0 230 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__2864_
timestamp 1728341909
transform -1 0 270 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__2865_
timestamp 1728341909
transform 1 0 4390 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2866_
timestamp 1728341909
transform 1 0 4410 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2867_
timestamp 1728341909
transform 1 0 5510 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2868_
timestamp 1728341909
transform -1 0 2890 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2869_
timestamp 1728341909
transform -1 0 3170 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2870_
timestamp 1728341909
transform -1 0 2230 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2871_
timestamp 1728341909
transform 1 0 2250 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2872_
timestamp 1728341909
transform -1 0 4530 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2873_
timestamp 1728341909
transform 1 0 4270 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2874_
timestamp 1728341909
transform -1 0 4070 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2875_
timestamp 1728341909
transform -1 0 1630 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2876_
timestamp 1728341909
transform -1 0 770 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2877_
timestamp 1728341909
transform -1 0 3430 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2878_
timestamp 1728341909
transform -1 0 3870 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2879_
timestamp 1728341909
transform -1 0 1210 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2880_
timestamp 1728341909
transform 1 0 1390 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2881_
timestamp 1728341909
transform -1 0 1710 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2882_
timestamp 1728341909
transform -1 0 2390 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2883_
timestamp 1728341909
transform 1 0 4390 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2884_
timestamp 1728341909
transform 1 0 4110 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2885_
timestamp 1728341909
transform 1 0 3050 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2886_
timestamp 1728341909
transform 1 0 4610 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2887_
timestamp 1728341909
transform 1 0 5070 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2888_
timestamp 1728341909
transform 1 0 3330 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2889_
timestamp 1728341909
transform 1 0 3550 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2890_
timestamp 1728341909
transform -1 0 4330 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2891_
timestamp 1728341909
transform -1 0 4070 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2892_
timestamp 1728341909
transform -1 0 1930 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2893_
timestamp 1728341909
transform 1 0 3610 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2894_
timestamp 1728341909
transform 1 0 3810 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2895_
timestamp 1728341909
transform 1 0 4390 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2896_
timestamp 1728341909
transform -1 0 3790 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2897_
timestamp 1728341909
transform -1 0 5790 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2898_
timestamp 1728341909
transform 1 0 5110 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2899_
timestamp 1728341909
transform 1 0 5070 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2900_
timestamp 1728341909
transform 1 0 5330 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2901_
timestamp 1728341909
transform -1 0 4810 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2902_
timestamp 1728341909
transform -1 0 1470 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2903_
timestamp 1728341909
transform 1 0 2130 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2904_
timestamp 1728341909
transform 1 0 2390 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2905_
timestamp 1728341909
transform 1 0 1190 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2906_
timestamp 1728341909
transform 1 0 970 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2907_
timestamp 1728341909
transform 1 0 1170 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2908_
timestamp 1728341909
transform -1 0 1490 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2909_
timestamp 1728341909
transform -1 0 1710 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2910_
timestamp 1728341909
transform -1 0 1490 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2911_
timestamp 1728341909
transform -1 0 1490 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2912_
timestamp 1728341909
transform -1 0 2410 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2913_
timestamp 1728341909
transform -1 0 1650 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2914_
timestamp 1728341909
transform 1 0 2170 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2915_
timestamp 1728341909
transform 1 0 1950 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2916_
timestamp 1728341909
transform 1 0 1630 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2917_
timestamp 1728341909
transform -1 0 1710 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2918_
timestamp 1728341909
transform 1 0 1650 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2919_
timestamp 1728341909
transform -1 0 2190 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2920_
timestamp 1728341909
transform -1 0 1910 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2921_
timestamp 1728341909
transform -1 0 1970 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2922_
timestamp 1728341909
transform -1 0 1890 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2923_
timestamp 1728341909
transform -1 0 1930 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2924_
timestamp 1728341909
transform -1 0 2890 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2925_
timestamp 1728341909
transform 1 0 3370 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2926_
timestamp 1728341909
transform -1 0 2350 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2927_
timestamp 1728341909
transform -1 0 2390 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2928_
timestamp 1728341909
transform 1 0 4530 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2929_
timestamp 1728341909
transform 1 0 3370 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2930_
timestamp 1728341909
transform -1 0 2650 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2931_
timestamp 1728341909
transform -1 0 2890 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2932_
timestamp 1728341909
transform 1 0 3090 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2933_
timestamp 1728341909
transform -1 0 2650 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2934_
timestamp 1728341909
transform 1 0 2870 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2935_
timestamp 1728341909
transform -1 0 1250 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2936_
timestamp 1728341909
transform -1 0 790 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2937_
timestamp 1728341909
transform 1 0 510 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2938_
timestamp 1728341909
transform 1 0 1670 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2939_
timestamp 1728341909
transform -1 0 1450 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2940_
timestamp 1728341909
transform 1 0 3110 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2941_
timestamp 1728341909
transform 1 0 3110 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2942_
timestamp 1728341909
transform -1 0 3330 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2943_
timestamp 1728341909
transform -1 0 3170 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2944_
timestamp 1728341909
transform -1 0 3670 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2945_
timestamp 1728341909
transform 1 0 3110 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2946_
timestamp 1728341909
transform 1 0 3550 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2947_
timestamp 1728341909
transform 1 0 3130 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2948_
timestamp 1728341909
transform -1 0 4130 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2949_
timestamp 1728341909
transform 1 0 3090 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2950_
timestamp 1728341909
transform 1 0 2410 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2951_
timestamp 1728341909
transform -1 0 2650 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2952_
timestamp 1728341909
transform -1 0 2930 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2953_
timestamp 1728341909
transform -1 0 2130 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2954_
timestamp 1728341909
transform -1 0 2370 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2955_
timestamp 1728341909
transform 1 0 2950 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2956_
timestamp 1728341909
transform 1 0 3190 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2957_
timestamp 1728341909
transform 1 0 3690 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2958_
timestamp 1728341909
transform 1 0 2130 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2959_
timestamp 1728341909
transform 1 0 3410 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2960_
timestamp 1728341909
transform 1 0 3530 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2961_
timestamp 1728341909
transform 1 0 2650 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2962_
timestamp 1728341909
transform 1 0 2390 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2963_
timestamp 1728341909
transform 1 0 2910 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2964_
timestamp 1728341909
transform 1 0 2650 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2965_
timestamp 1728341909
transform -1 0 5730 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2966_
timestamp 1728341909
transform 1 0 4050 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2967_
timestamp 1728341909
transform -1 0 4530 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2968_
timestamp 1728341909
transform -1 0 4770 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2969_
timestamp 1728341909
transform -1 0 1270 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2970_
timestamp 1728341909
transform -1 0 1450 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2971_
timestamp 1728341909
transform -1 0 1470 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2972_
timestamp 1728341909
transform -1 0 1210 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2973_
timestamp 1728341909
transform -1 0 970 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2974_
timestamp 1728341909
transform -1 0 1710 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2975_
timestamp 1728341909
transform -1 0 1930 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2976_
timestamp 1728341909
transform 1 0 3810 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2977_
timestamp 1728341909
transform -1 0 4370 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2978_
timestamp 1728341909
transform 1 0 4090 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2979_
timestamp 1728341909
transform 1 0 1470 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2980_
timestamp 1728341909
transform -1 0 950 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2981_
timestamp 1728341909
transform -1 0 710 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2982_
timestamp 1728341909
transform 1 0 2150 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2983_
timestamp 1728341909
transform -1 0 470 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2984_
timestamp 1728341909
transform -1 0 250 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2985_
timestamp 1728341909
transform -1 0 30 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2986_
timestamp 1728341909
transform -1 0 290 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2987_
timestamp 1728341909
transform -1 0 550 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2988_
timestamp 1728341909
transform -1 0 510 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2989_
timestamp 1728341909
transform 1 0 270 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2990_
timestamp 1728341909
transform 1 0 10 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2991_
timestamp 1728341909
transform -1 0 290 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2992_
timestamp 1728341909
transform -1 0 1950 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2993_
timestamp 1728341909
transform -1 0 990 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2994_
timestamp 1728341909
transform -1 0 750 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2995_
timestamp 1728341909
transform 1 0 530 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2996_
timestamp 1728341909
transform -1 0 470 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2997_
timestamp 1728341909
transform -1 0 790 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2998_
timestamp 1728341909
transform -1 0 30 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2999_
timestamp 1728341909
transform -1 0 270 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__3000_
timestamp 1728341909
transform -1 0 30 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__3001_
timestamp 1728341909
transform -1 0 30 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__3002_
timestamp 1728341909
transform -1 0 510 0 1 730
box -12 -8 32 252
use FILL  FILL_0__3003_
timestamp 1728341909
transform -1 0 30 0 1 730
box -12 -8 32 252
use FILL  FILL_0__3004_
timestamp 1728341909
transform -1 0 770 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__3005_
timestamp 1728341909
transform 1 0 730 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__3006_
timestamp 1728341909
transform -1 0 30 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__3007_
timestamp 1728341909
transform 1 0 1730 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3008_
timestamp 1728341909
transform -1 0 990 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__3009_
timestamp 1728341909
transform -1 0 1250 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__3010_
timestamp 1728341909
transform -1 0 1250 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__3011_
timestamp 1728341909
transform -1 0 1010 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__3012_
timestamp 1728341909
transform -1 0 1390 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__3013_
timestamp 1728341909
transform -1 0 1170 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__3014_
timestamp 1728341909
transform 1 0 970 0 1 250
box -12 -8 32 252
use FILL  FILL_0__3015_
timestamp 1728341909
transform -1 0 1470 0 1 250
box -12 -8 32 252
use FILL  FILL_0__3016_
timestamp 1728341909
transform -1 0 1230 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__3017_
timestamp 1728341909
transform -1 0 1210 0 1 250
box -12 -8 32 252
use FILL  FILL_0__3018_
timestamp 1728341909
transform 1 0 990 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__3019_
timestamp 1728341909
transform -1 0 990 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__3020_
timestamp 1728341909
transform -1 0 3630 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3021_
timestamp 1728341909
transform -1 0 5890 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__3022_
timestamp 1728341909
transform 1 0 2730 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3023_
timestamp 1728341909
transform 1 0 2750 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3024_
timestamp 1728341909
transform 1 0 3730 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3025_
timestamp 1728341909
transform -1 0 4150 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__3026_
timestamp 1728341909
transform -1 0 3010 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3027_
timestamp 1728341909
transform -1 0 3410 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__3028_
timestamp 1728341909
transform -1 0 3930 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3029_
timestamp 1728341909
transform -1 0 4430 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3030_
timestamp 1728341909
transform 1 0 3410 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__3031_
timestamp 1728341909
transform -1 0 3690 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__3032_
timestamp 1728341909
transform -1 0 2490 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3033_
timestamp 1728341909
transform -1 0 2510 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3034_
timestamp 1728341909
transform 1 0 2650 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__3035_
timestamp 1728341909
transform -1 0 2910 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__3036_
timestamp 1728341909
transform 1 0 3230 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3037_
timestamp 1728341909
transform -1 0 3670 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__3038_
timestamp 1728341909
transform -1 0 3230 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3039_
timestamp 1728341909
transform 1 0 2970 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3040_
timestamp 1728341909
transform 1 0 2110 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__3041_
timestamp 1728341909
transform 1 0 2650 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__3042_
timestamp 1728341909
transform 1 0 7410 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__3043_
timestamp 1728341909
transform 1 0 6250 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__3044_
timestamp 1728341909
transform 1 0 5270 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__3045_
timestamp 1728341909
transform 1 0 5690 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3046_
timestamp 1728341909
transform 1 0 5410 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__3047_
timestamp 1728341909
transform 1 0 4750 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__3048_
timestamp 1728341909
transform 1 0 5090 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__3049_
timestamp 1728341909
transform 1 0 5790 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3050_
timestamp 1728341909
transform -1 0 6810 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3051_
timestamp 1728341909
transform -1 0 6270 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__3052_
timestamp 1728341909
transform 1 0 6310 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3053_
timestamp 1728341909
transform 1 0 6050 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3054_
timestamp 1728341909
transform 1 0 5790 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3055_
timestamp 1728341909
transform -1 0 5890 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3056_
timestamp 1728341909
transform 1 0 4550 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__3057_
timestamp 1728341909
transform 1 0 4310 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__3058_
timestamp 1728341909
transform -1 0 4430 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3059_
timestamp 1728341909
transform 1 0 4250 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__3060_
timestamp 1728341909
transform -1 0 4230 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__3061_
timestamp 1728341909
transform 1 0 3930 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3062_
timestamp 1728341909
transform -1 0 4750 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__3063_
timestamp 1728341909
transform 1 0 4490 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__3064_
timestamp 1728341909
transform 1 0 5950 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__3065_
timestamp 1728341909
transform 1 0 5730 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__3066_
timestamp 1728341909
transform -1 0 5730 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3067_
timestamp 1728341909
transform -1 0 5870 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__3068_
timestamp 1728341909
transform -1 0 6910 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3069_
timestamp 1728341909
transform -1 0 6410 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3070_
timestamp 1728341909
transform 1 0 6050 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3071_
timestamp 1728341909
transform -1 0 6330 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3072_
timestamp 1728341909
transform 1 0 6530 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__3073_
timestamp 1728341909
transform 1 0 6290 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__3074_
timestamp 1728341909
transform 1 0 350 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__3075_
timestamp 1728341909
transform -1 0 510 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__3076_
timestamp 1728341909
transform -1 0 4210 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3077_
timestamp 1728341909
transform 1 0 1950 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3078_
timestamp 1728341909
transform -1 0 5450 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3079_
timestamp 1728341909
transform 1 0 4990 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3080_
timestamp 1728341909
transform 1 0 4190 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3081_
timestamp 1728341909
transform 1 0 5830 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__3082_
timestamp 1728341909
transform -1 0 6830 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__3083_
timestamp 1728341909
transform 1 0 5990 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__3084_
timestamp 1728341909
transform -1 0 5670 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3085_
timestamp 1728341909
transform -1 0 4950 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3086_
timestamp 1728341909
transform 1 0 5430 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3087_
timestamp 1728341909
transform -1 0 5030 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__3088_
timestamp 1728341909
transform -1 0 5570 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__3089_
timestamp 1728341909
transform -1 0 5530 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__3090_
timestamp 1728341909
transform 1 0 4710 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3091_
timestamp 1728341909
transform -1 0 4670 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3092_
timestamp 1728341909
transform 1 0 5530 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__3093_
timestamp 1728341909
transform -1 0 3930 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__3094_
timestamp 1728341909
transform 1 0 4370 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__3095_
timestamp 1728341909
transform 1 0 4670 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__3096_
timestamp 1728341909
transform 1 0 4650 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__3097_
timestamp 1728341909
transform 1 0 4890 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__3098_
timestamp 1728341909
transform -1 0 4990 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__3099_
timestamp 1728341909
transform 1 0 5130 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__3100_
timestamp 1728341909
transform -1 0 5530 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__3101_
timestamp 1728341909
transform 1 0 5070 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__3102_
timestamp 1728341909
transform 1 0 4590 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__3103_
timestamp 1728341909
transform 1 0 4810 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__3104_
timestamp 1728341909
transform -1 0 4950 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3105_
timestamp 1728341909
transform 1 0 5270 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__3106_
timestamp 1728341909
transform 1 0 8450 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__3107_
timestamp 1728341909
transform 1 0 8210 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__3108_
timestamp 1728341909
transform 1 0 7970 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__3109_
timestamp 1728341909
transform -1 0 8510 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3110_
timestamp 1728341909
transform -1 0 8270 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3111_
timestamp 1728341909
transform 1 0 4450 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3112_
timestamp 1728341909
transform 1 0 4690 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3113_
timestamp 1728341909
transform -1 0 1210 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3114_
timestamp 1728341909
transform 1 0 710 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3115_
timestamp 1728341909
transform 1 0 4390 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__3116_
timestamp 1728341909
transform -1 0 4010 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3117_
timestamp 1728341909
transform -1 0 270 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__3118_
timestamp 1728341909
transform -1 0 30 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__3119_
timestamp 1728341909
transform -1 0 4870 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__3120_
timestamp 1728341909
transform 1 0 4370 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3121_
timestamp 1728341909
transform 1 0 5110 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__3122_
timestamp 1728341909
transform -1 0 4410 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3123_
timestamp 1728341909
transform -1 0 3670 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3124_
timestamp 1728341909
transform -1 0 3890 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3125_
timestamp 1728341909
transform -1 0 3630 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3126_
timestamp 1728341909
transform 1 0 4650 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3127_
timestamp 1728341909
transform 1 0 4670 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3128_
timestamp 1728341909
transform 1 0 4590 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__3129_
timestamp 1728341909
transform 1 0 3670 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__3130_
timestamp 1728341909
transform -1 0 1770 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3131_
timestamp 1728341909
transform -1 0 1270 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3132_
timestamp 1728341909
transform 1 0 990 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3133_
timestamp 1728341909
transform 1 0 3850 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3134_
timestamp 1728341909
transform 1 0 3430 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3135_
timestamp 1728341909
transform 1 0 3170 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3136_
timestamp 1728341909
transform 1 0 3650 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3137_
timestamp 1728341909
transform 1 0 3910 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3138_
timestamp 1728341909
transform -1 0 3950 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3139_
timestamp 1728341909
transform 1 0 1010 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3140_
timestamp 1728341909
transform 1 0 750 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3141_
timestamp 1728341909
transform -1 0 3930 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3142_
timestamp 1728341909
transform 1 0 3690 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3143_
timestamp 1728341909
transform -1 0 4130 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3144_
timestamp 1728341909
transform -1 0 3410 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3145_
timestamp 1728341909
transform 1 0 3150 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3146_
timestamp 1728341909
transform -1 0 3230 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3147_
timestamp 1728341909
transform 1 0 3470 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3148_
timestamp 1728341909
transform -1 0 3430 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3149_
timestamp 1728341909
transform -1 0 3410 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__3150_
timestamp 1728341909
transform 1 0 1990 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3151_
timestamp 1728341909
transform -1 0 2230 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3152_
timestamp 1728341909
transform 1 0 7470 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3153_
timestamp 1728341909
transform 1 0 4390 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3154_
timestamp 1728341909
transform -1 0 730 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3155_
timestamp 1728341909
transform 1 0 950 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3156_
timestamp 1728341909
transform 1 0 2910 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3157_
timestamp 1728341909
transform -1 0 2690 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3158_
timestamp 1728341909
transform 1 0 1910 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3159_
timestamp 1728341909
transform 1 0 2450 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3160_
timestamp 1728341909
transform 1 0 3070 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3161_
timestamp 1728341909
transform -1 0 2610 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3162_
timestamp 1728341909
transform -1 0 2390 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3163_
timestamp 1728341909
transform -1 0 1490 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3164_
timestamp 1728341909
transform 1 0 1190 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3165_
timestamp 1728341909
transform -1 0 270 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3166_
timestamp 1728341909
transform -1 0 30 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3167_
timestamp 1728341909
transform 1 0 1990 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3168_
timestamp 1728341909
transform 1 0 1930 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3169_
timestamp 1728341909
transform -1 0 2230 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3170_
timestamp 1728341909
transform 1 0 1970 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3171_
timestamp 1728341909
transform -1 0 2170 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3172_
timestamp 1728341909
transform 1 0 1830 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__3173_
timestamp 1728341909
transform -1 0 1710 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3174_
timestamp 1728341909
transform -1 0 1730 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3175_
timestamp 1728341909
transform -1 0 2970 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3176_
timestamp 1728341909
transform -1 0 2770 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3177_
timestamp 1728341909
transform 1 0 2210 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3178_
timestamp 1728341909
transform 1 0 2550 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3179_
timestamp 1728341909
transform 1 0 2210 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3180_
timestamp 1728341909
transform 1 0 3150 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3181_
timestamp 1728341909
transform -1 0 2870 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3182_
timestamp 1728341909
transform -1 0 2950 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3183_
timestamp 1728341909
transform 1 0 2710 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3184_
timestamp 1728341909
transform -1 0 2470 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3185_
timestamp 1728341909
transform -1 0 2470 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3186_
timestamp 1728341909
transform 1 0 1950 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3187_
timestamp 1728341909
transform -1 0 290 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3188_
timestamp 1728341909
transform -1 0 30 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3189_
timestamp 1728341909
transform 1 0 970 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3190_
timestamp 1728341909
transform -1 0 770 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3191_
timestamp 1728341909
transform -1 0 1030 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3192_
timestamp 1728341909
transform 1 0 1650 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3193_
timestamp 1728341909
transform 1 0 1390 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3194_
timestamp 1728341909
transform 1 0 3190 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3195_
timestamp 1728341909
transform 1 0 3150 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__3196_
timestamp 1728341909
transform 1 0 1890 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3197_
timestamp 1728341909
transform -1 0 2470 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__3198_
timestamp 1728341909
transform -1 0 2050 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3199_
timestamp 1728341909
transform -1 0 2310 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3200_
timestamp 1728341909
transform 1 0 750 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3201_
timestamp 1728341909
transform -1 0 990 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3202_
timestamp 1728341909
transform 1 0 990 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3203_
timestamp 1728341909
transform -1 0 1250 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3204_
timestamp 1728341909
transform -1 0 510 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3205_
timestamp 1728341909
transform -1 0 510 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3206_
timestamp 1728341909
transform 1 0 1010 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__3207_
timestamp 1728341909
transform -1 0 270 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3208_
timestamp 1728341909
transform -1 0 30 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3209_
timestamp 1728341909
transform 1 0 250 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3210_
timestamp 1728341909
transform -1 0 30 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3211_
timestamp 1728341909
transform -1 0 1510 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3212_
timestamp 1728341909
transform -1 0 1250 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3213_
timestamp 1728341909
transform 1 0 1530 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3214_
timestamp 1728341909
transform 1 0 1270 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3215_
timestamp 1728341909
transform -1 0 1230 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3216_
timestamp 1728341909
transform 1 0 970 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3217_
timestamp 1728341909
transform -1 0 270 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3218_
timestamp 1728341909
transform -1 0 30 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3219_
timestamp 1728341909
transform -1 0 1550 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3220_
timestamp 1728341909
transform 1 0 1770 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3221_
timestamp 1728341909
transform -1 0 290 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3222_
timestamp 1728341909
transform -1 0 30 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3223_
timestamp 1728341909
transform -1 0 770 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__3224_
timestamp 1728341909
transform 1 0 490 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3225_
timestamp 1728341909
transform -1 0 270 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3226_
timestamp 1728341909
transform -1 0 30 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3227_
timestamp 1728341909
transform -1 0 290 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__3228_
timestamp 1728341909
transform -1 0 30 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__3229_
timestamp 1728341909
transform -1 0 1950 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__3230_
timestamp 1728341909
transform 1 0 1670 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__3231_
timestamp 1728341909
transform 1 0 1470 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__3232_
timestamp 1728341909
transform -1 0 1730 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__3233_
timestamp 1728341909
transform 1 0 1030 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3234_
timestamp 1728341909
transform -1 0 1310 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3235_
timestamp 1728341909
transform 1 0 990 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3236_
timestamp 1728341909
transform 1 0 1250 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3237_
timestamp 1728341909
transform 1 0 2170 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__3238_
timestamp 1728341909
transform 1 0 2410 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__3239_
timestamp 1728341909
transform -1 0 510 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3240_
timestamp 1728341909
transform -1 0 750 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3241_
timestamp 1728341909
transform 1 0 9650 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__3242_
timestamp 1728341909
transform -1 0 8990 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__3243_
timestamp 1728341909
transform 1 0 9410 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__3244_
timestamp 1728341909
transform 1 0 8710 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__3245_
timestamp 1728341909
transform 1 0 9010 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3246_
timestamp 1728341909
transform -1 0 9530 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3247_
timestamp 1728341909
transform 1 0 10430 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3248_
timestamp 1728341909
transform 1 0 10690 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3249_
timestamp 1728341909
transform -1 0 9430 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__3250_
timestamp 1728341909
transform 1 0 9350 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3251_
timestamp 1728341909
transform 1 0 9190 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__3252_
timestamp 1728341909
transform -1 0 9210 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__3253_
timestamp 1728341909
transform -1 0 7830 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3254_
timestamp 1728341909
transform -1 0 8090 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3255_
timestamp 1728341909
transform -1 0 9270 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3256_
timestamp 1728341909
transform 1 0 8210 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3257_
timestamp 1728341909
transform 1 0 7970 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3258_
timestamp 1728341909
transform 1 0 8510 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3259_
timestamp 1728341909
transform 1 0 9450 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3260_
timestamp 1728341909
transform -1 0 10810 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__3261_
timestamp 1728341909
transform -1 0 10350 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3262_
timestamp 1728341909
transform 1 0 9930 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3263_
timestamp 1728341909
transform 1 0 9610 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__3264_
timestamp 1728341909
transform 1 0 8950 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__3265_
timestamp 1728341909
transform -1 0 9690 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3266_
timestamp 1728341909
transform 1 0 9710 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3267_
timestamp 1728341909
transform -1 0 9610 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3268_
timestamp 1728341909
transform -1 0 9950 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3269_
timestamp 1728341909
transform -1 0 10450 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3270_
timestamp 1728341909
transform 1 0 10170 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3271_
timestamp 1728341909
transform -1 0 9990 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__3272_
timestamp 1728341909
transform 1 0 10210 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__3273_
timestamp 1728341909
transform -1 0 10110 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__3274_
timestamp 1728341909
transform -1 0 10210 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3275_
timestamp 1728341909
transform 1 0 9530 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__3276_
timestamp 1728341909
transform -1 0 9150 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3277_
timestamp 1728341909
transform -1 0 10610 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3278_
timestamp 1728341909
transform 1 0 10070 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3279_
timestamp 1728341909
transform -1 0 9850 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3280_
timestamp 1728341909
transform 1 0 9190 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__3281_
timestamp 1728341909
transform 1 0 8950 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__3282_
timestamp 1728341909
transform -1 0 6830 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__3283_
timestamp 1728341909
transform -1 0 6770 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3284_
timestamp 1728341909
transform 1 0 6530 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__3285_
timestamp 1728341909
transform 1 0 6970 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3286_
timestamp 1728341909
transform -1 0 7230 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3287_
timestamp 1728341909
transform -1 0 6590 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3288_
timestamp 1728341909
transform -1 0 6810 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3289_
timestamp 1728341909
transform -1 0 6770 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__3290_
timestamp 1728341909
transform 1 0 6490 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__3291_
timestamp 1728341909
transform 1 0 6990 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3292_
timestamp 1728341909
transform -1 0 7250 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3293_
timestamp 1728341909
transform 1 0 7090 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3294_
timestamp 1728341909
transform 1 0 6830 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3295_
timestamp 1728341909
transform 1 0 6030 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3296_
timestamp 1728341909
transform 1 0 5770 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3297_
timestamp 1728341909
transform 1 0 5390 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3298_
timestamp 1728341909
transform 1 0 5130 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3299_
timestamp 1728341909
transform 1 0 5570 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3300_
timestamp 1728341909
transform 1 0 5330 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3301_
timestamp 1728341909
transform 1 0 6830 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__3302_
timestamp 1728341909
transform 1 0 2910 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3303_
timestamp 1728341909
transform -1 0 2970 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3304_
timestamp 1728341909
transform 1 0 1910 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3305_
timestamp 1728341909
transform -1 0 2170 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3306_
timestamp 1728341909
transform 1 0 3830 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3307_
timestamp 1728341909
transform -1 0 4770 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3308_
timestamp 1728341909
transform -1 0 30 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__3309_
timestamp 1728341909
transform -1 0 30 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3310_
timestamp 1728341909
transform -1 0 710 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__3311_
timestamp 1728341909
transform -1 0 750 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3312_
timestamp 1728341909
transform -1 0 250 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__3313_
timestamp 1728341909
transform -1 0 290 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3314_
timestamp 1728341909
transform -1 0 30 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3315_
timestamp 1728341909
transform -1 0 30 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3316_
timestamp 1728341909
transform -1 0 530 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3317_
timestamp 1728341909
transform -1 0 750 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3449_
timestamp 1728341909
transform -1 0 3770 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3450_
timestamp 1728341909
transform 1 0 2930 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3451_
timestamp 1728341909
transform 1 0 3050 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3452_
timestamp 1728341909
transform -1 0 3310 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3453_
timestamp 1728341909
transform 1 0 3170 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3454_
timestamp 1728341909
transform -1 0 3530 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3455_
timestamp 1728341909
transform 1 0 9910 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3456_
timestamp 1728341909
transform 1 0 9470 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3457_
timestamp 1728341909
transform -1 0 9750 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3458_
timestamp 1728341909
transform -1 0 9910 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3459_
timestamp 1728341909
transform 1 0 10350 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3460_
timestamp 1728341909
transform -1 0 10650 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3461_
timestamp 1728341909
transform -1 0 10410 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3462_
timestamp 1728341909
transform -1 0 9970 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3463_
timestamp 1728341909
transform 1 0 10370 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3464_
timestamp 1728341909
transform -1 0 10170 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3465_
timestamp 1728341909
transform 1 0 10130 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0__3466_
timestamp 1728341909
transform -1 0 10150 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3467_
timestamp 1728341909
transform 1 0 8210 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3468_
timestamp 1728341909
transform 1 0 9050 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__3469_
timestamp 1728341909
transform 1 0 8510 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3470_
timestamp 1728341909
transform -1 0 8450 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3471_
timestamp 1728341909
transform 1 0 8590 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__3472_
timestamp 1728341909
transform 1 0 8830 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__3473_
timestamp 1728341909
transform -1 0 8650 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3474_
timestamp 1728341909
transform -1 0 8770 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3475_
timestamp 1728341909
transform -1 0 8890 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3476_
timestamp 1728341909
transform 1 0 9690 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3477_
timestamp 1728341909
transform 1 0 9130 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3478_
timestamp 1728341909
transform -1 0 9010 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3479_
timestamp 1728341909
transform 1 0 10490 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__3480_
timestamp 1728341909
transform -1 0 10050 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__3481_
timestamp 1728341909
transform -1 0 9910 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3482_
timestamp 1728341909
transform -1 0 9710 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__3483_
timestamp 1728341909
transform 1 0 10850 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3484_
timestamp 1728341909
transform 1 0 10830 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3485_
timestamp 1728341909
transform 1 0 11110 0 1 6490
box -12 -8 32 252
use FILL  FILL_0__3486_
timestamp 1728341909
transform 1 0 11070 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3487_
timestamp 1728341909
transform 1 0 10830 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3488_
timestamp 1728341909
transform 1 0 9470 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3489_
timestamp 1728341909
transform 1 0 9370 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3490_
timestamp 1728341909
transform -1 0 9630 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3491_
timestamp 1728341909
transform -1 0 9650 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3492_
timestamp 1728341909
transform 1 0 9850 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3493_
timestamp 1728341909
transform 1 0 10110 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3494_
timestamp 1728341909
transform 1 0 10250 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__3495_
timestamp 1728341909
transform -1 0 8750 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3496_
timestamp 1728341909
transform 1 0 9370 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3497_
timestamp 1728341909
transform 1 0 9890 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3498_
timestamp 1728341909
transform 1 0 9750 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__3499_
timestamp 1728341909
transform 1 0 9170 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3500_
timestamp 1728341909
transform -1 0 9430 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3501_
timestamp 1728341909
transform -1 0 9670 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3502_
timestamp 1728341909
transform 1 0 9510 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__3503_
timestamp 1728341909
transform 1 0 9990 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__3504_
timestamp 1728341909
transform -1 0 9950 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3505_
timestamp 1728341909
transform 1 0 10190 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3506_
timestamp 1728341909
transform 1 0 10710 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__3507_
timestamp 1728341909
transform -1 0 9330 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__3508_
timestamp 1728341909
transform -1 0 8450 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3509_
timestamp 1728341909
transform 1 0 8370 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__3510_
timestamp 1728341909
transform 1 0 9150 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3511_
timestamp 1728341909
transform -1 0 8910 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3512_
timestamp 1728341909
transform 1 0 8650 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3513_
timestamp 1728341909
transform -1 0 8930 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3514_
timestamp 1728341909
transform -1 0 8690 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3515_
timestamp 1728341909
transform -1 0 9090 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__3516_
timestamp 1728341909
transform 1 0 10930 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__3517_
timestamp 1728341909
transform -1 0 10250 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__3518_
timestamp 1728341909
transform 1 0 10330 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3519_
timestamp 1728341909
transform 1 0 10810 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3520_
timestamp 1728341909
transform -1 0 11110 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3521_
timestamp 1728341909
transform 1 0 7430 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3522_
timestamp 1728341909
transform -1 0 7950 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3523_
timestamp 1728341909
transform 1 0 8690 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3524_
timestamp 1728341909
transform 1 0 8470 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3525_
timestamp 1728341909
transform 1 0 8890 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3526_
timestamp 1728341909
transform -1 0 9170 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3527_
timestamp 1728341909
transform -1 0 8230 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3528_
timestamp 1728341909
transform -1 0 9870 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3529_
timestamp 1728341909
transform 1 0 9970 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__3530_
timestamp 1728341909
transform 1 0 10070 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3531_
timestamp 1728341909
transform -1 0 10110 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3532_
timestamp 1728341909
transform 1 0 10250 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__3533_
timestamp 1728341909
transform -1 0 8170 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3534_
timestamp 1728341909
transform -1 0 8430 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3535_
timestamp 1728341909
transform -1 0 7990 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3536_
timestamp 1728341909
transform -1 0 8210 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3537_
timestamp 1728341909
transform 1 0 8310 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__3538_
timestamp 1728341909
transform -1 0 8590 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__3539_
timestamp 1728341909
transform -1 0 9490 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__3540_
timestamp 1728341909
transform 1 0 9710 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__3541_
timestamp 1728341909
transform -1 0 9790 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__3542_
timestamp 1728341909
transform -1 0 7450 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3543_
timestamp 1728341909
transform -1 0 7710 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3544_
timestamp 1728341909
transform 1 0 7930 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3545_
timestamp 1728341909
transform 1 0 8790 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__3546_
timestamp 1728341909
transform -1 0 8230 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3547_
timestamp 1728341909
transform 1 0 8650 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3548_
timestamp 1728341909
transform -1 0 8910 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3549_
timestamp 1728341909
transform -1 0 8870 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__3550_
timestamp 1728341909
transform 1 0 8850 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3551_
timestamp 1728341909
transform 1 0 9130 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3552_
timestamp 1728341909
transform 1 0 9270 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__3553_
timestamp 1728341909
transform 1 0 9010 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__3554_
timestamp 1728341909
transform 1 0 8930 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__3555_
timestamp 1728341909
transform -1 0 8510 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3556_
timestamp 1728341909
transform 1 0 8410 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3557_
timestamp 1728341909
transform -1 0 8070 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__3558_
timestamp 1728341909
transform -1 0 7710 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3559_
timestamp 1728341909
transform 1 0 7670 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3560_
timestamp 1728341909
transform 1 0 8190 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3561_
timestamp 1728341909
transform -1 0 7930 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3562_
timestamp 1728341909
transform -1 0 8930 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3563_
timestamp 1728341909
transform -1 0 8910 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__3564_
timestamp 1728341909
transform 1 0 10010 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__3565_
timestamp 1728341909
transform -1 0 9930 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__3566_
timestamp 1728341909
transform 1 0 9850 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3567_
timestamp 1728341909
transform 1 0 9930 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__3568_
timestamp 1728341909
transform 1 0 10150 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__3569_
timestamp 1728341909
transform 1 0 10150 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__3570_
timestamp 1728341909
transform 1 0 10610 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__3571_
timestamp 1728341909
transform -1 0 10590 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3572_
timestamp 1728341909
transform -1 0 11090 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3573_
timestamp 1728341909
transform 1 0 10970 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__3574_
timestamp 1728341909
transform 1 0 10710 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__3575_
timestamp 1728341909
transform 1 0 11110 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__3576_
timestamp 1728341909
transform 1 0 9890 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__3577_
timestamp 1728341909
transform -1 0 11130 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__3578_
timestamp 1728341909
transform 1 0 10730 0 -1 9850
box -12 -8 32 252
use FILL  FILL_0__3579_
timestamp 1728341909
transform -1 0 10430 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__3580_
timestamp 1728341909
transform -1 0 9130 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3581_
timestamp 1728341909
transform -1 0 8830 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__3582_
timestamp 1728341909
transform 1 0 8670 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__3583_
timestamp 1728341909
transform -1 0 8990 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__3584_
timestamp 1728341909
transform 1 0 8730 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__3585_
timestamp 1728341909
transform -1 0 9470 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__3586_
timestamp 1728341909
transform 1 0 9050 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__3587_
timestamp 1728341909
transform -1 0 9190 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__3588_
timestamp 1728341909
transform 1 0 9210 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__3589_
timestamp 1728341909
transform 1 0 9930 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__3590_
timestamp 1728341909
transform -1 0 10190 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__3591_
timestamp 1728341909
transform 1 0 9670 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__3592_
timestamp 1728341909
transform 1 0 9690 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__3593_
timestamp 1728341909
transform -1 0 9470 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__3594_
timestamp 1728341909
transform 1 0 10310 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3595_
timestamp 1728341909
transform 1 0 10870 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__3596_
timestamp 1728341909
transform -1 0 10830 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3597_
timestamp 1728341909
transform 1 0 10470 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__3598_
timestamp 1728341909
transform 1 0 11110 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__3599_
timestamp 1728341909
transform 1 0 11070 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3600_
timestamp 1728341909
transform 1 0 10950 0 -1 9370
box -12 -8 32 252
use FILL  FILL_0__3601_
timestamp 1728341909
transform 1 0 10130 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3602_
timestamp 1728341909
transform 1 0 10370 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3603_
timestamp 1728341909
transform 1 0 10430 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3604_
timestamp 1728341909
transform 1 0 10650 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3605_
timestamp 1728341909
transform 1 0 11130 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3606_
timestamp 1728341909
transform 1 0 10610 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3607_
timestamp 1728341909
transform -1 0 9910 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3608_
timestamp 1728341909
transform -1 0 10150 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3609_
timestamp 1728341909
transform 1 0 10650 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3610_
timestamp 1728341909
transform 1 0 9470 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3611_
timestamp 1728341909
transform 1 0 9270 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__3612_
timestamp 1728341909
transform 1 0 9530 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__3613_
timestamp 1728341909
transform 1 0 9390 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3614_
timestamp 1728341909
transform -1 0 9790 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__3615_
timestamp 1728341909
transform -1 0 9670 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3616_
timestamp 1728341909
transform -1 0 8970 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3617_
timestamp 1728341909
transform -1 0 9230 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3618_
timestamp 1728341909
transform 1 0 9710 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3619_
timestamp 1728341909
transform 1 0 10870 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3620_
timestamp 1728341909
transform -1 0 10610 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3621_
timestamp 1728341909
transform -1 0 10390 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3622_
timestamp 1728341909
transform 1 0 10630 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3623_
timestamp 1728341909
transform 1 0 9930 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3624_
timestamp 1728341909
transform 1 0 10650 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3625_
timestamp 1728341909
transform 1 0 10750 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__3626_
timestamp 1728341909
transform -1 0 10650 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3627_
timestamp 1728341909
transform -1 0 9630 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3628_
timestamp 1728341909
transform -1 0 10370 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3629_
timestamp 1728341909
transform 1 0 10590 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3630_
timestamp 1728341909
transform 1 0 10390 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3631_
timestamp 1728341909
transform -1 0 10550 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__3632_
timestamp 1728341909
transform -1 0 10890 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__3633_
timestamp 1728341909
transform 1 0 10850 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__3634_
timestamp 1728341909
transform -1 0 10670 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__3635_
timestamp 1728341909
transform -1 0 10390 0 1 10810
box -12 -8 32 252
use FILL  FILL_0__3636_
timestamp 1728341909
transform -1 0 10490 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__3637_
timestamp 1728341909
transform -1 0 10650 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__3638_
timestamp 1728341909
transform -1 0 10570 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3639_
timestamp 1728341909
transform -1 0 10410 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__3640_
timestamp 1728341909
transform -1 0 10870 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3641_
timestamp 1728341909
transform -1 0 10610 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3642_
timestamp 1728341909
transform -1 0 10930 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3643_
timestamp 1728341909
transform 1 0 10850 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3644_
timestamp 1728341909
transform -1 0 10410 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3645_
timestamp 1728341909
transform -1 0 10150 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3646_
timestamp 1728341909
transform -1 0 10910 0 -1 8890
box -12 -8 32 252
use FILL  FILL_0__3647_
timestamp 1728341909
transform 1 0 11010 0 1 250
box -12 -8 32 252
use FILL  FILL_0__3648_
timestamp 1728341909
transform 1 0 11090 0 1 8410
box -12 -8 32 252
use FILL  FILL_0__3649_
timestamp 1728341909
transform 1 0 10170 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3650_
timestamp 1728341909
transform 1 0 10290 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__3651_
timestamp 1728341909
transform 1 0 10390 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3652_
timestamp 1728341909
transform -1 0 10350 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3653_
timestamp 1728341909
transform 1 0 10570 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3654_
timestamp 1728341909
transform 1 0 8370 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3655_
timestamp 1728341909
transform -1 0 8630 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3656_
timestamp 1728341909
transform 1 0 8210 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__3657_
timestamp 1728341909
transform -1 0 8590 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__3658_
timestamp 1728341909
transform -1 0 8490 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__3659_
timestamp 1728341909
transform -1 0 8230 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0__3660_
timestamp 1728341909
transform -1 0 8350 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__3661_
timestamp 1728341909
transform -1 0 9210 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__3662_
timestamp 1728341909
transform -1 0 9450 0 1 10330
box -12 -8 32 252
use FILL  FILL_0__3663_
timestamp 1728341909
transform 1 0 9370 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3664_
timestamp 1728341909
transform -1 0 9610 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3665_
timestamp 1728341909
transform 1 0 8210 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3666_
timestamp 1728341909
transform -1 0 8450 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3667_
timestamp 1728341909
transform -1 0 9170 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3668_
timestamp 1728341909
transform -1 0 10390 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3669_
timestamp 1728341909
transform -1 0 10130 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3670_
timestamp 1728341909
transform -1 0 9890 0 1 9370
box -12 -8 32 252
use FILL  FILL_0__3671_
timestamp 1728341909
transform 1 0 8250 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3672_
timestamp 1728341909
transform 1 0 8490 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3673_
timestamp 1728341909
transform -1 0 9410 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3674_
timestamp 1728341909
transform -1 0 9870 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3675_
timestamp 1728341909
transform 1 0 10090 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3676_
timestamp 1728341909
transform -1 0 10130 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3677_
timestamp 1728341909
transform 1 0 9370 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3678_
timestamp 1728341909
transform -1 0 9210 0 -1 6970
box -12 -8 32 252
use FILL  FILL_0__3691_
timestamp 1728341909
transform 1 0 7690 0 1 250
box -12 -8 32 252
use FILL  FILL_0__3692_
timestamp 1728341909
transform -1 0 7950 0 1 250
box -12 -8 32 252
use FILL  FILL_0__3693_
timestamp 1728341909
transform -1 0 1930 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3694_
timestamp 1728341909
transform -1 0 30 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3695_
timestamp 1728341909
transform 1 0 530 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3696_
timestamp 1728341909
transform -1 0 30 0 1 9850
box -12 -8 32 252
use FILL  FILL_0__3697_
timestamp 1728341909
transform -1 0 30 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__3698_
timestamp 1728341909
transform -1 0 270 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0__3699_
timestamp 1728341909
transform 1 0 6090 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__3700_
timestamp 1728341909
transform -1 0 6250 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__3701_
timestamp 1728341909
transform -1 0 6230 0 1 250
box -12 -8 32 252
use FILL  FILL_0__3702_
timestamp 1728341909
transform -1 0 5210 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__3703_
timestamp 1728341909
transform -1 0 3450 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__3704_
timestamp 1728341909
transform -1 0 3230 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__3705_
timestamp 1728341909
transform -1 0 30 0 1 8890
box -12 -8 32 252
use FILL  FILL_0__3706_
timestamp 1728341909
transform -1 0 1270 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0__3707_
timestamp 1728341909
transform 1 0 11090 0 1 6970
box -12 -8 32 252
use FILL  FILL_0__3708_
timestamp 1728341909
transform 1 0 11090 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0__3709_
timestamp 1728341909
transform 1 0 11110 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3710_
timestamp 1728341909
transform 1 0 10870 0 1 7450
box -12 -8 32 252
use FILL  FILL_0__3711_
timestamp 1728341909
transform 1 0 11090 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0__3712_
timestamp 1728341909
transform 1 0 10870 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3713_
timestamp 1728341909
transform 1 0 10990 0 1 7930
box -12 -8 32 252
use FILL  FILL_0__3714_
timestamp 1728341909
transform 1 0 11110 0 -1 8410
box -12 -8 32 252
use FILL  FILL_0__3715_
timestamp 1728341909
transform 1 0 11090 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert0
timestamp 1728341909
transform 1 0 7730 0 1 10810
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert1
timestamp 1728341909
transform 1 0 8950 0 1 1690
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert2
timestamp 1728341909
transform 1 0 9150 0 1 6970
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert3
timestamp 1728341909
transform 1 0 5630 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert4
timestamp 1728341909
transform 1 0 6730 0 1 1690
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert5
timestamp 1728341909
transform -1 0 3990 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert6
timestamp 1728341909
transform 1 0 7150 0 1 10330
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert7
timestamp 1728341909
transform -1 0 4070 0 1 4090
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert8
timestamp 1728341909
transform -1 0 7510 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert9
timestamp 1728341909
transform 1 0 4430 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert10
timestamp 1728341909
transform -1 0 550 0 1 4090
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert11
timestamp 1728341909
transform -1 0 4750 0 1 2650
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert12
timestamp 1728341909
transform 1 0 710 0 1 5530
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert13
timestamp 1728341909
transform -1 0 5850 0 1 7450
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert14
timestamp 1728341909
transform 1 0 4490 0 1 2650
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert15
timestamp 1728341909
transform 1 0 5570 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert16
timestamp 1728341909
transform 1 0 2650 0 1 8410
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert17
timestamp 1728341909
transform 1 0 4150 0 1 6490
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert18
timestamp 1728341909
transform -1 0 30 0 1 2650
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert19
timestamp 1728341909
transform -1 0 290 0 1 8410
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert20
timestamp 1728341909
transform 1 0 490 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert21
timestamp 1728341909
transform -1 0 7030 0 1 4570
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert22
timestamp 1728341909
transform -1 0 10410 0 1 4090
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert23
timestamp 1728341909
transform -1 0 8750 0 1 4090
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert24
timestamp 1728341909
transform 1 0 8470 0 1 3130
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert25
timestamp 1728341909
transform -1 0 7030 0 1 3130
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert37
timestamp 1728341909
transform -1 0 950 0 1 5530
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert38
timestamp 1728341909
transform 1 0 1230 0 1 4570
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert39
timestamp 1728341909
transform -1 0 990 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert40
timestamp 1728341909
transform -1 0 2690 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert41
timestamp 1728341909
transform 1 0 9490 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert42
timestamp 1728341909
transform 1 0 8810 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert43
timestamp 1728341909
transform -1 0 8730 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert44
timestamp 1728341909
transform -1 0 8950 0 1 4570
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert45
timestamp 1728341909
transform 1 0 3810 0 1 4090
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert46
timestamp 1728341909
transform 1 0 5170 0 1 4090
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert47
timestamp 1728341909
transform 1 0 4270 0 1 2650
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert48
timestamp 1728341909
transform 1 0 5390 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert49
timestamp 1728341909
transform -1 0 2190 0 1 2650
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert50
timestamp 1728341909
transform 1 0 8270 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert51
timestamp 1728341909
transform -1 0 10370 0 1 4570
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert52
timestamp 1728341909
transform -1 0 9410 0 1 4570
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert53
timestamp 1728341909
transform -1 0 9490 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert54
timestamp 1728341909
transform -1 0 8330 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert55
timestamp 1728341909
transform -1 0 290 0 1 730
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert56
timestamp 1728341909
transform 1 0 4970 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert57
timestamp 1728341909
transform 1 0 4570 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert58
timestamp 1728341909
transform 1 0 1890 0 1 1690
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert59
timestamp 1728341909
transform 1 0 4330 0 1 730
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert60
timestamp 1728341909
transform -1 0 8710 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert61
timestamp 1728341909
transform 1 0 10110 0 -1 7450
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert62
timestamp 1728341909
transform 1 0 9150 0 -1 10330
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert63
timestamp 1728341909
transform 1 0 9230 0 1 7450
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert64
timestamp 1728341909
transform 1 0 8570 0 1 1210
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert65
timestamp 1728341909
transform -1 0 4970 0 1 4090
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert66
timestamp 1728341909
transform 1 0 5710 0 1 2650
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert67
timestamp 1728341909
transform 1 0 6550 0 1 5050
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert68
timestamp 1728341909
transform 1 0 7550 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert69
timestamp 1728341909
transform -1 0 6030 0 1 1690
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert70
timestamp 1728341909
transform 1 0 8710 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert71
timestamp 1728341909
transform 1 0 2410 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert72
timestamp 1728341909
transform 1 0 3850 0 1 1210
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert73
timestamp 1728341909
transform 1 0 2650 0 1 2650
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert74
timestamp 1728341909
transform -1 0 3650 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert75
timestamp 1728341909
transform -1 0 730 0 1 2170
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert76
timestamp 1728341909
transform 1 0 8710 0 1 4570
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert77
timestamp 1728341909
transform -1 0 8450 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert78
timestamp 1728341909
transform 1 0 8910 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert79
timestamp 1728341909
transform -1 0 9170 0 1 4570
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert80
timestamp 1728341909
transform 1 0 4150 0 -1 6490
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert81
timestamp 1728341909
transform 1 0 3290 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert82
timestamp 1728341909
transform 1 0 2150 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert83
timestamp 1728341909
transform -1 0 2630 0 -1 7930
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert26
timestamp 1728341909
transform -1 0 1370 0 1 3130
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert27
timestamp 1728341909
transform 1 0 3610 0 1 3130
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert28
timestamp 1728341909
transform 1 0 10 0 1 3130
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert29
timestamp 1728341909
transform 1 0 490 0 1 7930
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert30
timestamp 1728341909
transform 1 0 8170 0 1 5530
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert31
timestamp 1728341909
transform -1 0 7530 0 -1 10810
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert32
timestamp 1728341909
transform -1 0 3150 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert33
timestamp 1728341909
transform -1 0 7890 0 1 10330
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert34
timestamp 1728341909
transform -1 0 30 0 -1 11290
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert35
timestamp 1728341909
transform -1 0 5450 0 1 5050
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert36
timestamp 1728341909
transform -1 0 2830 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__1744_
timestamp 1728341909
transform -1 0 4430 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__1745_
timestamp 1728341909
transform 1 0 4210 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__1746_
timestamp 1728341909
transform -1 0 4190 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__1747_
timestamp 1728341909
transform -1 0 5650 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__1748_
timestamp 1728341909
transform 1 0 6570 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__1749_
timestamp 1728341909
transform 1 0 6330 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__1750_
timestamp 1728341909
transform 1 0 5170 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__1751_
timestamp 1728341909
transform 1 0 6810 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__1752_
timestamp 1728341909
transform 1 0 5390 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__1753_
timestamp 1728341909
transform 1 0 7530 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__1754_
timestamp 1728341909
transform -1 0 7070 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__1755_
timestamp 1728341909
transform -1 0 7290 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__1756_
timestamp 1728341909
transform -1 0 6370 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1757_
timestamp 1728341909
transform 1 0 7030 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__1758_
timestamp 1728341909
transform 1 0 6790 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__1759_
timestamp 1728341909
transform -1 0 3050 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__1760_
timestamp 1728341909
transform 1 0 2350 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__1761_
timestamp 1728341909
transform 1 0 7270 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__1762_
timestamp 1728341909
transform 1 0 2550 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__1763_
timestamp 1728341909
transform -1 0 8190 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__1764_
timestamp 1728341909
transform -1 0 8010 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__1765_
timestamp 1728341909
transform -1 0 8010 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__1766_
timestamp 1728341909
transform -1 0 7810 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__1767_
timestamp 1728341909
transform -1 0 7810 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__1768_
timestamp 1728341909
transform -1 0 5690 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1769_
timestamp 1728341909
transform 1 0 3130 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1770_
timestamp 1728341909
transform 1 0 10790 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1771_
timestamp 1728341909
transform 1 0 11030 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1772_
timestamp 1728341909
transform 1 0 10770 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1773_
timestamp 1728341909
transform 1 0 10310 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1774_
timestamp 1728341909
transform 1 0 10670 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1775_
timestamp 1728341909
transform -1 0 9490 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1776_
timestamp 1728341909
transform 1 0 9530 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1777_
timestamp 1728341909
transform -1 0 8710 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__1778_
timestamp 1728341909
transform -1 0 10910 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1779_
timestamp 1728341909
transform 1 0 10130 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1780_
timestamp 1728341909
transform 1 0 10890 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__1781_
timestamp 1728341909
transform -1 0 10910 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1782_
timestamp 1728341909
transform -1 0 11150 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1783_
timestamp 1728341909
transform -1 0 9950 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1784_
timestamp 1728341909
transform 1 0 10530 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1785_
timestamp 1728341909
transform 1 0 10870 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1786_
timestamp 1728341909
transform -1 0 10210 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1787_
timestamp 1728341909
transform 1 0 9210 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1788_
timestamp 1728341909
transform 1 0 10490 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1789_
timestamp 1728341909
transform -1 0 9350 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1790_
timestamp 1728341909
transform -1 0 10710 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1791_
timestamp 1728341909
transform 1 0 10930 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1792_
timestamp 1728341909
transform 1 0 5630 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1793_
timestamp 1728341909
transform 1 0 5350 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1794_
timestamp 1728341909
transform -1 0 4930 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1795_
timestamp 1728341909
transform 1 0 3710 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1796_
timestamp 1728341909
transform 1 0 4170 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1797_
timestamp 1728341909
transform -1 0 4690 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1798_
timestamp 1728341909
transform -1 0 11010 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1799_
timestamp 1728341909
transform -1 0 10910 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1800_
timestamp 1728341909
transform -1 0 10430 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1801_
timestamp 1728341909
transform -1 0 10090 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1802_
timestamp 1728341909
transform 1 0 9970 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1803_
timestamp 1728341909
transform 1 0 10210 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1804_
timestamp 1728341909
transform 1 0 10210 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1805_
timestamp 1728341909
transform -1 0 10010 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1806_
timestamp 1728341909
transform 1 0 9950 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1807_
timestamp 1728341909
transform -1 0 10070 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1808_
timestamp 1728341909
transform -1 0 10370 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1809_
timestamp 1728341909
transform -1 0 11030 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1810_
timestamp 1728341909
transform -1 0 6210 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1811_
timestamp 1728341909
transform -1 0 11110 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__1812_
timestamp 1728341909
transform -1 0 10190 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1813_
timestamp 1728341909
transform -1 0 7670 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1814_
timestamp 1728341909
transform -1 0 7510 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1815_
timestamp 1728341909
transform -1 0 10930 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1816_
timestamp 1728341909
transform -1 0 7570 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1817_
timestamp 1728341909
transform 1 0 6690 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1818_
timestamp 1728341909
transform 1 0 6630 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1819_
timestamp 1728341909
transform 1 0 6130 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1820_
timestamp 1728341909
transform 1 0 10330 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1821_
timestamp 1728341909
transform -1 0 6690 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1822_
timestamp 1728341909
transform 1 0 11110 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1823_
timestamp 1728341909
transform -1 0 9970 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1824_
timestamp 1728341909
transform 1 0 7270 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1825_
timestamp 1728341909
transform 1 0 6490 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1826_
timestamp 1728341909
transform 1 0 10910 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1827_
timestamp 1728341909
transform -1 0 7350 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1828_
timestamp 1728341909
transform 1 0 11110 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__1829_
timestamp 1728341909
transform -1 0 7370 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__1830_
timestamp 1728341909
transform 1 0 7510 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1831_
timestamp 1728341909
transform 1 0 10650 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__1832_
timestamp 1728341909
transform 1 0 10630 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1833_
timestamp 1728341909
transform 1 0 7190 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1834_
timestamp 1728341909
transform -1 0 6990 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1835_
timestamp 1728341909
transform -1 0 6430 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1836_
timestamp 1728341909
transform -1 0 5990 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1837_
timestamp 1728341909
transform -1 0 5510 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1838_
timestamp 1728341909
transform 1 0 5230 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1839_
timestamp 1728341909
transform 1 0 5810 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1840_
timestamp 1728341909
transform -1 0 8010 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__1841_
timestamp 1728341909
transform -1 0 4950 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__1842_
timestamp 1728341909
transform -1 0 6810 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1843_
timestamp 1728341909
transform 1 0 7130 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1844_
timestamp 1728341909
transform -1 0 10210 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1845_
timestamp 1728341909
transform 1 0 11110 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1846_
timestamp 1728341909
transform 1 0 11130 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1847_
timestamp 1728341909
transform -1 0 8050 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1848_
timestamp 1728341909
transform 1 0 10650 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1849_
timestamp 1728341909
transform -1 0 10570 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1850_
timestamp 1728341909
transform -1 0 8510 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1851_
timestamp 1728341909
transform -1 0 11130 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1852_
timestamp 1728341909
transform 1 0 9690 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1853_
timestamp 1728341909
transform 1 0 9210 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1854_
timestamp 1728341909
transform 1 0 9010 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1855_
timestamp 1728341909
transform 1 0 8770 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1856_
timestamp 1728341909
transform 1 0 9290 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1857_
timestamp 1728341909
transform 1 0 9070 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1858_
timestamp 1728341909
transform 1 0 7250 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1859_
timestamp 1728341909
transform -1 0 10670 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__1860_
timestamp 1728341909
transform 1 0 7050 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1861_
timestamp 1728341909
transform 1 0 7290 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1862_
timestamp 1728341909
transform -1 0 9790 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1863_
timestamp 1728341909
transform 1 0 8530 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1864_
timestamp 1728341909
transform 1 0 9830 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1865_
timestamp 1728341909
transform 1 0 7690 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1866_
timestamp 1728341909
transform -1 0 8870 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1867_
timestamp 1728341909
transform 1 0 9250 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1868_
timestamp 1728341909
transform 1 0 10810 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1869_
timestamp 1728341909
transform 1 0 9270 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1870_
timestamp 1728341909
transform -1 0 9050 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1871_
timestamp 1728341909
transform 1 0 8490 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1872_
timestamp 1728341909
transform 1 0 7770 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1873_
timestamp 1728341909
transform 1 0 6330 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1874_
timestamp 1728341909
transform -1 0 6790 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1875_
timestamp 1728341909
transform -1 0 6550 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1876_
timestamp 1728341909
transform 1 0 6610 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1877_
timestamp 1728341909
transform -1 0 8030 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1878_
timestamp 1728341909
transform -1 0 8290 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1879_
timestamp 1728341909
transform -1 0 8030 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1880_
timestamp 1728341909
transform -1 0 6970 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__1881_
timestamp 1728341909
transform -1 0 6290 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__1882_
timestamp 1728341909
transform 1 0 3450 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__1883_
timestamp 1728341909
transform -1 0 6990 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__1884_
timestamp 1728341909
transform -1 0 6510 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__1885_
timestamp 1728341909
transform 1 0 5790 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__1886_
timestamp 1728341909
transform -1 0 6190 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__1887_
timestamp 1728341909
transform 1 0 6810 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__1888_
timestamp 1728341909
transform 1 0 3570 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__1889_
timestamp 1728341909
transform -1 0 5930 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__1890_
timestamp 1728341909
transform 1 0 6390 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__1891_
timestamp 1728341909
transform -1 0 6030 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__1892_
timestamp 1728341909
transform 1 0 5590 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__1893_
timestamp 1728341909
transform 1 0 990 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__1894_
timestamp 1728341909
transform 1 0 5930 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__1895_
timestamp 1728341909
transform 1 0 6810 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__1896_
timestamp 1728341909
transform 1 0 5130 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__1897_
timestamp 1728341909
transform 1 0 5970 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__1898_
timestamp 1728341909
transform 1 0 6390 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__1899_
timestamp 1728341909
transform 1 0 6490 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__1900_
timestamp 1728341909
transform 1 0 510 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1901_
timestamp 1728341909
transform 1 0 7950 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__1902_
timestamp 1728341909
transform 1 0 8490 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1903_
timestamp 1728341909
transform 1 0 7850 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1904_
timestamp 1728341909
transform -1 0 10010 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1905_
timestamp 1728341909
transform 1 0 7510 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1906_
timestamp 1728341909
transform 1 0 7490 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1907_
timestamp 1728341909
transform 1 0 8630 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1908_
timestamp 1728341909
transform -1 0 7690 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1909_
timestamp 1728341909
transform 1 0 1790 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1910_
timestamp 1728341909
transform -1 0 9750 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1911_
timestamp 1728341909
transform 1 0 9470 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1912_
timestamp 1728341909
transform 1 0 6090 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1913_
timestamp 1728341909
transform 1 0 10610 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1914_
timestamp 1728341909
transform 1 0 10670 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1915_
timestamp 1728341909
transform -1 0 10230 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1916_
timestamp 1728341909
transform -1 0 5850 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1917_
timestamp 1728341909
transform 1 0 3990 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1918_
timestamp 1728341909
transform -1 0 770 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1919_
timestamp 1728341909
transform -1 0 50 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1920_
timestamp 1728341909
transform 1 0 990 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1921_
timestamp 1728341909
transform -1 0 1170 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1922_
timestamp 1728341909
transform -1 0 910 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1923_
timestamp 1728341909
transform 1 0 510 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1924_
timestamp 1728341909
transform -1 0 4450 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1925_
timestamp 1728341909
transform -1 0 290 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__1926_
timestamp 1728341909
transform 1 0 750 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1927_
timestamp 1728341909
transform -1 0 2050 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1928_
timestamp 1728341909
transform -1 0 1570 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1929_
timestamp 1728341909
transform 1 0 250 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1930_
timestamp 1728341909
transform 1 0 630 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1931_
timestamp 1728341909
transform 1 0 510 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1932_
timestamp 1728341909
transform -1 0 530 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1933_
timestamp 1728341909
transform 1 0 510 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1934_
timestamp 1728341909
transform -1 0 530 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1935_
timestamp 1728341909
transform -1 0 1510 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1936_
timestamp 1728341909
transform 1 0 770 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1937_
timestamp 1728341909
transform -1 0 530 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1938_
timestamp 1728341909
transform -1 0 50 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1939_
timestamp 1728341909
transform 1 0 270 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1940_
timestamp 1728341909
transform 1 0 790 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1941_
timestamp 1728341909
transform 1 0 510 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__1942_
timestamp 1728341909
transform 1 0 510 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__1943_
timestamp 1728341909
transform 1 0 8070 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__1944_
timestamp 1728341909
transform -1 0 7610 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1945_
timestamp 1728341909
transform -1 0 7390 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1946_
timestamp 1728341909
transform 1 0 8410 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1947_
timestamp 1728341909
transform -1 0 7590 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1948_
timestamp 1728341909
transform -1 0 6930 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1949_
timestamp 1728341909
transform -1 0 7170 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1950_
timestamp 1728341909
transform 1 0 8270 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1951_
timestamp 1728341909
transform 1 0 8270 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1952_
timestamp 1728341909
transform 1 0 9790 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1953_
timestamp 1728341909
transform -1 0 8350 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1954_
timestamp 1728341909
transform 1 0 8190 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1955_
timestamp 1728341909
transform 1 0 6390 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1956_
timestamp 1728341909
transform -1 0 7950 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1957_
timestamp 1728341909
transform 1 0 8030 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__1958_
timestamp 1728341909
transform 1 0 10390 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1959_
timestamp 1728341909
transform 1 0 7750 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1960_
timestamp 1728341909
transform 1 0 7830 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1961_
timestamp 1728341909
transform 1 0 10650 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1962_
timestamp 1728341909
transform 1 0 10450 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1963_
timestamp 1728341909
transform 1 0 9790 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1964_
timestamp 1728341909
transform -1 0 7330 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1965_
timestamp 1728341909
transform -1 0 7610 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1966_
timestamp 1728341909
transform -1 0 3470 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__1967_
timestamp 1728341909
transform -1 0 6930 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__1968_
timestamp 1728341909
transform 1 0 7470 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__1969_
timestamp 1728341909
transform -1 0 7730 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__1970_
timestamp 1728341909
transform 1 0 1470 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1971_
timestamp 1728341909
transform -1 0 770 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1972_
timestamp 1728341909
transform 1 0 1290 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1973_
timestamp 1728341909
transform 1 0 1550 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1974_
timestamp 1728341909
transform 1 0 8310 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__1975_
timestamp 1728341909
transform 1 0 2930 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__1976_
timestamp 1728341909
transform -1 0 7090 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1977_
timestamp 1728341909
transform -1 0 2790 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__1978_
timestamp 1728341909
transform -1 0 3770 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__1979_
timestamp 1728341909
transform -1 0 6470 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__1980_
timestamp 1728341909
transform 1 0 7730 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__1981_
timestamp 1728341909
transform 1 0 8250 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__1982_
timestamp 1728341909
transform -1 0 2990 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__1983_
timestamp 1728341909
transform 1 0 1670 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__1984_
timestamp 1728341909
transform 1 0 1750 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__1985_
timestamp 1728341909
transform 1 0 2410 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__1986_
timestamp 1728341909
transform -1 0 7090 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__1987_
timestamp 1728341909
transform 1 0 5030 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__1988_
timestamp 1728341909
transform -1 0 4930 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__1989_
timestamp 1728341909
transform 1 0 6690 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__1990_
timestamp 1728341909
transform -1 0 7210 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__1991_
timestamp 1728341909
transform -1 0 2010 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1992_
timestamp 1728341909
transform -1 0 1510 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1993_
timestamp 1728341909
transform -1 0 1790 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1994_
timestamp 1728341909
transform 1 0 2030 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1995_
timestamp 1728341909
transform 1 0 7990 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__1996_
timestamp 1728341909
transform -1 0 2210 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__1997_
timestamp 1728341909
transform -1 0 3930 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__1998_
timestamp 1728341909
transform -1 0 6450 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__1999_
timestamp 1728341909
transform -1 0 8170 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2000_
timestamp 1728341909
transform 1 0 1770 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2001_
timestamp 1728341909
transform 1 0 1250 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2002_
timestamp 1728341909
transform 1 0 1490 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2003_
timestamp 1728341909
transform 1 0 1510 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2004_
timestamp 1728341909
transform 1 0 7790 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2005_
timestamp 1728341909
transform 1 0 1950 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2006_
timestamp 1728341909
transform -1 0 6210 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2007_
timestamp 1728341909
transform 1 0 7490 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2008_
timestamp 1728341909
transform -1 0 8010 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2009_
timestamp 1728341909
transform 1 0 750 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2010_
timestamp 1728341909
transform -1 0 810 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2011_
timestamp 1728341909
transform 1 0 510 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2012_
timestamp 1728341909
transform 1 0 770 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2013_
timestamp 1728341909
transform 1 0 5410 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2014_
timestamp 1728341909
transform 1 0 1710 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2015_
timestamp 1728341909
transform -1 0 3910 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2016_
timestamp 1728341909
transform 1 0 6710 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2017_
timestamp 1728341909
transform -1 0 7250 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2018_
timestamp 1728341909
transform -1 0 1490 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2019_
timestamp 1728341909
transform -1 0 1550 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2020_
timestamp 1728341909
transform 1 0 1730 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2021_
timestamp 1728341909
transform 1 0 1690 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2022_
timestamp 1728341909
transform 1 0 4470 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2023_
timestamp 1728341909
transform 1 0 510 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2024_
timestamp 1728341909
transform 1 0 1410 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2025_
timestamp 1728341909
transform 1 0 2470 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2026_
timestamp 1728341909
transform -1 0 4670 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2027_
timestamp 1728341909
transform 1 0 7170 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2028_
timestamp 1728341909
transform -1 0 7450 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2029_
timestamp 1728341909
transform -1 0 50 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2030_
timestamp 1728341909
transform -1 0 530 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2031_
timestamp 1728341909
transform -1 0 290 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2032_
timestamp 1728341909
transform 1 0 510 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2033_
timestamp 1728341909
transform 1 0 7590 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2034_
timestamp 1728341909
transform 1 0 1190 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2035_
timestamp 1728341909
transform 1 0 2070 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2036_
timestamp 1728341909
transform 1 0 2870 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2037_
timestamp 1728341909
transform -1 0 4070 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2038_
timestamp 1728341909
transform 1 0 7510 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2039_
timestamp 1728341909
transform -1 0 7790 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2040_
timestamp 1728341909
transform -1 0 2910 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2041_
timestamp 1728341909
transform -1 0 530 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2042_
timestamp 1728341909
transform 1 0 1690 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2043_
timestamp 1728341909
transform -1 0 3790 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__2044_
timestamp 1728341909
transform 1 0 5330 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2045_
timestamp 1728341909
transform -1 0 4030 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2046_
timestamp 1728341909
transform 1 0 2830 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2047_
timestamp 1728341909
transform 1 0 2590 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2048_
timestamp 1728341909
transform -1 0 3530 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2049_
timestamp 1728341909
transform -1 0 2930 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2050_
timestamp 1728341909
transform -1 0 2410 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2051_
timestamp 1728341909
transform -1 0 2390 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2052_
timestamp 1728341909
transform -1 0 810 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2053_
timestamp 1728341909
transform -1 0 3370 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2054_
timestamp 1728341909
transform 1 0 3090 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2055_
timestamp 1728341909
transform -1 0 2730 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2056_
timestamp 1728341909
transform 1 0 4350 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2057_
timestamp 1728341909
transform -1 0 3910 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2058_
timestamp 1728341909
transform 1 0 4570 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2059_
timestamp 1728341909
transform -1 0 1930 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2060_
timestamp 1728341909
transform -1 0 3750 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2061_
timestamp 1728341909
transform 1 0 3490 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2062_
timestamp 1728341909
transform -1 0 3510 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2063_
timestamp 1728341909
transform 1 0 2450 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2064_
timestamp 1728341909
transform -1 0 2550 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2065_
timestamp 1728341909
transform -1 0 2350 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2066_
timestamp 1728341909
transform 1 0 2410 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2067_
timestamp 1728341909
transform -1 0 2730 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2068_
timestamp 1728341909
transform -1 0 2970 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2069_
timestamp 1728341909
transform 1 0 2510 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2070_
timestamp 1728341909
transform -1 0 1050 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2071_
timestamp 1728341909
transform -1 0 2770 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2072_
timestamp 1728341909
transform -1 0 2510 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2073_
timestamp 1728341909
transform -1 0 1250 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2074_
timestamp 1728341909
transform 1 0 3190 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2075_
timestamp 1728341909
transform -1 0 2670 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2076_
timestamp 1728341909
transform 1 0 2370 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2077_
timestamp 1728341909
transform -1 0 3230 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2078_
timestamp 1728341909
transform 1 0 2750 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2079_
timestamp 1728341909
transform -1 0 3870 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2080_
timestamp 1728341909
transform 1 0 4090 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2081_
timestamp 1728341909
transform -1 0 3650 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2082_
timestamp 1728341909
transform 1 0 5730 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2083_
timestamp 1728341909
transform -1 0 6470 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2084_
timestamp 1728341909
transform 1 0 9890 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2085_
timestamp 1728341909
transform -1 0 10410 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2086_
timestamp 1728341909
transform 1 0 10430 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2087_
timestamp 1728341909
transform 1 0 10970 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2088_
timestamp 1728341909
transform 1 0 10170 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2089_
timestamp 1728341909
transform -1 0 9470 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2090_
timestamp 1728341909
transform 1 0 10650 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2091_
timestamp 1728341909
transform 1 0 11150 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2092_
timestamp 1728341909
transform -1 0 10110 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2093_
timestamp 1728341909
transform 1 0 10170 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2094_
timestamp 1728341909
transform -1 0 10670 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2095_
timestamp 1728341909
transform 1 0 10730 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2096_
timestamp 1728341909
transform -1 0 11130 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2097_
timestamp 1728341909
transform -1 0 11070 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2098_
timestamp 1728341909
transform 1 0 10150 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2099_
timestamp 1728341909
transform 1 0 10630 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2100_
timestamp 1728341909
transform 1 0 10850 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2101_
timestamp 1728341909
transform 1 0 11090 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2102_
timestamp 1728341909
transform 1 0 3970 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2103_
timestamp 1728341909
transform 1 0 4210 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2104_
timestamp 1728341909
transform 1 0 3830 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2105_
timestamp 1728341909
transform -1 0 1730 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2106_
timestamp 1728341909
transform -1 0 2110 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2107_
timestamp 1728341909
transform -1 0 2630 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2108_
timestamp 1728341909
transform 1 0 1430 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2109_
timestamp 1728341909
transform -1 0 2850 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2110_
timestamp 1728341909
transform 1 0 3070 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2111_
timestamp 1728341909
transform 1 0 5270 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2112_
timestamp 1728341909
transform 1 0 11150 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2113_
timestamp 1728341909
transform -1 0 9730 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2114_
timestamp 1728341909
transform 1 0 9730 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2115_
timestamp 1728341909
transform -1 0 11050 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2116_
timestamp 1728341909
transform -1 0 10990 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2117_
timestamp 1728341909
transform -1 0 10590 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2118_
timestamp 1728341909
transform 1 0 8990 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2119_
timestamp 1728341909
transform -1 0 11070 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2120_
timestamp 1728341909
transform 1 0 11010 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2121_
timestamp 1728341909
transform 1 0 11110 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2122_
timestamp 1728341909
transform 1 0 10810 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2123_
timestamp 1728341909
transform 1 0 10870 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2124_
timestamp 1728341909
transform 1 0 9330 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2125_
timestamp 1728341909
transform 1 0 9450 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2126_
timestamp 1728341909
transform -1 0 9890 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2127_
timestamp 1728341909
transform 1 0 9710 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2128_
timestamp 1728341909
transform 1 0 9670 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2129_
timestamp 1728341909
transform -1 0 8890 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2130_
timestamp 1728341909
transform 1 0 9570 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2131_
timestamp 1728341909
transform 1 0 9670 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2132_
timestamp 1728341909
transform 1 0 10130 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2133_
timestamp 1728341909
transform 1 0 10290 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2134_
timestamp 1728341909
transform -1 0 10070 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2135_
timestamp 1728341909
transform 1 0 10570 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2136_
timestamp 1728341909
transform -1 0 10530 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2137_
timestamp 1728341909
transform 1 0 10770 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2138_
timestamp 1728341909
transform -1 0 10870 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2139_
timestamp 1728341909
transform -1 0 10810 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2140_
timestamp 1728341909
transform -1 0 8290 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2141_
timestamp 1728341909
transform 1 0 8530 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2142_
timestamp 1728341909
transform 1 0 1850 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2143_
timestamp 1728341909
transform -1 0 2890 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2144_
timestamp 1728341909
transform -1 0 5990 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2145_
timestamp 1728341909
transform -1 0 6190 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2146_
timestamp 1728341909
transform 1 0 5490 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2147_
timestamp 1728341909
transform -1 0 6730 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2148_
timestamp 1728341909
transform 1 0 9630 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2149_
timestamp 1728341909
transform 1 0 8710 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2150_
timestamp 1728341909
transform -1 0 8470 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2151_
timestamp 1728341909
transform 1 0 8130 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2152_
timestamp 1728341909
transform -1 0 8970 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2153_
timestamp 1728341909
transform -1 0 9070 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2154_
timestamp 1728341909
transform 1 0 8810 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2155_
timestamp 1728341909
transform 1 0 7970 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2156_
timestamp 1728341909
transform -1 0 8250 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2157_
timestamp 1728341909
transform -1 0 8370 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2158_
timestamp 1728341909
transform 1 0 10290 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2159_
timestamp 1728341909
transform 1 0 5990 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2160_
timestamp 1728341909
transform -1 0 6350 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2161_
timestamp 1728341909
transform 1 0 6550 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2162_
timestamp 1728341909
transform -1 0 7890 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2163_
timestamp 1728341909
transform -1 0 8310 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2164_
timestamp 1728341909
transform 1 0 7070 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2165_
timestamp 1728341909
transform -1 0 7050 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2166_
timestamp 1728341909
transform -1 0 8110 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2167_
timestamp 1728341909
transform -1 0 7810 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2168_
timestamp 1728341909
transform -1 0 8070 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2169_
timestamp 1728341909
transform 1 0 8110 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2170_
timestamp 1728341909
transform -1 0 8330 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2171_
timestamp 1728341909
transform 1 0 8530 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2172_
timestamp 1728341909
transform -1 0 10390 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2173_
timestamp 1728341909
transform 1 0 10130 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2174_
timestamp 1728341909
transform 1 0 4350 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2175_
timestamp 1728341909
transform -1 0 3910 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2176_
timestamp 1728341909
transform -1 0 5370 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2177_
timestamp 1728341909
transform -1 0 6030 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2178_
timestamp 1728341909
transform -1 0 6290 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2179_
timestamp 1728341909
transform 1 0 6330 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2180_
timestamp 1728341909
transform 1 0 7130 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2181_
timestamp 1728341909
transform 1 0 7270 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2182_
timestamp 1728341909
transform -1 0 7130 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2183_
timestamp 1728341909
transform 1 0 6110 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2184_
timestamp 1728341909
transform 1 0 6430 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2185_
timestamp 1728341909
transform -1 0 6570 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2186_
timestamp 1728341909
transform -1 0 9010 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2187_
timestamp 1728341909
transform -1 0 9410 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2188_
timestamp 1728341909
transform 1 0 9010 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2189_
timestamp 1728341909
transform -1 0 8790 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2190_
timestamp 1728341909
transform 1 0 8470 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2191_
timestamp 1728341909
transform 1 0 8710 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2192_
timestamp 1728341909
transform 1 0 7270 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2193_
timestamp 1728341909
transform 1 0 7490 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2194_
timestamp 1728341909
transform -1 0 8610 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2195_
timestamp 1728341909
transform -1 0 8530 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2196_
timestamp 1728341909
transform 1 0 8570 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2197_
timestamp 1728341909
transform 1 0 8610 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2198_
timestamp 1728341909
transform -1 0 7210 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2199_
timestamp 1728341909
transform -1 0 7470 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2200_
timestamp 1728341909
transform 1 0 8990 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2201_
timestamp 1728341909
transform 1 0 8850 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2202_
timestamp 1728341909
transform -1 0 8650 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2203_
timestamp 1728341909
transform 1 0 8370 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2204_
timestamp 1728341909
transform -1 0 8370 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2205_
timestamp 1728341909
transform 1 0 8110 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2206_
timestamp 1728341909
transform -1 0 7990 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2207_
timestamp 1728341909
transform 1 0 8490 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2208_
timestamp 1728341909
transform -1 0 8250 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2209_
timestamp 1728341909
transform -1 0 7770 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2210_
timestamp 1728341909
transform 1 0 2710 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2211_
timestamp 1728341909
transform -1 0 7170 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2212_
timestamp 1728341909
transform -1 0 7430 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2213_
timestamp 1728341909
transform -1 0 7950 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2214_
timestamp 1728341909
transform 1 0 8510 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2215_
timestamp 1728341909
transform 1 0 9210 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2216_
timestamp 1728341909
transform 1 0 9190 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2217_
timestamp 1728341909
transform -1 0 9450 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2218_
timestamp 1728341909
transform 1 0 3890 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2219_
timestamp 1728341909
transform -1 0 2210 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2220_
timestamp 1728341909
transform -1 0 3630 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2221_
timestamp 1728341909
transform 1 0 4070 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2222_
timestamp 1728341909
transform 1 0 4290 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2223_
timestamp 1728341909
transform 1 0 4110 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2224_
timestamp 1728341909
transform -1 0 2790 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2225_
timestamp 1728341909
transform -1 0 5850 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2226_
timestamp 1728341909
transform 1 0 5970 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2227_
timestamp 1728341909
transform -1 0 6950 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2228_
timestamp 1728341909
transform 1 0 6690 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2229_
timestamp 1728341909
transform 1 0 7750 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2230_
timestamp 1728341909
transform -1 0 6150 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2231_
timestamp 1728341909
transform -1 0 6390 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2232_
timestamp 1728341909
transform 1 0 6810 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2233_
timestamp 1728341909
transform 1 0 7390 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2234_
timestamp 1728341909
transform 1 0 7290 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2235_
timestamp 1728341909
transform 1 0 9370 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2236_
timestamp 1728341909
transform 1 0 10430 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2237_
timestamp 1728341909
transform 1 0 9910 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2238_
timestamp 1728341909
transform -1 0 9830 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2239_
timestamp 1728341909
transform -1 0 5790 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2240_
timestamp 1728341909
transform 1 0 2650 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2241_
timestamp 1728341909
transform -1 0 4330 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2242_
timestamp 1728341909
transform -1 0 4550 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2243_
timestamp 1728341909
transform 1 0 3330 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2244_
timestamp 1728341909
transform 1 0 5090 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2245_
timestamp 1728341909
transform 1 0 7230 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2246_
timestamp 1728341909
transform 1 0 7250 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2247_
timestamp 1728341909
transform -1 0 3210 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2248_
timestamp 1728341909
transform 1 0 3390 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2249_
timestamp 1728341909
transform 1 0 5370 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2250_
timestamp 1728341909
transform 1 0 6630 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2251_
timestamp 1728341909
transform 1 0 7150 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2252_
timestamp 1728341909
transform -1 0 9590 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2253_
timestamp 1728341909
transform 1 0 9310 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2254_
timestamp 1728341909
transform 1 0 5590 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2255_
timestamp 1728341909
transform -1 0 6930 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2256_
timestamp 1728341909
transform 1 0 7090 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2257_
timestamp 1728341909
transform -1 0 3030 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2258_
timestamp 1728341909
transform -1 0 2990 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2259_
timestamp 1728341909
transform 1 0 3410 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2260_
timestamp 1728341909
transform 1 0 4590 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2261_
timestamp 1728341909
transform -1 0 5590 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2262_
timestamp 1728341909
transform 1 0 4770 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2263_
timestamp 1728341909
transform 1 0 4830 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2264_
timestamp 1728341909
transform -1 0 6130 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2265_
timestamp 1728341909
transform 1 0 3430 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2266_
timestamp 1728341909
transform 1 0 7470 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2267_
timestamp 1728341909
transform -1 0 5370 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2268_
timestamp 1728341909
transform -1 0 5610 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2269_
timestamp 1728341909
transform 1 0 5370 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2270_
timestamp 1728341909
transform -1 0 6210 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2271_
timestamp 1728341909
transform 1 0 5930 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2272_
timestamp 1728341909
transform 1 0 5530 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2273_
timestamp 1728341909
transform 1 0 5350 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2274_
timestamp 1728341909
transform 1 0 5110 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2275_
timestamp 1728341909
transform 1 0 5590 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2276_
timestamp 1728341909
transform -1 0 6230 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2277_
timestamp 1728341909
transform 1 0 7730 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2278_
timestamp 1728341909
transform -1 0 7670 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2279_
timestamp 1728341909
transform 1 0 6430 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2280_
timestamp 1728341909
transform -1 0 6450 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2281_
timestamp 1728341909
transform -1 0 6210 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2282_
timestamp 1728341909
transform 1 0 6490 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2283_
timestamp 1728341909
transform 1 0 7190 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2284_
timestamp 1728341909
transform 1 0 9150 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2285_
timestamp 1728341909
transform 1 0 9590 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2286_
timestamp 1728341909
transform -1 0 2490 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2287_
timestamp 1728341909
transform -1 0 1750 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2288_
timestamp 1728341909
transform -1 0 2190 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2289_
timestamp 1728341909
transform 1 0 2150 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2290_
timestamp 1728341909
transform -1 0 1710 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2291_
timestamp 1728341909
transform 1 0 1930 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2292_
timestamp 1728341909
transform 1 0 4050 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2293_
timestamp 1728341909
transform 1 0 4790 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2294_
timestamp 1728341909
transform 1 0 6010 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2295_
timestamp 1728341909
transform -1 0 2190 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2296_
timestamp 1728341909
transform 1 0 3630 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2297_
timestamp 1728341909
transform 1 0 2170 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2298_
timestamp 1728341909
transform 1 0 1930 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2299_
timestamp 1728341909
transform 1 0 3390 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2300_
timestamp 1728341909
transform 1 0 3130 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2301_
timestamp 1728341909
transform -1 0 3590 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2302_
timestamp 1728341909
transform 1 0 5070 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2303_
timestamp 1728341909
transform -1 0 5050 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2304_
timestamp 1728341909
transform 1 0 5290 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2305_
timestamp 1728341909
transform -1 0 1490 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2306_
timestamp 1728341909
transform 1 0 2390 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2307_
timestamp 1728341909
transform -1 0 5550 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2308_
timestamp 1728341909
transform -1 0 5550 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2309_
timestamp 1728341909
transform 1 0 4550 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2310_
timestamp 1728341909
transform 1 0 4310 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2311_
timestamp 1728341909
transform -1 0 3710 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2312_
timestamp 1728341909
transform -1 0 3950 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2313_
timestamp 1728341909
transform 1 0 5230 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2314_
timestamp 1728341909
transform 1 0 4410 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2315_
timestamp 1728341909
transform 1 0 5370 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2316_
timestamp 1728341909
transform -1 0 9810 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2317_
timestamp 1728341909
transform 1 0 11110 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2318_
timestamp 1728341909
transform -1 0 10810 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2319_
timestamp 1728341909
transform -1 0 10430 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2320_
timestamp 1728341909
transform 1 0 10590 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2321_
timestamp 1728341909
transform 1 0 10530 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2322_
timestamp 1728341909
transform 1 0 10430 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2323_
timestamp 1728341909
transform 1 0 6690 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2324_
timestamp 1728341909
transform 1 0 6890 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2325_
timestamp 1728341909
transform 1 0 9250 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2326_
timestamp 1728341909
transform -1 0 8790 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2327_
timestamp 1728341909
transform -1 0 9250 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2328_
timestamp 1728341909
transform -1 0 9490 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2329_
timestamp 1728341909
transform 1 0 9210 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2330_
timestamp 1728341909
transform -1 0 8970 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2331_
timestamp 1728341909
transform -1 0 9130 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2332_
timestamp 1728341909
transform 1 0 9110 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2333_
timestamp 1728341909
transform 1 0 9370 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2334_
timestamp 1728341909
transform -1 0 9570 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2335_
timestamp 1728341909
transform 1 0 5610 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2336_
timestamp 1728341909
transform 1 0 6130 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2337_
timestamp 1728341909
transform -1 0 5910 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2338_
timestamp 1728341909
transform -1 0 5850 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2339_
timestamp 1728341909
transform 1 0 10330 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2340_
timestamp 1728341909
transform -1 0 9210 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2341_
timestamp 1728341909
transform 1 0 9210 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2342_
timestamp 1728341909
transform 1 0 10070 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2343_
timestamp 1728341909
transform -1 0 9570 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2344_
timestamp 1728341909
transform 1 0 9670 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2345_
timestamp 1728341909
transform -1 0 6850 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2346_
timestamp 1728341909
transform 1 0 6710 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2347_
timestamp 1728341909
transform -1 0 7050 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2348_
timestamp 1728341909
transform 1 0 8050 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2349_
timestamp 1728341909
transform -1 0 7750 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2350_
timestamp 1728341909
transform 1 0 7470 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2351_
timestamp 1728341909
transform -1 0 5170 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2352_
timestamp 1728341909
transform 1 0 5770 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2353_
timestamp 1728341909
transform -1 0 4190 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2354_
timestamp 1728341909
transform 1 0 4670 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2355_
timestamp 1728341909
transform -1 0 4930 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2356_
timestamp 1728341909
transform 1 0 5870 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2357_
timestamp 1728341909
transform -1 0 5630 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2358_
timestamp 1728341909
transform 1 0 6910 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2359_
timestamp 1728341909
transform 1 0 6270 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2360_
timestamp 1728341909
transform 1 0 6510 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2361_
timestamp 1728341909
transform 1 0 7810 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2362_
timestamp 1728341909
transform 1 0 7330 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2363_
timestamp 1728341909
transform -1 0 7430 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2364_
timestamp 1728341909
transform 1 0 8050 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2365_
timestamp 1728341909
transform -1 0 7930 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2366_
timestamp 1728341909
transform 1 0 7690 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2367_
timestamp 1728341909
transform 1 0 7970 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2368_
timestamp 1728341909
transform 1 0 8190 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2369_
timestamp 1728341909
transform -1 0 9910 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2370_
timestamp 1728341909
transform 1 0 5330 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2371_
timestamp 1728341909
transform -1 0 8730 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2372_
timestamp 1728341909
transform -1 0 8470 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2373_
timestamp 1728341909
transform -1 0 8050 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2374_
timestamp 1728341909
transform 1 0 8050 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2375_
timestamp 1728341909
transform 1 0 6450 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2376_
timestamp 1728341909
transform 1 0 8410 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2377_
timestamp 1728341909
transform -1 0 8670 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2378_
timestamp 1728341909
transform -1 0 8970 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2379_
timestamp 1728341909
transform -1 0 6830 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2380_
timestamp 1728341909
transform -1 0 6970 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2381_
timestamp 1728341909
transform -1 0 6830 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2382_
timestamp 1728341909
transform -1 0 7910 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2383_
timestamp 1728341909
transform 1 0 7630 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2384_
timestamp 1728341909
transform 1 0 7730 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2385_
timestamp 1728341909
transform -1 0 7470 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2386_
timestamp 1728341909
transform -1 0 6590 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2387_
timestamp 1728341909
transform -1 0 6350 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2388_
timestamp 1728341909
transform -1 0 8910 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2389_
timestamp 1728341909
transform -1 0 8290 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2390_
timestamp 1728341909
transform -1 0 8230 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2391_
timestamp 1728341909
transform -1 0 9470 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2392_
timestamp 1728341909
transform 1 0 8230 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2393_
timestamp 1728341909
transform 1 0 8190 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2394_
timestamp 1728341909
transform 1 0 8830 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2395_
timestamp 1728341909
transform 1 0 8790 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2396_
timestamp 1728341909
transform 1 0 9070 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2397_
timestamp 1728341909
transform -1 0 9330 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2398_
timestamp 1728341909
transform 1 0 8710 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2399_
timestamp 1728341909
transform -1 0 7590 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2400_
timestamp 1728341909
transform 1 0 7330 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2401_
timestamp 1728341909
transform 1 0 8450 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2402_
timestamp 1728341909
transform -1 0 6390 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2403_
timestamp 1728341909
transform -1 0 6590 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2404_
timestamp 1728341909
transform -1 0 7550 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2405_
timestamp 1728341909
transform -1 0 7330 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2406_
timestamp 1728341909
transform 1 0 7050 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2407_
timestamp 1728341909
transform -1 0 6590 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2408_
timestamp 1728341909
transform -1 0 5890 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2409_
timestamp 1728341909
transform 1 0 6970 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2410_
timestamp 1728341909
transform -1 0 7250 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2411_
timestamp 1728341909
transform -1 0 6810 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2412_
timestamp 1728341909
transform -1 0 7470 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2413_
timestamp 1728341909
transform 1 0 6990 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2414_
timestamp 1728341909
transform 1 0 6810 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2415_
timestamp 1728341909
transform -1 0 8010 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2416_
timestamp 1728341909
transform 1 0 7750 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2417_
timestamp 1728341909
transform -1 0 8990 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2418_
timestamp 1728341909
transform -1 0 8770 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2419_
timestamp 1728341909
transform 1 0 7030 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2420_
timestamp 1728341909
transform 1 0 2190 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2421_
timestamp 1728341909
transform -1 0 9650 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2422_
timestamp 1728341909
transform 1 0 8230 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2423_
timestamp 1728341909
transform 1 0 8950 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2424_
timestamp 1728341909
transform 1 0 8730 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2425_
timestamp 1728341909
transform 1 0 3130 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2426_
timestamp 1728341909
transform 1 0 8710 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2427_
timestamp 1728341909
transform 1 0 8790 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2428_
timestamp 1728341909
transform 1 0 9190 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2429_
timestamp 1728341909
transform 1 0 9410 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2430_
timestamp 1728341909
transform 1 0 8770 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2431_
timestamp 1728341909
transform -1 0 9230 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2432_
timestamp 1728341909
transform 1 0 9450 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2433_
timestamp 1728341909
transform -1 0 9870 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2434_
timestamp 1728341909
transform -1 0 9950 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2435_
timestamp 1728341909
transform 1 0 4410 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2436_
timestamp 1728341909
transform 1 0 9170 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2437_
timestamp 1728341909
transform 1 0 10850 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2438_
timestamp 1728341909
transform -1 0 10910 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2439_
timestamp 1728341909
transform -1 0 10890 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2440_
timestamp 1728341909
transform 1 0 9010 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2441_
timestamp 1728341909
transform -1 0 6150 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2442_
timestamp 1728341909
transform -1 0 8230 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2443_
timestamp 1728341909
transform 1 0 3790 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2444_
timestamp 1728341909
transform -1 0 4670 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2445_
timestamp 1728341909
transform -1 0 8570 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2446_
timestamp 1728341909
transform 1 0 8210 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2447_
timestamp 1728341909
transform 1 0 8050 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2448_
timestamp 1728341909
transform 1 0 8450 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2449_
timestamp 1728341909
transform -1 0 8730 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2450_
timestamp 1728341909
transform -1 0 8930 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2451_
timestamp 1728341909
transform 1 0 3790 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2452_
timestamp 1728341909
transform 1 0 7570 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2453_
timestamp 1728341909
transform -1 0 6590 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2454_
timestamp 1728341909
transform -1 0 6310 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2455_
timestamp 1728341909
transform -1 0 6590 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2456_
timestamp 1728341909
transform -1 0 8710 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2457_
timestamp 1728341909
transform -1 0 8930 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2458_
timestamp 1728341909
transform -1 0 6770 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2459_
timestamp 1728341909
transform -1 0 3550 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2460_
timestamp 1728341909
transform 1 0 7070 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2461_
timestamp 1728341909
transform 1 0 6990 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2462_
timestamp 1728341909
transform -1 0 7270 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2463_
timestamp 1728341909
transform -1 0 7290 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2464_
timestamp 1728341909
transform 1 0 4450 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2465_
timestamp 1728341909
transform -1 0 7350 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2466_
timestamp 1728341909
transform -1 0 3330 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2467_
timestamp 1728341909
transform 1 0 6150 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2468_
timestamp 1728341909
transform -1 0 6270 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2469_
timestamp 1728341909
transform -1 0 6110 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2470_
timestamp 1728341909
transform -1 0 6370 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2471_
timestamp 1728341909
transform -1 0 8030 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2472_
timestamp 1728341909
transform -1 0 6050 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2473_
timestamp 1728341909
transform -1 0 5390 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2474_
timestamp 1728341909
transform -1 0 5310 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2475_
timestamp 1728341909
transform -1 0 7770 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2476_
timestamp 1728341909
transform -1 0 2690 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2477_
timestamp 1728341909
transform -1 0 5170 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2478_
timestamp 1728341909
transform 1 0 5250 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2479_
timestamp 1728341909
transform -1 0 7990 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2480_
timestamp 1728341909
transform 1 0 5890 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2481_
timestamp 1728341909
transform 1 0 4150 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2482_
timestamp 1728341909
transform -1 0 2430 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2483_
timestamp 1728341909
transform -1 0 4670 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2484_
timestamp 1728341909
transform -1 0 5710 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2485_
timestamp 1728341909
transform -1 0 6950 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2486_
timestamp 1728341909
transform 1 0 3070 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2487_
timestamp 1728341909
transform -1 0 5650 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2488_
timestamp 1728341909
transform 1 0 6410 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2489_
timestamp 1728341909
transform -1 0 6690 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2490_
timestamp 1728341909
transform 1 0 7670 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2491_
timestamp 1728341909
transform -1 0 7910 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2492_
timestamp 1728341909
transform -1 0 2850 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2493_
timestamp 1728341909
transform -1 0 5490 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2494_
timestamp 1728341909
transform -1 0 6570 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2495_
timestamp 1728341909
transform 1 0 6810 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2496_
timestamp 1728341909
transform 1 0 7530 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2497_
timestamp 1728341909
transform -1 0 7770 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2498_
timestamp 1728341909
transform -1 0 8750 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2499_
timestamp 1728341909
transform 1 0 8990 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2500_
timestamp 1728341909
transform -1 0 7610 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2501_
timestamp 1728341909
transform -1 0 6730 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2502_
timestamp 1728341909
transform -1 0 7590 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2503_
timestamp 1728341909
transform 1 0 11090 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2504_
timestamp 1728341909
transform -1 0 4530 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2505_
timestamp 1728341909
transform -1 0 5670 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2506_
timestamp 1728341909
transform -1 0 6690 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2507_
timestamp 1728341909
transform 1 0 5830 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2508_
timestamp 1728341909
transform 1 0 5630 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2509_
timestamp 1728341909
transform -1 0 8790 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2510_
timestamp 1728341909
transform -1 0 8050 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2511_
timestamp 1728341909
transform -1 0 7370 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2512_
timestamp 1728341909
transform 1 0 7070 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2513_
timestamp 1728341909
transform 1 0 6850 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2514_
timestamp 1728341909
transform 1 0 7010 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2515_
timestamp 1728341909
transform 1 0 10350 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2516_
timestamp 1728341909
transform 1 0 8490 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2517_
timestamp 1728341909
transform 1 0 10590 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2518_
timestamp 1728341909
transform -1 0 9690 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2519_
timestamp 1728341909
transform 1 0 9930 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2520_
timestamp 1728341909
transform -1 0 10390 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2521_
timestamp 1728341909
transform -1 0 8490 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2522_
timestamp 1728341909
transform 1 0 6050 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2523_
timestamp 1728341909
transform 1 0 5870 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2524_
timestamp 1728341909
transform 1 0 8250 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2525_
timestamp 1728341909
transform 1 0 6750 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2526_
timestamp 1728341909
transform -1 0 7750 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2527_
timestamp 1728341909
transform 1 0 7970 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2528_
timestamp 1728341909
transform -1 0 8030 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2529_
timestamp 1728341909
transform 1 0 7810 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2530_
timestamp 1728341909
transform -1 0 7770 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2531_
timestamp 1728341909
transform -1 0 7790 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2532_
timestamp 1728341909
transform 1 0 7790 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2533_
timestamp 1728341909
transform -1 0 5450 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2534_
timestamp 1728341909
transform -1 0 5870 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2535_
timestamp 1728341909
transform -1 0 7550 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2536_
timestamp 1728341909
transform 1 0 7350 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2537_
timestamp 1728341909
transform 1 0 7270 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2538_
timestamp 1728341909
transform 1 0 7990 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2539_
timestamp 1728341909
transform 1 0 5850 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2540_
timestamp 1728341909
transform 1 0 5570 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2541_
timestamp 1728341909
transform 1 0 6090 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2542_
timestamp 1728341909
transform -1 0 6630 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2543_
timestamp 1728341909
transform -1 0 6590 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2544_
timestamp 1728341909
transform 1 0 6130 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2545_
timestamp 1728341909
transform 1 0 6830 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2546_
timestamp 1728341909
transform 1 0 6090 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2547_
timestamp 1728341909
transform 1 0 6310 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2548_
timestamp 1728341909
transform 1 0 7090 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2549_
timestamp 1728341909
transform 1 0 7350 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2550_
timestamp 1728341909
transform -1 0 7510 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2551_
timestamp 1728341909
transform -1 0 6230 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2552_
timestamp 1728341909
transform -1 0 4790 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2553_
timestamp 1728341909
transform -1 0 5830 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2554_
timestamp 1728341909
transform -1 0 5550 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2555_
timestamp 1728341909
transform 1 0 5610 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2556_
timestamp 1728341909
transform 1 0 4990 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2557_
timestamp 1728341909
transform 1 0 5730 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2558_
timestamp 1728341909
transform -1 0 6370 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2559_
timestamp 1728341909
transform 1 0 6050 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2560_
timestamp 1728341909
transform 1 0 4310 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2561_
timestamp 1728341909
transform -1 0 5370 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2562_
timestamp 1728341909
transform 1 0 4990 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2563_
timestamp 1728341909
transform -1 0 4890 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2564_
timestamp 1728341909
transform -1 0 4550 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2565_
timestamp 1728341909
transform 1 0 4690 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2566_
timestamp 1728341909
transform -1 0 4910 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2567_
timestamp 1728341909
transform 1 0 5110 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2568_
timestamp 1728341909
transform 1 0 5250 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2569_
timestamp 1728341909
transform -1 0 4130 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2570_
timestamp 1728341909
transform 1 0 5150 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2571_
timestamp 1728341909
transform 1 0 4270 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2572_
timestamp 1728341909
transform -1 0 4390 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2573_
timestamp 1728341909
transform 1 0 4630 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2574_
timestamp 1728341909
transform 1 0 5350 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2575_
timestamp 1728341909
transform -1 0 4910 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2576_
timestamp 1728341909
transform 1 0 5090 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2577_
timestamp 1728341909
transform 1 0 4830 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2578_
timestamp 1728341909
transform -1 0 4770 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2579_
timestamp 1728341909
transform 1 0 4630 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__2580_
timestamp 1728341909
transform 1 0 4670 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2581_
timestamp 1728341909
transform -1 0 4110 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2582_
timestamp 1728341909
transform -1 0 3250 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2583_
timestamp 1728341909
transform 1 0 2190 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2584_
timestamp 1728341909
transform 1 0 3150 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2585_
timestamp 1728341909
transform -1 0 6310 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2586_
timestamp 1728341909
transform -1 0 3670 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2587_
timestamp 1728341909
transform -1 0 3410 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2588_
timestamp 1728341909
transform -1 0 2930 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2589_
timestamp 1728341909
transform -1 0 2930 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2590_
timestamp 1728341909
transform 1 0 3550 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__2591_
timestamp 1728341909
transform -1 0 3030 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2592_
timestamp 1728341909
transform 1 0 2530 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2593_
timestamp 1728341909
transform -1 0 2630 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2594_
timestamp 1728341909
transform -1 0 2650 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2595_
timestamp 1728341909
transform -1 0 3730 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__2596_
timestamp 1728341909
transform 1 0 3330 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2597_
timestamp 1728341909
transform 1 0 3270 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2598_
timestamp 1728341909
transform -1 0 3150 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2599_
timestamp 1728341909
transform -1 0 3150 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2600_
timestamp 1728341909
transform 1 0 2870 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2601_
timestamp 1728341909
transform -1 0 2430 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2602_
timestamp 1728341909
transform -1 0 2690 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2603_
timestamp 1728341909
transform -1 0 2290 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2604_
timestamp 1728341909
transform 1 0 2430 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2605_
timestamp 1728341909
transform -1 0 2430 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2606_
timestamp 1728341909
transform 1 0 2150 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2607_
timestamp 1728341909
transform -1 0 1510 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2608_
timestamp 1728341909
transform -1 0 1030 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2609_
timestamp 1728341909
transform 1 0 1990 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2610_
timestamp 1728341909
transform 1 0 1230 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2611_
timestamp 1728341909
transform -1 0 1210 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2612_
timestamp 1728341909
transform -1 0 950 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2613_
timestamp 1728341909
transform -1 0 1930 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2614_
timestamp 1728341909
transform -1 0 550 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2615_
timestamp 1728341909
transform 1 0 1730 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2616_
timestamp 1728341909
transform 1 0 1470 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2617_
timestamp 1728341909
transform -1 0 1470 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2618_
timestamp 1728341909
transform -1 0 1710 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2619_
timestamp 1728341909
transform 1 0 750 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2620_
timestamp 1728341909
transform -1 0 1270 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2621_
timestamp 1728341909
transform 1 0 1010 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2622_
timestamp 1728341909
transform -1 0 1230 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2623_
timestamp 1728341909
transform 1 0 970 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2624_
timestamp 1728341909
transform -1 0 510 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2625_
timestamp 1728341909
transform -1 0 2590 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2626_
timestamp 1728341909
transform 1 0 1610 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2627_
timestamp 1728341909
transform 1 0 1350 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2628_
timestamp 1728341909
transform 1 0 750 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2629_
timestamp 1728341909
transform -1 0 3350 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2630_
timestamp 1728341909
transform 1 0 4210 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2631_
timestamp 1728341909
transform -1 0 4870 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2632_
timestamp 1728341909
transform 1 0 10850 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2633_
timestamp 1728341909
transform 1 0 3850 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2634_
timestamp 1728341909
transform 1 0 8950 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2635_
timestamp 1728341909
transform -1 0 2230 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2636_
timestamp 1728341909
transform -1 0 9110 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2637_
timestamp 1728341909
transform 1 0 4310 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2638_
timestamp 1728341909
transform 1 0 4810 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2639_
timestamp 1728341909
transform -1 0 9890 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2640_
timestamp 1728341909
transform -1 0 9830 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2641_
timestamp 1728341909
transform 1 0 10130 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2642_
timestamp 1728341909
transform -1 0 9470 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2643_
timestamp 1728341909
transform 1 0 10870 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2644_
timestamp 1728341909
transform -1 0 9710 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2645_
timestamp 1728341909
transform -1 0 9670 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__2646_
timestamp 1728341909
transform 1 0 10070 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2647_
timestamp 1728341909
transform -1 0 8550 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2648_
timestamp 1728341909
transform -1 0 4130 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__2649_
timestamp 1728341909
transform -1 0 5770 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2650_
timestamp 1728341909
transform 1 0 9270 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2651_
timestamp 1728341909
transform -1 0 5650 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2652_
timestamp 1728341909
transform -1 0 7810 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2653_
timestamp 1728341909
transform -1 0 7710 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2654_
timestamp 1728341909
transform 1 0 4630 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2655_
timestamp 1728341909
transform -1 0 5410 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2656_
timestamp 1728341909
transform -1 0 5990 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2657_
timestamp 1728341909
transform -1 0 6730 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2658_
timestamp 1728341909
transform 1 0 6230 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2659_
timestamp 1728341909
transform 1 0 6930 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2660_
timestamp 1728341909
transform -1 0 7210 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2661_
timestamp 1728341909
transform -1 0 4430 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2662_
timestamp 1728341909
transform 1 0 4390 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2663_
timestamp 1728341909
transform 1 0 6310 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2664_
timestamp 1728341909
transform -1 0 6570 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2665_
timestamp 1728341909
transform 1 0 7070 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2666_
timestamp 1728341909
transform 1 0 6810 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2667_
timestamp 1728341909
transform 1 0 7550 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2668_
timestamp 1728341909
transform 1 0 7290 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2669_
timestamp 1728341909
transform 1 0 7950 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2670_
timestamp 1728341909
transform -1 0 4170 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2671_
timestamp 1728341909
transform -1 0 5290 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__2672_
timestamp 1728341909
transform 1 0 5190 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2673_
timestamp 1728341909
transform 1 0 7150 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2674_
timestamp 1728341909
transform -1 0 7370 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2675_
timestamp 1728341909
transform 1 0 7610 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2676_
timestamp 1728341909
transform -1 0 7550 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2677_
timestamp 1728341909
transform 1 0 7730 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2678_
timestamp 1728341909
transform 1 0 7690 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2679_
timestamp 1728341909
transform 1 0 4130 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2680_
timestamp 1728341909
transform -1 0 4390 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2681_
timestamp 1728341909
transform 1 0 6090 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2682_
timestamp 1728341909
transform 1 0 6710 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2683_
timestamp 1728341909
transform 1 0 4050 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2684_
timestamp 1728341909
transform -1 0 5710 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2685_
timestamp 1728341909
transform 1 0 5430 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2686_
timestamp 1728341909
transform -1 0 6850 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2687_
timestamp 1728341909
transform 1 0 7310 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2688_
timestamp 1728341909
transform -1 0 7450 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2689_
timestamp 1728341909
transform 1 0 6470 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2690_
timestamp 1728341909
transform 1 0 6550 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2691_
timestamp 1728341909
transform 1 0 7050 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2692_
timestamp 1728341909
transform -1 0 7190 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2693_
timestamp 1728341909
transform 1 0 5030 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2694_
timestamp 1728341909
transform -1 0 5170 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2695_
timestamp 1728341909
transform 1 0 6610 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2696_
timestamp 1728341909
transform 1 0 6550 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2697_
timestamp 1728341909
transform 1 0 6970 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2698_
timestamp 1728341909
transform 1 0 6870 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2699_
timestamp 1728341909
transform -1 0 6310 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2700_
timestamp 1728341909
transform 1 0 5370 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2701_
timestamp 1728341909
transform -1 0 5450 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2702_
timestamp 1728341909
transform -1 0 5530 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2703_
timestamp 1728341909
transform -1 0 5550 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2704_
timestamp 1728341909
transform 1 0 5610 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2705_
timestamp 1728341909
transform 1 0 5870 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2706_
timestamp 1728341909
transform -1 0 6130 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2707_
timestamp 1728341909
transform -1 0 5870 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2708_
timestamp 1728341909
transform -1 0 2270 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2709_
timestamp 1728341909
transform -1 0 4930 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2710_
timestamp 1728341909
transform -1 0 4850 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2711_
timestamp 1728341909
transform -1 0 5050 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2712_
timestamp 1728341909
transform -1 0 5630 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2713_
timestamp 1728341909
transform -1 0 5770 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2714_
timestamp 1728341909
transform -1 0 6070 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2715_
timestamp 1728341909
transform 1 0 5790 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2716_
timestamp 1728341909
transform -1 0 6630 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2717_
timestamp 1728341909
transform 1 0 6570 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2718_
timestamp 1728341909
transform 1 0 6150 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2719_
timestamp 1728341909
transform -1 0 6310 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2720_
timestamp 1728341909
transform 1 0 4610 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2721_
timestamp 1728341909
transform 1 0 4890 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2722_
timestamp 1728341909
transform 1 0 5130 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2723_
timestamp 1728341909
transform -1 0 5390 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2724_
timestamp 1728341909
transform 1 0 6110 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2725_
timestamp 1728341909
transform 1 0 6350 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2726_
timestamp 1728341909
transform -1 0 6110 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__2727_
timestamp 1728341909
transform 1 0 5810 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__2728_
timestamp 1728341909
transform -1 0 4290 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2729_
timestamp 1728341909
transform -1 0 4150 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2730_
timestamp 1728341909
transform -1 0 5190 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2731_
timestamp 1728341909
transform -1 0 5310 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2732_
timestamp 1728341909
transform -1 0 5610 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2733_
timestamp 1728341909
transform -1 0 5870 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2734_
timestamp 1728341909
transform -1 0 5190 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2735_
timestamp 1728341909
transform 1 0 5390 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2736_
timestamp 1728341909
transform -1 0 8310 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__2737_
timestamp 1728341909
transform 1 0 3710 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2738_
timestamp 1728341909
transform 1 0 3890 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2739_
timestamp 1728341909
transform -1 0 3710 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2740_
timestamp 1728341909
transform -1 0 3650 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2741_
timestamp 1728341909
transform -1 0 3990 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2742_
timestamp 1728341909
transform -1 0 4130 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2743_
timestamp 1728341909
transform 1 0 4870 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2744_
timestamp 1728341909
transform 1 0 4610 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__2745_
timestamp 1728341909
transform 1 0 5090 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2746_
timestamp 1728341909
transform 1 0 4590 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2747_
timestamp 1728341909
transform 1 0 5510 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2748_
timestamp 1728341909
transform -1 0 4910 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2749_
timestamp 1728341909
transform -1 0 5270 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2750_
timestamp 1728341909
transform -1 0 5370 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2751_
timestamp 1728341909
transform 1 0 4350 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2752_
timestamp 1728341909
transform 1 0 3850 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2753_
timestamp 1728341909
transform -1 0 3390 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2754_
timestamp 1728341909
transform -1 0 2970 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2755_
timestamp 1728341909
transform 1 0 3230 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2756_
timestamp 1728341909
transform -1 0 3610 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2757_
timestamp 1728341909
transform -1 0 3630 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2758_
timestamp 1728341909
transform -1 0 3610 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2759_
timestamp 1728341909
transform -1 0 3490 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2760_
timestamp 1728341909
transform -1 0 3530 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2761_
timestamp 1728341909
transform -1 0 3670 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2762_
timestamp 1728341909
transform -1 0 3430 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2763_
timestamp 1728341909
transform 1 0 2990 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__2764_
timestamp 1728341909
transform 1 0 3270 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__2765_
timestamp 1728341909
transform -1 0 2590 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2766_
timestamp 1728341909
transform 1 0 3670 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__2767_
timestamp 1728341909
transform -1 0 4370 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2768_
timestamp 1728341909
transform 1 0 4450 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2769_
timestamp 1728341909
transform 1 0 5110 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2770_
timestamp 1728341909
transform -1 0 4610 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2771_
timestamp 1728341909
transform -1 0 4890 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2772_
timestamp 1728341909
transform -1 0 4870 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2773_
timestamp 1728341909
transform 1 0 2630 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2774_
timestamp 1728341909
transform -1 0 2490 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__2775_
timestamp 1728341909
transform 1 0 3850 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2776_
timestamp 1728341909
transform 1 0 4370 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2777_
timestamp 1728341909
transform 1 0 5110 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2778_
timestamp 1728341909
transform -1 0 4610 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2779_
timestamp 1728341909
transform 1 0 3930 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__2780_
timestamp 1728341909
transform 1 0 2710 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__2781_
timestamp 1728341909
transform -1 0 3930 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2782_
timestamp 1728341909
transform -1 0 2730 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2783_
timestamp 1728341909
transform 1 0 2430 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2784_
timestamp 1728341909
transform 1 0 510 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2785_
timestamp 1728341909
transform -1 0 2210 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2786_
timestamp 1728341909
transform 1 0 2470 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2787_
timestamp 1728341909
transform -1 0 2890 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2788_
timestamp 1728341909
transform -1 0 2390 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2789_
timestamp 1728341909
transform -1 0 3690 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2790_
timestamp 1728341909
transform 1 0 3170 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2791_
timestamp 1728341909
transform -1 0 2910 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2792_
timestamp 1728341909
transform -1 0 2810 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2793_
timestamp 1728341909
transform -1 0 2230 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__2794_
timestamp 1728341909
transform 1 0 2110 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2795_
timestamp 1728341909
transform 1 0 750 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2796_
timestamp 1728341909
transform 1 0 1690 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2797_
timestamp 1728341909
transform -1 0 1970 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2798_
timestamp 1728341909
transform 1 0 1190 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2799_
timestamp 1728341909
transform -1 0 1470 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2800_
timestamp 1728341909
transform -1 0 1730 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2801_
timestamp 1728341909
transform 1 0 1690 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2802_
timestamp 1728341909
transform 1 0 1770 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2803_
timestamp 1728341909
transform 1 0 3250 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2804_
timestamp 1728341909
transform -1 0 410 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__2805_
timestamp 1728341909
transform 1 0 6950 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2806_
timestamp 1728341909
transform -1 0 5370 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2807_
timestamp 1728341909
transform -1 0 4970 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2808_
timestamp 1728341909
transform 1 0 3890 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2809_
timestamp 1728341909
transform -1 0 4350 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2810_
timestamp 1728341909
transform -1 0 4710 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2811_
timestamp 1728341909
transform -1 0 4570 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2812_
timestamp 1728341909
transform 1 0 4190 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2813_
timestamp 1728341909
transform 1 0 3950 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__2814_
timestamp 1728341909
transform 1 0 4070 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__2815_
timestamp 1728341909
transform -1 0 4150 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2816_
timestamp 1728341909
transform 1 0 2450 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2817_
timestamp 1728341909
transform -1 0 2730 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__2818_
timestamp 1728341909
transform 1 0 2690 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2819_
timestamp 1728341909
transform 1 0 3130 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2820_
timestamp 1728341909
transform 1 0 3370 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2821_
timestamp 1728341909
transform -1 0 3910 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2822_
timestamp 1728341909
transform -1 0 4710 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2823_
timestamp 1728341909
transform -1 0 1690 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2824_
timestamp 1728341909
transform 1 0 510 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__2825_
timestamp 1728341909
transform 1 0 490 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2826_
timestamp 1728341909
transform -1 0 650 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__2827_
timestamp 1728341909
transform 1 0 1690 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2828_
timestamp 1728341909
transform -1 0 1970 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2829_
timestamp 1728341909
transform 1 0 1210 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2830_
timestamp 1728341909
transform -1 0 1470 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2831_
timestamp 1728341909
transform -1 0 1490 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__2832_
timestamp 1728341909
transform 1 0 1990 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2833_
timestamp 1728341909
transform -1 0 1010 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__2834_
timestamp 1728341909
transform 1 0 830 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__2835_
timestamp 1728341909
transform 1 0 1070 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__2836_
timestamp 1728341909
transform 1 0 1290 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__2837_
timestamp 1728341909
transform 1 0 1610 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__2838_
timestamp 1728341909
transform -1 0 1490 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__2839_
timestamp 1728341909
transform 1 0 770 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__2840_
timestamp 1728341909
transform 1 0 1210 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2841_
timestamp 1728341909
transform 1 0 2010 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2842_
timestamp 1728341909
transform -1 0 1670 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2843_
timestamp 1728341909
transform -1 0 1770 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2844_
timestamp 1728341909
transform -1 0 1530 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__2845_
timestamp 1728341909
transform -1 0 1470 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2846_
timestamp 1728341909
transform 1 0 1250 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2847_
timestamp 1728341909
transform -1 0 1250 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__2848_
timestamp 1728341909
transform -1 0 1230 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2849_
timestamp 1728341909
transform -1 0 1530 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2850_
timestamp 1728341909
transform -1 0 1450 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2851_
timestamp 1728341909
transform -1 0 990 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2852_
timestamp 1728341909
transform -1 0 1050 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2853_
timestamp 1728341909
transform -1 0 2250 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2854_
timestamp 1728341909
transform 1 0 730 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__2855_
timestamp 1728341909
transform 1 0 2410 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__2856_
timestamp 1728341909
transform -1 0 1930 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__2857_
timestamp 1728341909
transform -1 0 2330 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__2858_
timestamp 1728341909
transform -1 0 2230 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__2859_
timestamp 1728341909
transform -1 0 810 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2860_
timestamp 1728341909
transform 1 0 490 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2861_
timestamp 1728341909
transform -1 0 50 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2862_
timestamp 1728341909
transform -1 0 1010 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__2863_
timestamp 1728341909
transform 1 0 250 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__2864_
timestamp 1728341909
transform -1 0 290 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__2865_
timestamp 1728341909
transform 1 0 4410 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2866_
timestamp 1728341909
transform 1 0 4430 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2867_
timestamp 1728341909
transform 1 0 5530 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2868_
timestamp 1728341909
transform -1 0 2910 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2869_
timestamp 1728341909
transform -1 0 3190 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2870_
timestamp 1728341909
transform -1 0 2250 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2871_
timestamp 1728341909
transform 1 0 2270 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2872_
timestamp 1728341909
transform -1 0 4550 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2873_
timestamp 1728341909
transform 1 0 4290 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2874_
timestamp 1728341909
transform -1 0 4090 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2875_
timestamp 1728341909
transform -1 0 1650 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2876_
timestamp 1728341909
transform -1 0 790 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2877_
timestamp 1728341909
transform -1 0 3450 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2878_
timestamp 1728341909
transform -1 0 3890 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2879_
timestamp 1728341909
transform -1 0 1230 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2880_
timestamp 1728341909
transform 1 0 1410 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2881_
timestamp 1728341909
transform -1 0 1730 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2882_
timestamp 1728341909
transform -1 0 2410 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2883_
timestamp 1728341909
transform 1 0 4410 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2884_
timestamp 1728341909
transform 1 0 4130 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2885_
timestamp 1728341909
transform 1 0 3070 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2886_
timestamp 1728341909
transform 1 0 4630 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2887_
timestamp 1728341909
transform 1 0 5090 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2888_
timestamp 1728341909
transform 1 0 3350 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2889_
timestamp 1728341909
transform 1 0 3570 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2890_
timestamp 1728341909
transform -1 0 4350 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2891_
timestamp 1728341909
transform -1 0 4090 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2892_
timestamp 1728341909
transform -1 0 1950 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2893_
timestamp 1728341909
transform 1 0 3630 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2894_
timestamp 1728341909
transform 1 0 3830 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2895_
timestamp 1728341909
transform 1 0 4410 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2896_
timestamp 1728341909
transform -1 0 3810 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2897_
timestamp 1728341909
transform -1 0 5810 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2898_
timestamp 1728341909
transform 1 0 5130 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2899_
timestamp 1728341909
transform 1 0 5090 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2900_
timestamp 1728341909
transform 1 0 5350 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2901_
timestamp 1728341909
transform -1 0 4830 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2902_
timestamp 1728341909
transform -1 0 1490 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2903_
timestamp 1728341909
transform 1 0 2150 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2904_
timestamp 1728341909
transform 1 0 2410 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2905_
timestamp 1728341909
transform 1 0 1210 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2906_
timestamp 1728341909
transform 1 0 990 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2907_
timestamp 1728341909
transform 1 0 1190 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2908_
timestamp 1728341909
transform -1 0 1510 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2909_
timestamp 1728341909
transform -1 0 1730 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2910_
timestamp 1728341909
transform -1 0 1510 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2911_
timestamp 1728341909
transform -1 0 1510 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2912_
timestamp 1728341909
transform -1 0 2430 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2913_
timestamp 1728341909
transform -1 0 1670 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2914_
timestamp 1728341909
transform 1 0 2190 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2915_
timestamp 1728341909
transform 1 0 1970 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2916_
timestamp 1728341909
transform 1 0 1650 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2917_
timestamp 1728341909
transform -1 0 1730 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2918_
timestamp 1728341909
transform 1 0 1670 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2919_
timestamp 1728341909
transform -1 0 2210 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2920_
timestamp 1728341909
transform -1 0 1930 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2921_
timestamp 1728341909
transform -1 0 1990 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2922_
timestamp 1728341909
transform -1 0 1910 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2923_
timestamp 1728341909
transform -1 0 1950 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2924_
timestamp 1728341909
transform -1 0 2910 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2925_
timestamp 1728341909
transform 1 0 3390 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2926_
timestamp 1728341909
transform -1 0 2370 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2927_
timestamp 1728341909
transform -1 0 2410 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2928_
timestamp 1728341909
transform 1 0 4550 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2929_
timestamp 1728341909
transform 1 0 3390 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2930_
timestamp 1728341909
transform -1 0 2670 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2931_
timestamp 1728341909
transform -1 0 2910 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2932_
timestamp 1728341909
transform 1 0 3110 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2933_
timestamp 1728341909
transform -1 0 2670 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2934_
timestamp 1728341909
transform 1 0 2890 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2935_
timestamp 1728341909
transform -1 0 1270 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2936_
timestamp 1728341909
transform -1 0 810 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2937_
timestamp 1728341909
transform 1 0 530 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2938_
timestamp 1728341909
transform 1 0 1690 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2939_
timestamp 1728341909
transform -1 0 1470 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2940_
timestamp 1728341909
transform 1 0 3130 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2941_
timestamp 1728341909
transform 1 0 3130 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2942_
timestamp 1728341909
transform -1 0 3350 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2943_
timestamp 1728341909
transform -1 0 3190 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2944_
timestamp 1728341909
transform -1 0 3690 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2945_
timestamp 1728341909
transform 1 0 3130 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2946_
timestamp 1728341909
transform 1 0 3570 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2947_
timestamp 1728341909
transform 1 0 3150 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2948_
timestamp 1728341909
transform -1 0 4150 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2949_
timestamp 1728341909
transform 1 0 3110 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2950_
timestamp 1728341909
transform 1 0 2430 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2951_
timestamp 1728341909
transform -1 0 2670 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2952_
timestamp 1728341909
transform -1 0 2950 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2953_
timestamp 1728341909
transform -1 0 2150 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2954_
timestamp 1728341909
transform -1 0 2390 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2955_
timestamp 1728341909
transform 1 0 2970 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2956_
timestamp 1728341909
transform 1 0 3210 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2957_
timestamp 1728341909
transform 1 0 3710 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2958_
timestamp 1728341909
transform 1 0 2150 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2959_
timestamp 1728341909
transform 1 0 3430 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2960_
timestamp 1728341909
transform 1 0 3550 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2961_
timestamp 1728341909
transform 1 0 2670 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2962_
timestamp 1728341909
transform 1 0 2410 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2963_
timestamp 1728341909
transform 1 0 2930 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2964_
timestamp 1728341909
transform 1 0 2670 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2965_
timestamp 1728341909
transform -1 0 5750 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2966_
timestamp 1728341909
transform 1 0 4070 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2967_
timestamp 1728341909
transform -1 0 4550 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2968_
timestamp 1728341909
transform -1 0 4790 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2969_
timestamp 1728341909
transform -1 0 1290 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2970_
timestamp 1728341909
transform -1 0 1470 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2971_
timestamp 1728341909
transform -1 0 1490 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2972_
timestamp 1728341909
transform -1 0 1230 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2973_
timestamp 1728341909
transform -1 0 990 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2974_
timestamp 1728341909
transform -1 0 1730 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2975_
timestamp 1728341909
transform -1 0 1950 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2976_
timestamp 1728341909
transform 1 0 3830 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2977_
timestamp 1728341909
transform -1 0 4390 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2978_
timestamp 1728341909
transform 1 0 4110 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2979_
timestamp 1728341909
transform 1 0 1490 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2980_
timestamp 1728341909
transform -1 0 970 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2981_
timestamp 1728341909
transform -1 0 730 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2982_
timestamp 1728341909
transform 1 0 2170 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2983_
timestamp 1728341909
transform -1 0 490 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2984_
timestamp 1728341909
transform -1 0 270 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2985_
timestamp 1728341909
transform -1 0 50 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2986_
timestamp 1728341909
transform -1 0 310 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2987_
timestamp 1728341909
transform -1 0 570 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2988_
timestamp 1728341909
transform -1 0 530 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2989_
timestamp 1728341909
transform 1 0 290 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2990_
timestamp 1728341909
transform 1 0 30 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2991_
timestamp 1728341909
transform -1 0 310 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2992_
timestamp 1728341909
transform -1 0 1970 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2993_
timestamp 1728341909
transform -1 0 1010 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2994_
timestamp 1728341909
transform -1 0 770 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2995_
timestamp 1728341909
transform 1 0 550 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2996_
timestamp 1728341909
transform -1 0 490 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2997_
timestamp 1728341909
transform -1 0 810 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2998_
timestamp 1728341909
transform -1 0 50 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2999_
timestamp 1728341909
transform -1 0 290 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__3000_
timestamp 1728341909
transform -1 0 50 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__3001_
timestamp 1728341909
transform -1 0 50 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__3002_
timestamp 1728341909
transform -1 0 530 0 1 730
box -12 -8 32 252
use FILL  FILL_1__3003_
timestamp 1728341909
transform -1 0 50 0 1 730
box -12 -8 32 252
use FILL  FILL_1__3004_
timestamp 1728341909
transform -1 0 790 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__3005_
timestamp 1728341909
transform 1 0 750 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__3006_
timestamp 1728341909
transform -1 0 50 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__3007_
timestamp 1728341909
transform 1 0 1750 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3008_
timestamp 1728341909
transform -1 0 1010 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__3009_
timestamp 1728341909
transform -1 0 1270 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__3010_
timestamp 1728341909
transform -1 0 1270 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__3011_
timestamp 1728341909
transform -1 0 1030 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__3012_
timestamp 1728341909
transform -1 0 1410 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__3013_
timestamp 1728341909
transform -1 0 1190 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__3014_
timestamp 1728341909
transform 1 0 990 0 1 250
box -12 -8 32 252
use FILL  FILL_1__3015_
timestamp 1728341909
transform -1 0 1490 0 1 250
box -12 -8 32 252
use FILL  FILL_1__3016_
timestamp 1728341909
transform -1 0 1250 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__3017_
timestamp 1728341909
transform -1 0 1230 0 1 250
box -12 -8 32 252
use FILL  FILL_1__3018_
timestamp 1728341909
transform 1 0 1010 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__3019_
timestamp 1728341909
transform -1 0 1010 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__3020_
timestamp 1728341909
transform -1 0 3650 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3021_
timestamp 1728341909
transform -1 0 5910 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__3022_
timestamp 1728341909
transform 1 0 2750 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3023_
timestamp 1728341909
transform 1 0 2770 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3024_
timestamp 1728341909
transform 1 0 3750 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3025_
timestamp 1728341909
transform -1 0 4170 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__3026_
timestamp 1728341909
transform -1 0 3030 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3027_
timestamp 1728341909
transform -1 0 3430 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__3028_
timestamp 1728341909
transform -1 0 3950 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3029_
timestamp 1728341909
transform -1 0 4450 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3030_
timestamp 1728341909
transform 1 0 3430 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__3031_
timestamp 1728341909
transform -1 0 3710 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__3032_
timestamp 1728341909
transform -1 0 2510 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3033_
timestamp 1728341909
transform -1 0 2530 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3034_
timestamp 1728341909
transform 1 0 2670 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__3035_
timestamp 1728341909
transform -1 0 2930 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__3036_
timestamp 1728341909
transform 1 0 3250 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3037_
timestamp 1728341909
transform -1 0 3690 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__3038_
timestamp 1728341909
transform -1 0 3250 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3039_
timestamp 1728341909
transform 1 0 2990 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3040_
timestamp 1728341909
transform 1 0 2130 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__3041_
timestamp 1728341909
transform 1 0 2670 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__3042_
timestamp 1728341909
transform 1 0 7430 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__3043_
timestamp 1728341909
transform 1 0 6270 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__3044_
timestamp 1728341909
transform 1 0 5290 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__3045_
timestamp 1728341909
transform 1 0 5710 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3046_
timestamp 1728341909
transform 1 0 5430 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__3047_
timestamp 1728341909
transform 1 0 4770 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__3048_
timestamp 1728341909
transform 1 0 5110 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__3049_
timestamp 1728341909
transform 1 0 5810 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3050_
timestamp 1728341909
transform -1 0 6830 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3051_
timestamp 1728341909
transform -1 0 6290 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__3052_
timestamp 1728341909
transform 1 0 6330 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3053_
timestamp 1728341909
transform 1 0 6070 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3054_
timestamp 1728341909
transform 1 0 5810 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3055_
timestamp 1728341909
transform -1 0 5910 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3056_
timestamp 1728341909
transform 1 0 4570 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__3057_
timestamp 1728341909
transform 1 0 4330 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__3058_
timestamp 1728341909
transform -1 0 4450 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3059_
timestamp 1728341909
transform 1 0 4270 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__3060_
timestamp 1728341909
transform -1 0 4250 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__3061_
timestamp 1728341909
transform 1 0 3950 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3062_
timestamp 1728341909
transform -1 0 4770 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__3063_
timestamp 1728341909
transform 1 0 4510 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__3064_
timestamp 1728341909
transform 1 0 5970 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__3065_
timestamp 1728341909
transform 1 0 5750 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__3066_
timestamp 1728341909
transform -1 0 5750 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3067_
timestamp 1728341909
transform -1 0 5890 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__3068_
timestamp 1728341909
transform -1 0 6930 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3069_
timestamp 1728341909
transform -1 0 6430 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3070_
timestamp 1728341909
transform 1 0 6070 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3071_
timestamp 1728341909
transform -1 0 6350 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3072_
timestamp 1728341909
transform 1 0 6550 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__3073_
timestamp 1728341909
transform 1 0 6310 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__3074_
timestamp 1728341909
transform 1 0 370 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__3075_
timestamp 1728341909
transform -1 0 530 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__3076_
timestamp 1728341909
transform -1 0 4230 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3077_
timestamp 1728341909
transform 1 0 1970 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3078_
timestamp 1728341909
transform -1 0 5470 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3079_
timestamp 1728341909
transform 1 0 5010 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3080_
timestamp 1728341909
transform 1 0 4210 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3081_
timestamp 1728341909
transform 1 0 5850 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__3082_
timestamp 1728341909
transform -1 0 6850 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__3083_
timestamp 1728341909
transform 1 0 6010 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__3084_
timestamp 1728341909
transform -1 0 5690 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3085_
timestamp 1728341909
transform -1 0 4970 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3086_
timestamp 1728341909
transform 1 0 5450 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3087_
timestamp 1728341909
transform -1 0 5050 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__3088_
timestamp 1728341909
transform -1 0 5590 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__3089_
timestamp 1728341909
transform -1 0 5550 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__3090_
timestamp 1728341909
transform 1 0 4730 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3091_
timestamp 1728341909
transform -1 0 4690 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3092_
timestamp 1728341909
transform 1 0 5550 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__3093_
timestamp 1728341909
transform -1 0 3950 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__3094_
timestamp 1728341909
transform 1 0 4390 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__3095_
timestamp 1728341909
transform 1 0 4690 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__3096_
timestamp 1728341909
transform 1 0 4670 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__3097_
timestamp 1728341909
transform 1 0 4910 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__3098_
timestamp 1728341909
transform -1 0 5010 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__3099_
timestamp 1728341909
transform 1 0 5150 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__3100_
timestamp 1728341909
transform -1 0 5550 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__3101_
timestamp 1728341909
transform 1 0 5090 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__3102_
timestamp 1728341909
transform 1 0 4610 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__3103_
timestamp 1728341909
transform 1 0 4830 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__3104_
timestamp 1728341909
transform -1 0 4970 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3105_
timestamp 1728341909
transform 1 0 5290 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__3106_
timestamp 1728341909
transform 1 0 8470 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__3107_
timestamp 1728341909
transform 1 0 8230 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__3108_
timestamp 1728341909
transform 1 0 7990 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__3109_
timestamp 1728341909
transform -1 0 8530 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3110_
timestamp 1728341909
transform -1 0 8290 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3111_
timestamp 1728341909
transform 1 0 4470 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3112_
timestamp 1728341909
transform 1 0 4710 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3113_
timestamp 1728341909
transform -1 0 1230 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3114_
timestamp 1728341909
transform 1 0 730 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3115_
timestamp 1728341909
transform 1 0 4410 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__3116_
timestamp 1728341909
transform -1 0 4030 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3117_
timestamp 1728341909
transform -1 0 290 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__3118_
timestamp 1728341909
transform -1 0 50 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__3119_
timestamp 1728341909
transform -1 0 4890 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__3120_
timestamp 1728341909
transform 1 0 4390 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3121_
timestamp 1728341909
transform 1 0 5130 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__3122_
timestamp 1728341909
transform -1 0 4430 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3123_
timestamp 1728341909
transform -1 0 3690 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3124_
timestamp 1728341909
transform -1 0 3910 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3125_
timestamp 1728341909
transform -1 0 3650 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3126_
timestamp 1728341909
transform 1 0 4670 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3127_
timestamp 1728341909
transform 1 0 4690 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3128_
timestamp 1728341909
transform 1 0 4610 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__3129_
timestamp 1728341909
transform 1 0 3690 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__3130_
timestamp 1728341909
transform -1 0 1790 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3131_
timestamp 1728341909
transform -1 0 1290 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3132_
timestamp 1728341909
transform 1 0 1010 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3133_
timestamp 1728341909
transform 1 0 3870 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3134_
timestamp 1728341909
transform 1 0 3450 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3135_
timestamp 1728341909
transform 1 0 3190 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3136_
timestamp 1728341909
transform 1 0 3670 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3137_
timestamp 1728341909
transform 1 0 3930 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3138_
timestamp 1728341909
transform -1 0 3970 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3139_
timestamp 1728341909
transform 1 0 1030 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3140_
timestamp 1728341909
transform 1 0 770 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3141_
timestamp 1728341909
transform -1 0 3950 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3142_
timestamp 1728341909
transform 1 0 3710 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3143_
timestamp 1728341909
transform -1 0 4150 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3144_
timestamp 1728341909
transform -1 0 3430 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3145_
timestamp 1728341909
transform 1 0 3170 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3146_
timestamp 1728341909
transform -1 0 3250 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3147_
timestamp 1728341909
transform 1 0 3490 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3148_
timestamp 1728341909
transform -1 0 3450 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3149_
timestamp 1728341909
transform -1 0 3430 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__3150_
timestamp 1728341909
transform 1 0 2010 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3151_
timestamp 1728341909
transform -1 0 2250 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3152_
timestamp 1728341909
transform 1 0 7490 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3153_
timestamp 1728341909
transform 1 0 4410 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3154_
timestamp 1728341909
transform -1 0 750 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3155_
timestamp 1728341909
transform 1 0 970 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3156_
timestamp 1728341909
transform 1 0 2930 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3157_
timestamp 1728341909
transform -1 0 2710 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3158_
timestamp 1728341909
transform 1 0 1930 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3159_
timestamp 1728341909
transform 1 0 2470 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3160_
timestamp 1728341909
transform 1 0 3090 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3161_
timestamp 1728341909
transform -1 0 2630 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3162_
timestamp 1728341909
transform -1 0 2410 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3163_
timestamp 1728341909
transform -1 0 1510 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3164_
timestamp 1728341909
transform 1 0 1210 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3165_
timestamp 1728341909
transform -1 0 290 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3166_
timestamp 1728341909
transform -1 0 50 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3167_
timestamp 1728341909
transform 1 0 2010 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3168_
timestamp 1728341909
transform 1 0 1950 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3169_
timestamp 1728341909
transform -1 0 2250 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3170_
timestamp 1728341909
transform 1 0 1990 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3171_
timestamp 1728341909
transform -1 0 2190 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3172_
timestamp 1728341909
transform 1 0 1850 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__3173_
timestamp 1728341909
transform -1 0 1730 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3174_
timestamp 1728341909
transform -1 0 1750 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3175_
timestamp 1728341909
transform -1 0 2990 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3176_
timestamp 1728341909
transform -1 0 2790 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3177_
timestamp 1728341909
transform 1 0 2230 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3178_
timestamp 1728341909
transform 1 0 2570 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3179_
timestamp 1728341909
transform 1 0 2230 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3180_
timestamp 1728341909
transform 1 0 3170 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3181_
timestamp 1728341909
transform -1 0 2890 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3182_
timestamp 1728341909
transform -1 0 2970 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3183_
timestamp 1728341909
transform 1 0 2730 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3184_
timestamp 1728341909
transform -1 0 2490 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3185_
timestamp 1728341909
transform -1 0 2490 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3186_
timestamp 1728341909
transform 1 0 1970 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3187_
timestamp 1728341909
transform -1 0 310 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3188_
timestamp 1728341909
transform -1 0 50 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3189_
timestamp 1728341909
transform 1 0 990 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3190_
timestamp 1728341909
transform -1 0 790 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3191_
timestamp 1728341909
transform -1 0 1050 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3192_
timestamp 1728341909
transform 1 0 1670 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3193_
timestamp 1728341909
transform 1 0 1410 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3194_
timestamp 1728341909
transform 1 0 3210 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3195_
timestamp 1728341909
transform 1 0 3170 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__3196_
timestamp 1728341909
transform 1 0 1910 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3197_
timestamp 1728341909
transform -1 0 2490 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__3198_
timestamp 1728341909
transform -1 0 2070 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3199_
timestamp 1728341909
transform -1 0 2330 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3200_
timestamp 1728341909
transform 1 0 770 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3201_
timestamp 1728341909
transform -1 0 1010 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3202_
timestamp 1728341909
transform 1 0 1010 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3203_
timestamp 1728341909
transform -1 0 1270 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3204_
timestamp 1728341909
transform -1 0 530 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3205_
timestamp 1728341909
transform -1 0 530 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3206_
timestamp 1728341909
transform 1 0 1030 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__3207_
timestamp 1728341909
transform -1 0 290 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3208_
timestamp 1728341909
transform -1 0 50 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3209_
timestamp 1728341909
transform 1 0 270 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3210_
timestamp 1728341909
transform -1 0 50 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3211_
timestamp 1728341909
transform -1 0 1530 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3212_
timestamp 1728341909
transform -1 0 1270 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3213_
timestamp 1728341909
transform 1 0 1550 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3214_
timestamp 1728341909
transform 1 0 1290 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3215_
timestamp 1728341909
transform -1 0 1250 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3216_
timestamp 1728341909
transform 1 0 990 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3217_
timestamp 1728341909
transform -1 0 290 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3218_
timestamp 1728341909
transform -1 0 50 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3219_
timestamp 1728341909
transform -1 0 1570 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3220_
timestamp 1728341909
transform 1 0 1790 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3221_
timestamp 1728341909
transform -1 0 310 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3222_
timestamp 1728341909
transform -1 0 50 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3223_
timestamp 1728341909
transform -1 0 790 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__3224_
timestamp 1728341909
transform 1 0 510 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3225_
timestamp 1728341909
transform -1 0 290 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3226_
timestamp 1728341909
transform -1 0 50 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3227_
timestamp 1728341909
transform -1 0 310 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__3228_
timestamp 1728341909
transform -1 0 50 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__3229_
timestamp 1728341909
transform -1 0 1970 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__3230_
timestamp 1728341909
transform 1 0 1690 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__3231_
timestamp 1728341909
transform 1 0 1490 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__3232_
timestamp 1728341909
transform -1 0 1750 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__3233_
timestamp 1728341909
transform 1 0 1050 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3234_
timestamp 1728341909
transform -1 0 1330 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3235_
timestamp 1728341909
transform 1 0 1010 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3236_
timestamp 1728341909
transform 1 0 1270 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3237_
timestamp 1728341909
transform 1 0 2190 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__3238_
timestamp 1728341909
transform 1 0 2430 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__3239_
timestamp 1728341909
transform -1 0 530 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3240_
timestamp 1728341909
transform -1 0 770 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3241_
timestamp 1728341909
transform 1 0 9670 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__3242_
timestamp 1728341909
transform -1 0 9010 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__3243_
timestamp 1728341909
transform 1 0 9430 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__3244_
timestamp 1728341909
transform 1 0 8730 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__3245_
timestamp 1728341909
transform 1 0 9030 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3246_
timestamp 1728341909
transform -1 0 9550 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3247_
timestamp 1728341909
transform 1 0 10450 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3248_
timestamp 1728341909
transform 1 0 10710 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3249_
timestamp 1728341909
transform -1 0 9450 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__3250_
timestamp 1728341909
transform 1 0 9370 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3251_
timestamp 1728341909
transform 1 0 9210 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__3252_
timestamp 1728341909
transform -1 0 9230 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__3253_
timestamp 1728341909
transform -1 0 7850 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3254_
timestamp 1728341909
transform -1 0 8110 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3255_
timestamp 1728341909
transform -1 0 9290 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3256_
timestamp 1728341909
transform 1 0 8230 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3257_
timestamp 1728341909
transform 1 0 7990 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3258_
timestamp 1728341909
transform 1 0 8530 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3259_
timestamp 1728341909
transform 1 0 9470 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3260_
timestamp 1728341909
transform -1 0 10830 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__3261_
timestamp 1728341909
transform -1 0 10370 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3262_
timestamp 1728341909
transform 1 0 9950 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3263_
timestamp 1728341909
transform 1 0 9630 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__3264_
timestamp 1728341909
transform 1 0 8970 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__3265_
timestamp 1728341909
transform -1 0 9710 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3266_
timestamp 1728341909
transform 1 0 9730 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3267_
timestamp 1728341909
transform -1 0 9630 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3268_
timestamp 1728341909
transform -1 0 9970 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3269_
timestamp 1728341909
transform -1 0 10470 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3270_
timestamp 1728341909
transform 1 0 10190 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3271_
timestamp 1728341909
transform -1 0 10010 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__3272_
timestamp 1728341909
transform 1 0 10230 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__3273_
timestamp 1728341909
transform -1 0 10130 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__3274_
timestamp 1728341909
transform -1 0 10230 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3275_
timestamp 1728341909
transform 1 0 9550 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__3276_
timestamp 1728341909
transform -1 0 9170 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3277_
timestamp 1728341909
transform -1 0 10630 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3278_
timestamp 1728341909
transform 1 0 10090 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3279_
timestamp 1728341909
transform -1 0 9870 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3280_
timestamp 1728341909
transform 1 0 9210 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__3281_
timestamp 1728341909
transform 1 0 8970 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__3282_
timestamp 1728341909
transform -1 0 6850 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__3283_
timestamp 1728341909
transform -1 0 6790 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3284_
timestamp 1728341909
transform 1 0 6550 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__3285_
timestamp 1728341909
transform 1 0 6990 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3286_
timestamp 1728341909
transform -1 0 7250 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3287_
timestamp 1728341909
transform -1 0 6610 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3288_
timestamp 1728341909
transform -1 0 6830 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3289_
timestamp 1728341909
transform -1 0 6790 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__3290_
timestamp 1728341909
transform 1 0 6510 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__3291_
timestamp 1728341909
transform 1 0 7010 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3292_
timestamp 1728341909
transform -1 0 7270 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3293_
timestamp 1728341909
transform 1 0 7110 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3294_
timestamp 1728341909
transform 1 0 6850 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3295_
timestamp 1728341909
transform 1 0 6050 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3296_
timestamp 1728341909
transform 1 0 5790 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3297_
timestamp 1728341909
transform 1 0 5410 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3298_
timestamp 1728341909
transform 1 0 5150 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3299_
timestamp 1728341909
transform 1 0 5590 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3300_
timestamp 1728341909
transform 1 0 5350 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3301_
timestamp 1728341909
transform 1 0 6850 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__3302_
timestamp 1728341909
transform 1 0 2930 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3303_
timestamp 1728341909
transform -1 0 2990 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3304_
timestamp 1728341909
transform 1 0 1930 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3305_
timestamp 1728341909
transform -1 0 2190 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3306_
timestamp 1728341909
transform 1 0 3850 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3307_
timestamp 1728341909
transform -1 0 4790 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3308_
timestamp 1728341909
transform -1 0 50 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__3309_
timestamp 1728341909
transform -1 0 50 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3310_
timestamp 1728341909
transform -1 0 730 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__3311_
timestamp 1728341909
transform -1 0 770 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3312_
timestamp 1728341909
transform -1 0 270 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__3313_
timestamp 1728341909
transform -1 0 310 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3314_
timestamp 1728341909
transform -1 0 50 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3315_
timestamp 1728341909
transform -1 0 50 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3316_
timestamp 1728341909
transform -1 0 550 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3317_
timestamp 1728341909
transform -1 0 770 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3449_
timestamp 1728341909
transform -1 0 3790 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3450_
timestamp 1728341909
transform 1 0 2950 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3451_
timestamp 1728341909
transform 1 0 3070 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3452_
timestamp 1728341909
transform -1 0 3330 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3453_
timestamp 1728341909
transform 1 0 3190 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3454_
timestamp 1728341909
transform -1 0 3550 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3455_
timestamp 1728341909
transform 1 0 9930 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3456_
timestamp 1728341909
transform 1 0 9490 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3457_
timestamp 1728341909
transform -1 0 9770 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3458_
timestamp 1728341909
transform -1 0 9930 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3459_
timestamp 1728341909
transform 1 0 10370 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3460_
timestamp 1728341909
transform -1 0 10670 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3461_
timestamp 1728341909
transform -1 0 10430 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3462_
timestamp 1728341909
transform -1 0 9990 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3463_
timestamp 1728341909
transform 1 0 10390 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3464_
timestamp 1728341909
transform -1 0 10190 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3465_
timestamp 1728341909
transform 1 0 10150 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1__3466_
timestamp 1728341909
transform -1 0 10170 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3467_
timestamp 1728341909
transform 1 0 8230 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__3468_
timestamp 1728341909
transform 1 0 9070 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__3469_
timestamp 1728341909
transform 1 0 8530 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3470_
timestamp 1728341909
transform -1 0 8470 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3471_
timestamp 1728341909
transform 1 0 8610 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__3472_
timestamp 1728341909
transform 1 0 8850 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__3473_
timestamp 1728341909
transform -1 0 8670 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3474_
timestamp 1728341909
transform -1 0 8790 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3475_
timestamp 1728341909
transform -1 0 8910 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3476_
timestamp 1728341909
transform 1 0 9710 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3477_
timestamp 1728341909
transform 1 0 9150 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3478_
timestamp 1728341909
transform -1 0 9030 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3479_
timestamp 1728341909
transform 1 0 10510 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__3480_
timestamp 1728341909
transform -1 0 10070 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__3481_
timestamp 1728341909
transform -1 0 9930 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3482_
timestamp 1728341909
transform -1 0 9730 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__3483_
timestamp 1728341909
transform 1 0 10870 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3484_
timestamp 1728341909
transform 1 0 10850 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3485_
timestamp 1728341909
transform 1 0 11130 0 1 6490
box -12 -8 32 252
use FILL  FILL_1__3486_
timestamp 1728341909
transform 1 0 11090 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3487_
timestamp 1728341909
transform 1 0 10850 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3488_
timestamp 1728341909
transform 1 0 9490 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3489_
timestamp 1728341909
transform 1 0 9390 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3490_
timestamp 1728341909
transform -1 0 9650 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3491_
timestamp 1728341909
transform -1 0 9670 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3492_
timestamp 1728341909
transform 1 0 9870 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3493_
timestamp 1728341909
transform 1 0 10130 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3494_
timestamp 1728341909
transform 1 0 10270 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__3495_
timestamp 1728341909
transform -1 0 8770 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3496_
timestamp 1728341909
transform 1 0 9390 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3497_
timestamp 1728341909
transform 1 0 9910 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3498_
timestamp 1728341909
transform 1 0 9770 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__3499_
timestamp 1728341909
transform 1 0 9190 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3500_
timestamp 1728341909
transform -1 0 9450 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3501_
timestamp 1728341909
transform -1 0 9690 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3502_
timestamp 1728341909
transform 1 0 9530 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__3503_
timestamp 1728341909
transform 1 0 10010 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__3504_
timestamp 1728341909
transform -1 0 9970 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3505_
timestamp 1728341909
transform 1 0 10210 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3506_
timestamp 1728341909
transform 1 0 10730 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__3507_
timestamp 1728341909
transform -1 0 9350 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__3508_
timestamp 1728341909
transform -1 0 8470 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3509_
timestamp 1728341909
transform 1 0 8390 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__3510_
timestamp 1728341909
transform 1 0 9170 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3511_
timestamp 1728341909
transform -1 0 8930 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3512_
timestamp 1728341909
transform 1 0 8670 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3513_
timestamp 1728341909
transform -1 0 8950 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3514_
timestamp 1728341909
transform -1 0 8710 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3515_
timestamp 1728341909
transform -1 0 9110 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__3516_
timestamp 1728341909
transform 1 0 10950 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__3517_
timestamp 1728341909
transform -1 0 10270 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__3518_
timestamp 1728341909
transform 1 0 10350 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3519_
timestamp 1728341909
transform 1 0 10830 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3520_
timestamp 1728341909
transform -1 0 11130 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3521_
timestamp 1728341909
transform 1 0 7450 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3522_
timestamp 1728341909
transform -1 0 7970 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3523_
timestamp 1728341909
transform 1 0 8710 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3524_
timestamp 1728341909
transform 1 0 8490 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3525_
timestamp 1728341909
transform 1 0 8910 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3526_
timestamp 1728341909
transform -1 0 9190 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3527_
timestamp 1728341909
transform -1 0 8250 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3528_
timestamp 1728341909
transform -1 0 9890 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3529_
timestamp 1728341909
transform 1 0 9990 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__3530_
timestamp 1728341909
transform 1 0 10090 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3531_
timestamp 1728341909
transform -1 0 10130 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3532_
timestamp 1728341909
transform 1 0 10270 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__3533_
timestamp 1728341909
transform -1 0 8190 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3534_
timestamp 1728341909
transform -1 0 8450 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3535_
timestamp 1728341909
transform -1 0 8010 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3536_
timestamp 1728341909
transform -1 0 8230 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3537_
timestamp 1728341909
transform 1 0 8330 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__3538_
timestamp 1728341909
transform -1 0 8610 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__3539_
timestamp 1728341909
transform -1 0 9510 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__3540_
timestamp 1728341909
transform 1 0 9730 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__3541_
timestamp 1728341909
transform -1 0 9810 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__3542_
timestamp 1728341909
transform -1 0 7470 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3543_
timestamp 1728341909
transform -1 0 7730 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3544_
timestamp 1728341909
transform 1 0 7950 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3545_
timestamp 1728341909
transform 1 0 8810 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__3546_
timestamp 1728341909
transform -1 0 8250 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3547_
timestamp 1728341909
transform 1 0 8670 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3548_
timestamp 1728341909
transform -1 0 8930 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3549_
timestamp 1728341909
transform -1 0 8890 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__3550_
timestamp 1728341909
transform 1 0 8870 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3551_
timestamp 1728341909
transform 1 0 9150 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3552_
timestamp 1728341909
transform 1 0 9290 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__3553_
timestamp 1728341909
transform 1 0 9030 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__3554_
timestamp 1728341909
transform 1 0 8950 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__3555_
timestamp 1728341909
transform -1 0 8530 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3556_
timestamp 1728341909
transform 1 0 8430 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3557_
timestamp 1728341909
transform -1 0 8090 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__3558_
timestamp 1728341909
transform -1 0 7730 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3559_
timestamp 1728341909
transform 1 0 7690 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3560_
timestamp 1728341909
transform 1 0 8210 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3561_
timestamp 1728341909
transform -1 0 7950 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3562_
timestamp 1728341909
transform -1 0 8950 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3563_
timestamp 1728341909
transform -1 0 8930 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__3564_
timestamp 1728341909
transform 1 0 10030 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__3565_
timestamp 1728341909
transform -1 0 9950 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__3566_
timestamp 1728341909
transform 1 0 9870 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3567_
timestamp 1728341909
transform 1 0 9950 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__3568_
timestamp 1728341909
transform 1 0 10170 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__3569_
timestamp 1728341909
transform 1 0 10170 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__3570_
timestamp 1728341909
transform 1 0 10630 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__3571_
timestamp 1728341909
transform -1 0 10610 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3572_
timestamp 1728341909
transform -1 0 11110 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3573_
timestamp 1728341909
transform 1 0 10990 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__3574_
timestamp 1728341909
transform 1 0 10730 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__3575_
timestamp 1728341909
transform 1 0 11130 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__3576_
timestamp 1728341909
transform 1 0 9910 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__3577_
timestamp 1728341909
transform -1 0 11150 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__3578_
timestamp 1728341909
transform 1 0 10750 0 -1 9850
box -12 -8 32 252
use FILL  FILL_1__3579_
timestamp 1728341909
transform -1 0 10450 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__3580_
timestamp 1728341909
transform -1 0 9150 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3581_
timestamp 1728341909
transform -1 0 8850 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__3582_
timestamp 1728341909
transform 1 0 8690 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__3583_
timestamp 1728341909
transform -1 0 9010 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__3584_
timestamp 1728341909
transform 1 0 8750 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__3585_
timestamp 1728341909
transform -1 0 9490 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__3586_
timestamp 1728341909
transform 1 0 9070 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__3587_
timestamp 1728341909
transform -1 0 9210 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__3588_
timestamp 1728341909
transform 1 0 9230 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__3589_
timestamp 1728341909
transform 1 0 9950 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__3590_
timestamp 1728341909
transform -1 0 10210 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__3591_
timestamp 1728341909
transform 1 0 9690 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__3592_
timestamp 1728341909
transform 1 0 9710 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__3593_
timestamp 1728341909
transform -1 0 9490 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__3594_
timestamp 1728341909
transform 1 0 10330 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3595_
timestamp 1728341909
transform 1 0 10890 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__3596_
timestamp 1728341909
transform -1 0 10850 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3597_
timestamp 1728341909
transform 1 0 10490 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__3598_
timestamp 1728341909
transform 1 0 11130 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__3599_
timestamp 1728341909
transform 1 0 11090 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3600_
timestamp 1728341909
transform 1 0 10970 0 -1 9370
box -12 -8 32 252
use FILL  FILL_1__3601_
timestamp 1728341909
transform 1 0 10150 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3602_
timestamp 1728341909
transform 1 0 10390 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3603_
timestamp 1728341909
transform 1 0 10450 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3604_
timestamp 1728341909
transform 1 0 10670 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3605_
timestamp 1728341909
transform 1 0 11150 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3606_
timestamp 1728341909
transform 1 0 10630 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3607_
timestamp 1728341909
transform -1 0 9930 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3608_
timestamp 1728341909
transform -1 0 10170 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3609_
timestamp 1728341909
transform 1 0 10670 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3610_
timestamp 1728341909
transform 1 0 9490 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3611_
timestamp 1728341909
transform 1 0 9290 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__3612_
timestamp 1728341909
transform 1 0 9550 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__3613_
timestamp 1728341909
transform 1 0 9410 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3614_
timestamp 1728341909
transform -1 0 9810 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__3615_
timestamp 1728341909
transform -1 0 9690 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3616_
timestamp 1728341909
transform -1 0 8990 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3617_
timestamp 1728341909
transform -1 0 9250 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3618_
timestamp 1728341909
transform 1 0 9730 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3619_
timestamp 1728341909
transform 1 0 10890 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3620_
timestamp 1728341909
transform -1 0 10630 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3621_
timestamp 1728341909
transform -1 0 10410 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3622_
timestamp 1728341909
transform 1 0 10650 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3623_
timestamp 1728341909
transform 1 0 9950 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3624_
timestamp 1728341909
transform 1 0 10670 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3625_
timestamp 1728341909
transform 1 0 10770 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__3626_
timestamp 1728341909
transform -1 0 10670 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3627_
timestamp 1728341909
transform -1 0 9650 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3628_
timestamp 1728341909
transform -1 0 10390 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3629_
timestamp 1728341909
transform 1 0 10610 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3630_
timestamp 1728341909
transform 1 0 10410 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3631_
timestamp 1728341909
transform -1 0 10570 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__3632_
timestamp 1728341909
transform -1 0 10910 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__3633_
timestamp 1728341909
transform 1 0 10870 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__3634_
timestamp 1728341909
transform -1 0 10690 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__3635_
timestamp 1728341909
transform -1 0 10410 0 1 10810
box -12 -8 32 252
use FILL  FILL_1__3636_
timestamp 1728341909
transform -1 0 10510 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__3637_
timestamp 1728341909
transform -1 0 10670 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__3638_
timestamp 1728341909
transform -1 0 10590 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3639_
timestamp 1728341909
transform -1 0 10430 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__3640_
timestamp 1728341909
transform -1 0 10890 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3641_
timestamp 1728341909
transform -1 0 10630 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3642_
timestamp 1728341909
transform -1 0 10950 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3643_
timestamp 1728341909
transform 1 0 10870 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3644_
timestamp 1728341909
transform -1 0 10430 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3645_
timestamp 1728341909
transform -1 0 10170 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3646_
timestamp 1728341909
transform -1 0 10930 0 -1 8890
box -12 -8 32 252
use FILL  FILL_1__3647_
timestamp 1728341909
transform 1 0 11030 0 1 250
box -12 -8 32 252
use FILL  FILL_1__3648_
timestamp 1728341909
transform 1 0 11110 0 1 8410
box -12 -8 32 252
use FILL  FILL_1__3649_
timestamp 1728341909
transform 1 0 10190 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3650_
timestamp 1728341909
transform 1 0 10310 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__3651_
timestamp 1728341909
transform 1 0 10410 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3652_
timestamp 1728341909
transform -1 0 10370 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3653_
timestamp 1728341909
transform 1 0 10590 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3654_
timestamp 1728341909
transform 1 0 8390 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3655_
timestamp 1728341909
transform -1 0 8650 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3656_
timestamp 1728341909
transform 1 0 8230 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__3657_
timestamp 1728341909
transform -1 0 8610 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__3658_
timestamp 1728341909
transform -1 0 8510 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__3659_
timestamp 1728341909
transform -1 0 8250 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1__3660_
timestamp 1728341909
transform -1 0 8370 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__3661_
timestamp 1728341909
transform -1 0 9230 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__3662_
timestamp 1728341909
transform -1 0 9470 0 1 10330
box -12 -8 32 252
use FILL  FILL_1__3663_
timestamp 1728341909
transform 1 0 9390 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3664_
timestamp 1728341909
transform -1 0 9630 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3665_
timestamp 1728341909
transform 1 0 8230 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3666_
timestamp 1728341909
transform -1 0 8470 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3667_
timestamp 1728341909
transform -1 0 9190 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3668_
timestamp 1728341909
transform -1 0 10410 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3669_
timestamp 1728341909
transform -1 0 10150 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3670_
timestamp 1728341909
transform -1 0 9910 0 1 9370
box -12 -8 32 252
use FILL  FILL_1__3671_
timestamp 1728341909
transform 1 0 8270 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3672_
timestamp 1728341909
transform 1 0 8510 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3673_
timestamp 1728341909
transform -1 0 9430 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3674_
timestamp 1728341909
transform -1 0 9890 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3675_
timestamp 1728341909
transform 1 0 10110 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3676_
timestamp 1728341909
transform -1 0 10150 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3677_
timestamp 1728341909
transform 1 0 9390 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3678_
timestamp 1728341909
transform -1 0 9230 0 -1 6970
box -12 -8 32 252
use FILL  FILL_1__3691_
timestamp 1728341909
transform 1 0 7710 0 1 250
box -12 -8 32 252
use FILL  FILL_1__3692_
timestamp 1728341909
transform -1 0 7970 0 1 250
box -12 -8 32 252
use FILL  FILL_1__3693_
timestamp 1728341909
transform -1 0 1950 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3694_
timestamp 1728341909
transform -1 0 50 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3695_
timestamp 1728341909
transform 1 0 550 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3696_
timestamp 1728341909
transform -1 0 50 0 1 9850
box -12 -8 32 252
use FILL  FILL_1__3697_
timestamp 1728341909
transform -1 0 50 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__3698_
timestamp 1728341909
transform -1 0 290 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1__3699_
timestamp 1728341909
transform 1 0 6110 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__3700_
timestamp 1728341909
transform -1 0 6270 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__3701_
timestamp 1728341909
transform -1 0 6250 0 1 250
box -12 -8 32 252
use FILL  FILL_1__3702_
timestamp 1728341909
transform -1 0 5230 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__3703_
timestamp 1728341909
transform -1 0 3470 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__3704_
timestamp 1728341909
transform -1 0 3250 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__3705_
timestamp 1728341909
transform -1 0 50 0 1 8890
box -12 -8 32 252
use FILL  FILL_1__3706_
timestamp 1728341909
transform -1 0 1290 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1__3707_
timestamp 1728341909
transform 1 0 11110 0 1 6970
box -12 -8 32 252
use FILL  FILL_1__3708_
timestamp 1728341909
transform 1 0 11110 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1__3709_
timestamp 1728341909
transform 1 0 11130 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3710_
timestamp 1728341909
transform 1 0 10890 0 1 7450
box -12 -8 32 252
use FILL  FILL_1__3711_
timestamp 1728341909
transform 1 0 11110 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1__3712_
timestamp 1728341909
transform 1 0 10890 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3713_
timestamp 1728341909
transform 1 0 11010 0 1 7930
box -12 -8 32 252
use FILL  FILL_1__3714_
timestamp 1728341909
transform 1 0 11130 0 -1 8410
box -12 -8 32 252
use FILL  FILL_1__3715_
timestamp 1728341909
transform 1 0 11110 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert0
timestamp 1728341909
transform 1 0 7750 0 1 10810
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert1
timestamp 1728341909
transform 1 0 8970 0 1 1690
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert2
timestamp 1728341909
transform 1 0 9170 0 1 6970
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert3
timestamp 1728341909
transform 1 0 5650 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert4
timestamp 1728341909
transform 1 0 6750 0 1 1690
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert5
timestamp 1728341909
transform -1 0 4010 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert6
timestamp 1728341909
transform 1 0 7170 0 1 10330
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert7
timestamp 1728341909
transform -1 0 4090 0 1 4090
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert8
timestamp 1728341909
transform -1 0 7530 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert9
timestamp 1728341909
transform 1 0 4450 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert10
timestamp 1728341909
transform -1 0 570 0 1 4090
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert11
timestamp 1728341909
transform -1 0 4770 0 1 2650
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert12
timestamp 1728341909
transform 1 0 730 0 1 5530
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert13
timestamp 1728341909
transform -1 0 5870 0 1 7450
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert14
timestamp 1728341909
transform 1 0 4510 0 1 2650
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert15
timestamp 1728341909
transform 1 0 5590 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert16
timestamp 1728341909
transform 1 0 2670 0 1 8410
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert17
timestamp 1728341909
transform 1 0 4170 0 1 6490
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert18
timestamp 1728341909
transform -1 0 50 0 1 2650
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert19
timestamp 1728341909
transform -1 0 310 0 1 8410
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert20
timestamp 1728341909
transform 1 0 510 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert21
timestamp 1728341909
transform -1 0 7050 0 1 4570
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert22
timestamp 1728341909
transform -1 0 10430 0 1 4090
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert23
timestamp 1728341909
transform -1 0 8770 0 1 4090
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert24
timestamp 1728341909
transform 1 0 8490 0 1 3130
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert25
timestamp 1728341909
transform -1 0 7050 0 1 3130
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert37
timestamp 1728341909
transform -1 0 970 0 1 5530
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert38
timestamp 1728341909
transform 1 0 1250 0 1 4570
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert39
timestamp 1728341909
transform -1 0 1010 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert40
timestamp 1728341909
transform -1 0 2710 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert41
timestamp 1728341909
transform 1 0 9510 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert42
timestamp 1728341909
transform 1 0 8830 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert43
timestamp 1728341909
transform -1 0 8750 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert44
timestamp 1728341909
transform -1 0 8970 0 1 4570
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert45
timestamp 1728341909
transform 1 0 3830 0 1 4090
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert46
timestamp 1728341909
transform 1 0 5190 0 1 4090
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert47
timestamp 1728341909
transform 1 0 4290 0 1 2650
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert48
timestamp 1728341909
transform 1 0 5410 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert49
timestamp 1728341909
transform -1 0 2210 0 1 2650
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert50
timestamp 1728341909
transform 1 0 8290 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert51
timestamp 1728341909
transform -1 0 10390 0 1 4570
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert52
timestamp 1728341909
transform -1 0 9430 0 1 4570
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert53
timestamp 1728341909
transform -1 0 9510 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert54
timestamp 1728341909
transform -1 0 8350 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert55
timestamp 1728341909
transform -1 0 310 0 1 730
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert56
timestamp 1728341909
transform 1 0 4990 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert57
timestamp 1728341909
transform 1 0 4590 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert58
timestamp 1728341909
transform 1 0 1910 0 1 1690
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert59
timestamp 1728341909
transform 1 0 4350 0 1 730
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert60
timestamp 1728341909
transform -1 0 8730 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert61
timestamp 1728341909
transform 1 0 10130 0 -1 7450
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert62
timestamp 1728341909
transform 1 0 9170 0 -1 10330
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert63
timestamp 1728341909
transform 1 0 9250 0 1 7450
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert64
timestamp 1728341909
transform 1 0 8590 0 1 1210
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert65
timestamp 1728341909
transform -1 0 4990 0 1 4090
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert66
timestamp 1728341909
transform 1 0 5730 0 1 2650
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert67
timestamp 1728341909
transform 1 0 6570 0 1 5050
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert68
timestamp 1728341909
transform 1 0 7570 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert69
timestamp 1728341909
transform -1 0 6050 0 1 1690
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert70
timestamp 1728341909
transform 1 0 8730 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert71
timestamp 1728341909
transform 1 0 2430 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert72
timestamp 1728341909
transform 1 0 3870 0 1 1210
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert73
timestamp 1728341909
transform 1 0 2670 0 1 2650
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert74
timestamp 1728341909
transform -1 0 3670 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert75
timestamp 1728341909
transform -1 0 750 0 1 2170
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert76
timestamp 1728341909
transform 1 0 8730 0 1 4570
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert77
timestamp 1728341909
transform -1 0 8470 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert78
timestamp 1728341909
transform 1 0 8930 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert79
timestamp 1728341909
transform -1 0 9190 0 1 4570
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert80
timestamp 1728341909
transform 1 0 4170 0 -1 6490
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert81
timestamp 1728341909
transform 1 0 3310 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert82
timestamp 1728341909
transform 1 0 2170 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert83
timestamp 1728341909
transform -1 0 2650 0 -1 7930
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert26
timestamp 1728341909
transform -1 0 1390 0 1 3130
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert27
timestamp 1728341909
transform 1 0 3630 0 1 3130
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert28
timestamp 1728341909
transform 1 0 30 0 1 3130
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert29
timestamp 1728341909
transform 1 0 510 0 1 7930
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert30
timestamp 1728341909
transform 1 0 8190 0 1 5530
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert31
timestamp 1728341909
transform -1 0 7550 0 -1 10810
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert32
timestamp 1728341909
transform -1 0 3170 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert33
timestamp 1728341909
transform -1 0 7910 0 1 10330
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert34
timestamp 1728341909
transform -1 0 50 0 -1 11290
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert35
timestamp 1728341909
transform -1 0 5470 0 1 5050
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert36
timestamp 1728341909
transform -1 0 2850 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__1744_
timestamp 1728341909
transform -1 0 4450 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__1745_
timestamp 1728341909
transform 1 0 4230 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__1746_
timestamp 1728341909
transform -1 0 4210 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__1747_
timestamp 1728341909
transform -1 0 5670 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__1748_
timestamp 1728341909
transform 1 0 6590 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__1749_
timestamp 1728341909
transform 1 0 6350 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__1750_
timestamp 1728341909
transform 1 0 5190 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__1751_
timestamp 1728341909
transform 1 0 6830 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__1752_
timestamp 1728341909
transform 1 0 5410 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__1753_
timestamp 1728341909
transform 1 0 7550 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__1754_
timestamp 1728341909
transform -1 0 7090 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__1755_
timestamp 1728341909
transform -1 0 7310 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__1756_
timestamp 1728341909
transform -1 0 6390 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__1757_
timestamp 1728341909
transform 1 0 7050 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__1758_
timestamp 1728341909
transform 1 0 6810 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__1759_
timestamp 1728341909
transform -1 0 3070 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__1760_
timestamp 1728341909
transform 1 0 2370 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__1761_
timestamp 1728341909
transform 1 0 7290 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__1762_
timestamp 1728341909
transform 1 0 2570 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__1763_
timestamp 1728341909
transform -1 0 8210 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__1764_
timestamp 1728341909
transform -1 0 8030 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__1765_
timestamp 1728341909
transform -1 0 8030 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__1766_
timestamp 1728341909
transform -1 0 7830 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__1767_
timestamp 1728341909
transform -1 0 7830 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__1768_
timestamp 1728341909
transform -1 0 5710 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__1769_
timestamp 1728341909
transform 1 0 3150 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__1770_
timestamp 1728341909
transform 1 0 10810 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__1771_
timestamp 1728341909
transform 1 0 11050 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__1772_
timestamp 1728341909
transform 1 0 10790 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__1773_
timestamp 1728341909
transform 1 0 10330 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__1774_
timestamp 1728341909
transform 1 0 10690 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1775_
timestamp 1728341909
transform -1 0 9510 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__1776_
timestamp 1728341909
transform 1 0 9550 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__1777_
timestamp 1728341909
transform -1 0 8730 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__1778_
timestamp 1728341909
transform -1 0 10930 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__1779_
timestamp 1728341909
transform 1 0 10150 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__1780_
timestamp 1728341909
transform 1 0 10910 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__1781_
timestamp 1728341909
transform -1 0 10930 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__1782_
timestamp 1728341909
transform -1 0 11170 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1783_
timestamp 1728341909
transform -1 0 9970 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1784_
timestamp 1728341909
transform 1 0 10550 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__1785_
timestamp 1728341909
transform 1 0 10890 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__1786_
timestamp 1728341909
transform -1 0 10230 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__1787_
timestamp 1728341909
transform 1 0 9230 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__1788_
timestamp 1728341909
transform 1 0 10510 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__1789_
timestamp 1728341909
transform -1 0 9370 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1790_
timestamp 1728341909
transform -1 0 10730 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1791_
timestamp 1728341909
transform 1 0 10950 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1792_
timestamp 1728341909
transform 1 0 5650 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1793_
timestamp 1728341909
transform 1 0 5370 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1794_
timestamp 1728341909
transform -1 0 4950 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1795_
timestamp 1728341909
transform 1 0 3730 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1796_
timestamp 1728341909
transform 1 0 4190 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1797_
timestamp 1728341909
transform -1 0 4710 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1798_
timestamp 1728341909
transform -1 0 11030 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__1799_
timestamp 1728341909
transform -1 0 10930 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__1800_
timestamp 1728341909
transform -1 0 10450 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__1801_
timestamp 1728341909
transform -1 0 10110 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__1802_
timestamp 1728341909
transform 1 0 9990 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__1803_
timestamp 1728341909
transform 1 0 10230 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1804_
timestamp 1728341909
transform 1 0 10230 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__1805_
timestamp 1728341909
transform -1 0 10030 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__1806_
timestamp 1728341909
transform 1 0 9970 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1807_
timestamp 1728341909
transform -1 0 10090 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1808_
timestamp 1728341909
transform -1 0 10390 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__1809_
timestamp 1728341909
transform -1 0 11050 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1810_
timestamp 1728341909
transform -1 0 6230 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1811_
timestamp 1728341909
transform -1 0 11130 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__1812_
timestamp 1728341909
transform -1 0 10210 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__1813_
timestamp 1728341909
transform -1 0 7690 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__1814_
timestamp 1728341909
transform -1 0 7530 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1815_
timestamp 1728341909
transform -1 0 10950 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1816_
timestamp 1728341909
transform -1 0 7590 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__1817_
timestamp 1728341909
transform 1 0 6710 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__1818_
timestamp 1728341909
transform 1 0 6650 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1819_
timestamp 1728341909
transform 1 0 6150 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1820_
timestamp 1728341909
transform 1 0 10350 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__1821_
timestamp 1728341909
transform -1 0 6710 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1822_
timestamp 1728341909
transform 1 0 11130 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__1823_
timestamp 1728341909
transform -1 0 9990 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__1824_
timestamp 1728341909
transform 1 0 7290 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__1825_
timestamp 1728341909
transform 1 0 6510 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1826_
timestamp 1728341909
transform 1 0 10930 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1827_
timestamp 1728341909
transform -1 0 7370 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1828_
timestamp 1728341909
transform 1 0 11130 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__1829_
timestamp 1728341909
transform -1 0 7390 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__1830_
timestamp 1728341909
transform 1 0 7530 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__1831_
timestamp 1728341909
transform 1 0 10670 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__1832_
timestamp 1728341909
transform 1 0 10650 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__1833_
timestamp 1728341909
transform 1 0 7210 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1834_
timestamp 1728341909
transform -1 0 7010 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1835_
timestamp 1728341909
transform -1 0 6450 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1836_
timestamp 1728341909
transform -1 0 6010 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1837_
timestamp 1728341909
transform -1 0 5530 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1838_
timestamp 1728341909
transform 1 0 5250 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1839_
timestamp 1728341909
transform 1 0 5830 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1840_
timestamp 1728341909
transform -1 0 8030 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__1841_
timestamp 1728341909
transform -1 0 4970 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__1842_
timestamp 1728341909
transform -1 0 6830 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__1843_
timestamp 1728341909
transform 1 0 7150 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__1844_
timestamp 1728341909
transform -1 0 10230 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__1845_
timestamp 1728341909
transform 1 0 11130 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__1846_
timestamp 1728341909
transform 1 0 11150 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1847_
timestamp 1728341909
transform -1 0 8070 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__1848_
timestamp 1728341909
transform 1 0 10670 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__1849_
timestamp 1728341909
transform -1 0 10590 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__1850_
timestamp 1728341909
transform -1 0 8530 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__1851_
timestamp 1728341909
transform -1 0 11150 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__1852_
timestamp 1728341909
transform 1 0 9710 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__1853_
timestamp 1728341909
transform 1 0 9230 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__1854_
timestamp 1728341909
transform 1 0 9030 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__1855_
timestamp 1728341909
transform 1 0 8790 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__1856_
timestamp 1728341909
transform 1 0 9310 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__1857_
timestamp 1728341909
transform 1 0 9090 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__1858_
timestamp 1728341909
transform 1 0 7270 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__1859_
timestamp 1728341909
transform -1 0 10690 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__1860_
timestamp 1728341909
transform 1 0 7070 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__1861_
timestamp 1728341909
transform 1 0 7310 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__1862_
timestamp 1728341909
transform -1 0 9810 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__1863_
timestamp 1728341909
transform 1 0 8550 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__1864_
timestamp 1728341909
transform 1 0 9850 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__1865_
timestamp 1728341909
transform 1 0 7710 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__1866_
timestamp 1728341909
transform -1 0 8890 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1867_
timestamp 1728341909
transform 1 0 9270 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__1868_
timestamp 1728341909
transform 1 0 10830 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__1869_
timestamp 1728341909
transform 1 0 9290 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__1870_
timestamp 1728341909
transform -1 0 9070 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__1871_
timestamp 1728341909
transform 1 0 8510 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__1872_
timestamp 1728341909
transform 1 0 7790 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__1873_
timestamp 1728341909
transform 1 0 6350 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1874_
timestamp 1728341909
transform -1 0 6810 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1875_
timestamp 1728341909
transform -1 0 6570 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1876_
timestamp 1728341909
transform 1 0 6630 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__1877_
timestamp 1728341909
transform -1 0 8050 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__1878_
timestamp 1728341909
transform -1 0 8310 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__1879_
timestamp 1728341909
transform -1 0 8050 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__1880_
timestamp 1728341909
transform -1 0 6990 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__1881_
timestamp 1728341909
transform -1 0 6310 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__1882_
timestamp 1728341909
transform 1 0 3470 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__1883_
timestamp 1728341909
transform -1 0 7010 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__1884_
timestamp 1728341909
transform -1 0 6530 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__1885_
timestamp 1728341909
transform 1 0 5810 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__1886_
timestamp 1728341909
transform -1 0 6210 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__1887_
timestamp 1728341909
transform 1 0 6830 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__1888_
timestamp 1728341909
transform 1 0 3590 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__1889_
timestamp 1728341909
transform -1 0 5950 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__1890_
timestamp 1728341909
transform 1 0 6410 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__1891_
timestamp 1728341909
transform -1 0 6050 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__1892_
timestamp 1728341909
transform 1 0 5610 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__1893_
timestamp 1728341909
transform 1 0 1010 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__1894_
timestamp 1728341909
transform 1 0 5950 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__1895_
timestamp 1728341909
transform 1 0 6830 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__1896_
timestamp 1728341909
transform 1 0 5150 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__1897_
timestamp 1728341909
transform 1 0 5990 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__1898_
timestamp 1728341909
transform 1 0 6410 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__1899_
timestamp 1728341909
transform 1 0 6510 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__1900_
timestamp 1728341909
transform 1 0 530 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__1901_
timestamp 1728341909
transform 1 0 7970 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__1902_
timestamp 1728341909
transform 1 0 8510 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__1903_
timestamp 1728341909
transform 1 0 7870 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__1904_
timestamp 1728341909
transform -1 0 10030 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1905_
timestamp 1728341909
transform 1 0 7530 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__1906_
timestamp 1728341909
transform 1 0 7510 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__1907_
timestamp 1728341909
transform 1 0 8650 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1908_
timestamp 1728341909
transform -1 0 7710 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1909_
timestamp 1728341909
transform 1 0 1810 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1910_
timestamp 1728341909
transform -1 0 9770 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__1911_
timestamp 1728341909
transform 1 0 9490 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1912_
timestamp 1728341909
transform 1 0 6110 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1913_
timestamp 1728341909
transform 1 0 10630 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__1914_
timestamp 1728341909
transform 1 0 10690 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1915_
timestamp 1728341909
transform -1 0 10250 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1916_
timestamp 1728341909
transform -1 0 5870 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1917_
timestamp 1728341909
transform 1 0 4010 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1918_
timestamp 1728341909
transform -1 0 790 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__1919_
timestamp 1728341909
transform -1 0 70 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__1920_
timestamp 1728341909
transform 1 0 1010 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__1921_
timestamp 1728341909
transform -1 0 1190 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1922_
timestamp 1728341909
transform -1 0 930 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1923_
timestamp 1728341909
transform 1 0 530 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__1924_
timestamp 1728341909
transform -1 0 4470 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1925_
timestamp 1728341909
transform -1 0 310 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__1926_
timestamp 1728341909
transform 1 0 770 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__1927_
timestamp 1728341909
transform -1 0 2070 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1928_
timestamp 1728341909
transform -1 0 1590 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1929_
timestamp 1728341909
transform 1 0 270 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__1930_
timestamp 1728341909
transform 1 0 650 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1931_
timestamp 1728341909
transform 1 0 530 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__1932_
timestamp 1728341909
transform -1 0 550 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1933_
timestamp 1728341909
transform 1 0 530 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__1934_
timestamp 1728341909
transform -1 0 550 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1935_
timestamp 1728341909
transform -1 0 1530 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1936_
timestamp 1728341909
transform 1 0 790 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1937_
timestamp 1728341909
transform -1 0 550 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__1938_
timestamp 1728341909
transform -1 0 70 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__1939_
timestamp 1728341909
transform 1 0 290 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__1940_
timestamp 1728341909
transform 1 0 810 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1941_
timestamp 1728341909
transform 1 0 530 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__1942_
timestamp 1728341909
transform 1 0 530 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__1943_
timestamp 1728341909
transform 1 0 8090 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__1944_
timestamp 1728341909
transform -1 0 7630 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1945_
timestamp 1728341909
transform -1 0 7410 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1946_
timestamp 1728341909
transform 1 0 8430 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1947_
timestamp 1728341909
transform -1 0 7610 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1948_
timestamp 1728341909
transform -1 0 6950 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1949_
timestamp 1728341909
transform -1 0 7190 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1950_
timestamp 1728341909
transform 1 0 8290 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__1951_
timestamp 1728341909
transform 1 0 8290 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__1952_
timestamp 1728341909
transform 1 0 9810 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1953_
timestamp 1728341909
transform -1 0 8370 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__1954_
timestamp 1728341909
transform 1 0 8210 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1955_
timestamp 1728341909
transform 1 0 6410 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__1956_
timestamp 1728341909
transform -1 0 7970 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1957_
timestamp 1728341909
transform 1 0 8050 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__1958_
timestamp 1728341909
transform 1 0 10410 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__1959_
timestamp 1728341909
transform 1 0 7770 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__1960_
timestamp 1728341909
transform 1 0 7850 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__1961_
timestamp 1728341909
transform 1 0 10670 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__1962_
timestamp 1728341909
transform 1 0 10470 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__1963_
timestamp 1728341909
transform 1 0 9810 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1964_
timestamp 1728341909
transform -1 0 7350 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__1965_
timestamp 1728341909
transform -1 0 7630 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__1966_
timestamp 1728341909
transform -1 0 3490 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__1967_
timestamp 1728341909
transform -1 0 6950 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__1968_
timestamp 1728341909
transform 1 0 7490 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__1969_
timestamp 1728341909
transform -1 0 7750 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__1970_
timestamp 1728341909
transform 1 0 1490 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__1971_
timestamp 1728341909
transform -1 0 790 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1972_
timestamp 1728341909
transform 1 0 1310 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1973_
timestamp 1728341909
transform 1 0 1570 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__1974_
timestamp 1728341909
transform 1 0 8330 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__1975_
timestamp 1728341909
transform 1 0 2950 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__1976_
timestamp 1728341909
transform -1 0 7110 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__1977_
timestamp 1728341909
transform -1 0 2810 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__1978_
timestamp 1728341909
transform -1 0 3790 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__1979_
timestamp 1728341909
transform -1 0 6490 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__1980_
timestamp 1728341909
transform 1 0 7750 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__1981_
timestamp 1728341909
transform 1 0 8270 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__1982_
timestamp 1728341909
transform -1 0 3010 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__1983_
timestamp 1728341909
transform 1 0 1690 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__1984_
timestamp 1728341909
transform 1 0 1770 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__1985_
timestamp 1728341909
transform 1 0 2430 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__1986_
timestamp 1728341909
transform -1 0 7110 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__1987_
timestamp 1728341909
transform 1 0 5050 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__1988_
timestamp 1728341909
transform -1 0 4950 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__1989_
timestamp 1728341909
transform 1 0 6710 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__1990_
timestamp 1728341909
transform -1 0 7230 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__1991_
timestamp 1728341909
transform -1 0 2030 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__1992_
timestamp 1728341909
transform -1 0 1530 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__1993_
timestamp 1728341909
transform -1 0 1810 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__1994_
timestamp 1728341909
transform 1 0 2050 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__1995_
timestamp 1728341909
transform 1 0 8010 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__1996_
timestamp 1728341909
transform -1 0 2230 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__1997_
timestamp 1728341909
transform -1 0 3950 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__1998_
timestamp 1728341909
transform -1 0 6470 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__1999_
timestamp 1728341909
transform -1 0 8190 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2000_
timestamp 1728341909
transform 1 0 1790 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2001_
timestamp 1728341909
transform 1 0 1270 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2002_
timestamp 1728341909
transform 1 0 1510 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2003_
timestamp 1728341909
transform 1 0 1530 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2004_
timestamp 1728341909
transform 1 0 7810 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2005_
timestamp 1728341909
transform 1 0 1970 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2006_
timestamp 1728341909
transform -1 0 6230 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2007_
timestamp 1728341909
transform 1 0 7510 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2008_
timestamp 1728341909
transform -1 0 8030 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2009_
timestamp 1728341909
transform 1 0 770 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2010_
timestamp 1728341909
transform -1 0 830 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2011_
timestamp 1728341909
transform 1 0 530 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2012_
timestamp 1728341909
transform 1 0 790 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2013_
timestamp 1728341909
transform 1 0 5430 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2014_
timestamp 1728341909
transform 1 0 1730 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2015_
timestamp 1728341909
transform -1 0 3930 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2016_
timestamp 1728341909
transform 1 0 6730 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2017_
timestamp 1728341909
transform -1 0 7270 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2018_
timestamp 1728341909
transform -1 0 1510 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2019_
timestamp 1728341909
transform -1 0 1570 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2020_
timestamp 1728341909
transform 1 0 1750 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2021_
timestamp 1728341909
transform 1 0 1710 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2022_
timestamp 1728341909
transform 1 0 4490 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2023_
timestamp 1728341909
transform 1 0 530 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2024_
timestamp 1728341909
transform 1 0 1430 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2025_
timestamp 1728341909
transform 1 0 2490 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2026_
timestamp 1728341909
transform -1 0 4690 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2027_
timestamp 1728341909
transform 1 0 7190 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2028_
timestamp 1728341909
transform -1 0 7470 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2029_
timestamp 1728341909
transform -1 0 70 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2030_
timestamp 1728341909
transform -1 0 550 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2031_
timestamp 1728341909
transform -1 0 310 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2032_
timestamp 1728341909
transform 1 0 530 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2033_
timestamp 1728341909
transform 1 0 7610 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2034_
timestamp 1728341909
transform 1 0 1210 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2035_
timestamp 1728341909
transform 1 0 2090 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2036_
timestamp 1728341909
transform 1 0 2890 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2037_
timestamp 1728341909
transform -1 0 4090 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2038_
timestamp 1728341909
transform 1 0 7530 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2039_
timestamp 1728341909
transform -1 0 7810 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2040_
timestamp 1728341909
transform -1 0 2930 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2041_
timestamp 1728341909
transform -1 0 550 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2042_
timestamp 1728341909
transform 1 0 1710 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__2043_
timestamp 1728341909
transform -1 0 3810 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__2044_
timestamp 1728341909
transform 1 0 5350 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2045_
timestamp 1728341909
transform -1 0 4050 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2046_
timestamp 1728341909
transform 1 0 2850 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__2047_
timestamp 1728341909
transform 1 0 2610 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__2048_
timestamp 1728341909
transform -1 0 3550 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__2049_
timestamp 1728341909
transform -1 0 2950 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__2050_
timestamp 1728341909
transform -1 0 2430 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__2051_
timestamp 1728341909
transform -1 0 2410 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2052_
timestamp 1728341909
transform -1 0 830 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2053_
timestamp 1728341909
transform -1 0 3390 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__2054_
timestamp 1728341909
transform 1 0 3110 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__2055_
timestamp 1728341909
transform -1 0 2750 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__2056_
timestamp 1728341909
transform 1 0 4370 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2057_
timestamp 1728341909
transform -1 0 3930 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2058_
timestamp 1728341909
transform 1 0 4590 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2059_
timestamp 1728341909
transform -1 0 1950 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__2060_
timestamp 1728341909
transform -1 0 3770 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__2061_
timestamp 1728341909
transform 1 0 3510 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__2062_
timestamp 1728341909
transform -1 0 3530 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__2063_
timestamp 1728341909
transform 1 0 2470 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__2064_
timestamp 1728341909
transform -1 0 2570 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2065_
timestamp 1728341909
transform -1 0 2370 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2066_
timestamp 1728341909
transform 1 0 2430 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2067_
timestamp 1728341909
transform -1 0 2750 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__2068_
timestamp 1728341909
transform -1 0 2990 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__2069_
timestamp 1728341909
transform 1 0 2530 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__2070_
timestamp 1728341909
transform -1 0 1070 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2071_
timestamp 1728341909
transform -1 0 2790 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__2072_
timestamp 1728341909
transform -1 0 2530 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__2073_
timestamp 1728341909
transform -1 0 1270 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2074_
timestamp 1728341909
transform 1 0 3210 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__2075_
timestamp 1728341909
transform -1 0 2690 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__2076_
timestamp 1728341909
transform 1 0 2390 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__2077_
timestamp 1728341909
transform -1 0 3250 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__2078_
timestamp 1728341909
transform 1 0 2770 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__2079_
timestamp 1728341909
transform -1 0 3890 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2080_
timestamp 1728341909
transform 1 0 4110 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2081_
timestamp 1728341909
transform -1 0 3670 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2082_
timestamp 1728341909
transform 1 0 5750 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2083_
timestamp 1728341909
transform -1 0 6490 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2084_
timestamp 1728341909
transform 1 0 9910 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2085_
timestamp 1728341909
transform -1 0 10430 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2086_
timestamp 1728341909
transform 1 0 10450 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2087_
timestamp 1728341909
transform 1 0 10990 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__2088_
timestamp 1728341909
transform 1 0 10190 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2089_
timestamp 1728341909
transform -1 0 9490 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2090_
timestamp 1728341909
transform 1 0 10670 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__2091_
timestamp 1728341909
transform 1 0 11170 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__2092_
timestamp 1728341909
transform -1 0 10130 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2093_
timestamp 1728341909
transform 1 0 10190 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__2094_
timestamp 1728341909
transform -1 0 10690 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__2095_
timestamp 1728341909
transform 1 0 10750 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__2096_
timestamp 1728341909
transform -1 0 11150 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__2097_
timestamp 1728341909
transform -1 0 11090 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2098_
timestamp 1728341909
transform 1 0 10170 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2099_
timestamp 1728341909
transform 1 0 10650 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2100_
timestamp 1728341909
transform 1 0 10870 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2101_
timestamp 1728341909
transform 1 0 11110 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2102_
timestamp 1728341909
transform 1 0 3990 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__2103_
timestamp 1728341909
transform 1 0 4230 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__2104_
timestamp 1728341909
transform 1 0 3850 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2105_
timestamp 1728341909
transform -1 0 1750 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2106_
timestamp 1728341909
transform -1 0 2130 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2107_
timestamp 1728341909
transform -1 0 2650 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2108_
timestamp 1728341909
transform 1 0 1450 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2109_
timestamp 1728341909
transform -1 0 2870 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2110_
timestamp 1728341909
transform 1 0 3090 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2111_
timestamp 1728341909
transform 1 0 5290 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2112_
timestamp 1728341909
transform 1 0 11170 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__2113_
timestamp 1728341909
transform -1 0 9750 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__2114_
timestamp 1728341909
transform 1 0 9750 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2115_
timestamp 1728341909
transform -1 0 11070 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2116_
timestamp 1728341909
transform -1 0 11010 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__2117_
timestamp 1728341909
transform -1 0 10610 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__2118_
timestamp 1728341909
transform 1 0 9010 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__2119_
timestamp 1728341909
transform -1 0 11090 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__2120_
timestamp 1728341909
transform 1 0 11030 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2121_
timestamp 1728341909
transform 1 0 11130 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2122_
timestamp 1728341909
transform 1 0 10830 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2123_
timestamp 1728341909
transform 1 0 10890 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2124_
timestamp 1728341909
transform 1 0 9350 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2125_
timestamp 1728341909
transform 1 0 9470 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2126_
timestamp 1728341909
transform -1 0 9910 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2127_
timestamp 1728341909
transform 1 0 9730 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2128_
timestamp 1728341909
transform 1 0 9690 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2129_
timestamp 1728341909
transform -1 0 8910 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2130_
timestamp 1728341909
transform 1 0 9590 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2131_
timestamp 1728341909
transform 1 0 9690 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2132_
timestamp 1728341909
transform 1 0 10150 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2133_
timestamp 1728341909
transform 1 0 10310 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2134_
timestamp 1728341909
transform -1 0 10090 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2135_
timestamp 1728341909
transform 1 0 10590 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2136_
timestamp 1728341909
transform -1 0 10550 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2137_
timestamp 1728341909
transform 1 0 10790 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2138_
timestamp 1728341909
transform -1 0 10890 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2139_
timestamp 1728341909
transform -1 0 10830 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2140_
timestamp 1728341909
transform -1 0 8310 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2141_
timestamp 1728341909
transform 1 0 8550 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2142_
timestamp 1728341909
transform 1 0 1870 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2143_
timestamp 1728341909
transform -1 0 2910 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2144_
timestamp 1728341909
transform -1 0 6010 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2145_
timestamp 1728341909
transform -1 0 6210 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2146_
timestamp 1728341909
transform 1 0 5510 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2147_
timestamp 1728341909
transform -1 0 6750 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2148_
timestamp 1728341909
transform 1 0 9650 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2149_
timestamp 1728341909
transform 1 0 8730 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2150_
timestamp 1728341909
transform -1 0 8490 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2151_
timestamp 1728341909
transform 1 0 8150 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2152_
timestamp 1728341909
transform -1 0 8990 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2153_
timestamp 1728341909
transform -1 0 9090 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2154_
timestamp 1728341909
transform 1 0 8830 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__2155_
timestamp 1728341909
transform 1 0 7990 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__2156_
timestamp 1728341909
transform -1 0 8270 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__2157_
timestamp 1728341909
transform -1 0 8390 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2158_
timestamp 1728341909
transform 1 0 10310 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__2159_
timestamp 1728341909
transform 1 0 6010 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2160_
timestamp 1728341909
transform -1 0 6370 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2161_
timestamp 1728341909
transform 1 0 6570 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2162_
timestamp 1728341909
transform -1 0 7910 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2163_
timestamp 1728341909
transform -1 0 8330 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__2164_
timestamp 1728341909
transform 1 0 7090 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2165_
timestamp 1728341909
transform -1 0 7070 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2166_
timestamp 1728341909
transform -1 0 8130 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2167_
timestamp 1728341909
transform -1 0 7830 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2168_
timestamp 1728341909
transform -1 0 8090 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2169_
timestamp 1728341909
transform 1 0 8130 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2170_
timestamp 1728341909
transform -1 0 8350 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2171_
timestamp 1728341909
transform 1 0 8550 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2172_
timestamp 1728341909
transform -1 0 10410 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2173_
timestamp 1728341909
transform 1 0 10150 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2174_
timestamp 1728341909
transform 1 0 4370 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2175_
timestamp 1728341909
transform -1 0 3930 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2176_
timestamp 1728341909
transform -1 0 5390 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2177_
timestamp 1728341909
transform -1 0 6050 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2178_
timestamp 1728341909
transform -1 0 6310 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2179_
timestamp 1728341909
transform 1 0 6350 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2180_
timestamp 1728341909
transform 1 0 7150 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2181_
timestamp 1728341909
transform 1 0 7290 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__2182_
timestamp 1728341909
transform -1 0 7150 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__2183_
timestamp 1728341909
transform 1 0 6130 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2184_
timestamp 1728341909
transform 1 0 6450 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2185_
timestamp 1728341909
transform -1 0 6590 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2186_
timestamp 1728341909
transform -1 0 9030 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2187_
timestamp 1728341909
transform -1 0 9430 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2188_
timestamp 1728341909
transform 1 0 9030 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2189_
timestamp 1728341909
transform -1 0 8810 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2190_
timestamp 1728341909
transform 1 0 8490 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2191_
timestamp 1728341909
transform 1 0 8730 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2192_
timestamp 1728341909
transform 1 0 7290 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2193_
timestamp 1728341909
transform 1 0 7510 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2194_
timestamp 1728341909
transform -1 0 8630 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__2195_
timestamp 1728341909
transform -1 0 8550 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__2196_
timestamp 1728341909
transform 1 0 8590 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2197_
timestamp 1728341909
transform 1 0 8630 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2198_
timestamp 1728341909
transform -1 0 7230 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2199_
timestamp 1728341909
transform -1 0 7490 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2200_
timestamp 1728341909
transform 1 0 9010 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__2201_
timestamp 1728341909
transform 1 0 8870 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2202_
timestamp 1728341909
transform -1 0 8670 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2203_
timestamp 1728341909
transform 1 0 8390 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2204_
timestamp 1728341909
transform -1 0 8390 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2205_
timestamp 1728341909
transform 1 0 8130 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2206_
timestamp 1728341909
transform -1 0 8010 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2207_
timestamp 1728341909
transform 1 0 8510 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2208_
timestamp 1728341909
transform -1 0 8270 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2209_
timestamp 1728341909
transform -1 0 7790 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2210_
timestamp 1728341909
transform 1 0 2730 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2211_
timestamp 1728341909
transform -1 0 7190 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2212_
timestamp 1728341909
transform -1 0 7450 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2213_
timestamp 1728341909
transform -1 0 7970 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2214_
timestamp 1728341909
transform 1 0 8530 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2215_
timestamp 1728341909
transform 1 0 9230 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2216_
timestamp 1728341909
transform 1 0 9210 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2217_
timestamp 1728341909
transform -1 0 9470 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2218_
timestamp 1728341909
transform 1 0 3910 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2219_
timestamp 1728341909
transform -1 0 2230 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__2220_
timestamp 1728341909
transform -1 0 3650 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2221_
timestamp 1728341909
transform 1 0 4090 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2222_
timestamp 1728341909
transform 1 0 4310 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2223_
timestamp 1728341909
transform 1 0 4130 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2224_
timestamp 1728341909
transform -1 0 2810 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2225_
timestamp 1728341909
transform -1 0 5870 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2226_
timestamp 1728341909
transform 1 0 5990 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2227_
timestamp 1728341909
transform -1 0 6970 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2228_
timestamp 1728341909
transform 1 0 6710 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2229_
timestamp 1728341909
transform 1 0 7770 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__2230_
timestamp 1728341909
transform -1 0 6170 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__2231_
timestamp 1728341909
transform -1 0 6410 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__2232_
timestamp 1728341909
transform 1 0 6830 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2233_
timestamp 1728341909
transform 1 0 7410 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2234_
timestamp 1728341909
transform 1 0 7310 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2235_
timestamp 1728341909
transform 1 0 9390 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2236_
timestamp 1728341909
transform 1 0 10450 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2237_
timestamp 1728341909
transform 1 0 9930 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2238_
timestamp 1728341909
transform -1 0 9850 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2239_
timestamp 1728341909
transform -1 0 5810 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2240_
timestamp 1728341909
transform 1 0 2670 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2241_
timestamp 1728341909
transform -1 0 4350 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2242_
timestamp 1728341909
transform -1 0 4570 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2243_
timestamp 1728341909
transform 1 0 3350 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2244_
timestamp 1728341909
transform 1 0 5110 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2245_
timestamp 1728341909
transform 1 0 7250 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2246_
timestamp 1728341909
transform 1 0 7270 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2247_
timestamp 1728341909
transform -1 0 3230 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2248_
timestamp 1728341909
transform 1 0 3410 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2249_
timestamp 1728341909
transform 1 0 5390 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2250_
timestamp 1728341909
transform 1 0 6650 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2251_
timestamp 1728341909
transform 1 0 7170 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2252_
timestamp 1728341909
transform -1 0 9610 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__2253_
timestamp 1728341909
transform 1 0 9330 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2254_
timestamp 1728341909
transform 1 0 5610 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2255_
timestamp 1728341909
transform -1 0 6950 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2256_
timestamp 1728341909
transform 1 0 7110 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2257_
timestamp 1728341909
transform -1 0 3050 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2258_
timestamp 1728341909
transform -1 0 3010 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__2259_
timestamp 1728341909
transform 1 0 3430 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2260_
timestamp 1728341909
transform 1 0 4610 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2261_
timestamp 1728341909
transform -1 0 5610 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2262_
timestamp 1728341909
transform 1 0 4790 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2263_
timestamp 1728341909
transform 1 0 4850 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2264_
timestamp 1728341909
transform -1 0 6150 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2265_
timestamp 1728341909
transform 1 0 3450 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__2266_
timestamp 1728341909
transform 1 0 7490 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__2267_
timestamp 1728341909
transform -1 0 5390 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__2268_
timestamp 1728341909
transform -1 0 5630 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__2269_
timestamp 1728341909
transform 1 0 5390 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__2270_
timestamp 1728341909
transform -1 0 6230 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__2271_
timestamp 1728341909
transform 1 0 5950 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__2272_
timestamp 1728341909
transform 1 0 5550 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__2273_
timestamp 1728341909
transform 1 0 5370 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__2274_
timestamp 1728341909
transform 1 0 5130 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__2275_
timestamp 1728341909
transform 1 0 5610 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__2276_
timestamp 1728341909
transform -1 0 6250 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2277_
timestamp 1728341909
transform 1 0 7750 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__2278_
timestamp 1728341909
transform -1 0 7690 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2279_
timestamp 1728341909
transform 1 0 6450 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2280_
timestamp 1728341909
transform -1 0 6470 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2281_
timestamp 1728341909
transform -1 0 6230 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2282_
timestamp 1728341909
transform 1 0 6510 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2283_
timestamp 1728341909
transform 1 0 7210 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2284_
timestamp 1728341909
transform 1 0 9170 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2285_
timestamp 1728341909
transform 1 0 9610 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2286_
timestamp 1728341909
transform -1 0 2510 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__2287_
timestamp 1728341909
transform -1 0 1770 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2288_
timestamp 1728341909
transform -1 0 2210 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2289_
timestamp 1728341909
transform 1 0 2170 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2290_
timestamp 1728341909
transform -1 0 1730 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2291_
timestamp 1728341909
transform 1 0 1950 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2292_
timestamp 1728341909
transform 1 0 4070 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2293_
timestamp 1728341909
transform 1 0 4810 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2294_
timestamp 1728341909
transform 1 0 6030 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2295_
timestamp 1728341909
transform -1 0 2210 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2296_
timestamp 1728341909
transform 1 0 3650 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2297_
timestamp 1728341909
transform 1 0 2190 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2298_
timestamp 1728341909
transform 1 0 1950 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2299_
timestamp 1728341909
transform 1 0 3410 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2300_
timestamp 1728341909
transform 1 0 3150 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2301_
timestamp 1728341909
transform -1 0 3610 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2302_
timestamp 1728341909
transform 1 0 5090 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2303_
timestamp 1728341909
transform -1 0 5070 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2304_
timestamp 1728341909
transform 1 0 5310 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2305_
timestamp 1728341909
transform -1 0 1510 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2306_
timestamp 1728341909
transform 1 0 2410 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2307_
timestamp 1728341909
transform -1 0 5570 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2308_
timestamp 1728341909
transform -1 0 5570 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2309_
timestamp 1728341909
transform 1 0 4570 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2310_
timestamp 1728341909
transform 1 0 4330 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2311_
timestamp 1728341909
transform -1 0 3730 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2312_
timestamp 1728341909
transform -1 0 3970 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2313_
timestamp 1728341909
transform 1 0 5250 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2314_
timestamp 1728341909
transform 1 0 4430 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2315_
timestamp 1728341909
transform 1 0 5390 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2316_
timestamp 1728341909
transform -1 0 9830 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2317_
timestamp 1728341909
transform 1 0 11130 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2318_
timestamp 1728341909
transform -1 0 10830 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__2319_
timestamp 1728341909
transform -1 0 10450 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__2320_
timestamp 1728341909
transform 1 0 10610 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2321_
timestamp 1728341909
transform 1 0 10550 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__2322_
timestamp 1728341909
transform 1 0 10450 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__2323_
timestamp 1728341909
transform 1 0 6710 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2324_
timestamp 1728341909
transform 1 0 6910 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2325_
timestamp 1728341909
transform 1 0 9270 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2326_
timestamp 1728341909
transform -1 0 8810 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2327_
timestamp 1728341909
transform -1 0 9270 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2328_
timestamp 1728341909
transform -1 0 9510 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2329_
timestamp 1728341909
transform 1 0 9230 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2330_
timestamp 1728341909
transform -1 0 8990 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2331_
timestamp 1728341909
transform -1 0 9150 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2332_
timestamp 1728341909
transform 1 0 9130 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2333_
timestamp 1728341909
transform 1 0 9390 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2334_
timestamp 1728341909
transform -1 0 9590 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2335_
timestamp 1728341909
transform 1 0 5630 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2336_
timestamp 1728341909
transform 1 0 6150 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2337_
timestamp 1728341909
transform -1 0 5930 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2338_
timestamp 1728341909
transform -1 0 5870 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2339_
timestamp 1728341909
transform 1 0 10350 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2340_
timestamp 1728341909
transform -1 0 9230 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2341_
timestamp 1728341909
transform 1 0 9230 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2342_
timestamp 1728341909
transform 1 0 10090 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2343_
timestamp 1728341909
transform -1 0 9590 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2344_
timestamp 1728341909
transform 1 0 9690 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2345_
timestamp 1728341909
transform -1 0 6870 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2346_
timestamp 1728341909
transform 1 0 6730 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2347_
timestamp 1728341909
transform -1 0 7070 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2348_
timestamp 1728341909
transform 1 0 8070 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2349_
timestamp 1728341909
transform -1 0 7770 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2350_
timestamp 1728341909
transform 1 0 7490 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2351_
timestamp 1728341909
transform -1 0 5190 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2352_
timestamp 1728341909
transform 1 0 5790 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2353_
timestamp 1728341909
transform -1 0 4210 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2354_
timestamp 1728341909
transform 1 0 4690 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2355_
timestamp 1728341909
transform -1 0 4950 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2356_
timestamp 1728341909
transform 1 0 5890 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2357_
timestamp 1728341909
transform -1 0 5650 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2358_
timestamp 1728341909
transform 1 0 6930 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2359_
timestamp 1728341909
transform 1 0 6290 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2360_
timestamp 1728341909
transform 1 0 6530 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2361_
timestamp 1728341909
transform 1 0 7830 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__2362_
timestamp 1728341909
transform 1 0 7350 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2363_
timestamp 1728341909
transform -1 0 7450 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2364_
timestamp 1728341909
transform 1 0 8070 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__2365_
timestamp 1728341909
transform -1 0 7950 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2366_
timestamp 1728341909
transform 1 0 7710 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2367_
timestamp 1728341909
transform 1 0 7990 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2368_
timestamp 1728341909
transform 1 0 8210 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2369_
timestamp 1728341909
transform -1 0 9930 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2370_
timestamp 1728341909
transform 1 0 5350 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2371_
timestamp 1728341909
transform -1 0 8750 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2372_
timestamp 1728341909
transform -1 0 8490 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2373_
timestamp 1728341909
transform -1 0 8070 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2374_
timestamp 1728341909
transform 1 0 8070 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2375_
timestamp 1728341909
transform 1 0 6470 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2376_
timestamp 1728341909
transform 1 0 8430 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2377_
timestamp 1728341909
transform -1 0 8690 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2378_
timestamp 1728341909
transform -1 0 8990 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2379_
timestamp 1728341909
transform -1 0 6850 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2380_
timestamp 1728341909
transform -1 0 6990 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2381_
timestamp 1728341909
transform -1 0 6850 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2382_
timestamp 1728341909
transform -1 0 7930 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2383_
timestamp 1728341909
transform 1 0 7650 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2384_
timestamp 1728341909
transform 1 0 7750 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2385_
timestamp 1728341909
transform -1 0 7490 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2386_
timestamp 1728341909
transform -1 0 6610 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2387_
timestamp 1728341909
transform -1 0 6370 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2388_
timestamp 1728341909
transform -1 0 8930 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2389_
timestamp 1728341909
transform -1 0 8310 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2390_
timestamp 1728341909
transform -1 0 8250 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2391_
timestamp 1728341909
transform -1 0 9490 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2392_
timestamp 1728341909
transform 1 0 8250 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2393_
timestamp 1728341909
transform 1 0 8210 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2394_
timestamp 1728341909
transform 1 0 8850 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2395_
timestamp 1728341909
transform 1 0 8810 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2396_
timestamp 1728341909
transform 1 0 9090 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2397_
timestamp 1728341909
transform -1 0 9350 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2398_
timestamp 1728341909
transform 1 0 8730 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2399_
timestamp 1728341909
transform -1 0 7610 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2400_
timestamp 1728341909
transform 1 0 7350 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2401_
timestamp 1728341909
transform 1 0 8470 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2402_
timestamp 1728341909
transform -1 0 6410 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2403_
timestamp 1728341909
transform -1 0 6610 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2404_
timestamp 1728341909
transform -1 0 7570 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2405_
timestamp 1728341909
transform -1 0 7350 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2406_
timestamp 1728341909
transform 1 0 7070 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2407_
timestamp 1728341909
transform -1 0 6610 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2408_
timestamp 1728341909
transform -1 0 5910 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2409_
timestamp 1728341909
transform 1 0 6990 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2410_
timestamp 1728341909
transform -1 0 7270 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2411_
timestamp 1728341909
transform -1 0 6830 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2412_
timestamp 1728341909
transform -1 0 7490 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2413_
timestamp 1728341909
transform 1 0 7010 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2414_
timestamp 1728341909
transform 1 0 6830 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2415_
timestamp 1728341909
transform -1 0 8030 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2416_
timestamp 1728341909
transform 1 0 7770 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2417_
timestamp 1728341909
transform -1 0 9010 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2418_
timestamp 1728341909
transform -1 0 8790 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2419_
timestamp 1728341909
transform 1 0 7050 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2420_
timestamp 1728341909
transform 1 0 2210 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2421_
timestamp 1728341909
transform -1 0 9670 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2422_
timestamp 1728341909
transform 1 0 8250 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__2423_
timestamp 1728341909
transform 1 0 8970 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2424_
timestamp 1728341909
transform 1 0 8750 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2425_
timestamp 1728341909
transform 1 0 3150 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2426_
timestamp 1728341909
transform 1 0 8730 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2427_
timestamp 1728341909
transform 1 0 8810 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__2428_
timestamp 1728341909
transform 1 0 9210 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2429_
timestamp 1728341909
transform 1 0 9430 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2430_
timestamp 1728341909
transform 1 0 8790 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2431_
timestamp 1728341909
transform -1 0 9250 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2432_
timestamp 1728341909
transform 1 0 9470 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2433_
timestamp 1728341909
transform -1 0 9890 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2434_
timestamp 1728341909
transform -1 0 9970 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2435_
timestamp 1728341909
transform 1 0 4430 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__2436_
timestamp 1728341909
transform 1 0 9190 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2437_
timestamp 1728341909
transform 1 0 10870 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__2438_
timestamp 1728341909
transform -1 0 10930 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__2439_
timestamp 1728341909
transform -1 0 10910 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__2440_
timestamp 1728341909
transform 1 0 9030 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__2441_
timestamp 1728341909
transform -1 0 6170 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__2442_
timestamp 1728341909
transform -1 0 8250 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2443_
timestamp 1728341909
transform 1 0 3810 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2444_
timestamp 1728341909
transform -1 0 4690 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__2445_
timestamp 1728341909
transform -1 0 8590 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__2446_
timestamp 1728341909
transform 1 0 8230 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2447_
timestamp 1728341909
transform 1 0 8070 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2448_
timestamp 1728341909
transform 1 0 8470 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2449_
timestamp 1728341909
transform -1 0 8750 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2450_
timestamp 1728341909
transform -1 0 8950 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2451_
timestamp 1728341909
transform 1 0 3810 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2452_
timestamp 1728341909
transform 1 0 7590 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2453_
timestamp 1728341909
transform -1 0 6610 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2454_
timestamp 1728341909
transform -1 0 6330 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2455_
timestamp 1728341909
transform -1 0 6610 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2456_
timestamp 1728341909
transform -1 0 8730 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2457_
timestamp 1728341909
transform -1 0 8950 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2458_
timestamp 1728341909
transform -1 0 6790 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2459_
timestamp 1728341909
transform -1 0 3570 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2460_
timestamp 1728341909
transform 1 0 7090 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2461_
timestamp 1728341909
transform 1 0 7010 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2462_
timestamp 1728341909
transform -1 0 7290 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2463_
timestamp 1728341909
transform -1 0 7310 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2464_
timestamp 1728341909
transform 1 0 4470 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__2465_
timestamp 1728341909
transform -1 0 7370 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2466_
timestamp 1728341909
transform -1 0 3350 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2467_
timestamp 1728341909
transform 1 0 6170 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2468_
timestamp 1728341909
transform -1 0 6290 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2469_
timestamp 1728341909
transform -1 0 6130 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2470_
timestamp 1728341909
transform -1 0 6390 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2471_
timestamp 1728341909
transform -1 0 8050 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2472_
timestamp 1728341909
transform -1 0 6070 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2473_
timestamp 1728341909
transform -1 0 5410 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2474_
timestamp 1728341909
transform -1 0 5330 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2475_
timestamp 1728341909
transform -1 0 7790 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__2476_
timestamp 1728341909
transform -1 0 2710 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2477_
timestamp 1728341909
transform -1 0 5190 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2478_
timestamp 1728341909
transform 1 0 5270 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2479_
timestamp 1728341909
transform -1 0 8010 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2480_
timestamp 1728341909
transform 1 0 5910 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2481_
timestamp 1728341909
transform 1 0 4170 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2482_
timestamp 1728341909
transform -1 0 2450 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2483_
timestamp 1728341909
transform -1 0 4690 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2484_
timestamp 1728341909
transform -1 0 5730 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2485_
timestamp 1728341909
transform -1 0 6970 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2486_
timestamp 1728341909
transform 1 0 3090 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2487_
timestamp 1728341909
transform -1 0 5670 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2488_
timestamp 1728341909
transform 1 0 6430 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2489_
timestamp 1728341909
transform -1 0 6710 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2490_
timestamp 1728341909
transform 1 0 7690 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2491_
timestamp 1728341909
transform -1 0 7930 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2492_
timestamp 1728341909
transform -1 0 2870 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2493_
timestamp 1728341909
transform -1 0 5510 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2494_
timestamp 1728341909
transform -1 0 6590 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2495_
timestamp 1728341909
transform 1 0 6830 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2496_
timestamp 1728341909
transform 1 0 7550 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2497_
timestamp 1728341909
transform -1 0 7790 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2498_
timestamp 1728341909
transform -1 0 8770 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__2499_
timestamp 1728341909
transform 1 0 9010 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2500_
timestamp 1728341909
transform -1 0 7630 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2501_
timestamp 1728341909
transform -1 0 6750 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__2502_
timestamp 1728341909
transform -1 0 7610 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__2503_
timestamp 1728341909
transform 1 0 11110 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2504_
timestamp 1728341909
transform -1 0 4550 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2505_
timestamp 1728341909
transform -1 0 5690 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2506_
timestamp 1728341909
transform -1 0 6710 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__2507_
timestamp 1728341909
transform 1 0 5850 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2508_
timestamp 1728341909
transform 1 0 5650 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2509_
timestamp 1728341909
transform -1 0 8810 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__2510_
timestamp 1728341909
transform -1 0 8070 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__2511_
timestamp 1728341909
transform -1 0 7390 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__2512_
timestamp 1728341909
transform 1 0 7090 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__2513_
timestamp 1728341909
transform 1 0 6870 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__2514_
timestamp 1728341909
transform 1 0 7030 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__2515_
timestamp 1728341909
transform 1 0 10370 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__2516_
timestamp 1728341909
transform 1 0 8510 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2517_
timestamp 1728341909
transform 1 0 10610 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2518_
timestamp 1728341909
transform -1 0 9710 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__2519_
timestamp 1728341909
transform 1 0 9950 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__2520_
timestamp 1728341909
transform -1 0 10410 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2521_
timestamp 1728341909
transform -1 0 8510 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2522_
timestamp 1728341909
transform 1 0 6070 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2523_
timestamp 1728341909
transform 1 0 5890 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2524_
timestamp 1728341909
transform 1 0 8270 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2525_
timestamp 1728341909
transform 1 0 6770 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2526_
timestamp 1728341909
transform -1 0 7770 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2527_
timestamp 1728341909
transform 1 0 7990 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2528_
timestamp 1728341909
transform -1 0 8050 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2529_
timestamp 1728341909
transform 1 0 7830 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2530_
timestamp 1728341909
transform -1 0 7790 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2531_
timestamp 1728341909
transform -1 0 7810 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2532_
timestamp 1728341909
transform 1 0 7810 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2533_
timestamp 1728341909
transform -1 0 5470 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2534_
timestamp 1728341909
transform -1 0 5890 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2535_
timestamp 1728341909
transform -1 0 7570 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2536_
timestamp 1728341909
transform 1 0 7370 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2537_
timestamp 1728341909
transform 1 0 7290 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2538_
timestamp 1728341909
transform 1 0 8010 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2539_
timestamp 1728341909
transform 1 0 5870 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2540_
timestamp 1728341909
transform 1 0 5590 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2541_
timestamp 1728341909
transform 1 0 6110 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2542_
timestamp 1728341909
transform -1 0 6650 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2543_
timestamp 1728341909
transform -1 0 6610 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2544_
timestamp 1728341909
transform 1 0 6150 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2545_
timestamp 1728341909
transform 1 0 6850 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2546_
timestamp 1728341909
transform 1 0 6110 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2547_
timestamp 1728341909
transform 1 0 6330 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2548_
timestamp 1728341909
transform 1 0 7110 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2549_
timestamp 1728341909
transform 1 0 7370 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2550_
timestamp 1728341909
transform -1 0 7530 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2551_
timestamp 1728341909
transform -1 0 6250 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2552_
timestamp 1728341909
transform -1 0 4810 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2553_
timestamp 1728341909
transform -1 0 5850 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2554_
timestamp 1728341909
transform -1 0 5570 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2555_
timestamp 1728341909
transform 1 0 5630 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2556_
timestamp 1728341909
transform 1 0 5010 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2557_
timestamp 1728341909
transform 1 0 5750 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2558_
timestamp 1728341909
transform -1 0 6390 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2559_
timestamp 1728341909
transform 1 0 6070 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__2560_
timestamp 1728341909
transform 1 0 4330 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2561_
timestamp 1728341909
transform -1 0 5390 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2562_
timestamp 1728341909
transform 1 0 5010 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2563_
timestamp 1728341909
transform -1 0 4910 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2564_
timestamp 1728341909
transform -1 0 4570 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2565_
timestamp 1728341909
transform 1 0 4710 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2566_
timestamp 1728341909
transform -1 0 4930 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2567_
timestamp 1728341909
transform 1 0 5130 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2568_
timestamp 1728341909
transform 1 0 5270 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__2569_
timestamp 1728341909
transform -1 0 4150 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2570_
timestamp 1728341909
transform 1 0 5170 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2571_
timestamp 1728341909
transform 1 0 4290 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2572_
timestamp 1728341909
transform -1 0 4410 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2573_
timestamp 1728341909
transform 1 0 4650 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2574_
timestamp 1728341909
transform 1 0 5370 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2575_
timestamp 1728341909
transform -1 0 4930 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2576_
timestamp 1728341909
transform 1 0 5110 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2577_
timestamp 1728341909
transform 1 0 4850 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2578_
timestamp 1728341909
transform -1 0 4790 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2579_
timestamp 1728341909
transform 1 0 4650 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__2580_
timestamp 1728341909
transform 1 0 4690 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__2581_
timestamp 1728341909
transform -1 0 4130 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2582_
timestamp 1728341909
transform -1 0 3270 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2583_
timestamp 1728341909
transform 1 0 2210 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2584_
timestamp 1728341909
transform 1 0 3170 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2585_
timestamp 1728341909
transform -1 0 6330 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2586_
timestamp 1728341909
transform -1 0 3690 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2587_
timestamp 1728341909
transform -1 0 3430 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2588_
timestamp 1728341909
transform -1 0 2950 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2589_
timestamp 1728341909
transform -1 0 2950 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2590_
timestamp 1728341909
transform 1 0 3570 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__2591_
timestamp 1728341909
transform -1 0 3050 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2592_
timestamp 1728341909
transform 1 0 2550 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2593_
timestamp 1728341909
transform -1 0 2650 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2594_
timestamp 1728341909
transform -1 0 2670 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2595_
timestamp 1728341909
transform -1 0 3750 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__2596_
timestamp 1728341909
transform 1 0 3350 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2597_
timestamp 1728341909
transform 1 0 3290 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2598_
timestamp 1728341909
transform -1 0 3170 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2599_
timestamp 1728341909
transform -1 0 3170 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2600_
timestamp 1728341909
transform 1 0 2890 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2601_
timestamp 1728341909
transform -1 0 2450 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2602_
timestamp 1728341909
transform -1 0 2710 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2603_
timestamp 1728341909
transform -1 0 2310 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2604_
timestamp 1728341909
transform 1 0 2450 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2605_
timestamp 1728341909
transform -1 0 2450 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2606_
timestamp 1728341909
transform 1 0 2170 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2607_
timestamp 1728341909
transform -1 0 1530 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2608_
timestamp 1728341909
transform -1 0 1050 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2609_
timestamp 1728341909
transform 1 0 2010 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2610_
timestamp 1728341909
transform 1 0 1250 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2611_
timestamp 1728341909
transform -1 0 1230 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2612_
timestamp 1728341909
transform -1 0 970 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2613_
timestamp 1728341909
transform -1 0 1950 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2614_
timestamp 1728341909
transform -1 0 570 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2615_
timestamp 1728341909
transform 1 0 1750 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2616_
timestamp 1728341909
transform 1 0 1490 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2617_
timestamp 1728341909
transform -1 0 1490 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2618_
timestamp 1728341909
transform -1 0 1730 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2619_
timestamp 1728341909
transform 1 0 770 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2620_
timestamp 1728341909
transform -1 0 1290 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2621_
timestamp 1728341909
transform 1 0 1030 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2622_
timestamp 1728341909
transform -1 0 1250 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2623_
timestamp 1728341909
transform 1 0 990 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2624_
timestamp 1728341909
transform -1 0 530 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2625_
timestamp 1728341909
transform -1 0 2610 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2626_
timestamp 1728341909
transform 1 0 1630 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2627_
timestamp 1728341909
transform 1 0 1370 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2628_
timestamp 1728341909
transform 1 0 770 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2629_
timestamp 1728341909
transform -1 0 3370 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__2630_
timestamp 1728341909
transform 1 0 4230 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__2631_
timestamp 1728341909
transform -1 0 4890 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__2632_
timestamp 1728341909
transform 1 0 10870 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2633_
timestamp 1728341909
transform 1 0 3870 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2634_
timestamp 1728341909
transform 1 0 8970 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2635_
timestamp 1728341909
transform -1 0 2250 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__2636_
timestamp 1728341909
transform -1 0 9130 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__2637_
timestamp 1728341909
transform 1 0 4330 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2638_
timestamp 1728341909
transform 1 0 4830 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2639_
timestamp 1728341909
transform -1 0 9910 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__2640_
timestamp 1728341909
transform -1 0 9850 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__2641_
timestamp 1728341909
transform 1 0 10150 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2642_
timestamp 1728341909
transform -1 0 9490 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__2643_
timestamp 1728341909
transform 1 0 10890 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2644_
timestamp 1728341909
transform -1 0 9730 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2645_
timestamp 1728341909
transform -1 0 9690 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__2646_
timestamp 1728341909
transform 1 0 10090 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__2647_
timestamp 1728341909
transform -1 0 8570 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2648_
timestamp 1728341909
transform -1 0 4150 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__2649_
timestamp 1728341909
transform -1 0 5790 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2650_
timestamp 1728341909
transform 1 0 9290 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__2651_
timestamp 1728341909
transform -1 0 5670 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2652_
timestamp 1728341909
transform -1 0 7830 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__2653_
timestamp 1728341909
transform -1 0 7730 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__2654_
timestamp 1728341909
transform 1 0 4650 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2655_
timestamp 1728341909
transform -1 0 5430 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2656_
timestamp 1728341909
transform -1 0 6010 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2657_
timestamp 1728341909
transform -1 0 6750 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2658_
timestamp 1728341909
transform 1 0 6250 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2659_
timestamp 1728341909
transform 1 0 6950 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2660_
timestamp 1728341909
transform -1 0 7230 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2661_
timestamp 1728341909
transform -1 0 4450 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2662_
timestamp 1728341909
transform 1 0 4410 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2663_
timestamp 1728341909
transform 1 0 6330 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2664_
timestamp 1728341909
transform -1 0 6590 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2665_
timestamp 1728341909
transform 1 0 7090 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2666_
timestamp 1728341909
transform 1 0 6830 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2667_
timestamp 1728341909
transform 1 0 7570 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2668_
timestamp 1728341909
transform 1 0 7310 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2669_
timestamp 1728341909
transform 1 0 7970 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2670_
timestamp 1728341909
transform -1 0 4190 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2671_
timestamp 1728341909
transform -1 0 5310 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__2672_
timestamp 1728341909
transform 1 0 5210 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2673_
timestamp 1728341909
transform 1 0 7170 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2674_
timestamp 1728341909
transform -1 0 7390 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2675_
timestamp 1728341909
transform 1 0 7630 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2676_
timestamp 1728341909
transform -1 0 7570 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2677_
timestamp 1728341909
transform 1 0 7750 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2678_
timestamp 1728341909
transform 1 0 7710 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2679_
timestamp 1728341909
transform 1 0 4150 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2680_
timestamp 1728341909
transform -1 0 4410 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2681_
timestamp 1728341909
transform 1 0 6110 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2682_
timestamp 1728341909
transform 1 0 6730 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2683_
timestamp 1728341909
transform 1 0 4070 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2684_
timestamp 1728341909
transform -1 0 5730 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2685_
timestamp 1728341909
transform 1 0 5450 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2686_
timestamp 1728341909
transform -1 0 6870 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2687_
timestamp 1728341909
transform 1 0 7330 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2688_
timestamp 1728341909
transform -1 0 7470 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2689_
timestamp 1728341909
transform 1 0 6490 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2690_
timestamp 1728341909
transform 1 0 6570 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2691_
timestamp 1728341909
transform 1 0 7070 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2692_
timestamp 1728341909
transform -1 0 7210 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2693_
timestamp 1728341909
transform 1 0 5050 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2694_
timestamp 1728341909
transform -1 0 5190 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2695_
timestamp 1728341909
transform 1 0 6630 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2696_
timestamp 1728341909
transform 1 0 6570 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2697_
timestamp 1728341909
transform 1 0 6990 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2698_
timestamp 1728341909
transform 1 0 6890 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2699_
timestamp 1728341909
transform -1 0 6330 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2700_
timestamp 1728341909
transform 1 0 5390 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2701_
timestamp 1728341909
transform -1 0 5470 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2702_
timestamp 1728341909
transform -1 0 5550 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2703_
timestamp 1728341909
transform -1 0 5570 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2704_
timestamp 1728341909
transform 1 0 5630 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2705_
timestamp 1728341909
transform 1 0 5890 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2706_
timestamp 1728341909
transform -1 0 6150 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2707_
timestamp 1728341909
transform -1 0 5890 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2708_
timestamp 1728341909
transform -1 0 2290 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2709_
timestamp 1728341909
transform -1 0 4950 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2710_
timestamp 1728341909
transform -1 0 4870 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2711_
timestamp 1728341909
transform -1 0 5070 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2712_
timestamp 1728341909
transform -1 0 5650 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2713_
timestamp 1728341909
transform -1 0 5790 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2714_
timestamp 1728341909
transform -1 0 6090 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2715_
timestamp 1728341909
transform 1 0 5810 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2716_
timestamp 1728341909
transform -1 0 6650 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2717_
timestamp 1728341909
transform 1 0 6590 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2718_
timestamp 1728341909
transform 1 0 6170 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2719_
timestamp 1728341909
transform -1 0 6330 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2720_
timestamp 1728341909
transform 1 0 4630 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2721_
timestamp 1728341909
transform 1 0 4910 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2722_
timestamp 1728341909
transform 1 0 5150 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2723_
timestamp 1728341909
transform -1 0 5410 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2724_
timestamp 1728341909
transform 1 0 6130 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2725_
timestamp 1728341909
transform 1 0 6370 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2726_
timestamp 1728341909
transform -1 0 6130 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__2727_
timestamp 1728341909
transform 1 0 5830 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__2728_
timestamp 1728341909
transform -1 0 4310 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2729_
timestamp 1728341909
transform -1 0 4170 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2730_
timestamp 1728341909
transform -1 0 5210 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2731_
timestamp 1728341909
transform -1 0 5330 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2732_
timestamp 1728341909
transform -1 0 5630 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2733_
timestamp 1728341909
transform -1 0 5890 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2734_
timestamp 1728341909
transform -1 0 5210 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2735_
timestamp 1728341909
transform 1 0 5410 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2736_
timestamp 1728341909
transform -1 0 8330 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__2737_
timestamp 1728341909
transform 1 0 3730 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2738_
timestamp 1728341909
transform 1 0 3910 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2739_
timestamp 1728341909
transform -1 0 3730 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2740_
timestamp 1728341909
transform -1 0 3670 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2741_
timestamp 1728341909
transform -1 0 4010 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2742_
timestamp 1728341909
transform -1 0 4150 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2743_
timestamp 1728341909
transform 1 0 4890 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2744_
timestamp 1728341909
transform 1 0 4630 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__2745_
timestamp 1728341909
transform 1 0 5110 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2746_
timestamp 1728341909
transform 1 0 4610 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2747_
timestamp 1728341909
transform 1 0 5530 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2748_
timestamp 1728341909
transform -1 0 4930 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2749_
timestamp 1728341909
transform -1 0 5290 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2750_
timestamp 1728341909
transform -1 0 5390 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2751_
timestamp 1728341909
transform 1 0 4370 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2752_
timestamp 1728341909
transform 1 0 3870 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2753_
timestamp 1728341909
transform -1 0 3410 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2754_
timestamp 1728341909
transform -1 0 2990 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2755_
timestamp 1728341909
transform 1 0 3250 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2756_
timestamp 1728341909
transform -1 0 3630 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2757_
timestamp 1728341909
transform -1 0 3650 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2758_
timestamp 1728341909
transform -1 0 3630 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2759_
timestamp 1728341909
transform -1 0 3510 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2760_
timestamp 1728341909
transform -1 0 3550 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2761_
timestamp 1728341909
transform -1 0 3690 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2762_
timestamp 1728341909
transform -1 0 3450 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2763_
timestamp 1728341909
transform 1 0 3010 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__2764_
timestamp 1728341909
transform 1 0 3290 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__2765_
timestamp 1728341909
transform -1 0 2610 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2766_
timestamp 1728341909
transform 1 0 3690 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__2767_
timestamp 1728341909
transform -1 0 4390 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2768_
timestamp 1728341909
transform 1 0 4470 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2769_
timestamp 1728341909
transform 1 0 5130 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2770_
timestamp 1728341909
transform -1 0 4630 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2771_
timestamp 1728341909
transform -1 0 4910 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2772_
timestamp 1728341909
transform -1 0 4890 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2773_
timestamp 1728341909
transform 1 0 2650 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2774_
timestamp 1728341909
transform -1 0 2510 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__2775_
timestamp 1728341909
transform 1 0 3870 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2776_
timestamp 1728341909
transform 1 0 4390 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2777_
timestamp 1728341909
transform 1 0 5130 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2778_
timestamp 1728341909
transform -1 0 4630 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2779_
timestamp 1728341909
transform 1 0 3950 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__2780_
timestamp 1728341909
transform 1 0 2730 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__2781_
timestamp 1728341909
transform -1 0 3950 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2782_
timestamp 1728341909
transform -1 0 2750 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2783_
timestamp 1728341909
transform 1 0 2450 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2784_
timestamp 1728341909
transform 1 0 530 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2785_
timestamp 1728341909
transform -1 0 2230 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2786_
timestamp 1728341909
transform 1 0 2490 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2787_
timestamp 1728341909
transform -1 0 2910 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2788_
timestamp 1728341909
transform -1 0 2410 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2789_
timestamp 1728341909
transform -1 0 3710 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2790_
timestamp 1728341909
transform 1 0 3190 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2791_
timestamp 1728341909
transform -1 0 2930 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2792_
timestamp 1728341909
transform -1 0 2830 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2793_
timestamp 1728341909
transform -1 0 2250 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__2794_
timestamp 1728341909
transform 1 0 2130 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2795_
timestamp 1728341909
transform 1 0 770 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2796_
timestamp 1728341909
transform 1 0 1710 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2797_
timestamp 1728341909
transform -1 0 1990 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2798_
timestamp 1728341909
transform 1 0 1210 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2799_
timestamp 1728341909
transform -1 0 1490 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2800_
timestamp 1728341909
transform -1 0 1750 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2801_
timestamp 1728341909
transform 1 0 1710 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2802_
timestamp 1728341909
transform 1 0 1790 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2803_
timestamp 1728341909
transform 1 0 3270 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2804_
timestamp 1728341909
transform -1 0 430 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__2805_
timestamp 1728341909
transform 1 0 6970 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2806_
timestamp 1728341909
transform -1 0 5390 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2807_
timestamp 1728341909
transform -1 0 4990 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2808_
timestamp 1728341909
transform 1 0 3910 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2809_
timestamp 1728341909
transform -1 0 4370 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2810_
timestamp 1728341909
transform -1 0 4730 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2811_
timestamp 1728341909
transform -1 0 4590 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2812_
timestamp 1728341909
transform 1 0 4210 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2813_
timestamp 1728341909
transform 1 0 3970 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__2814_
timestamp 1728341909
transform 1 0 4090 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__2815_
timestamp 1728341909
transform -1 0 4170 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2816_
timestamp 1728341909
transform 1 0 2470 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2817_
timestamp 1728341909
transform -1 0 2750 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__2818_
timestamp 1728341909
transform 1 0 2710 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2819_
timestamp 1728341909
transform 1 0 3150 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2820_
timestamp 1728341909
transform 1 0 3390 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2821_
timestamp 1728341909
transform -1 0 3930 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2822_
timestamp 1728341909
transform -1 0 4730 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2823_
timestamp 1728341909
transform -1 0 1710 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2824_
timestamp 1728341909
transform 1 0 530 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__2825_
timestamp 1728341909
transform 1 0 510 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2826_
timestamp 1728341909
transform -1 0 670 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__2827_
timestamp 1728341909
transform 1 0 1710 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2828_
timestamp 1728341909
transform -1 0 1990 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2829_
timestamp 1728341909
transform 1 0 1230 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2830_
timestamp 1728341909
transform -1 0 1490 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2831_
timestamp 1728341909
transform -1 0 1510 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__2832_
timestamp 1728341909
transform 1 0 2010 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2833_
timestamp 1728341909
transform -1 0 1030 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__2834_
timestamp 1728341909
transform 1 0 850 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__2835_
timestamp 1728341909
transform 1 0 1090 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__2836_
timestamp 1728341909
transform 1 0 1310 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__2837_
timestamp 1728341909
transform 1 0 1630 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__2838_
timestamp 1728341909
transform -1 0 1510 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__2839_
timestamp 1728341909
transform 1 0 790 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__2840_
timestamp 1728341909
transform 1 0 1230 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2841_
timestamp 1728341909
transform 1 0 2030 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2842_
timestamp 1728341909
transform -1 0 1690 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2843_
timestamp 1728341909
transform -1 0 1790 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2844_
timestamp 1728341909
transform -1 0 1550 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__2845_
timestamp 1728341909
transform -1 0 1490 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2846_
timestamp 1728341909
transform 1 0 1270 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2847_
timestamp 1728341909
transform -1 0 1270 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__2848_
timestamp 1728341909
transform -1 0 1250 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2849_
timestamp 1728341909
transform -1 0 1550 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2850_
timestamp 1728341909
transform -1 0 1470 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2851_
timestamp 1728341909
transform -1 0 1010 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2852_
timestamp 1728341909
transform -1 0 1070 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2853_
timestamp 1728341909
transform -1 0 2270 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2854_
timestamp 1728341909
transform 1 0 750 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__2855_
timestamp 1728341909
transform 1 0 2430 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__2856_
timestamp 1728341909
transform -1 0 1950 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__2857_
timestamp 1728341909
transform -1 0 2350 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__2858_
timestamp 1728341909
transform -1 0 2250 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__2859_
timestamp 1728341909
transform -1 0 830 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2860_
timestamp 1728341909
transform 1 0 510 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2861_
timestamp 1728341909
transform -1 0 70 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2862_
timestamp 1728341909
transform -1 0 1030 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__2863_
timestamp 1728341909
transform 1 0 270 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__2864_
timestamp 1728341909
transform -1 0 310 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__2865_
timestamp 1728341909
transform 1 0 4430 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__2866_
timestamp 1728341909
transform 1 0 4450 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2867_
timestamp 1728341909
transform 1 0 5550 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__2868_
timestamp 1728341909
transform -1 0 2930 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2869_
timestamp 1728341909
transform -1 0 3210 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__2870_
timestamp 1728341909
transform -1 0 2270 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__2871_
timestamp 1728341909
transform 1 0 2290 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__2872_
timestamp 1728341909
transform -1 0 4570 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__2873_
timestamp 1728341909
transform 1 0 4310 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__2874_
timestamp 1728341909
transform -1 0 4110 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2875_
timestamp 1728341909
transform -1 0 1670 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2876_
timestamp 1728341909
transform -1 0 810 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2877_
timestamp 1728341909
transform -1 0 3470 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2878_
timestamp 1728341909
transform -1 0 3910 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2879_
timestamp 1728341909
transform -1 0 1250 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2880_
timestamp 1728341909
transform 1 0 1430 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2881_
timestamp 1728341909
transform -1 0 1750 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2882_
timestamp 1728341909
transform -1 0 2430 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2883_
timestamp 1728341909
transform 1 0 4430 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2884_
timestamp 1728341909
transform 1 0 4150 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2885_
timestamp 1728341909
transform 1 0 3090 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2886_
timestamp 1728341909
transform 1 0 4650 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2887_
timestamp 1728341909
transform 1 0 5110 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2888_
timestamp 1728341909
transform 1 0 3370 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2889_
timestamp 1728341909
transform 1 0 3590 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2890_
timestamp 1728341909
transform -1 0 4370 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2891_
timestamp 1728341909
transform -1 0 4110 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2892_
timestamp 1728341909
transform -1 0 1970 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2893_
timestamp 1728341909
transform 1 0 3650 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2894_
timestamp 1728341909
transform 1 0 3850 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2895_
timestamp 1728341909
transform 1 0 4430 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2896_
timestamp 1728341909
transform -1 0 3830 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2897_
timestamp 1728341909
transform -1 0 5830 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2898_
timestamp 1728341909
transform 1 0 5150 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2899_
timestamp 1728341909
transform 1 0 5110 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2900_
timestamp 1728341909
transform 1 0 5370 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2901_
timestamp 1728341909
transform -1 0 4850 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2902_
timestamp 1728341909
transform -1 0 1510 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2903_
timestamp 1728341909
transform 1 0 2170 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2904_
timestamp 1728341909
transform 1 0 2430 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2905_
timestamp 1728341909
transform 1 0 1230 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2906_
timestamp 1728341909
transform 1 0 1010 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2907_
timestamp 1728341909
transform 1 0 1210 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2908_
timestamp 1728341909
transform -1 0 1530 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2909_
timestamp 1728341909
transform -1 0 1750 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2910_
timestamp 1728341909
transform -1 0 1530 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2911_
timestamp 1728341909
transform -1 0 1530 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2912_
timestamp 1728341909
transform -1 0 2450 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2913_
timestamp 1728341909
transform -1 0 1690 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2914_
timestamp 1728341909
transform 1 0 2210 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2915_
timestamp 1728341909
transform 1 0 1990 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2916_
timestamp 1728341909
transform 1 0 1670 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2917_
timestamp 1728341909
transform -1 0 1750 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2918_
timestamp 1728341909
transform 1 0 1690 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2919_
timestamp 1728341909
transform -1 0 2230 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2920_
timestamp 1728341909
transform -1 0 1950 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2921_
timestamp 1728341909
transform -1 0 2010 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2922_
timestamp 1728341909
transform -1 0 1930 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2923_
timestamp 1728341909
transform -1 0 1970 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2924_
timestamp 1728341909
transform -1 0 2930 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2925_
timestamp 1728341909
transform 1 0 3410 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2926_
timestamp 1728341909
transform -1 0 2390 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2927_
timestamp 1728341909
transform -1 0 2430 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2928_
timestamp 1728341909
transform 1 0 4570 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2929_
timestamp 1728341909
transform 1 0 3410 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2930_
timestamp 1728341909
transform -1 0 2690 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2931_
timestamp 1728341909
transform -1 0 2930 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2932_
timestamp 1728341909
transform 1 0 3130 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2933_
timestamp 1728341909
transform -1 0 2690 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2934_
timestamp 1728341909
transform 1 0 2910 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2935_
timestamp 1728341909
transform -1 0 1290 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2936_
timestamp 1728341909
transform -1 0 830 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2937_
timestamp 1728341909
transform 1 0 550 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2938_
timestamp 1728341909
transform 1 0 1710 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2939_
timestamp 1728341909
transform -1 0 1490 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2940_
timestamp 1728341909
transform 1 0 3150 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2941_
timestamp 1728341909
transform 1 0 3150 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2942_
timestamp 1728341909
transform -1 0 3370 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2943_
timestamp 1728341909
transform -1 0 3210 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2944_
timestamp 1728341909
transform -1 0 3710 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2945_
timestamp 1728341909
transform 1 0 3150 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__2946_
timestamp 1728341909
transform 1 0 3590 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__2947_
timestamp 1728341909
transform 1 0 3170 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2948_
timestamp 1728341909
transform -1 0 4170 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2949_
timestamp 1728341909
transform 1 0 3130 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__2950_
timestamp 1728341909
transform 1 0 2450 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2951_
timestamp 1728341909
transform -1 0 2690 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2952_
timestamp 1728341909
transform -1 0 2970 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2953_
timestamp 1728341909
transform -1 0 2170 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2954_
timestamp 1728341909
transform -1 0 2410 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2955_
timestamp 1728341909
transform 1 0 2990 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__2956_
timestamp 1728341909
transform 1 0 3230 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__2957_
timestamp 1728341909
transform 1 0 3730 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__2958_
timestamp 1728341909
transform 1 0 2170 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__2959_
timestamp 1728341909
transform 1 0 3450 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__2960_
timestamp 1728341909
transform 1 0 3570 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__2961_
timestamp 1728341909
transform 1 0 2690 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2962_
timestamp 1728341909
transform 1 0 2430 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2963_
timestamp 1728341909
transform 1 0 2950 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2964_
timestamp 1728341909
transform 1 0 2690 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2965_
timestamp 1728341909
transform -1 0 5770 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2966_
timestamp 1728341909
transform 1 0 4090 0 1 1690
box -12 -8 32 252
use FILL  FILL_2__2967_
timestamp 1728341909
transform -1 0 4570 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2968_
timestamp 1728341909
transform -1 0 4810 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2969_
timestamp 1728341909
transform -1 0 1310 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__2970_
timestamp 1728341909
transform -1 0 1490 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__2971_
timestamp 1728341909
transform -1 0 1510 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2972_
timestamp 1728341909
transform -1 0 1250 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2973_
timestamp 1728341909
transform -1 0 1010 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__2974_
timestamp 1728341909
transform -1 0 1750 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2975_
timestamp 1728341909
transform -1 0 1970 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2976_
timestamp 1728341909
transform 1 0 3850 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2977_
timestamp 1728341909
transform -1 0 4410 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2978_
timestamp 1728341909
transform 1 0 4130 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2979_
timestamp 1728341909
transform 1 0 1510 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2980_
timestamp 1728341909
transform -1 0 990 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2981_
timestamp 1728341909
transform -1 0 750 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2982_
timestamp 1728341909
transform 1 0 2190 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2983_
timestamp 1728341909
transform -1 0 510 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2984_
timestamp 1728341909
transform -1 0 290 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2985_
timestamp 1728341909
transform -1 0 70 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__2986_
timestamp 1728341909
transform -1 0 330 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2987_
timestamp 1728341909
transform -1 0 590 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2988_
timestamp 1728341909
transform -1 0 550 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2989_
timestamp 1728341909
transform 1 0 310 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2990_
timestamp 1728341909
transform 1 0 50 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2991_
timestamp 1728341909
transform -1 0 330 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2992_
timestamp 1728341909
transform -1 0 1990 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__2993_
timestamp 1728341909
transform -1 0 1030 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2994_
timestamp 1728341909
transform -1 0 790 0 1 730
box -12 -8 32 252
use FILL  FILL_2__2995_
timestamp 1728341909
transform 1 0 570 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__2996_
timestamp 1728341909
transform -1 0 510 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__2997_
timestamp 1728341909
transform -1 0 830 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__2998_
timestamp 1728341909
transform -1 0 70 0 1 250
box -12 -8 32 252
use FILL  FILL_2__2999_
timestamp 1728341909
transform -1 0 310 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__3000_
timestamp 1728341909
transform -1 0 70 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__3001_
timestamp 1728341909
transform -1 0 70 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__3002_
timestamp 1728341909
transform -1 0 550 0 1 730
box -12 -8 32 252
use FILL  FILL_2__3003_
timestamp 1728341909
transform -1 0 70 0 1 730
box -12 -8 32 252
use FILL  FILL_2__3004_
timestamp 1728341909
transform -1 0 810 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__3005_
timestamp 1728341909
transform 1 0 770 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__3006_
timestamp 1728341909
transform -1 0 70 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__3007_
timestamp 1728341909
transform 1 0 1770 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3008_
timestamp 1728341909
transform -1 0 1030 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__3009_
timestamp 1728341909
transform -1 0 1290 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__3010_
timestamp 1728341909
transform -1 0 1290 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__3011_
timestamp 1728341909
transform -1 0 1050 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2__3012_
timestamp 1728341909
transform -1 0 1430 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__3013_
timestamp 1728341909
transform -1 0 1210 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__3014_
timestamp 1728341909
transform 1 0 1010 0 1 250
box -12 -8 32 252
use FILL  FILL_2__3015_
timestamp 1728341909
transform -1 0 1510 0 1 250
box -12 -8 32 252
use FILL  FILL_2__3016_
timestamp 1728341909
transform -1 0 1270 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__3017_
timestamp 1728341909
transform -1 0 1250 0 1 250
box -12 -8 32 252
use FILL  FILL_2__3018_
timestamp 1728341909
transform 1 0 1030 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2__3019_
timestamp 1728341909
transform -1 0 1030 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__3020_
timestamp 1728341909
transform -1 0 3670 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3021_
timestamp 1728341909
transform -1 0 5930 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__3022_
timestamp 1728341909
transform 1 0 2770 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3023_
timestamp 1728341909
transform 1 0 2790 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3024_
timestamp 1728341909
transform 1 0 3770 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3025_
timestamp 1728341909
transform -1 0 4190 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__3026_
timestamp 1728341909
transform -1 0 3050 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3027_
timestamp 1728341909
transform -1 0 3450 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__3028_
timestamp 1728341909
transform -1 0 3970 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3029_
timestamp 1728341909
transform -1 0 4470 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3030_
timestamp 1728341909
transform 1 0 3450 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__3031_
timestamp 1728341909
transform -1 0 3730 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__3032_
timestamp 1728341909
transform -1 0 2530 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3033_
timestamp 1728341909
transform -1 0 2550 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3034_
timestamp 1728341909
transform 1 0 2690 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__3035_
timestamp 1728341909
transform -1 0 2950 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__3036_
timestamp 1728341909
transform 1 0 3270 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3037_
timestamp 1728341909
transform -1 0 3710 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__3038_
timestamp 1728341909
transform -1 0 3270 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3039_
timestamp 1728341909
transform 1 0 3010 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3040_
timestamp 1728341909
transform 1 0 2150 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__3041_
timestamp 1728341909
transform 1 0 2690 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__3042_
timestamp 1728341909
transform 1 0 7450 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__3043_
timestamp 1728341909
transform 1 0 6290 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__3044_
timestamp 1728341909
transform 1 0 5310 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__3045_
timestamp 1728341909
transform 1 0 5730 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3046_
timestamp 1728341909
transform 1 0 5450 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__3047_
timestamp 1728341909
transform 1 0 4790 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__3048_
timestamp 1728341909
transform 1 0 5130 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__3049_
timestamp 1728341909
transform 1 0 5830 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3050_
timestamp 1728341909
transform -1 0 6850 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3051_
timestamp 1728341909
transform -1 0 6310 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__3052_
timestamp 1728341909
transform 1 0 6350 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3053_
timestamp 1728341909
transform 1 0 6090 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3054_
timestamp 1728341909
transform 1 0 5830 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3055_
timestamp 1728341909
transform -1 0 5930 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3056_
timestamp 1728341909
transform 1 0 4590 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__3057_
timestamp 1728341909
transform 1 0 4350 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__3058_
timestamp 1728341909
transform -1 0 4470 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3059_
timestamp 1728341909
transform 1 0 4290 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__3060_
timestamp 1728341909
transform -1 0 4270 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__3061_
timestamp 1728341909
transform 1 0 3970 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3062_
timestamp 1728341909
transform -1 0 4790 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__3063_
timestamp 1728341909
transform 1 0 4530 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__3064_
timestamp 1728341909
transform 1 0 5990 0 1 2170
box -12 -8 32 252
use FILL  FILL_2__3065_
timestamp 1728341909
transform 1 0 5770 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__3066_
timestamp 1728341909
transform -1 0 5770 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3067_
timestamp 1728341909
transform -1 0 5910 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__3068_
timestamp 1728341909
transform -1 0 6950 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3069_
timestamp 1728341909
transform -1 0 6450 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3070_
timestamp 1728341909
transform 1 0 6090 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3071_
timestamp 1728341909
transform -1 0 6370 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3072_
timestamp 1728341909
transform 1 0 6570 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__3073_
timestamp 1728341909
transform 1 0 6330 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__3074_
timestamp 1728341909
transform 1 0 390 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__3075_
timestamp 1728341909
transform -1 0 550 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__3076_
timestamp 1728341909
transform -1 0 4250 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3077_
timestamp 1728341909
transform 1 0 1990 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3078_
timestamp 1728341909
transform -1 0 5490 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3079_
timestamp 1728341909
transform 1 0 5030 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3080_
timestamp 1728341909
transform 1 0 4230 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3081_
timestamp 1728341909
transform 1 0 5870 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__3082_
timestamp 1728341909
transform -1 0 6870 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__3083_
timestamp 1728341909
transform 1 0 6030 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__3084_
timestamp 1728341909
transform -1 0 5710 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3085_
timestamp 1728341909
transform -1 0 4990 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3086_
timestamp 1728341909
transform 1 0 5470 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3087_
timestamp 1728341909
transform -1 0 5070 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__3088_
timestamp 1728341909
transform -1 0 5610 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__3089_
timestamp 1728341909
transform -1 0 5570 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__3090_
timestamp 1728341909
transform 1 0 4750 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3091_
timestamp 1728341909
transform -1 0 4710 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3092_
timestamp 1728341909
transform 1 0 5570 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2__3093_
timestamp 1728341909
transform -1 0 3970 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__3094_
timestamp 1728341909
transform 1 0 4410 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__3095_
timestamp 1728341909
transform 1 0 4710 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__3096_
timestamp 1728341909
transform 1 0 4690 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__3097_
timestamp 1728341909
transform 1 0 4930 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__3098_
timestamp 1728341909
transform -1 0 5030 0 1 2650
box -12 -8 32 252
use FILL  FILL_2__3099_
timestamp 1728341909
transform 1 0 5170 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__3100_
timestamp 1728341909
transform -1 0 5570 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__3101_
timestamp 1728341909
transform 1 0 5110 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__3102_
timestamp 1728341909
transform 1 0 4630 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__3103_
timestamp 1728341909
transform 1 0 4850 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__3104_
timestamp 1728341909
transform -1 0 4990 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3105_
timestamp 1728341909
transform 1 0 5310 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__3106_
timestamp 1728341909
transform 1 0 8490 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__3107_
timestamp 1728341909
transform 1 0 8250 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__3108_
timestamp 1728341909
transform 1 0 8010 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__3109_
timestamp 1728341909
transform -1 0 8550 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3110_
timestamp 1728341909
transform -1 0 8310 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3111_
timestamp 1728341909
transform 1 0 4490 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3112_
timestamp 1728341909
transform 1 0 4730 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3113_
timestamp 1728341909
transform -1 0 1250 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3114_
timestamp 1728341909
transform 1 0 750 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3115_
timestamp 1728341909
transform 1 0 4430 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__3116_
timestamp 1728341909
transform -1 0 4050 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3117_
timestamp 1728341909
transform -1 0 310 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__3118_
timestamp 1728341909
transform -1 0 70 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__3119_
timestamp 1728341909
transform -1 0 4910 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__3120_
timestamp 1728341909
transform 1 0 4410 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3121_
timestamp 1728341909
transform 1 0 5150 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__3122_
timestamp 1728341909
transform -1 0 4450 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3123_
timestamp 1728341909
transform -1 0 3710 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3124_
timestamp 1728341909
transform -1 0 3930 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3125_
timestamp 1728341909
transform -1 0 3670 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3126_
timestamp 1728341909
transform 1 0 4690 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3127_
timestamp 1728341909
transform 1 0 4710 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3128_
timestamp 1728341909
transform 1 0 4630 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__3129_
timestamp 1728341909
transform 1 0 3710 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__3130_
timestamp 1728341909
transform -1 0 1810 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3131_
timestamp 1728341909
transform -1 0 1310 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3132_
timestamp 1728341909
transform 1 0 1030 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3133_
timestamp 1728341909
transform 1 0 3890 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3134_
timestamp 1728341909
transform 1 0 3470 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3135_
timestamp 1728341909
transform 1 0 3210 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3136_
timestamp 1728341909
transform 1 0 3690 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3137_
timestamp 1728341909
transform 1 0 3950 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3138_
timestamp 1728341909
transform -1 0 3990 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3139_
timestamp 1728341909
transform 1 0 1050 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3140_
timestamp 1728341909
transform 1 0 790 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3141_
timestamp 1728341909
transform -1 0 3970 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3142_
timestamp 1728341909
transform 1 0 3730 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3143_
timestamp 1728341909
transform -1 0 4170 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3144_
timestamp 1728341909
transform -1 0 3450 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3145_
timestamp 1728341909
transform 1 0 3190 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3146_
timestamp 1728341909
transform -1 0 3270 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3147_
timestamp 1728341909
transform 1 0 3510 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3148_
timestamp 1728341909
transform -1 0 3470 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3149_
timestamp 1728341909
transform -1 0 3450 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__3150_
timestamp 1728341909
transform 1 0 2030 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3151_
timestamp 1728341909
transform -1 0 2270 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3152_
timestamp 1728341909
transform 1 0 7510 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3153_
timestamp 1728341909
transform 1 0 4430 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3154_
timestamp 1728341909
transform -1 0 770 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3155_
timestamp 1728341909
transform 1 0 990 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3156_
timestamp 1728341909
transform 1 0 2950 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3157_
timestamp 1728341909
transform -1 0 2730 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3158_
timestamp 1728341909
transform 1 0 1950 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3159_
timestamp 1728341909
transform 1 0 2490 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3160_
timestamp 1728341909
transform 1 0 3110 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3161_
timestamp 1728341909
transform -1 0 2650 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3162_
timestamp 1728341909
transform -1 0 2430 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3163_
timestamp 1728341909
transform -1 0 1530 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3164_
timestamp 1728341909
transform 1 0 1230 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3165_
timestamp 1728341909
transform -1 0 310 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3166_
timestamp 1728341909
transform -1 0 70 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3167_
timestamp 1728341909
transform 1 0 2030 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3168_
timestamp 1728341909
transform 1 0 1970 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3169_
timestamp 1728341909
transform -1 0 2270 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3170_
timestamp 1728341909
transform 1 0 2010 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3171_
timestamp 1728341909
transform -1 0 2210 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3172_
timestamp 1728341909
transform 1 0 1870 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__3173_
timestamp 1728341909
transform -1 0 1750 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3174_
timestamp 1728341909
transform -1 0 1770 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3175_
timestamp 1728341909
transform -1 0 3010 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3176_
timestamp 1728341909
transform -1 0 2810 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3177_
timestamp 1728341909
transform 1 0 2250 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3178_
timestamp 1728341909
transform 1 0 2590 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3179_
timestamp 1728341909
transform 1 0 2250 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3180_
timestamp 1728341909
transform 1 0 3190 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3181_
timestamp 1728341909
transform -1 0 2910 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3182_
timestamp 1728341909
transform -1 0 2990 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3183_
timestamp 1728341909
transform 1 0 2750 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3184_
timestamp 1728341909
transform -1 0 2510 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3185_
timestamp 1728341909
transform -1 0 2510 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3186_
timestamp 1728341909
transform 1 0 1990 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3187_
timestamp 1728341909
transform -1 0 330 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3188_
timestamp 1728341909
transform -1 0 70 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3189_
timestamp 1728341909
transform 1 0 1010 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3190_
timestamp 1728341909
transform -1 0 810 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3191_
timestamp 1728341909
transform -1 0 1070 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3192_
timestamp 1728341909
transform 1 0 1690 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3193_
timestamp 1728341909
transform 1 0 1430 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3194_
timestamp 1728341909
transform 1 0 3230 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3195_
timestamp 1728341909
transform 1 0 3190 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__3196_
timestamp 1728341909
transform 1 0 1930 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3197_
timestamp 1728341909
transform -1 0 2510 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__3198_
timestamp 1728341909
transform -1 0 2090 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3199_
timestamp 1728341909
transform -1 0 2350 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3200_
timestamp 1728341909
transform 1 0 790 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3201_
timestamp 1728341909
transform -1 0 1030 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3202_
timestamp 1728341909
transform 1 0 1030 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3203_
timestamp 1728341909
transform -1 0 1290 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3204_
timestamp 1728341909
transform -1 0 550 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3205_
timestamp 1728341909
transform -1 0 550 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3206_
timestamp 1728341909
transform 1 0 1050 0 -1 4090
box -12 -8 32 252
use FILL  FILL_2__3207_
timestamp 1728341909
transform -1 0 310 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3208_
timestamp 1728341909
transform -1 0 70 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3209_
timestamp 1728341909
transform 1 0 290 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3210_
timestamp 1728341909
transform -1 0 70 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3211_
timestamp 1728341909
transform -1 0 1550 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3212_
timestamp 1728341909
transform -1 0 1290 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3213_
timestamp 1728341909
transform 1 0 1570 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3214_
timestamp 1728341909
transform 1 0 1310 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3215_
timestamp 1728341909
transform -1 0 1270 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3216_
timestamp 1728341909
transform 1 0 1010 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3217_
timestamp 1728341909
transform -1 0 310 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3218_
timestamp 1728341909
transform -1 0 70 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3219_
timestamp 1728341909
transform -1 0 1590 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3220_
timestamp 1728341909
transform 1 0 1810 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3221_
timestamp 1728341909
transform -1 0 330 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3222_
timestamp 1728341909
transform -1 0 70 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3223_
timestamp 1728341909
transform -1 0 810 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__3224_
timestamp 1728341909
transform 1 0 530 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3225_
timestamp 1728341909
transform -1 0 310 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3226_
timestamp 1728341909
transform -1 0 70 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3227_
timestamp 1728341909
transform -1 0 330 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__3228_
timestamp 1728341909
transform -1 0 70 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__3229_
timestamp 1728341909
transform -1 0 1990 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__3230_
timestamp 1728341909
transform 1 0 1710 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__3231_
timestamp 1728341909
transform 1 0 1510 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__3232_
timestamp 1728341909
transform -1 0 1770 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__3233_
timestamp 1728341909
transform 1 0 1070 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3234_
timestamp 1728341909
transform -1 0 1350 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3235_
timestamp 1728341909
transform 1 0 1030 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3236_
timestamp 1728341909
transform 1 0 1290 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3237_
timestamp 1728341909
transform 1 0 2210 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__3238_
timestamp 1728341909
transform 1 0 2450 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2__3239_
timestamp 1728341909
transform -1 0 550 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3240_
timestamp 1728341909
transform -1 0 790 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3241_
timestamp 1728341909
transform 1 0 9690 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__3242_
timestamp 1728341909
transform -1 0 9030 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2__3243_
timestamp 1728341909
transform 1 0 9450 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__3244_
timestamp 1728341909
transform 1 0 8750 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__3245_
timestamp 1728341909
transform 1 0 9050 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3246_
timestamp 1728341909
transform -1 0 9570 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3247_
timestamp 1728341909
transform 1 0 10470 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3248_
timestamp 1728341909
transform 1 0 10730 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3249_
timestamp 1728341909
transform -1 0 9470 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__3250_
timestamp 1728341909
transform 1 0 9390 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3251_
timestamp 1728341909
transform 1 0 9230 0 1 3130
box -12 -8 32 252
use FILL  FILL_2__3252_
timestamp 1728341909
transform -1 0 9250 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__3253_
timestamp 1728341909
transform -1 0 7870 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3254_
timestamp 1728341909
transform -1 0 8130 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3255_
timestamp 1728341909
transform -1 0 9310 0 1 3610
box -12 -8 32 252
use FILL  FILL_2__3256_
timestamp 1728341909
transform 1 0 8250 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3257_
timestamp 1728341909
transform 1 0 8010 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3258_
timestamp 1728341909
transform 1 0 8550 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3259_
timestamp 1728341909
transform 1 0 9490 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3260_
timestamp 1728341909
transform -1 0 10850 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__3261_
timestamp 1728341909
transform -1 0 10390 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3262_
timestamp 1728341909
transform 1 0 9970 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3263_
timestamp 1728341909
transform 1 0 9650 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__3264_
timestamp 1728341909
transform 1 0 8990 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2__3265_
timestamp 1728341909
transform -1 0 9730 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3266_
timestamp 1728341909
transform 1 0 9750 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3267_
timestamp 1728341909
transform -1 0 9650 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3268_
timestamp 1728341909
transform -1 0 9990 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3269_
timestamp 1728341909
transform -1 0 10490 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3270_
timestamp 1728341909
transform 1 0 10210 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3271_
timestamp 1728341909
transform -1 0 10030 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2__3272_
timestamp 1728341909
transform 1 0 10250 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2__3273_
timestamp 1728341909
transform -1 0 10150 0 1 4570
box -12 -8 32 252
use FILL  FILL_2__3274_
timestamp 1728341909
transform -1 0 10250 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3275_
timestamp 1728341909
transform 1 0 9570 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__3276_
timestamp 1728341909
transform -1 0 9190 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3277_
timestamp 1728341909
transform -1 0 10650 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3278_
timestamp 1728341909
transform 1 0 10110 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3279_
timestamp 1728341909
transform -1 0 9890 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3280_
timestamp 1728341909
transform 1 0 9230 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__3281_
timestamp 1728341909
transform 1 0 8990 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__3282_
timestamp 1728341909
transform -1 0 6870 0 1 4090
box -12 -8 32 252
use FILL  FILL_2__3283_
timestamp 1728341909
transform -1 0 6810 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3284_
timestamp 1728341909
transform 1 0 6570 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2__3285_
timestamp 1728341909
transform 1 0 7010 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3286_
timestamp 1728341909
transform -1 0 7270 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3287_
timestamp 1728341909
transform -1 0 6630 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3288_
timestamp 1728341909
transform -1 0 6850 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3289_
timestamp 1728341909
transform -1 0 6810 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__3290_
timestamp 1728341909
transform 1 0 6530 0 1 5530
box -12 -8 32 252
use FILL  FILL_2__3291_
timestamp 1728341909
transform 1 0 7030 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3292_
timestamp 1728341909
transform -1 0 7290 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3293_
timestamp 1728341909
transform 1 0 7130 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3294_
timestamp 1728341909
transform 1 0 6870 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3295_
timestamp 1728341909
transform 1 0 6070 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3296_
timestamp 1728341909
transform 1 0 5810 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3297_
timestamp 1728341909
transform 1 0 5430 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3298_
timestamp 1728341909
transform 1 0 5170 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3299_
timestamp 1728341909
transform 1 0 5610 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3300_
timestamp 1728341909
transform 1 0 5370 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3301_
timestamp 1728341909
transform 1 0 6870 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2__3302_
timestamp 1728341909
transform 1 0 2950 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3303_
timestamp 1728341909
transform -1 0 3010 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3304_
timestamp 1728341909
transform 1 0 1950 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3305_
timestamp 1728341909
transform -1 0 2210 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3306_
timestamp 1728341909
transform 1 0 3870 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3307_
timestamp 1728341909
transform -1 0 4810 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3308_
timestamp 1728341909
transform -1 0 70 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__3309_
timestamp 1728341909
transform -1 0 70 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3310_
timestamp 1728341909
transform -1 0 750 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__3311_
timestamp 1728341909
transform -1 0 790 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3312_
timestamp 1728341909
transform -1 0 290 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__3313_
timestamp 1728341909
transform -1 0 330 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3314_
timestamp 1728341909
transform -1 0 70 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3315_
timestamp 1728341909
transform -1 0 70 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3316_
timestamp 1728341909
transform -1 0 570 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3317_
timestamp 1728341909
transform -1 0 790 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3449_
timestamp 1728341909
transform -1 0 3810 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3450_
timestamp 1728341909
transform 1 0 2970 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3451_
timestamp 1728341909
transform 1 0 3090 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3452_
timestamp 1728341909
transform -1 0 3350 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3453_
timestamp 1728341909
transform 1 0 3210 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3454_
timestamp 1728341909
transform -1 0 3570 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3455_
timestamp 1728341909
transform 1 0 9950 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3456_
timestamp 1728341909
transform 1 0 9510 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3457_
timestamp 1728341909
transform -1 0 9790 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3458_
timestamp 1728341909
transform -1 0 9950 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3459_
timestamp 1728341909
transform 1 0 10390 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3460_
timestamp 1728341909
transform -1 0 10690 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3461_
timestamp 1728341909
transform -1 0 10450 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3462_
timestamp 1728341909
transform -1 0 10010 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3463_
timestamp 1728341909
transform 1 0 10410 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3464_
timestamp 1728341909
transform -1 0 10210 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3465_
timestamp 1728341909
transform 1 0 10170 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2__3466_
timestamp 1728341909
transform -1 0 10190 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3467_
timestamp 1728341909
transform 1 0 8250 0 1 6010
box -12 -8 32 252
use FILL  FILL_2__3468_
timestamp 1728341909
transform 1 0 9090 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__3469_
timestamp 1728341909
transform 1 0 8550 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3470_
timestamp 1728341909
transform -1 0 8490 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3471_
timestamp 1728341909
transform 1 0 8630 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__3472_
timestamp 1728341909
transform 1 0 8870 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__3473_
timestamp 1728341909
transform -1 0 8690 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3474_
timestamp 1728341909
transform -1 0 8810 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3475_
timestamp 1728341909
transform -1 0 8930 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3476_
timestamp 1728341909
transform 1 0 9730 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3477_
timestamp 1728341909
transform 1 0 9170 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3478_
timestamp 1728341909
transform -1 0 9050 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3479_
timestamp 1728341909
transform 1 0 10530 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__3480_
timestamp 1728341909
transform -1 0 10090 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__3481_
timestamp 1728341909
transform -1 0 9950 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3482_
timestamp 1728341909
transform -1 0 9750 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__3483_
timestamp 1728341909
transform 1 0 10890 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3484_
timestamp 1728341909
transform 1 0 10870 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3485_
timestamp 1728341909
transform 1 0 11150 0 1 6490
box -12 -8 32 252
use FILL  FILL_2__3486_
timestamp 1728341909
transform 1 0 11110 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3487_
timestamp 1728341909
transform 1 0 10870 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3488_
timestamp 1728341909
transform 1 0 9510 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3489_
timestamp 1728341909
transform 1 0 9410 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3490_
timestamp 1728341909
transform -1 0 9670 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3491_
timestamp 1728341909
transform -1 0 9690 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3492_
timestamp 1728341909
transform 1 0 9890 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3493_
timestamp 1728341909
transform 1 0 10150 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3494_
timestamp 1728341909
transform 1 0 10290 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__3495_
timestamp 1728341909
transform -1 0 8790 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3496_
timestamp 1728341909
transform 1 0 9410 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3497_
timestamp 1728341909
transform 1 0 9930 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3498_
timestamp 1728341909
transform 1 0 9790 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__3499_
timestamp 1728341909
transform 1 0 9210 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3500_
timestamp 1728341909
transform -1 0 9470 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3501_
timestamp 1728341909
transform -1 0 9710 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3502_
timestamp 1728341909
transform 1 0 9550 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__3503_
timestamp 1728341909
transform 1 0 10030 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__3504_
timestamp 1728341909
transform -1 0 9990 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3505_
timestamp 1728341909
transform 1 0 10230 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3506_
timestamp 1728341909
transform 1 0 10750 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__3507_
timestamp 1728341909
transform -1 0 9370 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__3508_
timestamp 1728341909
transform -1 0 8490 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3509_
timestamp 1728341909
transform 1 0 8410 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__3510_
timestamp 1728341909
transform 1 0 9190 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3511_
timestamp 1728341909
transform -1 0 8950 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3512_
timestamp 1728341909
transform 1 0 8690 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3513_
timestamp 1728341909
transform -1 0 8970 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3514_
timestamp 1728341909
transform -1 0 8730 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3515_
timestamp 1728341909
transform -1 0 9130 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__3516_
timestamp 1728341909
transform 1 0 10970 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__3517_
timestamp 1728341909
transform -1 0 10290 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__3518_
timestamp 1728341909
transform 1 0 10370 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3519_
timestamp 1728341909
transform 1 0 10850 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3520_
timestamp 1728341909
transform -1 0 11150 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3521_
timestamp 1728341909
transform 1 0 7470 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3522_
timestamp 1728341909
transform -1 0 7990 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3523_
timestamp 1728341909
transform 1 0 8730 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3524_
timestamp 1728341909
transform 1 0 8510 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3525_
timestamp 1728341909
transform 1 0 8930 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3526_
timestamp 1728341909
transform -1 0 9210 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3527_
timestamp 1728341909
transform -1 0 8270 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3528_
timestamp 1728341909
transform -1 0 9910 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3529_
timestamp 1728341909
transform 1 0 10010 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__3530_
timestamp 1728341909
transform 1 0 10110 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3531_
timestamp 1728341909
transform -1 0 10150 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3532_
timestamp 1728341909
transform 1 0 10290 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__3533_
timestamp 1728341909
transform -1 0 8210 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3534_
timestamp 1728341909
transform -1 0 8470 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3535_
timestamp 1728341909
transform -1 0 8030 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3536_
timestamp 1728341909
transform -1 0 8250 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3537_
timestamp 1728341909
transform 1 0 8350 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__3538_
timestamp 1728341909
transform -1 0 8630 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__3539_
timestamp 1728341909
transform -1 0 9530 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__3540_
timestamp 1728341909
transform 1 0 9750 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__3541_
timestamp 1728341909
transform -1 0 9830 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__3542_
timestamp 1728341909
transform -1 0 7490 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3543_
timestamp 1728341909
transform -1 0 7750 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3544_
timestamp 1728341909
transform 1 0 7970 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3545_
timestamp 1728341909
transform 1 0 8830 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__3546_
timestamp 1728341909
transform -1 0 8270 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3547_
timestamp 1728341909
transform 1 0 8690 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3548_
timestamp 1728341909
transform -1 0 8950 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3549_
timestamp 1728341909
transform -1 0 8910 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__3550_
timestamp 1728341909
transform 1 0 8890 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3551_
timestamp 1728341909
transform 1 0 9170 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3552_
timestamp 1728341909
transform 1 0 9310 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__3553_
timestamp 1728341909
transform 1 0 9050 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__3554_
timestamp 1728341909
transform 1 0 8970 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__3555_
timestamp 1728341909
transform -1 0 8550 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3556_
timestamp 1728341909
transform 1 0 8450 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3557_
timestamp 1728341909
transform -1 0 8110 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__3558_
timestamp 1728341909
transform -1 0 7750 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3559_
timestamp 1728341909
transform 1 0 7710 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3560_
timestamp 1728341909
transform 1 0 8230 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3561_
timestamp 1728341909
transform -1 0 7970 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3562_
timestamp 1728341909
transform -1 0 8970 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3563_
timestamp 1728341909
transform -1 0 8950 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__3564_
timestamp 1728341909
transform 1 0 10050 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__3565_
timestamp 1728341909
transform -1 0 9970 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__3566_
timestamp 1728341909
transform 1 0 9890 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3567_
timestamp 1728341909
transform 1 0 9970 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__3568_
timestamp 1728341909
transform 1 0 10190 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__3569_
timestamp 1728341909
transform 1 0 10190 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__3570_
timestamp 1728341909
transform 1 0 10650 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__3571_
timestamp 1728341909
transform -1 0 10630 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3572_
timestamp 1728341909
transform -1 0 11130 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3573_
timestamp 1728341909
transform 1 0 11010 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__3574_
timestamp 1728341909
transform 1 0 10750 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__3575_
timestamp 1728341909
transform 1 0 11150 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__3576_
timestamp 1728341909
transform 1 0 9930 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__3577_
timestamp 1728341909
transform -1 0 11170 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__3578_
timestamp 1728341909
transform 1 0 10770 0 -1 9850
box -12 -8 32 252
use FILL  FILL_2__3579_
timestamp 1728341909
transform -1 0 10470 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__3580_
timestamp 1728341909
transform -1 0 9170 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3581_
timestamp 1728341909
transform -1 0 8870 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__3582_
timestamp 1728341909
transform 1 0 8710 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__3583_
timestamp 1728341909
transform -1 0 9030 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__3584_
timestamp 1728341909
transform 1 0 8770 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__3585_
timestamp 1728341909
transform -1 0 9510 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__3586_
timestamp 1728341909
transform 1 0 9090 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__3587_
timestamp 1728341909
transform -1 0 9230 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__3588_
timestamp 1728341909
transform 1 0 9250 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__3589_
timestamp 1728341909
transform 1 0 9970 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__3590_
timestamp 1728341909
transform -1 0 10230 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__3591_
timestamp 1728341909
transform 1 0 9710 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__3592_
timestamp 1728341909
transform 1 0 9730 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__3593_
timestamp 1728341909
transform -1 0 9510 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__3594_
timestamp 1728341909
transform 1 0 10350 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3595_
timestamp 1728341909
transform 1 0 10910 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__3596_
timestamp 1728341909
transform -1 0 10870 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3597_
timestamp 1728341909
transform 1 0 10510 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__3598_
timestamp 1728341909
transform 1 0 11150 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__3599_
timestamp 1728341909
transform 1 0 11110 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3600_
timestamp 1728341909
transform 1 0 10990 0 -1 9370
box -12 -8 32 252
use FILL  FILL_2__3601_
timestamp 1728341909
transform 1 0 10170 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3602_
timestamp 1728341909
transform 1 0 10410 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3603_
timestamp 1728341909
transform 1 0 10470 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3604_
timestamp 1728341909
transform 1 0 10690 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3605_
timestamp 1728341909
transform 1 0 11170 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3606_
timestamp 1728341909
transform 1 0 10650 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3607_
timestamp 1728341909
transform -1 0 9950 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3608_
timestamp 1728341909
transform -1 0 10190 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3609_
timestamp 1728341909
transform 1 0 10690 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3610_
timestamp 1728341909
transform 1 0 9510 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3611_
timestamp 1728341909
transform 1 0 9310 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__3612_
timestamp 1728341909
transform 1 0 9570 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__3613_
timestamp 1728341909
transform 1 0 9430 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3614_
timestamp 1728341909
transform -1 0 9830 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__3615_
timestamp 1728341909
transform -1 0 9710 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3616_
timestamp 1728341909
transform -1 0 9010 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3617_
timestamp 1728341909
transform -1 0 9270 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3618_
timestamp 1728341909
transform 1 0 9750 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3619_
timestamp 1728341909
transform 1 0 10910 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3620_
timestamp 1728341909
transform -1 0 10650 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3621_
timestamp 1728341909
transform -1 0 10430 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3622_
timestamp 1728341909
transform 1 0 10670 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3623_
timestamp 1728341909
transform 1 0 9970 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3624_
timestamp 1728341909
transform 1 0 10690 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3625_
timestamp 1728341909
transform 1 0 10790 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__3626_
timestamp 1728341909
transform -1 0 10690 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3627_
timestamp 1728341909
transform -1 0 9670 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3628_
timestamp 1728341909
transform -1 0 10410 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3629_
timestamp 1728341909
transform 1 0 10630 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3630_
timestamp 1728341909
transform 1 0 10430 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3631_
timestamp 1728341909
transform -1 0 10590 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__3632_
timestamp 1728341909
transform -1 0 10930 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__3633_
timestamp 1728341909
transform 1 0 10890 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__3634_
timestamp 1728341909
transform -1 0 10710 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__3635_
timestamp 1728341909
transform -1 0 10430 0 1 10810
box -12 -8 32 252
use FILL  FILL_2__3636_
timestamp 1728341909
transform -1 0 10530 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__3637_
timestamp 1728341909
transform -1 0 10690 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__3638_
timestamp 1728341909
transform -1 0 10610 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3639_
timestamp 1728341909
transform -1 0 10450 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__3640_
timestamp 1728341909
transform -1 0 10910 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3641_
timestamp 1728341909
transform -1 0 10650 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3642_
timestamp 1728341909
transform -1 0 10970 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3643_
timestamp 1728341909
transform 1 0 10890 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3644_
timestamp 1728341909
transform -1 0 10450 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3645_
timestamp 1728341909
transform -1 0 10190 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3646_
timestamp 1728341909
transform -1 0 10950 0 -1 8890
box -12 -8 32 252
use FILL  FILL_2__3647_
timestamp 1728341909
transform 1 0 11050 0 1 250
box -12 -8 32 252
use FILL  FILL_2__3648_
timestamp 1728341909
transform 1 0 11130 0 1 8410
box -12 -8 32 252
use FILL  FILL_2__3649_
timestamp 1728341909
transform 1 0 10210 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3650_
timestamp 1728341909
transform 1 0 10330 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__3651_
timestamp 1728341909
transform 1 0 10430 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3652_
timestamp 1728341909
transform -1 0 10390 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3653_
timestamp 1728341909
transform 1 0 10610 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3654_
timestamp 1728341909
transform 1 0 8410 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3655_
timestamp 1728341909
transform -1 0 8670 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3656_
timestamp 1728341909
transform 1 0 8250 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__3657_
timestamp 1728341909
transform -1 0 8630 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__3658_
timestamp 1728341909
transform -1 0 8530 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__3659_
timestamp 1728341909
transform -1 0 8270 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2__3660_
timestamp 1728341909
transform -1 0 8390 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__3661_
timestamp 1728341909
transform -1 0 9250 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__3662_
timestamp 1728341909
transform -1 0 9490 0 1 10330
box -12 -8 32 252
use FILL  FILL_2__3663_
timestamp 1728341909
transform 1 0 9410 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3664_
timestamp 1728341909
transform -1 0 9650 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3665_
timestamp 1728341909
transform 1 0 8250 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3666_
timestamp 1728341909
transform -1 0 8490 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3667_
timestamp 1728341909
transform -1 0 9210 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3668_
timestamp 1728341909
transform -1 0 10430 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3669_
timestamp 1728341909
transform -1 0 10170 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3670_
timestamp 1728341909
transform -1 0 9930 0 1 9370
box -12 -8 32 252
use FILL  FILL_2__3671_
timestamp 1728341909
transform 1 0 8290 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3672_
timestamp 1728341909
transform 1 0 8530 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3673_
timestamp 1728341909
transform -1 0 9450 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3674_
timestamp 1728341909
transform -1 0 9910 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3675_
timestamp 1728341909
transform 1 0 10130 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3676_
timestamp 1728341909
transform -1 0 10170 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3677_
timestamp 1728341909
transform 1 0 9410 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3678_
timestamp 1728341909
transform -1 0 9250 0 -1 6970
box -12 -8 32 252
use FILL  FILL_2__3691_
timestamp 1728341909
transform 1 0 7730 0 1 250
box -12 -8 32 252
use FILL  FILL_2__3692_
timestamp 1728341909
transform -1 0 7990 0 1 250
box -12 -8 32 252
use FILL  FILL_2__3693_
timestamp 1728341909
transform -1 0 1970 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3694_
timestamp 1728341909
transform -1 0 70 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3695_
timestamp 1728341909
transform 1 0 570 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3696_
timestamp 1728341909
transform -1 0 70 0 1 9850
box -12 -8 32 252
use FILL  FILL_2__3697_
timestamp 1728341909
transform -1 0 70 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__3698_
timestamp 1728341909
transform -1 0 310 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2__3699_
timestamp 1728341909
transform 1 0 6130 0 1 1210
box -12 -8 32 252
use FILL  FILL_2__3700_
timestamp 1728341909
transform -1 0 6290 0 -1 730
box -12 -8 32 252
use FILL  FILL_2__3701_
timestamp 1728341909
transform -1 0 6270 0 1 250
box -12 -8 32 252
use FILL  FILL_2__3702_
timestamp 1728341909
transform -1 0 5250 0 1 5050
box -12 -8 32 252
use FILL  FILL_2__3703_
timestamp 1728341909
transform -1 0 3490 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__3704_
timestamp 1728341909
transform -1 0 3270 0 -1 250
box -12 -8 32 252
use FILL  FILL_2__3705_
timestamp 1728341909
transform -1 0 70 0 1 8890
box -12 -8 32 252
use FILL  FILL_2__3706_
timestamp 1728341909
transform -1 0 1310 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2__3707_
timestamp 1728341909
transform 1 0 11130 0 1 6970
box -12 -8 32 252
use FILL  FILL_2__3708_
timestamp 1728341909
transform 1 0 11130 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2__3709_
timestamp 1728341909
transform 1 0 11150 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3710_
timestamp 1728341909
transform 1 0 10910 0 1 7450
box -12 -8 32 252
use FILL  FILL_2__3711_
timestamp 1728341909
transform 1 0 11130 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2__3712_
timestamp 1728341909
transform 1 0 10910 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3713_
timestamp 1728341909
transform 1 0 11030 0 1 7930
box -12 -8 32 252
use FILL  FILL_2__3714_
timestamp 1728341909
transform 1 0 11150 0 -1 8410
box -12 -8 32 252
use FILL  FILL_2__3715_
timestamp 1728341909
transform 1 0 11130 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert0
timestamp 1728341909
transform 1 0 7770 0 1 10810
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert1
timestamp 1728341909
transform 1 0 8990 0 1 1690
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert2
timestamp 1728341909
transform 1 0 9190 0 1 6970
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert3
timestamp 1728341909
transform 1 0 5670 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert4
timestamp 1728341909
transform 1 0 6770 0 1 1690
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert5
timestamp 1728341909
transform -1 0 4030 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert6
timestamp 1728341909
transform 1 0 7190 0 1 10330
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert7
timestamp 1728341909
transform -1 0 4110 0 1 4090
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert8
timestamp 1728341909
transform -1 0 7550 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert9
timestamp 1728341909
transform 1 0 4470 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert10
timestamp 1728341909
transform -1 0 590 0 1 4090
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert11
timestamp 1728341909
transform -1 0 4790 0 1 2650
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert12
timestamp 1728341909
transform 1 0 750 0 1 5530
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert13
timestamp 1728341909
transform -1 0 5890 0 1 7450
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert14
timestamp 1728341909
transform 1 0 4530 0 1 2650
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert15
timestamp 1728341909
transform 1 0 5610 0 -1 5050
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert16
timestamp 1728341909
transform 1 0 2690 0 1 8410
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert17
timestamp 1728341909
transform 1 0 4190 0 1 6490
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert18
timestamp 1728341909
transform -1 0 70 0 1 2650
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert19
timestamp 1728341909
transform -1 0 330 0 1 8410
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert20
timestamp 1728341909
transform 1 0 530 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert21
timestamp 1728341909
transform -1 0 7070 0 1 4570
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert22
timestamp 1728341909
transform -1 0 10450 0 1 4090
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert23
timestamp 1728341909
transform -1 0 8790 0 1 4090
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert24
timestamp 1728341909
transform 1 0 8510 0 1 3130
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert25
timestamp 1728341909
transform -1 0 7070 0 1 3130
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert37
timestamp 1728341909
transform -1 0 990 0 1 5530
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert38
timestamp 1728341909
transform 1 0 1270 0 1 4570
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert39
timestamp 1728341909
transform -1 0 1030 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert40
timestamp 1728341909
transform -1 0 2730 0 -1 6010
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert41
timestamp 1728341909
transform 1 0 9530 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert42
timestamp 1728341909
transform 1 0 8850 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert43
timestamp 1728341909
transform -1 0 8770 0 -1 3610
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert44
timestamp 1728341909
transform -1 0 8990 0 1 4570
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert45
timestamp 1728341909
transform 1 0 3850 0 1 4090
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert46
timestamp 1728341909
transform 1 0 5210 0 1 4090
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert47
timestamp 1728341909
transform 1 0 4310 0 1 2650
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert48
timestamp 1728341909
transform 1 0 5430 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert49
timestamp 1728341909
transform -1 0 2230 0 1 2650
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert50
timestamp 1728341909
transform 1 0 8310 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert51
timestamp 1728341909
transform -1 0 10410 0 1 4570
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert52
timestamp 1728341909
transform -1 0 9450 0 1 4570
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert53
timestamp 1728341909
transform -1 0 9530 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert54
timestamp 1728341909
transform -1 0 8370 0 -1 3130
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert55
timestamp 1728341909
transform -1 0 330 0 1 730
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert56
timestamp 1728341909
transform 1 0 5010 0 -1 1210
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert57
timestamp 1728341909
transform 1 0 4610 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert58
timestamp 1728341909
transform 1 0 1930 0 1 1690
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert59
timestamp 1728341909
transform 1 0 4370 0 1 730
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert60
timestamp 1728341909
transform -1 0 8750 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert61
timestamp 1728341909
transform 1 0 10150 0 -1 7450
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert62
timestamp 1728341909
transform 1 0 9190 0 -1 10330
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert63
timestamp 1728341909
transform 1 0 9270 0 1 7450
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert64
timestamp 1728341909
transform 1 0 8610 0 1 1210
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert65
timestamp 1728341909
transform -1 0 5010 0 1 4090
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert66
timestamp 1728341909
transform 1 0 5750 0 1 2650
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert67
timestamp 1728341909
transform 1 0 6590 0 1 5050
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert68
timestamp 1728341909
transform 1 0 7590 0 -1 2650
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert69
timestamp 1728341909
transform -1 0 6070 0 1 1690
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert70
timestamp 1728341909
transform 1 0 8750 0 -1 2170
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert71
timestamp 1728341909
transform 1 0 2450 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert72
timestamp 1728341909
transform 1 0 3890 0 1 1210
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert73
timestamp 1728341909
transform 1 0 2690 0 1 2650
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert74
timestamp 1728341909
transform -1 0 3690 0 -1 1690
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert75
timestamp 1728341909
transform -1 0 770 0 1 2170
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert76
timestamp 1728341909
transform 1 0 8750 0 1 4570
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert77
timestamp 1728341909
transform -1 0 8490 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert78
timestamp 1728341909
transform 1 0 8950 0 -1 5530
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert79
timestamp 1728341909
transform -1 0 9210 0 1 4570
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert80
timestamp 1728341909
transform 1 0 4190 0 -1 6490
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert81
timestamp 1728341909
transform 1 0 3330 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert82
timestamp 1728341909
transform 1 0 2190 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2_BUFX2_insert83
timestamp 1728341909
transform -1 0 2670 0 -1 7930
box -12 -8 32 252
use FILL  FILL_2_CLKBUF1_insert26
timestamp 1728341909
transform -1 0 1410 0 1 3130
box -12 -8 32 252
use FILL  FILL_2_CLKBUF1_insert27
timestamp 1728341909
transform 1 0 3650 0 1 3130
box -12 -8 32 252
use FILL  FILL_2_CLKBUF1_insert28
timestamp 1728341909
transform 1 0 50 0 1 3130
box -12 -8 32 252
use FILL  FILL_2_CLKBUF1_insert29
timestamp 1728341909
transform 1 0 530 0 1 7930
box -12 -8 32 252
use FILL  FILL_2_CLKBUF1_insert30
timestamp 1728341909
transform 1 0 8210 0 1 5530
box -12 -8 32 252
use FILL  FILL_2_CLKBUF1_insert31
timestamp 1728341909
transform -1 0 7570 0 -1 10810
box -12 -8 32 252
use FILL  FILL_2_CLKBUF1_insert32
timestamp 1728341909
transform -1 0 3190 0 -1 4570
box -12 -8 32 252
use FILL  FILL_2_CLKBUF1_insert33
timestamp 1728341909
transform -1 0 7930 0 1 10330
box -12 -8 32 252
use FILL  FILL_2_CLKBUF1_insert34
timestamp 1728341909
transform -1 0 70 0 -1 11290
box -12 -8 32 252
use FILL  FILL_2_CLKBUF1_insert35
timestamp 1728341909
transform -1 0 5490 0 1 5050
box -12 -8 32 252
use FILL  FILL_2_CLKBUF1_insert36
timestamp 1728341909
transform -1 0 2870 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__1744_
timestamp 1728341909
transform -1 0 4470 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__1745_
timestamp 1728341909
transform 1 0 4250 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__1746_
timestamp 1728341909
transform -1 0 4230 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__1747_
timestamp 1728341909
transform -1 0 5690 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__1748_
timestamp 1728341909
transform 1 0 6610 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__1749_
timestamp 1728341909
transform 1 0 6370 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__1750_
timestamp 1728341909
transform 1 0 5210 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__1751_
timestamp 1728341909
transform 1 0 6850 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__1752_
timestamp 1728341909
transform 1 0 5430 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__1753_
timestamp 1728341909
transform 1 0 7570 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__1754_
timestamp 1728341909
transform -1 0 7110 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__1755_
timestamp 1728341909
transform -1 0 7330 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__1756_
timestamp 1728341909
transform -1 0 6410 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__1757_
timestamp 1728341909
transform 1 0 7070 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__1758_
timestamp 1728341909
transform 1 0 6830 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__1759_
timestamp 1728341909
transform -1 0 3090 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__1760_
timestamp 1728341909
transform 1 0 2390 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__1761_
timestamp 1728341909
transform 1 0 7310 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__1762_
timestamp 1728341909
transform 1 0 2590 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__1763_
timestamp 1728341909
transform -1 0 8230 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__1764_
timestamp 1728341909
transform -1 0 8050 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__1765_
timestamp 1728341909
transform -1 0 8050 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__1766_
timestamp 1728341909
transform -1 0 7850 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__1767_
timestamp 1728341909
transform -1 0 7850 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__1768_
timestamp 1728341909
transform -1 0 5730 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__1769_
timestamp 1728341909
transform 1 0 3170 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__1770_
timestamp 1728341909
transform 1 0 10830 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__1771_
timestamp 1728341909
transform 1 0 11070 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__1772_
timestamp 1728341909
transform 1 0 10810 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__1773_
timestamp 1728341909
transform 1 0 10350 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__1774_
timestamp 1728341909
transform 1 0 10710 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1775_
timestamp 1728341909
transform -1 0 9530 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__1776_
timestamp 1728341909
transform 1 0 9570 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__1777_
timestamp 1728341909
transform -1 0 8750 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__1778_
timestamp 1728341909
transform -1 0 10950 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__1779_
timestamp 1728341909
transform 1 0 10170 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__1780_
timestamp 1728341909
transform 1 0 10930 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__1781_
timestamp 1728341909
transform -1 0 10950 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__1782_
timestamp 1728341909
transform -1 0 11190 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1783_
timestamp 1728341909
transform -1 0 9990 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1784_
timestamp 1728341909
transform 1 0 10570 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__1785_
timestamp 1728341909
transform 1 0 10910 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__1786_
timestamp 1728341909
transform -1 0 10250 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__1787_
timestamp 1728341909
transform 1 0 9250 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__1788_
timestamp 1728341909
transform 1 0 10530 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__1789_
timestamp 1728341909
transform -1 0 9390 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1790_
timestamp 1728341909
transform -1 0 10750 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1791_
timestamp 1728341909
transform 1 0 10970 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1792_
timestamp 1728341909
transform 1 0 5670 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1793_
timestamp 1728341909
transform 1 0 5390 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1794_
timestamp 1728341909
transform -1 0 4970 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1795_
timestamp 1728341909
transform 1 0 3750 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1796_
timestamp 1728341909
transform 1 0 4210 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1797_
timestamp 1728341909
transform -1 0 4730 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1798_
timestamp 1728341909
transform -1 0 11050 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__1799_
timestamp 1728341909
transform -1 0 10950 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__1800_
timestamp 1728341909
transform -1 0 10470 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__1801_
timestamp 1728341909
transform -1 0 10130 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__1802_
timestamp 1728341909
transform 1 0 10010 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__1803_
timestamp 1728341909
transform 1 0 10250 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1804_
timestamp 1728341909
transform 1 0 10250 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__1805_
timestamp 1728341909
transform -1 0 10050 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__1806_
timestamp 1728341909
transform 1 0 9990 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1807_
timestamp 1728341909
transform -1 0 10110 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1808_
timestamp 1728341909
transform -1 0 10410 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__1809_
timestamp 1728341909
transform -1 0 11070 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1810_
timestamp 1728341909
transform -1 0 6250 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1811_
timestamp 1728341909
transform -1 0 11150 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__1812_
timestamp 1728341909
transform -1 0 10230 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__1813_
timestamp 1728341909
transform -1 0 7710 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__1814_
timestamp 1728341909
transform -1 0 7550 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1815_
timestamp 1728341909
transform -1 0 10970 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1816_
timestamp 1728341909
transform -1 0 7610 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__1817_
timestamp 1728341909
transform 1 0 6730 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__1818_
timestamp 1728341909
transform 1 0 6670 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1819_
timestamp 1728341909
transform 1 0 6170 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1820_
timestamp 1728341909
transform 1 0 10370 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__1821_
timestamp 1728341909
transform -1 0 6730 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1822_
timestamp 1728341909
transform 1 0 11150 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__1823_
timestamp 1728341909
transform -1 0 10010 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__1824_
timestamp 1728341909
transform 1 0 7310 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__1825_
timestamp 1728341909
transform 1 0 6530 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1826_
timestamp 1728341909
transform 1 0 10950 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1827_
timestamp 1728341909
transform -1 0 7390 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1828_
timestamp 1728341909
transform 1 0 11150 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__1829_
timestamp 1728341909
transform -1 0 7410 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__1830_
timestamp 1728341909
transform 1 0 7550 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__1831_
timestamp 1728341909
transform 1 0 10690 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__1832_
timestamp 1728341909
transform 1 0 10670 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__1833_
timestamp 1728341909
transform 1 0 7230 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1834_
timestamp 1728341909
transform -1 0 7030 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1835_
timestamp 1728341909
transform -1 0 6470 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1836_
timestamp 1728341909
transform -1 0 6030 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1837_
timestamp 1728341909
transform -1 0 5550 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1838_
timestamp 1728341909
transform 1 0 5270 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1839_
timestamp 1728341909
transform 1 0 5850 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1840_
timestamp 1728341909
transform -1 0 8050 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__1841_
timestamp 1728341909
transform -1 0 4990 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__1842_
timestamp 1728341909
transform -1 0 6850 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__1843_
timestamp 1728341909
transform 1 0 7170 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__1844_
timestamp 1728341909
transform -1 0 10250 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__1845_
timestamp 1728341909
transform 1 0 11150 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__1846_
timestamp 1728341909
transform 1 0 11170 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1847_
timestamp 1728341909
transform -1 0 8090 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__1848_
timestamp 1728341909
transform 1 0 10690 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__1849_
timestamp 1728341909
transform -1 0 10610 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__1850_
timestamp 1728341909
transform -1 0 8550 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__1851_
timestamp 1728341909
transform -1 0 11170 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__1852_
timestamp 1728341909
transform 1 0 9730 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__1853_
timestamp 1728341909
transform 1 0 9250 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__1854_
timestamp 1728341909
transform 1 0 9050 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__1855_
timestamp 1728341909
transform 1 0 8810 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__1856_
timestamp 1728341909
transform 1 0 9330 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__1857_
timestamp 1728341909
transform 1 0 9110 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__1858_
timestamp 1728341909
transform 1 0 7290 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__1859_
timestamp 1728341909
transform -1 0 10710 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__1860_
timestamp 1728341909
transform 1 0 7090 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__1861_
timestamp 1728341909
transform 1 0 7330 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__1862_
timestamp 1728341909
transform -1 0 9830 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__1863_
timestamp 1728341909
transform 1 0 8570 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__1864_
timestamp 1728341909
transform 1 0 9870 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__1865_
timestamp 1728341909
transform 1 0 7730 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__1866_
timestamp 1728341909
transform -1 0 8910 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1867_
timestamp 1728341909
transform 1 0 9290 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__1868_
timestamp 1728341909
transform 1 0 10850 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__1869_
timestamp 1728341909
transform 1 0 9310 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__1870_
timestamp 1728341909
transform -1 0 9090 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__1871_
timestamp 1728341909
transform 1 0 8530 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__1872_
timestamp 1728341909
transform 1 0 7810 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__1873_
timestamp 1728341909
transform 1 0 6370 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1874_
timestamp 1728341909
transform -1 0 6830 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1875_
timestamp 1728341909
transform -1 0 6590 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1876_
timestamp 1728341909
transform 1 0 6650 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__1877_
timestamp 1728341909
transform -1 0 8070 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__1878_
timestamp 1728341909
transform -1 0 8330 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__1879_
timestamp 1728341909
transform -1 0 8070 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__1880_
timestamp 1728341909
transform -1 0 7010 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__1881_
timestamp 1728341909
transform -1 0 6330 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__1882_
timestamp 1728341909
transform 1 0 3490 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__1883_
timestamp 1728341909
transform -1 0 7030 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__1884_
timestamp 1728341909
transform -1 0 6550 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__1885_
timestamp 1728341909
transform 1 0 5830 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__1886_
timestamp 1728341909
transform -1 0 6230 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__1887_
timestamp 1728341909
transform 1 0 6850 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__1888_
timestamp 1728341909
transform 1 0 3610 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__1889_
timestamp 1728341909
transform -1 0 5970 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__1890_
timestamp 1728341909
transform 1 0 6430 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__1891_
timestamp 1728341909
transform -1 0 6070 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__1892_
timestamp 1728341909
transform 1 0 5630 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__1893_
timestamp 1728341909
transform 1 0 1030 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__1894_
timestamp 1728341909
transform 1 0 5970 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__1895_
timestamp 1728341909
transform 1 0 6850 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__1896_
timestamp 1728341909
transform 1 0 5170 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__1897_
timestamp 1728341909
transform 1 0 6010 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__1898_
timestamp 1728341909
transform 1 0 6430 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__1899_
timestamp 1728341909
transform 1 0 6530 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__1900_
timestamp 1728341909
transform 1 0 550 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__1901_
timestamp 1728341909
transform 1 0 7990 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__1902_
timestamp 1728341909
transform 1 0 8530 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__1903_
timestamp 1728341909
transform 1 0 7890 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__1904_
timestamp 1728341909
transform -1 0 10050 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1905_
timestamp 1728341909
transform 1 0 7550 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__1906_
timestamp 1728341909
transform 1 0 7530 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__1907_
timestamp 1728341909
transform 1 0 8670 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1908_
timestamp 1728341909
transform -1 0 7730 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1909_
timestamp 1728341909
transform 1 0 1830 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1910_
timestamp 1728341909
transform -1 0 9790 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__1911_
timestamp 1728341909
transform 1 0 9510 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1912_
timestamp 1728341909
transform 1 0 6130 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1913_
timestamp 1728341909
transform 1 0 10650 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__1914_
timestamp 1728341909
transform 1 0 10710 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1915_
timestamp 1728341909
transform -1 0 10270 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1916_
timestamp 1728341909
transform -1 0 5890 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1917_
timestamp 1728341909
transform 1 0 4030 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1918_
timestamp 1728341909
transform -1 0 810 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__1919_
timestamp 1728341909
transform -1 0 90 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__1920_
timestamp 1728341909
transform 1 0 1030 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__1921_
timestamp 1728341909
transform -1 0 1210 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1922_
timestamp 1728341909
transform -1 0 950 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1923_
timestamp 1728341909
transform 1 0 550 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__1924_
timestamp 1728341909
transform -1 0 4490 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1925_
timestamp 1728341909
transform -1 0 330 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__1926_
timestamp 1728341909
transform 1 0 790 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__1927_
timestamp 1728341909
transform -1 0 2090 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1928_
timestamp 1728341909
transform -1 0 1610 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1929_
timestamp 1728341909
transform 1 0 290 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__1930_
timestamp 1728341909
transform 1 0 670 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1931_
timestamp 1728341909
transform 1 0 550 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__1932_
timestamp 1728341909
transform -1 0 570 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1933_
timestamp 1728341909
transform 1 0 550 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__1934_
timestamp 1728341909
transform -1 0 570 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1935_
timestamp 1728341909
transform -1 0 1550 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1936_
timestamp 1728341909
transform 1 0 810 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1937_
timestamp 1728341909
transform -1 0 570 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__1938_
timestamp 1728341909
transform -1 0 90 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__1939_
timestamp 1728341909
transform 1 0 310 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__1940_
timestamp 1728341909
transform 1 0 830 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1941_
timestamp 1728341909
transform 1 0 550 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__1942_
timestamp 1728341909
transform 1 0 550 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__1943_
timestamp 1728341909
transform 1 0 8110 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__1944_
timestamp 1728341909
transform -1 0 7650 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1945_
timestamp 1728341909
transform -1 0 7430 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1946_
timestamp 1728341909
transform 1 0 8450 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1947_
timestamp 1728341909
transform -1 0 7630 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1948_
timestamp 1728341909
transform -1 0 6970 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1949_
timestamp 1728341909
transform -1 0 7210 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1950_
timestamp 1728341909
transform 1 0 8310 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__1951_
timestamp 1728341909
transform 1 0 8310 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__1952_
timestamp 1728341909
transform 1 0 9830 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1953_
timestamp 1728341909
transform -1 0 8390 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__1954_
timestamp 1728341909
transform 1 0 8230 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1955_
timestamp 1728341909
transform 1 0 6430 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__1956_
timestamp 1728341909
transform -1 0 7990 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1957_
timestamp 1728341909
transform 1 0 8070 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__1958_
timestamp 1728341909
transform 1 0 10430 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__1959_
timestamp 1728341909
transform 1 0 7790 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__1960_
timestamp 1728341909
transform 1 0 7870 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__1961_
timestamp 1728341909
transform 1 0 10690 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__1962_
timestamp 1728341909
transform 1 0 10490 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__1963_
timestamp 1728341909
transform 1 0 9830 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1964_
timestamp 1728341909
transform -1 0 7370 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__1965_
timestamp 1728341909
transform -1 0 7650 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__1966_
timestamp 1728341909
transform -1 0 3510 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__1967_
timestamp 1728341909
transform -1 0 6970 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__1968_
timestamp 1728341909
transform 1 0 7510 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__1969_
timestamp 1728341909
transform -1 0 7770 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__1970_
timestamp 1728341909
transform 1 0 1510 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__1971_
timestamp 1728341909
transform -1 0 810 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1972_
timestamp 1728341909
transform 1 0 1330 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1973_
timestamp 1728341909
transform 1 0 1590 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__1974_
timestamp 1728341909
transform 1 0 8350 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__1975_
timestamp 1728341909
transform 1 0 2970 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__1976_
timestamp 1728341909
transform -1 0 7130 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__1977_
timestamp 1728341909
transform -1 0 2830 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__1978_
timestamp 1728341909
transform -1 0 3810 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__1979_
timestamp 1728341909
transform -1 0 6510 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__1980_
timestamp 1728341909
transform 1 0 7770 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__1981_
timestamp 1728341909
transform 1 0 8290 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__1982_
timestamp 1728341909
transform -1 0 3030 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__1983_
timestamp 1728341909
transform 1 0 1710 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__1984_
timestamp 1728341909
transform 1 0 1790 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__1985_
timestamp 1728341909
transform 1 0 2450 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__1986_
timestamp 1728341909
transform -1 0 7130 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__1987_
timestamp 1728341909
transform 1 0 5070 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__1988_
timestamp 1728341909
transform -1 0 4970 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__1989_
timestamp 1728341909
transform 1 0 6730 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__1990_
timestamp 1728341909
transform -1 0 7250 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__1991_
timestamp 1728341909
transform -1 0 2050 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__1992_
timestamp 1728341909
transform -1 0 1550 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__1993_
timestamp 1728341909
transform -1 0 1830 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__1994_
timestamp 1728341909
transform 1 0 2070 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__1995_
timestamp 1728341909
transform 1 0 8030 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__1996_
timestamp 1728341909
transform -1 0 2250 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__1997_
timestamp 1728341909
transform -1 0 3970 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__1998_
timestamp 1728341909
transform -1 0 6490 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__1999_
timestamp 1728341909
transform -1 0 8210 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2000_
timestamp 1728341909
transform 1 0 1810 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2001_
timestamp 1728341909
transform 1 0 1290 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2002_
timestamp 1728341909
transform 1 0 1530 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2003_
timestamp 1728341909
transform 1 0 1550 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2004_
timestamp 1728341909
transform 1 0 7830 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2005_
timestamp 1728341909
transform 1 0 1990 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2006_
timestamp 1728341909
transform -1 0 6250 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2007_
timestamp 1728341909
transform 1 0 7530 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2008_
timestamp 1728341909
transform -1 0 8050 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2009_
timestamp 1728341909
transform 1 0 790 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2010_
timestamp 1728341909
transform -1 0 850 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2011_
timestamp 1728341909
transform 1 0 550 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2012_
timestamp 1728341909
transform 1 0 810 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2013_
timestamp 1728341909
transform 1 0 5450 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2014_
timestamp 1728341909
transform 1 0 1750 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2015_
timestamp 1728341909
transform -1 0 3950 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2016_
timestamp 1728341909
transform 1 0 6750 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2017_
timestamp 1728341909
transform -1 0 7290 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2018_
timestamp 1728341909
transform -1 0 1530 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2019_
timestamp 1728341909
transform -1 0 1590 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2020_
timestamp 1728341909
transform 1 0 1770 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2021_
timestamp 1728341909
transform 1 0 1730 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2022_
timestamp 1728341909
transform 1 0 4510 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2023_
timestamp 1728341909
transform 1 0 550 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2024_
timestamp 1728341909
transform 1 0 1450 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2025_
timestamp 1728341909
transform 1 0 2510 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2026_
timestamp 1728341909
transform -1 0 4710 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2027_
timestamp 1728341909
transform 1 0 7210 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2028_
timestamp 1728341909
transform -1 0 7490 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2029_
timestamp 1728341909
transform -1 0 90 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2030_
timestamp 1728341909
transform -1 0 570 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2031_
timestamp 1728341909
transform -1 0 330 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2032_
timestamp 1728341909
transform 1 0 550 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2033_
timestamp 1728341909
transform 1 0 7630 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2034_
timestamp 1728341909
transform 1 0 1230 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2035_
timestamp 1728341909
transform 1 0 2110 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2036_
timestamp 1728341909
transform 1 0 2910 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2037_
timestamp 1728341909
transform -1 0 4110 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2038_
timestamp 1728341909
transform 1 0 7550 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2039_
timestamp 1728341909
transform -1 0 7830 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2040_
timestamp 1728341909
transform -1 0 2950 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2041_
timestamp 1728341909
transform -1 0 570 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2042_
timestamp 1728341909
transform 1 0 1730 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__2043_
timestamp 1728341909
transform -1 0 3830 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__2044_
timestamp 1728341909
transform 1 0 5370 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2045_
timestamp 1728341909
transform -1 0 4070 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2046_
timestamp 1728341909
transform 1 0 2870 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__2047_
timestamp 1728341909
transform 1 0 2630 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__2048_
timestamp 1728341909
transform -1 0 3570 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__2049_
timestamp 1728341909
transform -1 0 2970 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__2050_
timestamp 1728341909
transform -1 0 2450 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__2051_
timestamp 1728341909
transform -1 0 2430 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2052_
timestamp 1728341909
transform -1 0 850 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2053_
timestamp 1728341909
transform -1 0 3410 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__2054_
timestamp 1728341909
transform 1 0 3130 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__2055_
timestamp 1728341909
transform -1 0 2770 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__2056_
timestamp 1728341909
transform 1 0 4390 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2057_
timestamp 1728341909
transform -1 0 3950 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2058_
timestamp 1728341909
transform 1 0 4610 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2059_
timestamp 1728341909
transform -1 0 1970 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__2060_
timestamp 1728341909
transform -1 0 3790 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__2061_
timestamp 1728341909
transform 1 0 3530 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__2062_
timestamp 1728341909
transform -1 0 3550 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__2063_
timestamp 1728341909
transform 1 0 2490 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__2064_
timestamp 1728341909
transform -1 0 2590 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2065_
timestamp 1728341909
transform -1 0 2390 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2066_
timestamp 1728341909
transform 1 0 2450 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2067_
timestamp 1728341909
transform -1 0 2770 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__2068_
timestamp 1728341909
transform -1 0 3010 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__2069_
timestamp 1728341909
transform 1 0 2550 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__2070_
timestamp 1728341909
transform -1 0 1090 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2071_
timestamp 1728341909
transform -1 0 2810 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__2072_
timestamp 1728341909
transform -1 0 2550 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__2073_
timestamp 1728341909
transform -1 0 1290 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2074_
timestamp 1728341909
transform 1 0 3230 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__2075_
timestamp 1728341909
transform -1 0 2710 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__2076_
timestamp 1728341909
transform 1 0 2410 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__2077_
timestamp 1728341909
transform -1 0 3270 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__2078_
timestamp 1728341909
transform 1 0 2790 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__2079_
timestamp 1728341909
transform -1 0 3910 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2080_
timestamp 1728341909
transform 1 0 4130 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2081_
timestamp 1728341909
transform -1 0 3690 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2082_
timestamp 1728341909
transform 1 0 5770 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2083_
timestamp 1728341909
transform -1 0 6510 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2084_
timestamp 1728341909
transform 1 0 9930 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2085_
timestamp 1728341909
transform -1 0 10450 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2086_
timestamp 1728341909
transform 1 0 10470 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2087_
timestamp 1728341909
transform 1 0 11010 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__2088_
timestamp 1728341909
transform 1 0 10210 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2089_
timestamp 1728341909
transform -1 0 9510 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2090_
timestamp 1728341909
transform 1 0 10690 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__2091_
timestamp 1728341909
transform 1 0 11190 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__2092_
timestamp 1728341909
transform -1 0 10150 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2093_
timestamp 1728341909
transform 1 0 10210 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__2094_
timestamp 1728341909
transform -1 0 10710 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__2095_
timestamp 1728341909
transform 1 0 10770 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__2096_
timestamp 1728341909
transform -1 0 11170 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__2097_
timestamp 1728341909
transform -1 0 11110 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2098_
timestamp 1728341909
transform 1 0 10190 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2099_
timestamp 1728341909
transform 1 0 10670 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2100_
timestamp 1728341909
transform 1 0 10890 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2101_
timestamp 1728341909
transform 1 0 11130 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2102_
timestamp 1728341909
transform 1 0 4010 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__2103_
timestamp 1728341909
transform 1 0 4250 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__2104_
timestamp 1728341909
transform 1 0 3870 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2105_
timestamp 1728341909
transform -1 0 1770 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2106_
timestamp 1728341909
transform -1 0 2150 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2107_
timestamp 1728341909
transform -1 0 2670 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2108_
timestamp 1728341909
transform 1 0 1470 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2109_
timestamp 1728341909
transform -1 0 2890 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2110_
timestamp 1728341909
transform 1 0 3110 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2111_
timestamp 1728341909
transform 1 0 5310 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2112_
timestamp 1728341909
transform 1 0 11190 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__2113_
timestamp 1728341909
transform -1 0 9770 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__2114_
timestamp 1728341909
transform 1 0 9770 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2115_
timestamp 1728341909
transform -1 0 11090 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2116_
timestamp 1728341909
transform -1 0 11030 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__2117_
timestamp 1728341909
transform -1 0 10630 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__2118_
timestamp 1728341909
transform 1 0 9030 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__2119_
timestamp 1728341909
transform -1 0 11110 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__2120_
timestamp 1728341909
transform 1 0 11050 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2121_
timestamp 1728341909
transform 1 0 11150 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2122_
timestamp 1728341909
transform 1 0 10850 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2123_
timestamp 1728341909
transform 1 0 10910 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2124_
timestamp 1728341909
transform 1 0 9370 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2125_
timestamp 1728341909
transform 1 0 9490 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2126_
timestamp 1728341909
transform -1 0 9930 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2127_
timestamp 1728341909
transform 1 0 9750 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2128_
timestamp 1728341909
transform 1 0 9710 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2129_
timestamp 1728341909
transform -1 0 8930 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2130_
timestamp 1728341909
transform 1 0 9610 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2131_
timestamp 1728341909
transform 1 0 9710 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2132_
timestamp 1728341909
transform 1 0 10170 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2133_
timestamp 1728341909
transform 1 0 10330 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2134_
timestamp 1728341909
transform -1 0 10110 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2135_
timestamp 1728341909
transform 1 0 10610 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2136_
timestamp 1728341909
transform -1 0 10570 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2137_
timestamp 1728341909
transform 1 0 10810 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2138_
timestamp 1728341909
transform -1 0 10910 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2139_
timestamp 1728341909
transform -1 0 10850 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2140_
timestamp 1728341909
transform -1 0 8330 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2141_
timestamp 1728341909
transform 1 0 8570 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2142_
timestamp 1728341909
transform 1 0 1890 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2143_
timestamp 1728341909
transform -1 0 2930 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2144_
timestamp 1728341909
transform -1 0 6030 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2145_
timestamp 1728341909
transform -1 0 6230 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2146_
timestamp 1728341909
transform 1 0 5530 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2147_
timestamp 1728341909
transform -1 0 6770 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2148_
timestamp 1728341909
transform 1 0 9670 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2149_
timestamp 1728341909
transform 1 0 8750 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2150_
timestamp 1728341909
transform -1 0 8510 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2151_
timestamp 1728341909
transform 1 0 8170 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2152_
timestamp 1728341909
transform -1 0 9010 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2153_
timestamp 1728341909
transform -1 0 9110 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2154_
timestamp 1728341909
transform 1 0 8850 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__2155_
timestamp 1728341909
transform 1 0 8010 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__2156_
timestamp 1728341909
transform -1 0 8290 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__2157_
timestamp 1728341909
transform -1 0 8410 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2158_
timestamp 1728341909
transform 1 0 10330 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__2159_
timestamp 1728341909
transform 1 0 6030 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2160_
timestamp 1728341909
transform -1 0 6390 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2161_
timestamp 1728341909
transform 1 0 6590 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2162_
timestamp 1728341909
transform -1 0 7930 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2163_
timestamp 1728341909
transform -1 0 8350 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__2164_
timestamp 1728341909
transform 1 0 7110 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2165_
timestamp 1728341909
transform -1 0 7090 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2166_
timestamp 1728341909
transform -1 0 8150 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2167_
timestamp 1728341909
transform -1 0 7850 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2168_
timestamp 1728341909
transform -1 0 8110 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2169_
timestamp 1728341909
transform 1 0 8150 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2170_
timestamp 1728341909
transform -1 0 8370 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2171_
timestamp 1728341909
transform 1 0 8570 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2172_
timestamp 1728341909
transform -1 0 10430 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2173_
timestamp 1728341909
transform 1 0 10170 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2174_
timestamp 1728341909
transform 1 0 4390 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2175_
timestamp 1728341909
transform -1 0 3950 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2176_
timestamp 1728341909
transform -1 0 5410 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2177_
timestamp 1728341909
transform -1 0 6070 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2178_
timestamp 1728341909
transform -1 0 6330 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2179_
timestamp 1728341909
transform 1 0 6370 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2180_
timestamp 1728341909
transform 1 0 7170 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2181_
timestamp 1728341909
transform 1 0 7310 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__2182_
timestamp 1728341909
transform -1 0 7170 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__2183_
timestamp 1728341909
transform 1 0 6150 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2184_
timestamp 1728341909
transform 1 0 6470 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2185_
timestamp 1728341909
transform -1 0 6610 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2186_
timestamp 1728341909
transform -1 0 9050 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2187_
timestamp 1728341909
transform -1 0 9450 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2188_
timestamp 1728341909
transform 1 0 9050 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2189_
timestamp 1728341909
transform -1 0 8830 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2190_
timestamp 1728341909
transform 1 0 8510 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2191_
timestamp 1728341909
transform 1 0 8750 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2192_
timestamp 1728341909
transform 1 0 7310 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2193_
timestamp 1728341909
transform 1 0 7530 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2194_
timestamp 1728341909
transform -1 0 8650 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__2195_
timestamp 1728341909
transform -1 0 8570 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__2196_
timestamp 1728341909
transform 1 0 8610 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2197_
timestamp 1728341909
transform 1 0 8650 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2198_
timestamp 1728341909
transform -1 0 7250 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2199_
timestamp 1728341909
transform -1 0 7510 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2200_
timestamp 1728341909
transform 1 0 9030 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__2201_
timestamp 1728341909
transform 1 0 8890 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2202_
timestamp 1728341909
transform -1 0 8690 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2203_
timestamp 1728341909
transform 1 0 8410 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2204_
timestamp 1728341909
transform -1 0 8410 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2205_
timestamp 1728341909
transform 1 0 8150 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2206_
timestamp 1728341909
transform -1 0 8030 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2207_
timestamp 1728341909
transform 1 0 8530 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2208_
timestamp 1728341909
transform -1 0 8290 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2209_
timestamp 1728341909
transform -1 0 7810 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2210_
timestamp 1728341909
transform 1 0 2750 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2211_
timestamp 1728341909
transform -1 0 7210 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2212_
timestamp 1728341909
transform -1 0 7470 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2213_
timestamp 1728341909
transform -1 0 7990 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2214_
timestamp 1728341909
transform 1 0 8550 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2215_
timestamp 1728341909
transform 1 0 9250 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2216_
timestamp 1728341909
transform 1 0 9230 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2217_
timestamp 1728341909
transform -1 0 9490 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2218_
timestamp 1728341909
transform 1 0 3930 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2219_
timestamp 1728341909
transform -1 0 2250 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__2220_
timestamp 1728341909
transform -1 0 3670 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2221_
timestamp 1728341909
transform 1 0 4110 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2222_
timestamp 1728341909
transform 1 0 4330 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2223_
timestamp 1728341909
transform 1 0 4150 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2224_
timestamp 1728341909
transform -1 0 2830 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2225_
timestamp 1728341909
transform -1 0 5890 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2226_
timestamp 1728341909
transform 1 0 6010 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2227_
timestamp 1728341909
transform -1 0 6990 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2228_
timestamp 1728341909
transform 1 0 6730 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2229_
timestamp 1728341909
transform 1 0 7790 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__2230_
timestamp 1728341909
transform -1 0 6190 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__2231_
timestamp 1728341909
transform -1 0 6430 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__2232_
timestamp 1728341909
transform 1 0 6850 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2233_
timestamp 1728341909
transform 1 0 7430 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2234_
timestamp 1728341909
transform 1 0 7330 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2235_
timestamp 1728341909
transform 1 0 9410 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2236_
timestamp 1728341909
transform 1 0 10470 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2237_
timestamp 1728341909
transform 1 0 9950 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2238_
timestamp 1728341909
transform -1 0 9870 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2239_
timestamp 1728341909
transform -1 0 5830 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2240_
timestamp 1728341909
transform 1 0 2690 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2241_
timestamp 1728341909
transform -1 0 4370 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2242_
timestamp 1728341909
transform -1 0 4590 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2243_
timestamp 1728341909
transform 1 0 3370 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2244_
timestamp 1728341909
transform 1 0 5130 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2245_
timestamp 1728341909
transform 1 0 7270 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2246_
timestamp 1728341909
transform 1 0 7290 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2247_
timestamp 1728341909
transform -1 0 3250 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2248_
timestamp 1728341909
transform 1 0 3430 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2249_
timestamp 1728341909
transform 1 0 5410 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2250_
timestamp 1728341909
transform 1 0 6670 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2251_
timestamp 1728341909
transform 1 0 7190 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2252_
timestamp 1728341909
transform -1 0 9630 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__2253_
timestamp 1728341909
transform 1 0 9350 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2254_
timestamp 1728341909
transform 1 0 5630 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2255_
timestamp 1728341909
transform -1 0 6970 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2256_
timestamp 1728341909
transform 1 0 7130 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2257_
timestamp 1728341909
transform -1 0 3070 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2258_
timestamp 1728341909
transform -1 0 3030 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__2259_
timestamp 1728341909
transform 1 0 3450 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2260_
timestamp 1728341909
transform 1 0 4630 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2261_
timestamp 1728341909
transform -1 0 5630 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2262_
timestamp 1728341909
transform 1 0 4810 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2263_
timestamp 1728341909
transform 1 0 4870 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2264_
timestamp 1728341909
transform -1 0 6170 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2265_
timestamp 1728341909
transform 1 0 3470 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__2266_
timestamp 1728341909
transform 1 0 7510 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__2267_
timestamp 1728341909
transform -1 0 5410 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__2268_
timestamp 1728341909
transform -1 0 5650 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__2269_
timestamp 1728341909
transform 1 0 5410 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__2270_
timestamp 1728341909
transform -1 0 6250 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__2271_
timestamp 1728341909
transform 1 0 5970 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__2272_
timestamp 1728341909
transform 1 0 5570 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__2273_
timestamp 1728341909
transform 1 0 5390 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__2274_
timestamp 1728341909
transform 1 0 5150 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__2275_
timestamp 1728341909
transform 1 0 5630 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__2276_
timestamp 1728341909
transform -1 0 6270 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2277_
timestamp 1728341909
transform 1 0 7770 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__2278_
timestamp 1728341909
transform -1 0 7710 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2279_
timestamp 1728341909
transform 1 0 6470 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2280_
timestamp 1728341909
transform -1 0 6490 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2281_
timestamp 1728341909
transform -1 0 6250 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2282_
timestamp 1728341909
transform 1 0 6530 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2283_
timestamp 1728341909
transform 1 0 7230 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2284_
timestamp 1728341909
transform 1 0 9190 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2285_
timestamp 1728341909
transform 1 0 9630 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2286_
timestamp 1728341909
transform -1 0 2530 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__2287_
timestamp 1728341909
transform -1 0 1790 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2288_
timestamp 1728341909
transform -1 0 2230 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2289_
timestamp 1728341909
transform 1 0 2190 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2290_
timestamp 1728341909
transform -1 0 1750 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2291_
timestamp 1728341909
transform 1 0 1970 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2292_
timestamp 1728341909
transform 1 0 4090 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2293_
timestamp 1728341909
transform 1 0 4830 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2294_
timestamp 1728341909
transform 1 0 6050 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2295_
timestamp 1728341909
transform -1 0 2230 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2296_
timestamp 1728341909
transform 1 0 3670 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2297_
timestamp 1728341909
transform 1 0 2210 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2298_
timestamp 1728341909
transform 1 0 1970 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2299_
timestamp 1728341909
transform 1 0 3430 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2300_
timestamp 1728341909
transform 1 0 3170 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2301_
timestamp 1728341909
transform -1 0 3630 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2302_
timestamp 1728341909
transform 1 0 5110 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2303_
timestamp 1728341909
transform -1 0 5090 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2304_
timestamp 1728341909
transform 1 0 5330 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2305_
timestamp 1728341909
transform -1 0 1530 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2306_
timestamp 1728341909
transform 1 0 2430 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2307_
timestamp 1728341909
transform -1 0 5590 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2308_
timestamp 1728341909
transform -1 0 5590 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2309_
timestamp 1728341909
transform 1 0 4590 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2310_
timestamp 1728341909
transform 1 0 4350 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2311_
timestamp 1728341909
transform -1 0 3750 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2312_
timestamp 1728341909
transform -1 0 3990 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2313_
timestamp 1728341909
transform 1 0 5270 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2314_
timestamp 1728341909
transform 1 0 4450 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2315_
timestamp 1728341909
transform 1 0 5410 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2316_
timestamp 1728341909
transform -1 0 9850 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2317_
timestamp 1728341909
transform 1 0 11150 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2318_
timestamp 1728341909
transform -1 0 10850 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__2319_
timestamp 1728341909
transform -1 0 10470 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__2320_
timestamp 1728341909
transform 1 0 10630 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2321_
timestamp 1728341909
transform 1 0 10570 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__2322_
timestamp 1728341909
transform 1 0 10470 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__2323_
timestamp 1728341909
transform 1 0 6730 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2324_
timestamp 1728341909
transform 1 0 6930 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2325_
timestamp 1728341909
transform 1 0 9290 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2326_
timestamp 1728341909
transform -1 0 8830 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2327_
timestamp 1728341909
transform -1 0 9290 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2328_
timestamp 1728341909
transform -1 0 9530 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2329_
timestamp 1728341909
transform 1 0 9250 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2330_
timestamp 1728341909
transform -1 0 9010 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2331_
timestamp 1728341909
transform -1 0 9170 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2332_
timestamp 1728341909
transform 1 0 9150 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2333_
timestamp 1728341909
transform 1 0 9410 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2334_
timestamp 1728341909
transform -1 0 9610 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2335_
timestamp 1728341909
transform 1 0 5650 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2336_
timestamp 1728341909
transform 1 0 6170 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2337_
timestamp 1728341909
transform -1 0 5950 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2338_
timestamp 1728341909
transform -1 0 5890 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2339_
timestamp 1728341909
transform 1 0 10370 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2340_
timestamp 1728341909
transform -1 0 9250 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2341_
timestamp 1728341909
transform 1 0 9250 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2342_
timestamp 1728341909
transform 1 0 10110 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2343_
timestamp 1728341909
transform -1 0 9610 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2344_
timestamp 1728341909
transform 1 0 9710 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2345_
timestamp 1728341909
transform -1 0 6890 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2346_
timestamp 1728341909
transform 1 0 6750 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2347_
timestamp 1728341909
transform -1 0 7090 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2348_
timestamp 1728341909
transform 1 0 8090 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2349_
timestamp 1728341909
transform -1 0 7790 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2350_
timestamp 1728341909
transform 1 0 7510 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2351_
timestamp 1728341909
transform -1 0 5210 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2352_
timestamp 1728341909
transform 1 0 5810 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2353_
timestamp 1728341909
transform -1 0 4230 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2354_
timestamp 1728341909
transform 1 0 4710 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2355_
timestamp 1728341909
transform -1 0 4970 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2356_
timestamp 1728341909
transform 1 0 5910 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2357_
timestamp 1728341909
transform -1 0 5670 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2358_
timestamp 1728341909
transform 1 0 6950 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2359_
timestamp 1728341909
transform 1 0 6310 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2360_
timestamp 1728341909
transform 1 0 6550 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2361_
timestamp 1728341909
transform 1 0 7850 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__2362_
timestamp 1728341909
transform 1 0 7370 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2363_
timestamp 1728341909
transform -1 0 7470 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2364_
timestamp 1728341909
transform 1 0 8090 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__2365_
timestamp 1728341909
transform -1 0 7970 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2366_
timestamp 1728341909
transform 1 0 7730 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2367_
timestamp 1728341909
transform 1 0 8010 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2368_
timestamp 1728341909
transform 1 0 8230 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2369_
timestamp 1728341909
transform -1 0 9950 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2370_
timestamp 1728341909
transform 1 0 5370 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2371_
timestamp 1728341909
transform -1 0 8770 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2372_
timestamp 1728341909
transform -1 0 8510 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2373_
timestamp 1728341909
transform -1 0 8090 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2374_
timestamp 1728341909
transform 1 0 8090 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2375_
timestamp 1728341909
transform 1 0 6490 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2376_
timestamp 1728341909
transform 1 0 8450 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2377_
timestamp 1728341909
transform -1 0 8710 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2378_
timestamp 1728341909
transform -1 0 9010 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2379_
timestamp 1728341909
transform -1 0 6870 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2380_
timestamp 1728341909
transform -1 0 7010 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2381_
timestamp 1728341909
transform -1 0 6870 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2382_
timestamp 1728341909
transform -1 0 7950 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2383_
timestamp 1728341909
transform 1 0 7670 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2384_
timestamp 1728341909
transform 1 0 7770 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2385_
timestamp 1728341909
transform -1 0 7510 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2386_
timestamp 1728341909
transform -1 0 6630 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2387_
timestamp 1728341909
transform -1 0 6390 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2388_
timestamp 1728341909
transform -1 0 8950 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2389_
timestamp 1728341909
transform -1 0 8330 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2390_
timestamp 1728341909
transform -1 0 8270 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2391_
timestamp 1728341909
transform -1 0 9510 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2392_
timestamp 1728341909
transform 1 0 8270 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2393_
timestamp 1728341909
transform 1 0 8230 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2394_
timestamp 1728341909
transform 1 0 8870 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2395_
timestamp 1728341909
transform 1 0 8830 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2396_
timestamp 1728341909
transform 1 0 9110 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2397_
timestamp 1728341909
transform -1 0 9370 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2398_
timestamp 1728341909
transform 1 0 8750 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2399_
timestamp 1728341909
transform -1 0 7630 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2400_
timestamp 1728341909
transform 1 0 7370 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2401_
timestamp 1728341909
transform 1 0 8490 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2402_
timestamp 1728341909
transform -1 0 6430 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2403_
timestamp 1728341909
transform -1 0 6630 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2404_
timestamp 1728341909
transform -1 0 7590 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2405_
timestamp 1728341909
transform -1 0 7370 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2406_
timestamp 1728341909
transform 1 0 7090 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2407_
timestamp 1728341909
transform -1 0 6630 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2408_
timestamp 1728341909
transform -1 0 5930 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2409_
timestamp 1728341909
transform 1 0 7010 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2410_
timestamp 1728341909
transform -1 0 7290 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2411_
timestamp 1728341909
transform -1 0 6850 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2412_
timestamp 1728341909
transform -1 0 7510 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2413_
timestamp 1728341909
transform 1 0 7030 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2414_
timestamp 1728341909
transform 1 0 6850 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2415_
timestamp 1728341909
transform -1 0 8050 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2416_
timestamp 1728341909
transform 1 0 7790 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2417_
timestamp 1728341909
transform -1 0 9030 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2418_
timestamp 1728341909
transform -1 0 8810 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2419_
timestamp 1728341909
transform 1 0 7070 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2420_
timestamp 1728341909
transform 1 0 2230 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2421_
timestamp 1728341909
transform -1 0 9690 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2422_
timestamp 1728341909
transform 1 0 8270 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__2423_
timestamp 1728341909
transform 1 0 8990 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2424_
timestamp 1728341909
transform 1 0 8770 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2425_
timestamp 1728341909
transform 1 0 3170 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2426_
timestamp 1728341909
transform 1 0 8750 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2427_
timestamp 1728341909
transform 1 0 8830 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__2428_
timestamp 1728341909
transform 1 0 9230 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2429_
timestamp 1728341909
transform 1 0 9450 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2430_
timestamp 1728341909
transform 1 0 8810 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2431_
timestamp 1728341909
transform -1 0 9270 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2432_
timestamp 1728341909
transform 1 0 9490 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2433_
timestamp 1728341909
transform -1 0 9910 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2434_
timestamp 1728341909
transform -1 0 9990 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2435_
timestamp 1728341909
transform 1 0 4450 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__2436_
timestamp 1728341909
transform 1 0 9210 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2437_
timestamp 1728341909
transform 1 0 10890 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__2438_
timestamp 1728341909
transform -1 0 10950 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__2439_
timestamp 1728341909
transform -1 0 10930 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__2440_
timestamp 1728341909
transform 1 0 9050 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__2441_
timestamp 1728341909
transform -1 0 6190 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__2442_
timestamp 1728341909
transform -1 0 8270 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2443_
timestamp 1728341909
transform 1 0 3830 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2444_
timestamp 1728341909
transform -1 0 4710 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__2445_
timestamp 1728341909
transform -1 0 8610 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__2446_
timestamp 1728341909
transform 1 0 8250 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2447_
timestamp 1728341909
transform 1 0 8090 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2448_
timestamp 1728341909
transform 1 0 8490 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2449_
timestamp 1728341909
transform -1 0 8770 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2450_
timestamp 1728341909
transform -1 0 8970 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2451_
timestamp 1728341909
transform 1 0 3830 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2452_
timestamp 1728341909
transform 1 0 7610 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2453_
timestamp 1728341909
transform -1 0 6630 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2454_
timestamp 1728341909
transform -1 0 6350 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2455_
timestamp 1728341909
transform -1 0 6630 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2456_
timestamp 1728341909
transform -1 0 8750 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2457_
timestamp 1728341909
transform -1 0 8970 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2458_
timestamp 1728341909
transform -1 0 6810 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2459_
timestamp 1728341909
transform -1 0 3590 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2460_
timestamp 1728341909
transform 1 0 7110 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2461_
timestamp 1728341909
transform 1 0 7030 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2462_
timestamp 1728341909
transform -1 0 7310 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2463_
timestamp 1728341909
transform -1 0 7330 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2464_
timestamp 1728341909
transform 1 0 4490 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__2465_
timestamp 1728341909
transform -1 0 7390 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2466_
timestamp 1728341909
transform -1 0 3370 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2467_
timestamp 1728341909
transform 1 0 6190 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2468_
timestamp 1728341909
transform -1 0 6310 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2469_
timestamp 1728341909
transform -1 0 6150 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2470_
timestamp 1728341909
transform -1 0 6410 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2471_
timestamp 1728341909
transform -1 0 8070 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2472_
timestamp 1728341909
transform -1 0 6090 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2473_
timestamp 1728341909
transform -1 0 5430 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2474_
timestamp 1728341909
transform -1 0 5350 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2475_
timestamp 1728341909
transform -1 0 7810 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__2476_
timestamp 1728341909
transform -1 0 2730 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2477_
timestamp 1728341909
transform -1 0 5210 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2478_
timestamp 1728341909
transform 1 0 5290 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2479_
timestamp 1728341909
transform -1 0 8030 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2480_
timestamp 1728341909
transform 1 0 5930 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2481_
timestamp 1728341909
transform 1 0 4190 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2482_
timestamp 1728341909
transform -1 0 2470 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2483_
timestamp 1728341909
transform -1 0 4710 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2484_
timestamp 1728341909
transform -1 0 5750 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2485_
timestamp 1728341909
transform -1 0 6990 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2486_
timestamp 1728341909
transform 1 0 3110 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2487_
timestamp 1728341909
transform -1 0 5690 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2488_
timestamp 1728341909
transform 1 0 6450 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2489_
timestamp 1728341909
transform -1 0 6730 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2490_
timestamp 1728341909
transform 1 0 7710 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2491_
timestamp 1728341909
transform -1 0 7950 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2492_
timestamp 1728341909
transform -1 0 2890 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2493_
timestamp 1728341909
transform -1 0 5530 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2494_
timestamp 1728341909
transform -1 0 6610 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2495_
timestamp 1728341909
transform 1 0 6850 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2496_
timestamp 1728341909
transform 1 0 7570 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2497_
timestamp 1728341909
transform -1 0 7810 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2498_
timestamp 1728341909
transform -1 0 8790 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__2499_
timestamp 1728341909
transform 1 0 9030 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2500_
timestamp 1728341909
transform -1 0 7650 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2501_
timestamp 1728341909
transform -1 0 6770 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__2502_
timestamp 1728341909
transform -1 0 7630 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__2503_
timestamp 1728341909
transform 1 0 11130 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2504_
timestamp 1728341909
transform -1 0 4570 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2505_
timestamp 1728341909
transform -1 0 5710 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2506_
timestamp 1728341909
transform -1 0 6730 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__2507_
timestamp 1728341909
transform 1 0 5870 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2508_
timestamp 1728341909
transform 1 0 5670 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2509_
timestamp 1728341909
transform -1 0 8830 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__2510_
timestamp 1728341909
transform -1 0 8090 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__2511_
timestamp 1728341909
transform -1 0 7410 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__2512_
timestamp 1728341909
transform 1 0 7110 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__2513_
timestamp 1728341909
transform 1 0 6890 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__2514_
timestamp 1728341909
transform 1 0 7050 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__2515_
timestamp 1728341909
transform 1 0 10390 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__2516_
timestamp 1728341909
transform 1 0 8530 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2517_
timestamp 1728341909
transform 1 0 10630 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2518_
timestamp 1728341909
transform -1 0 9730 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__2519_
timestamp 1728341909
transform 1 0 9970 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__2520_
timestamp 1728341909
transform -1 0 10430 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2521_
timestamp 1728341909
transform -1 0 8530 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2522_
timestamp 1728341909
transform 1 0 6090 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2523_
timestamp 1728341909
transform 1 0 5910 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2524_
timestamp 1728341909
transform 1 0 8290 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2525_
timestamp 1728341909
transform 1 0 6790 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2526_
timestamp 1728341909
transform -1 0 7790 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2527_
timestamp 1728341909
transform 1 0 8010 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2528_
timestamp 1728341909
transform -1 0 8070 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2529_
timestamp 1728341909
transform 1 0 7850 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2530_
timestamp 1728341909
transform -1 0 7810 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2531_
timestamp 1728341909
transform -1 0 7830 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2532_
timestamp 1728341909
transform 1 0 7830 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2533_
timestamp 1728341909
transform -1 0 5490 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2534_
timestamp 1728341909
transform -1 0 5910 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2535_
timestamp 1728341909
transform -1 0 7590 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2536_
timestamp 1728341909
transform 1 0 7390 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2537_
timestamp 1728341909
transform 1 0 7310 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2538_
timestamp 1728341909
transform 1 0 8030 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2539_
timestamp 1728341909
transform 1 0 5890 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2540_
timestamp 1728341909
transform 1 0 5610 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2541_
timestamp 1728341909
transform 1 0 6130 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2542_
timestamp 1728341909
transform -1 0 6670 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2543_
timestamp 1728341909
transform -1 0 6630 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2544_
timestamp 1728341909
transform 1 0 6170 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2545_
timestamp 1728341909
transform 1 0 6870 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2546_
timestamp 1728341909
transform 1 0 6130 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2547_
timestamp 1728341909
transform 1 0 6350 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2548_
timestamp 1728341909
transform 1 0 7130 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2549_
timestamp 1728341909
transform 1 0 7390 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2550_
timestamp 1728341909
transform -1 0 7550 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2551_
timestamp 1728341909
transform -1 0 6270 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2552_
timestamp 1728341909
transform -1 0 4830 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2553_
timestamp 1728341909
transform -1 0 5870 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2554_
timestamp 1728341909
transform -1 0 5590 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2555_
timestamp 1728341909
transform 1 0 5650 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2556_
timestamp 1728341909
transform 1 0 5030 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2557_
timestamp 1728341909
transform 1 0 5770 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2558_
timestamp 1728341909
transform -1 0 6410 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2559_
timestamp 1728341909
transform 1 0 6090 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__2560_
timestamp 1728341909
transform 1 0 4350 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2561_
timestamp 1728341909
transform -1 0 5410 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2562_
timestamp 1728341909
transform 1 0 5030 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2563_
timestamp 1728341909
transform -1 0 4930 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2564_
timestamp 1728341909
transform -1 0 4590 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2565_
timestamp 1728341909
transform 1 0 4730 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2566_
timestamp 1728341909
transform -1 0 4950 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2567_
timestamp 1728341909
transform 1 0 5150 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2568_
timestamp 1728341909
transform 1 0 5290 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__2569_
timestamp 1728341909
transform -1 0 4170 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2570_
timestamp 1728341909
transform 1 0 5190 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2571_
timestamp 1728341909
transform 1 0 4310 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2572_
timestamp 1728341909
transform -1 0 4430 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2573_
timestamp 1728341909
transform 1 0 4670 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2574_
timestamp 1728341909
transform 1 0 5390 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2575_
timestamp 1728341909
transform -1 0 4950 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2576_
timestamp 1728341909
transform 1 0 5130 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2577_
timestamp 1728341909
transform 1 0 4870 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2578_
timestamp 1728341909
transform -1 0 4810 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2579_
timestamp 1728341909
transform 1 0 4670 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__2580_
timestamp 1728341909
transform 1 0 4710 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__2581_
timestamp 1728341909
transform -1 0 4150 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2582_
timestamp 1728341909
transform -1 0 3290 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2583_
timestamp 1728341909
transform 1 0 2230 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2584_
timestamp 1728341909
transform 1 0 3190 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2585_
timestamp 1728341909
transform -1 0 6350 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2586_
timestamp 1728341909
transform -1 0 3710 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2587_
timestamp 1728341909
transform -1 0 3450 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2588_
timestamp 1728341909
transform -1 0 2970 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2589_
timestamp 1728341909
transform -1 0 2970 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2590_
timestamp 1728341909
transform 1 0 3590 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__2591_
timestamp 1728341909
transform -1 0 3070 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2592_
timestamp 1728341909
transform 1 0 2570 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2593_
timestamp 1728341909
transform -1 0 2670 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2594_
timestamp 1728341909
transform -1 0 2690 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2595_
timestamp 1728341909
transform -1 0 3770 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__2596_
timestamp 1728341909
transform 1 0 3370 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2597_
timestamp 1728341909
transform 1 0 3310 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2598_
timestamp 1728341909
transform -1 0 3190 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2599_
timestamp 1728341909
transform -1 0 3190 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2600_
timestamp 1728341909
transform 1 0 2910 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2601_
timestamp 1728341909
transform -1 0 2470 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2602_
timestamp 1728341909
transform -1 0 2730 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2603_
timestamp 1728341909
transform -1 0 2330 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2604_
timestamp 1728341909
transform 1 0 2470 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2605_
timestamp 1728341909
transform -1 0 2470 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2606_
timestamp 1728341909
transform 1 0 2190 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2607_
timestamp 1728341909
transform -1 0 1550 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2608_
timestamp 1728341909
transform -1 0 1070 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2609_
timestamp 1728341909
transform 1 0 2030 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2610_
timestamp 1728341909
transform 1 0 1270 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2611_
timestamp 1728341909
transform -1 0 1250 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2612_
timestamp 1728341909
transform -1 0 990 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2613_
timestamp 1728341909
transform -1 0 1970 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2614_
timestamp 1728341909
transform -1 0 590 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2615_
timestamp 1728341909
transform 1 0 1770 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2616_
timestamp 1728341909
transform 1 0 1510 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2617_
timestamp 1728341909
transform -1 0 1510 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2618_
timestamp 1728341909
transform -1 0 1750 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2619_
timestamp 1728341909
transform 1 0 790 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2620_
timestamp 1728341909
transform -1 0 1310 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2621_
timestamp 1728341909
transform 1 0 1050 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2622_
timestamp 1728341909
transform -1 0 1270 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2623_
timestamp 1728341909
transform 1 0 1010 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2624_
timestamp 1728341909
transform -1 0 550 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2625_
timestamp 1728341909
transform -1 0 2630 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2626_
timestamp 1728341909
transform 1 0 1650 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2627_
timestamp 1728341909
transform 1 0 1390 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2628_
timestamp 1728341909
transform 1 0 790 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2629_
timestamp 1728341909
transform -1 0 3390 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__2630_
timestamp 1728341909
transform 1 0 4250 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__2631_
timestamp 1728341909
transform -1 0 4910 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__2632_
timestamp 1728341909
transform 1 0 10890 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2633_
timestamp 1728341909
transform 1 0 3890 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2634_
timestamp 1728341909
transform 1 0 8990 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2635_
timestamp 1728341909
transform -1 0 2270 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__2636_
timestamp 1728341909
transform -1 0 9150 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__2637_
timestamp 1728341909
transform 1 0 4350 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2638_
timestamp 1728341909
transform 1 0 4850 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2639_
timestamp 1728341909
transform -1 0 9930 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__2640_
timestamp 1728341909
transform -1 0 9870 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__2641_
timestamp 1728341909
transform 1 0 10170 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2642_
timestamp 1728341909
transform -1 0 9510 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__2643_
timestamp 1728341909
transform 1 0 10910 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2644_
timestamp 1728341909
transform -1 0 9750 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2645_
timestamp 1728341909
transform -1 0 9710 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__2646_
timestamp 1728341909
transform 1 0 10110 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__2647_
timestamp 1728341909
transform -1 0 8590 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2648_
timestamp 1728341909
transform -1 0 4170 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__2649_
timestamp 1728341909
transform -1 0 5810 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2650_
timestamp 1728341909
transform 1 0 9310 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__2651_
timestamp 1728341909
transform -1 0 5690 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2652_
timestamp 1728341909
transform -1 0 7850 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__2653_
timestamp 1728341909
transform -1 0 7750 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__2654_
timestamp 1728341909
transform 1 0 4670 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2655_
timestamp 1728341909
transform -1 0 5450 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2656_
timestamp 1728341909
transform -1 0 6030 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2657_
timestamp 1728341909
transform -1 0 6770 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2658_
timestamp 1728341909
transform 1 0 6270 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2659_
timestamp 1728341909
transform 1 0 6970 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2660_
timestamp 1728341909
transform -1 0 7250 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2661_
timestamp 1728341909
transform -1 0 4470 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2662_
timestamp 1728341909
transform 1 0 4430 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2663_
timestamp 1728341909
transform 1 0 6350 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2664_
timestamp 1728341909
transform -1 0 6610 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2665_
timestamp 1728341909
transform 1 0 7110 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2666_
timestamp 1728341909
transform 1 0 6850 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2667_
timestamp 1728341909
transform 1 0 7590 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2668_
timestamp 1728341909
transform 1 0 7330 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2669_
timestamp 1728341909
transform 1 0 7990 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2670_
timestamp 1728341909
transform -1 0 4210 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2671_
timestamp 1728341909
transform -1 0 5330 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__2672_
timestamp 1728341909
transform 1 0 5230 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2673_
timestamp 1728341909
transform 1 0 7190 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2674_
timestamp 1728341909
transform -1 0 7410 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2675_
timestamp 1728341909
transform 1 0 7650 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2676_
timestamp 1728341909
transform -1 0 7590 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2677_
timestamp 1728341909
transform 1 0 7770 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2678_
timestamp 1728341909
transform 1 0 7730 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2679_
timestamp 1728341909
transform 1 0 4170 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2680_
timestamp 1728341909
transform -1 0 4430 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2681_
timestamp 1728341909
transform 1 0 6130 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2682_
timestamp 1728341909
transform 1 0 6750 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2683_
timestamp 1728341909
transform 1 0 4090 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2684_
timestamp 1728341909
transform -1 0 5750 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2685_
timestamp 1728341909
transform 1 0 5470 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2686_
timestamp 1728341909
transform -1 0 6890 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2687_
timestamp 1728341909
transform 1 0 7350 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2688_
timestamp 1728341909
transform -1 0 7490 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2689_
timestamp 1728341909
transform 1 0 6510 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2690_
timestamp 1728341909
transform 1 0 6590 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2691_
timestamp 1728341909
transform 1 0 7090 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2692_
timestamp 1728341909
transform -1 0 7230 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2693_
timestamp 1728341909
transform 1 0 5070 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2694_
timestamp 1728341909
transform -1 0 5210 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2695_
timestamp 1728341909
transform 1 0 6650 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2696_
timestamp 1728341909
transform 1 0 6590 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2697_
timestamp 1728341909
transform 1 0 7010 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2698_
timestamp 1728341909
transform 1 0 6910 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2699_
timestamp 1728341909
transform -1 0 6350 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2700_
timestamp 1728341909
transform 1 0 5410 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2701_
timestamp 1728341909
transform -1 0 5490 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2702_
timestamp 1728341909
transform -1 0 5570 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2703_
timestamp 1728341909
transform -1 0 5590 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2704_
timestamp 1728341909
transform 1 0 5650 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2705_
timestamp 1728341909
transform 1 0 5910 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2706_
timestamp 1728341909
transform -1 0 6170 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2707_
timestamp 1728341909
transform -1 0 5910 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2708_
timestamp 1728341909
transform -1 0 2310 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2709_
timestamp 1728341909
transform -1 0 4970 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2710_
timestamp 1728341909
transform -1 0 4890 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2711_
timestamp 1728341909
transform -1 0 5090 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2712_
timestamp 1728341909
transform -1 0 5670 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2713_
timestamp 1728341909
transform -1 0 5810 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2714_
timestamp 1728341909
transform -1 0 6110 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2715_
timestamp 1728341909
transform 1 0 5830 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2716_
timestamp 1728341909
transform -1 0 6670 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2717_
timestamp 1728341909
transform 1 0 6610 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2718_
timestamp 1728341909
transform 1 0 6190 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2719_
timestamp 1728341909
transform -1 0 6350 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2720_
timestamp 1728341909
transform 1 0 4650 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2721_
timestamp 1728341909
transform 1 0 4930 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2722_
timestamp 1728341909
transform 1 0 5170 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2723_
timestamp 1728341909
transform -1 0 5430 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2724_
timestamp 1728341909
transform 1 0 6150 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2725_
timestamp 1728341909
transform 1 0 6390 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2726_
timestamp 1728341909
transform -1 0 6150 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__2727_
timestamp 1728341909
transform 1 0 5850 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__2728_
timestamp 1728341909
transform -1 0 4330 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2729_
timestamp 1728341909
transform -1 0 4190 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2730_
timestamp 1728341909
transform -1 0 5230 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2731_
timestamp 1728341909
transform -1 0 5350 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2732_
timestamp 1728341909
transform -1 0 5650 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2733_
timestamp 1728341909
transform -1 0 5910 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2734_
timestamp 1728341909
transform -1 0 5230 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2735_
timestamp 1728341909
transform 1 0 5430 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2736_
timestamp 1728341909
transform -1 0 8350 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__2737_
timestamp 1728341909
transform 1 0 3750 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2738_
timestamp 1728341909
transform 1 0 3930 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2739_
timestamp 1728341909
transform -1 0 3750 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2740_
timestamp 1728341909
transform -1 0 3690 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2741_
timestamp 1728341909
transform -1 0 4030 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2742_
timestamp 1728341909
transform -1 0 4170 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2743_
timestamp 1728341909
transform 1 0 4910 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2744_
timestamp 1728341909
transform 1 0 4650 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__2745_
timestamp 1728341909
transform 1 0 5130 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2746_
timestamp 1728341909
transform 1 0 4630 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2747_
timestamp 1728341909
transform 1 0 5550 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2748_
timestamp 1728341909
transform -1 0 4950 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2749_
timestamp 1728341909
transform -1 0 5310 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2750_
timestamp 1728341909
transform -1 0 5410 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2751_
timestamp 1728341909
transform 1 0 4390 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2752_
timestamp 1728341909
transform 1 0 3890 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2753_
timestamp 1728341909
transform -1 0 3430 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2754_
timestamp 1728341909
transform -1 0 3010 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2755_
timestamp 1728341909
transform 1 0 3270 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2756_
timestamp 1728341909
transform -1 0 3650 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2757_
timestamp 1728341909
transform -1 0 3670 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2758_
timestamp 1728341909
transform -1 0 3650 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2759_
timestamp 1728341909
transform -1 0 3530 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2760_
timestamp 1728341909
transform -1 0 3570 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2761_
timestamp 1728341909
transform -1 0 3710 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2762_
timestamp 1728341909
transform -1 0 3470 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2763_
timestamp 1728341909
transform 1 0 3030 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__2764_
timestamp 1728341909
transform 1 0 3310 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__2765_
timestamp 1728341909
transform -1 0 2630 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2766_
timestamp 1728341909
transform 1 0 3710 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__2767_
timestamp 1728341909
transform -1 0 4410 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2768_
timestamp 1728341909
transform 1 0 4490 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2769_
timestamp 1728341909
transform 1 0 5150 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2770_
timestamp 1728341909
transform -1 0 4650 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2771_
timestamp 1728341909
transform -1 0 4930 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2772_
timestamp 1728341909
transform -1 0 4910 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2773_
timestamp 1728341909
transform 1 0 2670 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2774_
timestamp 1728341909
transform -1 0 2530 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__2775_
timestamp 1728341909
transform 1 0 3890 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2776_
timestamp 1728341909
transform 1 0 4410 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2777_
timestamp 1728341909
transform 1 0 5150 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2778_
timestamp 1728341909
transform -1 0 4650 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2779_
timestamp 1728341909
transform 1 0 3970 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__2780_
timestamp 1728341909
transform 1 0 2750 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__2781_
timestamp 1728341909
transform -1 0 3970 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2782_
timestamp 1728341909
transform -1 0 2770 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2783_
timestamp 1728341909
transform 1 0 2470 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2784_
timestamp 1728341909
transform 1 0 550 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2785_
timestamp 1728341909
transform -1 0 2250 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2786_
timestamp 1728341909
transform 1 0 2510 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2787_
timestamp 1728341909
transform -1 0 2930 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2788_
timestamp 1728341909
transform -1 0 2430 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2789_
timestamp 1728341909
transform -1 0 3730 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2790_
timestamp 1728341909
transform 1 0 3210 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2791_
timestamp 1728341909
transform -1 0 2950 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2792_
timestamp 1728341909
transform -1 0 2850 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2793_
timestamp 1728341909
transform -1 0 2270 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__2794_
timestamp 1728341909
transform 1 0 2150 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2795_
timestamp 1728341909
transform 1 0 790 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2796_
timestamp 1728341909
transform 1 0 1730 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2797_
timestamp 1728341909
transform -1 0 2010 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2798_
timestamp 1728341909
transform 1 0 1230 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2799_
timestamp 1728341909
transform -1 0 1510 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2800_
timestamp 1728341909
transform -1 0 1770 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2801_
timestamp 1728341909
transform 1 0 1730 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2802_
timestamp 1728341909
transform 1 0 1810 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2803_
timestamp 1728341909
transform 1 0 3290 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2804_
timestamp 1728341909
transform -1 0 450 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__2805_
timestamp 1728341909
transform 1 0 6990 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2806_
timestamp 1728341909
transform -1 0 5410 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2807_
timestamp 1728341909
transform -1 0 5010 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2808_
timestamp 1728341909
transform 1 0 3930 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2809_
timestamp 1728341909
transform -1 0 4390 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2810_
timestamp 1728341909
transform -1 0 4750 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2811_
timestamp 1728341909
transform -1 0 4610 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2812_
timestamp 1728341909
transform 1 0 4230 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2813_
timestamp 1728341909
transform 1 0 3990 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__2814_
timestamp 1728341909
transform 1 0 4110 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__2815_
timestamp 1728341909
transform -1 0 4190 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2816_
timestamp 1728341909
transform 1 0 2490 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2817_
timestamp 1728341909
transform -1 0 2770 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__2818_
timestamp 1728341909
transform 1 0 2730 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2819_
timestamp 1728341909
transform 1 0 3170 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2820_
timestamp 1728341909
transform 1 0 3410 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2821_
timestamp 1728341909
transform -1 0 3950 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2822_
timestamp 1728341909
transform -1 0 4750 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2823_
timestamp 1728341909
transform -1 0 1730 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2824_
timestamp 1728341909
transform 1 0 550 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__2825_
timestamp 1728341909
transform 1 0 530 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2826_
timestamp 1728341909
transform -1 0 690 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__2827_
timestamp 1728341909
transform 1 0 1730 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2828_
timestamp 1728341909
transform -1 0 2010 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2829_
timestamp 1728341909
transform 1 0 1250 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2830_
timestamp 1728341909
transform -1 0 1510 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2831_
timestamp 1728341909
transform -1 0 1530 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__2832_
timestamp 1728341909
transform 1 0 2030 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2833_
timestamp 1728341909
transform -1 0 1050 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__2834_
timestamp 1728341909
transform 1 0 870 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__2835_
timestamp 1728341909
transform 1 0 1110 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__2836_
timestamp 1728341909
transform 1 0 1330 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__2837_
timestamp 1728341909
transform 1 0 1650 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__2838_
timestamp 1728341909
transform -1 0 1530 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__2839_
timestamp 1728341909
transform 1 0 810 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__2840_
timestamp 1728341909
transform 1 0 1250 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2841_
timestamp 1728341909
transform 1 0 2050 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2842_
timestamp 1728341909
transform -1 0 1710 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2843_
timestamp 1728341909
transform -1 0 1810 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2844_
timestamp 1728341909
transform -1 0 1570 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__2845_
timestamp 1728341909
transform -1 0 1510 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2846_
timestamp 1728341909
transform 1 0 1290 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2847_
timestamp 1728341909
transform -1 0 1290 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__2848_
timestamp 1728341909
transform -1 0 1270 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2849_
timestamp 1728341909
transform -1 0 1570 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2850_
timestamp 1728341909
transform -1 0 1490 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2851_
timestamp 1728341909
transform -1 0 1030 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2852_
timestamp 1728341909
transform -1 0 1090 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2853_
timestamp 1728341909
transform -1 0 2290 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2854_
timestamp 1728341909
transform 1 0 770 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__2855_
timestamp 1728341909
transform 1 0 2450 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__2856_
timestamp 1728341909
transform -1 0 1970 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__2857_
timestamp 1728341909
transform -1 0 2370 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__2858_
timestamp 1728341909
transform -1 0 2270 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__2859_
timestamp 1728341909
transform -1 0 850 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2860_
timestamp 1728341909
transform 1 0 530 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2861_
timestamp 1728341909
transform -1 0 90 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2862_
timestamp 1728341909
transform -1 0 1050 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__2863_
timestamp 1728341909
transform 1 0 290 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__2864_
timestamp 1728341909
transform -1 0 330 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__2865_
timestamp 1728341909
transform 1 0 4450 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__2866_
timestamp 1728341909
transform 1 0 4470 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2867_
timestamp 1728341909
transform 1 0 5570 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__2868_
timestamp 1728341909
transform -1 0 2950 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2869_
timestamp 1728341909
transform -1 0 3230 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__2870_
timestamp 1728341909
transform -1 0 2290 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__2871_
timestamp 1728341909
transform 1 0 2310 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__2872_
timestamp 1728341909
transform -1 0 4590 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__2873_
timestamp 1728341909
transform 1 0 4330 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__2874_
timestamp 1728341909
transform -1 0 4130 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2875_
timestamp 1728341909
transform -1 0 1690 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2876_
timestamp 1728341909
transform -1 0 830 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2877_
timestamp 1728341909
transform -1 0 3490 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2878_
timestamp 1728341909
transform -1 0 3930 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2879_
timestamp 1728341909
transform -1 0 1270 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2880_
timestamp 1728341909
transform 1 0 1450 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2881_
timestamp 1728341909
transform -1 0 1770 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2882_
timestamp 1728341909
transform -1 0 2450 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2883_
timestamp 1728341909
transform 1 0 4450 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2884_
timestamp 1728341909
transform 1 0 4170 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2885_
timestamp 1728341909
transform 1 0 3110 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2886_
timestamp 1728341909
transform 1 0 4670 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2887_
timestamp 1728341909
transform 1 0 5130 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2888_
timestamp 1728341909
transform 1 0 3390 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2889_
timestamp 1728341909
transform 1 0 3610 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2890_
timestamp 1728341909
transform -1 0 4390 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2891_
timestamp 1728341909
transform -1 0 4130 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2892_
timestamp 1728341909
transform -1 0 1990 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2893_
timestamp 1728341909
transform 1 0 3670 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2894_
timestamp 1728341909
transform 1 0 3870 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2895_
timestamp 1728341909
transform 1 0 4450 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2896_
timestamp 1728341909
transform -1 0 3850 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2897_
timestamp 1728341909
transform -1 0 5850 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2898_
timestamp 1728341909
transform 1 0 5170 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2899_
timestamp 1728341909
transform 1 0 5130 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2900_
timestamp 1728341909
transform 1 0 5390 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2901_
timestamp 1728341909
transform -1 0 4870 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2902_
timestamp 1728341909
transform -1 0 1530 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2903_
timestamp 1728341909
transform 1 0 2190 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2904_
timestamp 1728341909
transform 1 0 2450 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2905_
timestamp 1728341909
transform 1 0 1250 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2906_
timestamp 1728341909
transform 1 0 1030 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2907_
timestamp 1728341909
transform 1 0 1230 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2908_
timestamp 1728341909
transform -1 0 1550 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2909_
timestamp 1728341909
transform -1 0 1770 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2910_
timestamp 1728341909
transform -1 0 1550 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2911_
timestamp 1728341909
transform -1 0 1550 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2912_
timestamp 1728341909
transform -1 0 2470 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2913_
timestamp 1728341909
transform -1 0 1710 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2914_
timestamp 1728341909
transform 1 0 2230 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2915_
timestamp 1728341909
transform 1 0 2010 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2916_
timestamp 1728341909
transform 1 0 1690 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2917_
timestamp 1728341909
transform -1 0 1770 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2918_
timestamp 1728341909
transform 1 0 1710 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2919_
timestamp 1728341909
transform -1 0 2250 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2920_
timestamp 1728341909
transform -1 0 1970 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2921_
timestamp 1728341909
transform -1 0 2030 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2922_
timestamp 1728341909
transform -1 0 1950 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2923_
timestamp 1728341909
transform -1 0 1990 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2924_
timestamp 1728341909
transform -1 0 2950 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2925_
timestamp 1728341909
transform 1 0 3430 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2926_
timestamp 1728341909
transform -1 0 2410 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2927_
timestamp 1728341909
transform -1 0 2450 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2928_
timestamp 1728341909
transform 1 0 4590 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2929_
timestamp 1728341909
transform 1 0 3430 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2930_
timestamp 1728341909
transform -1 0 2710 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2931_
timestamp 1728341909
transform -1 0 2950 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2932_
timestamp 1728341909
transform 1 0 3150 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2933_
timestamp 1728341909
transform -1 0 2710 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2934_
timestamp 1728341909
transform 1 0 2930 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2935_
timestamp 1728341909
transform -1 0 1310 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2936_
timestamp 1728341909
transform -1 0 850 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2937_
timestamp 1728341909
transform 1 0 570 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2938_
timestamp 1728341909
transform 1 0 1730 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2939_
timestamp 1728341909
transform -1 0 1510 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2940_
timestamp 1728341909
transform 1 0 3170 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2941_
timestamp 1728341909
transform 1 0 3170 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2942_
timestamp 1728341909
transform -1 0 3390 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2943_
timestamp 1728341909
transform -1 0 3230 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2944_
timestamp 1728341909
transform -1 0 3730 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2945_
timestamp 1728341909
transform 1 0 3170 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__2946_
timestamp 1728341909
transform 1 0 3610 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__2947_
timestamp 1728341909
transform 1 0 3190 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2948_
timestamp 1728341909
transform -1 0 4190 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2949_
timestamp 1728341909
transform 1 0 3150 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__2950_
timestamp 1728341909
transform 1 0 2470 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2951_
timestamp 1728341909
transform -1 0 2710 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2952_
timestamp 1728341909
transform -1 0 2990 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2953_
timestamp 1728341909
transform -1 0 2190 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2954_
timestamp 1728341909
transform -1 0 2430 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2955_
timestamp 1728341909
transform 1 0 3010 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__2956_
timestamp 1728341909
transform 1 0 3250 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__2957_
timestamp 1728341909
transform 1 0 3750 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__2958_
timestamp 1728341909
transform 1 0 2190 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__2959_
timestamp 1728341909
transform 1 0 3470 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__2960_
timestamp 1728341909
transform 1 0 3590 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__2961_
timestamp 1728341909
transform 1 0 2710 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2962_
timestamp 1728341909
transform 1 0 2450 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2963_
timestamp 1728341909
transform 1 0 2970 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2964_
timestamp 1728341909
transform 1 0 2710 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2965_
timestamp 1728341909
transform -1 0 5790 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2966_
timestamp 1728341909
transform 1 0 4110 0 1 1690
box -12 -8 32 252
use FILL  FILL_3__2967_
timestamp 1728341909
transform -1 0 4590 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2968_
timestamp 1728341909
transform -1 0 4830 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2969_
timestamp 1728341909
transform -1 0 1330 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__2970_
timestamp 1728341909
transform -1 0 1510 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__2971_
timestamp 1728341909
transform -1 0 1530 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2972_
timestamp 1728341909
transform -1 0 1270 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2973_
timestamp 1728341909
transform -1 0 1030 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__2974_
timestamp 1728341909
transform -1 0 1770 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2975_
timestamp 1728341909
transform -1 0 1990 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2976_
timestamp 1728341909
transform 1 0 3870 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2977_
timestamp 1728341909
transform -1 0 4430 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2978_
timestamp 1728341909
transform 1 0 4150 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2979_
timestamp 1728341909
transform 1 0 1530 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2980_
timestamp 1728341909
transform -1 0 1010 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2981_
timestamp 1728341909
transform -1 0 770 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2982_
timestamp 1728341909
transform 1 0 2210 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2983_
timestamp 1728341909
transform -1 0 530 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2984_
timestamp 1728341909
transform -1 0 310 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2985_
timestamp 1728341909
transform -1 0 90 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__2986_
timestamp 1728341909
transform -1 0 350 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2987_
timestamp 1728341909
transform -1 0 610 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2988_
timestamp 1728341909
transform -1 0 570 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2989_
timestamp 1728341909
transform 1 0 330 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2990_
timestamp 1728341909
transform 1 0 70 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2991_
timestamp 1728341909
transform -1 0 350 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2992_
timestamp 1728341909
transform -1 0 2010 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__2993_
timestamp 1728341909
transform -1 0 1050 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2994_
timestamp 1728341909
transform -1 0 810 0 1 730
box -12 -8 32 252
use FILL  FILL_3__2995_
timestamp 1728341909
transform 1 0 590 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__2996_
timestamp 1728341909
transform -1 0 530 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__2997_
timestamp 1728341909
transform -1 0 850 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__2998_
timestamp 1728341909
transform -1 0 90 0 1 250
box -12 -8 32 252
use FILL  FILL_3__2999_
timestamp 1728341909
transform -1 0 330 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__3000_
timestamp 1728341909
transform -1 0 90 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__3001_
timestamp 1728341909
transform -1 0 90 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__3002_
timestamp 1728341909
transform -1 0 570 0 1 730
box -12 -8 32 252
use FILL  FILL_3__3003_
timestamp 1728341909
transform -1 0 90 0 1 730
box -12 -8 32 252
use FILL  FILL_3__3004_
timestamp 1728341909
transform -1 0 830 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__3005_
timestamp 1728341909
transform 1 0 790 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__3006_
timestamp 1728341909
transform -1 0 90 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__3007_
timestamp 1728341909
transform 1 0 1790 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3008_
timestamp 1728341909
transform -1 0 1050 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__3009_
timestamp 1728341909
transform -1 0 1310 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__3010_
timestamp 1728341909
transform -1 0 1310 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__3011_
timestamp 1728341909
transform -1 0 1070 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3__3012_
timestamp 1728341909
transform -1 0 1450 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__3013_
timestamp 1728341909
transform -1 0 1230 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__3014_
timestamp 1728341909
transform 1 0 1030 0 1 250
box -12 -8 32 252
use FILL  FILL_3__3015_
timestamp 1728341909
transform -1 0 1530 0 1 250
box -12 -8 32 252
use FILL  FILL_3__3016_
timestamp 1728341909
transform -1 0 1290 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__3017_
timestamp 1728341909
transform -1 0 1270 0 1 250
box -12 -8 32 252
use FILL  FILL_3__3018_
timestamp 1728341909
transform 1 0 1050 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3__3019_
timestamp 1728341909
transform -1 0 1050 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__3020_
timestamp 1728341909
transform -1 0 3690 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3021_
timestamp 1728341909
transform -1 0 5950 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__3022_
timestamp 1728341909
transform 1 0 2790 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3023_
timestamp 1728341909
transform 1 0 2810 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3024_
timestamp 1728341909
transform 1 0 3790 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3025_
timestamp 1728341909
transform -1 0 4210 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__3026_
timestamp 1728341909
transform -1 0 3070 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3027_
timestamp 1728341909
transform -1 0 3470 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__3028_
timestamp 1728341909
transform -1 0 3990 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3029_
timestamp 1728341909
transform -1 0 4490 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3030_
timestamp 1728341909
transform 1 0 3470 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__3031_
timestamp 1728341909
transform -1 0 3750 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__3032_
timestamp 1728341909
transform -1 0 2550 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3033_
timestamp 1728341909
transform -1 0 2570 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3034_
timestamp 1728341909
transform 1 0 2710 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__3035_
timestamp 1728341909
transform -1 0 2970 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__3036_
timestamp 1728341909
transform 1 0 3290 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3037_
timestamp 1728341909
transform -1 0 3730 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__3038_
timestamp 1728341909
transform -1 0 3290 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3039_
timestamp 1728341909
transform 1 0 3030 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3040_
timestamp 1728341909
transform 1 0 2170 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__3041_
timestamp 1728341909
transform 1 0 2710 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__3042_
timestamp 1728341909
transform 1 0 7470 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__3043_
timestamp 1728341909
transform 1 0 6310 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__3044_
timestamp 1728341909
transform 1 0 5330 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__3045_
timestamp 1728341909
transform 1 0 5750 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3046_
timestamp 1728341909
transform 1 0 5470 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__3047_
timestamp 1728341909
transform 1 0 4810 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__3048_
timestamp 1728341909
transform 1 0 5150 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__3049_
timestamp 1728341909
transform 1 0 5850 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3050_
timestamp 1728341909
transform -1 0 6870 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3051_
timestamp 1728341909
transform -1 0 6330 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__3052_
timestamp 1728341909
transform 1 0 6370 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3053_
timestamp 1728341909
transform 1 0 6110 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3054_
timestamp 1728341909
transform 1 0 5850 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3055_
timestamp 1728341909
transform -1 0 5950 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3056_
timestamp 1728341909
transform 1 0 4610 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__3057_
timestamp 1728341909
transform 1 0 4370 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__3058_
timestamp 1728341909
transform -1 0 4490 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3059_
timestamp 1728341909
transform 1 0 4310 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__3060_
timestamp 1728341909
transform -1 0 4290 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__3061_
timestamp 1728341909
transform 1 0 3990 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3062_
timestamp 1728341909
transform -1 0 4810 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__3063_
timestamp 1728341909
transform 1 0 4550 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__3064_
timestamp 1728341909
transform 1 0 6010 0 1 2170
box -12 -8 32 252
use FILL  FILL_3__3065_
timestamp 1728341909
transform 1 0 5790 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__3066_
timestamp 1728341909
transform -1 0 5790 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3067_
timestamp 1728341909
transform -1 0 5930 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__3068_
timestamp 1728341909
transform -1 0 6970 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3069_
timestamp 1728341909
transform -1 0 6470 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3070_
timestamp 1728341909
transform 1 0 6110 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3071_
timestamp 1728341909
transform -1 0 6390 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3072_
timestamp 1728341909
transform 1 0 6590 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__3073_
timestamp 1728341909
transform 1 0 6350 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__3074_
timestamp 1728341909
transform 1 0 410 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__3075_
timestamp 1728341909
transform -1 0 570 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__3076_
timestamp 1728341909
transform -1 0 4270 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3077_
timestamp 1728341909
transform 1 0 2010 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3078_
timestamp 1728341909
transform -1 0 5510 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3079_
timestamp 1728341909
transform 1 0 5050 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3080_
timestamp 1728341909
transform 1 0 4250 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3081_
timestamp 1728341909
transform 1 0 5890 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__3082_
timestamp 1728341909
transform -1 0 6890 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__3083_
timestamp 1728341909
transform 1 0 6050 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__3084_
timestamp 1728341909
transform -1 0 5730 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3085_
timestamp 1728341909
transform -1 0 5010 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3086_
timestamp 1728341909
transform 1 0 5490 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3087_
timestamp 1728341909
transform -1 0 5090 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__3088_
timestamp 1728341909
transform -1 0 5630 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__3089_
timestamp 1728341909
transform -1 0 5590 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__3090_
timestamp 1728341909
transform 1 0 4770 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3091_
timestamp 1728341909
transform -1 0 4730 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3092_
timestamp 1728341909
transform 1 0 5590 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3__3093_
timestamp 1728341909
transform -1 0 3990 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__3094_
timestamp 1728341909
transform 1 0 4430 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__3095_
timestamp 1728341909
transform 1 0 4730 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__3096_
timestamp 1728341909
transform 1 0 4710 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__3097_
timestamp 1728341909
transform 1 0 4950 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__3098_
timestamp 1728341909
transform -1 0 5050 0 1 2650
box -12 -8 32 252
use FILL  FILL_3__3099_
timestamp 1728341909
transform 1 0 5190 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__3100_
timestamp 1728341909
transform -1 0 5590 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__3101_
timestamp 1728341909
transform 1 0 5130 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__3102_
timestamp 1728341909
transform 1 0 4650 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__3103_
timestamp 1728341909
transform 1 0 4870 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__3104_
timestamp 1728341909
transform -1 0 5010 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3105_
timestamp 1728341909
transform 1 0 5330 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__3106_
timestamp 1728341909
transform 1 0 8510 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__3107_
timestamp 1728341909
transform 1 0 8270 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__3108_
timestamp 1728341909
transform 1 0 8030 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__3109_
timestamp 1728341909
transform -1 0 8570 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3110_
timestamp 1728341909
transform -1 0 8330 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3111_
timestamp 1728341909
transform 1 0 4510 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3112_
timestamp 1728341909
transform 1 0 4750 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3113_
timestamp 1728341909
transform -1 0 1270 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3114_
timestamp 1728341909
transform 1 0 770 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3115_
timestamp 1728341909
transform 1 0 4450 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__3116_
timestamp 1728341909
transform -1 0 4070 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3117_
timestamp 1728341909
transform -1 0 330 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__3118_
timestamp 1728341909
transform -1 0 90 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__3119_
timestamp 1728341909
transform -1 0 4930 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__3120_
timestamp 1728341909
transform 1 0 4430 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3121_
timestamp 1728341909
transform 1 0 5170 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__3122_
timestamp 1728341909
transform -1 0 4470 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3123_
timestamp 1728341909
transform -1 0 3730 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3124_
timestamp 1728341909
transform -1 0 3950 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3125_
timestamp 1728341909
transform -1 0 3690 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3126_
timestamp 1728341909
transform 1 0 4710 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3127_
timestamp 1728341909
transform 1 0 4730 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3128_
timestamp 1728341909
transform 1 0 4650 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__3129_
timestamp 1728341909
transform 1 0 3730 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__3130_
timestamp 1728341909
transform -1 0 1830 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3131_
timestamp 1728341909
transform -1 0 1330 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3132_
timestamp 1728341909
transform 1 0 1050 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3133_
timestamp 1728341909
transform 1 0 3910 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3134_
timestamp 1728341909
transform 1 0 3490 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3135_
timestamp 1728341909
transform 1 0 3230 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3136_
timestamp 1728341909
transform 1 0 3710 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3137_
timestamp 1728341909
transform 1 0 3970 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3138_
timestamp 1728341909
transform -1 0 4010 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3139_
timestamp 1728341909
transform 1 0 1070 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3140_
timestamp 1728341909
transform 1 0 810 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3141_
timestamp 1728341909
transform -1 0 3990 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3142_
timestamp 1728341909
transform 1 0 3750 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3143_
timestamp 1728341909
transform -1 0 4190 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3144_
timestamp 1728341909
transform -1 0 3470 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3145_
timestamp 1728341909
transform 1 0 3210 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3146_
timestamp 1728341909
transform -1 0 3290 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3147_
timestamp 1728341909
transform 1 0 3530 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3148_
timestamp 1728341909
transform -1 0 3490 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3149_
timestamp 1728341909
transform -1 0 3470 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__3150_
timestamp 1728341909
transform 1 0 2050 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3151_
timestamp 1728341909
transform -1 0 2290 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3152_
timestamp 1728341909
transform 1 0 7530 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3153_
timestamp 1728341909
transform 1 0 4450 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3154_
timestamp 1728341909
transform -1 0 790 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3155_
timestamp 1728341909
transform 1 0 1010 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3156_
timestamp 1728341909
transform 1 0 2970 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3157_
timestamp 1728341909
transform -1 0 2750 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3158_
timestamp 1728341909
transform 1 0 1970 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3159_
timestamp 1728341909
transform 1 0 2510 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3160_
timestamp 1728341909
transform 1 0 3130 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3161_
timestamp 1728341909
transform -1 0 2670 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3162_
timestamp 1728341909
transform -1 0 2450 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3163_
timestamp 1728341909
transform -1 0 1550 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3164_
timestamp 1728341909
transform 1 0 1250 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3165_
timestamp 1728341909
transform -1 0 330 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3166_
timestamp 1728341909
transform -1 0 90 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3167_
timestamp 1728341909
transform 1 0 2050 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3168_
timestamp 1728341909
transform 1 0 1990 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3169_
timestamp 1728341909
transform -1 0 2290 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3170_
timestamp 1728341909
transform 1 0 2030 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3171_
timestamp 1728341909
transform -1 0 2230 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3172_
timestamp 1728341909
transform 1 0 1890 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__3173_
timestamp 1728341909
transform -1 0 1770 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3174_
timestamp 1728341909
transform -1 0 1790 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3175_
timestamp 1728341909
transform -1 0 3030 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3176_
timestamp 1728341909
transform -1 0 2830 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3177_
timestamp 1728341909
transform 1 0 2270 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3178_
timestamp 1728341909
transform 1 0 2610 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3179_
timestamp 1728341909
transform 1 0 2270 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3180_
timestamp 1728341909
transform 1 0 3210 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3181_
timestamp 1728341909
transform -1 0 2930 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3182_
timestamp 1728341909
transform -1 0 3010 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3183_
timestamp 1728341909
transform 1 0 2770 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3184_
timestamp 1728341909
transform -1 0 2530 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3185_
timestamp 1728341909
transform -1 0 2530 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3186_
timestamp 1728341909
transform 1 0 2010 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3187_
timestamp 1728341909
transform -1 0 350 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3188_
timestamp 1728341909
transform -1 0 90 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3189_
timestamp 1728341909
transform 1 0 1030 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3190_
timestamp 1728341909
transform -1 0 830 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3191_
timestamp 1728341909
transform -1 0 1090 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3192_
timestamp 1728341909
transform 1 0 1710 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3193_
timestamp 1728341909
transform 1 0 1450 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3194_
timestamp 1728341909
transform 1 0 3250 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3195_
timestamp 1728341909
transform 1 0 3210 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__3196_
timestamp 1728341909
transform 1 0 1950 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3197_
timestamp 1728341909
transform -1 0 2530 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__3198_
timestamp 1728341909
transform -1 0 2110 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3199_
timestamp 1728341909
transform -1 0 2370 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3200_
timestamp 1728341909
transform 1 0 810 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3201_
timestamp 1728341909
transform -1 0 1050 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3202_
timestamp 1728341909
transform 1 0 1050 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3203_
timestamp 1728341909
transform -1 0 1310 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3204_
timestamp 1728341909
transform -1 0 570 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3205_
timestamp 1728341909
transform -1 0 570 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3206_
timestamp 1728341909
transform 1 0 1070 0 -1 4090
box -12 -8 32 252
use FILL  FILL_3__3207_
timestamp 1728341909
transform -1 0 330 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3208_
timestamp 1728341909
transform -1 0 90 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3209_
timestamp 1728341909
transform 1 0 310 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3210_
timestamp 1728341909
transform -1 0 90 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3211_
timestamp 1728341909
transform -1 0 1570 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3212_
timestamp 1728341909
transform -1 0 1310 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3213_
timestamp 1728341909
transform 1 0 1590 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3214_
timestamp 1728341909
transform 1 0 1330 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3215_
timestamp 1728341909
transform -1 0 1290 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3216_
timestamp 1728341909
transform 1 0 1030 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3217_
timestamp 1728341909
transform -1 0 330 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3218_
timestamp 1728341909
transform -1 0 90 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3219_
timestamp 1728341909
transform -1 0 1610 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3220_
timestamp 1728341909
transform 1 0 1830 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3221_
timestamp 1728341909
transform -1 0 350 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3222_
timestamp 1728341909
transform -1 0 90 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3223_
timestamp 1728341909
transform -1 0 830 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__3224_
timestamp 1728341909
transform 1 0 550 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3225_
timestamp 1728341909
transform -1 0 330 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3226_
timestamp 1728341909
transform -1 0 90 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3227_
timestamp 1728341909
transform -1 0 350 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__3228_
timestamp 1728341909
transform -1 0 90 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__3229_
timestamp 1728341909
transform -1 0 2010 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__3230_
timestamp 1728341909
transform 1 0 1730 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__3231_
timestamp 1728341909
transform 1 0 1530 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__3232_
timestamp 1728341909
transform -1 0 1790 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__3233_
timestamp 1728341909
transform 1 0 1090 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3234_
timestamp 1728341909
transform -1 0 1370 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3235_
timestamp 1728341909
transform 1 0 1050 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3236_
timestamp 1728341909
transform 1 0 1310 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3237_
timestamp 1728341909
transform 1 0 2230 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__3238_
timestamp 1728341909
transform 1 0 2470 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3__3239_
timestamp 1728341909
transform -1 0 570 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3240_
timestamp 1728341909
transform -1 0 810 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3241_
timestamp 1728341909
transform 1 0 9710 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__3242_
timestamp 1728341909
transform -1 0 9050 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3__3243_
timestamp 1728341909
transform 1 0 9470 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__3244_
timestamp 1728341909
transform 1 0 8770 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__3245_
timestamp 1728341909
transform 1 0 9070 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3246_
timestamp 1728341909
transform -1 0 9590 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3247_
timestamp 1728341909
transform 1 0 10490 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3248_
timestamp 1728341909
transform 1 0 10750 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3249_
timestamp 1728341909
transform -1 0 9490 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__3250_
timestamp 1728341909
transform 1 0 9410 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3251_
timestamp 1728341909
transform 1 0 9250 0 1 3130
box -12 -8 32 252
use FILL  FILL_3__3252_
timestamp 1728341909
transform -1 0 9270 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__3253_
timestamp 1728341909
transform -1 0 7890 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3254_
timestamp 1728341909
transform -1 0 8150 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3255_
timestamp 1728341909
transform -1 0 9330 0 1 3610
box -12 -8 32 252
use FILL  FILL_3__3256_
timestamp 1728341909
transform 1 0 8270 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3257_
timestamp 1728341909
transform 1 0 8030 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3258_
timestamp 1728341909
transform 1 0 8570 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3259_
timestamp 1728341909
transform 1 0 9510 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3260_
timestamp 1728341909
transform -1 0 10870 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__3261_
timestamp 1728341909
transform -1 0 10410 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3262_
timestamp 1728341909
transform 1 0 9990 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3263_
timestamp 1728341909
transform 1 0 9670 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__3264_
timestamp 1728341909
transform 1 0 9010 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3__3265_
timestamp 1728341909
transform -1 0 9750 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3266_
timestamp 1728341909
transform 1 0 9770 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3267_
timestamp 1728341909
transform -1 0 9670 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3268_
timestamp 1728341909
transform -1 0 10010 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3269_
timestamp 1728341909
transform -1 0 10510 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3270_
timestamp 1728341909
transform 1 0 10230 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3271_
timestamp 1728341909
transform -1 0 10050 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3__3272_
timestamp 1728341909
transform 1 0 10270 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3__3273_
timestamp 1728341909
transform -1 0 10170 0 1 4570
box -12 -8 32 252
use FILL  FILL_3__3274_
timestamp 1728341909
transform -1 0 10270 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3275_
timestamp 1728341909
transform 1 0 9590 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__3276_
timestamp 1728341909
transform -1 0 9210 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3277_
timestamp 1728341909
transform -1 0 10670 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3278_
timestamp 1728341909
transform 1 0 10130 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3279_
timestamp 1728341909
transform -1 0 9910 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3280_
timestamp 1728341909
transform 1 0 9250 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__3281_
timestamp 1728341909
transform 1 0 9010 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__3282_
timestamp 1728341909
transform -1 0 6890 0 1 4090
box -12 -8 32 252
use FILL  FILL_3__3283_
timestamp 1728341909
transform -1 0 6830 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3284_
timestamp 1728341909
transform 1 0 6590 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3__3285_
timestamp 1728341909
transform 1 0 7030 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3286_
timestamp 1728341909
transform -1 0 7290 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3287_
timestamp 1728341909
transform -1 0 6650 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3288_
timestamp 1728341909
transform -1 0 6870 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3289_
timestamp 1728341909
transform -1 0 6830 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__3290_
timestamp 1728341909
transform 1 0 6550 0 1 5530
box -12 -8 32 252
use FILL  FILL_3__3291_
timestamp 1728341909
transform 1 0 7050 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3292_
timestamp 1728341909
transform -1 0 7310 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3293_
timestamp 1728341909
transform 1 0 7150 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3294_
timestamp 1728341909
transform 1 0 6890 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3295_
timestamp 1728341909
transform 1 0 6090 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3296_
timestamp 1728341909
transform 1 0 5830 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3297_
timestamp 1728341909
transform 1 0 5450 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3298_
timestamp 1728341909
transform 1 0 5190 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3299_
timestamp 1728341909
transform 1 0 5630 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3300_
timestamp 1728341909
transform 1 0 5390 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3301_
timestamp 1728341909
transform 1 0 6890 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3__3302_
timestamp 1728341909
transform 1 0 2970 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3303_
timestamp 1728341909
transform -1 0 3030 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3304_
timestamp 1728341909
transform 1 0 1970 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3305_
timestamp 1728341909
transform -1 0 2230 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3306_
timestamp 1728341909
transform 1 0 3890 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3307_
timestamp 1728341909
transform -1 0 4830 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3308_
timestamp 1728341909
transform -1 0 90 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__3309_
timestamp 1728341909
transform -1 0 90 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3310_
timestamp 1728341909
transform -1 0 770 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__3311_
timestamp 1728341909
transform -1 0 810 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3312_
timestamp 1728341909
transform -1 0 310 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__3313_
timestamp 1728341909
transform -1 0 350 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3314_
timestamp 1728341909
transform -1 0 90 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3315_
timestamp 1728341909
transform -1 0 90 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3316_
timestamp 1728341909
transform -1 0 590 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3317_
timestamp 1728341909
transform -1 0 810 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3449_
timestamp 1728341909
transform -1 0 3830 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3450_
timestamp 1728341909
transform 1 0 2990 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3451_
timestamp 1728341909
transform 1 0 3110 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3452_
timestamp 1728341909
transform -1 0 3370 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3453_
timestamp 1728341909
transform 1 0 3230 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3454_
timestamp 1728341909
transform -1 0 3590 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3455_
timestamp 1728341909
transform 1 0 9970 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3456_
timestamp 1728341909
transform 1 0 9530 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3457_
timestamp 1728341909
transform -1 0 9810 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3458_
timestamp 1728341909
transform -1 0 9970 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3459_
timestamp 1728341909
transform 1 0 10410 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3460_
timestamp 1728341909
transform -1 0 10710 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3461_
timestamp 1728341909
transform -1 0 10470 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3462_
timestamp 1728341909
transform -1 0 10030 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3463_
timestamp 1728341909
transform 1 0 10430 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3464_
timestamp 1728341909
transform -1 0 10230 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3465_
timestamp 1728341909
transform 1 0 10190 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3__3466_
timestamp 1728341909
transform -1 0 10210 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3467_
timestamp 1728341909
transform 1 0 8270 0 1 6010
box -12 -8 32 252
use FILL  FILL_3__3468_
timestamp 1728341909
transform 1 0 9110 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__3469_
timestamp 1728341909
transform 1 0 8570 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3470_
timestamp 1728341909
transform -1 0 8510 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3471_
timestamp 1728341909
transform 1 0 8650 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__3472_
timestamp 1728341909
transform 1 0 8890 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__3473_
timestamp 1728341909
transform -1 0 8710 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3474_
timestamp 1728341909
transform -1 0 8830 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3475_
timestamp 1728341909
transform -1 0 8950 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3476_
timestamp 1728341909
transform 1 0 9750 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3477_
timestamp 1728341909
transform 1 0 9190 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3478_
timestamp 1728341909
transform -1 0 9070 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3479_
timestamp 1728341909
transform 1 0 10550 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__3480_
timestamp 1728341909
transform -1 0 10110 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__3481_
timestamp 1728341909
transform -1 0 9970 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3482_
timestamp 1728341909
transform -1 0 9770 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__3483_
timestamp 1728341909
transform 1 0 10910 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3484_
timestamp 1728341909
transform 1 0 10890 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3485_
timestamp 1728341909
transform 1 0 11170 0 1 6490
box -12 -8 32 252
use FILL  FILL_3__3486_
timestamp 1728341909
transform 1 0 11130 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3487_
timestamp 1728341909
transform 1 0 10890 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3488_
timestamp 1728341909
transform 1 0 9530 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3489_
timestamp 1728341909
transform 1 0 9430 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3490_
timestamp 1728341909
transform -1 0 9690 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3491_
timestamp 1728341909
transform -1 0 9710 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3492_
timestamp 1728341909
transform 1 0 9910 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3493_
timestamp 1728341909
transform 1 0 10170 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3494_
timestamp 1728341909
transform 1 0 10310 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__3495_
timestamp 1728341909
transform -1 0 8810 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3496_
timestamp 1728341909
transform 1 0 9430 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3497_
timestamp 1728341909
transform 1 0 9950 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3498_
timestamp 1728341909
transform 1 0 9810 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__3499_
timestamp 1728341909
transform 1 0 9230 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3500_
timestamp 1728341909
transform -1 0 9490 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3501_
timestamp 1728341909
transform -1 0 9730 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3502_
timestamp 1728341909
transform 1 0 9570 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__3503_
timestamp 1728341909
transform 1 0 10050 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__3504_
timestamp 1728341909
transform -1 0 10010 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3505_
timestamp 1728341909
transform 1 0 10250 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3506_
timestamp 1728341909
transform 1 0 10770 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__3507_
timestamp 1728341909
transform -1 0 9390 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__3508_
timestamp 1728341909
transform -1 0 8510 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3509_
timestamp 1728341909
transform 1 0 8430 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__3510_
timestamp 1728341909
transform 1 0 9210 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3511_
timestamp 1728341909
transform -1 0 8970 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3512_
timestamp 1728341909
transform 1 0 8710 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3513_
timestamp 1728341909
transform -1 0 8990 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3514_
timestamp 1728341909
transform -1 0 8750 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3515_
timestamp 1728341909
transform -1 0 9150 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__3516_
timestamp 1728341909
transform 1 0 10990 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__3517_
timestamp 1728341909
transform -1 0 10310 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__3518_
timestamp 1728341909
transform 1 0 10390 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3519_
timestamp 1728341909
transform 1 0 10870 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3520_
timestamp 1728341909
transform -1 0 11170 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3521_
timestamp 1728341909
transform 1 0 7490 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3522_
timestamp 1728341909
transform -1 0 8010 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3523_
timestamp 1728341909
transform 1 0 8750 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3524_
timestamp 1728341909
transform 1 0 8530 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3525_
timestamp 1728341909
transform 1 0 8950 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3526_
timestamp 1728341909
transform -1 0 9230 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3527_
timestamp 1728341909
transform -1 0 8290 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3528_
timestamp 1728341909
transform -1 0 9930 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3529_
timestamp 1728341909
transform 1 0 10030 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__3530_
timestamp 1728341909
transform 1 0 10130 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3531_
timestamp 1728341909
transform -1 0 10170 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3532_
timestamp 1728341909
transform 1 0 10310 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__3533_
timestamp 1728341909
transform -1 0 8230 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3534_
timestamp 1728341909
transform -1 0 8490 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3535_
timestamp 1728341909
transform -1 0 8050 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3536_
timestamp 1728341909
transform -1 0 8270 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3537_
timestamp 1728341909
transform 1 0 8370 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__3538_
timestamp 1728341909
transform -1 0 8650 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__3539_
timestamp 1728341909
transform -1 0 9550 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__3540_
timestamp 1728341909
transform 1 0 9770 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__3541_
timestamp 1728341909
transform -1 0 9850 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__3542_
timestamp 1728341909
transform -1 0 7510 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3543_
timestamp 1728341909
transform -1 0 7770 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3544_
timestamp 1728341909
transform 1 0 7990 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3545_
timestamp 1728341909
transform 1 0 8850 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__3546_
timestamp 1728341909
transform -1 0 8290 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3547_
timestamp 1728341909
transform 1 0 8710 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3548_
timestamp 1728341909
transform -1 0 8970 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3549_
timestamp 1728341909
transform -1 0 8930 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__3550_
timestamp 1728341909
transform 1 0 8910 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3551_
timestamp 1728341909
transform 1 0 9190 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3552_
timestamp 1728341909
transform 1 0 9330 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__3553_
timestamp 1728341909
transform 1 0 9070 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__3554_
timestamp 1728341909
transform 1 0 8990 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__3555_
timestamp 1728341909
transform -1 0 8570 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3556_
timestamp 1728341909
transform 1 0 8470 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3557_
timestamp 1728341909
transform -1 0 8130 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__3558_
timestamp 1728341909
transform -1 0 7770 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3559_
timestamp 1728341909
transform 1 0 7730 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3560_
timestamp 1728341909
transform 1 0 8250 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3561_
timestamp 1728341909
transform -1 0 7990 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3562_
timestamp 1728341909
transform -1 0 8990 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3563_
timestamp 1728341909
transform -1 0 8970 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__3564_
timestamp 1728341909
transform 1 0 10070 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__3565_
timestamp 1728341909
transform -1 0 9990 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__3566_
timestamp 1728341909
transform 1 0 9910 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3567_
timestamp 1728341909
transform 1 0 9990 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__3568_
timestamp 1728341909
transform 1 0 10210 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__3569_
timestamp 1728341909
transform 1 0 10210 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__3570_
timestamp 1728341909
transform 1 0 10670 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__3571_
timestamp 1728341909
transform -1 0 10650 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3572_
timestamp 1728341909
transform -1 0 11150 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3573_
timestamp 1728341909
transform 1 0 11030 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__3574_
timestamp 1728341909
transform 1 0 10770 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__3575_
timestamp 1728341909
transform 1 0 11170 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__3576_
timestamp 1728341909
transform 1 0 9950 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__3577_
timestamp 1728341909
transform -1 0 11190 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__3578_
timestamp 1728341909
transform 1 0 10790 0 -1 9850
box -12 -8 32 252
use FILL  FILL_3__3579_
timestamp 1728341909
transform -1 0 10490 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__3580_
timestamp 1728341909
transform -1 0 9190 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3581_
timestamp 1728341909
transform -1 0 8890 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__3582_
timestamp 1728341909
transform 1 0 8730 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__3583_
timestamp 1728341909
transform -1 0 9050 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__3584_
timestamp 1728341909
transform 1 0 8790 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__3585_
timestamp 1728341909
transform -1 0 9530 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__3586_
timestamp 1728341909
transform 1 0 9110 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__3587_
timestamp 1728341909
transform -1 0 9250 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__3588_
timestamp 1728341909
transform 1 0 9270 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__3589_
timestamp 1728341909
transform 1 0 9990 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__3590_
timestamp 1728341909
transform -1 0 10250 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__3591_
timestamp 1728341909
transform 1 0 9730 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__3592_
timestamp 1728341909
transform 1 0 9750 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__3593_
timestamp 1728341909
transform -1 0 9530 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__3594_
timestamp 1728341909
transform 1 0 10370 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3595_
timestamp 1728341909
transform 1 0 10930 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__3596_
timestamp 1728341909
transform -1 0 10890 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3597_
timestamp 1728341909
transform 1 0 10530 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__3598_
timestamp 1728341909
transform 1 0 11170 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__3599_
timestamp 1728341909
transform 1 0 11130 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3600_
timestamp 1728341909
transform 1 0 11010 0 -1 9370
box -12 -8 32 252
use FILL  FILL_3__3601_
timestamp 1728341909
transform 1 0 10190 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3602_
timestamp 1728341909
transform 1 0 10430 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3603_
timestamp 1728341909
transform 1 0 10490 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3604_
timestamp 1728341909
transform 1 0 10710 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3605_
timestamp 1728341909
transform 1 0 11190 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3606_
timestamp 1728341909
transform 1 0 10670 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3607_
timestamp 1728341909
transform -1 0 9970 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3608_
timestamp 1728341909
transform -1 0 10210 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3609_
timestamp 1728341909
transform 1 0 10710 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3610_
timestamp 1728341909
transform 1 0 9530 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3611_
timestamp 1728341909
transform 1 0 9330 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__3612_
timestamp 1728341909
transform 1 0 9590 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__3613_
timestamp 1728341909
transform 1 0 9450 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3614_
timestamp 1728341909
transform -1 0 9850 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__3615_
timestamp 1728341909
transform -1 0 9730 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3616_
timestamp 1728341909
transform -1 0 9030 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3617_
timestamp 1728341909
transform -1 0 9290 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3618_
timestamp 1728341909
transform 1 0 9770 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3619_
timestamp 1728341909
transform 1 0 10930 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3620_
timestamp 1728341909
transform -1 0 10670 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3621_
timestamp 1728341909
transform -1 0 10450 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3622_
timestamp 1728341909
transform 1 0 10690 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3623_
timestamp 1728341909
transform 1 0 9990 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3624_
timestamp 1728341909
transform 1 0 10710 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3625_
timestamp 1728341909
transform 1 0 10810 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__3626_
timestamp 1728341909
transform -1 0 10710 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3627_
timestamp 1728341909
transform -1 0 9690 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3628_
timestamp 1728341909
transform -1 0 10430 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3629_
timestamp 1728341909
transform 1 0 10650 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3630_
timestamp 1728341909
transform 1 0 10450 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3631_
timestamp 1728341909
transform -1 0 10610 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__3632_
timestamp 1728341909
transform -1 0 10950 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__3633_
timestamp 1728341909
transform 1 0 10910 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__3634_
timestamp 1728341909
transform -1 0 10730 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__3635_
timestamp 1728341909
transform -1 0 10450 0 1 10810
box -12 -8 32 252
use FILL  FILL_3__3636_
timestamp 1728341909
transform -1 0 10550 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__3637_
timestamp 1728341909
transform -1 0 10710 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__3638_
timestamp 1728341909
transform -1 0 10630 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3639_
timestamp 1728341909
transform -1 0 10470 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__3640_
timestamp 1728341909
transform -1 0 10930 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3641_
timestamp 1728341909
transform -1 0 10670 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3642_
timestamp 1728341909
transform -1 0 10990 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3643_
timestamp 1728341909
transform 1 0 10910 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3644_
timestamp 1728341909
transform -1 0 10470 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3645_
timestamp 1728341909
transform -1 0 10210 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3646_
timestamp 1728341909
transform -1 0 10970 0 -1 8890
box -12 -8 32 252
use FILL  FILL_3__3647_
timestamp 1728341909
transform 1 0 11070 0 1 250
box -12 -8 32 252
use FILL  FILL_3__3648_
timestamp 1728341909
transform 1 0 11150 0 1 8410
box -12 -8 32 252
use FILL  FILL_3__3649_
timestamp 1728341909
transform 1 0 10230 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3650_
timestamp 1728341909
transform 1 0 10350 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__3651_
timestamp 1728341909
transform 1 0 10450 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3652_
timestamp 1728341909
transform -1 0 10410 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3653_
timestamp 1728341909
transform 1 0 10630 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3654_
timestamp 1728341909
transform 1 0 8430 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3655_
timestamp 1728341909
transform -1 0 8690 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3656_
timestamp 1728341909
transform 1 0 8270 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__3657_
timestamp 1728341909
transform -1 0 8650 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__3658_
timestamp 1728341909
transform -1 0 8550 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__3659_
timestamp 1728341909
transform -1 0 8290 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3__3660_
timestamp 1728341909
transform -1 0 8410 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__3661_
timestamp 1728341909
transform -1 0 9270 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__3662_
timestamp 1728341909
transform -1 0 9510 0 1 10330
box -12 -8 32 252
use FILL  FILL_3__3663_
timestamp 1728341909
transform 1 0 9430 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3664_
timestamp 1728341909
transform -1 0 9670 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3665_
timestamp 1728341909
transform 1 0 8270 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3666_
timestamp 1728341909
transform -1 0 8510 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3667_
timestamp 1728341909
transform -1 0 9230 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3668_
timestamp 1728341909
transform -1 0 10450 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3669_
timestamp 1728341909
transform -1 0 10190 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3670_
timestamp 1728341909
transform -1 0 9950 0 1 9370
box -12 -8 32 252
use FILL  FILL_3__3671_
timestamp 1728341909
transform 1 0 8310 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3672_
timestamp 1728341909
transform 1 0 8550 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3673_
timestamp 1728341909
transform -1 0 9470 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3674_
timestamp 1728341909
transform -1 0 9930 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3675_
timestamp 1728341909
transform 1 0 10150 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3676_
timestamp 1728341909
transform -1 0 10190 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3677_
timestamp 1728341909
transform 1 0 9430 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3678_
timestamp 1728341909
transform -1 0 9270 0 -1 6970
box -12 -8 32 252
use FILL  FILL_3__3691_
timestamp 1728341909
transform 1 0 7750 0 1 250
box -12 -8 32 252
use FILL  FILL_3__3692_
timestamp 1728341909
transform -1 0 8010 0 1 250
box -12 -8 32 252
use FILL  FILL_3__3693_
timestamp 1728341909
transform -1 0 1990 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3694_
timestamp 1728341909
transform -1 0 90 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3695_
timestamp 1728341909
transform 1 0 590 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3696_
timestamp 1728341909
transform -1 0 90 0 1 9850
box -12 -8 32 252
use FILL  FILL_3__3697_
timestamp 1728341909
transform -1 0 90 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__3698_
timestamp 1728341909
transform -1 0 330 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3__3699_
timestamp 1728341909
transform 1 0 6150 0 1 1210
box -12 -8 32 252
use FILL  FILL_3__3700_
timestamp 1728341909
transform -1 0 6310 0 -1 730
box -12 -8 32 252
use FILL  FILL_3__3701_
timestamp 1728341909
transform -1 0 6290 0 1 250
box -12 -8 32 252
use FILL  FILL_3__3702_
timestamp 1728341909
transform -1 0 5270 0 1 5050
box -12 -8 32 252
use FILL  FILL_3__3703_
timestamp 1728341909
transform -1 0 3510 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__3704_
timestamp 1728341909
transform -1 0 3290 0 -1 250
box -12 -8 32 252
use FILL  FILL_3__3705_
timestamp 1728341909
transform -1 0 90 0 1 8890
box -12 -8 32 252
use FILL  FILL_3__3706_
timestamp 1728341909
transform -1 0 1330 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3__3707_
timestamp 1728341909
transform 1 0 11150 0 1 6970
box -12 -8 32 252
use FILL  FILL_3__3708_
timestamp 1728341909
transform 1 0 11150 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3__3709_
timestamp 1728341909
transform 1 0 11170 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3710_
timestamp 1728341909
transform 1 0 10930 0 1 7450
box -12 -8 32 252
use FILL  FILL_3__3711_
timestamp 1728341909
transform 1 0 11150 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3__3712_
timestamp 1728341909
transform 1 0 10930 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3713_
timestamp 1728341909
transform 1 0 11050 0 1 7930
box -12 -8 32 252
use FILL  FILL_3__3714_
timestamp 1728341909
transform 1 0 11170 0 -1 8410
box -12 -8 32 252
use FILL  FILL_3__3715_
timestamp 1728341909
transform 1 0 11150 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert0
timestamp 1728341909
transform 1 0 7790 0 1 10810
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert1
timestamp 1728341909
transform 1 0 9010 0 1 1690
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert2
timestamp 1728341909
transform 1 0 9210 0 1 6970
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert3
timestamp 1728341909
transform 1 0 5690 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert4
timestamp 1728341909
transform 1 0 6790 0 1 1690
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert5
timestamp 1728341909
transform -1 0 4050 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert6
timestamp 1728341909
transform 1 0 7210 0 1 10330
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert7
timestamp 1728341909
transform -1 0 4130 0 1 4090
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert8
timestamp 1728341909
transform -1 0 7570 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert9
timestamp 1728341909
transform 1 0 4490 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert10
timestamp 1728341909
transform -1 0 610 0 1 4090
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert11
timestamp 1728341909
transform -1 0 4810 0 1 2650
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert12
timestamp 1728341909
transform 1 0 770 0 1 5530
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert13
timestamp 1728341909
transform -1 0 5910 0 1 7450
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert14
timestamp 1728341909
transform 1 0 4550 0 1 2650
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert15
timestamp 1728341909
transform 1 0 5630 0 -1 5050
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert16
timestamp 1728341909
transform 1 0 2710 0 1 8410
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert17
timestamp 1728341909
transform 1 0 4210 0 1 6490
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert18
timestamp 1728341909
transform -1 0 90 0 1 2650
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert19
timestamp 1728341909
transform -1 0 350 0 1 8410
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert20
timestamp 1728341909
transform 1 0 550 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert21
timestamp 1728341909
transform -1 0 7090 0 1 4570
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert22
timestamp 1728341909
transform -1 0 10470 0 1 4090
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert23
timestamp 1728341909
transform -1 0 8810 0 1 4090
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert24
timestamp 1728341909
transform 1 0 8530 0 1 3130
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert25
timestamp 1728341909
transform -1 0 7090 0 1 3130
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert37
timestamp 1728341909
transform -1 0 1010 0 1 5530
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert38
timestamp 1728341909
transform 1 0 1290 0 1 4570
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert39
timestamp 1728341909
transform -1 0 1050 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert40
timestamp 1728341909
transform -1 0 2750 0 -1 6010
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert41
timestamp 1728341909
transform 1 0 9550 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert42
timestamp 1728341909
transform 1 0 8870 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert43
timestamp 1728341909
transform -1 0 8790 0 -1 3610
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert44
timestamp 1728341909
transform -1 0 9010 0 1 4570
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert45
timestamp 1728341909
transform 1 0 3870 0 1 4090
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert46
timestamp 1728341909
transform 1 0 5230 0 1 4090
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert47
timestamp 1728341909
transform 1 0 4330 0 1 2650
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert48
timestamp 1728341909
transform 1 0 5450 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert49
timestamp 1728341909
transform -1 0 2250 0 1 2650
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert50
timestamp 1728341909
transform 1 0 8330 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert51
timestamp 1728341909
transform -1 0 10430 0 1 4570
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert52
timestamp 1728341909
transform -1 0 9470 0 1 4570
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert53
timestamp 1728341909
transform -1 0 9550 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert54
timestamp 1728341909
transform -1 0 8390 0 -1 3130
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert55
timestamp 1728341909
transform -1 0 350 0 1 730
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert56
timestamp 1728341909
transform 1 0 5030 0 -1 1210
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert57
timestamp 1728341909
transform 1 0 4630 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert58
timestamp 1728341909
transform 1 0 1950 0 1 1690
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert59
timestamp 1728341909
transform 1 0 4390 0 1 730
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert60
timestamp 1728341909
transform -1 0 8770 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert61
timestamp 1728341909
transform 1 0 10170 0 -1 7450
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert62
timestamp 1728341909
transform 1 0 9210 0 -1 10330
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert63
timestamp 1728341909
transform 1 0 9290 0 1 7450
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert64
timestamp 1728341909
transform 1 0 8630 0 1 1210
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert65
timestamp 1728341909
transform -1 0 5030 0 1 4090
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert66
timestamp 1728341909
transform 1 0 5770 0 1 2650
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert67
timestamp 1728341909
transform 1 0 6610 0 1 5050
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert68
timestamp 1728341909
transform 1 0 7610 0 -1 2650
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert69
timestamp 1728341909
transform -1 0 6090 0 1 1690
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert70
timestamp 1728341909
transform 1 0 8770 0 -1 2170
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert71
timestamp 1728341909
transform 1 0 2470 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert72
timestamp 1728341909
transform 1 0 3910 0 1 1210
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert73
timestamp 1728341909
transform 1 0 2710 0 1 2650
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert74
timestamp 1728341909
transform -1 0 3710 0 -1 1690
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert75
timestamp 1728341909
transform -1 0 790 0 1 2170
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert76
timestamp 1728341909
transform 1 0 8770 0 1 4570
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert77
timestamp 1728341909
transform -1 0 8510 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert78
timestamp 1728341909
transform 1 0 8970 0 -1 5530
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert79
timestamp 1728341909
transform -1 0 9230 0 1 4570
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert80
timestamp 1728341909
transform 1 0 4210 0 -1 6490
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert81
timestamp 1728341909
transform 1 0 3350 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert82
timestamp 1728341909
transform 1 0 2210 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3_BUFX2_insert83
timestamp 1728341909
transform -1 0 2690 0 -1 7930
box -12 -8 32 252
use FILL  FILL_3_CLKBUF1_insert26
timestamp 1728341909
transform -1 0 1430 0 1 3130
box -12 -8 32 252
use FILL  FILL_3_CLKBUF1_insert27
timestamp 1728341909
transform 1 0 3670 0 1 3130
box -12 -8 32 252
use FILL  FILL_3_CLKBUF1_insert28
timestamp 1728341909
transform 1 0 70 0 1 3130
box -12 -8 32 252
use FILL  FILL_3_CLKBUF1_insert29
timestamp 1728341909
transform 1 0 550 0 1 7930
box -12 -8 32 252
use FILL  FILL_3_CLKBUF1_insert30
timestamp 1728341909
transform 1 0 8230 0 1 5530
box -12 -8 32 252
use FILL  FILL_3_CLKBUF1_insert31
timestamp 1728341909
transform -1 0 7590 0 -1 10810
box -12 -8 32 252
use FILL  FILL_3_CLKBUF1_insert32
timestamp 1728341909
transform -1 0 3210 0 -1 4570
box -12 -8 32 252
use FILL  FILL_3_CLKBUF1_insert33
timestamp 1728341909
transform -1 0 7950 0 1 10330
box -12 -8 32 252
use FILL  FILL_3_CLKBUF1_insert34
timestamp 1728341909
transform -1 0 90 0 -1 11290
box -12 -8 32 252
use FILL  FILL_3_CLKBUF1_insert35
timestamp 1728341909
transform -1 0 5510 0 1 5050
box -12 -8 32 252
use FILL  FILL_3_CLKBUF1_insert36
timestamp 1728341909
transform -1 0 2890 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__1744_
timestamp 1728341909
transform -1 0 4490 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__1745_
timestamp 1728341909
transform 1 0 4270 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__1746_
timestamp 1728341909
transform -1 0 4250 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__1747_
timestamp 1728341909
transform -1 0 5710 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__1748_
timestamp 1728341909
transform 1 0 6630 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__1749_
timestamp 1728341909
transform 1 0 6390 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__1750_
timestamp 1728341909
transform 1 0 5230 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__1751_
timestamp 1728341909
transform 1 0 6870 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__1752_
timestamp 1728341909
transform 1 0 5450 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__1753_
timestamp 1728341909
transform 1 0 7590 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__1754_
timestamp 1728341909
transform -1 0 7130 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__1755_
timestamp 1728341909
transform -1 0 7350 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__1756_
timestamp 1728341909
transform -1 0 6430 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__1757_
timestamp 1728341909
transform 1 0 7090 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__1758_
timestamp 1728341909
transform 1 0 6850 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__1759_
timestamp 1728341909
transform -1 0 3110 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__1760_
timestamp 1728341909
transform 1 0 2410 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__1761_
timestamp 1728341909
transform 1 0 7330 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__1762_
timestamp 1728341909
transform 1 0 2610 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__1763_
timestamp 1728341909
transform -1 0 8250 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__1764_
timestamp 1728341909
transform -1 0 8070 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__1765_
timestamp 1728341909
transform -1 0 8070 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__1766_
timestamp 1728341909
transform -1 0 7870 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__1767_
timestamp 1728341909
transform -1 0 7870 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__1768_
timestamp 1728341909
transform -1 0 5750 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__1769_
timestamp 1728341909
transform 1 0 3190 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__1770_
timestamp 1728341909
transform 1 0 10850 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__1771_
timestamp 1728341909
transform 1 0 11090 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__1772_
timestamp 1728341909
transform 1 0 10830 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__1773_
timestamp 1728341909
transform 1 0 10370 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__1774_
timestamp 1728341909
transform 1 0 10730 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1775_
timestamp 1728341909
transform -1 0 9550 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__1776_
timestamp 1728341909
transform 1 0 9590 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__1777_
timestamp 1728341909
transform -1 0 8770 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__1778_
timestamp 1728341909
transform -1 0 10970 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__1779_
timestamp 1728341909
transform 1 0 10190 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__1780_
timestamp 1728341909
transform 1 0 10950 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__1781_
timestamp 1728341909
transform -1 0 10970 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__1782_
timestamp 1728341909
transform -1 0 11210 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1783_
timestamp 1728341909
transform -1 0 10010 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1784_
timestamp 1728341909
transform 1 0 10590 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__1785_
timestamp 1728341909
transform 1 0 10930 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__1786_
timestamp 1728341909
transform -1 0 10270 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__1787_
timestamp 1728341909
transform 1 0 9270 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__1788_
timestamp 1728341909
transform 1 0 10550 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__1789_
timestamp 1728341909
transform -1 0 9410 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1790_
timestamp 1728341909
transform -1 0 10770 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1791_
timestamp 1728341909
transform 1 0 10990 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1792_
timestamp 1728341909
transform 1 0 5690 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1793_
timestamp 1728341909
transform 1 0 5410 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1794_
timestamp 1728341909
transform -1 0 4990 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1795_
timestamp 1728341909
transform 1 0 3770 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1796_
timestamp 1728341909
transform 1 0 4230 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1797_
timestamp 1728341909
transform -1 0 4750 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1798_
timestamp 1728341909
transform -1 0 11070 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__1799_
timestamp 1728341909
transform -1 0 10970 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__1800_
timestamp 1728341909
transform -1 0 10490 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__1801_
timestamp 1728341909
transform -1 0 10150 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__1802_
timestamp 1728341909
transform 1 0 10030 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__1803_
timestamp 1728341909
transform 1 0 10270 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1804_
timestamp 1728341909
transform 1 0 10270 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__1805_
timestamp 1728341909
transform -1 0 10070 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__1806_
timestamp 1728341909
transform 1 0 10010 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1807_
timestamp 1728341909
transform -1 0 10130 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1808_
timestamp 1728341909
transform -1 0 10430 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__1809_
timestamp 1728341909
transform -1 0 11090 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1810_
timestamp 1728341909
transform -1 0 6270 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1811_
timestamp 1728341909
transform -1 0 11170 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__1812_
timestamp 1728341909
transform -1 0 10250 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__1813_
timestamp 1728341909
transform -1 0 7730 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__1814_
timestamp 1728341909
transform -1 0 7570 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1815_
timestamp 1728341909
transform -1 0 10990 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1816_
timestamp 1728341909
transform -1 0 7630 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__1817_
timestamp 1728341909
transform 1 0 6750 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__1818_
timestamp 1728341909
transform 1 0 6690 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1819_
timestamp 1728341909
transform 1 0 6190 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1820_
timestamp 1728341909
transform 1 0 10390 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__1821_
timestamp 1728341909
transform -1 0 6750 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1822_
timestamp 1728341909
transform 1 0 11170 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__1823_
timestamp 1728341909
transform -1 0 10030 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__1824_
timestamp 1728341909
transform 1 0 7330 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__1825_
timestamp 1728341909
transform 1 0 6550 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1826_
timestamp 1728341909
transform 1 0 10970 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1827_
timestamp 1728341909
transform -1 0 7410 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1828_
timestamp 1728341909
transform 1 0 11170 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__1829_
timestamp 1728341909
transform -1 0 7430 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__1830_
timestamp 1728341909
transform 1 0 7570 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__1831_
timestamp 1728341909
transform 1 0 10710 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__1832_
timestamp 1728341909
transform 1 0 10690 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__1833_
timestamp 1728341909
transform 1 0 7250 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1834_
timestamp 1728341909
transform -1 0 7050 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1835_
timestamp 1728341909
transform -1 0 6490 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1836_
timestamp 1728341909
transform -1 0 6050 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1837_
timestamp 1728341909
transform -1 0 5570 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1838_
timestamp 1728341909
transform 1 0 5290 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1839_
timestamp 1728341909
transform 1 0 5870 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1840_
timestamp 1728341909
transform -1 0 8070 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__1841_
timestamp 1728341909
transform -1 0 5010 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__1842_
timestamp 1728341909
transform -1 0 6870 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__1843_
timestamp 1728341909
transform 1 0 7190 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__1844_
timestamp 1728341909
transform -1 0 10270 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__1845_
timestamp 1728341909
transform 1 0 11170 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__1846_
timestamp 1728341909
transform 1 0 11190 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1847_
timestamp 1728341909
transform -1 0 8110 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__1848_
timestamp 1728341909
transform 1 0 10710 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__1849_
timestamp 1728341909
transform -1 0 10630 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__1850_
timestamp 1728341909
transform -1 0 8570 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__1851_
timestamp 1728341909
transform -1 0 11190 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__1852_
timestamp 1728341909
transform 1 0 9750 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__1853_
timestamp 1728341909
transform 1 0 9270 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__1854_
timestamp 1728341909
transform 1 0 9070 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__1855_
timestamp 1728341909
transform 1 0 8830 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__1856_
timestamp 1728341909
transform 1 0 9350 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__1857_
timestamp 1728341909
transform 1 0 9130 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__1858_
timestamp 1728341909
transform 1 0 7310 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__1859_
timestamp 1728341909
transform -1 0 10730 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__1860_
timestamp 1728341909
transform 1 0 7110 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__1861_
timestamp 1728341909
transform 1 0 7350 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__1862_
timestamp 1728341909
transform -1 0 9850 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__1863_
timestamp 1728341909
transform 1 0 8590 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__1864_
timestamp 1728341909
transform 1 0 9890 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__1865_
timestamp 1728341909
transform 1 0 7750 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__1866_
timestamp 1728341909
transform -1 0 8930 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1867_
timestamp 1728341909
transform 1 0 9310 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__1868_
timestamp 1728341909
transform 1 0 10870 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__1869_
timestamp 1728341909
transform 1 0 9330 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__1870_
timestamp 1728341909
transform -1 0 9110 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__1871_
timestamp 1728341909
transform 1 0 8550 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__1872_
timestamp 1728341909
transform 1 0 7830 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__1873_
timestamp 1728341909
transform 1 0 6390 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1874_
timestamp 1728341909
transform -1 0 6850 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1875_
timestamp 1728341909
transform -1 0 6610 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1876_
timestamp 1728341909
transform 1 0 6670 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__1877_
timestamp 1728341909
transform -1 0 8090 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__1878_
timestamp 1728341909
transform -1 0 8350 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__1879_
timestamp 1728341909
transform -1 0 8090 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__1880_
timestamp 1728341909
transform -1 0 7030 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__1881_
timestamp 1728341909
transform -1 0 6350 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__1882_
timestamp 1728341909
transform 1 0 3510 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__1883_
timestamp 1728341909
transform -1 0 7050 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__1884_
timestamp 1728341909
transform -1 0 6570 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__1885_
timestamp 1728341909
transform 1 0 5850 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__1886_
timestamp 1728341909
transform -1 0 6250 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__1887_
timestamp 1728341909
transform 1 0 6870 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__1888_
timestamp 1728341909
transform 1 0 3630 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__1889_
timestamp 1728341909
transform -1 0 5990 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__1890_
timestamp 1728341909
transform 1 0 6450 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__1891_
timestamp 1728341909
transform -1 0 6090 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__1892_
timestamp 1728341909
transform 1 0 5650 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__1893_
timestamp 1728341909
transform 1 0 1050 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__1894_
timestamp 1728341909
transform 1 0 5990 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__1895_
timestamp 1728341909
transform 1 0 6870 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__1896_
timestamp 1728341909
transform 1 0 5190 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__1897_
timestamp 1728341909
transform 1 0 6030 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__1898_
timestamp 1728341909
transform 1 0 6450 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__1899_
timestamp 1728341909
transform 1 0 6550 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__1900_
timestamp 1728341909
transform 1 0 570 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__1901_
timestamp 1728341909
transform 1 0 8010 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__1902_
timestamp 1728341909
transform 1 0 8550 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__1903_
timestamp 1728341909
transform 1 0 7910 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__1904_
timestamp 1728341909
transform -1 0 10070 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1905_
timestamp 1728341909
transform 1 0 7570 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__1906_
timestamp 1728341909
transform 1 0 7550 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__1907_
timestamp 1728341909
transform 1 0 8690 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1908_
timestamp 1728341909
transform -1 0 7750 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1909_
timestamp 1728341909
transform 1 0 1850 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1910_
timestamp 1728341909
transform -1 0 9810 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__1911_
timestamp 1728341909
transform 1 0 9530 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1912_
timestamp 1728341909
transform 1 0 6150 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1913_
timestamp 1728341909
transform 1 0 10670 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__1914_
timestamp 1728341909
transform 1 0 10730 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1915_
timestamp 1728341909
transform -1 0 10290 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1916_
timestamp 1728341909
transform -1 0 5910 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1917_
timestamp 1728341909
transform 1 0 4050 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1918_
timestamp 1728341909
transform -1 0 830 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__1919_
timestamp 1728341909
transform -1 0 110 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__1920_
timestamp 1728341909
transform 1 0 1050 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__1921_
timestamp 1728341909
transform -1 0 1230 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1922_
timestamp 1728341909
transform -1 0 970 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1923_
timestamp 1728341909
transform 1 0 570 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__1924_
timestamp 1728341909
transform -1 0 4510 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1925_
timestamp 1728341909
transform -1 0 350 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__1926_
timestamp 1728341909
transform 1 0 810 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__1927_
timestamp 1728341909
transform -1 0 2110 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1928_
timestamp 1728341909
transform -1 0 1630 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1929_
timestamp 1728341909
transform 1 0 310 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__1930_
timestamp 1728341909
transform 1 0 690 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1931_
timestamp 1728341909
transform 1 0 570 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__1932_
timestamp 1728341909
transform -1 0 590 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1933_
timestamp 1728341909
transform 1 0 570 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__1934_
timestamp 1728341909
transform -1 0 590 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1935_
timestamp 1728341909
transform -1 0 1570 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1936_
timestamp 1728341909
transform 1 0 830 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1937_
timestamp 1728341909
transform -1 0 590 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__1938_
timestamp 1728341909
transform -1 0 110 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__1939_
timestamp 1728341909
transform 1 0 330 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__1940_
timestamp 1728341909
transform 1 0 850 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1941_
timestamp 1728341909
transform 1 0 570 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__1942_
timestamp 1728341909
transform 1 0 570 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__1943_
timestamp 1728341909
transform 1 0 8130 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__1944_
timestamp 1728341909
transform -1 0 7670 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1945_
timestamp 1728341909
transform -1 0 7450 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1946_
timestamp 1728341909
transform 1 0 8470 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1947_
timestamp 1728341909
transform -1 0 7650 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1948_
timestamp 1728341909
transform -1 0 6990 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1949_
timestamp 1728341909
transform -1 0 7230 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1950_
timestamp 1728341909
transform 1 0 8330 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__1951_
timestamp 1728341909
transform 1 0 8330 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__1952_
timestamp 1728341909
transform 1 0 9850 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1953_
timestamp 1728341909
transform -1 0 8410 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__1954_
timestamp 1728341909
transform 1 0 8250 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1955_
timestamp 1728341909
transform 1 0 6450 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__1956_
timestamp 1728341909
transform -1 0 8010 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1957_
timestamp 1728341909
transform 1 0 8090 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__1958_
timestamp 1728341909
transform 1 0 10450 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__1959_
timestamp 1728341909
transform 1 0 7810 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__1960_
timestamp 1728341909
transform 1 0 7890 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__1961_
timestamp 1728341909
transform 1 0 10710 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__1962_
timestamp 1728341909
transform 1 0 10510 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__1963_
timestamp 1728341909
transform 1 0 9850 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1964_
timestamp 1728341909
transform -1 0 7390 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__1965_
timestamp 1728341909
transform -1 0 7670 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__1966_
timestamp 1728341909
transform -1 0 3530 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__1967_
timestamp 1728341909
transform -1 0 6990 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__1968_
timestamp 1728341909
transform 1 0 7530 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__1969_
timestamp 1728341909
transform -1 0 7790 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__1970_
timestamp 1728341909
transform 1 0 1530 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__1971_
timestamp 1728341909
transform -1 0 830 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1972_
timestamp 1728341909
transform 1 0 1350 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1973_
timestamp 1728341909
transform 1 0 1610 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__1974_
timestamp 1728341909
transform 1 0 8370 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__1975_
timestamp 1728341909
transform 1 0 2990 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__1976_
timestamp 1728341909
transform -1 0 7150 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__1977_
timestamp 1728341909
transform -1 0 2850 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__1978_
timestamp 1728341909
transform -1 0 3830 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__1979_
timestamp 1728341909
transform -1 0 6530 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__1980_
timestamp 1728341909
transform 1 0 7790 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__1981_
timestamp 1728341909
transform 1 0 8310 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__1982_
timestamp 1728341909
transform -1 0 3050 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__1983_
timestamp 1728341909
transform 1 0 1730 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__1984_
timestamp 1728341909
transform 1 0 1810 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__1985_
timestamp 1728341909
transform 1 0 2470 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__1986_
timestamp 1728341909
transform -1 0 7150 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__1987_
timestamp 1728341909
transform 1 0 5090 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__1988_
timestamp 1728341909
transform -1 0 4990 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__1989_
timestamp 1728341909
transform 1 0 6750 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__1990_
timestamp 1728341909
transform -1 0 7270 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__1991_
timestamp 1728341909
transform -1 0 2070 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__1992_
timestamp 1728341909
transform -1 0 1570 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__1993_
timestamp 1728341909
transform -1 0 1850 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__1994_
timestamp 1728341909
transform 1 0 2090 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__1995_
timestamp 1728341909
transform 1 0 8050 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__1996_
timestamp 1728341909
transform -1 0 2270 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__1997_
timestamp 1728341909
transform -1 0 3990 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__1998_
timestamp 1728341909
transform -1 0 6510 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__1999_
timestamp 1728341909
transform -1 0 8230 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2000_
timestamp 1728341909
transform 1 0 1830 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2001_
timestamp 1728341909
transform 1 0 1310 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2002_
timestamp 1728341909
transform 1 0 1550 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2003_
timestamp 1728341909
transform 1 0 1570 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2004_
timestamp 1728341909
transform 1 0 7850 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2005_
timestamp 1728341909
transform 1 0 2010 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2006_
timestamp 1728341909
transform -1 0 6270 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2007_
timestamp 1728341909
transform 1 0 7550 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2008_
timestamp 1728341909
transform -1 0 8070 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2009_
timestamp 1728341909
transform 1 0 810 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2010_
timestamp 1728341909
transform -1 0 870 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2011_
timestamp 1728341909
transform 1 0 570 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2012_
timestamp 1728341909
transform 1 0 830 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2013_
timestamp 1728341909
transform 1 0 5470 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2014_
timestamp 1728341909
transform 1 0 1770 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2015_
timestamp 1728341909
transform -1 0 3970 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2016_
timestamp 1728341909
transform 1 0 6770 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2017_
timestamp 1728341909
transform -1 0 7310 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2018_
timestamp 1728341909
transform -1 0 1550 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2019_
timestamp 1728341909
transform -1 0 1610 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2020_
timestamp 1728341909
transform 1 0 1790 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2021_
timestamp 1728341909
transform 1 0 1750 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2022_
timestamp 1728341909
transform 1 0 4530 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2023_
timestamp 1728341909
transform 1 0 570 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2024_
timestamp 1728341909
transform 1 0 1470 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2025_
timestamp 1728341909
transform 1 0 2530 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2026_
timestamp 1728341909
transform -1 0 4730 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2027_
timestamp 1728341909
transform 1 0 7230 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2028_
timestamp 1728341909
transform -1 0 7510 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2029_
timestamp 1728341909
transform -1 0 110 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2030_
timestamp 1728341909
transform -1 0 590 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2031_
timestamp 1728341909
transform -1 0 350 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2032_
timestamp 1728341909
transform 1 0 570 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2033_
timestamp 1728341909
transform 1 0 7650 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2034_
timestamp 1728341909
transform 1 0 1250 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2035_
timestamp 1728341909
transform 1 0 2130 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2036_
timestamp 1728341909
transform 1 0 2930 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2037_
timestamp 1728341909
transform -1 0 4130 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2038_
timestamp 1728341909
transform 1 0 7570 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2039_
timestamp 1728341909
transform -1 0 7850 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2040_
timestamp 1728341909
transform -1 0 2970 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2041_
timestamp 1728341909
transform -1 0 590 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2042_
timestamp 1728341909
transform 1 0 1750 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__2043_
timestamp 1728341909
transform -1 0 3850 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__2044_
timestamp 1728341909
transform 1 0 5390 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2045_
timestamp 1728341909
transform -1 0 4090 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2046_
timestamp 1728341909
transform 1 0 2890 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__2047_
timestamp 1728341909
transform 1 0 2650 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__2048_
timestamp 1728341909
transform -1 0 3590 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__2049_
timestamp 1728341909
transform -1 0 2990 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__2050_
timestamp 1728341909
transform -1 0 2470 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__2051_
timestamp 1728341909
transform -1 0 2450 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2052_
timestamp 1728341909
transform -1 0 870 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2053_
timestamp 1728341909
transform -1 0 3430 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__2054_
timestamp 1728341909
transform 1 0 3150 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__2055_
timestamp 1728341909
transform -1 0 2790 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__2056_
timestamp 1728341909
transform 1 0 4410 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2057_
timestamp 1728341909
transform -1 0 3970 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2058_
timestamp 1728341909
transform 1 0 4630 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2059_
timestamp 1728341909
transform -1 0 1990 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__2060_
timestamp 1728341909
transform -1 0 3810 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__2061_
timestamp 1728341909
transform 1 0 3550 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__2062_
timestamp 1728341909
transform -1 0 3570 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__2063_
timestamp 1728341909
transform 1 0 2510 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__2064_
timestamp 1728341909
transform -1 0 2610 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2065_
timestamp 1728341909
transform -1 0 2410 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2066_
timestamp 1728341909
transform 1 0 2470 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2067_
timestamp 1728341909
transform -1 0 2790 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__2068_
timestamp 1728341909
transform -1 0 3030 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__2069_
timestamp 1728341909
transform 1 0 2570 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__2070_
timestamp 1728341909
transform -1 0 1110 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2071_
timestamp 1728341909
transform -1 0 2830 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__2072_
timestamp 1728341909
transform -1 0 2570 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__2073_
timestamp 1728341909
transform -1 0 1310 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2074_
timestamp 1728341909
transform 1 0 3250 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__2075_
timestamp 1728341909
transform -1 0 2730 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__2076_
timestamp 1728341909
transform 1 0 2430 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__2077_
timestamp 1728341909
transform -1 0 3290 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__2078_
timestamp 1728341909
transform 1 0 2810 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__2079_
timestamp 1728341909
transform -1 0 3930 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2080_
timestamp 1728341909
transform 1 0 4150 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2081_
timestamp 1728341909
transform -1 0 3710 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2082_
timestamp 1728341909
transform 1 0 5790 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2083_
timestamp 1728341909
transform -1 0 6530 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2084_
timestamp 1728341909
transform 1 0 9950 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2085_
timestamp 1728341909
transform -1 0 10470 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2086_
timestamp 1728341909
transform 1 0 10490 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2087_
timestamp 1728341909
transform 1 0 11030 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__2088_
timestamp 1728341909
transform 1 0 10230 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2089_
timestamp 1728341909
transform -1 0 9530 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2090_
timestamp 1728341909
transform 1 0 10710 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__2091_
timestamp 1728341909
transform 1 0 11210 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__2092_
timestamp 1728341909
transform -1 0 10170 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2093_
timestamp 1728341909
transform 1 0 10230 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__2094_
timestamp 1728341909
transform -1 0 10730 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__2095_
timestamp 1728341909
transform 1 0 10790 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__2096_
timestamp 1728341909
transform -1 0 11190 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__2097_
timestamp 1728341909
transform -1 0 11130 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2098_
timestamp 1728341909
transform 1 0 10210 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2099_
timestamp 1728341909
transform 1 0 10690 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2100_
timestamp 1728341909
transform 1 0 10910 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2101_
timestamp 1728341909
transform 1 0 11150 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2102_
timestamp 1728341909
transform 1 0 4030 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__2103_
timestamp 1728341909
transform 1 0 4270 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__2104_
timestamp 1728341909
transform 1 0 3890 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2105_
timestamp 1728341909
transform -1 0 1790 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2106_
timestamp 1728341909
transform -1 0 2170 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2107_
timestamp 1728341909
transform -1 0 2690 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2108_
timestamp 1728341909
transform 1 0 1490 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2109_
timestamp 1728341909
transform -1 0 2910 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2110_
timestamp 1728341909
transform 1 0 3130 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2111_
timestamp 1728341909
transform 1 0 5330 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2112_
timestamp 1728341909
transform 1 0 11210 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__2113_
timestamp 1728341909
transform -1 0 9790 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__2114_
timestamp 1728341909
transform 1 0 9790 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2115_
timestamp 1728341909
transform -1 0 11110 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2116_
timestamp 1728341909
transform -1 0 11050 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__2117_
timestamp 1728341909
transform -1 0 10650 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__2118_
timestamp 1728341909
transform 1 0 9050 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__2119_
timestamp 1728341909
transform -1 0 11130 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__2120_
timestamp 1728341909
transform 1 0 11070 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2121_
timestamp 1728341909
transform 1 0 11170 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2122_
timestamp 1728341909
transform 1 0 10870 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2123_
timestamp 1728341909
transform 1 0 10930 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2124_
timestamp 1728341909
transform 1 0 9390 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2125_
timestamp 1728341909
transform 1 0 9510 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2126_
timestamp 1728341909
transform -1 0 9950 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2127_
timestamp 1728341909
transform 1 0 9770 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2128_
timestamp 1728341909
transform 1 0 9730 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2129_
timestamp 1728341909
transform -1 0 8950 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2130_
timestamp 1728341909
transform 1 0 9630 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2131_
timestamp 1728341909
transform 1 0 9730 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2132_
timestamp 1728341909
transform 1 0 10190 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2133_
timestamp 1728341909
transform 1 0 10350 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2134_
timestamp 1728341909
transform -1 0 10130 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2135_
timestamp 1728341909
transform 1 0 10630 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2136_
timestamp 1728341909
transform -1 0 10590 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2137_
timestamp 1728341909
transform 1 0 10830 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2138_
timestamp 1728341909
transform -1 0 10930 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2139_
timestamp 1728341909
transform -1 0 10870 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2140_
timestamp 1728341909
transform -1 0 8350 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2141_
timestamp 1728341909
transform 1 0 8590 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2142_
timestamp 1728341909
transform 1 0 1910 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2143_
timestamp 1728341909
transform -1 0 2950 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2144_
timestamp 1728341909
transform -1 0 6050 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2145_
timestamp 1728341909
transform -1 0 6250 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2146_
timestamp 1728341909
transform 1 0 5550 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2147_
timestamp 1728341909
transform -1 0 6790 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2148_
timestamp 1728341909
transform 1 0 9690 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2149_
timestamp 1728341909
transform 1 0 8770 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2150_
timestamp 1728341909
transform -1 0 8530 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2151_
timestamp 1728341909
transform 1 0 8190 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2152_
timestamp 1728341909
transform -1 0 9030 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2153_
timestamp 1728341909
transform -1 0 9130 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2154_
timestamp 1728341909
transform 1 0 8870 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__2155_
timestamp 1728341909
transform 1 0 8030 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__2156_
timestamp 1728341909
transform -1 0 8310 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__2157_
timestamp 1728341909
transform -1 0 8430 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2158_
timestamp 1728341909
transform 1 0 10350 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__2159_
timestamp 1728341909
transform 1 0 6050 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2160_
timestamp 1728341909
transform -1 0 6410 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2161_
timestamp 1728341909
transform 1 0 6610 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2162_
timestamp 1728341909
transform -1 0 7950 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2163_
timestamp 1728341909
transform -1 0 8370 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__2164_
timestamp 1728341909
transform 1 0 7130 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2165_
timestamp 1728341909
transform -1 0 7110 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2166_
timestamp 1728341909
transform -1 0 8170 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2167_
timestamp 1728341909
transform -1 0 7870 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2168_
timestamp 1728341909
transform -1 0 8130 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2169_
timestamp 1728341909
transform 1 0 8170 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2170_
timestamp 1728341909
transform -1 0 8390 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2171_
timestamp 1728341909
transform 1 0 8590 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2172_
timestamp 1728341909
transform -1 0 10450 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2173_
timestamp 1728341909
transform 1 0 10190 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2174_
timestamp 1728341909
transform 1 0 4410 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2175_
timestamp 1728341909
transform -1 0 3970 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2176_
timestamp 1728341909
transform -1 0 5430 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2177_
timestamp 1728341909
transform -1 0 6090 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2178_
timestamp 1728341909
transform -1 0 6350 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2179_
timestamp 1728341909
transform 1 0 6390 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2180_
timestamp 1728341909
transform 1 0 7190 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2181_
timestamp 1728341909
transform 1 0 7330 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__2182_
timestamp 1728341909
transform -1 0 7190 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__2183_
timestamp 1728341909
transform 1 0 6170 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2184_
timestamp 1728341909
transform 1 0 6490 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2185_
timestamp 1728341909
transform -1 0 6630 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2186_
timestamp 1728341909
transform -1 0 9070 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2187_
timestamp 1728341909
transform -1 0 9470 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2188_
timestamp 1728341909
transform 1 0 9070 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2189_
timestamp 1728341909
transform -1 0 8850 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2190_
timestamp 1728341909
transform 1 0 8530 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2191_
timestamp 1728341909
transform 1 0 8770 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2192_
timestamp 1728341909
transform 1 0 7330 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2193_
timestamp 1728341909
transform 1 0 7550 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2194_
timestamp 1728341909
transform -1 0 8670 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__2195_
timestamp 1728341909
transform -1 0 8590 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__2196_
timestamp 1728341909
transform 1 0 8630 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2197_
timestamp 1728341909
transform 1 0 8670 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2198_
timestamp 1728341909
transform -1 0 7270 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2199_
timestamp 1728341909
transform -1 0 7530 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2200_
timestamp 1728341909
transform 1 0 9050 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__2201_
timestamp 1728341909
transform 1 0 8910 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2202_
timestamp 1728341909
transform -1 0 8710 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2203_
timestamp 1728341909
transform 1 0 8430 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2204_
timestamp 1728341909
transform -1 0 8430 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2205_
timestamp 1728341909
transform 1 0 8170 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2206_
timestamp 1728341909
transform -1 0 8050 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2207_
timestamp 1728341909
transform 1 0 8550 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2208_
timestamp 1728341909
transform -1 0 8310 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2209_
timestamp 1728341909
transform -1 0 7830 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2210_
timestamp 1728341909
transform 1 0 2770 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2211_
timestamp 1728341909
transform -1 0 7230 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2212_
timestamp 1728341909
transform -1 0 7490 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2213_
timestamp 1728341909
transform -1 0 8010 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2214_
timestamp 1728341909
transform 1 0 8570 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2215_
timestamp 1728341909
transform 1 0 9270 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2216_
timestamp 1728341909
transform 1 0 9250 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2217_
timestamp 1728341909
transform -1 0 9510 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2218_
timestamp 1728341909
transform 1 0 3950 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2219_
timestamp 1728341909
transform -1 0 2270 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__2220_
timestamp 1728341909
transform -1 0 3690 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2221_
timestamp 1728341909
transform 1 0 4130 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2222_
timestamp 1728341909
transform 1 0 4350 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2223_
timestamp 1728341909
transform 1 0 4170 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2224_
timestamp 1728341909
transform -1 0 2850 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2225_
timestamp 1728341909
transform -1 0 5910 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2226_
timestamp 1728341909
transform 1 0 6030 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2227_
timestamp 1728341909
transform -1 0 7010 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2228_
timestamp 1728341909
transform 1 0 6750 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2229_
timestamp 1728341909
transform 1 0 7810 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__2230_
timestamp 1728341909
transform -1 0 6210 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__2231_
timestamp 1728341909
transform -1 0 6450 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__2232_
timestamp 1728341909
transform 1 0 6870 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2233_
timestamp 1728341909
transform 1 0 7450 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2234_
timestamp 1728341909
transform 1 0 7350 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2235_
timestamp 1728341909
transform 1 0 9430 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2236_
timestamp 1728341909
transform 1 0 10490 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2237_
timestamp 1728341909
transform 1 0 9970 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2238_
timestamp 1728341909
transform -1 0 9890 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2239_
timestamp 1728341909
transform -1 0 5850 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2240_
timestamp 1728341909
transform 1 0 2710 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2241_
timestamp 1728341909
transform -1 0 4390 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2242_
timestamp 1728341909
transform -1 0 4610 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2243_
timestamp 1728341909
transform 1 0 3390 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2244_
timestamp 1728341909
transform 1 0 5150 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2245_
timestamp 1728341909
transform 1 0 7290 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2246_
timestamp 1728341909
transform 1 0 7310 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2247_
timestamp 1728341909
transform -1 0 3270 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2248_
timestamp 1728341909
transform 1 0 3450 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2249_
timestamp 1728341909
transform 1 0 5430 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2250_
timestamp 1728341909
transform 1 0 6690 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2251_
timestamp 1728341909
transform 1 0 7210 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2252_
timestamp 1728341909
transform -1 0 9650 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__2253_
timestamp 1728341909
transform 1 0 9370 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2254_
timestamp 1728341909
transform 1 0 5650 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2255_
timestamp 1728341909
transform -1 0 6990 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2256_
timestamp 1728341909
transform 1 0 7150 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2257_
timestamp 1728341909
transform -1 0 3090 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2258_
timestamp 1728341909
transform -1 0 3050 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__2259_
timestamp 1728341909
transform 1 0 3470 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2260_
timestamp 1728341909
transform 1 0 4650 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2261_
timestamp 1728341909
transform -1 0 5650 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2262_
timestamp 1728341909
transform 1 0 4830 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2263_
timestamp 1728341909
transform 1 0 4890 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2264_
timestamp 1728341909
transform -1 0 6190 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2265_
timestamp 1728341909
transform 1 0 3490 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__2266_
timestamp 1728341909
transform 1 0 7530 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__2267_
timestamp 1728341909
transform -1 0 5430 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__2268_
timestamp 1728341909
transform -1 0 5670 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__2269_
timestamp 1728341909
transform 1 0 5430 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__2270_
timestamp 1728341909
transform -1 0 6270 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__2271_
timestamp 1728341909
transform 1 0 5990 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__2272_
timestamp 1728341909
transform 1 0 5590 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__2273_
timestamp 1728341909
transform 1 0 5410 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__2274_
timestamp 1728341909
transform 1 0 5170 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__2275_
timestamp 1728341909
transform 1 0 5650 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__2276_
timestamp 1728341909
transform -1 0 6290 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2277_
timestamp 1728341909
transform 1 0 7790 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__2278_
timestamp 1728341909
transform -1 0 7730 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2279_
timestamp 1728341909
transform 1 0 6490 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2280_
timestamp 1728341909
transform -1 0 6510 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2281_
timestamp 1728341909
transform -1 0 6270 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2282_
timestamp 1728341909
transform 1 0 6550 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2283_
timestamp 1728341909
transform 1 0 7250 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2284_
timestamp 1728341909
transform 1 0 9210 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2285_
timestamp 1728341909
transform 1 0 9650 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2286_
timestamp 1728341909
transform -1 0 2550 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__2287_
timestamp 1728341909
transform -1 0 1810 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2288_
timestamp 1728341909
transform -1 0 2250 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2289_
timestamp 1728341909
transform 1 0 2210 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2290_
timestamp 1728341909
transform -1 0 1770 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2291_
timestamp 1728341909
transform 1 0 1990 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2292_
timestamp 1728341909
transform 1 0 4110 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2293_
timestamp 1728341909
transform 1 0 4850 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2294_
timestamp 1728341909
transform 1 0 6070 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2295_
timestamp 1728341909
transform -1 0 2250 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2296_
timestamp 1728341909
transform 1 0 3690 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2297_
timestamp 1728341909
transform 1 0 2230 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2298_
timestamp 1728341909
transform 1 0 1990 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2299_
timestamp 1728341909
transform 1 0 3450 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2300_
timestamp 1728341909
transform 1 0 3190 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2301_
timestamp 1728341909
transform -1 0 3650 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2302_
timestamp 1728341909
transform 1 0 5130 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2303_
timestamp 1728341909
transform -1 0 5110 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2304_
timestamp 1728341909
transform 1 0 5350 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2305_
timestamp 1728341909
transform -1 0 1550 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2306_
timestamp 1728341909
transform 1 0 2450 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2307_
timestamp 1728341909
transform -1 0 5610 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2308_
timestamp 1728341909
transform -1 0 5610 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2309_
timestamp 1728341909
transform 1 0 4610 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2310_
timestamp 1728341909
transform 1 0 4370 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2311_
timestamp 1728341909
transform -1 0 3770 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2312_
timestamp 1728341909
transform -1 0 4010 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2313_
timestamp 1728341909
transform 1 0 5290 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2314_
timestamp 1728341909
transform 1 0 4470 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2315_
timestamp 1728341909
transform 1 0 5430 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2316_
timestamp 1728341909
transform -1 0 9870 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2317_
timestamp 1728341909
transform 1 0 11170 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2318_
timestamp 1728341909
transform -1 0 10870 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__2319_
timestamp 1728341909
transform -1 0 10490 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__2320_
timestamp 1728341909
transform 1 0 10650 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2321_
timestamp 1728341909
transform 1 0 10590 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__2322_
timestamp 1728341909
transform 1 0 10490 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__2323_
timestamp 1728341909
transform 1 0 6750 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2324_
timestamp 1728341909
transform 1 0 6950 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2325_
timestamp 1728341909
transform 1 0 9310 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2326_
timestamp 1728341909
transform -1 0 8850 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2327_
timestamp 1728341909
transform -1 0 9310 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2328_
timestamp 1728341909
transform -1 0 9550 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2329_
timestamp 1728341909
transform 1 0 9270 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2330_
timestamp 1728341909
transform -1 0 9030 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2331_
timestamp 1728341909
transform -1 0 9190 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2332_
timestamp 1728341909
transform 1 0 9170 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2333_
timestamp 1728341909
transform 1 0 9430 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2334_
timestamp 1728341909
transform -1 0 9630 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2335_
timestamp 1728341909
transform 1 0 5670 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2336_
timestamp 1728341909
transform 1 0 6190 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2337_
timestamp 1728341909
transform -1 0 5970 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2338_
timestamp 1728341909
transform -1 0 5910 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2339_
timestamp 1728341909
transform 1 0 10390 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2340_
timestamp 1728341909
transform -1 0 9270 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2341_
timestamp 1728341909
transform 1 0 9270 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2342_
timestamp 1728341909
transform 1 0 10130 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2343_
timestamp 1728341909
transform -1 0 9630 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2344_
timestamp 1728341909
transform 1 0 9730 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2345_
timestamp 1728341909
transform -1 0 6910 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2346_
timestamp 1728341909
transform 1 0 6770 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2347_
timestamp 1728341909
transform -1 0 7110 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2348_
timestamp 1728341909
transform 1 0 8110 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2349_
timestamp 1728341909
transform -1 0 7810 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2350_
timestamp 1728341909
transform 1 0 7530 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2351_
timestamp 1728341909
transform -1 0 5230 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2352_
timestamp 1728341909
transform 1 0 5830 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2353_
timestamp 1728341909
transform -1 0 4250 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2354_
timestamp 1728341909
transform 1 0 4730 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2355_
timestamp 1728341909
transform -1 0 4990 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2356_
timestamp 1728341909
transform 1 0 5930 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2357_
timestamp 1728341909
transform -1 0 5690 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2358_
timestamp 1728341909
transform 1 0 6970 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2359_
timestamp 1728341909
transform 1 0 6330 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2360_
timestamp 1728341909
transform 1 0 6570 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2361_
timestamp 1728341909
transform 1 0 7870 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__2362_
timestamp 1728341909
transform 1 0 7390 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2363_
timestamp 1728341909
transform -1 0 7490 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2364_
timestamp 1728341909
transform 1 0 8110 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__2365_
timestamp 1728341909
transform -1 0 7990 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2366_
timestamp 1728341909
transform 1 0 7750 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2367_
timestamp 1728341909
transform 1 0 8030 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2368_
timestamp 1728341909
transform 1 0 8250 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2369_
timestamp 1728341909
transform -1 0 9970 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2370_
timestamp 1728341909
transform 1 0 5390 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2371_
timestamp 1728341909
transform -1 0 8790 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2372_
timestamp 1728341909
transform -1 0 8530 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2373_
timestamp 1728341909
transform -1 0 8110 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2374_
timestamp 1728341909
transform 1 0 8110 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2375_
timestamp 1728341909
transform 1 0 6510 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2376_
timestamp 1728341909
transform 1 0 8470 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2377_
timestamp 1728341909
transform -1 0 8730 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2378_
timestamp 1728341909
transform -1 0 9030 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2379_
timestamp 1728341909
transform -1 0 6890 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2380_
timestamp 1728341909
transform -1 0 7030 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2381_
timestamp 1728341909
transform -1 0 6890 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2382_
timestamp 1728341909
transform -1 0 7970 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2383_
timestamp 1728341909
transform 1 0 7690 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2384_
timestamp 1728341909
transform 1 0 7790 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2385_
timestamp 1728341909
transform -1 0 7530 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2386_
timestamp 1728341909
transform -1 0 6650 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2387_
timestamp 1728341909
transform -1 0 6410 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2388_
timestamp 1728341909
transform -1 0 8970 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2389_
timestamp 1728341909
transform -1 0 8350 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2390_
timestamp 1728341909
transform -1 0 8290 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2391_
timestamp 1728341909
transform -1 0 9530 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2392_
timestamp 1728341909
transform 1 0 8290 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2393_
timestamp 1728341909
transform 1 0 8250 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2394_
timestamp 1728341909
transform 1 0 8890 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2395_
timestamp 1728341909
transform 1 0 8850 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2396_
timestamp 1728341909
transform 1 0 9130 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2397_
timestamp 1728341909
transform -1 0 9390 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2398_
timestamp 1728341909
transform 1 0 8770 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2399_
timestamp 1728341909
transform -1 0 7650 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2400_
timestamp 1728341909
transform 1 0 7390 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2401_
timestamp 1728341909
transform 1 0 8510 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2402_
timestamp 1728341909
transform -1 0 6450 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2403_
timestamp 1728341909
transform -1 0 6650 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2404_
timestamp 1728341909
transform -1 0 7610 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2405_
timestamp 1728341909
transform -1 0 7390 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2406_
timestamp 1728341909
transform 1 0 7110 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2407_
timestamp 1728341909
transform -1 0 6650 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2408_
timestamp 1728341909
transform -1 0 5950 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2409_
timestamp 1728341909
transform 1 0 7030 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2410_
timestamp 1728341909
transform -1 0 7310 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2411_
timestamp 1728341909
transform -1 0 6870 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2412_
timestamp 1728341909
transform -1 0 7530 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2413_
timestamp 1728341909
transform 1 0 7050 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2414_
timestamp 1728341909
transform 1 0 6870 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2415_
timestamp 1728341909
transform -1 0 8070 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2416_
timestamp 1728341909
transform 1 0 7810 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2417_
timestamp 1728341909
transform -1 0 9050 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2418_
timestamp 1728341909
transform -1 0 8830 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2419_
timestamp 1728341909
transform 1 0 7090 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2420_
timestamp 1728341909
transform 1 0 2250 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2421_
timestamp 1728341909
transform -1 0 9710 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2422_
timestamp 1728341909
transform 1 0 8290 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__2423_
timestamp 1728341909
transform 1 0 9010 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2424_
timestamp 1728341909
transform 1 0 8790 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2425_
timestamp 1728341909
transform 1 0 3190 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2426_
timestamp 1728341909
transform 1 0 8770 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2427_
timestamp 1728341909
transform 1 0 8850 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__2428_
timestamp 1728341909
transform 1 0 9250 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2429_
timestamp 1728341909
transform 1 0 9470 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2430_
timestamp 1728341909
transform 1 0 8830 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2431_
timestamp 1728341909
transform -1 0 9290 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2432_
timestamp 1728341909
transform 1 0 9510 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2433_
timestamp 1728341909
transform -1 0 9930 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2434_
timestamp 1728341909
transform -1 0 10010 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2435_
timestamp 1728341909
transform 1 0 4470 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__2436_
timestamp 1728341909
transform 1 0 9230 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2437_
timestamp 1728341909
transform 1 0 10910 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__2438_
timestamp 1728341909
transform -1 0 10970 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__2439_
timestamp 1728341909
transform -1 0 10950 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__2440_
timestamp 1728341909
transform 1 0 9070 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__2441_
timestamp 1728341909
transform -1 0 6210 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__2442_
timestamp 1728341909
transform -1 0 8290 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2443_
timestamp 1728341909
transform 1 0 3850 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2444_
timestamp 1728341909
transform -1 0 4730 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__2445_
timestamp 1728341909
transform -1 0 8630 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__2446_
timestamp 1728341909
transform 1 0 8270 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2447_
timestamp 1728341909
transform 1 0 8110 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2448_
timestamp 1728341909
transform 1 0 8510 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2449_
timestamp 1728341909
transform -1 0 8790 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2450_
timestamp 1728341909
transform -1 0 8990 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2451_
timestamp 1728341909
transform 1 0 3850 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2452_
timestamp 1728341909
transform 1 0 7630 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2453_
timestamp 1728341909
transform -1 0 6650 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2454_
timestamp 1728341909
transform -1 0 6370 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2455_
timestamp 1728341909
transform -1 0 6650 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2456_
timestamp 1728341909
transform -1 0 8770 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2457_
timestamp 1728341909
transform -1 0 8990 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2458_
timestamp 1728341909
transform -1 0 6830 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2459_
timestamp 1728341909
transform -1 0 3610 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2460_
timestamp 1728341909
transform 1 0 7130 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2461_
timestamp 1728341909
transform 1 0 7050 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2462_
timestamp 1728341909
transform -1 0 7330 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2463_
timestamp 1728341909
transform -1 0 7350 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2464_
timestamp 1728341909
transform 1 0 4510 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__2465_
timestamp 1728341909
transform -1 0 7410 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2466_
timestamp 1728341909
transform -1 0 3390 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2467_
timestamp 1728341909
transform 1 0 6210 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2468_
timestamp 1728341909
transform -1 0 6330 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2469_
timestamp 1728341909
transform -1 0 6170 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2470_
timestamp 1728341909
transform -1 0 6430 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2471_
timestamp 1728341909
transform -1 0 8090 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2472_
timestamp 1728341909
transform -1 0 6110 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2473_
timestamp 1728341909
transform -1 0 5450 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2474_
timestamp 1728341909
transform -1 0 5370 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2475_
timestamp 1728341909
transform -1 0 7830 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__2476_
timestamp 1728341909
transform -1 0 2750 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2477_
timestamp 1728341909
transform -1 0 5230 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2478_
timestamp 1728341909
transform 1 0 5310 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2479_
timestamp 1728341909
transform -1 0 8050 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2480_
timestamp 1728341909
transform 1 0 5950 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2481_
timestamp 1728341909
transform 1 0 4210 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2482_
timestamp 1728341909
transform -1 0 2490 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2483_
timestamp 1728341909
transform -1 0 4730 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2484_
timestamp 1728341909
transform -1 0 5770 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2485_
timestamp 1728341909
transform -1 0 7010 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2486_
timestamp 1728341909
transform 1 0 3130 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2487_
timestamp 1728341909
transform -1 0 5710 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2488_
timestamp 1728341909
transform 1 0 6470 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2489_
timestamp 1728341909
transform -1 0 6750 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2490_
timestamp 1728341909
transform 1 0 7730 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2491_
timestamp 1728341909
transform -1 0 7970 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2492_
timestamp 1728341909
transform -1 0 2910 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2493_
timestamp 1728341909
transform -1 0 5550 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2494_
timestamp 1728341909
transform -1 0 6630 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2495_
timestamp 1728341909
transform 1 0 6870 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2496_
timestamp 1728341909
transform 1 0 7590 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2497_
timestamp 1728341909
transform -1 0 7830 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2498_
timestamp 1728341909
transform -1 0 8810 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__2499_
timestamp 1728341909
transform 1 0 9050 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2500_
timestamp 1728341909
transform -1 0 7670 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2501_
timestamp 1728341909
transform -1 0 6790 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__2502_
timestamp 1728341909
transform -1 0 7650 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__2503_
timestamp 1728341909
transform 1 0 11150 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2504_
timestamp 1728341909
transform -1 0 4590 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2505_
timestamp 1728341909
transform -1 0 5730 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2506_
timestamp 1728341909
transform -1 0 6750 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__2507_
timestamp 1728341909
transform 1 0 5890 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2508_
timestamp 1728341909
transform 1 0 5690 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2509_
timestamp 1728341909
transform -1 0 8850 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__2510_
timestamp 1728341909
transform -1 0 8110 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__2511_
timestamp 1728341909
transform -1 0 7430 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__2512_
timestamp 1728341909
transform 1 0 7130 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__2513_
timestamp 1728341909
transform 1 0 6910 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__2514_
timestamp 1728341909
transform 1 0 7070 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__2515_
timestamp 1728341909
transform 1 0 10410 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__2516_
timestamp 1728341909
transform 1 0 8550 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2517_
timestamp 1728341909
transform 1 0 10650 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2518_
timestamp 1728341909
transform -1 0 9750 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__2519_
timestamp 1728341909
transform 1 0 9990 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__2520_
timestamp 1728341909
transform -1 0 10450 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2521_
timestamp 1728341909
transform -1 0 8550 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2522_
timestamp 1728341909
transform 1 0 6110 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2523_
timestamp 1728341909
transform 1 0 5930 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2524_
timestamp 1728341909
transform 1 0 8310 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2525_
timestamp 1728341909
transform 1 0 6810 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2526_
timestamp 1728341909
transform -1 0 7810 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2527_
timestamp 1728341909
transform 1 0 8030 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2528_
timestamp 1728341909
transform -1 0 8090 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2529_
timestamp 1728341909
transform 1 0 7870 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2530_
timestamp 1728341909
transform -1 0 7830 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2531_
timestamp 1728341909
transform -1 0 7850 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2532_
timestamp 1728341909
transform 1 0 7850 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2533_
timestamp 1728341909
transform -1 0 5510 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2534_
timestamp 1728341909
transform -1 0 5930 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2535_
timestamp 1728341909
transform -1 0 7610 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2536_
timestamp 1728341909
transform 1 0 7410 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2537_
timestamp 1728341909
transform 1 0 7330 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2538_
timestamp 1728341909
transform 1 0 8050 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2539_
timestamp 1728341909
transform 1 0 5910 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2540_
timestamp 1728341909
transform 1 0 5630 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2541_
timestamp 1728341909
transform 1 0 6150 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2542_
timestamp 1728341909
transform -1 0 6690 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2543_
timestamp 1728341909
transform -1 0 6650 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2544_
timestamp 1728341909
transform 1 0 6190 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2545_
timestamp 1728341909
transform 1 0 6890 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2546_
timestamp 1728341909
transform 1 0 6150 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2547_
timestamp 1728341909
transform 1 0 6370 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2548_
timestamp 1728341909
transform 1 0 7150 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2549_
timestamp 1728341909
transform 1 0 7410 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2550_
timestamp 1728341909
transform -1 0 7570 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2551_
timestamp 1728341909
transform -1 0 6290 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2552_
timestamp 1728341909
transform -1 0 4850 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2553_
timestamp 1728341909
transform -1 0 5890 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2554_
timestamp 1728341909
transform -1 0 5610 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2555_
timestamp 1728341909
transform 1 0 5670 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2556_
timestamp 1728341909
transform 1 0 5050 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2557_
timestamp 1728341909
transform 1 0 5790 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2558_
timestamp 1728341909
transform -1 0 6430 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2559_
timestamp 1728341909
transform 1 0 6110 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__2560_
timestamp 1728341909
transform 1 0 4370 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2561_
timestamp 1728341909
transform -1 0 5430 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2562_
timestamp 1728341909
transform 1 0 5050 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2563_
timestamp 1728341909
transform -1 0 4950 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2564_
timestamp 1728341909
transform -1 0 4610 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2565_
timestamp 1728341909
transform 1 0 4750 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2566_
timestamp 1728341909
transform -1 0 4970 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2567_
timestamp 1728341909
transform 1 0 5170 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2568_
timestamp 1728341909
transform 1 0 5310 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__2569_
timestamp 1728341909
transform -1 0 4190 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2570_
timestamp 1728341909
transform 1 0 5210 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2571_
timestamp 1728341909
transform 1 0 4330 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2572_
timestamp 1728341909
transform -1 0 4450 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2573_
timestamp 1728341909
transform 1 0 4690 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2574_
timestamp 1728341909
transform 1 0 5410 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2575_
timestamp 1728341909
transform -1 0 4970 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2576_
timestamp 1728341909
transform 1 0 5150 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2577_
timestamp 1728341909
transform 1 0 4890 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2578_
timestamp 1728341909
transform -1 0 4830 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2579_
timestamp 1728341909
transform 1 0 4690 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__2580_
timestamp 1728341909
transform 1 0 4730 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__2581_
timestamp 1728341909
transform -1 0 4170 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2582_
timestamp 1728341909
transform -1 0 3310 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2583_
timestamp 1728341909
transform 1 0 2250 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2584_
timestamp 1728341909
transform 1 0 3210 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2585_
timestamp 1728341909
transform -1 0 6370 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2586_
timestamp 1728341909
transform -1 0 3730 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2587_
timestamp 1728341909
transform -1 0 3470 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2588_
timestamp 1728341909
transform -1 0 2990 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2589_
timestamp 1728341909
transform -1 0 2990 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2590_
timestamp 1728341909
transform 1 0 3610 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__2591_
timestamp 1728341909
transform -1 0 3090 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2592_
timestamp 1728341909
transform 1 0 2590 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2593_
timestamp 1728341909
transform -1 0 2690 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2594_
timestamp 1728341909
transform -1 0 2710 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2595_
timestamp 1728341909
transform -1 0 3790 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__2596_
timestamp 1728341909
transform 1 0 3390 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2597_
timestamp 1728341909
transform 1 0 3330 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2598_
timestamp 1728341909
transform -1 0 3210 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2599_
timestamp 1728341909
transform -1 0 3210 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2600_
timestamp 1728341909
transform 1 0 2930 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2601_
timestamp 1728341909
transform -1 0 2490 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2602_
timestamp 1728341909
transform -1 0 2750 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2603_
timestamp 1728341909
transform -1 0 2350 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2604_
timestamp 1728341909
transform 1 0 2490 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2605_
timestamp 1728341909
transform -1 0 2490 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2606_
timestamp 1728341909
transform 1 0 2210 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2607_
timestamp 1728341909
transform -1 0 1570 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2608_
timestamp 1728341909
transform -1 0 1090 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2609_
timestamp 1728341909
transform 1 0 2050 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2610_
timestamp 1728341909
transform 1 0 1290 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2611_
timestamp 1728341909
transform -1 0 1270 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2612_
timestamp 1728341909
transform -1 0 1010 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2613_
timestamp 1728341909
transform -1 0 1990 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2614_
timestamp 1728341909
transform -1 0 610 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2615_
timestamp 1728341909
transform 1 0 1790 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2616_
timestamp 1728341909
transform 1 0 1530 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2617_
timestamp 1728341909
transform -1 0 1530 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2618_
timestamp 1728341909
transform -1 0 1770 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2619_
timestamp 1728341909
transform 1 0 810 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2620_
timestamp 1728341909
transform -1 0 1330 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2621_
timestamp 1728341909
transform 1 0 1070 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2622_
timestamp 1728341909
transform -1 0 1290 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2623_
timestamp 1728341909
transform 1 0 1030 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2624_
timestamp 1728341909
transform -1 0 570 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2625_
timestamp 1728341909
transform -1 0 2650 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2626_
timestamp 1728341909
transform 1 0 1670 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2627_
timestamp 1728341909
transform 1 0 1410 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2628_
timestamp 1728341909
transform 1 0 810 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2629_
timestamp 1728341909
transform -1 0 3410 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__2630_
timestamp 1728341909
transform 1 0 4270 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__2631_
timestamp 1728341909
transform -1 0 4930 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__2632_
timestamp 1728341909
transform 1 0 10910 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2633_
timestamp 1728341909
transform 1 0 3910 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2634_
timestamp 1728341909
transform 1 0 9010 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2635_
timestamp 1728341909
transform -1 0 2290 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__2636_
timestamp 1728341909
transform -1 0 9170 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__2637_
timestamp 1728341909
transform 1 0 4370 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2638_
timestamp 1728341909
transform 1 0 4870 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2639_
timestamp 1728341909
transform -1 0 9950 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__2640_
timestamp 1728341909
transform -1 0 9890 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__2641_
timestamp 1728341909
transform 1 0 10190 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2642_
timestamp 1728341909
transform -1 0 9530 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__2643_
timestamp 1728341909
transform 1 0 10930 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2644_
timestamp 1728341909
transform -1 0 9770 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2645_
timestamp 1728341909
transform -1 0 9730 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__2646_
timestamp 1728341909
transform 1 0 10130 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__2647_
timestamp 1728341909
transform -1 0 8610 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2648_
timestamp 1728341909
transform -1 0 4190 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__2649_
timestamp 1728341909
transform -1 0 5830 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2650_
timestamp 1728341909
transform 1 0 9330 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__2651_
timestamp 1728341909
transform -1 0 5710 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2652_
timestamp 1728341909
transform -1 0 7870 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__2653_
timestamp 1728341909
transform -1 0 7770 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__2654_
timestamp 1728341909
transform 1 0 4690 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2655_
timestamp 1728341909
transform -1 0 5470 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2656_
timestamp 1728341909
transform -1 0 6050 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2657_
timestamp 1728341909
transform -1 0 6790 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2658_
timestamp 1728341909
transform 1 0 6290 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2659_
timestamp 1728341909
transform 1 0 6990 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2660_
timestamp 1728341909
transform -1 0 7270 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2661_
timestamp 1728341909
transform -1 0 4490 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2662_
timestamp 1728341909
transform 1 0 4450 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2663_
timestamp 1728341909
transform 1 0 6370 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2664_
timestamp 1728341909
transform -1 0 6630 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2665_
timestamp 1728341909
transform 1 0 7130 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2666_
timestamp 1728341909
transform 1 0 6870 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2667_
timestamp 1728341909
transform 1 0 7610 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2668_
timestamp 1728341909
transform 1 0 7350 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2669_
timestamp 1728341909
transform 1 0 8010 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2670_
timestamp 1728341909
transform -1 0 4230 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2671_
timestamp 1728341909
transform -1 0 5350 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__2672_
timestamp 1728341909
transform 1 0 5250 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2673_
timestamp 1728341909
transform 1 0 7210 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2674_
timestamp 1728341909
transform -1 0 7430 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2675_
timestamp 1728341909
transform 1 0 7670 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2676_
timestamp 1728341909
transform -1 0 7610 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2677_
timestamp 1728341909
transform 1 0 7790 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2678_
timestamp 1728341909
transform 1 0 7750 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2679_
timestamp 1728341909
transform 1 0 4190 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2680_
timestamp 1728341909
transform -1 0 4450 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2681_
timestamp 1728341909
transform 1 0 6150 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2682_
timestamp 1728341909
transform 1 0 6770 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2683_
timestamp 1728341909
transform 1 0 4110 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2684_
timestamp 1728341909
transform -1 0 5770 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2685_
timestamp 1728341909
transform 1 0 5490 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2686_
timestamp 1728341909
transform -1 0 6910 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2687_
timestamp 1728341909
transform 1 0 7370 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2688_
timestamp 1728341909
transform -1 0 7510 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2689_
timestamp 1728341909
transform 1 0 6530 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2690_
timestamp 1728341909
transform 1 0 6610 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2691_
timestamp 1728341909
transform 1 0 7110 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2692_
timestamp 1728341909
transform -1 0 7250 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2693_
timestamp 1728341909
transform 1 0 5090 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2694_
timestamp 1728341909
transform -1 0 5230 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2695_
timestamp 1728341909
transform 1 0 6670 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2696_
timestamp 1728341909
transform 1 0 6610 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2697_
timestamp 1728341909
transform 1 0 7030 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2698_
timestamp 1728341909
transform 1 0 6930 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2699_
timestamp 1728341909
transform -1 0 6370 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2700_
timestamp 1728341909
transform 1 0 5430 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2701_
timestamp 1728341909
transform -1 0 5510 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2702_
timestamp 1728341909
transform -1 0 5590 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2703_
timestamp 1728341909
transform -1 0 5610 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2704_
timestamp 1728341909
transform 1 0 5670 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2705_
timestamp 1728341909
transform 1 0 5930 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2706_
timestamp 1728341909
transform -1 0 6190 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2707_
timestamp 1728341909
transform -1 0 5930 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2708_
timestamp 1728341909
transform -1 0 2330 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2709_
timestamp 1728341909
transform -1 0 4990 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2710_
timestamp 1728341909
transform -1 0 4910 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2711_
timestamp 1728341909
transform -1 0 5110 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2712_
timestamp 1728341909
transform -1 0 5690 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2713_
timestamp 1728341909
transform -1 0 5830 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2714_
timestamp 1728341909
transform -1 0 6130 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2715_
timestamp 1728341909
transform 1 0 5850 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2716_
timestamp 1728341909
transform -1 0 6690 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2717_
timestamp 1728341909
transform 1 0 6630 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2718_
timestamp 1728341909
transform 1 0 6210 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2719_
timestamp 1728341909
transform -1 0 6370 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2720_
timestamp 1728341909
transform 1 0 4670 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2721_
timestamp 1728341909
transform 1 0 4950 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2722_
timestamp 1728341909
transform 1 0 5190 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2723_
timestamp 1728341909
transform -1 0 5450 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2724_
timestamp 1728341909
transform 1 0 6170 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2725_
timestamp 1728341909
transform 1 0 6410 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2726_
timestamp 1728341909
transform -1 0 6170 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__2727_
timestamp 1728341909
transform 1 0 5870 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__2728_
timestamp 1728341909
transform -1 0 4350 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2729_
timestamp 1728341909
transform -1 0 4210 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2730_
timestamp 1728341909
transform -1 0 5250 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2731_
timestamp 1728341909
transform -1 0 5370 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2732_
timestamp 1728341909
transform -1 0 5670 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2733_
timestamp 1728341909
transform -1 0 5930 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2734_
timestamp 1728341909
transform -1 0 5250 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2735_
timestamp 1728341909
transform 1 0 5450 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2736_
timestamp 1728341909
transform -1 0 8370 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__2737_
timestamp 1728341909
transform 1 0 3770 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2738_
timestamp 1728341909
transform 1 0 3950 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2739_
timestamp 1728341909
transform -1 0 3770 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2740_
timestamp 1728341909
transform -1 0 3710 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2741_
timestamp 1728341909
transform -1 0 4050 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2742_
timestamp 1728341909
transform -1 0 4190 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2743_
timestamp 1728341909
transform 1 0 4930 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2744_
timestamp 1728341909
transform 1 0 4670 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__2745_
timestamp 1728341909
transform 1 0 5150 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2746_
timestamp 1728341909
transform 1 0 4650 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2747_
timestamp 1728341909
transform 1 0 5570 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2748_
timestamp 1728341909
transform -1 0 4970 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2749_
timestamp 1728341909
transform -1 0 5330 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2750_
timestamp 1728341909
transform -1 0 5430 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2751_
timestamp 1728341909
transform 1 0 4410 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2752_
timestamp 1728341909
transform 1 0 3910 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2753_
timestamp 1728341909
transform -1 0 3450 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2754_
timestamp 1728341909
transform -1 0 3030 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2755_
timestamp 1728341909
transform 1 0 3290 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2756_
timestamp 1728341909
transform -1 0 3670 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2757_
timestamp 1728341909
transform -1 0 3690 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2758_
timestamp 1728341909
transform -1 0 3670 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2759_
timestamp 1728341909
transform -1 0 3550 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2760_
timestamp 1728341909
transform -1 0 3590 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2761_
timestamp 1728341909
transform -1 0 3730 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2762_
timestamp 1728341909
transform -1 0 3490 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2763_
timestamp 1728341909
transform 1 0 3050 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__2764_
timestamp 1728341909
transform 1 0 3330 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__2765_
timestamp 1728341909
transform -1 0 2650 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2766_
timestamp 1728341909
transform 1 0 3730 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__2767_
timestamp 1728341909
transform -1 0 4430 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2768_
timestamp 1728341909
transform 1 0 4510 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2769_
timestamp 1728341909
transform 1 0 5170 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2770_
timestamp 1728341909
transform -1 0 4670 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2771_
timestamp 1728341909
transform -1 0 4950 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2772_
timestamp 1728341909
transform -1 0 4930 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2773_
timestamp 1728341909
transform 1 0 2690 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2774_
timestamp 1728341909
transform -1 0 2550 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__2775_
timestamp 1728341909
transform 1 0 3910 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2776_
timestamp 1728341909
transform 1 0 4430 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2777_
timestamp 1728341909
transform 1 0 5170 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2778_
timestamp 1728341909
transform -1 0 4670 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2779_
timestamp 1728341909
transform 1 0 3990 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__2780_
timestamp 1728341909
transform 1 0 2770 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__2781_
timestamp 1728341909
transform -1 0 3990 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2782_
timestamp 1728341909
transform -1 0 2790 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2783_
timestamp 1728341909
transform 1 0 2490 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2784_
timestamp 1728341909
transform 1 0 570 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2785_
timestamp 1728341909
transform -1 0 2270 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2786_
timestamp 1728341909
transform 1 0 2530 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2787_
timestamp 1728341909
transform -1 0 2950 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2788_
timestamp 1728341909
transform -1 0 2450 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2789_
timestamp 1728341909
transform -1 0 3750 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2790_
timestamp 1728341909
transform 1 0 3230 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2791_
timestamp 1728341909
transform -1 0 2970 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2792_
timestamp 1728341909
transform -1 0 2870 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2793_
timestamp 1728341909
transform -1 0 2290 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__2794_
timestamp 1728341909
transform 1 0 2170 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2795_
timestamp 1728341909
transform 1 0 810 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2796_
timestamp 1728341909
transform 1 0 1750 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2797_
timestamp 1728341909
transform -1 0 2030 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2798_
timestamp 1728341909
transform 1 0 1250 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2799_
timestamp 1728341909
transform -1 0 1530 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2800_
timestamp 1728341909
transform -1 0 1790 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2801_
timestamp 1728341909
transform 1 0 1750 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2802_
timestamp 1728341909
transform 1 0 1830 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2803_
timestamp 1728341909
transform 1 0 3310 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2804_
timestamp 1728341909
transform -1 0 470 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__2805_
timestamp 1728341909
transform 1 0 7010 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2806_
timestamp 1728341909
transform -1 0 5430 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2807_
timestamp 1728341909
transform -1 0 5030 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2808_
timestamp 1728341909
transform 1 0 3950 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2809_
timestamp 1728341909
transform -1 0 4410 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2810_
timestamp 1728341909
transform -1 0 4770 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2811_
timestamp 1728341909
transform -1 0 4630 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2812_
timestamp 1728341909
transform 1 0 4250 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2813_
timestamp 1728341909
transform 1 0 4010 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__2814_
timestamp 1728341909
transform 1 0 4130 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__2815_
timestamp 1728341909
transform -1 0 4210 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2816_
timestamp 1728341909
transform 1 0 2510 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2817_
timestamp 1728341909
transform -1 0 2790 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__2818_
timestamp 1728341909
transform 1 0 2750 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2819_
timestamp 1728341909
transform 1 0 3190 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2820_
timestamp 1728341909
transform 1 0 3430 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2821_
timestamp 1728341909
transform -1 0 3970 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2822_
timestamp 1728341909
transform -1 0 4770 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2823_
timestamp 1728341909
transform -1 0 1750 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2824_
timestamp 1728341909
transform 1 0 570 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__2825_
timestamp 1728341909
transform 1 0 550 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2826_
timestamp 1728341909
transform -1 0 710 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__2827_
timestamp 1728341909
transform 1 0 1750 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2828_
timestamp 1728341909
transform -1 0 2030 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2829_
timestamp 1728341909
transform 1 0 1270 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2830_
timestamp 1728341909
transform -1 0 1530 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2831_
timestamp 1728341909
transform -1 0 1550 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__2832_
timestamp 1728341909
transform 1 0 2050 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2833_
timestamp 1728341909
transform -1 0 1070 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__2834_
timestamp 1728341909
transform 1 0 890 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__2835_
timestamp 1728341909
transform 1 0 1130 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__2836_
timestamp 1728341909
transform 1 0 1350 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__2837_
timestamp 1728341909
transform 1 0 1670 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__2838_
timestamp 1728341909
transform -1 0 1550 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__2839_
timestamp 1728341909
transform 1 0 830 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__2840_
timestamp 1728341909
transform 1 0 1270 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2841_
timestamp 1728341909
transform 1 0 2070 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2842_
timestamp 1728341909
transform -1 0 1730 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2843_
timestamp 1728341909
transform -1 0 1830 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2844_
timestamp 1728341909
transform -1 0 1590 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__2845_
timestamp 1728341909
transform -1 0 1530 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2846_
timestamp 1728341909
transform 1 0 1310 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2847_
timestamp 1728341909
transform -1 0 1310 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__2848_
timestamp 1728341909
transform -1 0 1290 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2849_
timestamp 1728341909
transform -1 0 1590 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2850_
timestamp 1728341909
transform -1 0 1510 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2851_
timestamp 1728341909
transform -1 0 1050 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2852_
timestamp 1728341909
transform -1 0 1110 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2853_
timestamp 1728341909
transform -1 0 2310 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2854_
timestamp 1728341909
transform 1 0 790 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__2855_
timestamp 1728341909
transform 1 0 2470 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__2856_
timestamp 1728341909
transform -1 0 1990 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__2857_
timestamp 1728341909
transform -1 0 2390 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__2858_
timestamp 1728341909
transform -1 0 2290 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__2859_
timestamp 1728341909
transform -1 0 870 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2860_
timestamp 1728341909
transform 1 0 550 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2861_
timestamp 1728341909
transform -1 0 110 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2862_
timestamp 1728341909
transform -1 0 1070 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__2863_
timestamp 1728341909
transform 1 0 310 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__2864_
timestamp 1728341909
transform -1 0 350 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__2865_
timestamp 1728341909
transform 1 0 4470 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__2866_
timestamp 1728341909
transform 1 0 4490 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2867_
timestamp 1728341909
transform 1 0 5590 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__2868_
timestamp 1728341909
transform -1 0 2970 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2869_
timestamp 1728341909
transform -1 0 3250 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__2870_
timestamp 1728341909
transform -1 0 2310 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__2871_
timestamp 1728341909
transform 1 0 2330 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__2872_
timestamp 1728341909
transform -1 0 4610 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__2873_
timestamp 1728341909
transform 1 0 4350 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__2874_
timestamp 1728341909
transform -1 0 4150 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2875_
timestamp 1728341909
transform -1 0 1710 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2876_
timestamp 1728341909
transform -1 0 850 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2877_
timestamp 1728341909
transform -1 0 3510 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2878_
timestamp 1728341909
transform -1 0 3950 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2879_
timestamp 1728341909
transform -1 0 1290 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2880_
timestamp 1728341909
transform 1 0 1470 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2881_
timestamp 1728341909
transform -1 0 1790 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2882_
timestamp 1728341909
transform -1 0 2470 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2883_
timestamp 1728341909
transform 1 0 4470 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2884_
timestamp 1728341909
transform 1 0 4190 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2885_
timestamp 1728341909
transform 1 0 3130 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2886_
timestamp 1728341909
transform 1 0 4690 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2887_
timestamp 1728341909
transform 1 0 5150 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2888_
timestamp 1728341909
transform 1 0 3410 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2889_
timestamp 1728341909
transform 1 0 3630 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2890_
timestamp 1728341909
transform -1 0 4410 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2891_
timestamp 1728341909
transform -1 0 4150 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2892_
timestamp 1728341909
transform -1 0 2010 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2893_
timestamp 1728341909
transform 1 0 3690 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2894_
timestamp 1728341909
transform 1 0 3890 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2895_
timestamp 1728341909
transform 1 0 4470 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2896_
timestamp 1728341909
transform -1 0 3870 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2897_
timestamp 1728341909
transform -1 0 5870 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2898_
timestamp 1728341909
transform 1 0 5190 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2899_
timestamp 1728341909
transform 1 0 5150 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2900_
timestamp 1728341909
transform 1 0 5410 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2901_
timestamp 1728341909
transform -1 0 4890 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2902_
timestamp 1728341909
transform -1 0 1550 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2903_
timestamp 1728341909
transform 1 0 2210 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2904_
timestamp 1728341909
transform 1 0 2470 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2905_
timestamp 1728341909
transform 1 0 1270 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2906_
timestamp 1728341909
transform 1 0 1050 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2907_
timestamp 1728341909
transform 1 0 1250 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2908_
timestamp 1728341909
transform -1 0 1570 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2909_
timestamp 1728341909
transform -1 0 1790 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2910_
timestamp 1728341909
transform -1 0 1570 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2911_
timestamp 1728341909
transform -1 0 1570 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2912_
timestamp 1728341909
transform -1 0 2490 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2913_
timestamp 1728341909
transform -1 0 1730 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2914_
timestamp 1728341909
transform 1 0 2250 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2915_
timestamp 1728341909
transform 1 0 2030 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2916_
timestamp 1728341909
transform 1 0 1710 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2917_
timestamp 1728341909
transform -1 0 1790 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2918_
timestamp 1728341909
transform 1 0 1730 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2919_
timestamp 1728341909
transform -1 0 2270 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2920_
timestamp 1728341909
transform -1 0 1990 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2921_
timestamp 1728341909
transform -1 0 2050 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2922_
timestamp 1728341909
transform -1 0 1970 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2923_
timestamp 1728341909
transform -1 0 2010 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2924_
timestamp 1728341909
transform -1 0 2970 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2925_
timestamp 1728341909
transform 1 0 3450 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2926_
timestamp 1728341909
transform -1 0 2430 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2927_
timestamp 1728341909
transform -1 0 2470 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2928_
timestamp 1728341909
transform 1 0 4610 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2929_
timestamp 1728341909
transform 1 0 3450 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2930_
timestamp 1728341909
transform -1 0 2730 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2931_
timestamp 1728341909
transform -1 0 2970 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2932_
timestamp 1728341909
transform 1 0 3170 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2933_
timestamp 1728341909
transform -1 0 2730 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2934_
timestamp 1728341909
transform 1 0 2950 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2935_
timestamp 1728341909
transform -1 0 1330 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2936_
timestamp 1728341909
transform -1 0 870 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2937_
timestamp 1728341909
transform 1 0 590 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2938_
timestamp 1728341909
transform 1 0 1750 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2939_
timestamp 1728341909
transform -1 0 1530 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2940_
timestamp 1728341909
transform 1 0 3190 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2941_
timestamp 1728341909
transform 1 0 3190 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2942_
timestamp 1728341909
transform -1 0 3410 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2943_
timestamp 1728341909
transform -1 0 3250 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2944_
timestamp 1728341909
transform -1 0 3750 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2945_
timestamp 1728341909
transform 1 0 3190 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__2946_
timestamp 1728341909
transform 1 0 3630 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__2947_
timestamp 1728341909
transform 1 0 3210 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2948_
timestamp 1728341909
transform -1 0 4210 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2949_
timestamp 1728341909
transform 1 0 3170 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__2950_
timestamp 1728341909
transform 1 0 2490 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2951_
timestamp 1728341909
transform -1 0 2730 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2952_
timestamp 1728341909
transform -1 0 3010 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2953_
timestamp 1728341909
transform -1 0 2210 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2954_
timestamp 1728341909
transform -1 0 2450 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2955_
timestamp 1728341909
transform 1 0 3030 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__2956_
timestamp 1728341909
transform 1 0 3270 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__2957_
timestamp 1728341909
transform 1 0 3770 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__2958_
timestamp 1728341909
transform 1 0 2210 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__2959_
timestamp 1728341909
transform 1 0 3490 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__2960_
timestamp 1728341909
transform 1 0 3610 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__2961_
timestamp 1728341909
transform 1 0 2730 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2962_
timestamp 1728341909
transform 1 0 2470 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2963_
timestamp 1728341909
transform 1 0 2990 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2964_
timestamp 1728341909
transform 1 0 2730 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2965_
timestamp 1728341909
transform -1 0 5810 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2966_
timestamp 1728341909
transform 1 0 4130 0 1 1690
box -12 -8 32 252
use FILL  FILL_4__2967_
timestamp 1728341909
transform -1 0 4610 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2968_
timestamp 1728341909
transform -1 0 4850 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2969_
timestamp 1728341909
transform -1 0 1350 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__2970_
timestamp 1728341909
transform -1 0 1530 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__2971_
timestamp 1728341909
transform -1 0 1550 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2972_
timestamp 1728341909
transform -1 0 1290 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2973_
timestamp 1728341909
transform -1 0 1050 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__2974_
timestamp 1728341909
transform -1 0 1790 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2975_
timestamp 1728341909
transform -1 0 2010 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2976_
timestamp 1728341909
transform 1 0 3890 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2977_
timestamp 1728341909
transform -1 0 4450 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2978_
timestamp 1728341909
transform 1 0 4170 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2979_
timestamp 1728341909
transform 1 0 1550 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2980_
timestamp 1728341909
transform -1 0 1030 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2981_
timestamp 1728341909
transform -1 0 790 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2982_
timestamp 1728341909
transform 1 0 2230 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2983_
timestamp 1728341909
transform -1 0 550 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2984_
timestamp 1728341909
transform -1 0 330 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2985_
timestamp 1728341909
transform -1 0 110 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__2986_
timestamp 1728341909
transform -1 0 370 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2987_
timestamp 1728341909
transform -1 0 630 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2988_
timestamp 1728341909
transform -1 0 590 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2989_
timestamp 1728341909
transform 1 0 350 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2990_
timestamp 1728341909
transform 1 0 90 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2991_
timestamp 1728341909
transform -1 0 370 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2992_
timestamp 1728341909
transform -1 0 2030 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__2993_
timestamp 1728341909
transform -1 0 1070 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2994_
timestamp 1728341909
transform -1 0 830 0 1 730
box -12 -8 32 252
use FILL  FILL_4__2995_
timestamp 1728341909
transform 1 0 610 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__2996_
timestamp 1728341909
transform -1 0 550 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__2997_
timestamp 1728341909
transform -1 0 870 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__2998_
timestamp 1728341909
transform -1 0 110 0 1 250
box -12 -8 32 252
use FILL  FILL_4__2999_
timestamp 1728341909
transform -1 0 350 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__3000_
timestamp 1728341909
transform -1 0 110 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__3001_
timestamp 1728341909
transform -1 0 110 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__3002_
timestamp 1728341909
transform -1 0 590 0 1 730
box -12 -8 32 252
use FILL  FILL_4__3003_
timestamp 1728341909
transform -1 0 110 0 1 730
box -12 -8 32 252
use FILL  FILL_4__3004_
timestamp 1728341909
transform -1 0 850 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__3005_
timestamp 1728341909
transform 1 0 810 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__3006_
timestamp 1728341909
transform -1 0 110 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__3007_
timestamp 1728341909
transform 1 0 1810 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3008_
timestamp 1728341909
transform -1 0 1070 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__3009_
timestamp 1728341909
transform -1 0 1330 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__3010_
timestamp 1728341909
transform -1 0 1330 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__3011_
timestamp 1728341909
transform -1 0 1090 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4__3012_
timestamp 1728341909
transform -1 0 1470 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__3013_
timestamp 1728341909
transform -1 0 1250 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__3014_
timestamp 1728341909
transform 1 0 1050 0 1 250
box -12 -8 32 252
use FILL  FILL_4__3015_
timestamp 1728341909
transform -1 0 1550 0 1 250
box -12 -8 32 252
use FILL  FILL_4__3016_
timestamp 1728341909
transform -1 0 1310 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__3017_
timestamp 1728341909
transform -1 0 1290 0 1 250
box -12 -8 32 252
use FILL  FILL_4__3018_
timestamp 1728341909
transform 1 0 1070 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4__3019_
timestamp 1728341909
transform -1 0 1070 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__3020_
timestamp 1728341909
transform -1 0 3710 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3021_
timestamp 1728341909
transform -1 0 5970 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__3022_
timestamp 1728341909
transform 1 0 2810 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3023_
timestamp 1728341909
transform 1 0 2830 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3024_
timestamp 1728341909
transform 1 0 3810 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3025_
timestamp 1728341909
transform -1 0 4230 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__3026_
timestamp 1728341909
transform -1 0 3090 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3027_
timestamp 1728341909
transform -1 0 3490 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__3028_
timestamp 1728341909
transform -1 0 4010 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3029_
timestamp 1728341909
transform -1 0 4510 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3030_
timestamp 1728341909
transform 1 0 3490 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__3031_
timestamp 1728341909
transform -1 0 3770 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__3032_
timestamp 1728341909
transform -1 0 2570 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3033_
timestamp 1728341909
transform -1 0 2590 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3034_
timestamp 1728341909
transform 1 0 2730 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__3035_
timestamp 1728341909
transform -1 0 2990 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__3036_
timestamp 1728341909
transform 1 0 3310 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3037_
timestamp 1728341909
transform -1 0 3750 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__3038_
timestamp 1728341909
transform -1 0 3310 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3039_
timestamp 1728341909
transform 1 0 3050 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3040_
timestamp 1728341909
transform 1 0 2190 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__3041_
timestamp 1728341909
transform 1 0 2730 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__3042_
timestamp 1728341909
transform 1 0 7490 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__3043_
timestamp 1728341909
transform 1 0 6330 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__3044_
timestamp 1728341909
transform 1 0 5350 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__3045_
timestamp 1728341909
transform 1 0 5770 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3046_
timestamp 1728341909
transform 1 0 5490 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__3047_
timestamp 1728341909
transform 1 0 4830 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__3048_
timestamp 1728341909
transform 1 0 5170 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__3049_
timestamp 1728341909
transform 1 0 5870 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3050_
timestamp 1728341909
transform -1 0 6890 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3051_
timestamp 1728341909
transform -1 0 6350 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__3052_
timestamp 1728341909
transform 1 0 6390 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3053_
timestamp 1728341909
transform 1 0 6130 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3054_
timestamp 1728341909
transform 1 0 5870 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3055_
timestamp 1728341909
transform -1 0 5970 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3056_
timestamp 1728341909
transform 1 0 4630 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__3057_
timestamp 1728341909
transform 1 0 4390 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__3058_
timestamp 1728341909
transform -1 0 4510 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3059_
timestamp 1728341909
transform 1 0 4330 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__3060_
timestamp 1728341909
transform -1 0 4310 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__3061_
timestamp 1728341909
transform 1 0 4010 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3062_
timestamp 1728341909
transform -1 0 4830 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__3063_
timestamp 1728341909
transform 1 0 4570 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__3064_
timestamp 1728341909
transform 1 0 6030 0 1 2170
box -12 -8 32 252
use FILL  FILL_4__3065_
timestamp 1728341909
transform 1 0 5810 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__3066_
timestamp 1728341909
transform -1 0 5810 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3067_
timestamp 1728341909
transform -1 0 5950 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__3068_
timestamp 1728341909
transform -1 0 6990 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3069_
timestamp 1728341909
transform -1 0 6490 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3070_
timestamp 1728341909
transform 1 0 6130 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3071_
timestamp 1728341909
transform -1 0 6410 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3072_
timestamp 1728341909
transform 1 0 6610 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__3073_
timestamp 1728341909
transform 1 0 6370 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__3074_
timestamp 1728341909
transform 1 0 430 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__3075_
timestamp 1728341909
transform -1 0 590 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__3076_
timestamp 1728341909
transform -1 0 4290 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3077_
timestamp 1728341909
transform 1 0 2030 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3078_
timestamp 1728341909
transform -1 0 5530 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3079_
timestamp 1728341909
transform 1 0 5070 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3080_
timestamp 1728341909
transform 1 0 4270 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3081_
timestamp 1728341909
transform 1 0 5910 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__3082_
timestamp 1728341909
transform -1 0 6910 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__3083_
timestamp 1728341909
transform 1 0 6070 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__3084_
timestamp 1728341909
transform -1 0 5750 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3085_
timestamp 1728341909
transform -1 0 5030 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3086_
timestamp 1728341909
transform 1 0 5510 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3087_
timestamp 1728341909
transform -1 0 5110 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__3088_
timestamp 1728341909
transform -1 0 5650 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__3089_
timestamp 1728341909
transform -1 0 5610 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__3090_
timestamp 1728341909
transform 1 0 4790 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3091_
timestamp 1728341909
transform -1 0 4750 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3092_
timestamp 1728341909
transform 1 0 5610 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4__3093_
timestamp 1728341909
transform -1 0 4010 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__3094_
timestamp 1728341909
transform 1 0 4450 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__3095_
timestamp 1728341909
transform 1 0 4750 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__3096_
timestamp 1728341909
transform 1 0 4730 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__3097_
timestamp 1728341909
transform 1 0 4970 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__3098_
timestamp 1728341909
transform -1 0 5070 0 1 2650
box -12 -8 32 252
use FILL  FILL_4__3099_
timestamp 1728341909
transform 1 0 5210 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__3100_
timestamp 1728341909
transform -1 0 5610 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__3101_
timestamp 1728341909
transform 1 0 5150 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__3102_
timestamp 1728341909
transform 1 0 4670 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__3103_
timestamp 1728341909
transform 1 0 4890 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__3104_
timestamp 1728341909
transform -1 0 5030 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3105_
timestamp 1728341909
transform 1 0 5350 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__3106_
timestamp 1728341909
transform 1 0 8530 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__3107_
timestamp 1728341909
transform 1 0 8290 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__3108_
timestamp 1728341909
transform 1 0 8050 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__3109_
timestamp 1728341909
transform -1 0 8590 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3110_
timestamp 1728341909
transform -1 0 8350 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3111_
timestamp 1728341909
transform 1 0 4530 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3112_
timestamp 1728341909
transform 1 0 4770 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3113_
timestamp 1728341909
transform -1 0 1290 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3114_
timestamp 1728341909
transform 1 0 790 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3115_
timestamp 1728341909
transform 1 0 4470 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__3116_
timestamp 1728341909
transform -1 0 4090 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3117_
timestamp 1728341909
transform -1 0 350 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__3118_
timestamp 1728341909
transform -1 0 110 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__3119_
timestamp 1728341909
transform -1 0 4950 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__3120_
timestamp 1728341909
transform 1 0 4450 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3121_
timestamp 1728341909
transform 1 0 5190 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__3122_
timestamp 1728341909
transform -1 0 4490 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3123_
timestamp 1728341909
transform -1 0 3750 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3124_
timestamp 1728341909
transform -1 0 3970 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3125_
timestamp 1728341909
transform -1 0 3710 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3126_
timestamp 1728341909
transform 1 0 4730 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3127_
timestamp 1728341909
transform 1 0 4750 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3128_
timestamp 1728341909
transform 1 0 4670 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__3129_
timestamp 1728341909
transform 1 0 3750 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__3130_
timestamp 1728341909
transform -1 0 1850 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3131_
timestamp 1728341909
transform -1 0 1350 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3132_
timestamp 1728341909
transform 1 0 1070 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3133_
timestamp 1728341909
transform 1 0 3930 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3134_
timestamp 1728341909
transform 1 0 3510 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3135_
timestamp 1728341909
transform 1 0 3250 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3136_
timestamp 1728341909
transform 1 0 3730 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3137_
timestamp 1728341909
transform 1 0 3990 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3138_
timestamp 1728341909
transform -1 0 4030 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3139_
timestamp 1728341909
transform 1 0 1090 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3140_
timestamp 1728341909
transform 1 0 830 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3141_
timestamp 1728341909
transform -1 0 4010 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3142_
timestamp 1728341909
transform 1 0 3770 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3143_
timestamp 1728341909
transform -1 0 4210 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3144_
timestamp 1728341909
transform -1 0 3490 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3145_
timestamp 1728341909
transform 1 0 3230 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3146_
timestamp 1728341909
transform -1 0 3310 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3147_
timestamp 1728341909
transform 1 0 3550 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3148_
timestamp 1728341909
transform -1 0 3510 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3149_
timestamp 1728341909
transform -1 0 3490 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__3150_
timestamp 1728341909
transform 1 0 2070 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3151_
timestamp 1728341909
transform -1 0 2310 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3152_
timestamp 1728341909
transform 1 0 7550 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3153_
timestamp 1728341909
transform 1 0 4470 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3154_
timestamp 1728341909
transform -1 0 810 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3155_
timestamp 1728341909
transform 1 0 1030 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3156_
timestamp 1728341909
transform 1 0 2990 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3157_
timestamp 1728341909
transform -1 0 2770 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3158_
timestamp 1728341909
transform 1 0 1990 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3159_
timestamp 1728341909
transform 1 0 2530 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3160_
timestamp 1728341909
transform 1 0 3150 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3161_
timestamp 1728341909
transform -1 0 2690 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3162_
timestamp 1728341909
transform -1 0 2470 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3163_
timestamp 1728341909
transform -1 0 1570 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3164_
timestamp 1728341909
transform 1 0 1270 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3165_
timestamp 1728341909
transform -1 0 350 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3166_
timestamp 1728341909
transform -1 0 110 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3167_
timestamp 1728341909
transform 1 0 2070 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3168_
timestamp 1728341909
transform 1 0 2010 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3169_
timestamp 1728341909
transform -1 0 2310 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3170_
timestamp 1728341909
transform 1 0 2050 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3171_
timestamp 1728341909
transform -1 0 2250 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3172_
timestamp 1728341909
transform 1 0 1910 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__3173_
timestamp 1728341909
transform -1 0 1790 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3174_
timestamp 1728341909
transform -1 0 1810 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3175_
timestamp 1728341909
transform -1 0 3050 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3176_
timestamp 1728341909
transform -1 0 2850 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3177_
timestamp 1728341909
transform 1 0 2290 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3178_
timestamp 1728341909
transform 1 0 2630 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3179_
timestamp 1728341909
transform 1 0 2290 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3180_
timestamp 1728341909
transform 1 0 3230 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3181_
timestamp 1728341909
transform -1 0 2950 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3182_
timestamp 1728341909
transform -1 0 3030 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3183_
timestamp 1728341909
transform 1 0 2790 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3184_
timestamp 1728341909
transform -1 0 2550 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3185_
timestamp 1728341909
transform -1 0 2550 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3186_
timestamp 1728341909
transform 1 0 2030 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3187_
timestamp 1728341909
transform -1 0 370 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3188_
timestamp 1728341909
transform -1 0 110 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3189_
timestamp 1728341909
transform 1 0 1050 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3190_
timestamp 1728341909
transform -1 0 850 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3191_
timestamp 1728341909
transform -1 0 1110 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3192_
timestamp 1728341909
transform 1 0 1730 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3193_
timestamp 1728341909
transform 1 0 1470 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3194_
timestamp 1728341909
transform 1 0 3270 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3195_
timestamp 1728341909
transform 1 0 3230 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__3196_
timestamp 1728341909
transform 1 0 1970 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3197_
timestamp 1728341909
transform -1 0 2550 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__3198_
timestamp 1728341909
transform -1 0 2130 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3199_
timestamp 1728341909
transform -1 0 2390 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3200_
timestamp 1728341909
transform 1 0 830 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3201_
timestamp 1728341909
transform -1 0 1070 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3202_
timestamp 1728341909
transform 1 0 1070 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3203_
timestamp 1728341909
transform -1 0 1330 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3204_
timestamp 1728341909
transform -1 0 590 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3205_
timestamp 1728341909
transform -1 0 590 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3206_
timestamp 1728341909
transform 1 0 1090 0 -1 4090
box -12 -8 32 252
use FILL  FILL_4__3207_
timestamp 1728341909
transform -1 0 350 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3208_
timestamp 1728341909
transform -1 0 110 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3209_
timestamp 1728341909
transform 1 0 330 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3210_
timestamp 1728341909
transform -1 0 110 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3211_
timestamp 1728341909
transform -1 0 1590 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3212_
timestamp 1728341909
transform -1 0 1330 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3213_
timestamp 1728341909
transform 1 0 1610 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3214_
timestamp 1728341909
transform 1 0 1350 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3215_
timestamp 1728341909
transform -1 0 1310 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3216_
timestamp 1728341909
transform 1 0 1050 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3217_
timestamp 1728341909
transform -1 0 350 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3218_
timestamp 1728341909
transform -1 0 110 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3219_
timestamp 1728341909
transform -1 0 1630 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3220_
timestamp 1728341909
transform 1 0 1850 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3221_
timestamp 1728341909
transform -1 0 370 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3222_
timestamp 1728341909
transform -1 0 110 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3223_
timestamp 1728341909
transform -1 0 850 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__3224_
timestamp 1728341909
transform 1 0 570 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3225_
timestamp 1728341909
transform -1 0 350 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3226_
timestamp 1728341909
transform -1 0 110 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3227_
timestamp 1728341909
transform -1 0 370 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__3228_
timestamp 1728341909
transform -1 0 110 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__3229_
timestamp 1728341909
transform -1 0 2030 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__3230_
timestamp 1728341909
transform 1 0 1750 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__3231_
timestamp 1728341909
transform 1 0 1550 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__3232_
timestamp 1728341909
transform -1 0 1810 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__3233_
timestamp 1728341909
transform 1 0 1110 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3234_
timestamp 1728341909
transform -1 0 1390 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3235_
timestamp 1728341909
transform 1 0 1070 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3236_
timestamp 1728341909
transform 1 0 1330 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3237_
timestamp 1728341909
transform 1 0 2250 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__3238_
timestamp 1728341909
transform 1 0 2490 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4__3239_
timestamp 1728341909
transform -1 0 590 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3240_
timestamp 1728341909
transform -1 0 830 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3241_
timestamp 1728341909
transform 1 0 9730 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__3242_
timestamp 1728341909
transform -1 0 9070 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4__3243_
timestamp 1728341909
transform 1 0 9490 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__3244_
timestamp 1728341909
transform 1 0 8790 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__3245_
timestamp 1728341909
transform 1 0 9090 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3246_
timestamp 1728341909
transform -1 0 9610 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3247_
timestamp 1728341909
transform 1 0 10510 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3248_
timestamp 1728341909
transform 1 0 10770 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3249_
timestamp 1728341909
transform -1 0 9510 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__3250_
timestamp 1728341909
transform 1 0 9430 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3251_
timestamp 1728341909
transform 1 0 9270 0 1 3130
box -12 -8 32 252
use FILL  FILL_4__3252_
timestamp 1728341909
transform -1 0 9290 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__3253_
timestamp 1728341909
transform -1 0 7910 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3254_
timestamp 1728341909
transform -1 0 8170 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3255_
timestamp 1728341909
transform -1 0 9350 0 1 3610
box -12 -8 32 252
use FILL  FILL_4__3256_
timestamp 1728341909
transform 1 0 8290 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3257_
timestamp 1728341909
transform 1 0 8050 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3258_
timestamp 1728341909
transform 1 0 8590 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3259_
timestamp 1728341909
transform 1 0 9530 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3260_
timestamp 1728341909
transform -1 0 10890 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__3261_
timestamp 1728341909
transform -1 0 10430 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3262_
timestamp 1728341909
transform 1 0 10010 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3263_
timestamp 1728341909
transform 1 0 9690 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__3264_
timestamp 1728341909
transform 1 0 9030 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4__3265_
timestamp 1728341909
transform -1 0 9770 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3266_
timestamp 1728341909
transform 1 0 9790 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3267_
timestamp 1728341909
transform -1 0 9690 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3268_
timestamp 1728341909
transform -1 0 10030 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3269_
timestamp 1728341909
transform -1 0 10530 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3270_
timestamp 1728341909
transform 1 0 10250 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3271_
timestamp 1728341909
transform -1 0 10070 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4__3272_
timestamp 1728341909
transform 1 0 10290 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4__3273_
timestamp 1728341909
transform -1 0 10190 0 1 4570
box -12 -8 32 252
use FILL  FILL_4__3274_
timestamp 1728341909
transform -1 0 10290 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3275_
timestamp 1728341909
transform 1 0 9610 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__3276_
timestamp 1728341909
transform -1 0 9230 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3277_
timestamp 1728341909
transform -1 0 10690 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3278_
timestamp 1728341909
transform 1 0 10150 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3279_
timestamp 1728341909
transform -1 0 9930 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3280_
timestamp 1728341909
transform 1 0 9270 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__3281_
timestamp 1728341909
transform 1 0 9030 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__3282_
timestamp 1728341909
transform -1 0 6910 0 1 4090
box -12 -8 32 252
use FILL  FILL_4__3283_
timestamp 1728341909
transform -1 0 6850 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3284_
timestamp 1728341909
transform 1 0 6610 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4__3285_
timestamp 1728341909
transform 1 0 7050 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3286_
timestamp 1728341909
transform -1 0 7310 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3287_
timestamp 1728341909
transform -1 0 6670 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3288_
timestamp 1728341909
transform -1 0 6890 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3289_
timestamp 1728341909
transform -1 0 6850 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__3290_
timestamp 1728341909
transform 1 0 6570 0 1 5530
box -12 -8 32 252
use FILL  FILL_4__3291_
timestamp 1728341909
transform 1 0 7070 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3292_
timestamp 1728341909
transform -1 0 7330 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3293_
timestamp 1728341909
transform 1 0 7170 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3294_
timestamp 1728341909
transform 1 0 6910 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3295_
timestamp 1728341909
transform 1 0 6110 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3296_
timestamp 1728341909
transform 1 0 5850 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3297_
timestamp 1728341909
transform 1 0 5470 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3298_
timestamp 1728341909
transform 1 0 5210 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3299_
timestamp 1728341909
transform 1 0 5650 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3300_
timestamp 1728341909
transform 1 0 5410 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3301_
timestamp 1728341909
transform 1 0 6910 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4__3302_
timestamp 1728341909
transform 1 0 2990 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3303_
timestamp 1728341909
transform -1 0 3050 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3304_
timestamp 1728341909
transform 1 0 1990 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3305_
timestamp 1728341909
transform -1 0 2250 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3306_
timestamp 1728341909
transform 1 0 3910 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3307_
timestamp 1728341909
transform -1 0 4850 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3308_
timestamp 1728341909
transform -1 0 110 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__3309_
timestamp 1728341909
transform -1 0 110 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3310_
timestamp 1728341909
transform -1 0 790 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__3311_
timestamp 1728341909
transform -1 0 830 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3312_
timestamp 1728341909
transform -1 0 330 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__3313_
timestamp 1728341909
transform -1 0 370 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3314_
timestamp 1728341909
transform -1 0 110 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3315_
timestamp 1728341909
transform -1 0 110 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3316_
timestamp 1728341909
transform -1 0 610 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3317_
timestamp 1728341909
transform -1 0 830 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3449_
timestamp 1728341909
transform -1 0 3850 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3450_
timestamp 1728341909
transform 1 0 3010 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3451_
timestamp 1728341909
transform 1 0 3130 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3452_
timestamp 1728341909
transform -1 0 3390 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3453_
timestamp 1728341909
transform 1 0 3250 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3454_
timestamp 1728341909
transform -1 0 3610 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3455_
timestamp 1728341909
transform 1 0 9990 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3456_
timestamp 1728341909
transform 1 0 9550 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3457_
timestamp 1728341909
transform -1 0 9830 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3458_
timestamp 1728341909
transform -1 0 9990 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3459_
timestamp 1728341909
transform 1 0 10430 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3460_
timestamp 1728341909
transform -1 0 10730 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3461_
timestamp 1728341909
transform -1 0 10490 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3462_
timestamp 1728341909
transform -1 0 10050 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3463_
timestamp 1728341909
transform 1 0 10450 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3464_
timestamp 1728341909
transform -1 0 10250 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3465_
timestamp 1728341909
transform 1 0 10210 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4__3466_
timestamp 1728341909
transform -1 0 10230 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3467_
timestamp 1728341909
transform 1 0 8290 0 1 6010
box -12 -8 32 252
use FILL  FILL_4__3468_
timestamp 1728341909
transform 1 0 9130 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__3469_
timestamp 1728341909
transform 1 0 8590 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3470_
timestamp 1728341909
transform -1 0 8530 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3471_
timestamp 1728341909
transform 1 0 8670 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__3472_
timestamp 1728341909
transform 1 0 8910 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__3473_
timestamp 1728341909
transform -1 0 8730 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3474_
timestamp 1728341909
transform -1 0 8850 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3475_
timestamp 1728341909
transform -1 0 8970 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3476_
timestamp 1728341909
transform 1 0 9770 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3477_
timestamp 1728341909
transform 1 0 9210 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3478_
timestamp 1728341909
transform -1 0 9090 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3479_
timestamp 1728341909
transform 1 0 10570 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__3480_
timestamp 1728341909
transform -1 0 10130 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__3481_
timestamp 1728341909
transform -1 0 9990 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3482_
timestamp 1728341909
transform -1 0 9790 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__3483_
timestamp 1728341909
transform 1 0 10930 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3484_
timestamp 1728341909
transform 1 0 10910 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3485_
timestamp 1728341909
transform 1 0 11190 0 1 6490
box -12 -8 32 252
use FILL  FILL_4__3486_
timestamp 1728341909
transform 1 0 11150 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3487_
timestamp 1728341909
transform 1 0 10910 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3488_
timestamp 1728341909
transform 1 0 9550 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3489_
timestamp 1728341909
transform 1 0 9450 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3490_
timestamp 1728341909
transform -1 0 9710 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3491_
timestamp 1728341909
transform -1 0 9730 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3492_
timestamp 1728341909
transform 1 0 9930 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3493_
timestamp 1728341909
transform 1 0 10190 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3494_
timestamp 1728341909
transform 1 0 10330 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__3495_
timestamp 1728341909
transform -1 0 8830 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3496_
timestamp 1728341909
transform 1 0 9450 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3497_
timestamp 1728341909
transform 1 0 9970 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3498_
timestamp 1728341909
transform 1 0 9830 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__3499_
timestamp 1728341909
transform 1 0 9250 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3500_
timestamp 1728341909
transform -1 0 9510 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3501_
timestamp 1728341909
transform -1 0 9750 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3502_
timestamp 1728341909
transform 1 0 9590 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__3503_
timestamp 1728341909
transform 1 0 10070 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__3504_
timestamp 1728341909
transform -1 0 10030 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3505_
timestamp 1728341909
transform 1 0 10270 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3506_
timestamp 1728341909
transform 1 0 10790 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__3507_
timestamp 1728341909
transform -1 0 9410 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__3508_
timestamp 1728341909
transform -1 0 8530 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3509_
timestamp 1728341909
transform 1 0 8450 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__3510_
timestamp 1728341909
transform 1 0 9230 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3511_
timestamp 1728341909
transform -1 0 8990 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3512_
timestamp 1728341909
transform 1 0 8730 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3513_
timestamp 1728341909
transform -1 0 9010 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3514_
timestamp 1728341909
transform -1 0 8770 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3515_
timestamp 1728341909
transform -1 0 9170 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__3516_
timestamp 1728341909
transform 1 0 11010 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__3517_
timestamp 1728341909
transform -1 0 10330 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__3518_
timestamp 1728341909
transform 1 0 10410 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3519_
timestamp 1728341909
transform 1 0 10890 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3520_
timestamp 1728341909
transform -1 0 11190 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3521_
timestamp 1728341909
transform 1 0 7510 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3522_
timestamp 1728341909
transform -1 0 8030 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3523_
timestamp 1728341909
transform 1 0 8770 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3524_
timestamp 1728341909
transform 1 0 8550 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3525_
timestamp 1728341909
transform 1 0 8970 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3526_
timestamp 1728341909
transform -1 0 9250 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3527_
timestamp 1728341909
transform -1 0 8310 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3528_
timestamp 1728341909
transform -1 0 9950 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3529_
timestamp 1728341909
transform 1 0 10050 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__3530_
timestamp 1728341909
transform 1 0 10150 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3531_
timestamp 1728341909
transform -1 0 10190 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3532_
timestamp 1728341909
transform 1 0 10330 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__3533_
timestamp 1728341909
transform -1 0 8250 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3534_
timestamp 1728341909
transform -1 0 8510 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3535_
timestamp 1728341909
transform -1 0 8070 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3536_
timestamp 1728341909
transform -1 0 8290 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3537_
timestamp 1728341909
transform 1 0 8390 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__3538_
timestamp 1728341909
transform -1 0 8670 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__3539_
timestamp 1728341909
transform -1 0 9570 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__3540_
timestamp 1728341909
transform 1 0 9790 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__3541_
timestamp 1728341909
transform -1 0 9870 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__3542_
timestamp 1728341909
transform -1 0 7530 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3543_
timestamp 1728341909
transform -1 0 7790 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3544_
timestamp 1728341909
transform 1 0 8010 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3545_
timestamp 1728341909
transform 1 0 8870 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__3546_
timestamp 1728341909
transform -1 0 8310 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3547_
timestamp 1728341909
transform 1 0 8730 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3548_
timestamp 1728341909
transform -1 0 8990 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3549_
timestamp 1728341909
transform -1 0 8950 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__3550_
timestamp 1728341909
transform 1 0 8930 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3551_
timestamp 1728341909
transform 1 0 9210 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3552_
timestamp 1728341909
transform 1 0 9350 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__3553_
timestamp 1728341909
transform 1 0 9090 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__3554_
timestamp 1728341909
transform 1 0 9010 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__3555_
timestamp 1728341909
transform -1 0 8590 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3556_
timestamp 1728341909
transform 1 0 8490 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3557_
timestamp 1728341909
transform -1 0 8150 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__3558_
timestamp 1728341909
transform -1 0 7790 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3559_
timestamp 1728341909
transform 1 0 7750 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3560_
timestamp 1728341909
transform 1 0 8270 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3561_
timestamp 1728341909
transform -1 0 8010 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3562_
timestamp 1728341909
transform -1 0 9010 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3563_
timestamp 1728341909
transform -1 0 8990 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__3564_
timestamp 1728341909
transform 1 0 10090 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__3565_
timestamp 1728341909
transform -1 0 10010 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__3566_
timestamp 1728341909
transform 1 0 9930 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3567_
timestamp 1728341909
transform 1 0 10010 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__3568_
timestamp 1728341909
transform 1 0 10230 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__3569_
timestamp 1728341909
transform 1 0 10230 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__3570_
timestamp 1728341909
transform 1 0 10690 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__3571_
timestamp 1728341909
transform -1 0 10670 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3572_
timestamp 1728341909
transform -1 0 11170 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3573_
timestamp 1728341909
transform 1 0 11050 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__3574_
timestamp 1728341909
transform 1 0 10790 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__3575_
timestamp 1728341909
transform 1 0 11190 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__3576_
timestamp 1728341909
transform 1 0 9970 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__3577_
timestamp 1728341909
transform -1 0 11210 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__3578_
timestamp 1728341909
transform 1 0 10810 0 -1 9850
box -12 -8 32 252
use FILL  FILL_4__3579_
timestamp 1728341909
transform -1 0 10510 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__3580_
timestamp 1728341909
transform -1 0 9210 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3581_
timestamp 1728341909
transform -1 0 8910 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__3582_
timestamp 1728341909
transform 1 0 8750 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__3583_
timestamp 1728341909
transform -1 0 9070 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__3584_
timestamp 1728341909
transform 1 0 8810 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__3585_
timestamp 1728341909
transform -1 0 9550 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__3586_
timestamp 1728341909
transform 1 0 9130 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__3587_
timestamp 1728341909
transform -1 0 9270 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__3588_
timestamp 1728341909
transform 1 0 9290 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__3589_
timestamp 1728341909
transform 1 0 10010 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__3590_
timestamp 1728341909
transform -1 0 10270 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__3591_
timestamp 1728341909
transform 1 0 9750 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__3592_
timestamp 1728341909
transform 1 0 9770 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__3593_
timestamp 1728341909
transform -1 0 9550 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__3594_
timestamp 1728341909
transform 1 0 10390 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3595_
timestamp 1728341909
transform 1 0 10950 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__3596_
timestamp 1728341909
transform -1 0 10910 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3597_
timestamp 1728341909
transform 1 0 10550 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__3598_
timestamp 1728341909
transform 1 0 11190 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__3599_
timestamp 1728341909
transform 1 0 11150 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3600_
timestamp 1728341909
transform 1 0 11030 0 -1 9370
box -12 -8 32 252
use FILL  FILL_4__3601_
timestamp 1728341909
transform 1 0 10210 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3602_
timestamp 1728341909
transform 1 0 10450 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3603_
timestamp 1728341909
transform 1 0 10510 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3604_
timestamp 1728341909
transform 1 0 10730 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3605_
timestamp 1728341909
transform 1 0 11210 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3606_
timestamp 1728341909
transform 1 0 10690 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3607_
timestamp 1728341909
transform -1 0 9990 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3608_
timestamp 1728341909
transform -1 0 10230 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3609_
timestamp 1728341909
transform 1 0 10730 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3610_
timestamp 1728341909
transform 1 0 9550 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3611_
timestamp 1728341909
transform 1 0 9350 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__3612_
timestamp 1728341909
transform 1 0 9610 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__3613_
timestamp 1728341909
transform 1 0 9470 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3614_
timestamp 1728341909
transform -1 0 9870 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__3615_
timestamp 1728341909
transform -1 0 9750 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3616_
timestamp 1728341909
transform -1 0 9050 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3617_
timestamp 1728341909
transform -1 0 9310 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3618_
timestamp 1728341909
transform 1 0 9790 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3619_
timestamp 1728341909
transform 1 0 10950 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3620_
timestamp 1728341909
transform -1 0 10690 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3621_
timestamp 1728341909
transform -1 0 10470 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3622_
timestamp 1728341909
transform 1 0 10710 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3623_
timestamp 1728341909
transform 1 0 10010 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3624_
timestamp 1728341909
transform 1 0 10730 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3625_
timestamp 1728341909
transform 1 0 10830 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__3626_
timestamp 1728341909
transform -1 0 10730 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3627_
timestamp 1728341909
transform -1 0 9710 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3628_
timestamp 1728341909
transform -1 0 10450 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3629_
timestamp 1728341909
transform 1 0 10670 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3630_
timestamp 1728341909
transform 1 0 10470 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3631_
timestamp 1728341909
transform -1 0 10630 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__3632_
timestamp 1728341909
transform -1 0 10970 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__3633_
timestamp 1728341909
transform 1 0 10930 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__3634_
timestamp 1728341909
transform -1 0 10750 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__3635_
timestamp 1728341909
transform -1 0 10470 0 1 10810
box -12 -8 32 252
use FILL  FILL_4__3636_
timestamp 1728341909
transform -1 0 10570 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__3637_
timestamp 1728341909
transform -1 0 10730 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__3638_
timestamp 1728341909
transform -1 0 10650 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3639_
timestamp 1728341909
transform -1 0 10490 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__3640_
timestamp 1728341909
transform -1 0 10950 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3641_
timestamp 1728341909
transform -1 0 10690 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3642_
timestamp 1728341909
transform -1 0 11010 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3643_
timestamp 1728341909
transform 1 0 10930 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3644_
timestamp 1728341909
transform -1 0 10490 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3645_
timestamp 1728341909
transform -1 0 10230 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3646_
timestamp 1728341909
transform -1 0 10990 0 -1 8890
box -12 -8 32 252
use FILL  FILL_4__3647_
timestamp 1728341909
transform 1 0 11090 0 1 250
box -12 -8 32 252
use FILL  FILL_4__3648_
timestamp 1728341909
transform 1 0 11170 0 1 8410
box -12 -8 32 252
use FILL  FILL_4__3649_
timestamp 1728341909
transform 1 0 10250 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3650_
timestamp 1728341909
transform 1 0 10370 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__3651_
timestamp 1728341909
transform 1 0 10470 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3652_
timestamp 1728341909
transform -1 0 10430 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3653_
timestamp 1728341909
transform 1 0 10650 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3654_
timestamp 1728341909
transform 1 0 8450 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3655_
timestamp 1728341909
transform -1 0 8710 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3656_
timestamp 1728341909
transform 1 0 8290 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__3657_
timestamp 1728341909
transform -1 0 8670 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__3658_
timestamp 1728341909
transform -1 0 8570 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__3659_
timestamp 1728341909
transform -1 0 8310 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4__3660_
timestamp 1728341909
transform -1 0 8430 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__3661_
timestamp 1728341909
transform -1 0 9290 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__3662_
timestamp 1728341909
transform -1 0 9530 0 1 10330
box -12 -8 32 252
use FILL  FILL_4__3663_
timestamp 1728341909
transform 1 0 9450 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3664_
timestamp 1728341909
transform -1 0 9690 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3665_
timestamp 1728341909
transform 1 0 8290 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3666_
timestamp 1728341909
transform -1 0 8530 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3667_
timestamp 1728341909
transform -1 0 9250 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3668_
timestamp 1728341909
transform -1 0 10470 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3669_
timestamp 1728341909
transform -1 0 10210 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3670_
timestamp 1728341909
transform -1 0 9970 0 1 9370
box -12 -8 32 252
use FILL  FILL_4__3671_
timestamp 1728341909
transform 1 0 8330 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3672_
timestamp 1728341909
transform 1 0 8570 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3673_
timestamp 1728341909
transform -1 0 9490 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3674_
timestamp 1728341909
transform -1 0 9950 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3675_
timestamp 1728341909
transform 1 0 10170 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3676_
timestamp 1728341909
transform -1 0 10210 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3677_
timestamp 1728341909
transform 1 0 9450 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3678_
timestamp 1728341909
transform -1 0 9290 0 -1 6970
box -12 -8 32 252
use FILL  FILL_4__3691_
timestamp 1728341909
transform 1 0 7770 0 1 250
box -12 -8 32 252
use FILL  FILL_4__3692_
timestamp 1728341909
transform -1 0 8030 0 1 250
box -12 -8 32 252
use FILL  FILL_4__3693_
timestamp 1728341909
transform -1 0 2010 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3694_
timestamp 1728341909
transform -1 0 110 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3695_
timestamp 1728341909
transform 1 0 610 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3696_
timestamp 1728341909
transform -1 0 110 0 1 9850
box -12 -8 32 252
use FILL  FILL_4__3697_
timestamp 1728341909
transform -1 0 110 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__3698_
timestamp 1728341909
transform -1 0 350 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4__3699_
timestamp 1728341909
transform 1 0 6170 0 1 1210
box -12 -8 32 252
use FILL  FILL_4__3700_
timestamp 1728341909
transform -1 0 6330 0 -1 730
box -12 -8 32 252
use FILL  FILL_4__3701_
timestamp 1728341909
transform -1 0 6310 0 1 250
box -12 -8 32 252
use FILL  FILL_4__3702_
timestamp 1728341909
transform -1 0 5290 0 1 5050
box -12 -8 32 252
use FILL  FILL_4__3703_
timestamp 1728341909
transform -1 0 3530 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__3704_
timestamp 1728341909
transform -1 0 3310 0 -1 250
box -12 -8 32 252
use FILL  FILL_4__3705_
timestamp 1728341909
transform -1 0 110 0 1 8890
box -12 -8 32 252
use FILL  FILL_4__3706_
timestamp 1728341909
transform -1 0 1350 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4__3707_
timestamp 1728341909
transform 1 0 11170 0 1 6970
box -12 -8 32 252
use FILL  FILL_4__3708_
timestamp 1728341909
transform 1 0 11170 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4__3709_
timestamp 1728341909
transform 1 0 11190 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3710_
timestamp 1728341909
transform 1 0 10950 0 1 7450
box -12 -8 32 252
use FILL  FILL_4__3711_
timestamp 1728341909
transform 1 0 11170 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4__3712_
timestamp 1728341909
transform 1 0 10950 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3713_
timestamp 1728341909
transform 1 0 11070 0 1 7930
box -12 -8 32 252
use FILL  FILL_4__3714_
timestamp 1728341909
transform 1 0 11190 0 -1 8410
box -12 -8 32 252
use FILL  FILL_4__3715_
timestamp 1728341909
transform 1 0 11170 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert0
timestamp 1728341909
transform 1 0 7810 0 1 10810
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert1
timestamp 1728341909
transform 1 0 9030 0 1 1690
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert2
timestamp 1728341909
transform 1 0 9230 0 1 6970
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert3
timestamp 1728341909
transform 1 0 5710 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert4
timestamp 1728341909
transform 1 0 6810 0 1 1690
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert5
timestamp 1728341909
transform -1 0 4070 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert6
timestamp 1728341909
transform 1 0 7230 0 1 10330
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert7
timestamp 1728341909
transform -1 0 4150 0 1 4090
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert8
timestamp 1728341909
transform -1 0 7590 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert9
timestamp 1728341909
transform 1 0 4510 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert10
timestamp 1728341909
transform -1 0 630 0 1 4090
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert11
timestamp 1728341909
transform -1 0 4830 0 1 2650
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert12
timestamp 1728341909
transform 1 0 790 0 1 5530
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert13
timestamp 1728341909
transform -1 0 5930 0 1 7450
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert14
timestamp 1728341909
transform 1 0 4570 0 1 2650
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert15
timestamp 1728341909
transform 1 0 5650 0 -1 5050
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert16
timestamp 1728341909
transform 1 0 2730 0 1 8410
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert17
timestamp 1728341909
transform 1 0 4230 0 1 6490
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert18
timestamp 1728341909
transform -1 0 110 0 1 2650
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert19
timestamp 1728341909
transform -1 0 370 0 1 8410
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert20
timestamp 1728341909
transform 1 0 570 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert21
timestamp 1728341909
transform -1 0 7110 0 1 4570
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert22
timestamp 1728341909
transform -1 0 10490 0 1 4090
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert23
timestamp 1728341909
transform -1 0 8830 0 1 4090
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert24
timestamp 1728341909
transform 1 0 8550 0 1 3130
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert25
timestamp 1728341909
transform -1 0 7110 0 1 3130
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert37
timestamp 1728341909
transform -1 0 1030 0 1 5530
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert38
timestamp 1728341909
transform 1 0 1310 0 1 4570
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert39
timestamp 1728341909
transform -1 0 1070 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert40
timestamp 1728341909
transform -1 0 2770 0 -1 6010
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert41
timestamp 1728341909
transform 1 0 9570 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert42
timestamp 1728341909
transform 1 0 8890 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert43
timestamp 1728341909
transform -1 0 8810 0 -1 3610
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert44
timestamp 1728341909
transform -1 0 9030 0 1 4570
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert45
timestamp 1728341909
transform 1 0 3890 0 1 4090
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert46
timestamp 1728341909
transform 1 0 5250 0 1 4090
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert47
timestamp 1728341909
transform 1 0 4350 0 1 2650
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert48
timestamp 1728341909
transform 1 0 5470 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert49
timestamp 1728341909
transform -1 0 2270 0 1 2650
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert50
timestamp 1728341909
transform 1 0 8350 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert51
timestamp 1728341909
transform -1 0 10450 0 1 4570
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert52
timestamp 1728341909
transform -1 0 9490 0 1 4570
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert53
timestamp 1728341909
transform -1 0 9570 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert54
timestamp 1728341909
transform -1 0 8410 0 -1 3130
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert55
timestamp 1728341909
transform -1 0 370 0 1 730
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert56
timestamp 1728341909
transform 1 0 5050 0 -1 1210
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert57
timestamp 1728341909
transform 1 0 4650 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert58
timestamp 1728341909
transform 1 0 1970 0 1 1690
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert59
timestamp 1728341909
transform 1 0 4410 0 1 730
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert60
timestamp 1728341909
transform -1 0 8790 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert61
timestamp 1728341909
transform 1 0 10190 0 -1 7450
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert62
timestamp 1728341909
transform 1 0 9230 0 -1 10330
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert63
timestamp 1728341909
transform 1 0 9310 0 1 7450
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert64
timestamp 1728341909
transform 1 0 8650 0 1 1210
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert65
timestamp 1728341909
transform -1 0 5050 0 1 4090
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert66
timestamp 1728341909
transform 1 0 5790 0 1 2650
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert67
timestamp 1728341909
transform 1 0 6630 0 1 5050
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert68
timestamp 1728341909
transform 1 0 7630 0 -1 2650
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert69
timestamp 1728341909
transform -1 0 6110 0 1 1690
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert70
timestamp 1728341909
transform 1 0 8790 0 -1 2170
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert71
timestamp 1728341909
transform 1 0 2490 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert72
timestamp 1728341909
transform 1 0 3930 0 1 1210
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert73
timestamp 1728341909
transform 1 0 2730 0 1 2650
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert74
timestamp 1728341909
transform -1 0 3730 0 -1 1690
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert75
timestamp 1728341909
transform -1 0 810 0 1 2170
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert76
timestamp 1728341909
transform 1 0 8790 0 1 4570
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert77
timestamp 1728341909
transform -1 0 8530 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert78
timestamp 1728341909
transform 1 0 8990 0 -1 5530
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert79
timestamp 1728341909
transform -1 0 9250 0 1 4570
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert80
timestamp 1728341909
transform 1 0 4230 0 -1 6490
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert81
timestamp 1728341909
transform 1 0 3370 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert82
timestamp 1728341909
transform 1 0 2230 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4_BUFX2_insert83
timestamp 1728341909
transform -1 0 2710 0 -1 7930
box -12 -8 32 252
use FILL  FILL_4_CLKBUF1_insert26
timestamp 1728341909
transform -1 0 1450 0 1 3130
box -12 -8 32 252
use FILL  FILL_4_CLKBUF1_insert27
timestamp 1728341909
transform 1 0 3690 0 1 3130
box -12 -8 32 252
use FILL  FILL_4_CLKBUF1_insert28
timestamp 1728341909
transform 1 0 90 0 1 3130
box -12 -8 32 252
use FILL  FILL_4_CLKBUF1_insert29
timestamp 1728341909
transform 1 0 570 0 1 7930
box -12 -8 32 252
use FILL  FILL_4_CLKBUF1_insert30
timestamp 1728341909
transform 1 0 8250 0 1 5530
box -12 -8 32 252
use FILL  FILL_4_CLKBUF1_insert31
timestamp 1728341909
transform -1 0 7610 0 -1 10810
box -12 -8 32 252
use FILL  FILL_4_CLKBUF1_insert32
timestamp 1728341909
transform -1 0 3230 0 -1 4570
box -12 -8 32 252
use FILL  FILL_4_CLKBUF1_insert33
timestamp 1728341909
transform -1 0 7970 0 1 10330
box -12 -8 32 252
use FILL  FILL_4_CLKBUF1_insert34
timestamp 1728341909
transform -1 0 110 0 -1 11290
box -12 -8 32 252
use FILL  FILL_4_CLKBUF1_insert35
timestamp 1728341909
transform -1 0 5530 0 1 5050
box -12 -8 32 252
use FILL  FILL_4_CLKBUF1_insert36
timestamp 1728341909
transform -1 0 2910 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__1744_
timestamp 1728341909
transform -1 0 4510 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__1745_
timestamp 1728341909
transform 1 0 4290 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__1746_
timestamp 1728341909
transform -1 0 4270 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__1747_
timestamp 1728341909
transform -1 0 5730 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__1748_
timestamp 1728341909
transform 1 0 6650 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__1749_
timestamp 1728341909
transform 1 0 6410 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__1750_
timestamp 1728341909
transform 1 0 5250 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__1751_
timestamp 1728341909
transform 1 0 6890 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__1752_
timestamp 1728341909
transform 1 0 5470 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__1753_
timestamp 1728341909
transform 1 0 7610 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__1754_
timestamp 1728341909
transform -1 0 7150 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__1755_
timestamp 1728341909
transform -1 0 7370 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__1756_
timestamp 1728341909
transform -1 0 6450 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__1757_
timestamp 1728341909
transform 1 0 7110 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__1758_
timestamp 1728341909
transform 1 0 6870 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__1759_
timestamp 1728341909
transform -1 0 3130 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__1760_
timestamp 1728341909
transform 1 0 2430 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__1761_
timestamp 1728341909
transform 1 0 7350 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__1762_
timestamp 1728341909
transform 1 0 2630 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__1763_
timestamp 1728341909
transform -1 0 8270 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__1764_
timestamp 1728341909
transform -1 0 8090 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__1765_
timestamp 1728341909
transform -1 0 8090 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__1766_
timestamp 1728341909
transform -1 0 7890 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__1767_
timestamp 1728341909
transform -1 0 7890 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__1768_
timestamp 1728341909
transform -1 0 5770 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__1769_
timestamp 1728341909
transform 1 0 3210 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__1770_
timestamp 1728341909
transform 1 0 10870 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__1771_
timestamp 1728341909
transform 1 0 11110 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__1772_
timestamp 1728341909
transform 1 0 10850 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__1773_
timestamp 1728341909
transform 1 0 10390 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__1774_
timestamp 1728341909
transform 1 0 10750 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1775_
timestamp 1728341909
transform -1 0 9570 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__1776_
timestamp 1728341909
transform 1 0 9610 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__1777_
timestamp 1728341909
transform -1 0 8790 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__1778_
timestamp 1728341909
transform -1 0 10990 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__1779_
timestamp 1728341909
transform 1 0 10210 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__1780_
timestamp 1728341909
transform 1 0 10970 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__1781_
timestamp 1728341909
transform -1 0 10990 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__1782_
timestamp 1728341909
transform -1 0 11230 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1783_
timestamp 1728341909
transform -1 0 10030 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1784_
timestamp 1728341909
transform 1 0 10610 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__1785_
timestamp 1728341909
transform 1 0 10950 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__1786_
timestamp 1728341909
transform -1 0 10290 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__1787_
timestamp 1728341909
transform 1 0 9290 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__1788_
timestamp 1728341909
transform 1 0 10570 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__1789_
timestamp 1728341909
transform -1 0 9430 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1790_
timestamp 1728341909
transform -1 0 10790 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1791_
timestamp 1728341909
transform 1 0 11010 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1792_
timestamp 1728341909
transform 1 0 5710 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1793_
timestamp 1728341909
transform 1 0 5430 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1794_
timestamp 1728341909
transform -1 0 5010 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1795_
timestamp 1728341909
transform 1 0 3790 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1796_
timestamp 1728341909
transform 1 0 4250 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1797_
timestamp 1728341909
transform -1 0 4770 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1798_
timestamp 1728341909
transform -1 0 11090 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__1799_
timestamp 1728341909
transform -1 0 10990 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__1800_
timestamp 1728341909
transform -1 0 10510 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__1801_
timestamp 1728341909
transform -1 0 10170 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__1802_
timestamp 1728341909
transform 1 0 10050 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__1803_
timestamp 1728341909
transform 1 0 10290 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1804_
timestamp 1728341909
transform 1 0 10290 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__1805_
timestamp 1728341909
transform -1 0 10090 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__1806_
timestamp 1728341909
transform 1 0 10030 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1807_
timestamp 1728341909
transform -1 0 10150 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1808_
timestamp 1728341909
transform -1 0 10450 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__1809_
timestamp 1728341909
transform -1 0 11110 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1810_
timestamp 1728341909
transform -1 0 6290 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1811_
timestamp 1728341909
transform -1 0 11190 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__1812_
timestamp 1728341909
transform -1 0 10270 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__1813_
timestamp 1728341909
transform -1 0 7750 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__1814_
timestamp 1728341909
transform -1 0 7590 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1815_
timestamp 1728341909
transform -1 0 11010 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1816_
timestamp 1728341909
transform -1 0 7650 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__1817_
timestamp 1728341909
transform 1 0 6770 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__1818_
timestamp 1728341909
transform 1 0 6710 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1819_
timestamp 1728341909
transform 1 0 6210 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1820_
timestamp 1728341909
transform 1 0 10410 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__1821_
timestamp 1728341909
transform -1 0 6770 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1822_
timestamp 1728341909
transform 1 0 11190 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__1823_
timestamp 1728341909
transform -1 0 10050 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__1824_
timestamp 1728341909
transform 1 0 7350 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__1825_
timestamp 1728341909
transform 1 0 6570 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1826_
timestamp 1728341909
transform 1 0 10990 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1827_
timestamp 1728341909
transform -1 0 7430 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1828_
timestamp 1728341909
transform 1 0 11190 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__1829_
timestamp 1728341909
transform -1 0 7450 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__1830_
timestamp 1728341909
transform 1 0 7590 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__1831_
timestamp 1728341909
transform 1 0 10730 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__1832_
timestamp 1728341909
transform 1 0 10710 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__1833_
timestamp 1728341909
transform 1 0 7270 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1834_
timestamp 1728341909
transform -1 0 7070 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1835_
timestamp 1728341909
transform -1 0 6510 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1836_
timestamp 1728341909
transform -1 0 6070 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1837_
timestamp 1728341909
transform -1 0 5590 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1838_
timestamp 1728341909
transform 1 0 5310 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1839_
timestamp 1728341909
transform 1 0 5890 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1840_
timestamp 1728341909
transform -1 0 8090 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__1841_
timestamp 1728341909
transform -1 0 5030 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__1842_
timestamp 1728341909
transform -1 0 6890 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__1843_
timestamp 1728341909
transform 1 0 7210 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__1844_
timestamp 1728341909
transform -1 0 10290 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__1845_
timestamp 1728341909
transform 1 0 11190 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__1846_
timestamp 1728341909
transform 1 0 11210 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1847_
timestamp 1728341909
transform -1 0 8130 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__1848_
timestamp 1728341909
transform 1 0 10730 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__1849_
timestamp 1728341909
transform -1 0 10650 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__1850_
timestamp 1728341909
transform -1 0 8590 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__1851_
timestamp 1728341909
transform -1 0 11210 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__1852_
timestamp 1728341909
transform 1 0 9770 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__1853_
timestamp 1728341909
transform 1 0 9290 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__1854_
timestamp 1728341909
transform 1 0 9090 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__1855_
timestamp 1728341909
transform 1 0 8850 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__1856_
timestamp 1728341909
transform 1 0 9370 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__1857_
timestamp 1728341909
transform 1 0 9150 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__1858_
timestamp 1728341909
transform 1 0 7330 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__1859_
timestamp 1728341909
transform -1 0 10750 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__1860_
timestamp 1728341909
transform 1 0 7130 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__1861_
timestamp 1728341909
transform 1 0 7370 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__1862_
timestamp 1728341909
transform -1 0 9870 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__1863_
timestamp 1728341909
transform 1 0 8610 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__1864_
timestamp 1728341909
transform 1 0 9910 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__1865_
timestamp 1728341909
transform 1 0 7770 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__1866_
timestamp 1728341909
transform -1 0 8950 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1867_
timestamp 1728341909
transform 1 0 9330 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__1868_
timestamp 1728341909
transform 1 0 10890 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__1869_
timestamp 1728341909
transform 1 0 9350 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__1870_
timestamp 1728341909
transform -1 0 9130 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__1871_
timestamp 1728341909
transform 1 0 8570 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__1872_
timestamp 1728341909
transform 1 0 7850 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__1873_
timestamp 1728341909
transform 1 0 6410 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1874_
timestamp 1728341909
transform -1 0 6870 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1875_
timestamp 1728341909
transform -1 0 6630 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1876_
timestamp 1728341909
transform 1 0 6690 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__1877_
timestamp 1728341909
transform -1 0 8110 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__1878_
timestamp 1728341909
transform -1 0 8370 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__1879_
timestamp 1728341909
transform -1 0 8110 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__1880_
timestamp 1728341909
transform -1 0 7050 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__1881_
timestamp 1728341909
transform -1 0 6370 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__1882_
timestamp 1728341909
transform 1 0 3530 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__1883_
timestamp 1728341909
transform -1 0 7070 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__1884_
timestamp 1728341909
transform -1 0 6590 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__1885_
timestamp 1728341909
transform 1 0 5870 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__1886_
timestamp 1728341909
transform -1 0 6270 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__1887_
timestamp 1728341909
transform 1 0 6890 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__1888_
timestamp 1728341909
transform 1 0 3650 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__1889_
timestamp 1728341909
transform -1 0 6010 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__1890_
timestamp 1728341909
transform 1 0 6470 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__1891_
timestamp 1728341909
transform -1 0 6110 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__1892_
timestamp 1728341909
transform 1 0 5670 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__1893_
timestamp 1728341909
transform 1 0 1070 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__1894_
timestamp 1728341909
transform 1 0 6010 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__1895_
timestamp 1728341909
transform 1 0 6890 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__1896_
timestamp 1728341909
transform 1 0 5210 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__1897_
timestamp 1728341909
transform 1 0 6050 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__1898_
timestamp 1728341909
transform 1 0 6470 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__1899_
timestamp 1728341909
transform 1 0 6570 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__1900_
timestamp 1728341909
transform 1 0 590 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__1901_
timestamp 1728341909
transform 1 0 8030 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__1902_
timestamp 1728341909
transform 1 0 8570 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__1903_
timestamp 1728341909
transform 1 0 7930 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__1904_
timestamp 1728341909
transform -1 0 10090 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1905_
timestamp 1728341909
transform 1 0 7590 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__1906_
timestamp 1728341909
transform 1 0 7570 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__1907_
timestamp 1728341909
transform 1 0 8710 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1908_
timestamp 1728341909
transform -1 0 7770 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1909_
timestamp 1728341909
transform 1 0 1870 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1910_
timestamp 1728341909
transform -1 0 9830 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__1911_
timestamp 1728341909
transform 1 0 9550 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1912_
timestamp 1728341909
transform 1 0 6170 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1913_
timestamp 1728341909
transform 1 0 10690 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__1914_
timestamp 1728341909
transform 1 0 10750 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1915_
timestamp 1728341909
transform -1 0 10310 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1916_
timestamp 1728341909
transform -1 0 5930 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1917_
timestamp 1728341909
transform 1 0 4070 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1918_
timestamp 1728341909
transform -1 0 850 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__1919_
timestamp 1728341909
transform -1 0 130 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__1920_
timestamp 1728341909
transform 1 0 1070 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__1921_
timestamp 1728341909
transform -1 0 1250 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1922_
timestamp 1728341909
transform -1 0 990 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1923_
timestamp 1728341909
transform 1 0 590 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__1924_
timestamp 1728341909
transform -1 0 4530 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1925_
timestamp 1728341909
transform -1 0 370 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__1926_
timestamp 1728341909
transform 1 0 830 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__1927_
timestamp 1728341909
transform -1 0 2130 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1928_
timestamp 1728341909
transform -1 0 1650 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1929_
timestamp 1728341909
transform 1 0 330 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__1930_
timestamp 1728341909
transform 1 0 710 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1931_
timestamp 1728341909
transform 1 0 590 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__1932_
timestamp 1728341909
transform -1 0 610 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1933_
timestamp 1728341909
transform 1 0 590 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__1934_
timestamp 1728341909
transform -1 0 610 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1935_
timestamp 1728341909
transform -1 0 1590 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1936_
timestamp 1728341909
transform 1 0 850 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1937_
timestamp 1728341909
transform -1 0 610 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__1938_
timestamp 1728341909
transform -1 0 130 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__1939_
timestamp 1728341909
transform 1 0 350 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__1940_
timestamp 1728341909
transform 1 0 870 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1941_
timestamp 1728341909
transform 1 0 590 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__1942_
timestamp 1728341909
transform 1 0 590 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__1943_
timestamp 1728341909
transform 1 0 8150 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__1944_
timestamp 1728341909
transform -1 0 7690 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1945_
timestamp 1728341909
transform -1 0 7470 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1946_
timestamp 1728341909
transform 1 0 8490 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1947_
timestamp 1728341909
transform -1 0 7670 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1948_
timestamp 1728341909
transform -1 0 7010 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1949_
timestamp 1728341909
transform -1 0 7250 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1950_
timestamp 1728341909
transform 1 0 8350 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__1951_
timestamp 1728341909
transform 1 0 8350 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__1952_
timestamp 1728341909
transform 1 0 9870 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1953_
timestamp 1728341909
transform -1 0 8430 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__1954_
timestamp 1728341909
transform 1 0 8270 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1955_
timestamp 1728341909
transform 1 0 6470 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__1956_
timestamp 1728341909
transform -1 0 8030 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1957_
timestamp 1728341909
transform 1 0 8110 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__1958_
timestamp 1728341909
transform 1 0 10470 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__1959_
timestamp 1728341909
transform 1 0 7830 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__1960_
timestamp 1728341909
transform 1 0 7910 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__1961_
timestamp 1728341909
transform 1 0 10730 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__1962_
timestamp 1728341909
transform 1 0 10530 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__1963_
timestamp 1728341909
transform 1 0 9870 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1964_
timestamp 1728341909
transform -1 0 7410 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__1965_
timestamp 1728341909
transform -1 0 7690 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__1966_
timestamp 1728341909
transform -1 0 3550 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__1967_
timestamp 1728341909
transform -1 0 7010 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__1968_
timestamp 1728341909
transform 1 0 7550 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__1969_
timestamp 1728341909
transform -1 0 7810 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__1970_
timestamp 1728341909
transform 1 0 1550 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__1971_
timestamp 1728341909
transform -1 0 850 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1972_
timestamp 1728341909
transform 1 0 1370 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1973_
timestamp 1728341909
transform 1 0 1630 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__1974_
timestamp 1728341909
transform 1 0 8390 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__1975_
timestamp 1728341909
transform 1 0 3010 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__1976_
timestamp 1728341909
transform -1 0 7170 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__1977_
timestamp 1728341909
transform -1 0 2870 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__1978_
timestamp 1728341909
transform -1 0 3850 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__1979_
timestamp 1728341909
transform -1 0 6550 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__1980_
timestamp 1728341909
transform 1 0 7810 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__1981_
timestamp 1728341909
transform 1 0 8330 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__1982_
timestamp 1728341909
transform -1 0 3070 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__1983_
timestamp 1728341909
transform 1 0 1750 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__1984_
timestamp 1728341909
transform 1 0 1830 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__1985_
timestamp 1728341909
transform 1 0 2490 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__1986_
timestamp 1728341909
transform -1 0 7170 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__1987_
timestamp 1728341909
transform 1 0 5110 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__1988_
timestamp 1728341909
transform -1 0 5010 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__1989_
timestamp 1728341909
transform 1 0 6770 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__1990_
timestamp 1728341909
transform -1 0 7290 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__1991_
timestamp 1728341909
transform -1 0 2090 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__1992_
timestamp 1728341909
transform -1 0 1590 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__1993_
timestamp 1728341909
transform -1 0 1870 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__1994_
timestamp 1728341909
transform 1 0 2110 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__1995_
timestamp 1728341909
transform 1 0 8070 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__1996_
timestamp 1728341909
transform -1 0 2290 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__1997_
timestamp 1728341909
transform -1 0 4010 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__1998_
timestamp 1728341909
transform -1 0 6530 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__1999_
timestamp 1728341909
transform -1 0 8250 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2000_
timestamp 1728341909
transform 1 0 1850 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2001_
timestamp 1728341909
transform 1 0 1330 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2002_
timestamp 1728341909
transform 1 0 1570 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2003_
timestamp 1728341909
transform 1 0 1590 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2004_
timestamp 1728341909
transform 1 0 7870 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2005_
timestamp 1728341909
transform 1 0 2030 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2006_
timestamp 1728341909
transform -1 0 6290 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2007_
timestamp 1728341909
transform 1 0 7570 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2008_
timestamp 1728341909
transform -1 0 8090 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2009_
timestamp 1728341909
transform 1 0 830 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2010_
timestamp 1728341909
transform -1 0 890 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2011_
timestamp 1728341909
transform 1 0 590 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2012_
timestamp 1728341909
transform 1 0 850 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2013_
timestamp 1728341909
transform 1 0 5490 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2014_
timestamp 1728341909
transform 1 0 1790 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2015_
timestamp 1728341909
transform -1 0 3990 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2016_
timestamp 1728341909
transform 1 0 6790 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2017_
timestamp 1728341909
transform -1 0 7330 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2018_
timestamp 1728341909
transform -1 0 1570 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2019_
timestamp 1728341909
transform -1 0 1630 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2020_
timestamp 1728341909
transform 1 0 1810 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2021_
timestamp 1728341909
transform 1 0 1770 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2022_
timestamp 1728341909
transform 1 0 4550 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2023_
timestamp 1728341909
transform 1 0 590 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2024_
timestamp 1728341909
transform 1 0 1490 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2025_
timestamp 1728341909
transform 1 0 2550 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2026_
timestamp 1728341909
transform -1 0 4750 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2027_
timestamp 1728341909
transform 1 0 7250 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2028_
timestamp 1728341909
transform -1 0 7530 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2029_
timestamp 1728341909
transform -1 0 130 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2030_
timestamp 1728341909
transform -1 0 610 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2031_
timestamp 1728341909
transform -1 0 370 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2032_
timestamp 1728341909
transform 1 0 590 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2033_
timestamp 1728341909
transform 1 0 7670 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2034_
timestamp 1728341909
transform 1 0 1270 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2035_
timestamp 1728341909
transform 1 0 2150 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2036_
timestamp 1728341909
transform 1 0 2950 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2037_
timestamp 1728341909
transform -1 0 4150 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2038_
timestamp 1728341909
transform 1 0 7590 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2039_
timestamp 1728341909
transform -1 0 7870 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2040_
timestamp 1728341909
transform -1 0 2990 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2041_
timestamp 1728341909
transform -1 0 610 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2042_
timestamp 1728341909
transform 1 0 1770 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__2043_
timestamp 1728341909
transform -1 0 3870 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__2044_
timestamp 1728341909
transform 1 0 5410 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2045_
timestamp 1728341909
transform -1 0 4110 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2046_
timestamp 1728341909
transform 1 0 2910 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__2047_
timestamp 1728341909
transform 1 0 2670 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__2048_
timestamp 1728341909
transform -1 0 3610 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__2049_
timestamp 1728341909
transform -1 0 3010 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__2050_
timestamp 1728341909
transform -1 0 2490 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__2051_
timestamp 1728341909
transform -1 0 2470 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2052_
timestamp 1728341909
transform -1 0 890 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2053_
timestamp 1728341909
transform -1 0 3450 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__2054_
timestamp 1728341909
transform 1 0 3170 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__2055_
timestamp 1728341909
transform -1 0 2810 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__2056_
timestamp 1728341909
transform 1 0 4430 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2057_
timestamp 1728341909
transform -1 0 3990 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2058_
timestamp 1728341909
transform 1 0 4650 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2059_
timestamp 1728341909
transform -1 0 2010 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__2060_
timestamp 1728341909
transform -1 0 3830 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__2061_
timestamp 1728341909
transform 1 0 3570 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__2062_
timestamp 1728341909
transform -1 0 3590 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__2063_
timestamp 1728341909
transform 1 0 2530 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__2064_
timestamp 1728341909
transform -1 0 2630 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2065_
timestamp 1728341909
transform -1 0 2430 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2066_
timestamp 1728341909
transform 1 0 2490 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2067_
timestamp 1728341909
transform -1 0 2810 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__2068_
timestamp 1728341909
transform -1 0 3050 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__2069_
timestamp 1728341909
transform 1 0 2590 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__2070_
timestamp 1728341909
transform -1 0 1130 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2071_
timestamp 1728341909
transform -1 0 2850 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__2072_
timestamp 1728341909
transform -1 0 2590 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__2073_
timestamp 1728341909
transform -1 0 1330 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2074_
timestamp 1728341909
transform 1 0 3270 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__2075_
timestamp 1728341909
transform -1 0 2750 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__2076_
timestamp 1728341909
transform 1 0 2450 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__2077_
timestamp 1728341909
transform -1 0 3310 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__2078_
timestamp 1728341909
transform 1 0 2830 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__2079_
timestamp 1728341909
transform -1 0 3950 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2080_
timestamp 1728341909
transform 1 0 4170 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2081_
timestamp 1728341909
transform -1 0 3730 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2082_
timestamp 1728341909
transform 1 0 5810 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2083_
timestamp 1728341909
transform -1 0 6550 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2084_
timestamp 1728341909
transform 1 0 9970 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2085_
timestamp 1728341909
transform -1 0 10490 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2086_
timestamp 1728341909
transform 1 0 10510 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2087_
timestamp 1728341909
transform 1 0 11050 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__2088_
timestamp 1728341909
transform 1 0 10250 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2089_
timestamp 1728341909
transform -1 0 9550 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2090_
timestamp 1728341909
transform 1 0 10730 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__2091_
timestamp 1728341909
transform 1 0 11230 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__2092_
timestamp 1728341909
transform -1 0 10190 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2093_
timestamp 1728341909
transform 1 0 10250 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__2094_
timestamp 1728341909
transform -1 0 10750 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__2095_
timestamp 1728341909
transform 1 0 10810 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__2096_
timestamp 1728341909
transform -1 0 11210 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__2097_
timestamp 1728341909
transform -1 0 11150 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2098_
timestamp 1728341909
transform 1 0 10230 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2099_
timestamp 1728341909
transform 1 0 10710 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2100_
timestamp 1728341909
transform 1 0 10930 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2101_
timestamp 1728341909
transform 1 0 11170 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2102_
timestamp 1728341909
transform 1 0 4050 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__2103_
timestamp 1728341909
transform 1 0 4290 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__2104_
timestamp 1728341909
transform 1 0 3910 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2105_
timestamp 1728341909
transform -1 0 1810 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2106_
timestamp 1728341909
transform -1 0 2190 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2107_
timestamp 1728341909
transform -1 0 2710 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2108_
timestamp 1728341909
transform 1 0 1510 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2109_
timestamp 1728341909
transform -1 0 2930 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2110_
timestamp 1728341909
transform 1 0 3150 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2111_
timestamp 1728341909
transform 1 0 5350 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2112_
timestamp 1728341909
transform 1 0 11230 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__2113_
timestamp 1728341909
transform -1 0 9810 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__2114_
timestamp 1728341909
transform 1 0 9810 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2115_
timestamp 1728341909
transform -1 0 11130 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2116_
timestamp 1728341909
transform -1 0 11070 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__2117_
timestamp 1728341909
transform -1 0 10670 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__2118_
timestamp 1728341909
transform 1 0 9070 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__2119_
timestamp 1728341909
transform -1 0 11150 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__2120_
timestamp 1728341909
transform 1 0 11090 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2121_
timestamp 1728341909
transform 1 0 11190 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2122_
timestamp 1728341909
transform 1 0 10890 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2123_
timestamp 1728341909
transform 1 0 10950 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2124_
timestamp 1728341909
transform 1 0 9410 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2125_
timestamp 1728341909
transform 1 0 9530 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2126_
timestamp 1728341909
transform -1 0 9970 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2127_
timestamp 1728341909
transform 1 0 9790 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2128_
timestamp 1728341909
transform 1 0 9750 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2129_
timestamp 1728341909
transform -1 0 8970 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2130_
timestamp 1728341909
transform 1 0 9650 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2131_
timestamp 1728341909
transform 1 0 9750 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2132_
timestamp 1728341909
transform 1 0 10210 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2133_
timestamp 1728341909
transform 1 0 10370 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2134_
timestamp 1728341909
transform -1 0 10150 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2135_
timestamp 1728341909
transform 1 0 10650 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2136_
timestamp 1728341909
transform -1 0 10610 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2137_
timestamp 1728341909
transform 1 0 10850 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2138_
timestamp 1728341909
transform -1 0 10950 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2139_
timestamp 1728341909
transform -1 0 10890 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2140_
timestamp 1728341909
transform -1 0 8370 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2141_
timestamp 1728341909
transform 1 0 8610 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2142_
timestamp 1728341909
transform 1 0 1930 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2143_
timestamp 1728341909
transform -1 0 2970 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2144_
timestamp 1728341909
transform -1 0 6070 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2145_
timestamp 1728341909
transform -1 0 6270 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2146_
timestamp 1728341909
transform 1 0 5570 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2147_
timestamp 1728341909
transform -1 0 6810 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2148_
timestamp 1728341909
transform 1 0 9710 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2149_
timestamp 1728341909
transform 1 0 8790 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2150_
timestamp 1728341909
transform -1 0 8550 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2151_
timestamp 1728341909
transform 1 0 8210 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2152_
timestamp 1728341909
transform -1 0 9050 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2153_
timestamp 1728341909
transform -1 0 9150 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2154_
timestamp 1728341909
transform 1 0 8890 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__2155_
timestamp 1728341909
transform 1 0 8050 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__2156_
timestamp 1728341909
transform -1 0 8330 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__2157_
timestamp 1728341909
transform -1 0 8450 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2158_
timestamp 1728341909
transform 1 0 10370 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__2159_
timestamp 1728341909
transform 1 0 6070 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2160_
timestamp 1728341909
transform -1 0 6430 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2161_
timestamp 1728341909
transform 1 0 6630 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2162_
timestamp 1728341909
transform -1 0 7970 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2163_
timestamp 1728341909
transform -1 0 8390 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__2164_
timestamp 1728341909
transform 1 0 7150 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2165_
timestamp 1728341909
transform -1 0 7130 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2166_
timestamp 1728341909
transform -1 0 8190 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2167_
timestamp 1728341909
transform -1 0 7890 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2168_
timestamp 1728341909
transform -1 0 8150 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2169_
timestamp 1728341909
transform 1 0 8190 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2170_
timestamp 1728341909
transform -1 0 8410 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2171_
timestamp 1728341909
transform 1 0 8610 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2172_
timestamp 1728341909
transform -1 0 10470 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2173_
timestamp 1728341909
transform 1 0 10210 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2174_
timestamp 1728341909
transform 1 0 4430 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2175_
timestamp 1728341909
transform -1 0 3990 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2176_
timestamp 1728341909
transform -1 0 5450 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2177_
timestamp 1728341909
transform -1 0 6110 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2178_
timestamp 1728341909
transform -1 0 6370 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2179_
timestamp 1728341909
transform 1 0 6410 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2180_
timestamp 1728341909
transform 1 0 7210 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2181_
timestamp 1728341909
transform 1 0 7350 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__2182_
timestamp 1728341909
transform -1 0 7210 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__2183_
timestamp 1728341909
transform 1 0 6190 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2184_
timestamp 1728341909
transform 1 0 6510 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2185_
timestamp 1728341909
transform -1 0 6650 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2186_
timestamp 1728341909
transform -1 0 9090 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2187_
timestamp 1728341909
transform -1 0 9490 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2188_
timestamp 1728341909
transform 1 0 9090 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2189_
timestamp 1728341909
transform -1 0 8870 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2190_
timestamp 1728341909
transform 1 0 8550 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2191_
timestamp 1728341909
transform 1 0 8790 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2192_
timestamp 1728341909
transform 1 0 7350 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2193_
timestamp 1728341909
transform 1 0 7570 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2194_
timestamp 1728341909
transform -1 0 8690 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__2195_
timestamp 1728341909
transform -1 0 8610 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__2196_
timestamp 1728341909
transform 1 0 8650 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2197_
timestamp 1728341909
transform 1 0 8690 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2198_
timestamp 1728341909
transform -1 0 7290 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2199_
timestamp 1728341909
transform -1 0 7550 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2200_
timestamp 1728341909
transform 1 0 9070 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__2201_
timestamp 1728341909
transform 1 0 8930 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2202_
timestamp 1728341909
transform -1 0 8730 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2203_
timestamp 1728341909
transform 1 0 8450 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2204_
timestamp 1728341909
transform -1 0 8450 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2205_
timestamp 1728341909
transform 1 0 8190 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2206_
timestamp 1728341909
transform -1 0 8070 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2207_
timestamp 1728341909
transform 1 0 8570 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2208_
timestamp 1728341909
transform -1 0 8330 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2209_
timestamp 1728341909
transform -1 0 7850 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2210_
timestamp 1728341909
transform 1 0 2790 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2211_
timestamp 1728341909
transform -1 0 7250 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2212_
timestamp 1728341909
transform -1 0 7510 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2213_
timestamp 1728341909
transform -1 0 8030 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2214_
timestamp 1728341909
transform 1 0 8590 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2215_
timestamp 1728341909
transform 1 0 9290 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2216_
timestamp 1728341909
transform 1 0 9270 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2217_
timestamp 1728341909
transform -1 0 9530 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2218_
timestamp 1728341909
transform 1 0 3970 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2219_
timestamp 1728341909
transform -1 0 2290 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__2220_
timestamp 1728341909
transform -1 0 3710 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2221_
timestamp 1728341909
transform 1 0 4150 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2222_
timestamp 1728341909
transform 1 0 4370 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2223_
timestamp 1728341909
transform 1 0 4190 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2224_
timestamp 1728341909
transform -1 0 2870 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2225_
timestamp 1728341909
transform -1 0 5930 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2226_
timestamp 1728341909
transform 1 0 6050 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2227_
timestamp 1728341909
transform -1 0 7030 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2228_
timestamp 1728341909
transform 1 0 6770 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2229_
timestamp 1728341909
transform 1 0 7830 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__2230_
timestamp 1728341909
transform -1 0 6230 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__2231_
timestamp 1728341909
transform -1 0 6470 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__2232_
timestamp 1728341909
transform 1 0 6890 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2233_
timestamp 1728341909
transform 1 0 7470 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2234_
timestamp 1728341909
transform 1 0 7370 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2235_
timestamp 1728341909
transform 1 0 9450 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2236_
timestamp 1728341909
transform 1 0 10510 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2237_
timestamp 1728341909
transform 1 0 9990 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2238_
timestamp 1728341909
transform -1 0 9910 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2239_
timestamp 1728341909
transform -1 0 5870 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2240_
timestamp 1728341909
transform 1 0 2730 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2241_
timestamp 1728341909
transform -1 0 4410 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2242_
timestamp 1728341909
transform -1 0 4630 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2243_
timestamp 1728341909
transform 1 0 3410 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2244_
timestamp 1728341909
transform 1 0 5170 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2245_
timestamp 1728341909
transform 1 0 7310 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2246_
timestamp 1728341909
transform 1 0 7330 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2247_
timestamp 1728341909
transform -1 0 3290 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2248_
timestamp 1728341909
transform 1 0 3470 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2249_
timestamp 1728341909
transform 1 0 5450 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2250_
timestamp 1728341909
transform 1 0 6710 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2251_
timestamp 1728341909
transform 1 0 7230 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2252_
timestamp 1728341909
transform -1 0 9670 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__2253_
timestamp 1728341909
transform 1 0 9390 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2254_
timestamp 1728341909
transform 1 0 5670 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2255_
timestamp 1728341909
transform -1 0 7010 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2256_
timestamp 1728341909
transform 1 0 7170 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2257_
timestamp 1728341909
transform -1 0 3110 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2258_
timestamp 1728341909
transform -1 0 3070 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__2259_
timestamp 1728341909
transform 1 0 3490 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2260_
timestamp 1728341909
transform 1 0 4670 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2261_
timestamp 1728341909
transform -1 0 5670 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2262_
timestamp 1728341909
transform 1 0 4850 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2263_
timestamp 1728341909
transform 1 0 4910 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2264_
timestamp 1728341909
transform -1 0 6210 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2265_
timestamp 1728341909
transform 1 0 3510 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__2266_
timestamp 1728341909
transform 1 0 7550 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__2267_
timestamp 1728341909
transform -1 0 5450 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__2268_
timestamp 1728341909
transform -1 0 5690 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__2269_
timestamp 1728341909
transform 1 0 5450 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__2270_
timestamp 1728341909
transform -1 0 6290 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__2271_
timestamp 1728341909
transform 1 0 6010 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__2272_
timestamp 1728341909
transform 1 0 5610 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__2273_
timestamp 1728341909
transform 1 0 5430 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__2274_
timestamp 1728341909
transform 1 0 5190 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__2275_
timestamp 1728341909
transform 1 0 5670 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__2276_
timestamp 1728341909
transform -1 0 6310 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2277_
timestamp 1728341909
transform 1 0 7810 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__2278_
timestamp 1728341909
transform -1 0 7750 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2279_
timestamp 1728341909
transform 1 0 6510 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2280_
timestamp 1728341909
transform -1 0 6530 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2281_
timestamp 1728341909
transform -1 0 6290 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2282_
timestamp 1728341909
transform 1 0 6570 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2283_
timestamp 1728341909
transform 1 0 7270 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2284_
timestamp 1728341909
transform 1 0 9230 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2285_
timestamp 1728341909
transform 1 0 9670 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2286_
timestamp 1728341909
transform -1 0 2570 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__2287_
timestamp 1728341909
transform -1 0 1830 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2288_
timestamp 1728341909
transform -1 0 2270 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2289_
timestamp 1728341909
transform 1 0 2230 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2290_
timestamp 1728341909
transform -1 0 1790 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2291_
timestamp 1728341909
transform 1 0 2010 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2292_
timestamp 1728341909
transform 1 0 4130 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2293_
timestamp 1728341909
transform 1 0 4870 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2294_
timestamp 1728341909
transform 1 0 6090 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2295_
timestamp 1728341909
transform -1 0 2270 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2296_
timestamp 1728341909
transform 1 0 3710 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2297_
timestamp 1728341909
transform 1 0 2250 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2298_
timestamp 1728341909
transform 1 0 2010 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2299_
timestamp 1728341909
transform 1 0 3470 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2300_
timestamp 1728341909
transform 1 0 3210 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2301_
timestamp 1728341909
transform -1 0 3670 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2302_
timestamp 1728341909
transform 1 0 5150 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2303_
timestamp 1728341909
transform -1 0 5130 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2304_
timestamp 1728341909
transform 1 0 5370 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2305_
timestamp 1728341909
transform -1 0 1570 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2306_
timestamp 1728341909
transform 1 0 2470 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2307_
timestamp 1728341909
transform -1 0 5630 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2308_
timestamp 1728341909
transform -1 0 5630 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2309_
timestamp 1728341909
transform 1 0 4630 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2310_
timestamp 1728341909
transform 1 0 4390 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2311_
timestamp 1728341909
transform -1 0 3790 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2312_
timestamp 1728341909
transform -1 0 4030 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2313_
timestamp 1728341909
transform 1 0 5310 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2314_
timestamp 1728341909
transform 1 0 4490 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2315_
timestamp 1728341909
transform 1 0 5450 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2316_
timestamp 1728341909
transform -1 0 9890 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2317_
timestamp 1728341909
transform 1 0 11190 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2318_
timestamp 1728341909
transform -1 0 10890 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__2319_
timestamp 1728341909
transform -1 0 10510 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__2320_
timestamp 1728341909
transform 1 0 10670 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2321_
timestamp 1728341909
transform 1 0 10610 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__2322_
timestamp 1728341909
transform 1 0 10510 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__2323_
timestamp 1728341909
transform 1 0 6770 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2324_
timestamp 1728341909
transform 1 0 6970 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2325_
timestamp 1728341909
transform 1 0 9330 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2326_
timestamp 1728341909
transform -1 0 8870 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2327_
timestamp 1728341909
transform -1 0 9330 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2328_
timestamp 1728341909
transform -1 0 9570 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2329_
timestamp 1728341909
transform 1 0 9290 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2330_
timestamp 1728341909
transform -1 0 9050 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2331_
timestamp 1728341909
transform -1 0 9210 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2332_
timestamp 1728341909
transform 1 0 9190 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2333_
timestamp 1728341909
transform 1 0 9450 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2334_
timestamp 1728341909
transform -1 0 9650 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2335_
timestamp 1728341909
transform 1 0 5690 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2336_
timestamp 1728341909
transform 1 0 6210 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2337_
timestamp 1728341909
transform -1 0 5990 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2338_
timestamp 1728341909
transform -1 0 5930 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2339_
timestamp 1728341909
transform 1 0 10410 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2340_
timestamp 1728341909
transform -1 0 9290 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2341_
timestamp 1728341909
transform 1 0 9290 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2342_
timestamp 1728341909
transform 1 0 10150 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2343_
timestamp 1728341909
transform -1 0 9650 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2344_
timestamp 1728341909
transform 1 0 9750 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2345_
timestamp 1728341909
transform -1 0 6930 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2346_
timestamp 1728341909
transform 1 0 6790 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2347_
timestamp 1728341909
transform -1 0 7130 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2348_
timestamp 1728341909
transform 1 0 8130 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2349_
timestamp 1728341909
transform -1 0 7830 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2350_
timestamp 1728341909
transform 1 0 7550 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2351_
timestamp 1728341909
transform -1 0 5250 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2352_
timestamp 1728341909
transform 1 0 5850 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2353_
timestamp 1728341909
transform -1 0 4270 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2354_
timestamp 1728341909
transform 1 0 4750 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2355_
timestamp 1728341909
transform -1 0 5010 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2356_
timestamp 1728341909
transform 1 0 5950 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2357_
timestamp 1728341909
transform -1 0 5710 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2358_
timestamp 1728341909
transform 1 0 6990 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2359_
timestamp 1728341909
transform 1 0 6350 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2360_
timestamp 1728341909
transform 1 0 6590 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2361_
timestamp 1728341909
transform 1 0 7890 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__2362_
timestamp 1728341909
transform 1 0 7410 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2363_
timestamp 1728341909
transform -1 0 7510 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2364_
timestamp 1728341909
transform 1 0 8130 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__2365_
timestamp 1728341909
transform -1 0 8010 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2366_
timestamp 1728341909
transform 1 0 7770 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2367_
timestamp 1728341909
transform 1 0 8050 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2368_
timestamp 1728341909
transform 1 0 8270 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2369_
timestamp 1728341909
transform -1 0 9990 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2370_
timestamp 1728341909
transform 1 0 5410 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2371_
timestamp 1728341909
transform -1 0 8810 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2372_
timestamp 1728341909
transform -1 0 8550 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2373_
timestamp 1728341909
transform -1 0 8130 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2374_
timestamp 1728341909
transform 1 0 8130 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2375_
timestamp 1728341909
transform 1 0 6530 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2376_
timestamp 1728341909
transform 1 0 8490 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2377_
timestamp 1728341909
transform -1 0 8750 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2378_
timestamp 1728341909
transform -1 0 9050 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2379_
timestamp 1728341909
transform -1 0 6910 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2380_
timestamp 1728341909
transform -1 0 7050 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2381_
timestamp 1728341909
transform -1 0 6910 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2382_
timestamp 1728341909
transform -1 0 7990 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2383_
timestamp 1728341909
transform 1 0 7710 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2384_
timestamp 1728341909
transform 1 0 7810 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2385_
timestamp 1728341909
transform -1 0 7550 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2386_
timestamp 1728341909
transform -1 0 6670 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2387_
timestamp 1728341909
transform -1 0 6430 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2388_
timestamp 1728341909
transform -1 0 8990 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2389_
timestamp 1728341909
transform -1 0 8370 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2390_
timestamp 1728341909
transform -1 0 8310 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2391_
timestamp 1728341909
transform -1 0 9550 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2392_
timestamp 1728341909
transform 1 0 8310 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2393_
timestamp 1728341909
transform 1 0 8270 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2394_
timestamp 1728341909
transform 1 0 8910 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2395_
timestamp 1728341909
transform 1 0 8870 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2396_
timestamp 1728341909
transform 1 0 9150 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2397_
timestamp 1728341909
transform -1 0 9410 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2398_
timestamp 1728341909
transform 1 0 8790 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2399_
timestamp 1728341909
transform -1 0 7670 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2400_
timestamp 1728341909
transform 1 0 7410 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2401_
timestamp 1728341909
transform 1 0 8530 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2402_
timestamp 1728341909
transform -1 0 6470 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2403_
timestamp 1728341909
transform -1 0 6670 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2404_
timestamp 1728341909
transform -1 0 7630 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2405_
timestamp 1728341909
transform -1 0 7410 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2406_
timestamp 1728341909
transform 1 0 7130 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2407_
timestamp 1728341909
transform -1 0 6670 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2408_
timestamp 1728341909
transform -1 0 5970 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2409_
timestamp 1728341909
transform 1 0 7050 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2410_
timestamp 1728341909
transform -1 0 7330 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2411_
timestamp 1728341909
transform -1 0 6890 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2412_
timestamp 1728341909
transform -1 0 7550 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2413_
timestamp 1728341909
transform 1 0 7070 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2414_
timestamp 1728341909
transform 1 0 6890 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2415_
timestamp 1728341909
transform -1 0 8090 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2416_
timestamp 1728341909
transform 1 0 7830 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2417_
timestamp 1728341909
transform -1 0 9070 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2418_
timestamp 1728341909
transform -1 0 8850 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2419_
timestamp 1728341909
transform 1 0 7110 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2420_
timestamp 1728341909
transform 1 0 2270 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2421_
timestamp 1728341909
transform -1 0 9730 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2422_
timestamp 1728341909
transform 1 0 8310 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__2423_
timestamp 1728341909
transform 1 0 9030 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2424_
timestamp 1728341909
transform 1 0 8810 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2425_
timestamp 1728341909
transform 1 0 3210 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2426_
timestamp 1728341909
transform 1 0 8790 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2427_
timestamp 1728341909
transform 1 0 8870 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__2428_
timestamp 1728341909
transform 1 0 9270 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2429_
timestamp 1728341909
transform 1 0 9490 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2430_
timestamp 1728341909
transform 1 0 8850 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2431_
timestamp 1728341909
transform -1 0 9310 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2432_
timestamp 1728341909
transform 1 0 9530 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2433_
timestamp 1728341909
transform -1 0 9950 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2434_
timestamp 1728341909
transform -1 0 10030 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2435_
timestamp 1728341909
transform 1 0 4490 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__2436_
timestamp 1728341909
transform 1 0 9250 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2437_
timestamp 1728341909
transform 1 0 10930 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__2438_
timestamp 1728341909
transform -1 0 10990 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__2439_
timestamp 1728341909
transform -1 0 10970 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__2440_
timestamp 1728341909
transform 1 0 9090 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__2441_
timestamp 1728341909
transform -1 0 6230 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__2442_
timestamp 1728341909
transform -1 0 8310 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2443_
timestamp 1728341909
transform 1 0 3870 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2444_
timestamp 1728341909
transform -1 0 4750 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__2445_
timestamp 1728341909
transform -1 0 8650 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__2446_
timestamp 1728341909
transform 1 0 8290 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2447_
timestamp 1728341909
transform 1 0 8130 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2448_
timestamp 1728341909
transform 1 0 8530 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2449_
timestamp 1728341909
transform -1 0 8810 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2450_
timestamp 1728341909
transform -1 0 9010 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2451_
timestamp 1728341909
transform 1 0 3870 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2452_
timestamp 1728341909
transform 1 0 7650 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2453_
timestamp 1728341909
transform -1 0 6670 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2454_
timestamp 1728341909
transform -1 0 6390 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2455_
timestamp 1728341909
transform -1 0 6670 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2456_
timestamp 1728341909
transform -1 0 8790 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2457_
timestamp 1728341909
transform -1 0 9010 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2458_
timestamp 1728341909
transform -1 0 6850 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2459_
timestamp 1728341909
transform -1 0 3630 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2460_
timestamp 1728341909
transform 1 0 7150 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2461_
timestamp 1728341909
transform 1 0 7070 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2462_
timestamp 1728341909
transform -1 0 7350 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2463_
timestamp 1728341909
transform -1 0 7370 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2464_
timestamp 1728341909
transform 1 0 4530 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__2465_
timestamp 1728341909
transform -1 0 7430 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2466_
timestamp 1728341909
transform -1 0 3410 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2467_
timestamp 1728341909
transform 1 0 6230 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2468_
timestamp 1728341909
transform -1 0 6350 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2469_
timestamp 1728341909
transform -1 0 6190 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2470_
timestamp 1728341909
transform -1 0 6450 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2471_
timestamp 1728341909
transform -1 0 8110 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2472_
timestamp 1728341909
transform -1 0 6130 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2473_
timestamp 1728341909
transform -1 0 5470 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2474_
timestamp 1728341909
transform -1 0 5390 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2475_
timestamp 1728341909
transform -1 0 7850 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__2476_
timestamp 1728341909
transform -1 0 2770 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2477_
timestamp 1728341909
transform -1 0 5250 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2478_
timestamp 1728341909
transform 1 0 5330 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2479_
timestamp 1728341909
transform -1 0 8070 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2480_
timestamp 1728341909
transform 1 0 5970 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2481_
timestamp 1728341909
transform 1 0 4230 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2482_
timestamp 1728341909
transform -1 0 2510 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2483_
timestamp 1728341909
transform -1 0 4750 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2484_
timestamp 1728341909
transform -1 0 5790 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2485_
timestamp 1728341909
transform -1 0 7030 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2486_
timestamp 1728341909
transform 1 0 3150 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2487_
timestamp 1728341909
transform -1 0 5730 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2488_
timestamp 1728341909
transform 1 0 6490 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2489_
timestamp 1728341909
transform -1 0 6770 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2490_
timestamp 1728341909
transform 1 0 7750 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2491_
timestamp 1728341909
transform -1 0 7990 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2492_
timestamp 1728341909
transform -1 0 2930 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2493_
timestamp 1728341909
transform -1 0 5570 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2494_
timestamp 1728341909
transform -1 0 6650 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2495_
timestamp 1728341909
transform 1 0 6890 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2496_
timestamp 1728341909
transform 1 0 7610 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2497_
timestamp 1728341909
transform -1 0 7850 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2498_
timestamp 1728341909
transform -1 0 8830 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__2499_
timestamp 1728341909
transform 1 0 9070 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2500_
timestamp 1728341909
transform -1 0 7690 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2501_
timestamp 1728341909
transform -1 0 6810 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__2502_
timestamp 1728341909
transform -1 0 7670 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__2503_
timestamp 1728341909
transform 1 0 11170 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2504_
timestamp 1728341909
transform -1 0 4610 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2505_
timestamp 1728341909
transform -1 0 5750 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2506_
timestamp 1728341909
transform -1 0 6770 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__2507_
timestamp 1728341909
transform 1 0 5910 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2508_
timestamp 1728341909
transform 1 0 5710 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2509_
timestamp 1728341909
transform -1 0 8870 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__2510_
timestamp 1728341909
transform -1 0 8130 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__2511_
timestamp 1728341909
transform -1 0 7450 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__2512_
timestamp 1728341909
transform 1 0 7150 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__2513_
timestamp 1728341909
transform 1 0 6930 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__2514_
timestamp 1728341909
transform 1 0 7090 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__2515_
timestamp 1728341909
transform 1 0 10430 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__2516_
timestamp 1728341909
transform 1 0 8570 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2517_
timestamp 1728341909
transform 1 0 10670 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2518_
timestamp 1728341909
transform -1 0 9770 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__2519_
timestamp 1728341909
transform 1 0 10010 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__2520_
timestamp 1728341909
transform -1 0 10470 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2521_
timestamp 1728341909
transform -1 0 8570 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2522_
timestamp 1728341909
transform 1 0 6130 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2523_
timestamp 1728341909
transform 1 0 5950 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2524_
timestamp 1728341909
transform 1 0 8330 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2525_
timestamp 1728341909
transform 1 0 6830 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2526_
timestamp 1728341909
transform -1 0 7830 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2527_
timestamp 1728341909
transform 1 0 8050 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2528_
timestamp 1728341909
transform -1 0 8110 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2529_
timestamp 1728341909
transform 1 0 7890 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2530_
timestamp 1728341909
transform -1 0 7850 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2531_
timestamp 1728341909
transform -1 0 7870 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2532_
timestamp 1728341909
transform 1 0 7870 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2533_
timestamp 1728341909
transform -1 0 5530 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2534_
timestamp 1728341909
transform -1 0 5950 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2535_
timestamp 1728341909
transform -1 0 7630 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2536_
timestamp 1728341909
transform 1 0 7430 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2537_
timestamp 1728341909
transform 1 0 7350 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2538_
timestamp 1728341909
transform 1 0 8070 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2539_
timestamp 1728341909
transform 1 0 5930 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2540_
timestamp 1728341909
transform 1 0 5650 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2541_
timestamp 1728341909
transform 1 0 6170 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2542_
timestamp 1728341909
transform -1 0 6710 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2543_
timestamp 1728341909
transform -1 0 6670 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2544_
timestamp 1728341909
transform 1 0 6210 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2545_
timestamp 1728341909
transform 1 0 6910 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2546_
timestamp 1728341909
transform 1 0 6170 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2547_
timestamp 1728341909
transform 1 0 6390 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2548_
timestamp 1728341909
transform 1 0 7170 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2549_
timestamp 1728341909
transform 1 0 7430 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2550_
timestamp 1728341909
transform -1 0 7590 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2551_
timestamp 1728341909
transform -1 0 6310 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2552_
timestamp 1728341909
transform -1 0 4870 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2553_
timestamp 1728341909
transform -1 0 5910 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2554_
timestamp 1728341909
transform -1 0 5630 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2555_
timestamp 1728341909
transform 1 0 5690 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2556_
timestamp 1728341909
transform 1 0 5070 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2557_
timestamp 1728341909
transform 1 0 5810 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2558_
timestamp 1728341909
transform -1 0 6450 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2559_
timestamp 1728341909
transform 1 0 6130 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__2560_
timestamp 1728341909
transform 1 0 4390 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2561_
timestamp 1728341909
transform -1 0 5450 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2562_
timestamp 1728341909
transform 1 0 5070 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2563_
timestamp 1728341909
transform -1 0 4970 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2564_
timestamp 1728341909
transform -1 0 4630 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2565_
timestamp 1728341909
transform 1 0 4770 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2566_
timestamp 1728341909
transform -1 0 4990 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2567_
timestamp 1728341909
transform 1 0 5190 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2568_
timestamp 1728341909
transform 1 0 5330 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__2569_
timestamp 1728341909
transform -1 0 4210 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2570_
timestamp 1728341909
transform 1 0 5230 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2571_
timestamp 1728341909
transform 1 0 4350 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2572_
timestamp 1728341909
transform -1 0 4470 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2573_
timestamp 1728341909
transform 1 0 4710 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2574_
timestamp 1728341909
transform 1 0 5430 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2575_
timestamp 1728341909
transform -1 0 4990 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2576_
timestamp 1728341909
transform 1 0 5170 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2577_
timestamp 1728341909
transform 1 0 4910 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2578_
timestamp 1728341909
transform -1 0 4850 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2579_
timestamp 1728341909
transform 1 0 4710 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__2580_
timestamp 1728341909
transform 1 0 4750 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__2581_
timestamp 1728341909
transform -1 0 4190 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2582_
timestamp 1728341909
transform -1 0 3330 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2583_
timestamp 1728341909
transform 1 0 2270 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2584_
timestamp 1728341909
transform 1 0 3230 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2585_
timestamp 1728341909
transform -1 0 6390 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2586_
timestamp 1728341909
transform -1 0 3750 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2587_
timestamp 1728341909
transform -1 0 3490 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2588_
timestamp 1728341909
transform -1 0 3010 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2589_
timestamp 1728341909
transform -1 0 3010 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2590_
timestamp 1728341909
transform 1 0 3630 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__2591_
timestamp 1728341909
transform -1 0 3110 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2592_
timestamp 1728341909
transform 1 0 2610 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2593_
timestamp 1728341909
transform -1 0 2710 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2594_
timestamp 1728341909
transform -1 0 2730 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2595_
timestamp 1728341909
transform -1 0 3810 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__2596_
timestamp 1728341909
transform 1 0 3410 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2597_
timestamp 1728341909
transform 1 0 3350 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2598_
timestamp 1728341909
transform -1 0 3230 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2599_
timestamp 1728341909
transform -1 0 3230 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2600_
timestamp 1728341909
transform 1 0 2950 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2601_
timestamp 1728341909
transform -1 0 2510 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2602_
timestamp 1728341909
transform -1 0 2770 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2603_
timestamp 1728341909
transform -1 0 2370 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2604_
timestamp 1728341909
transform 1 0 2510 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2605_
timestamp 1728341909
transform -1 0 2510 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2606_
timestamp 1728341909
transform 1 0 2230 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2607_
timestamp 1728341909
transform -1 0 1590 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2608_
timestamp 1728341909
transform -1 0 1110 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2609_
timestamp 1728341909
transform 1 0 2070 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2610_
timestamp 1728341909
transform 1 0 1310 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2611_
timestamp 1728341909
transform -1 0 1290 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2612_
timestamp 1728341909
transform -1 0 1030 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2613_
timestamp 1728341909
transform -1 0 2010 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2614_
timestamp 1728341909
transform -1 0 630 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2615_
timestamp 1728341909
transform 1 0 1810 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2616_
timestamp 1728341909
transform 1 0 1550 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2617_
timestamp 1728341909
transform -1 0 1550 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2618_
timestamp 1728341909
transform -1 0 1790 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2619_
timestamp 1728341909
transform 1 0 830 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2620_
timestamp 1728341909
transform -1 0 1350 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2621_
timestamp 1728341909
transform 1 0 1090 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2622_
timestamp 1728341909
transform -1 0 1310 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2623_
timestamp 1728341909
transform 1 0 1050 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2624_
timestamp 1728341909
transform -1 0 590 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2625_
timestamp 1728341909
transform -1 0 2670 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2626_
timestamp 1728341909
transform 1 0 1690 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2627_
timestamp 1728341909
transform 1 0 1430 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2628_
timestamp 1728341909
transform 1 0 830 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2629_
timestamp 1728341909
transform -1 0 3430 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__2630_
timestamp 1728341909
transform 1 0 4290 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__2631_
timestamp 1728341909
transform -1 0 4950 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__2632_
timestamp 1728341909
transform 1 0 10930 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2633_
timestamp 1728341909
transform 1 0 3930 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2634_
timestamp 1728341909
transform 1 0 9030 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2635_
timestamp 1728341909
transform -1 0 2310 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__2636_
timestamp 1728341909
transform -1 0 9190 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__2637_
timestamp 1728341909
transform 1 0 4390 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2638_
timestamp 1728341909
transform 1 0 4890 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2639_
timestamp 1728341909
transform -1 0 9970 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__2640_
timestamp 1728341909
transform -1 0 9910 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__2641_
timestamp 1728341909
transform 1 0 10210 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2642_
timestamp 1728341909
transform -1 0 9550 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__2643_
timestamp 1728341909
transform 1 0 10950 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2644_
timestamp 1728341909
transform -1 0 9790 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2645_
timestamp 1728341909
transform -1 0 9750 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__2646_
timestamp 1728341909
transform 1 0 10150 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__2647_
timestamp 1728341909
transform -1 0 8630 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2648_
timestamp 1728341909
transform -1 0 4210 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__2649_
timestamp 1728341909
transform -1 0 5850 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2650_
timestamp 1728341909
transform 1 0 9350 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__2651_
timestamp 1728341909
transform -1 0 5730 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2652_
timestamp 1728341909
transform -1 0 7890 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__2653_
timestamp 1728341909
transform -1 0 7790 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__2654_
timestamp 1728341909
transform 1 0 4710 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2655_
timestamp 1728341909
transform -1 0 5490 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2656_
timestamp 1728341909
transform -1 0 6070 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2657_
timestamp 1728341909
transform -1 0 6810 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2658_
timestamp 1728341909
transform 1 0 6310 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2659_
timestamp 1728341909
transform 1 0 7010 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2660_
timestamp 1728341909
transform -1 0 7290 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2661_
timestamp 1728341909
transform -1 0 4510 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2662_
timestamp 1728341909
transform 1 0 4470 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2663_
timestamp 1728341909
transform 1 0 6390 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2664_
timestamp 1728341909
transform -1 0 6650 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2665_
timestamp 1728341909
transform 1 0 7150 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2666_
timestamp 1728341909
transform 1 0 6890 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2667_
timestamp 1728341909
transform 1 0 7630 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2668_
timestamp 1728341909
transform 1 0 7370 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2669_
timestamp 1728341909
transform 1 0 8030 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2670_
timestamp 1728341909
transform -1 0 4250 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2671_
timestamp 1728341909
transform -1 0 5370 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__2672_
timestamp 1728341909
transform 1 0 5270 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2673_
timestamp 1728341909
transform 1 0 7230 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2674_
timestamp 1728341909
transform -1 0 7450 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2675_
timestamp 1728341909
transform 1 0 7690 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2676_
timestamp 1728341909
transform -1 0 7630 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2677_
timestamp 1728341909
transform 1 0 7810 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2678_
timestamp 1728341909
transform 1 0 7770 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2679_
timestamp 1728341909
transform 1 0 4210 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2680_
timestamp 1728341909
transform -1 0 4470 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2681_
timestamp 1728341909
transform 1 0 6170 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2682_
timestamp 1728341909
transform 1 0 6790 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2683_
timestamp 1728341909
transform 1 0 4130 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2684_
timestamp 1728341909
transform -1 0 5790 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2685_
timestamp 1728341909
transform 1 0 5510 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2686_
timestamp 1728341909
transform -1 0 6930 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2687_
timestamp 1728341909
transform 1 0 7390 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2688_
timestamp 1728341909
transform -1 0 7530 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2689_
timestamp 1728341909
transform 1 0 6550 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2690_
timestamp 1728341909
transform 1 0 6630 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2691_
timestamp 1728341909
transform 1 0 7130 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2692_
timestamp 1728341909
transform -1 0 7270 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2693_
timestamp 1728341909
transform 1 0 5110 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2694_
timestamp 1728341909
transform -1 0 5250 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2695_
timestamp 1728341909
transform 1 0 6690 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2696_
timestamp 1728341909
transform 1 0 6630 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2697_
timestamp 1728341909
transform 1 0 7050 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2698_
timestamp 1728341909
transform 1 0 6950 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2699_
timestamp 1728341909
transform -1 0 6390 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2700_
timestamp 1728341909
transform 1 0 5450 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2701_
timestamp 1728341909
transform -1 0 5530 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2702_
timestamp 1728341909
transform -1 0 5610 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2703_
timestamp 1728341909
transform -1 0 5630 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2704_
timestamp 1728341909
transform 1 0 5690 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2705_
timestamp 1728341909
transform 1 0 5950 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2706_
timestamp 1728341909
transform -1 0 6210 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2707_
timestamp 1728341909
transform -1 0 5950 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2708_
timestamp 1728341909
transform -1 0 2350 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2709_
timestamp 1728341909
transform -1 0 5010 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2710_
timestamp 1728341909
transform -1 0 4930 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2711_
timestamp 1728341909
transform -1 0 5130 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2712_
timestamp 1728341909
transform -1 0 5710 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2713_
timestamp 1728341909
transform -1 0 5850 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2714_
timestamp 1728341909
transform -1 0 6150 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2715_
timestamp 1728341909
transform 1 0 5870 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2716_
timestamp 1728341909
transform -1 0 6710 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2717_
timestamp 1728341909
transform 1 0 6650 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2718_
timestamp 1728341909
transform 1 0 6230 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2719_
timestamp 1728341909
transform -1 0 6390 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2720_
timestamp 1728341909
transform 1 0 4690 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2721_
timestamp 1728341909
transform 1 0 4970 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2722_
timestamp 1728341909
transform 1 0 5210 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2723_
timestamp 1728341909
transform -1 0 5470 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2724_
timestamp 1728341909
transform 1 0 6190 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2725_
timestamp 1728341909
transform 1 0 6430 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2726_
timestamp 1728341909
transform -1 0 6190 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__2727_
timestamp 1728341909
transform 1 0 5890 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__2728_
timestamp 1728341909
transform -1 0 4370 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2729_
timestamp 1728341909
transform -1 0 4230 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2730_
timestamp 1728341909
transform -1 0 5270 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2731_
timestamp 1728341909
transform -1 0 5390 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2732_
timestamp 1728341909
transform -1 0 5690 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2733_
timestamp 1728341909
transform -1 0 5950 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2734_
timestamp 1728341909
transform -1 0 5270 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2735_
timestamp 1728341909
transform 1 0 5470 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2736_
timestamp 1728341909
transform -1 0 8390 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__2737_
timestamp 1728341909
transform 1 0 3790 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2738_
timestamp 1728341909
transform 1 0 3970 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2739_
timestamp 1728341909
transform -1 0 3790 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2740_
timestamp 1728341909
transform -1 0 3730 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2741_
timestamp 1728341909
transform -1 0 4070 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2742_
timestamp 1728341909
transform -1 0 4210 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2743_
timestamp 1728341909
transform 1 0 4950 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2744_
timestamp 1728341909
transform 1 0 4690 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__2745_
timestamp 1728341909
transform 1 0 5170 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2746_
timestamp 1728341909
transform 1 0 4670 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2747_
timestamp 1728341909
transform 1 0 5590 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2748_
timestamp 1728341909
transform -1 0 4990 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2749_
timestamp 1728341909
transform -1 0 5350 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2750_
timestamp 1728341909
transform -1 0 5450 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2751_
timestamp 1728341909
transform 1 0 4430 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2752_
timestamp 1728341909
transform 1 0 3930 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2753_
timestamp 1728341909
transform -1 0 3470 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2754_
timestamp 1728341909
transform -1 0 3050 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2755_
timestamp 1728341909
transform 1 0 3310 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2756_
timestamp 1728341909
transform -1 0 3690 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2757_
timestamp 1728341909
transform -1 0 3710 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2758_
timestamp 1728341909
transform -1 0 3690 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2759_
timestamp 1728341909
transform -1 0 3570 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2760_
timestamp 1728341909
transform -1 0 3610 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2761_
timestamp 1728341909
transform -1 0 3750 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2762_
timestamp 1728341909
transform -1 0 3510 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2763_
timestamp 1728341909
transform 1 0 3070 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__2764_
timestamp 1728341909
transform 1 0 3350 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__2765_
timestamp 1728341909
transform -1 0 2670 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2766_
timestamp 1728341909
transform 1 0 3750 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__2767_
timestamp 1728341909
transform -1 0 4450 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2768_
timestamp 1728341909
transform 1 0 4530 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2769_
timestamp 1728341909
transform 1 0 5190 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2770_
timestamp 1728341909
transform -1 0 4690 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2771_
timestamp 1728341909
transform -1 0 4970 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2772_
timestamp 1728341909
transform -1 0 4950 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2773_
timestamp 1728341909
transform 1 0 2710 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2774_
timestamp 1728341909
transform -1 0 2570 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__2775_
timestamp 1728341909
transform 1 0 3930 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2776_
timestamp 1728341909
transform 1 0 4450 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2777_
timestamp 1728341909
transform 1 0 5190 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2778_
timestamp 1728341909
transform -1 0 4690 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2779_
timestamp 1728341909
transform 1 0 4010 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__2780_
timestamp 1728341909
transform 1 0 2790 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__2781_
timestamp 1728341909
transform -1 0 4010 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2782_
timestamp 1728341909
transform -1 0 2810 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2783_
timestamp 1728341909
transform 1 0 2510 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2784_
timestamp 1728341909
transform 1 0 590 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2785_
timestamp 1728341909
transform -1 0 2290 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2786_
timestamp 1728341909
transform 1 0 2550 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2787_
timestamp 1728341909
transform -1 0 2970 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2788_
timestamp 1728341909
transform -1 0 2470 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2789_
timestamp 1728341909
transform -1 0 3770 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2790_
timestamp 1728341909
transform 1 0 3250 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2791_
timestamp 1728341909
transform -1 0 2990 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2792_
timestamp 1728341909
transform -1 0 2890 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2793_
timestamp 1728341909
transform -1 0 2310 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__2794_
timestamp 1728341909
transform 1 0 2190 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2795_
timestamp 1728341909
transform 1 0 830 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2796_
timestamp 1728341909
transform 1 0 1770 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2797_
timestamp 1728341909
transform -1 0 2050 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2798_
timestamp 1728341909
transform 1 0 1270 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2799_
timestamp 1728341909
transform -1 0 1550 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2800_
timestamp 1728341909
transform -1 0 1810 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2801_
timestamp 1728341909
transform 1 0 1770 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2802_
timestamp 1728341909
transform 1 0 1850 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2803_
timestamp 1728341909
transform 1 0 3330 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2804_
timestamp 1728341909
transform -1 0 490 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__2805_
timestamp 1728341909
transform 1 0 7030 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2806_
timestamp 1728341909
transform -1 0 5450 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2807_
timestamp 1728341909
transform -1 0 5050 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2808_
timestamp 1728341909
transform 1 0 3970 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2809_
timestamp 1728341909
transform -1 0 4430 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2810_
timestamp 1728341909
transform -1 0 4790 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2811_
timestamp 1728341909
transform -1 0 4650 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2812_
timestamp 1728341909
transform 1 0 4270 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2813_
timestamp 1728341909
transform 1 0 4030 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__2814_
timestamp 1728341909
transform 1 0 4150 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__2815_
timestamp 1728341909
transform -1 0 4230 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2816_
timestamp 1728341909
transform 1 0 2530 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2817_
timestamp 1728341909
transform -1 0 2810 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__2818_
timestamp 1728341909
transform 1 0 2770 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2819_
timestamp 1728341909
transform 1 0 3210 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2820_
timestamp 1728341909
transform 1 0 3450 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2821_
timestamp 1728341909
transform -1 0 3990 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2822_
timestamp 1728341909
transform -1 0 4790 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2823_
timestamp 1728341909
transform -1 0 1770 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2824_
timestamp 1728341909
transform 1 0 590 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__2825_
timestamp 1728341909
transform 1 0 570 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2826_
timestamp 1728341909
transform -1 0 730 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__2827_
timestamp 1728341909
transform 1 0 1770 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2828_
timestamp 1728341909
transform -1 0 2050 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2829_
timestamp 1728341909
transform 1 0 1290 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2830_
timestamp 1728341909
transform -1 0 1550 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2831_
timestamp 1728341909
transform -1 0 1570 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__2832_
timestamp 1728341909
transform 1 0 2070 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2833_
timestamp 1728341909
transform -1 0 1090 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__2834_
timestamp 1728341909
transform 1 0 910 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__2835_
timestamp 1728341909
transform 1 0 1150 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__2836_
timestamp 1728341909
transform 1 0 1370 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__2837_
timestamp 1728341909
transform 1 0 1690 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__2838_
timestamp 1728341909
transform -1 0 1570 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__2839_
timestamp 1728341909
transform 1 0 850 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__2840_
timestamp 1728341909
transform 1 0 1290 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2841_
timestamp 1728341909
transform 1 0 2090 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2842_
timestamp 1728341909
transform -1 0 1750 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2843_
timestamp 1728341909
transform -1 0 1850 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2844_
timestamp 1728341909
transform -1 0 1610 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__2845_
timestamp 1728341909
transform -1 0 1550 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2846_
timestamp 1728341909
transform 1 0 1330 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2847_
timestamp 1728341909
transform -1 0 1330 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__2848_
timestamp 1728341909
transform -1 0 1310 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2849_
timestamp 1728341909
transform -1 0 1610 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2850_
timestamp 1728341909
transform -1 0 1530 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2851_
timestamp 1728341909
transform -1 0 1070 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2852_
timestamp 1728341909
transform -1 0 1130 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2853_
timestamp 1728341909
transform -1 0 2330 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2854_
timestamp 1728341909
transform 1 0 810 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__2855_
timestamp 1728341909
transform 1 0 2490 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__2856_
timestamp 1728341909
transform -1 0 2010 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__2857_
timestamp 1728341909
transform -1 0 2410 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__2858_
timestamp 1728341909
transform -1 0 2310 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__2859_
timestamp 1728341909
transform -1 0 890 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2860_
timestamp 1728341909
transform 1 0 570 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2861_
timestamp 1728341909
transform -1 0 130 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2862_
timestamp 1728341909
transform -1 0 1090 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__2863_
timestamp 1728341909
transform 1 0 330 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__2864_
timestamp 1728341909
transform -1 0 370 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__2865_
timestamp 1728341909
transform 1 0 4490 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__2866_
timestamp 1728341909
transform 1 0 4510 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2867_
timestamp 1728341909
transform 1 0 5610 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__2868_
timestamp 1728341909
transform -1 0 2990 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2869_
timestamp 1728341909
transform -1 0 3270 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__2870_
timestamp 1728341909
transform -1 0 2330 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__2871_
timestamp 1728341909
transform 1 0 2350 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__2872_
timestamp 1728341909
transform -1 0 4630 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__2873_
timestamp 1728341909
transform 1 0 4370 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__2874_
timestamp 1728341909
transform -1 0 4170 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2875_
timestamp 1728341909
transform -1 0 1730 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2876_
timestamp 1728341909
transform -1 0 870 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2877_
timestamp 1728341909
transform -1 0 3530 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2878_
timestamp 1728341909
transform -1 0 3970 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2879_
timestamp 1728341909
transform -1 0 1310 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2880_
timestamp 1728341909
transform 1 0 1490 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2881_
timestamp 1728341909
transform -1 0 1810 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2882_
timestamp 1728341909
transform -1 0 2490 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2883_
timestamp 1728341909
transform 1 0 4490 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2884_
timestamp 1728341909
transform 1 0 4210 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2885_
timestamp 1728341909
transform 1 0 3150 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2886_
timestamp 1728341909
transform 1 0 4710 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2887_
timestamp 1728341909
transform 1 0 5170 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2888_
timestamp 1728341909
transform 1 0 3430 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2889_
timestamp 1728341909
transform 1 0 3650 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2890_
timestamp 1728341909
transform -1 0 4430 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2891_
timestamp 1728341909
transform -1 0 4170 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2892_
timestamp 1728341909
transform -1 0 2030 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2893_
timestamp 1728341909
transform 1 0 3710 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2894_
timestamp 1728341909
transform 1 0 3910 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2895_
timestamp 1728341909
transform 1 0 4490 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2896_
timestamp 1728341909
transform -1 0 3890 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2897_
timestamp 1728341909
transform -1 0 5890 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2898_
timestamp 1728341909
transform 1 0 5210 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2899_
timestamp 1728341909
transform 1 0 5170 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2900_
timestamp 1728341909
transform 1 0 5430 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2901_
timestamp 1728341909
transform -1 0 4910 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2902_
timestamp 1728341909
transform -1 0 1570 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2903_
timestamp 1728341909
transform 1 0 2230 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2904_
timestamp 1728341909
transform 1 0 2490 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2905_
timestamp 1728341909
transform 1 0 1290 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2906_
timestamp 1728341909
transform 1 0 1070 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2907_
timestamp 1728341909
transform 1 0 1270 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2908_
timestamp 1728341909
transform -1 0 1590 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2909_
timestamp 1728341909
transform -1 0 1810 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2910_
timestamp 1728341909
transform -1 0 1590 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2911_
timestamp 1728341909
transform -1 0 1590 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2912_
timestamp 1728341909
transform -1 0 2510 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2913_
timestamp 1728341909
transform -1 0 1750 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2914_
timestamp 1728341909
transform 1 0 2270 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2915_
timestamp 1728341909
transform 1 0 2050 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2916_
timestamp 1728341909
transform 1 0 1730 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2917_
timestamp 1728341909
transform -1 0 1810 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2918_
timestamp 1728341909
transform 1 0 1750 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2919_
timestamp 1728341909
transform -1 0 2290 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2920_
timestamp 1728341909
transform -1 0 2010 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2921_
timestamp 1728341909
transform -1 0 2070 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2922_
timestamp 1728341909
transform -1 0 1990 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2923_
timestamp 1728341909
transform -1 0 2030 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2924_
timestamp 1728341909
transform -1 0 2990 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2925_
timestamp 1728341909
transform 1 0 3470 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2926_
timestamp 1728341909
transform -1 0 2450 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2927_
timestamp 1728341909
transform -1 0 2490 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2928_
timestamp 1728341909
transform 1 0 4630 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2929_
timestamp 1728341909
transform 1 0 3470 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2930_
timestamp 1728341909
transform -1 0 2750 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2931_
timestamp 1728341909
transform -1 0 2990 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2932_
timestamp 1728341909
transform 1 0 3190 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2933_
timestamp 1728341909
transform -1 0 2750 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2934_
timestamp 1728341909
transform 1 0 2970 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2935_
timestamp 1728341909
transform -1 0 1350 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2936_
timestamp 1728341909
transform -1 0 890 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2937_
timestamp 1728341909
transform 1 0 610 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2938_
timestamp 1728341909
transform 1 0 1770 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2939_
timestamp 1728341909
transform -1 0 1550 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2940_
timestamp 1728341909
transform 1 0 3210 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2941_
timestamp 1728341909
transform 1 0 3210 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2942_
timestamp 1728341909
transform -1 0 3430 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2943_
timestamp 1728341909
transform -1 0 3270 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2944_
timestamp 1728341909
transform -1 0 3770 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2945_
timestamp 1728341909
transform 1 0 3210 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__2946_
timestamp 1728341909
transform 1 0 3650 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__2947_
timestamp 1728341909
transform 1 0 3230 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2948_
timestamp 1728341909
transform -1 0 4230 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2949_
timestamp 1728341909
transform 1 0 3190 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__2950_
timestamp 1728341909
transform 1 0 2510 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2951_
timestamp 1728341909
transform -1 0 2750 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2952_
timestamp 1728341909
transform -1 0 3030 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2953_
timestamp 1728341909
transform -1 0 2230 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2954_
timestamp 1728341909
transform -1 0 2470 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2955_
timestamp 1728341909
transform 1 0 3050 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__2956_
timestamp 1728341909
transform 1 0 3290 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__2957_
timestamp 1728341909
transform 1 0 3790 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__2958_
timestamp 1728341909
transform 1 0 2230 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__2959_
timestamp 1728341909
transform 1 0 3510 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__2960_
timestamp 1728341909
transform 1 0 3630 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__2961_
timestamp 1728341909
transform 1 0 2750 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2962_
timestamp 1728341909
transform 1 0 2490 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2963_
timestamp 1728341909
transform 1 0 3010 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2964_
timestamp 1728341909
transform 1 0 2750 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2965_
timestamp 1728341909
transform -1 0 5830 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2966_
timestamp 1728341909
transform 1 0 4150 0 1 1690
box -12 -8 32 252
use FILL  FILL_5__2967_
timestamp 1728341909
transform -1 0 4630 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2968_
timestamp 1728341909
transform -1 0 4870 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2969_
timestamp 1728341909
transform -1 0 1370 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__2970_
timestamp 1728341909
transform -1 0 1550 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__2971_
timestamp 1728341909
transform -1 0 1570 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2972_
timestamp 1728341909
transform -1 0 1310 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2973_
timestamp 1728341909
transform -1 0 1070 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__2974_
timestamp 1728341909
transform -1 0 1810 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2975_
timestamp 1728341909
transform -1 0 2030 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2976_
timestamp 1728341909
transform 1 0 3910 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2977_
timestamp 1728341909
transform -1 0 4470 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2978_
timestamp 1728341909
transform 1 0 4190 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2979_
timestamp 1728341909
transform 1 0 1570 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2980_
timestamp 1728341909
transform -1 0 1050 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2981_
timestamp 1728341909
transform -1 0 810 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2982_
timestamp 1728341909
transform 1 0 2250 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2983_
timestamp 1728341909
transform -1 0 570 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2984_
timestamp 1728341909
transform -1 0 350 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2985_
timestamp 1728341909
transform -1 0 130 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__2986_
timestamp 1728341909
transform -1 0 390 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2987_
timestamp 1728341909
transform -1 0 650 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2988_
timestamp 1728341909
transform -1 0 610 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2989_
timestamp 1728341909
transform 1 0 370 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2990_
timestamp 1728341909
transform 1 0 110 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2991_
timestamp 1728341909
transform -1 0 390 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2992_
timestamp 1728341909
transform -1 0 2050 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__2993_
timestamp 1728341909
transform -1 0 1090 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2994_
timestamp 1728341909
transform -1 0 850 0 1 730
box -12 -8 32 252
use FILL  FILL_5__2995_
timestamp 1728341909
transform 1 0 630 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__2996_
timestamp 1728341909
transform -1 0 570 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__2997_
timestamp 1728341909
transform -1 0 890 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__2998_
timestamp 1728341909
transform -1 0 130 0 1 250
box -12 -8 32 252
use FILL  FILL_5__2999_
timestamp 1728341909
transform -1 0 370 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__3000_
timestamp 1728341909
transform -1 0 130 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__3001_
timestamp 1728341909
transform -1 0 130 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__3002_
timestamp 1728341909
transform -1 0 610 0 1 730
box -12 -8 32 252
use FILL  FILL_5__3003_
timestamp 1728341909
transform -1 0 130 0 1 730
box -12 -8 32 252
use FILL  FILL_5__3004_
timestamp 1728341909
transform -1 0 870 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__3005_
timestamp 1728341909
transform 1 0 830 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__3006_
timestamp 1728341909
transform -1 0 130 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__3007_
timestamp 1728341909
transform 1 0 1830 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3008_
timestamp 1728341909
transform -1 0 1090 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__3009_
timestamp 1728341909
transform -1 0 1350 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__3010_
timestamp 1728341909
transform -1 0 1350 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__3011_
timestamp 1728341909
transform -1 0 1110 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5__3012_
timestamp 1728341909
transform -1 0 1490 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__3013_
timestamp 1728341909
transform -1 0 1270 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__3014_
timestamp 1728341909
transform 1 0 1070 0 1 250
box -12 -8 32 252
use FILL  FILL_5__3015_
timestamp 1728341909
transform -1 0 1570 0 1 250
box -12 -8 32 252
use FILL  FILL_5__3016_
timestamp 1728341909
transform -1 0 1330 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__3017_
timestamp 1728341909
transform -1 0 1310 0 1 250
box -12 -8 32 252
use FILL  FILL_5__3018_
timestamp 1728341909
transform 1 0 1090 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5__3019_
timestamp 1728341909
transform -1 0 1090 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__3020_
timestamp 1728341909
transform -1 0 3730 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3021_
timestamp 1728341909
transform -1 0 5990 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__3022_
timestamp 1728341909
transform 1 0 2830 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3023_
timestamp 1728341909
transform 1 0 2850 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3024_
timestamp 1728341909
transform 1 0 3830 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3025_
timestamp 1728341909
transform -1 0 4250 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__3026_
timestamp 1728341909
transform -1 0 3110 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3027_
timestamp 1728341909
transform -1 0 3510 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__3028_
timestamp 1728341909
transform -1 0 4030 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3029_
timestamp 1728341909
transform -1 0 4530 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3030_
timestamp 1728341909
transform 1 0 3510 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__3031_
timestamp 1728341909
transform -1 0 3790 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__3032_
timestamp 1728341909
transform -1 0 2590 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3033_
timestamp 1728341909
transform -1 0 2610 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3034_
timestamp 1728341909
transform 1 0 2750 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__3035_
timestamp 1728341909
transform -1 0 3010 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__3036_
timestamp 1728341909
transform 1 0 3330 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3037_
timestamp 1728341909
transform -1 0 3770 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__3038_
timestamp 1728341909
transform -1 0 3330 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3039_
timestamp 1728341909
transform 1 0 3070 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3040_
timestamp 1728341909
transform 1 0 2210 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__3041_
timestamp 1728341909
transform 1 0 2750 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__3042_
timestamp 1728341909
transform 1 0 7510 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__3043_
timestamp 1728341909
transform 1 0 6350 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__3044_
timestamp 1728341909
transform 1 0 5370 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__3045_
timestamp 1728341909
transform 1 0 5790 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3046_
timestamp 1728341909
transform 1 0 5510 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__3047_
timestamp 1728341909
transform 1 0 4850 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__3048_
timestamp 1728341909
transform 1 0 5190 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__3049_
timestamp 1728341909
transform 1 0 5890 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3050_
timestamp 1728341909
transform -1 0 6910 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3051_
timestamp 1728341909
transform -1 0 6370 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__3052_
timestamp 1728341909
transform 1 0 6410 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3053_
timestamp 1728341909
transform 1 0 6150 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3054_
timestamp 1728341909
transform 1 0 5890 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3055_
timestamp 1728341909
transform -1 0 5990 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3056_
timestamp 1728341909
transform 1 0 4650 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__3057_
timestamp 1728341909
transform 1 0 4410 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__3058_
timestamp 1728341909
transform -1 0 4530 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3059_
timestamp 1728341909
transform 1 0 4350 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__3060_
timestamp 1728341909
transform -1 0 4330 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__3061_
timestamp 1728341909
transform 1 0 4030 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3062_
timestamp 1728341909
transform -1 0 4850 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__3063_
timestamp 1728341909
transform 1 0 4590 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__3064_
timestamp 1728341909
transform 1 0 6050 0 1 2170
box -12 -8 32 252
use FILL  FILL_5__3065_
timestamp 1728341909
transform 1 0 5830 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__3066_
timestamp 1728341909
transform -1 0 5830 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3067_
timestamp 1728341909
transform -1 0 5970 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__3068_
timestamp 1728341909
transform -1 0 7010 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3069_
timestamp 1728341909
transform -1 0 6510 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3070_
timestamp 1728341909
transform 1 0 6150 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3071_
timestamp 1728341909
transform -1 0 6430 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3072_
timestamp 1728341909
transform 1 0 6630 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__3073_
timestamp 1728341909
transform 1 0 6390 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__3074_
timestamp 1728341909
transform 1 0 450 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__3075_
timestamp 1728341909
transform -1 0 610 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__3076_
timestamp 1728341909
transform -1 0 4310 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3077_
timestamp 1728341909
transform 1 0 2050 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3078_
timestamp 1728341909
transform -1 0 5550 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3079_
timestamp 1728341909
transform 1 0 5090 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3080_
timestamp 1728341909
transform 1 0 4290 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3081_
timestamp 1728341909
transform 1 0 5930 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__3082_
timestamp 1728341909
transform -1 0 6930 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__3083_
timestamp 1728341909
transform 1 0 6090 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__3084_
timestamp 1728341909
transform -1 0 5770 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3085_
timestamp 1728341909
transform -1 0 5050 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3086_
timestamp 1728341909
transform 1 0 5530 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3087_
timestamp 1728341909
transform -1 0 5130 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__3088_
timestamp 1728341909
transform -1 0 5670 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__3089_
timestamp 1728341909
transform -1 0 5630 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__3090_
timestamp 1728341909
transform 1 0 4810 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3091_
timestamp 1728341909
transform -1 0 4770 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3092_
timestamp 1728341909
transform 1 0 5630 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5__3093_
timestamp 1728341909
transform -1 0 4030 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__3094_
timestamp 1728341909
transform 1 0 4470 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__3095_
timestamp 1728341909
transform 1 0 4770 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__3096_
timestamp 1728341909
transform 1 0 4750 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__3097_
timestamp 1728341909
transform 1 0 4990 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__3098_
timestamp 1728341909
transform -1 0 5090 0 1 2650
box -12 -8 32 252
use FILL  FILL_5__3099_
timestamp 1728341909
transform 1 0 5230 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__3100_
timestamp 1728341909
transform -1 0 5630 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__3101_
timestamp 1728341909
transform 1 0 5170 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__3102_
timestamp 1728341909
transform 1 0 4690 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__3103_
timestamp 1728341909
transform 1 0 4910 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__3104_
timestamp 1728341909
transform -1 0 5050 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3105_
timestamp 1728341909
transform 1 0 5370 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__3106_
timestamp 1728341909
transform 1 0 8550 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__3107_
timestamp 1728341909
transform 1 0 8310 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__3108_
timestamp 1728341909
transform 1 0 8070 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__3109_
timestamp 1728341909
transform -1 0 8610 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3110_
timestamp 1728341909
transform -1 0 8370 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3111_
timestamp 1728341909
transform 1 0 4550 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3112_
timestamp 1728341909
transform 1 0 4790 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3113_
timestamp 1728341909
transform -1 0 1310 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3114_
timestamp 1728341909
transform 1 0 810 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3115_
timestamp 1728341909
transform 1 0 4490 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__3116_
timestamp 1728341909
transform -1 0 4110 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3117_
timestamp 1728341909
transform -1 0 370 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__3118_
timestamp 1728341909
transform -1 0 130 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__3119_
timestamp 1728341909
transform -1 0 4970 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__3120_
timestamp 1728341909
transform 1 0 4470 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3121_
timestamp 1728341909
transform 1 0 5210 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__3122_
timestamp 1728341909
transform -1 0 4510 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3123_
timestamp 1728341909
transform -1 0 3770 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3124_
timestamp 1728341909
transform -1 0 3990 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3125_
timestamp 1728341909
transform -1 0 3730 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3126_
timestamp 1728341909
transform 1 0 4750 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3127_
timestamp 1728341909
transform 1 0 4770 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3128_
timestamp 1728341909
transform 1 0 4690 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__3129_
timestamp 1728341909
transform 1 0 3770 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__3130_
timestamp 1728341909
transform -1 0 1870 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3131_
timestamp 1728341909
transform -1 0 1370 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3132_
timestamp 1728341909
transform 1 0 1090 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3133_
timestamp 1728341909
transform 1 0 3950 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3134_
timestamp 1728341909
transform 1 0 3530 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3135_
timestamp 1728341909
transform 1 0 3270 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3136_
timestamp 1728341909
transform 1 0 3750 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3137_
timestamp 1728341909
transform 1 0 4010 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3138_
timestamp 1728341909
transform -1 0 4050 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3139_
timestamp 1728341909
transform 1 0 1110 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3140_
timestamp 1728341909
transform 1 0 850 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3141_
timestamp 1728341909
transform -1 0 4030 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3142_
timestamp 1728341909
transform 1 0 3790 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3143_
timestamp 1728341909
transform -1 0 4230 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3144_
timestamp 1728341909
transform -1 0 3510 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3145_
timestamp 1728341909
transform 1 0 3250 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3146_
timestamp 1728341909
transform -1 0 3330 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3147_
timestamp 1728341909
transform 1 0 3570 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3148_
timestamp 1728341909
transform -1 0 3530 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3149_
timestamp 1728341909
transform -1 0 3510 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__3150_
timestamp 1728341909
transform 1 0 2090 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3151_
timestamp 1728341909
transform -1 0 2330 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3152_
timestamp 1728341909
transform 1 0 7570 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3153_
timestamp 1728341909
transform 1 0 4490 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3154_
timestamp 1728341909
transform -1 0 830 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3155_
timestamp 1728341909
transform 1 0 1050 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3156_
timestamp 1728341909
transform 1 0 3010 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3157_
timestamp 1728341909
transform -1 0 2790 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3158_
timestamp 1728341909
transform 1 0 2010 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3159_
timestamp 1728341909
transform 1 0 2550 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3160_
timestamp 1728341909
transform 1 0 3170 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3161_
timestamp 1728341909
transform -1 0 2710 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3162_
timestamp 1728341909
transform -1 0 2490 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3163_
timestamp 1728341909
transform -1 0 1590 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3164_
timestamp 1728341909
transform 1 0 1290 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3165_
timestamp 1728341909
transform -1 0 370 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3166_
timestamp 1728341909
transform -1 0 130 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3167_
timestamp 1728341909
transform 1 0 2090 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3168_
timestamp 1728341909
transform 1 0 2030 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3169_
timestamp 1728341909
transform -1 0 2330 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3170_
timestamp 1728341909
transform 1 0 2070 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3171_
timestamp 1728341909
transform -1 0 2270 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3172_
timestamp 1728341909
transform 1 0 1930 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__3173_
timestamp 1728341909
transform -1 0 1810 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3174_
timestamp 1728341909
transform -1 0 1830 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3175_
timestamp 1728341909
transform -1 0 3070 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3176_
timestamp 1728341909
transform -1 0 2870 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3177_
timestamp 1728341909
transform 1 0 2310 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3178_
timestamp 1728341909
transform 1 0 2650 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3179_
timestamp 1728341909
transform 1 0 2310 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3180_
timestamp 1728341909
transform 1 0 3250 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3181_
timestamp 1728341909
transform -1 0 2970 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3182_
timestamp 1728341909
transform -1 0 3050 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3183_
timestamp 1728341909
transform 1 0 2810 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3184_
timestamp 1728341909
transform -1 0 2570 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3185_
timestamp 1728341909
transform -1 0 2570 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3186_
timestamp 1728341909
transform 1 0 2050 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3187_
timestamp 1728341909
transform -1 0 390 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3188_
timestamp 1728341909
transform -1 0 130 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3189_
timestamp 1728341909
transform 1 0 1070 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3190_
timestamp 1728341909
transform -1 0 870 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3191_
timestamp 1728341909
transform -1 0 1130 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3192_
timestamp 1728341909
transform 1 0 1750 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3193_
timestamp 1728341909
transform 1 0 1490 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3194_
timestamp 1728341909
transform 1 0 3290 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3195_
timestamp 1728341909
transform 1 0 3250 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__3196_
timestamp 1728341909
transform 1 0 1990 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3197_
timestamp 1728341909
transform -1 0 2570 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__3198_
timestamp 1728341909
transform -1 0 2150 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3199_
timestamp 1728341909
transform -1 0 2410 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3200_
timestamp 1728341909
transform 1 0 850 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3201_
timestamp 1728341909
transform -1 0 1090 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3202_
timestamp 1728341909
transform 1 0 1090 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3203_
timestamp 1728341909
transform -1 0 1350 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3204_
timestamp 1728341909
transform -1 0 610 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3205_
timestamp 1728341909
transform -1 0 610 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3206_
timestamp 1728341909
transform 1 0 1110 0 -1 4090
box -12 -8 32 252
use FILL  FILL_5__3207_
timestamp 1728341909
transform -1 0 370 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3208_
timestamp 1728341909
transform -1 0 130 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3209_
timestamp 1728341909
transform 1 0 350 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3210_
timestamp 1728341909
transform -1 0 130 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3211_
timestamp 1728341909
transform -1 0 1610 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3212_
timestamp 1728341909
transform -1 0 1350 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3213_
timestamp 1728341909
transform 1 0 1630 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3214_
timestamp 1728341909
transform 1 0 1370 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3215_
timestamp 1728341909
transform -1 0 1330 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3216_
timestamp 1728341909
transform 1 0 1070 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3217_
timestamp 1728341909
transform -1 0 370 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3218_
timestamp 1728341909
transform -1 0 130 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3219_
timestamp 1728341909
transform -1 0 1650 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3220_
timestamp 1728341909
transform 1 0 1870 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3221_
timestamp 1728341909
transform -1 0 390 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3222_
timestamp 1728341909
transform -1 0 130 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3223_
timestamp 1728341909
transform -1 0 870 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__3224_
timestamp 1728341909
transform 1 0 590 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3225_
timestamp 1728341909
transform -1 0 370 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3226_
timestamp 1728341909
transform -1 0 130 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3227_
timestamp 1728341909
transform -1 0 390 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__3228_
timestamp 1728341909
transform -1 0 130 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__3229_
timestamp 1728341909
transform -1 0 2050 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__3230_
timestamp 1728341909
transform 1 0 1770 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__3231_
timestamp 1728341909
transform 1 0 1570 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__3232_
timestamp 1728341909
transform -1 0 1830 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__3233_
timestamp 1728341909
transform 1 0 1130 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3234_
timestamp 1728341909
transform -1 0 1410 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3235_
timestamp 1728341909
transform 1 0 1090 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3236_
timestamp 1728341909
transform 1 0 1350 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3237_
timestamp 1728341909
transform 1 0 2270 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__3238_
timestamp 1728341909
transform 1 0 2510 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5__3239_
timestamp 1728341909
transform -1 0 610 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3240_
timestamp 1728341909
transform -1 0 850 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3241_
timestamp 1728341909
transform 1 0 9750 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__3242_
timestamp 1728341909
transform -1 0 9090 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5__3243_
timestamp 1728341909
transform 1 0 9510 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__3244_
timestamp 1728341909
transform 1 0 8810 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__3245_
timestamp 1728341909
transform 1 0 9110 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3246_
timestamp 1728341909
transform -1 0 9630 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3247_
timestamp 1728341909
transform 1 0 10530 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3248_
timestamp 1728341909
transform 1 0 10790 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3249_
timestamp 1728341909
transform -1 0 9530 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__3250_
timestamp 1728341909
transform 1 0 9450 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3251_
timestamp 1728341909
transform 1 0 9290 0 1 3130
box -12 -8 32 252
use FILL  FILL_5__3252_
timestamp 1728341909
transform -1 0 9310 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__3253_
timestamp 1728341909
transform -1 0 7930 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3254_
timestamp 1728341909
transform -1 0 8190 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3255_
timestamp 1728341909
transform -1 0 9370 0 1 3610
box -12 -8 32 252
use FILL  FILL_5__3256_
timestamp 1728341909
transform 1 0 8310 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3257_
timestamp 1728341909
transform 1 0 8070 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3258_
timestamp 1728341909
transform 1 0 8610 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3259_
timestamp 1728341909
transform 1 0 9550 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3260_
timestamp 1728341909
transform -1 0 10910 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__3261_
timestamp 1728341909
transform -1 0 10450 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3262_
timestamp 1728341909
transform 1 0 10030 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3263_
timestamp 1728341909
transform 1 0 9710 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__3264_
timestamp 1728341909
transform 1 0 9050 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5__3265_
timestamp 1728341909
transform -1 0 9790 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3266_
timestamp 1728341909
transform 1 0 9810 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3267_
timestamp 1728341909
transform -1 0 9710 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3268_
timestamp 1728341909
transform -1 0 10050 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3269_
timestamp 1728341909
transform -1 0 10550 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3270_
timestamp 1728341909
transform 1 0 10270 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3271_
timestamp 1728341909
transform -1 0 10090 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5__3272_
timestamp 1728341909
transform 1 0 10310 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5__3273_
timestamp 1728341909
transform -1 0 10210 0 1 4570
box -12 -8 32 252
use FILL  FILL_5__3274_
timestamp 1728341909
transform -1 0 10310 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3275_
timestamp 1728341909
transform 1 0 9630 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__3276_
timestamp 1728341909
transform -1 0 9250 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3277_
timestamp 1728341909
transform -1 0 10710 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3278_
timestamp 1728341909
transform 1 0 10170 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3279_
timestamp 1728341909
transform -1 0 9950 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3280_
timestamp 1728341909
transform 1 0 9290 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__3281_
timestamp 1728341909
transform 1 0 9050 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__3282_
timestamp 1728341909
transform -1 0 6930 0 1 4090
box -12 -8 32 252
use FILL  FILL_5__3283_
timestamp 1728341909
transform -1 0 6870 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3284_
timestamp 1728341909
transform 1 0 6630 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5__3285_
timestamp 1728341909
transform 1 0 7070 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3286_
timestamp 1728341909
transform -1 0 7330 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3287_
timestamp 1728341909
transform -1 0 6690 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3288_
timestamp 1728341909
transform -1 0 6910 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3289_
timestamp 1728341909
transform -1 0 6870 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__3290_
timestamp 1728341909
transform 1 0 6590 0 1 5530
box -12 -8 32 252
use FILL  FILL_5__3291_
timestamp 1728341909
transform 1 0 7090 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3292_
timestamp 1728341909
transform -1 0 7350 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3293_
timestamp 1728341909
transform 1 0 7190 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3294_
timestamp 1728341909
transform 1 0 6930 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3295_
timestamp 1728341909
transform 1 0 6130 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3296_
timestamp 1728341909
transform 1 0 5870 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3297_
timestamp 1728341909
transform 1 0 5490 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3298_
timestamp 1728341909
transform 1 0 5230 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3299_
timestamp 1728341909
transform 1 0 5670 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3300_
timestamp 1728341909
transform 1 0 5430 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3301_
timestamp 1728341909
transform 1 0 6930 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5__3302_
timestamp 1728341909
transform 1 0 3010 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3303_
timestamp 1728341909
transform -1 0 3070 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3304_
timestamp 1728341909
transform 1 0 2010 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3305_
timestamp 1728341909
transform -1 0 2270 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3306_
timestamp 1728341909
transform 1 0 3930 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3307_
timestamp 1728341909
transform -1 0 4870 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3308_
timestamp 1728341909
transform -1 0 130 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__3309_
timestamp 1728341909
transform -1 0 130 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3310_
timestamp 1728341909
transform -1 0 810 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__3311_
timestamp 1728341909
transform -1 0 850 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3312_
timestamp 1728341909
transform -1 0 350 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__3313_
timestamp 1728341909
transform -1 0 390 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3314_
timestamp 1728341909
transform -1 0 130 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3315_
timestamp 1728341909
transform -1 0 130 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3316_
timestamp 1728341909
transform -1 0 630 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3317_
timestamp 1728341909
transform -1 0 850 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3449_
timestamp 1728341909
transform -1 0 3870 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3450_
timestamp 1728341909
transform 1 0 3030 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3451_
timestamp 1728341909
transform 1 0 3150 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3452_
timestamp 1728341909
transform -1 0 3410 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3453_
timestamp 1728341909
transform 1 0 3270 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3454_
timestamp 1728341909
transform -1 0 3630 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3455_
timestamp 1728341909
transform 1 0 10010 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3456_
timestamp 1728341909
transform 1 0 9570 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3457_
timestamp 1728341909
transform -1 0 9850 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3458_
timestamp 1728341909
transform -1 0 10010 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3459_
timestamp 1728341909
transform 1 0 10450 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3460_
timestamp 1728341909
transform -1 0 10750 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3461_
timestamp 1728341909
transform -1 0 10510 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3462_
timestamp 1728341909
transform -1 0 10070 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3463_
timestamp 1728341909
transform 1 0 10470 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3464_
timestamp 1728341909
transform -1 0 10270 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3465_
timestamp 1728341909
transform 1 0 10230 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5__3466_
timestamp 1728341909
transform -1 0 10250 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3467_
timestamp 1728341909
transform 1 0 8310 0 1 6010
box -12 -8 32 252
use FILL  FILL_5__3468_
timestamp 1728341909
transform 1 0 9150 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__3469_
timestamp 1728341909
transform 1 0 8610 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3470_
timestamp 1728341909
transform -1 0 8550 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3471_
timestamp 1728341909
transform 1 0 8690 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__3472_
timestamp 1728341909
transform 1 0 8930 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__3473_
timestamp 1728341909
transform -1 0 8750 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3474_
timestamp 1728341909
transform -1 0 8870 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3475_
timestamp 1728341909
transform -1 0 8990 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3476_
timestamp 1728341909
transform 1 0 9790 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3477_
timestamp 1728341909
transform 1 0 9230 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3478_
timestamp 1728341909
transform -1 0 9110 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3479_
timestamp 1728341909
transform 1 0 10590 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__3480_
timestamp 1728341909
transform -1 0 10150 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__3481_
timestamp 1728341909
transform -1 0 10010 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3482_
timestamp 1728341909
transform -1 0 9810 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__3483_
timestamp 1728341909
transform 1 0 10950 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3484_
timestamp 1728341909
transform 1 0 10930 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3485_
timestamp 1728341909
transform 1 0 11210 0 1 6490
box -12 -8 32 252
use FILL  FILL_5__3486_
timestamp 1728341909
transform 1 0 11170 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3487_
timestamp 1728341909
transform 1 0 10930 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3488_
timestamp 1728341909
transform 1 0 9570 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3489_
timestamp 1728341909
transform 1 0 9470 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3490_
timestamp 1728341909
transform -1 0 9730 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3491_
timestamp 1728341909
transform -1 0 9750 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3492_
timestamp 1728341909
transform 1 0 9950 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3493_
timestamp 1728341909
transform 1 0 10210 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3494_
timestamp 1728341909
transform 1 0 10350 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__3495_
timestamp 1728341909
transform -1 0 8850 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3496_
timestamp 1728341909
transform 1 0 9470 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3497_
timestamp 1728341909
transform 1 0 9990 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3498_
timestamp 1728341909
transform 1 0 9850 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__3499_
timestamp 1728341909
transform 1 0 9270 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3500_
timestamp 1728341909
transform -1 0 9530 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3501_
timestamp 1728341909
transform -1 0 9770 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3502_
timestamp 1728341909
transform 1 0 9610 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__3503_
timestamp 1728341909
transform 1 0 10090 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__3504_
timestamp 1728341909
transform -1 0 10050 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3505_
timestamp 1728341909
transform 1 0 10290 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3506_
timestamp 1728341909
transform 1 0 10810 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__3507_
timestamp 1728341909
transform -1 0 9430 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__3508_
timestamp 1728341909
transform -1 0 8550 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3509_
timestamp 1728341909
transform 1 0 8470 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__3510_
timestamp 1728341909
transform 1 0 9250 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3511_
timestamp 1728341909
transform -1 0 9010 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3512_
timestamp 1728341909
transform 1 0 8750 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3513_
timestamp 1728341909
transform -1 0 9030 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3514_
timestamp 1728341909
transform -1 0 8790 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3515_
timestamp 1728341909
transform -1 0 9190 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__3516_
timestamp 1728341909
transform 1 0 11030 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__3517_
timestamp 1728341909
transform -1 0 10350 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__3518_
timestamp 1728341909
transform 1 0 10430 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3519_
timestamp 1728341909
transform 1 0 10910 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3520_
timestamp 1728341909
transform -1 0 11210 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3521_
timestamp 1728341909
transform 1 0 7530 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3522_
timestamp 1728341909
transform -1 0 8050 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3523_
timestamp 1728341909
transform 1 0 8790 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3524_
timestamp 1728341909
transform 1 0 8570 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3525_
timestamp 1728341909
transform 1 0 8990 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3526_
timestamp 1728341909
transform -1 0 9270 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3527_
timestamp 1728341909
transform -1 0 8330 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3528_
timestamp 1728341909
transform -1 0 9970 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3529_
timestamp 1728341909
transform 1 0 10070 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__3530_
timestamp 1728341909
transform 1 0 10170 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3531_
timestamp 1728341909
transform -1 0 10210 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3532_
timestamp 1728341909
transform 1 0 10350 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__3533_
timestamp 1728341909
transform -1 0 8270 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3534_
timestamp 1728341909
transform -1 0 8530 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3535_
timestamp 1728341909
transform -1 0 8090 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3536_
timestamp 1728341909
transform -1 0 8310 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3537_
timestamp 1728341909
transform 1 0 8410 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__3538_
timestamp 1728341909
transform -1 0 8690 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__3539_
timestamp 1728341909
transform -1 0 9590 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__3540_
timestamp 1728341909
transform 1 0 9810 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__3541_
timestamp 1728341909
transform -1 0 9890 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__3542_
timestamp 1728341909
transform -1 0 7550 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3543_
timestamp 1728341909
transform -1 0 7810 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3544_
timestamp 1728341909
transform 1 0 8030 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3545_
timestamp 1728341909
transform 1 0 8890 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__3546_
timestamp 1728341909
transform -1 0 8330 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3547_
timestamp 1728341909
transform 1 0 8750 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3548_
timestamp 1728341909
transform -1 0 9010 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3549_
timestamp 1728341909
transform -1 0 8970 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__3550_
timestamp 1728341909
transform 1 0 8950 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3551_
timestamp 1728341909
transform 1 0 9230 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3552_
timestamp 1728341909
transform 1 0 9370 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__3553_
timestamp 1728341909
transform 1 0 9110 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__3554_
timestamp 1728341909
transform 1 0 9030 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__3555_
timestamp 1728341909
transform -1 0 8610 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3556_
timestamp 1728341909
transform 1 0 8510 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3557_
timestamp 1728341909
transform -1 0 8170 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__3558_
timestamp 1728341909
transform -1 0 7810 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3559_
timestamp 1728341909
transform 1 0 7770 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3560_
timestamp 1728341909
transform 1 0 8290 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3561_
timestamp 1728341909
transform -1 0 8030 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3562_
timestamp 1728341909
transform -1 0 9030 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3563_
timestamp 1728341909
transform -1 0 9010 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__3564_
timestamp 1728341909
transform 1 0 10110 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__3565_
timestamp 1728341909
transform -1 0 10030 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__3566_
timestamp 1728341909
transform 1 0 9950 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3567_
timestamp 1728341909
transform 1 0 10030 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__3568_
timestamp 1728341909
transform 1 0 10250 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__3569_
timestamp 1728341909
transform 1 0 10250 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__3570_
timestamp 1728341909
transform 1 0 10710 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__3571_
timestamp 1728341909
transform -1 0 10690 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3572_
timestamp 1728341909
transform -1 0 11190 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3573_
timestamp 1728341909
transform 1 0 11070 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__3574_
timestamp 1728341909
transform 1 0 10810 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__3575_
timestamp 1728341909
transform 1 0 11210 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__3576_
timestamp 1728341909
transform 1 0 9990 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__3577_
timestamp 1728341909
transform -1 0 11230 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__3578_
timestamp 1728341909
transform 1 0 10830 0 -1 9850
box -12 -8 32 252
use FILL  FILL_5__3579_
timestamp 1728341909
transform -1 0 10530 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__3580_
timestamp 1728341909
transform -1 0 9230 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3581_
timestamp 1728341909
transform -1 0 8930 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__3582_
timestamp 1728341909
transform 1 0 8770 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__3583_
timestamp 1728341909
transform -1 0 9090 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__3584_
timestamp 1728341909
transform 1 0 8830 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__3585_
timestamp 1728341909
transform -1 0 9570 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__3586_
timestamp 1728341909
transform 1 0 9150 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__3587_
timestamp 1728341909
transform -1 0 9290 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__3588_
timestamp 1728341909
transform 1 0 9310 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__3589_
timestamp 1728341909
transform 1 0 10030 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__3590_
timestamp 1728341909
transform -1 0 10290 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__3591_
timestamp 1728341909
transform 1 0 9770 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__3592_
timestamp 1728341909
transform 1 0 9790 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__3593_
timestamp 1728341909
transform -1 0 9570 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__3594_
timestamp 1728341909
transform 1 0 10410 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3595_
timestamp 1728341909
transform 1 0 10970 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__3596_
timestamp 1728341909
transform -1 0 10930 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3597_
timestamp 1728341909
transform 1 0 10570 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__3598_
timestamp 1728341909
transform 1 0 11210 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__3599_
timestamp 1728341909
transform 1 0 11170 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3600_
timestamp 1728341909
transform 1 0 11050 0 -1 9370
box -12 -8 32 252
use FILL  FILL_5__3601_
timestamp 1728341909
transform 1 0 10230 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3602_
timestamp 1728341909
transform 1 0 10470 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3603_
timestamp 1728341909
transform 1 0 10530 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3604_
timestamp 1728341909
transform 1 0 10750 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3605_
timestamp 1728341909
transform 1 0 11230 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3606_
timestamp 1728341909
transform 1 0 10710 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3607_
timestamp 1728341909
transform -1 0 10010 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3608_
timestamp 1728341909
transform -1 0 10250 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3609_
timestamp 1728341909
transform 1 0 10750 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3610_
timestamp 1728341909
transform 1 0 9570 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3611_
timestamp 1728341909
transform 1 0 9370 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__3612_
timestamp 1728341909
transform 1 0 9630 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__3613_
timestamp 1728341909
transform 1 0 9490 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3614_
timestamp 1728341909
transform -1 0 9890 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__3615_
timestamp 1728341909
transform -1 0 9770 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3616_
timestamp 1728341909
transform -1 0 9070 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3617_
timestamp 1728341909
transform -1 0 9330 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3618_
timestamp 1728341909
transform 1 0 9810 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3619_
timestamp 1728341909
transform 1 0 10970 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3620_
timestamp 1728341909
transform -1 0 10710 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3621_
timestamp 1728341909
transform -1 0 10490 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3622_
timestamp 1728341909
transform 1 0 10730 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3623_
timestamp 1728341909
transform 1 0 10030 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3624_
timestamp 1728341909
transform 1 0 10750 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3625_
timestamp 1728341909
transform 1 0 10850 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__3626_
timestamp 1728341909
transform -1 0 10750 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3627_
timestamp 1728341909
transform -1 0 9730 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3628_
timestamp 1728341909
transform -1 0 10470 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3629_
timestamp 1728341909
transform 1 0 10690 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3630_
timestamp 1728341909
transform 1 0 10490 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3631_
timestamp 1728341909
transform -1 0 10650 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__3632_
timestamp 1728341909
transform -1 0 10990 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__3633_
timestamp 1728341909
transform 1 0 10950 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__3634_
timestamp 1728341909
transform -1 0 10770 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__3635_
timestamp 1728341909
transform -1 0 10490 0 1 10810
box -12 -8 32 252
use FILL  FILL_5__3636_
timestamp 1728341909
transform -1 0 10590 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__3637_
timestamp 1728341909
transform -1 0 10750 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__3638_
timestamp 1728341909
transform -1 0 10670 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3639_
timestamp 1728341909
transform -1 0 10510 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__3640_
timestamp 1728341909
transform -1 0 10970 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3641_
timestamp 1728341909
transform -1 0 10710 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3642_
timestamp 1728341909
transform -1 0 11030 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3643_
timestamp 1728341909
transform 1 0 10950 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3644_
timestamp 1728341909
transform -1 0 10510 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3645_
timestamp 1728341909
transform -1 0 10250 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3646_
timestamp 1728341909
transform -1 0 11010 0 -1 8890
box -12 -8 32 252
use FILL  FILL_5__3647_
timestamp 1728341909
transform 1 0 11110 0 1 250
box -12 -8 32 252
use FILL  FILL_5__3648_
timestamp 1728341909
transform 1 0 11190 0 1 8410
box -12 -8 32 252
use FILL  FILL_5__3649_
timestamp 1728341909
transform 1 0 10270 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3650_
timestamp 1728341909
transform 1 0 10390 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__3651_
timestamp 1728341909
transform 1 0 10490 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3652_
timestamp 1728341909
transform -1 0 10450 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3653_
timestamp 1728341909
transform 1 0 10670 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3654_
timestamp 1728341909
transform 1 0 8470 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3655_
timestamp 1728341909
transform -1 0 8730 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3656_
timestamp 1728341909
transform 1 0 8310 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__3657_
timestamp 1728341909
transform -1 0 8690 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__3658_
timestamp 1728341909
transform -1 0 8590 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__3659_
timestamp 1728341909
transform -1 0 8330 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5__3660_
timestamp 1728341909
transform -1 0 8450 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__3661_
timestamp 1728341909
transform -1 0 9310 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__3662_
timestamp 1728341909
transform -1 0 9550 0 1 10330
box -12 -8 32 252
use FILL  FILL_5__3663_
timestamp 1728341909
transform 1 0 9470 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3664_
timestamp 1728341909
transform -1 0 9710 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3665_
timestamp 1728341909
transform 1 0 8310 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3666_
timestamp 1728341909
transform -1 0 8550 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3667_
timestamp 1728341909
transform -1 0 9270 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3668_
timestamp 1728341909
transform -1 0 10490 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3669_
timestamp 1728341909
transform -1 0 10230 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3670_
timestamp 1728341909
transform -1 0 9990 0 1 9370
box -12 -8 32 252
use FILL  FILL_5__3671_
timestamp 1728341909
transform 1 0 8350 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3672_
timestamp 1728341909
transform 1 0 8590 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3673_
timestamp 1728341909
transform -1 0 9510 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3674_
timestamp 1728341909
transform -1 0 9970 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3675_
timestamp 1728341909
transform 1 0 10190 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3676_
timestamp 1728341909
transform -1 0 10230 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3677_
timestamp 1728341909
transform 1 0 9470 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3678_
timestamp 1728341909
transform -1 0 9310 0 -1 6970
box -12 -8 32 252
use FILL  FILL_5__3691_
timestamp 1728341909
transform 1 0 7790 0 1 250
box -12 -8 32 252
use FILL  FILL_5__3692_
timestamp 1728341909
transform -1 0 8050 0 1 250
box -12 -8 32 252
use FILL  FILL_5__3693_
timestamp 1728341909
transform -1 0 2030 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3694_
timestamp 1728341909
transform -1 0 130 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3695_
timestamp 1728341909
transform 1 0 630 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3696_
timestamp 1728341909
transform -1 0 130 0 1 9850
box -12 -8 32 252
use FILL  FILL_5__3697_
timestamp 1728341909
transform -1 0 130 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__3698_
timestamp 1728341909
transform -1 0 370 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5__3699_
timestamp 1728341909
transform 1 0 6190 0 1 1210
box -12 -8 32 252
use FILL  FILL_5__3700_
timestamp 1728341909
transform -1 0 6350 0 -1 730
box -12 -8 32 252
use FILL  FILL_5__3701_
timestamp 1728341909
transform -1 0 6330 0 1 250
box -12 -8 32 252
use FILL  FILL_5__3702_
timestamp 1728341909
transform -1 0 5310 0 1 5050
box -12 -8 32 252
use FILL  FILL_5__3703_
timestamp 1728341909
transform -1 0 3550 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__3704_
timestamp 1728341909
transform -1 0 3330 0 -1 250
box -12 -8 32 252
use FILL  FILL_5__3705_
timestamp 1728341909
transform -1 0 130 0 1 8890
box -12 -8 32 252
use FILL  FILL_5__3706_
timestamp 1728341909
transform -1 0 1370 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5__3707_
timestamp 1728341909
transform 1 0 11190 0 1 6970
box -12 -8 32 252
use FILL  FILL_5__3708_
timestamp 1728341909
transform 1 0 11190 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5__3709_
timestamp 1728341909
transform 1 0 11210 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3710_
timestamp 1728341909
transform 1 0 10970 0 1 7450
box -12 -8 32 252
use FILL  FILL_5__3711_
timestamp 1728341909
transform 1 0 11190 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5__3712_
timestamp 1728341909
transform 1 0 10970 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3713_
timestamp 1728341909
transform 1 0 11090 0 1 7930
box -12 -8 32 252
use FILL  FILL_5__3714_
timestamp 1728341909
transform 1 0 11210 0 -1 8410
box -12 -8 32 252
use FILL  FILL_5__3715_
timestamp 1728341909
transform 1 0 11190 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert0
timestamp 1728341909
transform 1 0 7830 0 1 10810
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert1
timestamp 1728341909
transform 1 0 9050 0 1 1690
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert2
timestamp 1728341909
transform 1 0 9250 0 1 6970
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert3
timestamp 1728341909
transform 1 0 5730 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert4
timestamp 1728341909
transform 1 0 6830 0 1 1690
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert5
timestamp 1728341909
transform -1 0 4090 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert6
timestamp 1728341909
transform 1 0 7250 0 1 10330
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert7
timestamp 1728341909
transform -1 0 4170 0 1 4090
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert8
timestamp 1728341909
transform -1 0 7610 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert9
timestamp 1728341909
transform 1 0 4530 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert10
timestamp 1728341909
transform -1 0 650 0 1 4090
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert11
timestamp 1728341909
transform -1 0 4850 0 1 2650
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert12
timestamp 1728341909
transform 1 0 810 0 1 5530
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert13
timestamp 1728341909
transform -1 0 5950 0 1 7450
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert14
timestamp 1728341909
transform 1 0 4590 0 1 2650
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert15
timestamp 1728341909
transform 1 0 5670 0 -1 5050
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert16
timestamp 1728341909
transform 1 0 2750 0 1 8410
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert17
timestamp 1728341909
transform 1 0 4250 0 1 6490
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert18
timestamp 1728341909
transform -1 0 130 0 1 2650
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert19
timestamp 1728341909
transform -1 0 390 0 1 8410
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert20
timestamp 1728341909
transform 1 0 590 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert21
timestamp 1728341909
transform -1 0 7130 0 1 4570
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert22
timestamp 1728341909
transform -1 0 10510 0 1 4090
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert23
timestamp 1728341909
transform -1 0 8850 0 1 4090
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert24
timestamp 1728341909
transform 1 0 8570 0 1 3130
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert25
timestamp 1728341909
transform -1 0 7130 0 1 3130
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert37
timestamp 1728341909
transform -1 0 1050 0 1 5530
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert38
timestamp 1728341909
transform 1 0 1330 0 1 4570
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert39
timestamp 1728341909
transform -1 0 1090 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert40
timestamp 1728341909
transform -1 0 2790 0 -1 6010
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert41
timestamp 1728341909
transform 1 0 9590 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert42
timestamp 1728341909
transform 1 0 8910 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert43
timestamp 1728341909
transform -1 0 8830 0 -1 3610
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert44
timestamp 1728341909
transform -1 0 9050 0 1 4570
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert45
timestamp 1728341909
transform 1 0 3910 0 1 4090
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert46
timestamp 1728341909
transform 1 0 5270 0 1 4090
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert47
timestamp 1728341909
transform 1 0 4370 0 1 2650
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert48
timestamp 1728341909
transform 1 0 5490 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert49
timestamp 1728341909
transform -1 0 2290 0 1 2650
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert50
timestamp 1728341909
transform 1 0 8370 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert51
timestamp 1728341909
transform -1 0 10470 0 1 4570
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert52
timestamp 1728341909
transform -1 0 9510 0 1 4570
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert53
timestamp 1728341909
transform -1 0 9590 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert54
timestamp 1728341909
transform -1 0 8430 0 -1 3130
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert55
timestamp 1728341909
transform -1 0 390 0 1 730
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert56
timestamp 1728341909
transform 1 0 5070 0 -1 1210
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert57
timestamp 1728341909
transform 1 0 4670 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert58
timestamp 1728341909
transform 1 0 1990 0 1 1690
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert59
timestamp 1728341909
transform 1 0 4430 0 1 730
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert60
timestamp 1728341909
transform -1 0 8810 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert61
timestamp 1728341909
transform 1 0 10210 0 -1 7450
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert62
timestamp 1728341909
transform 1 0 9250 0 -1 10330
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert63
timestamp 1728341909
transform 1 0 9330 0 1 7450
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert64
timestamp 1728341909
transform 1 0 8670 0 1 1210
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert65
timestamp 1728341909
transform -1 0 5070 0 1 4090
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert66
timestamp 1728341909
transform 1 0 5810 0 1 2650
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert67
timestamp 1728341909
transform 1 0 6650 0 1 5050
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert68
timestamp 1728341909
transform 1 0 7650 0 -1 2650
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert69
timestamp 1728341909
transform -1 0 6130 0 1 1690
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert70
timestamp 1728341909
transform 1 0 8810 0 -1 2170
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert71
timestamp 1728341909
transform 1 0 2510 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert72
timestamp 1728341909
transform 1 0 3950 0 1 1210
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert73
timestamp 1728341909
transform 1 0 2750 0 1 2650
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert74
timestamp 1728341909
transform -1 0 3750 0 -1 1690
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert75
timestamp 1728341909
transform -1 0 830 0 1 2170
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert76
timestamp 1728341909
transform 1 0 8810 0 1 4570
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert77
timestamp 1728341909
transform -1 0 8550 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert78
timestamp 1728341909
transform 1 0 9010 0 -1 5530
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert79
timestamp 1728341909
transform -1 0 9270 0 1 4570
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert80
timestamp 1728341909
transform 1 0 4250 0 -1 6490
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert81
timestamp 1728341909
transform 1 0 3390 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert82
timestamp 1728341909
transform 1 0 2250 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5_BUFX2_insert83
timestamp 1728341909
transform -1 0 2730 0 -1 7930
box -12 -8 32 252
use FILL  FILL_5_CLKBUF1_insert26
timestamp 1728341909
transform -1 0 1470 0 1 3130
box -12 -8 32 252
use FILL  FILL_5_CLKBUF1_insert27
timestamp 1728341909
transform 1 0 3710 0 1 3130
box -12 -8 32 252
use FILL  FILL_5_CLKBUF1_insert28
timestamp 1728341909
transform 1 0 110 0 1 3130
box -12 -8 32 252
use FILL  FILL_5_CLKBUF1_insert29
timestamp 1728341909
transform 1 0 590 0 1 7930
box -12 -8 32 252
use FILL  FILL_5_CLKBUF1_insert30
timestamp 1728341909
transform 1 0 8270 0 1 5530
box -12 -8 32 252
use FILL  FILL_5_CLKBUF1_insert31
timestamp 1728341909
transform -1 0 7630 0 -1 10810
box -12 -8 32 252
use FILL  FILL_5_CLKBUF1_insert32
timestamp 1728341909
transform -1 0 3250 0 -1 4570
box -12 -8 32 252
use FILL  FILL_5_CLKBUF1_insert33
timestamp 1728341909
transform -1 0 7990 0 1 10330
box -12 -8 32 252
use FILL  FILL_5_CLKBUF1_insert34
timestamp 1728341909
transform -1 0 130 0 -1 11290
box -12 -8 32 252
use FILL  FILL_5_CLKBUF1_insert35
timestamp 1728341909
transform -1 0 5550 0 1 5050
box -12 -8 32 252
use FILL  FILL_5_CLKBUF1_insert36
timestamp 1728341909
transform -1 0 2930 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__1744_
timestamp 1728341909
transform -1 0 4530 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__1745_
timestamp 1728341909
transform 1 0 4310 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__1746_
timestamp 1728341909
transform -1 0 4290 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__1747_
timestamp 1728341909
transform -1 0 5750 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__1748_
timestamp 1728341909
transform 1 0 6670 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__1749_
timestamp 1728341909
transform 1 0 6430 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__1750_
timestamp 1728341909
transform 1 0 5270 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__1751_
timestamp 1728341909
transform 1 0 6910 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__1752_
timestamp 1728341909
transform 1 0 5490 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__1753_
timestamp 1728341909
transform 1 0 7630 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__1754_
timestamp 1728341909
transform -1 0 7170 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__1755_
timestamp 1728341909
transform -1 0 7390 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__1756_
timestamp 1728341909
transform -1 0 6470 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__1757_
timestamp 1728341909
transform 1 0 7130 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__1758_
timestamp 1728341909
transform 1 0 6890 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__1759_
timestamp 1728341909
transform -1 0 3150 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__1760_
timestamp 1728341909
transform 1 0 2450 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__1761_
timestamp 1728341909
transform 1 0 7370 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__1762_
timestamp 1728341909
transform 1 0 2650 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__1763_
timestamp 1728341909
transform -1 0 8290 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__1764_
timestamp 1728341909
transform -1 0 8110 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__1765_
timestamp 1728341909
transform -1 0 8110 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__1766_
timestamp 1728341909
transform -1 0 7910 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__1767_
timestamp 1728341909
transform -1 0 7910 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__1768_
timestamp 1728341909
transform -1 0 5790 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__1769_
timestamp 1728341909
transform 1 0 3230 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__1770_
timestamp 1728341909
transform 1 0 10890 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__1771_
timestamp 1728341909
transform 1 0 11130 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__1772_
timestamp 1728341909
transform 1 0 10870 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__1773_
timestamp 1728341909
transform 1 0 10410 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__1774_
timestamp 1728341909
transform 1 0 10770 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1775_
timestamp 1728341909
transform -1 0 9590 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__1776_
timestamp 1728341909
transform 1 0 9630 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__1777_
timestamp 1728341909
transform -1 0 8810 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__1778_
timestamp 1728341909
transform -1 0 11010 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__1779_
timestamp 1728341909
transform 1 0 10230 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__1780_
timestamp 1728341909
transform 1 0 10990 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__1781_
timestamp 1728341909
transform -1 0 11010 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__1782_
timestamp 1728341909
transform -1 0 11250 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1783_
timestamp 1728341909
transform -1 0 10050 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1784_
timestamp 1728341909
transform 1 0 10630 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__1785_
timestamp 1728341909
transform 1 0 10970 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__1786_
timestamp 1728341909
transform -1 0 10310 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__1787_
timestamp 1728341909
transform 1 0 9310 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__1788_
timestamp 1728341909
transform 1 0 10590 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__1789_
timestamp 1728341909
transform -1 0 9450 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1790_
timestamp 1728341909
transform -1 0 10810 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1791_
timestamp 1728341909
transform 1 0 11030 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1792_
timestamp 1728341909
transform 1 0 5730 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1793_
timestamp 1728341909
transform 1 0 5450 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1794_
timestamp 1728341909
transform -1 0 5030 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1795_
timestamp 1728341909
transform 1 0 3810 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1796_
timestamp 1728341909
transform 1 0 4270 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1797_
timestamp 1728341909
transform -1 0 4790 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1798_
timestamp 1728341909
transform -1 0 11110 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__1799_
timestamp 1728341909
transform -1 0 11010 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__1800_
timestamp 1728341909
transform -1 0 10530 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__1801_
timestamp 1728341909
transform -1 0 10190 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__1802_
timestamp 1728341909
transform 1 0 10070 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__1803_
timestamp 1728341909
transform 1 0 10310 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1804_
timestamp 1728341909
transform 1 0 10310 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__1805_
timestamp 1728341909
transform -1 0 10110 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__1806_
timestamp 1728341909
transform 1 0 10050 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1807_
timestamp 1728341909
transform -1 0 10170 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1808_
timestamp 1728341909
transform -1 0 10470 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__1809_
timestamp 1728341909
transform -1 0 11130 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1810_
timestamp 1728341909
transform -1 0 6310 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1811_
timestamp 1728341909
transform -1 0 11210 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__1812_
timestamp 1728341909
transform -1 0 10290 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__1813_
timestamp 1728341909
transform -1 0 7770 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__1814_
timestamp 1728341909
transform -1 0 7610 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1815_
timestamp 1728341909
transform -1 0 11030 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1816_
timestamp 1728341909
transform -1 0 7670 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__1817_
timestamp 1728341909
transform 1 0 6790 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__1818_
timestamp 1728341909
transform 1 0 6730 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1819_
timestamp 1728341909
transform 1 0 6230 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1820_
timestamp 1728341909
transform 1 0 10430 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__1821_
timestamp 1728341909
transform -1 0 6790 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1822_
timestamp 1728341909
transform 1 0 11210 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__1823_
timestamp 1728341909
transform -1 0 10070 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__1824_
timestamp 1728341909
transform 1 0 7370 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__1825_
timestamp 1728341909
transform 1 0 6590 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1826_
timestamp 1728341909
transform 1 0 11010 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1827_
timestamp 1728341909
transform -1 0 7450 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1828_
timestamp 1728341909
transform 1 0 11210 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__1829_
timestamp 1728341909
transform -1 0 7470 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__1830_
timestamp 1728341909
transform 1 0 7610 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__1831_
timestamp 1728341909
transform 1 0 10750 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__1832_
timestamp 1728341909
transform 1 0 10730 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__1833_
timestamp 1728341909
transform 1 0 7290 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1834_
timestamp 1728341909
transform -1 0 7090 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1835_
timestamp 1728341909
transform -1 0 6530 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1836_
timestamp 1728341909
transform -1 0 6090 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1837_
timestamp 1728341909
transform -1 0 5610 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1838_
timestamp 1728341909
transform 1 0 5330 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1839_
timestamp 1728341909
transform 1 0 5910 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1840_
timestamp 1728341909
transform -1 0 8110 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__1841_
timestamp 1728341909
transform -1 0 5050 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__1842_
timestamp 1728341909
transform -1 0 6910 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__1843_
timestamp 1728341909
transform 1 0 7230 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__1844_
timestamp 1728341909
transform -1 0 10310 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__1845_
timestamp 1728341909
transform 1 0 11210 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__1846_
timestamp 1728341909
transform 1 0 11230 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1847_
timestamp 1728341909
transform -1 0 8150 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__1848_
timestamp 1728341909
transform 1 0 10750 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__1849_
timestamp 1728341909
transform -1 0 10670 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__1850_
timestamp 1728341909
transform -1 0 8610 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__1851_
timestamp 1728341909
transform -1 0 11230 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__1852_
timestamp 1728341909
transform 1 0 9790 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__1853_
timestamp 1728341909
transform 1 0 9310 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__1854_
timestamp 1728341909
transform 1 0 9110 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__1855_
timestamp 1728341909
transform 1 0 8870 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__1856_
timestamp 1728341909
transform 1 0 9390 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__1857_
timestamp 1728341909
transform 1 0 9170 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__1858_
timestamp 1728341909
transform 1 0 7350 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__1859_
timestamp 1728341909
transform -1 0 10770 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__1860_
timestamp 1728341909
transform 1 0 7150 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__1861_
timestamp 1728341909
transform 1 0 7390 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__1862_
timestamp 1728341909
transform -1 0 9890 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__1863_
timestamp 1728341909
transform 1 0 8630 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__1864_
timestamp 1728341909
transform 1 0 9930 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__1865_
timestamp 1728341909
transform 1 0 7790 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__1866_
timestamp 1728341909
transform -1 0 8970 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1867_
timestamp 1728341909
transform 1 0 9350 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__1868_
timestamp 1728341909
transform 1 0 10910 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__1869_
timestamp 1728341909
transform 1 0 9370 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__1870_
timestamp 1728341909
transform -1 0 9150 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__1871_
timestamp 1728341909
transform 1 0 8590 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__1872_
timestamp 1728341909
transform 1 0 7870 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__1873_
timestamp 1728341909
transform 1 0 6430 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1874_
timestamp 1728341909
transform -1 0 6890 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1875_
timestamp 1728341909
transform -1 0 6650 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1876_
timestamp 1728341909
transform 1 0 6710 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__1877_
timestamp 1728341909
transform -1 0 8130 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__1878_
timestamp 1728341909
transform -1 0 8390 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__1879_
timestamp 1728341909
transform -1 0 8130 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__1880_
timestamp 1728341909
transform -1 0 7070 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__1881_
timestamp 1728341909
transform -1 0 6390 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__1882_
timestamp 1728341909
transform 1 0 3550 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__1883_
timestamp 1728341909
transform -1 0 7090 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__1884_
timestamp 1728341909
transform -1 0 6610 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__1885_
timestamp 1728341909
transform 1 0 5890 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__1886_
timestamp 1728341909
transform -1 0 6290 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__1887_
timestamp 1728341909
transform 1 0 6910 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__1888_
timestamp 1728341909
transform 1 0 3670 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__1889_
timestamp 1728341909
transform -1 0 6030 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__1890_
timestamp 1728341909
transform 1 0 6490 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__1891_
timestamp 1728341909
transform -1 0 6130 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__1892_
timestamp 1728341909
transform 1 0 5690 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__1893_
timestamp 1728341909
transform 1 0 1090 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__1894_
timestamp 1728341909
transform 1 0 6030 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__1895_
timestamp 1728341909
transform 1 0 6910 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__1896_
timestamp 1728341909
transform 1 0 5230 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__1897_
timestamp 1728341909
transform 1 0 6070 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__1898_
timestamp 1728341909
transform 1 0 6490 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__1899_
timestamp 1728341909
transform 1 0 6590 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__1900_
timestamp 1728341909
transform 1 0 610 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__1901_
timestamp 1728341909
transform 1 0 8050 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__1902_
timestamp 1728341909
transform 1 0 8590 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__1903_
timestamp 1728341909
transform 1 0 7950 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__1904_
timestamp 1728341909
transform -1 0 10110 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1905_
timestamp 1728341909
transform 1 0 7610 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__1906_
timestamp 1728341909
transform 1 0 7590 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__1907_
timestamp 1728341909
transform 1 0 8730 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1908_
timestamp 1728341909
transform -1 0 7790 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1909_
timestamp 1728341909
transform 1 0 1890 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1910_
timestamp 1728341909
transform -1 0 9850 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__1911_
timestamp 1728341909
transform 1 0 9570 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1912_
timestamp 1728341909
transform 1 0 6190 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1913_
timestamp 1728341909
transform 1 0 10710 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__1914_
timestamp 1728341909
transform 1 0 10770 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1915_
timestamp 1728341909
transform -1 0 10330 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1916_
timestamp 1728341909
transform -1 0 5950 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1917_
timestamp 1728341909
transform 1 0 4090 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1918_
timestamp 1728341909
transform -1 0 870 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__1919_
timestamp 1728341909
transform -1 0 150 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__1920_
timestamp 1728341909
transform 1 0 1090 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__1921_
timestamp 1728341909
transform -1 0 1270 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1922_
timestamp 1728341909
transform -1 0 1010 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1923_
timestamp 1728341909
transform 1 0 610 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__1924_
timestamp 1728341909
transform -1 0 4550 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1925_
timestamp 1728341909
transform -1 0 390 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__1926_
timestamp 1728341909
transform 1 0 850 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__1927_
timestamp 1728341909
transform -1 0 2150 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1928_
timestamp 1728341909
transform -1 0 1670 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1929_
timestamp 1728341909
transform 1 0 350 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__1930_
timestamp 1728341909
transform 1 0 730 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1931_
timestamp 1728341909
transform 1 0 610 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__1932_
timestamp 1728341909
transform -1 0 630 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1933_
timestamp 1728341909
transform 1 0 610 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__1934_
timestamp 1728341909
transform -1 0 630 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1935_
timestamp 1728341909
transform -1 0 1610 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1936_
timestamp 1728341909
transform 1 0 870 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1937_
timestamp 1728341909
transform -1 0 630 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__1938_
timestamp 1728341909
transform -1 0 150 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__1939_
timestamp 1728341909
transform 1 0 370 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__1940_
timestamp 1728341909
transform 1 0 890 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1941_
timestamp 1728341909
transform 1 0 610 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__1942_
timestamp 1728341909
transform 1 0 610 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__1943_
timestamp 1728341909
transform 1 0 8170 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__1944_
timestamp 1728341909
transform -1 0 7710 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1945_
timestamp 1728341909
transform -1 0 7490 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1946_
timestamp 1728341909
transform 1 0 8510 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1947_
timestamp 1728341909
transform -1 0 7690 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1948_
timestamp 1728341909
transform -1 0 7030 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1949_
timestamp 1728341909
transform -1 0 7270 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1950_
timestamp 1728341909
transform 1 0 8370 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__1951_
timestamp 1728341909
transform 1 0 8370 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__1952_
timestamp 1728341909
transform 1 0 9890 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1953_
timestamp 1728341909
transform -1 0 8450 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__1954_
timestamp 1728341909
transform 1 0 8290 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1955_
timestamp 1728341909
transform 1 0 6490 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__1956_
timestamp 1728341909
transform -1 0 8050 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1957_
timestamp 1728341909
transform 1 0 8130 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__1958_
timestamp 1728341909
transform 1 0 10490 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__1959_
timestamp 1728341909
transform 1 0 7850 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__1960_
timestamp 1728341909
transform 1 0 7930 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__1961_
timestamp 1728341909
transform 1 0 10750 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__1962_
timestamp 1728341909
transform 1 0 10550 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__1963_
timestamp 1728341909
transform 1 0 9890 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1964_
timestamp 1728341909
transform -1 0 7430 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__1965_
timestamp 1728341909
transform -1 0 7710 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__1966_
timestamp 1728341909
transform -1 0 3570 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__1967_
timestamp 1728341909
transform -1 0 7030 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__1968_
timestamp 1728341909
transform 1 0 7570 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__1969_
timestamp 1728341909
transform -1 0 7830 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__1970_
timestamp 1728341909
transform 1 0 1570 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__1971_
timestamp 1728341909
transform -1 0 870 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1972_
timestamp 1728341909
transform 1 0 1390 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1973_
timestamp 1728341909
transform 1 0 1650 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__1974_
timestamp 1728341909
transform 1 0 8410 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__1975_
timestamp 1728341909
transform 1 0 3030 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__1976_
timestamp 1728341909
transform -1 0 7190 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__1977_
timestamp 1728341909
transform -1 0 2890 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__1978_
timestamp 1728341909
transform -1 0 3870 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__1979_
timestamp 1728341909
transform -1 0 6570 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__1980_
timestamp 1728341909
transform 1 0 7830 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__1981_
timestamp 1728341909
transform 1 0 8350 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__1982_
timestamp 1728341909
transform -1 0 3090 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__1983_
timestamp 1728341909
transform 1 0 1770 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__1984_
timestamp 1728341909
transform 1 0 1850 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__1985_
timestamp 1728341909
transform 1 0 2510 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__1986_
timestamp 1728341909
transform -1 0 7190 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__1987_
timestamp 1728341909
transform 1 0 5130 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__1988_
timestamp 1728341909
transform -1 0 5030 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__1989_
timestamp 1728341909
transform 1 0 6790 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__1990_
timestamp 1728341909
transform -1 0 7310 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__1991_
timestamp 1728341909
transform -1 0 2110 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__1992_
timestamp 1728341909
transform -1 0 1610 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__1993_
timestamp 1728341909
transform -1 0 1890 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__1994_
timestamp 1728341909
transform 1 0 2130 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__1995_
timestamp 1728341909
transform 1 0 8090 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__1996_
timestamp 1728341909
transform -1 0 2310 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__1997_
timestamp 1728341909
transform -1 0 4030 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__1998_
timestamp 1728341909
transform -1 0 6550 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__1999_
timestamp 1728341909
transform -1 0 8270 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2000_
timestamp 1728341909
transform 1 0 1870 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2001_
timestamp 1728341909
transform 1 0 1350 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2002_
timestamp 1728341909
transform 1 0 1590 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2003_
timestamp 1728341909
transform 1 0 1610 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2004_
timestamp 1728341909
transform 1 0 7890 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2005_
timestamp 1728341909
transform 1 0 2050 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2006_
timestamp 1728341909
transform -1 0 6310 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2007_
timestamp 1728341909
transform 1 0 7590 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2008_
timestamp 1728341909
transform -1 0 8110 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2009_
timestamp 1728341909
transform 1 0 850 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2010_
timestamp 1728341909
transform -1 0 910 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2011_
timestamp 1728341909
transform 1 0 610 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2012_
timestamp 1728341909
transform 1 0 870 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2013_
timestamp 1728341909
transform 1 0 5510 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2014_
timestamp 1728341909
transform 1 0 1810 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2015_
timestamp 1728341909
transform -1 0 4010 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2016_
timestamp 1728341909
transform 1 0 6810 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2017_
timestamp 1728341909
transform -1 0 7350 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2018_
timestamp 1728341909
transform -1 0 1590 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2019_
timestamp 1728341909
transform -1 0 1650 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2020_
timestamp 1728341909
transform 1 0 1830 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2021_
timestamp 1728341909
transform 1 0 1790 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2022_
timestamp 1728341909
transform 1 0 4570 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2023_
timestamp 1728341909
transform 1 0 610 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2024_
timestamp 1728341909
transform 1 0 1510 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2025_
timestamp 1728341909
transform 1 0 2570 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2026_
timestamp 1728341909
transform -1 0 4770 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2027_
timestamp 1728341909
transform 1 0 7270 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2028_
timestamp 1728341909
transform -1 0 7550 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2029_
timestamp 1728341909
transform -1 0 150 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2030_
timestamp 1728341909
transform -1 0 630 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2031_
timestamp 1728341909
transform -1 0 390 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2032_
timestamp 1728341909
transform 1 0 610 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2033_
timestamp 1728341909
transform 1 0 7690 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2034_
timestamp 1728341909
transform 1 0 1290 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2035_
timestamp 1728341909
transform 1 0 2170 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2036_
timestamp 1728341909
transform 1 0 2970 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2037_
timestamp 1728341909
transform -1 0 4170 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2038_
timestamp 1728341909
transform 1 0 7610 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2039_
timestamp 1728341909
transform -1 0 7890 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2040_
timestamp 1728341909
transform -1 0 3010 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2041_
timestamp 1728341909
transform -1 0 630 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2042_
timestamp 1728341909
transform 1 0 1790 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__2043_
timestamp 1728341909
transform -1 0 3890 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__2044_
timestamp 1728341909
transform 1 0 5430 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2045_
timestamp 1728341909
transform -1 0 4130 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2046_
timestamp 1728341909
transform 1 0 2930 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__2047_
timestamp 1728341909
transform 1 0 2690 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__2048_
timestamp 1728341909
transform -1 0 3630 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__2049_
timestamp 1728341909
transform -1 0 3030 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__2050_
timestamp 1728341909
transform -1 0 2510 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__2051_
timestamp 1728341909
transform -1 0 2490 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2052_
timestamp 1728341909
transform -1 0 910 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2053_
timestamp 1728341909
transform -1 0 3470 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__2054_
timestamp 1728341909
transform 1 0 3190 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__2055_
timestamp 1728341909
transform -1 0 2830 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__2056_
timestamp 1728341909
transform 1 0 4450 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2057_
timestamp 1728341909
transform -1 0 4010 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2058_
timestamp 1728341909
transform 1 0 4670 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2059_
timestamp 1728341909
transform -1 0 2030 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__2060_
timestamp 1728341909
transform -1 0 3850 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__2061_
timestamp 1728341909
transform 1 0 3590 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__2062_
timestamp 1728341909
transform -1 0 3610 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__2063_
timestamp 1728341909
transform 1 0 2550 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__2064_
timestamp 1728341909
transform -1 0 2650 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2065_
timestamp 1728341909
transform -1 0 2450 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2066_
timestamp 1728341909
transform 1 0 2510 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2067_
timestamp 1728341909
transform -1 0 2830 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__2068_
timestamp 1728341909
transform -1 0 3070 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__2069_
timestamp 1728341909
transform 1 0 2610 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__2070_
timestamp 1728341909
transform -1 0 1150 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2071_
timestamp 1728341909
transform -1 0 2870 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__2072_
timestamp 1728341909
transform -1 0 2610 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__2073_
timestamp 1728341909
transform -1 0 1350 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2074_
timestamp 1728341909
transform 1 0 3290 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__2075_
timestamp 1728341909
transform -1 0 2770 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__2076_
timestamp 1728341909
transform 1 0 2470 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__2077_
timestamp 1728341909
transform -1 0 3330 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__2078_
timestamp 1728341909
transform 1 0 2850 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__2079_
timestamp 1728341909
transform -1 0 3970 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2080_
timestamp 1728341909
transform 1 0 4190 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2081_
timestamp 1728341909
transform -1 0 3750 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2082_
timestamp 1728341909
transform 1 0 5830 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2083_
timestamp 1728341909
transform -1 0 6570 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2084_
timestamp 1728341909
transform 1 0 9990 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2085_
timestamp 1728341909
transform -1 0 10510 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2086_
timestamp 1728341909
transform 1 0 10530 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2087_
timestamp 1728341909
transform 1 0 11070 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__2088_
timestamp 1728341909
transform 1 0 10270 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2089_
timestamp 1728341909
transform -1 0 9570 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2090_
timestamp 1728341909
transform 1 0 10750 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__2091_
timestamp 1728341909
transform 1 0 11250 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__2092_
timestamp 1728341909
transform -1 0 10210 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2093_
timestamp 1728341909
transform 1 0 10270 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__2094_
timestamp 1728341909
transform -1 0 10770 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__2095_
timestamp 1728341909
transform 1 0 10830 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__2096_
timestamp 1728341909
transform -1 0 11230 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__2097_
timestamp 1728341909
transform -1 0 11170 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2098_
timestamp 1728341909
transform 1 0 10250 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2099_
timestamp 1728341909
transform 1 0 10730 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2100_
timestamp 1728341909
transform 1 0 10950 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2101_
timestamp 1728341909
transform 1 0 11190 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2102_
timestamp 1728341909
transform 1 0 4070 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__2103_
timestamp 1728341909
transform 1 0 4310 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__2104_
timestamp 1728341909
transform 1 0 3930 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2105_
timestamp 1728341909
transform -1 0 1830 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2106_
timestamp 1728341909
transform -1 0 2210 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2107_
timestamp 1728341909
transform -1 0 2730 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2108_
timestamp 1728341909
transform 1 0 1530 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2109_
timestamp 1728341909
transform -1 0 2950 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2110_
timestamp 1728341909
transform 1 0 3170 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2111_
timestamp 1728341909
transform 1 0 5370 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2112_
timestamp 1728341909
transform 1 0 11250 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__2113_
timestamp 1728341909
transform -1 0 9830 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__2114_
timestamp 1728341909
transform 1 0 9830 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2115_
timestamp 1728341909
transform -1 0 11150 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2116_
timestamp 1728341909
transform -1 0 11090 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__2117_
timestamp 1728341909
transform -1 0 10690 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__2118_
timestamp 1728341909
transform 1 0 9090 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__2119_
timestamp 1728341909
transform -1 0 11170 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__2120_
timestamp 1728341909
transform 1 0 11110 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2121_
timestamp 1728341909
transform 1 0 11210 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2122_
timestamp 1728341909
transform 1 0 10910 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2123_
timestamp 1728341909
transform 1 0 10970 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2124_
timestamp 1728341909
transform 1 0 9430 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2125_
timestamp 1728341909
transform 1 0 9550 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2126_
timestamp 1728341909
transform -1 0 9990 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2127_
timestamp 1728341909
transform 1 0 9810 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2128_
timestamp 1728341909
transform 1 0 9770 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2129_
timestamp 1728341909
transform -1 0 8990 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2130_
timestamp 1728341909
transform 1 0 9670 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2131_
timestamp 1728341909
transform 1 0 9770 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2132_
timestamp 1728341909
transform 1 0 10230 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2133_
timestamp 1728341909
transform 1 0 10390 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2134_
timestamp 1728341909
transform -1 0 10170 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2135_
timestamp 1728341909
transform 1 0 10670 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2136_
timestamp 1728341909
transform -1 0 10630 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2137_
timestamp 1728341909
transform 1 0 10870 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2138_
timestamp 1728341909
transform -1 0 10970 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2139_
timestamp 1728341909
transform -1 0 10910 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2140_
timestamp 1728341909
transform -1 0 8390 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2141_
timestamp 1728341909
transform 1 0 8630 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2142_
timestamp 1728341909
transform 1 0 1950 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2143_
timestamp 1728341909
transform -1 0 2990 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2144_
timestamp 1728341909
transform -1 0 6090 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2145_
timestamp 1728341909
transform -1 0 6290 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2146_
timestamp 1728341909
transform 1 0 5590 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2147_
timestamp 1728341909
transform -1 0 6830 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2148_
timestamp 1728341909
transform 1 0 9730 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2149_
timestamp 1728341909
transform 1 0 8810 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2150_
timestamp 1728341909
transform -1 0 8570 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2151_
timestamp 1728341909
transform 1 0 8230 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2152_
timestamp 1728341909
transform -1 0 9070 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2153_
timestamp 1728341909
transform -1 0 9170 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2154_
timestamp 1728341909
transform 1 0 8910 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__2155_
timestamp 1728341909
transform 1 0 8070 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__2156_
timestamp 1728341909
transform -1 0 8350 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__2157_
timestamp 1728341909
transform -1 0 8470 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2158_
timestamp 1728341909
transform 1 0 10390 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__2159_
timestamp 1728341909
transform 1 0 6090 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2160_
timestamp 1728341909
transform -1 0 6450 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2161_
timestamp 1728341909
transform 1 0 6650 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2162_
timestamp 1728341909
transform -1 0 7990 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2163_
timestamp 1728341909
transform -1 0 8410 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__2164_
timestamp 1728341909
transform 1 0 7170 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2165_
timestamp 1728341909
transform -1 0 7150 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2166_
timestamp 1728341909
transform -1 0 8210 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2167_
timestamp 1728341909
transform -1 0 7910 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2168_
timestamp 1728341909
transform -1 0 8170 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2169_
timestamp 1728341909
transform 1 0 8210 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2170_
timestamp 1728341909
transform -1 0 8430 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2171_
timestamp 1728341909
transform 1 0 8630 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2172_
timestamp 1728341909
transform -1 0 10490 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2173_
timestamp 1728341909
transform 1 0 10230 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2174_
timestamp 1728341909
transform 1 0 4450 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2175_
timestamp 1728341909
transform -1 0 4010 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2176_
timestamp 1728341909
transform -1 0 5470 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2177_
timestamp 1728341909
transform -1 0 6130 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2178_
timestamp 1728341909
transform -1 0 6390 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2179_
timestamp 1728341909
transform 1 0 6430 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2180_
timestamp 1728341909
transform 1 0 7230 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2181_
timestamp 1728341909
transform 1 0 7370 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__2182_
timestamp 1728341909
transform -1 0 7230 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__2183_
timestamp 1728341909
transform 1 0 6210 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2184_
timestamp 1728341909
transform 1 0 6530 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2185_
timestamp 1728341909
transform -1 0 6670 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2186_
timestamp 1728341909
transform -1 0 9110 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2187_
timestamp 1728341909
transform -1 0 9510 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2188_
timestamp 1728341909
transform 1 0 9110 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2189_
timestamp 1728341909
transform -1 0 8890 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2190_
timestamp 1728341909
transform 1 0 8570 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2191_
timestamp 1728341909
transform 1 0 8810 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2192_
timestamp 1728341909
transform 1 0 7370 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2193_
timestamp 1728341909
transform 1 0 7590 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2194_
timestamp 1728341909
transform -1 0 8710 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__2195_
timestamp 1728341909
transform -1 0 8630 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__2196_
timestamp 1728341909
transform 1 0 8670 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2197_
timestamp 1728341909
transform 1 0 8710 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2198_
timestamp 1728341909
transform -1 0 7310 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2199_
timestamp 1728341909
transform -1 0 7570 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2200_
timestamp 1728341909
transform 1 0 9090 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__2201_
timestamp 1728341909
transform 1 0 8950 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2202_
timestamp 1728341909
transform -1 0 8750 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2203_
timestamp 1728341909
transform 1 0 8470 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2204_
timestamp 1728341909
transform -1 0 8470 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2205_
timestamp 1728341909
transform 1 0 8210 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2206_
timestamp 1728341909
transform -1 0 8090 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2207_
timestamp 1728341909
transform 1 0 8590 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2208_
timestamp 1728341909
transform -1 0 8350 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2209_
timestamp 1728341909
transform -1 0 7870 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2210_
timestamp 1728341909
transform 1 0 2810 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2211_
timestamp 1728341909
transform -1 0 7270 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2212_
timestamp 1728341909
transform -1 0 7530 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2213_
timestamp 1728341909
transform -1 0 8050 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2214_
timestamp 1728341909
transform 1 0 8610 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2215_
timestamp 1728341909
transform 1 0 9310 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2216_
timestamp 1728341909
transform 1 0 9290 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2217_
timestamp 1728341909
transform -1 0 9550 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2218_
timestamp 1728341909
transform 1 0 3990 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2219_
timestamp 1728341909
transform -1 0 2310 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__2220_
timestamp 1728341909
transform -1 0 3730 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2221_
timestamp 1728341909
transform 1 0 4170 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2222_
timestamp 1728341909
transform 1 0 4390 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2223_
timestamp 1728341909
transform 1 0 4210 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2224_
timestamp 1728341909
transform -1 0 2890 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2225_
timestamp 1728341909
transform -1 0 5950 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2226_
timestamp 1728341909
transform 1 0 6070 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2227_
timestamp 1728341909
transform -1 0 7050 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2228_
timestamp 1728341909
transform 1 0 6790 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2229_
timestamp 1728341909
transform 1 0 7850 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__2230_
timestamp 1728341909
transform -1 0 6250 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__2231_
timestamp 1728341909
transform -1 0 6490 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__2232_
timestamp 1728341909
transform 1 0 6910 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2233_
timestamp 1728341909
transform 1 0 7490 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2234_
timestamp 1728341909
transform 1 0 7390 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2235_
timestamp 1728341909
transform 1 0 9470 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2236_
timestamp 1728341909
transform 1 0 10530 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2237_
timestamp 1728341909
transform 1 0 10010 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2238_
timestamp 1728341909
transform -1 0 9930 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2239_
timestamp 1728341909
transform -1 0 5890 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2240_
timestamp 1728341909
transform 1 0 2750 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2241_
timestamp 1728341909
transform -1 0 4430 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2242_
timestamp 1728341909
transform -1 0 4650 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2243_
timestamp 1728341909
transform 1 0 3430 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2244_
timestamp 1728341909
transform 1 0 5190 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2245_
timestamp 1728341909
transform 1 0 7330 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2246_
timestamp 1728341909
transform 1 0 7350 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2247_
timestamp 1728341909
transform -1 0 3310 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2248_
timestamp 1728341909
transform 1 0 3490 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2249_
timestamp 1728341909
transform 1 0 5470 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2250_
timestamp 1728341909
transform 1 0 6730 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2251_
timestamp 1728341909
transform 1 0 7250 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2252_
timestamp 1728341909
transform -1 0 9690 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__2253_
timestamp 1728341909
transform 1 0 9410 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2254_
timestamp 1728341909
transform 1 0 5690 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2255_
timestamp 1728341909
transform -1 0 7030 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2256_
timestamp 1728341909
transform 1 0 7190 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2257_
timestamp 1728341909
transform -1 0 3130 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2258_
timestamp 1728341909
transform -1 0 3090 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__2259_
timestamp 1728341909
transform 1 0 3510 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2260_
timestamp 1728341909
transform 1 0 4690 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2261_
timestamp 1728341909
transform -1 0 5690 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2262_
timestamp 1728341909
transform 1 0 4870 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2263_
timestamp 1728341909
transform 1 0 4930 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2264_
timestamp 1728341909
transform -1 0 6230 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2265_
timestamp 1728341909
transform 1 0 3530 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__2266_
timestamp 1728341909
transform 1 0 7570 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__2267_
timestamp 1728341909
transform -1 0 5470 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__2268_
timestamp 1728341909
transform -1 0 5710 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__2269_
timestamp 1728341909
transform 1 0 5470 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__2270_
timestamp 1728341909
transform -1 0 6310 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__2271_
timestamp 1728341909
transform 1 0 6030 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__2272_
timestamp 1728341909
transform 1 0 5630 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__2273_
timestamp 1728341909
transform 1 0 5450 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__2274_
timestamp 1728341909
transform 1 0 5210 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__2275_
timestamp 1728341909
transform 1 0 5690 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__2276_
timestamp 1728341909
transform -1 0 6330 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2277_
timestamp 1728341909
transform 1 0 7830 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__2278_
timestamp 1728341909
transform -1 0 7770 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2279_
timestamp 1728341909
transform 1 0 6530 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2280_
timestamp 1728341909
transform -1 0 6550 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2281_
timestamp 1728341909
transform -1 0 6310 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2282_
timestamp 1728341909
transform 1 0 6590 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2283_
timestamp 1728341909
transform 1 0 7290 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2284_
timestamp 1728341909
transform 1 0 9250 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2285_
timestamp 1728341909
transform 1 0 9690 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2286_
timestamp 1728341909
transform -1 0 2590 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__2287_
timestamp 1728341909
transform -1 0 1850 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2288_
timestamp 1728341909
transform -1 0 2290 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2289_
timestamp 1728341909
transform 1 0 2250 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2290_
timestamp 1728341909
transform -1 0 1810 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2291_
timestamp 1728341909
transform 1 0 2030 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2292_
timestamp 1728341909
transform 1 0 4150 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2293_
timestamp 1728341909
transform 1 0 4890 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2294_
timestamp 1728341909
transform 1 0 6110 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2295_
timestamp 1728341909
transform -1 0 2290 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2296_
timestamp 1728341909
transform 1 0 3730 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2297_
timestamp 1728341909
transform 1 0 2270 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2298_
timestamp 1728341909
transform 1 0 2030 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2299_
timestamp 1728341909
transform 1 0 3490 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2300_
timestamp 1728341909
transform 1 0 3230 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2301_
timestamp 1728341909
transform -1 0 3690 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2302_
timestamp 1728341909
transform 1 0 5170 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2303_
timestamp 1728341909
transform -1 0 5150 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2304_
timestamp 1728341909
transform 1 0 5390 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2305_
timestamp 1728341909
transform -1 0 1590 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2306_
timestamp 1728341909
transform 1 0 2490 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2307_
timestamp 1728341909
transform -1 0 5650 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2308_
timestamp 1728341909
transform -1 0 5650 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2309_
timestamp 1728341909
transform 1 0 4650 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2310_
timestamp 1728341909
transform 1 0 4410 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2311_
timestamp 1728341909
transform -1 0 3810 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2312_
timestamp 1728341909
transform -1 0 4050 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2313_
timestamp 1728341909
transform 1 0 5330 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2314_
timestamp 1728341909
transform 1 0 4510 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2315_
timestamp 1728341909
transform 1 0 5470 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2316_
timestamp 1728341909
transform -1 0 9910 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2317_
timestamp 1728341909
transform 1 0 11210 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2318_
timestamp 1728341909
transform -1 0 10910 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__2319_
timestamp 1728341909
transform -1 0 10530 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__2320_
timestamp 1728341909
transform 1 0 10690 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2321_
timestamp 1728341909
transform 1 0 10630 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__2322_
timestamp 1728341909
transform 1 0 10530 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__2323_
timestamp 1728341909
transform 1 0 6790 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2324_
timestamp 1728341909
transform 1 0 6990 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2325_
timestamp 1728341909
transform 1 0 9350 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2326_
timestamp 1728341909
transform -1 0 8890 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2327_
timestamp 1728341909
transform -1 0 9350 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2328_
timestamp 1728341909
transform -1 0 9590 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2329_
timestamp 1728341909
transform 1 0 9310 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2330_
timestamp 1728341909
transform -1 0 9070 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2331_
timestamp 1728341909
transform -1 0 9230 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2332_
timestamp 1728341909
transform 1 0 9210 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2333_
timestamp 1728341909
transform 1 0 9470 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2334_
timestamp 1728341909
transform -1 0 9670 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2335_
timestamp 1728341909
transform 1 0 5710 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2336_
timestamp 1728341909
transform 1 0 6230 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2337_
timestamp 1728341909
transform -1 0 6010 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2338_
timestamp 1728341909
transform -1 0 5950 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2339_
timestamp 1728341909
transform 1 0 10430 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2340_
timestamp 1728341909
transform -1 0 9310 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2341_
timestamp 1728341909
transform 1 0 9310 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2342_
timestamp 1728341909
transform 1 0 10170 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2343_
timestamp 1728341909
transform -1 0 9670 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2344_
timestamp 1728341909
transform 1 0 9770 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2345_
timestamp 1728341909
transform -1 0 6950 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2346_
timestamp 1728341909
transform 1 0 6810 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2347_
timestamp 1728341909
transform -1 0 7150 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2348_
timestamp 1728341909
transform 1 0 8150 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2349_
timestamp 1728341909
transform -1 0 7850 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2350_
timestamp 1728341909
transform 1 0 7570 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2351_
timestamp 1728341909
transform -1 0 5270 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2352_
timestamp 1728341909
transform 1 0 5870 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2353_
timestamp 1728341909
transform -1 0 4290 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2354_
timestamp 1728341909
transform 1 0 4770 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2355_
timestamp 1728341909
transform -1 0 5030 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2356_
timestamp 1728341909
transform 1 0 5970 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2357_
timestamp 1728341909
transform -1 0 5730 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2358_
timestamp 1728341909
transform 1 0 7010 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2359_
timestamp 1728341909
transform 1 0 6370 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2360_
timestamp 1728341909
transform 1 0 6610 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2361_
timestamp 1728341909
transform 1 0 7910 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__2362_
timestamp 1728341909
transform 1 0 7430 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2363_
timestamp 1728341909
transform -1 0 7530 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2364_
timestamp 1728341909
transform 1 0 8150 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__2365_
timestamp 1728341909
transform -1 0 8030 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2366_
timestamp 1728341909
transform 1 0 7790 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2367_
timestamp 1728341909
transform 1 0 8070 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2368_
timestamp 1728341909
transform 1 0 8290 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2369_
timestamp 1728341909
transform -1 0 10010 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2370_
timestamp 1728341909
transform 1 0 5430 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2371_
timestamp 1728341909
transform -1 0 8830 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2372_
timestamp 1728341909
transform -1 0 8570 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2373_
timestamp 1728341909
transform -1 0 8150 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2374_
timestamp 1728341909
transform 1 0 8150 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2375_
timestamp 1728341909
transform 1 0 6550 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2376_
timestamp 1728341909
transform 1 0 8510 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2377_
timestamp 1728341909
transform -1 0 8770 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2378_
timestamp 1728341909
transform -1 0 9070 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2379_
timestamp 1728341909
transform -1 0 6930 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2380_
timestamp 1728341909
transform -1 0 7070 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2381_
timestamp 1728341909
transform -1 0 6930 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2382_
timestamp 1728341909
transform -1 0 8010 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2383_
timestamp 1728341909
transform 1 0 7730 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2384_
timestamp 1728341909
transform 1 0 7830 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2385_
timestamp 1728341909
transform -1 0 7570 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2386_
timestamp 1728341909
transform -1 0 6690 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2387_
timestamp 1728341909
transform -1 0 6450 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2388_
timestamp 1728341909
transform -1 0 9010 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2389_
timestamp 1728341909
transform -1 0 8390 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2390_
timestamp 1728341909
transform -1 0 8330 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2391_
timestamp 1728341909
transform -1 0 9570 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2392_
timestamp 1728341909
transform 1 0 8330 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2393_
timestamp 1728341909
transform 1 0 8290 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2394_
timestamp 1728341909
transform 1 0 8930 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2395_
timestamp 1728341909
transform 1 0 8890 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2396_
timestamp 1728341909
transform 1 0 9170 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2397_
timestamp 1728341909
transform -1 0 9430 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2398_
timestamp 1728341909
transform 1 0 8810 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2399_
timestamp 1728341909
transform -1 0 7690 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2400_
timestamp 1728341909
transform 1 0 7430 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2401_
timestamp 1728341909
transform 1 0 8550 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2402_
timestamp 1728341909
transform -1 0 6490 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2403_
timestamp 1728341909
transform -1 0 6690 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2404_
timestamp 1728341909
transform -1 0 7650 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2405_
timestamp 1728341909
transform -1 0 7430 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2406_
timestamp 1728341909
transform 1 0 7150 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2407_
timestamp 1728341909
transform -1 0 6690 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2408_
timestamp 1728341909
transform -1 0 5990 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2409_
timestamp 1728341909
transform 1 0 7070 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2410_
timestamp 1728341909
transform -1 0 7350 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2411_
timestamp 1728341909
transform -1 0 6910 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2412_
timestamp 1728341909
transform -1 0 7570 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2413_
timestamp 1728341909
transform 1 0 7090 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2414_
timestamp 1728341909
transform 1 0 6910 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2415_
timestamp 1728341909
transform -1 0 8110 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2416_
timestamp 1728341909
transform 1 0 7850 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2417_
timestamp 1728341909
transform -1 0 9090 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2418_
timestamp 1728341909
transform -1 0 8870 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2419_
timestamp 1728341909
transform 1 0 7130 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2420_
timestamp 1728341909
transform 1 0 2290 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2421_
timestamp 1728341909
transform -1 0 9750 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2422_
timestamp 1728341909
transform 1 0 8330 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__2423_
timestamp 1728341909
transform 1 0 9050 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2424_
timestamp 1728341909
transform 1 0 8830 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2425_
timestamp 1728341909
transform 1 0 3230 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2426_
timestamp 1728341909
transform 1 0 8810 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2427_
timestamp 1728341909
transform 1 0 8890 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__2428_
timestamp 1728341909
transform 1 0 9290 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2429_
timestamp 1728341909
transform 1 0 9510 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2430_
timestamp 1728341909
transform 1 0 8870 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2431_
timestamp 1728341909
transform -1 0 9330 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2432_
timestamp 1728341909
transform 1 0 9550 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2433_
timestamp 1728341909
transform -1 0 9970 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2434_
timestamp 1728341909
transform -1 0 10050 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2435_
timestamp 1728341909
transform 1 0 4510 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__2436_
timestamp 1728341909
transform 1 0 9270 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2437_
timestamp 1728341909
transform 1 0 10950 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__2438_
timestamp 1728341909
transform -1 0 11010 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__2439_
timestamp 1728341909
transform -1 0 10990 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__2440_
timestamp 1728341909
transform 1 0 9110 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__2441_
timestamp 1728341909
transform -1 0 6250 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__2442_
timestamp 1728341909
transform -1 0 8330 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2443_
timestamp 1728341909
transform 1 0 3890 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2444_
timestamp 1728341909
transform -1 0 4770 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__2445_
timestamp 1728341909
transform -1 0 8670 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__2446_
timestamp 1728341909
transform 1 0 8310 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2447_
timestamp 1728341909
transform 1 0 8150 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2448_
timestamp 1728341909
transform 1 0 8550 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2449_
timestamp 1728341909
transform -1 0 8830 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2450_
timestamp 1728341909
transform -1 0 9030 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2451_
timestamp 1728341909
transform 1 0 3890 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2452_
timestamp 1728341909
transform 1 0 7670 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2453_
timestamp 1728341909
transform -1 0 6690 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2454_
timestamp 1728341909
transform -1 0 6410 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2455_
timestamp 1728341909
transform -1 0 6690 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2456_
timestamp 1728341909
transform -1 0 8810 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2457_
timestamp 1728341909
transform -1 0 9030 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2458_
timestamp 1728341909
transform -1 0 6870 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2459_
timestamp 1728341909
transform -1 0 3650 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2460_
timestamp 1728341909
transform 1 0 7170 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2461_
timestamp 1728341909
transform 1 0 7090 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2462_
timestamp 1728341909
transform -1 0 7370 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2463_
timestamp 1728341909
transform -1 0 7390 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2464_
timestamp 1728341909
transform 1 0 4550 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__2465_
timestamp 1728341909
transform -1 0 7450 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2466_
timestamp 1728341909
transform -1 0 3430 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2467_
timestamp 1728341909
transform 1 0 6250 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2468_
timestamp 1728341909
transform -1 0 6370 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2469_
timestamp 1728341909
transform -1 0 6210 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2470_
timestamp 1728341909
transform -1 0 6470 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2471_
timestamp 1728341909
transform -1 0 8130 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2472_
timestamp 1728341909
transform -1 0 6150 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2473_
timestamp 1728341909
transform -1 0 5490 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2474_
timestamp 1728341909
transform -1 0 5410 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2475_
timestamp 1728341909
transform -1 0 7870 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__2476_
timestamp 1728341909
transform -1 0 2790 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2477_
timestamp 1728341909
transform -1 0 5270 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2478_
timestamp 1728341909
transform 1 0 5350 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2479_
timestamp 1728341909
transform -1 0 8090 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2480_
timestamp 1728341909
transform 1 0 5990 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2481_
timestamp 1728341909
transform 1 0 4250 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2482_
timestamp 1728341909
transform -1 0 2530 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2483_
timestamp 1728341909
transform -1 0 4770 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2484_
timestamp 1728341909
transform -1 0 5810 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2485_
timestamp 1728341909
transform -1 0 7050 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2486_
timestamp 1728341909
transform 1 0 3170 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2487_
timestamp 1728341909
transform -1 0 5750 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2488_
timestamp 1728341909
transform 1 0 6510 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2489_
timestamp 1728341909
transform -1 0 6790 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2490_
timestamp 1728341909
transform 1 0 7770 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2491_
timestamp 1728341909
transform -1 0 8010 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2492_
timestamp 1728341909
transform -1 0 2950 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2493_
timestamp 1728341909
transform -1 0 5590 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2494_
timestamp 1728341909
transform -1 0 6670 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2495_
timestamp 1728341909
transform 1 0 6910 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2496_
timestamp 1728341909
transform 1 0 7630 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2497_
timestamp 1728341909
transform -1 0 7870 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2498_
timestamp 1728341909
transform -1 0 8850 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__2499_
timestamp 1728341909
transform 1 0 9090 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2500_
timestamp 1728341909
transform -1 0 7710 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2501_
timestamp 1728341909
transform -1 0 6830 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__2502_
timestamp 1728341909
transform -1 0 7690 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__2503_
timestamp 1728341909
transform 1 0 11190 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2504_
timestamp 1728341909
transform -1 0 4630 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2505_
timestamp 1728341909
transform -1 0 5770 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2506_
timestamp 1728341909
transform -1 0 6790 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__2507_
timestamp 1728341909
transform 1 0 5930 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2508_
timestamp 1728341909
transform 1 0 5730 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2509_
timestamp 1728341909
transform -1 0 8890 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__2510_
timestamp 1728341909
transform -1 0 8150 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__2511_
timestamp 1728341909
transform -1 0 7470 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__2512_
timestamp 1728341909
transform 1 0 7170 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__2513_
timestamp 1728341909
transform 1 0 6950 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__2514_
timestamp 1728341909
transform 1 0 7110 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__2515_
timestamp 1728341909
transform 1 0 10450 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__2516_
timestamp 1728341909
transform 1 0 8590 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2517_
timestamp 1728341909
transform 1 0 10690 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2518_
timestamp 1728341909
transform -1 0 9790 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__2519_
timestamp 1728341909
transform 1 0 10030 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__2520_
timestamp 1728341909
transform -1 0 10490 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2521_
timestamp 1728341909
transform -1 0 8590 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2522_
timestamp 1728341909
transform 1 0 6150 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2523_
timestamp 1728341909
transform 1 0 5970 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2524_
timestamp 1728341909
transform 1 0 8350 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2525_
timestamp 1728341909
transform 1 0 6850 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2526_
timestamp 1728341909
transform -1 0 7850 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2527_
timestamp 1728341909
transform 1 0 8070 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2528_
timestamp 1728341909
transform -1 0 8130 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2529_
timestamp 1728341909
transform 1 0 7910 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2530_
timestamp 1728341909
transform -1 0 7870 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2531_
timestamp 1728341909
transform -1 0 7890 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2532_
timestamp 1728341909
transform 1 0 7890 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2533_
timestamp 1728341909
transform -1 0 5550 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2534_
timestamp 1728341909
transform -1 0 5970 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2535_
timestamp 1728341909
transform -1 0 7650 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2536_
timestamp 1728341909
transform 1 0 7450 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2537_
timestamp 1728341909
transform 1 0 7370 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2538_
timestamp 1728341909
transform 1 0 8090 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2539_
timestamp 1728341909
transform 1 0 5950 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2540_
timestamp 1728341909
transform 1 0 5670 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2541_
timestamp 1728341909
transform 1 0 6190 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2542_
timestamp 1728341909
transform -1 0 6730 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2543_
timestamp 1728341909
transform -1 0 6690 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2544_
timestamp 1728341909
transform 1 0 6230 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2545_
timestamp 1728341909
transform 1 0 6930 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2546_
timestamp 1728341909
transform 1 0 6190 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2547_
timestamp 1728341909
transform 1 0 6410 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2548_
timestamp 1728341909
transform 1 0 7190 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2549_
timestamp 1728341909
transform 1 0 7450 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2550_
timestamp 1728341909
transform -1 0 7610 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2551_
timestamp 1728341909
transform -1 0 6330 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2552_
timestamp 1728341909
transform -1 0 4890 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2553_
timestamp 1728341909
transform -1 0 5930 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2554_
timestamp 1728341909
transform -1 0 5650 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2555_
timestamp 1728341909
transform 1 0 5710 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2556_
timestamp 1728341909
transform 1 0 5090 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2557_
timestamp 1728341909
transform 1 0 5830 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2558_
timestamp 1728341909
transform -1 0 6470 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2559_
timestamp 1728341909
transform 1 0 6150 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__2560_
timestamp 1728341909
transform 1 0 4410 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2561_
timestamp 1728341909
transform -1 0 5470 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2562_
timestamp 1728341909
transform 1 0 5090 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2563_
timestamp 1728341909
transform -1 0 4990 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2564_
timestamp 1728341909
transform -1 0 4650 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2565_
timestamp 1728341909
transform 1 0 4790 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2566_
timestamp 1728341909
transform -1 0 5010 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2567_
timestamp 1728341909
transform 1 0 5210 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2568_
timestamp 1728341909
transform 1 0 5350 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__2569_
timestamp 1728341909
transform -1 0 4230 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2570_
timestamp 1728341909
transform 1 0 5250 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2571_
timestamp 1728341909
transform 1 0 4370 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2572_
timestamp 1728341909
transform -1 0 4490 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2573_
timestamp 1728341909
transform 1 0 4730 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2574_
timestamp 1728341909
transform 1 0 5450 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2575_
timestamp 1728341909
transform -1 0 5010 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2576_
timestamp 1728341909
transform 1 0 5190 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2577_
timestamp 1728341909
transform 1 0 4930 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2578_
timestamp 1728341909
transform -1 0 4870 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2579_
timestamp 1728341909
transform 1 0 4730 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__2580_
timestamp 1728341909
transform 1 0 4770 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__2581_
timestamp 1728341909
transform -1 0 4210 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2582_
timestamp 1728341909
transform -1 0 3350 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2583_
timestamp 1728341909
transform 1 0 2290 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2584_
timestamp 1728341909
transform 1 0 3250 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2585_
timestamp 1728341909
transform -1 0 6410 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2586_
timestamp 1728341909
transform -1 0 3770 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2587_
timestamp 1728341909
transform -1 0 3510 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2588_
timestamp 1728341909
transform -1 0 3030 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2589_
timestamp 1728341909
transform -1 0 3030 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2590_
timestamp 1728341909
transform 1 0 3650 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__2591_
timestamp 1728341909
transform -1 0 3130 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2592_
timestamp 1728341909
transform 1 0 2630 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2593_
timestamp 1728341909
transform -1 0 2730 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2594_
timestamp 1728341909
transform -1 0 2750 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2595_
timestamp 1728341909
transform -1 0 3830 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__2596_
timestamp 1728341909
transform 1 0 3430 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2597_
timestamp 1728341909
transform 1 0 3370 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2598_
timestamp 1728341909
transform -1 0 3250 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2599_
timestamp 1728341909
transform -1 0 3250 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2600_
timestamp 1728341909
transform 1 0 2970 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2601_
timestamp 1728341909
transform -1 0 2530 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2602_
timestamp 1728341909
transform -1 0 2790 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2603_
timestamp 1728341909
transform -1 0 2390 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2604_
timestamp 1728341909
transform 1 0 2530 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2605_
timestamp 1728341909
transform -1 0 2530 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2606_
timestamp 1728341909
transform 1 0 2250 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2607_
timestamp 1728341909
transform -1 0 1610 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2608_
timestamp 1728341909
transform -1 0 1130 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2609_
timestamp 1728341909
transform 1 0 2090 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2610_
timestamp 1728341909
transform 1 0 1330 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2611_
timestamp 1728341909
transform -1 0 1310 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2612_
timestamp 1728341909
transform -1 0 1050 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2613_
timestamp 1728341909
transform -1 0 2030 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2614_
timestamp 1728341909
transform -1 0 650 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2615_
timestamp 1728341909
transform 1 0 1830 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2616_
timestamp 1728341909
transform 1 0 1570 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2617_
timestamp 1728341909
transform -1 0 1570 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2618_
timestamp 1728341909
transform -1 0 1810 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2619_
timestamp 1728341909
transform 1 0 850 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2620_
timestamp 1728341909
transform -1 0 1370 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2621_
timestamp 1728341909
transform 1 0 1110 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2622_
timestamp 1728341909
transform -1 0 1330 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2623_
timestamp 1728341909
transform 1 0 1070 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2624_
timestamp 1728341909
transform -1 0 610 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2625_
timestamp 1728341909
transform -1 0 2690 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2626_
timestamp 1728341909
transform 1 0 1710 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2627_
timestamp 1728341909
transform 1 0 1450 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2628_
timestamp 1728341909
transform 1 0 850 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2629_
timestamp 1728341909
transform -1 0 3450 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__2630_
timestamp 1728341909
transform 1 0 4310 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__2631_
timestamp 1728341909
transform -1 0 4970 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__2632_
timestamp 1728341909
transform 1 0 10950 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2633_
timestamp 1728341909
transform 1 0 3950 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2634_
timestamp 1728341909
transform 1 0 9050 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2635_
timestamp 1728341909
transform -1 0 2330 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__2636_
timestamp 1728341909
transform -1 0 9210 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__2637_
timestamp 1728341909
transform 1 0 4410 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2638_
timestamp 1728341909
transform 1 0 4910 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2639_
timestamp 1728341909
transform -1 0 9990 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__2640_
timestamp 1728341909
transform -1 0 9930 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__2641_
timestamp 1728341909
transform 1 0 10230 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2642_
timestamp 1728341909
transform -1 0 9570 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__2643_
timestamp 1728341909
transform 1 0 10970 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2644_
timestamp 1728341909
transform -1 0 9810 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2645_
timestamp 1728341909
transform -1 0 9770 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__2646_
timestamp 1728341909
transform 1 0 10170 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__2647_
timestamp 1728341909
transform -1 0 8650 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2648_
timestamp 1728341909
transform -1 0 4230 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__2649_
timestamp 1728341909
transform -1 0 5870 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2650_
timestamp 1728341909
transform 1 0 9370 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__2651_
timestamp 1728341909
transform -1 0 5750 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2652_
timestamp 1728341909
transform -1 0 7910 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__2653_
timestamp 1728341909
transform -1 0 7810 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__2654_
timestamp 1728341909
transform 1 0 4730 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2655_
timestamp 1728341909
transform -1 0 5510 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2656_
timestamp 1728341909
transform -1 0 6090 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2657_
timestamp 1728341909
transform -1 0 6830 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2658_
timestamp 1728341909
transform 1 0 6330 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2659_
timestamp 1728341909
transform 1 0 7030 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2660_
timestamp 1728341909
transform -1 0 7310 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2661_
timestamp 1728341909
transform -1 0 4530 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2662_
timestamp 1728341909
transform 1 0 4490 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2663_
timestamp 1728341909
transform 1 0 6410 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2664_
timestamp 1728341909
transform -1 0 6670 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2665_
timestamp 1728341909
transform 1 0 7170 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2666_
timestamp 1728341909
transform 1 0 6910 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2667_
timestamp 1728341909
transform 1 0 7650 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2668_
timestamp 1728341909
transform 1 0 7390 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2669_
timestamp 1728341909
transform 1 0 8050 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2670_
timestamp 1728341909
transform -1 0 4270 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2671_
timestamp 1728341909
transform -1 0 5390 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__2672_
timestamp 1728341909
transform 1 0 5290 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2673_
timestamp 1728341909
transform 1 0 7250 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2674_
timestamp 1728341909
transform -1 0 7470 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2675_
timestamp 1728341909
transform 1 0 7710 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2676_
timestamp 1728341909
transform -1 0 7650 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2677_
timestamp 1728341909
transform 1 0 7830 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2678_
timestamp 1728341909
transform 1 0 7790 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2679_
timestamp 1728341909
transform 1 0 4230 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2680_
timestamp 1728341909
transform -1 0 4490 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2681_
timestamp 1728341909
transform 1 0 6190 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2682_
timestamp 1728341909
transform 1 0 6810 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2683_
timestamp 1728341909
transform 1 0 4150 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2684_
timestamp 1728341909
transform -1 0 5810 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2685_
timestamp 1728341909
transform 1 0 5530 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2686_
timestamp 1728341909
transform -1 0 6950 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2687_
timestamp 1728341909
transform 1 0 7410 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2688_
timestamp 1728341909
transform -1 0 7550 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2689_
timestamp 1728341909
transform 1 0 6570 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2690_
timestamp 1728341909
transform 1 0 6650 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2691_
timestamp 1728341909
transform 1 0 7150 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2692_
timestamp 1728341909
transform -1 0 7290 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2693_
timestamp 1728341909
transform 1 0 5130 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2694_
timestamp 1728341909
transform -1 0 5270 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2695_
timestamp 1728341909
transform 1 0 6710 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2696_
timestamp 1728341909
transform 1 0 6650 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2697_
timestamp 1728341909
transform 1 0 7070 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2698_
timestamp 1728341909
transform 1 0 6970 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2699_
timestamp 1728341909
transform -1 0 6410 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2700_
timestamp 1728341909
transform 1 0 5470 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2701_
timestamp 1728341909
transform -1 0 5550 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2702_
timestamp 1728341909
transform -1 0 5630 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2703_
timestamp 1728341909
transform -1 0 5650 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2704_
timestamp 1728341909
transform 1 0 5710 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2705_
timestamp 1728341909
transform 1 0 5970 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2706_
timestamp 1728341909
transform -1 0 6230 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2707_
timestamp 1728341909
transform -1 0 5970 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2708_
timestamp 1728341909
transform -1 0 2370 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2709_
timestamp 1728341909
transform -1 0 5030 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2710_
timestamp 1728341909
transform -1 0 4950 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2711_
timestamp 1728341909
transform -1 0 5150 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2712_
timestamp 1728341909
transform -1 0 5730 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2713_
timestamp 1728341909
transform -1 0 5870 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2714_
timestamp 1728341909
transform -1 0 6170 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2715_
timestamp 1728341909
transform 1 0 5890 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2716_
timestamp 1728341909
transform -1 0 6730 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2717_
timestamp 1728341909
transform 1 0 6670 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2718_
timestamp 1728341909
transform 1 0 6250 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2719_
timestamp 1728341909
transform -1 0 6410 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2720_
timestamp 1728341909
transform 1 0 4710 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2721_
timestamp 1728341909
transform 1 0 4990 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2722_
timestamp 1728341909
transform 1 0 5230 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2723_
timestamp 1728341909
transform -1 0 5490 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2724_
timestamp 1728341909
transform 1 0 6210 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2725_
timestamp 1728341909
transform 1 0 6450 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2726_
timestamp 1728341909
transform -1 0 6210 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__2727_
timestamp 1728341909
transform 1 0 5910 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__2728_
timestamp 1728341909
transform -1 0 4390 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2729_
timestamp 1728341909
transform -1 0 4250 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2730_
timestamp 1728341909
transform -1 0 5290 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2731_
timestamp 1728341909
transform -1 0 5410 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2732_
timestamp 1728341909
transform -1 0 5710 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2733_
timestamp 1728341909
transform -1 0 5970 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2734_
timestamp 1728341909
transform -1 0 5290 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2735_
timestamp 1728341909
transform 1 0 5490 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2736_
timestamp 1728341909
transform -1 0 8410 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__2737_
timestamp 1728341909
transform 1 0 3810 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2738_
timestamp 1728341909
transform 1 0 3990 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2739_
timestamp 1728341909
transform -1 0 3810 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2740_
timestamp 1728341909
transform -1 0 3750 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2741_
timestamp 1728341909
transform -1 0 4090 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2742_
timestamp 1728341909
transform -1 0 4230 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2743_
timestamp 1728341909
transform 1 0 4970 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2744_
timestamp 1728341909
transform 1 0 4710 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__2745_
timestamp 1728341909
transform 1 0 5190 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2746_
timestamp 1728341909
transform 1 0 4690 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2747_
timestamp 1728341909
transform 1 0 5610 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2748_
timestamp 1728341909
transform -1 0 5010 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2749_
timestamp 1728341909
transform -1 0 5370 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2750_
timestamp 1728341909
transform -1 0 5470 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2751_
timestamp 1728341909
transform 1 0 4450 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2752_
timestamp 1728341909
transform 1 0 3950 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2753_
timestamp 1728341909
transform -1 0 3490 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2754_
timestamp 1728341909
transform -1 0 3070 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2755_
timestamp 1728341909
transform 1 0 3330 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2756_
timestamp 1728341909
transform -1 0 3710 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2757_
timestamp 1728341909
transform -1 0 3730 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2758_
timestamp 1728341909
transform -1 0 3710 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2759_
timestamp 1728341909
transform -1 0 3590 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2760_
timestamp 1728341909
transform -1 0 3630 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2761_
timestamp 1728341909
transform -1 0 3770 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2762_
timestamp 1728341909
transform -1 0 3530 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2763_
timestamp 1728341909
transform 1 0 3090 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__2764_
timestamp 1728341909
transform 1 0 3370 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__2765_
timestamp 1728341909
transform -1 0 2690 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2766_
timestamp 1728341909
transform 1 0 3770 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__2767_
timestamp 1728341909
transform -1 0 4470 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2768_
timestamp 1728341909
transform 1 0 4550 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2769_
timestamp 1728341909
transform 1 0 5210 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2770_
timestamp 1728341909
transform -1 0 4710 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2771_
timestamp 1728341909
transform -1 0 4990 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2772_
timestamp 1728341909
transform -1 0 4970 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2773_
timestamp 1728341909
transform 1 0 2730 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2774_
timestamp 1728341909
transform -1 0 2590 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__2775_
timestamp 1728341909
transform 1 0 3950 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2776_
timestamp 1728341909
transform 1 0 4470 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2777_
timestamp 1728341909
transform 1 0 5210 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2778_
timestamp 1728341909
transform -1 0 4710 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2779_
timestamp 1728341909
transform 1 0 4030 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__2780_
timestamp 1728341909
transform 1 0 2810 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__2781_
timestamp 1728341909
transform -1 0 4030 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2782_
timestamp 1728341909
transform -1 0 2830 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2783_
timestamp 1728341909
transform 1 0 2530 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2784_
timestamp 1728341909
transform 1 0 610 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2785_
timestamp 1728341909
transform -1 0 2310 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2786_
timestamp 1728341909
transform 1 0 2570 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2787_
timestamp 1728341909
transform -1 0 2990 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2788_
timestamp 1728341909
transform -1 0 2490 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2789_
timestamp 1728341909
transform -1 0 3790 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2790_
timestamp 1728341909
transform 1 0 3270 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2791_
timestamp 1728341909
transform -1 0 3010 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2792_
timestamp 1728341909
transform -1 0 2910 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2793_
timestamp 1728341909
transform -1 0 2330 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__2794_
timestamp 1728341909
transform 1 0 2210 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2795_
timestamp 1728341909
transform 1 0 850 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2796_
timestamp 1728341909
transform 1 0 1790 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2797_
timestamp 1728341909
transform -1 0 2070 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2798_
timestamp 1728341909
transform 1 0 1290 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2799_
timestamp 1728341909
transform -1 0 1570 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2800_
timestamp 1728341909
transform -1 0 1830 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2801_
timestamp 1728341909
transform 1 0 1790 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2802_
timestamp 1728341909
transform 1 0 1870 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2803_
timestamp 1728341909
transform 1 0 3350 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2804_
timestamp 1728341909
transform -1 0 510 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__2805_
timestamp 1728341909
transform 1 0 7050 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2806_
timestamp 1728341909
transform -1 0 5470 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2807_
timestamp 1728341909
transform -1 0 5070 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2808_
timestamp 1728341909
transform 1 0 3990 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2809_
timestamp 1728341909
transform -1 0 4450 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2810_
timestamp 1728341909
transform -1 0 4810 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2811_
timestamp 1728341909
transform -1 0 4670 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2812_
timestamp 1728341909
transform 1 0 4290 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2813_
timestamp 1728341909
transform 1 0 4050 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__2814_
timestamp 1728341909
transform 1 0 4170 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__2815_
timestamp 1728341909
transform -1 0 4250 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2816_
timestamp 1728341909
transform 1 0 2550 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2817_
timestamp 1728341909
transform -1 0 2830 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__2818_
timestamp 1728341909
transform 1 0 2790 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2819_
timestamp 1728341909
transform 1 0 3230 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2820_
timestamp 1728341909
transform 1 0 3470 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2821_
timestamp 1728341909
transform -1 0 4010 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2822_
timestamp 1728341909
transform -1 0 4810 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2823_
timestamp 1728341909
transform -1 0 1790 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2824_
timestamp 1728341909
transform 1 0 610 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__2825_
timestamp 1728341909
transform 1 0 590 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2826_
timestamp 1728341909
transform -1 0 750 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__2827_
timestamp 1728341909
transform 1 0 1790 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2828_
timestamp 1728341909
transform -1 0 2070 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2829_
timestamp 1728341909
transform 1 0 1310 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2830_
timestamp 1728341909
transform -1 0 1570 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2831_
timestamp 1728341909
transform -1 0 1590 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__2832_
timestamp 1728341909
transform 1 0 2090 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2833_
timestamp 1728341909
transform -1 0 1110 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__2834_
timestamp 1728341909
transform 1 0 930 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__2835_
timestamp 1728341909
transform 1 0 1170 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__2836_
timestamp 1728341909
transform 1 0 1390 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__2837_
timestamp 1728341909
transform 1 0 1710 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__2838_
timestamp 1728341909
transform -1 0 1590 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__2839_
timestamp 1728341909
transform 1 0 870 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__2840_
timestamp 1728341909
transform 1 0 1310 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2841_
timestamp 1728341909
transform 1 0 2110 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2842_
timestamp 1728341909
transform -1 0 1770 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2843_
timestamp 1728341909
transform -1 0 1870 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2844_
timestamp 1728341909
transform -1 0 1630 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__2845_
timestamp 1728341909
transform -1 0 1570 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2846_
timestamp 1728341909
transform 1 0 1350 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2847_
timestamp 1728341909
transform -1 0 1350 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__2848_
timestamp 1728341909
transform -1 0 1330 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2849_
timestamp 1728341909
transform -1 0 1630 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2850_
timestamp 1728341909
transform -1 0 1550 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2851_
timestamp 1728341909
transform -1 0 1090 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2852_
timestamp 1728341909
transform -1 0 1150 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2853_
timestamp 1728341909
transform -1 0 2350 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2854_
timestamp 1728341909
transform 1 0 830 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__2855_
timestamp 1728341909
transform 1 0 2510 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__2856_
timestamp 1728341909
transform -1 0 2030 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__2857_
timestamp 1728341909
transform -1 0 2430 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__2858_
timestamp 1728341909
transform -1 0 2330 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__2859_
timestamp 1728341909
transform -1 0 910 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2860_
timestamp 1728341909
transform 1 0 590 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2861_
timestamp 1728341909
transform -1 0 150 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2862_
timestamp 1728341909
transform -1 0 1110 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__2863_
timestamp 1728341909
transform 1 0 350 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__2864_
timestamp 1728341909
transform -1 0 390 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__2865_
timestamp 1728341909
transform 1 0 4510 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__2866_
timestamp 1728341909
transform 1 0 4530 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2867_
timestamp 1728341909
transform 1 0 5630 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__2868_
timestamp 1728341909
transform -1 0 3010 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2869_
timestamp 1728341909
transform -1 0 3290 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__2870_
timestamp 1728341909
transform -1 0 2350 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__2871_
timestamp 1728341909
transform 1 0 2370 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__2872_
timestamp 1728341909
transform -1 0 4650 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__2873_
timestamp 1728341909
transform 1 0 4390 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__2874_
timestamp 1728341909
transform -1 0 4190 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2875_
timestamp 1728341909
transform -1 0 1750 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2876_
timestamp 1728341909
transform -1 0 890 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2877_
timestamp 1728341909
transform -1 0 3550 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2878_
timestamp 1728341909
transform -1 0 3990 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2879_
timestamp 1728341909
transform -1 0 1330 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2880_
timestamp 1728341909
transform 1 0 1510 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2881_
timestamp 1728341909
transform -1 0 1830 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2882_
timestamp 1728341909
transform -1 0 2510 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2883_
timestamp 1728341909
transform 1 0 4510 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2884_
timestamp 1728341909
transform 1 0 4230 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2885_
timestamp 1728341909
transform 1 0 3170 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2886_
timestamp 1728341909
transform 1 0 4730 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2887_
timestamp 1728341909
transform 1 0 5190 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2888_
timestamp 1728341909
transform 1 0 3450 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2889_
timestamp 1728341909
transform 1 0 3670 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2890_
timestamp 1728341909
transform -1 0 4450 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2891_
timestamp 1728341909
transform -1 0 4190 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2892_
timestamp 1728341909
transform -1 0 2050 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2893_
timestamp 1728341909
transform 1 0 3730 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2894_
timestamp 1728341909
transform 1 0 3930 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2895_
timestamp 1728341909
transform 1 0 4510 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2896_
timestamp 1728341909
transform -1 0 3910 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2897_
timestamp 1728341909
transform -1 0 5910 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2898_
timestamp 1728341909
transform 1 0 5230 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2899_
timestamp 1728341909
transform 1 0 5190 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2900_
timestamp 1728341909
transform 1 0 5450 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2901_
timestamp 1728341909
transform -1 0 4930 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2902_
timestamp 1728341909
transform -1 0 1590 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2903_
timestamp 1728341909
transform 1 0 2250 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2904_
timestamp 1728341909
transform 1 0 2510 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2905_
timestamp 1728341909
transform 1 0 1310 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2906_
timestamp 1728341909
transform 1 0 1090 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2907_
timestamp 1728341909
transform 1 0 1290 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2908_
timestamp 1728341909
transform -1 0 1610 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2909_
timestamp 1728341909
transform -1 0 1830 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2910_
timestamp 1728341909
transform -1 0 1610 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2911_
timestamp 1728341909
transform -1 0 1610 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2912_
timestamp 1728341909
transform -1 0 2530 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2913_
timestamp 1728341909
transform -1 0 1770 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2914_
timestamp 1728341909
transform 1 0 2290 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2915_
timestamp 1728341909
transform 1 0 2070 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2916_
timestamp 1728341909
transform 1 0 1750 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2917_
timestamp 1728341909
transform -1 0 1830 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2918_
timestamp 1728341909
transform 1 0 1770 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2919_
timestamp 1728341909
transform -1 0 2310 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2920_
timestamp 1728341909
transform -1 0 2030 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2921_
timestamp 1728341909
transform -1 0 2090 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2922_
timestamp 1728341909
transform -1 0 2010 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2923_
timestamp 1728341909
transform -1 0 2050 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2924_
timestamp 1728341909
transform -1 0 3010 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2925_
timestamp 1728341909
transform 1 0 3490 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2926_
timestamp 1728341909
transform -1 0 2470 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2927_
timestamp 1728341909
transform -1 0 2510 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2928_
timestamp 1728341909
transform 1 0 4650 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2929_
timestamp 1728341909
transform 1 0 3490 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2930_
timestamp 1728341909
transform -1 0 2770 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2931_
timestamp 1728341909
transform -1 0 3010 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2932_
timestamp 1728341909
transform 1 0 3210 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2933_
timestamp 1728341909
transform -1 0 2770 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2934_
timestamp 1728341909
transform 1 0 2990 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2935_
timestamp 1728341909
transform -1 0 1370 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2936_
timestamp 1728341909
transform -1 0 910 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2937_
timestamp 1728341909
transform 1 0 630 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2938_
timestamp 1728341909
transform 1 0 1790 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2939_
timestamp 1728341909
transform -1 0 1570 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2940_
timestamp 1728341909
transform 1 0 3230 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2941_
timestamp 1728341909
transform 1 0 3230 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2942_
timestamp 1728341909
transform -1 0 3450 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2943_
timestamp 1728341909
transform -1 0 3290 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2944_
timestamp 1728341909
transform -1 0 3790 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2945_
timestamp 1728341909
transform 1 0 3230 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__2946_
timestamp 1728341909
transform 1 0 3670 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__2947_
timestamp 1728341909
transform 1 0 3250 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2948_
timestamp 1728341909
transform -1 0 4250 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2949_
timestamp 1728341909
transform 1 0 3210 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__2950_
timestamp 1728341909
transform 1 0 2530 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2951_
timestamp 1728341909
transform -1 0 2770 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2952_
timestamp 1728341909
transform -1 0 3050 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2953_
timestamp 1728341909
transform -1 0 2250 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2954_
timestamp 1728341909
transform -1 0 2490 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2955_
timestamp 1728341909
transform 1 0 3070 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__2956_
timestamp 1728341909
transform 1 0 3310 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__2957_
timestamp 1728341909
transform 1 0 3810 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__2958_
timestamp 1728341909
transform 1 0 2250 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__2959_
timestamp 1728341909
transform 1 0 3530 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__2960_
timestamp 1728341909
transform 1 0 3650 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__2961_
timestamp 1728341909
transform 1 0 2770 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2962_
timestamp 1728341909
transform 1 0 2510 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2963_
timestamp 1728341909
transform 1 0 3030 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2964_
timestamp 1728341909
transform 1 0 2770 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2965_
timestamp 1728341909
transform -1 0 5850 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2966_
timestamp 1728341909
transform 1 0 4170 0 1 1690
box -12 -8 32 252
use FILL  FILL_6__2967_
timestamp 1728341909
transform -1 0 4650 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2968_
timestamp 1728341909
transform -1 0 4890 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2969_
timestamp 1728341909
transform -1 0 1390 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__2970_
timestamp 1728341909
transform -1 0 1570 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__2971_
timestamp 1728341909
transform -1 0 1590 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2972_
timestamp 1728341909
transform -1 0 1330 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2973_
timestamp 1728341909
transform -1 0 1090 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__2974_
timestamp 1728341909
transform -1 0 1830 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2975_
timestamp 1728341909
transform -1 0 2050 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2976_
timestamp 1728341909
transform 1 0 3930 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2977_
timestamp 1728341909
transform -1 0 4490 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2978_
timestamp 1728341909
transform 1 0 4210 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2979_
timestamp 1728341909
transform 1 0 1590 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2980_
timestamp 1728341909
transform -1 0 1070 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2981_
timestamp 1728341909
transform -1 0 830 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2982_
timestamp 1728341909
transform 1 0 2270 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2983_
timestamp 1728341909
transform -1 0 590 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2984_
timestamp 1728341909
transform -1 0 370 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2985_
timestamp 1728341909
transform -1 0 150 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__2986_
timestamp 1728341909
transform -1 0 410 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2987_
timestamp 1728341909
transform -1 0 670 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2988_
timestamp 1728341909
transform -1 0 630 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2989_
timestamp 1728341909
transform 1 0 390 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2990_
timestamp 1728341909
transform 1 0 130 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2991_
timestamp 1728341909
transform -1 0 410 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2992_
timestamp 1728341909
transform -1 0 2070 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__2993_
timestamp 1728341909
transform -1 0 1110 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2994_
timestamp 1728341909
transform -1 0 870 0 1 730
box -12 -8 32 252
use FILL  FILL_6__2995_
timestamp 1728341909
transform 1 0 650 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__2996_
timestamp 1728341909
transform -1 0 590 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__2997_
timestamp 1728341909
transform -1 0 910 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__2998_
timestamp 1728341909
transform -1 0 150 0 1 250
box -12 -8 32 252
use FILL  FILL_6__2999_
timestamp 1728341909
transform -1 0 390 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__3000_
timestamp 1728341909
transform -1 0 150 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__3001_
timestamp 1728341909
transform -1 0 150 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__3002_
timestamp 1728341909
transform -1 0 630 0 1 730
box -12 -8 32 252
use FILL  FILL_6__3003_
timestamp 1728341909
transform -1 0 150 0 1 730
box -12 -8 32 252
use FILL  FILL_6__3004_
timestamp 1728341909
transform -1 0 890 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__3005_
timestamp 1728341909
transform 1 0 850 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__3006_
timestamp 1728341909
transform -1 0 150 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__3007_
timestamp 1728341909
transform 1 0 1850 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3008_
timestamp 1728341909
transform -1 0 1110 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__3009_
timestamp 1728341909
transform -1 0 1370 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__3010_
timestamp 1728341909
transform -1 0 1370 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__3011_
timestamp 1728341909
transform -1 0 1130 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6__3012_
timestamp 1728341909
transform -1 0 1510 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__3013_
timestamp 1728341909
transform -1 0 1290 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__3014_
timestamp 1728341909
transform 1 0 1090 0 1 250
box -12 -8 32 252
use FILL  FILL_6__3015_
timestamp 1728341909
transform -1 0 1590 0 1 250
box -12 -8 32 252
use FILL  FILL_6__3016_
timestamp 1728341909
transform -1 0 1350 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__3017_
timestamp 1728341909
transform -1 0 1330 0 1 250
box -12 -8 32 252
use FILL  FILL_6__3018_
timestamp 1728341909
transform 1 0 1110 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6__3019_
timestamp 1728341909
transform -1 0 1110 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__3020_
timestamp 1728341909
transform -1 0 3750 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3021_
timestamp 1728341909
transform -1 0 6010 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__3022_
timestamp 1728341909
transform 1 0 2850 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3023_
timestamp 1728341909
transform 1 0 2870 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3024_
timestamp 1728341909
transform 1 0 3850 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3025_
timestamp 1728341909
transform -1 0 4270 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__3026_
timestamp 1728341909
transform -1 0 3130 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3027_
timestamp 1728341909
transform -1 0 3530 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__3028_
timestamp 1728341909
transform -1 0 4050 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3029_
timestamp 1728341909
transform -1 0 4550 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3030_
timestamp 1728341909
transform 1 0 3530 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__3031_
timestamp 1728341909
transform -1 0 3810 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__3032_
timestamp 1728341909
transform -1 0 2610 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3033_
timestamp 1728341909
transform -1 0 2630 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3034_
timestamp 1728341909
transform 1 0 2770 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__3035_
timestamp 1728341909
transform -1 0 3030 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__3036_
timestamp 1728341909
transform 1 0 3350 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3037_
timestamp 1728341909
transform -1 0 3790 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__3038_
timestamp 1728341909
transform -1 0 3350 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3039_
timestamp 1728341909
transform 1 0 3090 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3040_
timestamp 1728341909
transform 1 0 2230 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__3041_
timestamp 1728341909
transform 1 0 2770 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__3042_
timestamp 1728341909
transform 1 0 7530 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__3043_
timestamp 1728341909
transform 1 0 6370 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__3044_
timestamp 1728341909
transform 1 0 5390 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__3045_
timestamp 1728341909
transform 1 0 5810 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3046_
timestamp 1728341909
transform 1 0 5530 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__3047_
timestamp 1728341909
transform 1 0 4870 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__3048_
timestamp 1728341909
transform 1 0 5210 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__3049_
timestamp 1728341909
transform 1 0 5910 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3050_
timestamp 1728341909
transform -1 0 6930 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3051_
timestamp 1728341909
transform -1 0 6390 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__3052_
timestamp 1728341909
transform 1 0 6430 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3053_
timestamp 1728341909
transform 1 0 6170 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3054_
timestamp 1728341909
transform 1 0 5910 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3055_
timestamp 1728341909
transform -1 0 6010 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3056_
timestamp 1728341909
transform 1 0 4670 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__3057_
timestamp 1728341909
transform 1 0 4430 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__3058_
timestamp 1728341909
transform -1 0 4550 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3059_
timestamp 1728341909
transform 1 0 4370 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__3060_
timestamp 1728341909
transform -1 0 4350 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__3061_
timestamp 1728341909
transform 1 0 4050 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3062_
timestamp 1728341909
transform -1 0 4870 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__3063_
timestamp 1728341909
transform 1 0 4610 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__3064_
timestamp 1728341909
transform 1 0 6070 0 1 2170
box -12 -8 32 252
use FILL  FILL_6__3065_
timestamp 1728341909
transform 1 0 5850 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__3066_
timestamp 1728341909
transform -1 0 5850 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3067_
timestamp 1728341909
transform -1 0 5990 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__3068_
timestamp 1728341909
transform -1 0 7030 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3069_
timestamp 1728341909
transform -1 0 6530 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3070_
timestamp 1728341909
transform 1 0 6170 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3071_
timestamp 1728341909
transform -1 0 6450 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3072_
timestamp 1728341909
transform 1 0 6650 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__3073_
timestamp 1728341909
transform 1 0 6410 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__3074_
timestamp 1728341909
transform 1 0 470 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__3075_
timestamp 1728341909
transform -1 0 630 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__3076_
timestamp 1728341909
transform -1 0 4330 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3077_
timestamp 1728341909
transform 1 0 2070 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3078_
timestamp 1728341909
transform -1 0 5570 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3079_
timestamp 1728341909
transform 1 0 5110 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3080_
timestamp 1728341909
transform 1 0 4310 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3081_
timestamp 1728341909
transform 1 0 5950 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__3082_
timestamp 1728341909
transform -1 0 6950 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__3083_
timestamp 1728341909
transform 1 0 6110 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__3084_
timestamp 1728341909
transform -1 0 5790 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3085_
timestamp 1728341909
transform -1 0 5070 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3086_
timestamp 1728341909
transform 1 0 5550 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3087_
timestamp 1728341909
transform -1 0 5150 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__3088_
timestamp 1728341909
transform -1 0 5690 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__3089_
timestamp 1728341909
transform -1 0 5650 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__3090_
timestamp 1728341909
transform 1 0 4830 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3091_
timestamp 1728341909
transform -1 0 4790 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3092_
timestamp 1728341909
transform 1 0 5650 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6__3093_
timestamp 1728341909
transform -1 0 4050 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__3094_
timestamp 1728341909
transform 1 0 4490 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__3095_
timestamp 1728341909
transform 1 0 4790 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__3096_
timestamp 1728341909
transform 1 0 4770 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__3097_
timestamp 1728341909
transform 1 0 5010 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__3098_
timestamp 1728341909
transform -1 0 5110 0 1 2650
box -12 -8 32 252
use FILL  FILL_6__3099_
timestamp 1728341909
transform 1 0 5250 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__3100_
timestamp 1728341909
transform -1 0 5650 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__3101_
timestamp 1728341909
transform 1 0 5190 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__3102_
timestamp 1728341909
transform 1 0 4710 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__3103_
timestamp 1728341909
transform 1 0 4930 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__3104_
timestamp 1728341909
transform -1 0 5070 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3105_
timestamp 1728341909
transform 1 0 5390 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__3106_
timestamp 1728341909
transform 1 0 8570 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__3107_
timestamp 1728341909
transform 1 0 8330 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__3108_
timestamp 1728341909
transform 1 0 8090 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__3109_
timestamp 1728341909
transform -1 0 8630 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3110_
timestamp 1728341909
transform -1 0 8390 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3111_
timestamp 1728341909
transform 1 0 4570 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3112_
timestamp 1728341909
transform 1 0 4810 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3113_
timestamp 1728341909
transform -1 0 1330 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3114_
timestamp 1728341909
transform 1 0 830 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3115_
timestamp 1728341909
transform 1 0 4510 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__3116_
timestamp 1728341909
transform -1 0 4130 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3117_
timestamp 1728341909
transform -1 0 390 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__3118_
timestamp 1728341909
transform -1 0 150 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__3119_
timestamp 1728341909
transform -1 0 4990 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__3120_
timestamp 1728341909
transform 1 0 4490 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3121_
timestamp 1728341909
transform 1 0 5230 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__3122_
timestamp 1728341909
transform -1 0 4530 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3123_
timestamp 1728341909
transform -1 0 3790 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3124_
timestamp 1728341909
transform -1 0 4010 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3125_
timestamp 1728341909
transform -1 0 3750 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3126_
timestamp 1728341909
transform 1 0 4770 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3127_
timestamp 1728341909
transform 1 0 4790 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3128_
timestamp 1728341909
transform 1 0 4710 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__3129_
timestamp 1728341909
transform 1 0 3790 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__3130_
timestamp 1728341909
transform -1 0 1890 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3131_
timestamp 1728341909
transform -1 0 1390 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3132_
timestamp 1728341909
transform 1 0 1110 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3133_
timestamp 1728341909
transform 1 0 3970 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3134_
timestamp 1728341909
transform 1 0 3550 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3135_
timestamp 1728341909
transform 1 0 3290 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3136_
timestamp 1728341909
transform 1 0 3770 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3137_
timestamp 1728341909
transform 1 0 4030 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3138_
timestamp 1728341909
transform -1 0 4070 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3139_
timestamp 1728341909
transform 1 0 1130 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3140_
timestamp 1728341909
transform 1 0 870 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3141_
timestamp 1728341909
transform -1 0 4050 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3142_
timestamp 1728341909
transform 1 0 3810 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3143_
timestamp 1728341909
transform -1 0 4250 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3144_
timestamp 1728341909
transform -1 0 3530 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3145_
timestamp 1728341909
transform 1 0 3270 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3146_
timestamp 1728341909
transform -1 0 3350 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3147_
timestamp 1728341909
transform 1 0 3590 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3148_
timestamp 1728341909
transform -1 0 3550 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3149_
timestamp 1728341909
transform -1 0 3530 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__3150_
timestamp 1728341909
transform 1 0 2110 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3151_
timestamp 1728341909
transform -1 0 2350 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3152_
timestamp 1728341909
transform 1 0 7590 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3153_
timestamp 1728341909
transform 1 0 4510 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3154_
timestamp 1728341909
transform -1 0 850 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3155_
timestamp 1728341909
transform 1 0 1070 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3156_
timestamp 1728341909
transform 1 0 3030 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3157_
timestamp 1728341909
transform -1 0 2810 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3158_
timestamp 1728341909
transform 1 0 2030 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3159_
timestamp 1728341909
transform 1 0 2570 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3160_
timestamp 1728341909
transform 1 0 3190 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3161_
timestamp 1728341909
transform -1 0 2730 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3162_
timestamp 1728341909
transform -1 0 2510 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3163_
timestamp 1728341909
transform -1 0 1610 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3164_
timestamp 1728341909
transform 1 0 1310 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3165_
timestamp 1728341909
transform -1 0 390 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3166_
timestamp 1728341909
transform -1 0 150 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3167_
timestamp 1728341909
transform 1 0 2110 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3168_
timestamp 1728341909
transform 1 0 2050 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3169_
timestamp 1728341909
transform -1 0 2350 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3170_
timestamp 1728341909
transform 1 0 2090 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3171_
timestamp 1728341909
transform -1 0 2290 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3172_
timestamp 1728341909
transform 1 0 1950 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__3173_
timestamp 1728341909
transform -1 0 1830 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3174_
timestamp 1728341909
transform -1 0 1850 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3175_
timestamp 1728341909
transform -1 0 3090 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3176_
timestamp 1728341909
transform -1 0 2890 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3177_
timestamp 1728341909
transform 1 0 2330 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3178_
timestamp 1728341909
transform 1 0 2670 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3179_
timestamp 1728341909
transform 1 0 2330 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3180_
timestamp 1728341909
transform 1 0 3270 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3181_
timestamp 1728341909
transform -1 0 2990 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3182_
timestamp 1728341909
transform -1 0 3070 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3183_
timestamp 1728341909
transform 1 0 2830 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3184_
timestamp 1728341909
transform -1 0 2590 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3185_
timestamp 1728341909
transform -1 0 2590 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3186_
timestamp 1728341909
transform 1 0 2070 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3187_
timestamp 1728341909
transform -1 0 410 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3188_
timestamp 1728341909
transform -1 0 150 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3189_
timestamp 1728341909
transform 1 0 1090 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3190_
timestamp 1728341909
transform -1 0 890 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3191_
timestamp 1728341909
transform -1 0 1150 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3192_
timestamp 1728341909
transform 1 0 1770 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3193_
timestamp 1728341909
transform 1 0 1510 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3194_
timestamp 1728341909
transform 1 0 3310 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3195_
timestamp 1728341909
transform 1 0 3270 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__3196_
timestamp 1728341909
transform 1 0 2010 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3197_
timestamp 1728341909
transform -1 0 2590 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__3198_
timestamp 1728341909
transform -1 0 2170 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3199_
timestamp 1728341909
transform -1 0 2430 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3200_
timestamp 1728341909
transform 1 0 870 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3201_
timestamp 1728341909
transform -1 0 1110 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3202_
timestamp 1728341909
transform 1 0 1110 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3203_
timestamp 1728341909
transform -1 0 1370 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3204_
timestamp 1728341909
transform -1 0 630 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3205_
timestamp 1728341909
transform -1 0 630 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3206_
timestamp 1728341909
transform 1 0 1130 0 -1 4090
box -12 -8 32 252
use FILL  FILL_6__3207_
timestamp 1728341909
transform -1 0 390 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3208_
timestamp 1728341909
transform -1 0 150 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3209_
timestamp 1728341909
transform 1 0 370 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3210_
timestamp 1728341909
transform -1 0 150 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3211_
timestamp 1728341909
transform -1 0 1630 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3212_
timestamp 1728341909
transform -1 0 1370 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3213_
timestamp 1728341909
transform 1 0 1650 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3214_
timestamp 1728341909
transform 1 0 1390 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3215_
timestamp 1728341909
transform -1 0 1350 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3216_
timestamp 1728341909
transform 1 0 1090 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3217_
timestamp 1728341909
transform -1 0 390 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3218_
timestamp 1728341909
transform -1 0 150 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3219_
timestamp 1728341909
transform -1 0 1670 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3220_
timestamp 1728341909
transform 1 0 1890 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3221_
timestamp 1728341909
transform -1 0 410 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3222_
timestamp 1728341909
transform -1 0 150 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3223_
timestamp 1728341909
transform -1 0 890 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__3224_
timestamp 1728341909
transform 1 0 610 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3225_
timestamp 1728341909
transform -1 0 390 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3226_
timestamp 1728341909
transform -1 0 150 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3227_
timestamp 1728341909
transform -1 0 410 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__3228_
timestamp 1728341909
transform -1 0 150 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__3229_
timestamp 1728341909
transform -1 0 2070 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__3230_
timestamp 1728341909
transform 1 0 1790 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__3231_
timestamp 1728341909
transform 1 0 1590 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__3232_
timestamp 1728341909
transform -1 0 1850 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__3233_
timestamp 1728341909
transform 1 0 1150 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3234_
timestamp 1728341909
transform -1 0 1430 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3235_
timestamp 1728341909
transform 1 0 1110 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3236_
timestamp 1728341909
transform 1 0 1370 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3237_
timestamp 1728341909
transform 1 0 2290 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__3238_
timestamp 1728341909
transform 1 0 2530 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6__3239_
timestamp 1728341909
transform -1 0 630 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3240_
timestamp 1728341909
transform -1 0 870 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3241_
timestamp 1728341909
transform 1 0 9770 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__3242_
timestamp 1728341909
transform -1 0 9110 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6__3243_
timestamp 1728341909
transform 1 0 9530 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__3244_
timestamp 1728341909
transform 1 0 8830 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__3245_
timestamp 1728341909
transform 1 0 9130 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3246_
timestamp 1728341909
transform -1 0 9650 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3247_
timestamp 1728341909
transform 1 0 10550 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3248_
timestamp 1728341909
transform 1 0 10810 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3249_
timestamp 1728341909
transform -1 0 9550 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__3250_
timestamp 1728341909
transform 1 0 9470 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3251_
timestamp 1728341909
transform 1 0 9310 0 1 3130
box -12 -8 32 252
use FILL  FILL_6__3252_
timestamp 1728341909
transform -1 0 9330 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__3253_
timestamp 1728341909
transform -1 0 7950 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3254_
timestamp 1728341909
transform -1 0 8210 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3255_
timestamp 1728341909
transform -1 0 9390 0 1 3610
box -12 -8 32 252
use FILL  FILL_6__3256_
timestamp 1728341909
transform 1 0 8330 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3257_
timestamp 1728341909
transform 1 0 8090 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3258_
timestamp 1728341909
transform 1 0 8630 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3259_
timestamp 1728341909
transform 1 0 9570 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3260_
timestamp 1728341909
transform -1 0 10930 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__3261_
timestamp 1728341909
transform -1 0 10470 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3262_
timestamp 1728341909
transform 1 0 10050 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3263_
timestamp 1728341909
transform 1 0 9730 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__3264_
timestamp 1728341909
transform 1 0 9070 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6__3265_
timestamp 1728341909
transform -1 0 9810 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3266_
timestamp 1728341909
transform 1 0 9830 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3267_
timestamp 1728341909
transform -1 0 9730 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3268_
timestamp 1728341909
transform -1 0 10070 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3269_
timestamp 1728341909
transform -1 0 10570 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3270_
timestamp 1728341909
transform 1 0 10290 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3271_
timestamp 1728341909
transform -1 0 10110 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6__3272_
timestamp 1728341909
transform 1 0 10330 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6__3273_
timestamp 1728341909
transform -1 0 10230 0 1 4570
box -12 -8 32 252
use FILL  FILL_6__3274_
timestamp 1728341909
transform -1 0 10330 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3275_
timestamp 1728341909
transform 1 0 9650 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__3276_
timestamp 1728341909
transform -1 0 9270 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3277_
timestamp 1728341909
transform -1 0 10730 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3278_
timestamp 1728341909
transform 1 0 10190 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3279_
timestamp 1728341909
transform -1 0 9970 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3280_
timestamp 1728341909
transform 1 0 9310 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__3281_
timestamp 1728341909
transform 1 0 9070 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__3282_
timestamp 1728341909
transform -1 0 6950 0 1 4090
box -12 -8 32 252
use FILL  FILL_6__3283_
timestamp 1728341909
transform -1 0 6890 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3284_
timestamp 1728341909
transform 1 0 6650 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6__3285_
timestamp 1728341909
transform 1 0 7090 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3286_
timestamp 1728341909
transform -1 0 7350 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3287_
timestamp 1728341909
transform -1 0 6710 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3288_
timestamp 1728341909
transform -1 0 6930 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3289_
timestamp 1728341909
transform -1 0 6890 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__3290_
timestamp 1728341909
transform 1 0 6610 0 1 5530
box -12 -8 32 252
use FILL  FILL_6__3291_
timestamp 1728341909
transform 1 0 7110 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3292_
timestamp 1728341909
transform -1 0 7370 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3293_
timestamp 1728341909
transform 1 0 7210 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3294_
timestamp 1728341909
transform 1 0 6950 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3295_
timestamp 1728341909
transform 1 0 6150 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3296_
timestamp 1728341909
transform 1 0 5890 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3297_
timestamp 1728341909
transform 1 0 5510 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3298_
timestamp 1728341909
transform 1 0 5250 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3299_
timestamp 1728341909
transform 1 0 5690 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3300_
timestamp 1728341909
transform 1 0 5450 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3301_
timestamp 1728341909
transform 1 0 6950 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6__3302_
timestamp 1728341909
transform 1 0 3030 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3303_
timestamp 1728341909
transform -1 0 3090 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3304_
timestamp 1728341909
transform 1 0 2030 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3305_
timestamp 1728341909
transform -1 0 2290 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3306_
timestamp 1728341909
transform 1 0 3950 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3307_
timestamp 1728341909
transform -1 0 4890 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3308_
timestamp 1728341909
transform -1 0 150 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__3309_
timestamp 1728341909
transform -1 0 150 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3310_
timestamp 1728341909
transform -1 0 830 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__3311_
timestamp 1728341909
transform -1 0 870 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3312_
timestamp 1728341909
transform -1 0 370 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__3313_
timestamp 1728341909
transform -1 0 410 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3314_
timestamp 1728341909
transform -1 0 150 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3315_
timestamp 1728341909
transform -1 0 150 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3316_
timestamp 1728341909
transform -1 0 650 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3317_
timestamp 1728341909
transform -1 0 870 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3449_
timestamp 1728341909
transform -1 0 3890 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3450_
timestamp 1728341909
transform 1 0 3050 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3451_
timestamp 1728341909
transform 1 0 3170 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3452_
timestamp 1728341909
transform -1 0 3430 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3453_
timestamp 1728341909
transform 1 0 3290 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3454_
timestamp 1728341909
transform -1 0 3650 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3455_
timestamp 1728341909
transform 1 0 10030 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3456_
timestamp 1728341909
transform 1 0 9590 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3457_
timestamp 1728341909
transform -1 0 9870 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3458_
timestamp 1728341909
transform -1 0 10030 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3459_
timestamp 1728341909
transform 1 0 10470 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3460_
timestamp 1728341909
transform -1 0 10770 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3461_
timestamp 1728341909
transform -1 0 10530 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3462_
timestamp 1728341909
transform -1 0 10090 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3463_
timestamp 1728341909
transform 1 0 10490 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3464_
timestamp 1728341909
transform -1 0 10290 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3465_
timestamp 1728341909
transform 1 0 10250 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6__3466_
timestamp 1728341909
transform -1 0 10270 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3467_
timestamp 1728341909
transform 1 0 8330 0 1 6010
box -12 -8 32 252
use FILL  FILL_6__3468_
timestamp 1728341909
transform 1 0 9170 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__3469_
timestamp 1728341909
transform 1 0 8630 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3470_
timestamp 1728341909
transform -1 0 8570 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3471_
timestamp 1728341909
transform 1 0 8710 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__3472_
timestamp 1728341909
transform 1 0 8950 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__3473_
timestamp 1728341909
transform -1 0 8770 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3474_
timestamp 1728341909
transform -1 0 8890 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3475_
timestamp 1728341909
transform -1 0 9010 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3476_
timestamp 1728341909
transform 1 0 9810 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3477_
timestamp 1728341909
transform 1 0 9250 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3478_
timestamp 1728341909
transform -1 0 9130 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3479_
timestamp 1728341909
transform 1 0 10610 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__3480_
timestamp 1728341909
transform -1 0 10170 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__3481_
timestamp 1728341909
transform -1 0 10030 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3482_
timestamp 1728341909
transform -1 0 9830 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__3483_
timestamp 1728341909
transform 1 0 10970 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3484_
timestamp 1728341909
transform 1 0 10950 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3485_
timestamp 1728341909
transform 1 0 11230 0 1 6490
box -12 -8 32 252
use FILL  FILL_6__3486_
timestamp 1728341909
transform 1 0 11190 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3487_
timestamp 1728341909
transform 1 0 10950 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3488_
timestamp 1728341909
transform 1 0 9590 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3489_
timestamp 1728341909
transform 1 0 9490 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3490_
timestamp 1728341909
transform -1 0 9750 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3491_
timestamp 1728341909
transform -1 0 9770 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3492_
timestamp 1728341909
transform 1 0 9970 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3493_
timestamp 1728341909
transform 1 0 10230 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3494_
timestamp 1728341909
transform 1 0 10370 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__3495_
timestamp 1728341909
transform -1 0 8870 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3496_
timestamp 1728341909
transform 1 0 9490 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3497_
timestamp 1728341909
transform 1 0 10010 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3498_
timestamp 1728341909
transform 1 0 9870 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__3499_
timestamp 1728341909
transform 1 0 9290 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3500_
timestamp 1728341909
transform -1 0 9550 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3501_
timestamp 1728341909
transform -1 0 9790 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3502_
timestamp 1728341909
transform 1 0 9630 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__3503_
timestamp 1728341909
transform 1 0 10110 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__3504_
timestamp 1728341909
transform -1 0 10070 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3505_
timestamp 1728341909
transform 1 0 10310 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3506_
timestamp 1728341909
transform 1 0 10830 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__3507_
timestamp 1728341909
transform -1 0 9450 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__3508_
timestamp 1728341909
transform -1 0 8570 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3509_
timestamp 1728341909
transform 1 0 8490 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__3510_
timestamp 1728341909
transform 1 0 9270 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3511_
timestamp 1728341909
transform -1 0 9030 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3512_
timestamp 1728341909
transform 1 0 8770 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3513_
timestamp 1728341909
transform -1 0 9050 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3514_
timestamp 1728341909
transform -1 0 8810 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3515_
timestamp 1728341909
transform -1 0 9210 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__3516_
timestamp 1728341909
transform 1 0 11050 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__3517_
timestamp 1728341909
transform -1 0 10370 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__3518_
timestamp 1728341909
transform 1 0 10450 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3519_
timestamp 1728341909
transform 1 0 10930 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3520_
timestamp 1728341909
transform -1 0 11230 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3521_
timestamp 1728341909
transform 1 0 7550 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3522_
timestamp 1728341909
transform -1 0 8070 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3523_
timestamp 1728341909
transform 1 0 8810 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3524_
timestamp 1728341909
transform 1 0 8590 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3525_
timestamp 1728341909
transform 1 0 9010 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3526_
timestamp 1728341909
transform -1 0 9290 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3527_
timestamp 1728341909
transform -1 0 8350 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3528_
timestamp 1728341909
transform -1 0 9990 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3529_
timestamp 1728341909
transform 1 0 10090 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__3530_
timestamp 1728341909
transform 1 0 10190 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3531_
timestamp 1728341909
transform -1 0 10230 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3532_
timestamp 1728341909
transform 1 0 10370 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__3533_
timestamp 1728341909
transform -1 0 8290 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3534_
timestamp 1728341909
transform -1 0 8550 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3535_
timestamp 1728341909
transform -1 0 8110 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3536_
timestamp 1728341909
transform -1 0 8330 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3537_
timestamp 1728341909
transform 1 0 8430 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__3538_
timestamp 1728341909
transform -1 0 8710 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__3539_
timestamp 1728341909
transform -1 0 9610 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__3540_
timestamp 1728341909
transform 1 0 9830 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__3541_
timestamp 1728341909
transform -1 0 9910 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__3542_
timestamp 1728341909
transform -1 0 7570 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3543_
timestamp 1728341909
transform -1 0 7830 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3544_
timestamp 1728341909
transform 1 0 8050 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3545_
timestamp 1728341909
transform 1 0 8910 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__3546_
timestamp 1728341909
transform -1 0 8350 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3547_
timestamp 1728341909
transform 1 0 8770 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3548_
timestamp 1728341909
transform -1 0 9030 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3549_
timestamp 1728341909
transform -1 0 8990 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__3550_
timestamp 1728341909
transform 1 0 8970 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3551_
timestamp 1728341909
transform 1 0 9250 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3552_
timestamp 1728341909
transform 1 0 9390 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__3553_
timestamp 1728341909
transform 1 0 9130 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__3554_
timestamp 1728341909
transform 1 0 9050 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__3555_
timestamp 1728341909
transform -1 0 8630 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3556_
timestamp 1728341909
transform 1 0 8530 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3557_
timestamp 1728341909
transform -1 0 8190 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__3558_
timestamp 1728341909
transform -1 0 7830 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3559_
timestamp 1728341909
transform 1 0 7790 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3560_
timestamp 1728341909
transform 1 0 8310 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3561_
timestamp 1728341909
transform -1 0 8050 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3562_
timestamp 1728341909
transform -1 0 9050 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3563_
timestamp 1728341909
transform -1 0 9030 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__3564_
timestamp 1728341909
transform 1 0 10130 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__3565_
timestamp 1728341909
transform -1 0 10050 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__3566_
timestamp 1728341909
transform 1 0 9970 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3567_
timestamp 1728341909
transform 1 0 10050 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__3568_
timestamp 1728341909
transform 1 0 10270 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__3569_
timestamp 1728341909
transform 1 0 10270 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__3570_
timestamp 1728341909
transform 1 0 10730 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__3571_
timestamp 1728341909
transform -1 0 10710 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3572_
timestamp 1728341909
transform -1 0 11210 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3573_
timestamp 1728341909
transform 1 0 11090 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__3574_
timestamp 1728341909
transform 1 0 10830 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__3575_
timestamp 1728341909
transform 1 0 11230 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__3576_
timestamp 1728341909
transform 1 0 10010 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__3577_
timestamp 1728341909
transform -1 0 11250 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__3578_
timestamp 1728341909
transform 1 0 10850 0 -1 9850
box -12 -8 32 252
use FILL  FILL_6__3579_
timestamp 1728341909
transform -1 0 10550 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__3580_
timestamp 1728341909
transform -1 0 9250 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3581_
timestamp 1728341909
transform -1 0 8950 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__3582_
timestamp 1728341909
transform 1 0 8790 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__3583_
timestamp 1728341909
transform -1 0 9110 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__3584_
timestamp 1728341909
transform 1 0 8850 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__3585_
timestamp 1728341909
transform -1 0 9590 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__3586_
timestamp 1728341909
transform 1 0 9170 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__3587_
timestamp 1728341909
transform -1 0 9310 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__3588_
timestamp 1728341909
transform 1 0 9330 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__3589_
timestamp 1728341909
transform 1 0 10050 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__3590_
timestamp 1728341909
transform -1 0 10310 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__3591_
timestamp 1728341909
transform 1 0 9790 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__3592_
timestamp 1728341909
transform 1 0 9810 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__3593_
timestamp 1728341909
transform -1 0 9590 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__3594_
timestamp 1728341909
transform 1 0 10430 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3595_
timestamp 1728341909
transform 1 0 10990 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__3596_
timestamp 1728341909
transform -1 0 10950 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3597_
timestamp 1728341909
transform 1 0 10590 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__3598_
timestamp 1728341909
transform 1 0 11230 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__3599_
timestamp 1728341909
transform 1 0 11190 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3600_
timestamp 1728341909
transform 1 0 11070 0 -1 9370
box -12 -8 32 252
use FILL  FILL_6__3601_
timestamp 1728341909
transform 1 0 10250 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3602_
timestamp 1728341909
transform 1 0 10490 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3603_
timestamp 1728341909
transform 1 0 10550 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3604_
timestamp 1728341909
transform 1 0 10770 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3605_
timestamp 1728341909
transform 1 0 11250 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3606_
timestamp 1728341909
transform 1 0 10730 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3607_
timestamp 1728341909
transform -1 0 10030 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3608_
timestamp 1728341909
transform -1 0 10270 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3609_
timestamp 1728341909
transform 1 0 10770 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3610_
timestamp 1728341909
transform 1 0 9590 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3611_
timestamp 1728341909
transform 1 0 9390 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__3612_
timestamp 1728341909
transform 1 0 9650 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__3613_
timestamp 1728341909
transform 1 0 9510 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3614_
timestamp 1728341909
transform -1 0 9910 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__3615_
timestamp 1728341909
transform -1 0 9790 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3616_
timestamp 1728341909
transform -1 0 9090 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3617_
timestamp 1728341909
transform -1 0 9350 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3618_
timestamp 1728341909
transform 1 0 9830 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3619_
timestamp 1728341909
transform 1 0 10990 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3620_
timestamp 1728341909
transform -1 0 10730 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3621_
timestamp 1728341909
transform -1 0 10510 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3622_
timestamp 1728341909
transform 1 0 10750 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3623_
timestamp 1728341909
transform 1 0 10050 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3624_
timestamp 1728341909
transform 1 0 10770 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3625_
timestamp 1728341909
transform 1 0 10870 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__3626_
timestamp 1728341909
transform -1 0 10770 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3627_
timestamp 1728341909
transform -1 0 9750 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3628_
timestamp 1728341909
transform -1 0 10490 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3629_
timestamp 1728341909
transform 1 0 10710 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3630_
timestamp 1728341909
transform 1 0 10510 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3631_
timestamp 1728341909
transform -1 0 10670 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__3632_
timestamp 1728341909
transform -1 0 11010 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__3633_
timestamp 1728341909
transform 1 0 10970 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__3634_
timestamp 1728341909
transform -1 0 10790 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__3635_
timestamp 1728341909
transform -1 0 10510 0 1 10810
box -12 -8 32 252
use FILL  FILL_6__3636_
timestamp 1728341909
transform -1 0 10610 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__3637_
timestamp 1728341909
transform -1 0 10770 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__3638_
timestamp 1728341909
transform -1 0 10690 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3639_
timestamp 1728341909
transform -1 0 10530 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__3640_
timestamp 1728341909
transform -1 0 10990 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3641_
timestamp 1728341909
transform -1 0 10730 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3642_
timestamp 1728341909
transform -1 0 11050 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3643_
timestamp 1728341909
transform 1 0 10970 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3644_
timestamp 1728341909
transform -1 0 10530 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3645_
timestamp 1728341909
transform -1 0 10270 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3646_
timestamp 1728341909
transform -1 0 11030 0 -1 8890
box -12 -8 32 252
use FILL  FILL_6__3647_
timestamp 1728341909
transform 1 0 11130 0 1 250
box -12 -8 32 252
use FILL  FILL_6__3648_
timestamp 1728341909
transform 1 0 11210 0 1 8410
box -12 -8 32 252
use FILL  FILL_6__3649_
timestamp 1728341909
transform 1 0 10290 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3650_
timestamp 1728341909
transform 1 0 10410 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__3651_
timestamp 1728341909
transform 1 0 10510 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3652_
timestamp 1728341909
transform -1 0 10470 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3653_
timestamp 1728341909
transform 1 0 10690 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3654_
timestamp 1728341909
transform 1 0 8490 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3655_
timestamp 1728341909
transform -1 0 8750 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3656_
timestamp 1728341909
transform 1 0 8330 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__3657_
timestamp 1728341909
transform -1 0 8710 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__3658_
timestamp 1728341909
transform -1 0 8610 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__3659_
timestamp 1728341909
transform -1 0 8350 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6__3660_
timestamp 1728341909
transform -1 0 8470 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__3661_
timestamp 1728341909
transform -1 0 9330 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__3662_
timestamp 1728341909
transform -1 0 9570 0 1 10330
box -12 -8 32 252
use FILL  FILL_6__3663_
timestamp 1728341909
transform 1 0 9490 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3664_
timestamp 1728341909
transform -1 0 9730 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3665_
timestamp 1728341909
transform 1 0 8330 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3666_
timestamp 1728341909
transform -1 0 8570 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3667_
timestamp 1728341909
transform -1 0 9290 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3668_
timestamp 1728341909
transform -1 0 10510 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3669_
timestamp 1728341909
transform -1 0 10250 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3670_
timestamp 1728341909
transform -1 0 10010 0 1 9370
box -12 -8 32 252
use FILL  FILL_6__3671_
timestamp 1728341909
transform 1 0 8370 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3672_
timestamp 1728341909
transform 1 0 8610 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3673_
timestamp 1728341909
transform -1 0 9530 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3674_
timestamp 1728341909
transform -1 0 9990 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3675_
timestamp 1728341909
transform 1 0 10210 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3676_
timestamp 1728341909
transform -1 0 10250 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3677_
timestamp 1728341909
transform 1 0 9490 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3678_
timestamp 1728341909
transform -1 0 9330 0 -1 6970
box -12 -8 32 252
use FILL  FILL_6__3691_
timestamp 1728341909
transform 1 0 7810 0 1 250
box -12 -8 32 252
use FILL  FILL_6__3692_
timestamp 1728341909
transform -1 0 8070 0 1 250
box -12 -8 32 252
use FILL  FILL_6__3693_
timestamp 1728341909
transform -1 0 2050 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3694_
timestamp 1728341909
transform -1 0 150 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3695_
timestamp 1728341909
transform 1 0 650 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3696_
timestamp 1728341909
transform -1 0 150 0 1 9850
box -12 -8 32 252
use FILL  FILL_6__3697_
timestamp 1728341909
transform -1 0 150 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__3698_
timestamp 1728341909
transform -1 0 390 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6__3699_
timestamp 1728341909
transform 1 0 6210 0 1 1210
box -12 -8 32 252
use FILL  FILL_6__3700_
timestamp 1728341909
transform -1 0 6370 0 -1 730
box -12 -8 32 252
use FILL  FILL_6__3701_
timestamp 1728341909
transform -1 0 6350 0 1 250
box -12 -8 32 252
use FILL  FILL_6__3702_
timestamp 1728341909
transform -1 0 5330 0 1 5050
box -12 -8 32 252
use FILL  FILL_6__3703_
timestamp 1728341909
transform -1 0 3570 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__3704_
timestamp 1728341909
transform -1 0 3350 0 -1 250
box -12 -8 32 252
use FILL  FILL_6__3705_
timestamp 1728341909
transform -1 0 150 0 1 8890
box -12 -8 32 252
use FILL  FILL_6__3706_
timestamp 1728341909
transform -1 0 1390 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6__3707_
timestamp 1728341909
transform 1 0 11210 0 1 6970
box -12 -8 32 252
use FILL  FILL_6__3708_
timestamp 1728341909
transform 1 0 11210 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6__3709_
timestamp 1728341909
transform 1 0 11230 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3710_
timestamp 1728341909
transform 1 0 10990 0 1 7450
box -12 -8 32 252
use FILL  FILL_6__3711_
timestamp 1728341909
transform 1 0 11210 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6__3712_
timestamp 1728341909
transform 1 0 10990 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3713_
timestamp 1728341909
transform 1 0 11110 0 1 7930
box -12 -8 32 252
use FILL  FILL_6__3714_
timestamp 1728341909
transform 1 0 11230 0 -1 8410
box -12 -8 32 252
use FILL  FILL_6__3715_
timestamp 1728341909
transform 1 0 11210 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert0
timestamp 1728341909
transform 1 0 7850 0 1 10810
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert1
timestamp 1728341909
transform 1 0 9070 0 1 1690
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert2
timestamp 1728341909
transform 1 0 9270 0 1 6970
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert3
timestamp 1728341909
transform 1 0 5750 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert4
timestamp 1728341909
transform 1 0 6850 0 1 1690
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert5
timestamp 1728341909
transform -1 0 4110 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert6
timestamp 1728341909
transform 1 0 7270 0 1 10330
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert7
timestamp 1728341909
transform -1 0 4190 0 1 4090
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert8
timestamp 1728341909
transform -1 0 7630 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert9
timestamp 1728341909
transform 1 0 4550 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert10
timestamp 1728341909
transform -1 0 670 0 1 4090
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert11
timestamp 1728341909
transform -1 0 4870 0 1 2650
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert12
timestamp 1728341909
transform 1 0 830 0 1 5530
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert13
timestamp 1728341909
transform -1 0 5970 0 1 7450
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert14
timestamp 1728341909
transform 1 0 4610 0 1 2650
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert15
timestamp 1728341909
transform 1 0 5690 0 -1 5050
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert16
timestamp 1728341909
transform 1 0 2770 0 1 8410
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert17
timestamp 1728341909
transform 1 0 4270 0 1 6490
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert18
timestamp 1728341909
transform -1 0 150 0 1 2650
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert19
timestamp 1728341909
transform -1 0 410 0 1 8410
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert20
timestamp 1728341909
transform 1 0 610 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert21
timestamp 1728341909
transform -1 0 7150 0 1 4570
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert22
timestamp 1728341909
transform -1 0 10530 0 1 4090
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert23
timestamp 1728341909
transform -1 0 8870 0 1 4090
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert24
timestamp 1728341909
transform 1 0 8590 0 1 3130
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert25
timestamp 1728341909
transform -1 0 7150 0 1 3130
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert37
timestamp 1728341909
transform -1 0 1070 0 1 5530
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert38
timestamp 1728341909
transform 1 0 1350 0 1 4570
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert39
timestamp 1728341909
transform -1 0 1110 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert40
timestamp 1728341909
transform -1 0 2810 0 -1 6010
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert41
timestamp 1728341909
transform 1 0 9610 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert42
timestamp 1728341909
transform 1 0 8930 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert43
timestamp 1728341909
transform -1 0 8850 0 -1 3610
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert44
timestamp 1728341909
transform -1 0 9070 0 1 4570
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert45
timestamp 1728341909
transform 1 0 3930 0 1 4090
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert46
timestamp 1728341909
transform 1 0 5290 0 1 4090
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert47
timestamp 1728341909
transform 1 0 4390 0 1 2650
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert48
timestamp 1728341909
transform 1 0 5510 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert49
timestamp 1728341909
transform -1 0 2310 0 1 2650
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert50
timestamp 1728341909
transform 1 0 8390 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert51
timestamp 1728341909
transform -1 0 10490 0 1 4570
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert52
timestamp 1728341909
transform -1 0 9530 0 1 4570
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert53
timestamp 1728341909
transform -1 0 9610 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert54
timestamp 1728341909
transform -1 0 8450 0 -1 3130
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert55
timestamp 1728341909
transform -1 0 410 0 1 730
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert56
timestamp 1728341909
transform 1 0 5090 0 -1 1210
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert57
timestamp 1728341909
transform 1 0 4690 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert58
timestamp 1728341909
transform 1 0 2010 0 1 1690
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert59
timestamp 1728341909
transform 1 0 4450 0 1 730
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert60
timestamp 1728341909
transform -1 0 8830 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert61
timestamp 1728341909
transform 1 0 10230 0 -1 7450
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert62
timestamp 1728341909
transform 1 0 9270 0 -1 10330
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert63
timestamp 1728341909
transform 1 0 9350 0 1 7450
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert64
timestamp 1728341909
transform 1 0 8690 0 1 1210
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert65
timestamp 1728341909
transform -1 0 5090 0 1 4090
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert66
timestamp 1728341909
transform 1 0 5830 0 1 2650
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert67
timestamp 1728341909
transform 1 0 6670 0 1 5050
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert68
timestamp 1728341909
transform 1 0 7670 0 -1 2650
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert69
timestamp 1728341909
transform -1 0 6150 0 1 1690
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert70
timestamp 1728341909
transform 1 0 8830 0 -1 2170
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert71
timestamp 1728341909
transform 1 0 2530 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert72
timestamp 1728341909
transform 1 0 3970 0 1 1210
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert73
timestamp 1728341909
transform 1 0 2770 0 1 2650
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert74
timestamp 1728341909
transform -1 0 3770 0 -1 1690
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert75
timestamp 1728341909
transform -1 0 850 0 1 2170
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert76
timestamp 1728341909
transform 1 0 8830 0 1 4570
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert77
timestamp 1728341909
transform -1 0 8570 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert78
timestamp 1728341909
transform 1 0 9030 0 -1 5530
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert79
timestamp 1728341909
transform -1 0 9290 0 1 4570
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert80
timestamp 1728341909
transform 1 0 4270 0 -1 6490
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert81
timestamp 1728341909
transform 1 0 3410 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert82
timestamp 1728341909
transform 1 0 2270 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6_BUFX2_insert83
timestamp 1728341909
transform -1 0 2750 0 -1 7930
box -12 -8 32 252
use FILL  FILL_6_CLKBUF1_insert26
timestamp 1728341909
transform -1 0 1490 0 1 3130
box -12 -8 32 252
use FILL  FILL_6_CLKBUF1_insert27
timestamp 1728341909
transform 1 0 3730 0 1 3130
box -12 -8 32 252
use FILL  FILL_6_CLKBUF1_insert28
timestamp 1728341909
transform 1 0 130 0 1 3130
box -12 -8 32 252
use FILL  FILL_6_CLKBUF1_insert29
timestamp 1728341909
transform 1 0 610 0 1 7930
box -12 -8 32 252
use FILL  FILL_6_CLKBUF1_insert30
timestamp 1728341909
transform 1 0 8290 0 1 5530
box -12 -8 32 252
use FILL  FILL_6_CLKBUF1_insert31
timestamp 1728341909
transform -1 0 7650 0 -1 10810
box -12 -8 32 252
use FILL  FILL_6_CLKBUF1_insert32
timestamp 1728341909
transform -1 0 3270 0 -1 4570
box -12 -8 32 252
use FILL  FILL_6_CLKBUF1_insert33
timestamp 1728341909
transform -1 0 8010 0 1 10330
box -12 -8 32 252
use FILL  FILL_6_CLKBUF1_insert34
timestamp 1728341909
transform -1 0 150 0 -1 11290
box -12 -8 32 252
use FILL  FILL_6_CLKBUF1_insert35
timestamp 1728341909
transform -1 0 5570 0 1 5050
box -12 -8 32 252
use FILL  FILL_6_CLKBUF1_insert36
timestamp 1728341909
transform -1 0 2950 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__1745_
timestamp 1728341909
transform 1 0 4330 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__1747_
timestamp 1728341909
transform -1 0 5770 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__1748_
timestamp 1728341909
transform 1 0 6690 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__1750_
timestamp 1728341909
transform 1 0 5290 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__1751_
timestamp 1728341909
transform 1 0 6930 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__1753_
timestamp 1728341909
transform 1 0 7650 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__1755_
timestamp 1728341909
transform -1 0 7410 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__1756_
timestamp 1728341909
transform -1 0 6490 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__1758_
timestamp 1728341909
transform 1 0 6910 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__1759_
timestamp 1728341909
transform -1 0 3170 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__1761_
timestamp 1728341909
transform 1 0 7390 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__1763_
timestamp 1728341909
transform -1 0 8310 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__1764_
timestamp 1728341909
transform -1 0 8130 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__1766_
timestamp 1728341909
transform -1 0 7930 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__1768_
timestamp 1728341909
transform -1 0 5810 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__1769_
timestamp 1728341909
transform 1 0 3250 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__1771_
timestamp 1728341909
transform 1 0 11150 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__1772_
timestamp 1728341909
transform 1 0 10890 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__1774_
timestamp 1728341909
transform 1 0 10790 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__1776_
timestamp 1728341909
transform 1 0 9650 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__1777_
timestamp 1728341909
transform -1 0 8830 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__1779_
timestamp 1728341909
transform 1 0 10250 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__1780_
timestamp 1728341909
transform 1 0 11010 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__1782_
timestamp 1728341909
transform -1 0 11270 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__1784_
timestamp 1728341909
transform 1 0 10650 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__1785_
timestamp 1728341909
transform 1 0 10990 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__1787_
timestamp 1728341909
transform 1 0 9330 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__1788_
timestamp 1728341909
transform 1 0 10610 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__1790_
timestamp 1728341909
transform -1 0 10830 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__1792_
timestamp 1728341909
transform 1 0 5750 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__1793_
timestamp 1728341909
transform 1 0 5470 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__1795_
timestamp 1728341909
transform 1 0 3830 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__1797_
timestamp 1728341909
transform -1 0 4810 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__1798_
timestamp 1728341909
transform -1 0 11130 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__1800_
timestamp 1728341909
transform -1 0 10550 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__1801_
timestamp 1728341909
transform -1 0 10210 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__1803_
timestamp 1728341909
transform 1 0 10330 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__1805_
timestamp 1728341909
transform -1 0 10130 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__1806_
timestamp 1728341909
transform 1 0 10070 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__1808_
timestamp 1728341909
transform -1 0 10490 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__1809_
timestamp 1728341909
transform -1 0 11150 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__1811_
timestamp 1728341909
transform -1 0 11230 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__1813_
timestamp 1728341909
transform -1 0 7790 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__1814_
timestamp 1728341909
transform -1 0 7630 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__1816_
timestamp 1728341909
transform -1 0 7690 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__1818_
timestamp 1728341909
transform 1 0 6750 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__1819_
timestamp 1728341909
transform 1 0 6250 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__1821_
timestamp 1728341909
transform -1 0 6810 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__1822_
timestamp 1728341909
transform 1 0 11230 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__1824_
timestamp 1728341909
transform 1 0 7390 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__1826_
timestamp 1728341909
transform 1 0 11030 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__1827_
timestamp 1728341909
transform -1 0 7470 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__1829_
timestamp 1728341909
transform -1 0 7490 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__1830_
timestamp 1728341909
transform 1 0 7630 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__1832_
timestamp 1728341909
transform 1 0 10750 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__1834_
timestamp 1728341909
transform -1 0 7110 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__1835_
timestamp 1728341909
transform -1 0 6550 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__1837_
timestamp 1728341909
transform -1 0 5630 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__1838_
timestamp 1728341909
transform 1 0 5350 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__1840_
timestamp 1728341909
transform -1 0 8130 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__1842_
timestamp 1728341909
transform -1 0 6930 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__1843_
timestamp 1728341909
transform 1 0 7250 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__1845_
timestamp 1728341909
transform 1 0 11230 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__1847_
timestamp 1728341909
transform -1 0 8170 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__1848_
timestamp 1728341909
transform 1 0 10770 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__1850_
timestamp 1728341909
transform -1 0 8630 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__1851_
timestamp 1728341909
transform -1 0 11250 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__1853_
timestamp 1728341909
transform 1 0 9330 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__1855_
timestamp 1728341909
transform 1 0 8890 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__1856_
timestamp 1728341909
transform 1 0 9410 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__1858_
timestamp 1728341909
transform 1 0 7370 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__1859_
timestamp 1728341909
transform -1 0 10790 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__1861_
timestamp 1728341909
transform 1 0 7410 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__1863_
timestamp 1728341909
transform 1 0 8650 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__1864_
timestamp 1728341909
transform 1 0 9950 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__1866_
timestamp 1728341909
transform -1 0 8990 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__1867_
timestamp 1728341909
transform 1 0 9370 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__1869_
timestamp 1728341909
transform 1 0 9390 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__1871_
timestamp 1728341909
transform 1 0 8610 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__1872_
timestamp 1728341909
transform 1 0 7890 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__1874_
timestamp 1728341909
transform -1 0 6910 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__1876_
timestamp 1728341909
transform 1 0 6730 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__1877_
timestamp 1728341909
transform -1 0 8150 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__1879_
timestamp 1728341909
transform -1 0 8150 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__1880_
timestamp 1728341909
transform -1 0 7090 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__1882_
timestamp 1728341909
transform 1 0 3570 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__1884_
timestamp 1728341909
transform -1 0 6630 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__1885_
timestamp 1728341909
transform 1 0 5910 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__1887_
timestamp 1728341909
transform 1 0 6930 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__1888_
timestamp 1728341909
transform 1 0 3690 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__1890_
timestamp 1728341909
transform 1 0 6510 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__1892_
timestamp 1728341909
transform 1 0 5710 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__1893_
timestamp 1728341909
transform 1 0 1110 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__1895_
timestamp 1728341909
transform 1 0 6930 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__1897_
timestamp 1728341909
transform 1 0 6090 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__1898_
timestamp 1728341909
transform 1 0 6510 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__1900_
timestamp 1728341909
transform 1 0 630 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__1901_
timestamp 1728341909
transform 1 0 8070 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__1903_
timestamp 1728341909
transform 1 0 7970 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__1905_
timestamp 1728341909
transform 1 0 7630 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__1906_
timestamp 1728341909
transform 1 0 7610 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__1908_
timestamp 1728341909
transform -1 0 7810 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__1909_
timestamp 1728341909
transform 1 0 1910 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__1911_
timestamp 1728341909
transform 1 0 9590 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__1913_
timestamp 1728341909
transform 1 0 10730 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__1914_
timestamp 1728341909
transform 1 0 10790 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__1916_
timestamp 1728341909
transform -1 0 5970 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__1917_
timestamp 1728341909
transform 1 0 4110 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__1919_
timestamp 1728341909
transform -1 0 170 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__1921_
timestamp 1728341909
transform -1 0 1290 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__1922_
timestamp 1728341909
transform -1 0 1030 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__1924_
timestamp 1728341909
transform -1 0 4570 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__1926_
timestamp 1728341909
transform 1 0 870 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__1927_
timestamp 1728341909
transform -1 0 2170 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__1929_
timestamp 1728341909
transform 1 0 370 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__1930_
timestamp 1728341909
transform 1 0 750 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__1932_
timestamp 1728341909
transform -1 0 650 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__1934_
timestamp 1728341909
transform -1 0 650 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__1935_
timestamp 1728341909
transform -1 0 1630 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__1937_
timestamp 1728341909
transform -1 0 650 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__1938_
timestamp 1728341909
transform -1 0 170 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__1940_
timestamp 1728341909
transform 1 0 910 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__1942_
timestamp 1728341909
transform 1 0 630 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__1943_
timestamp 1728341909
transform 1 0 8190 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__1945_
timestamp 1728341909
transform -1 0 7510 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__1947_
timestamp 1728341909
transform -1 0 7710 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__1948_
timestamp 1728341909
transform -1 0 7050 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__1950_
timestamp 1728341909
transform 1 0 8390 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__1951_
timestamp 1728341909
transform 1 0 8390 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__1953_
timestamp 1728341909
transform -1 0 8470 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__1955_
timestamp 1728341909
transform 1 0 6510 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__1956_
timestamp 1728341909
transform -1 0 8070 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__1958_
timestamp 1728341909
transform 1 0 10510 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__1959_
timestamp 1728341909
transform 1 0 7870 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__1961_
timestamp 1728341909
transform 1 0 10770 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__1963_
timestamp 1728341909
transform 1 0 9910 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__1964_
timestamp 1728341909
transform -1 0 7450 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__1966_
timestamp 1728341909
transform -1 0 3590 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__1967_
timestamp 1728341909
transform -1 0 7050 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__1969_
timestamp 1728341909
transform -1 0 7850 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__1971_
timestamp 1728341909
transform -1 0 890 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__1972_
timestamp 1728341909
transform 1 0 1410 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__1974_
timestamp 1728341909
transform 1 0 8430 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__1976_
timestamp 1728341909
transform -1 0 7210 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__1977_
timestamp 1728341909
transform -1 0 2910 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__1979_
timestamp 1728341909
transform -1 0 6590 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__1980_
timestamp 1728341909
transform 1 0 7850 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__1982_
timestamp 1728341909
transform -1 0 3110 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__1984_
timestamp 1728341909
transform 1 0 1870 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__1985_
timestamp 1728341909
transform 1 0 2530 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__1987_
timestamp 1728341909
transform 1 0 5150 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__1988_
timestamp 1728341909
transform -1 0 5050 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__1990_
timestamp 1728341909
transform -1 0 7330 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__1992_
timestamp 1728341909
transform -1 0 1630 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__1993_
timestamp 1728341909
transform -1 0 1910 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__1995_
timestamp 1728341909
transform 1 0 8110 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__1996_
timestamp 1728341909
transform -1 0 2330 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__1998_
timestamp 1728341909
transform -1 0 6570 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__2000_
timestamp 1728341909
transform 1 0 1890 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__2001_
timestamp 1728341909
transform 1 0 1370 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__2003_
timestamp 1728341909
transform 1 0 1630 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__2005_
timestamp 1728341909
transform 1 0 2070 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2006_
timestamp 1728341909
transform -1 0 6330 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__2008_
timestamp 1728341909
transform -1 0 8130 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__2009_
timestamp 1728341909
transform 1 0 870 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__2011_
timestamp 1728341909
transform 1 0 630 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__2013_
timestamp 1728341909
transform 1 0 5530 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2014_
timestamp 1728341909
transform 1 0 1830 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__2016_
timestamp 1728341909
transform 1 0 6830 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__2017_
timestamp 1728341909
transform -1 0 7370 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__2019_
timestamp 1728341909
transform -1 0 1670 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__2021_
timestamp 1728341909
transform 1 0 1810 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__2022_
timestamp 1728341909
transform 1 0 4590 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2024_
timestamp 1728341909
transform 1 0 1530 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__2026_
timestamp 1728341909
transform -1 0 4790 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__2027_
timestamp 1728341909
transform 1 0 7290 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2029_
timestamp 1728341909
transform -1 0 170 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__2030_
timestamp 1728341909
transform -1 0 650 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__2032_
timestamp 1728341909
transform 1 0 630 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__2034_
timestamp 1728341909
transform 1 0 1310 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__2035_
timestamp 1728341909
transform 1 0 2190 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2037_
timestamp 1728341909
transform -1 0 4190 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__2038_
timestamp 1728341909
transform 1 0 7630 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__2040_
timestamp 1728341909
transform -1 0 3030 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2042_
timestamp 1728341909
transform 1 0 1810 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__2043_
timestamp 1728341909
transform -1 0 3910 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__2045_
timestamp 1728341909
transform -1 0 4150 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__2046_
timestamp 1728341909
transform 1 0 2950 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__2048_
timestamp 1728341909
transform -1 0 3650 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__2050_
timestamp 1728341909
transform -1 0 2530 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__2051_
timestamp 1728341909
transform -1 0 2510 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2053_
timestamp 1728341909
transform -1 0 3490 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__2055_
timestamp 1728341909
transform -1 0 2850 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__2056_
timestamp 1728341909
transform 1 0 4470 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__2058_
timestamp 1728341909
transform 1 0 4690 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__2059_
timestamp 1728341909
transform -1 0 2050 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__2061_
timestamp 1728341909
transform 1 0 3610 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__2063_
timestamp 1728341909
transform 1 0 2570 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__2064_
timestamp 1728341909
transform -1 0 2670 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2066_
timestamp 1728341909
transform 1 0 2530 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2067_
timestamp 1728341909
transform -1 0 2850 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__2069_
timestamp 1728341909
transform 1 0 2630 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__2071_
timestamp 1728341909
transform -1 0 2890 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__2072_
timestamp 1728341909
transform -1 0 2630 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__2074_
timestamp 1728341909
transform 1 0 3310 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__2075_
timestamp 1728341909
transform -1 0 2790 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__2077_
timestamp 1728341909
transform -1 0 3350 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__2079_
timestamp 1728341909
transform -1 0 3990 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2080_
timestamp 1728341909
transform 1 0 4210 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2082_
timestamp 1728341909
transform 1 0 5850 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2084_
timestamp 1728341909
transform 1 0 10010 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2085_
timestamp 1728341909
transform -1 0 10530 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2087_
timestamp 1728341909
transform 1 0 11090 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__2088_
timestamp 1728341909
transform 1 0 10290 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2090_
timestamp 1728341909
transform 1 0 10770 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__2092_
timestamp 1728341909
transform -1 0 10230 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2093_
timestamp 1728341909
transform 1 0 10290 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__2095_
timestamp 1728341909
transform 1 0 10850 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__2096_
timestamp 1728341909
transform -1 0 11250 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__2098_
timestamp 1728341909
transform 1 0 10270 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2100_
timestamp 1728341909
transform 1 0 10970 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2101_
timestamp 1728341909
transform 1 0 11210 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2103_
timestamp 1728341909
transform 1 0 4330 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__2105_
timestamp 1728341909
transform -1 0 1850 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2106_
timestamp 1728341909
transform -1 0 2230 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2108_
timestamp 1728341909
transform 1 0 1550 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2109_
timestamp 1728341909
transform -1 0 2970 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2111_
timestamp 1728341909
transform 1 0 5390 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2113_
timestamp 1728341909
transform -1 0 9850 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__2114_
timestamp 1728341909
transform 1 0 9850 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__2116_
timestamp 1728341909
transform -1 0 11110 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__2117_
timestamp 1728341909
transform -1 0 10710 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__2119_
timestamp 1728341909
transform -1 0 11190 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__2121_
timestamp 1728341909
transform 1 0 11230 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2122_
timestamp 1728341909
transform 1 0 10930 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2124_
timestamp 1728341909
transform 1 0 9450 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__2125_
timestamp 1728341909
transform 1 0 9570 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2127_
timestamp 1728341909
transform 1 0 9830 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2129_
timestamp 1728341909
transform -1 0 9010 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__2130_
timestamp 1728341909
transform 1 0 9690 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__2132_
timestamp 1728341909
transform 1 0 10250 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2134_
timestamp 1728341909
transform -1 0 10190 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2135_
timestamp 1728341909
transform 1 0 10690 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2137_
timestamp 1728341909
transform 1 0 10890 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2138_
timestamp 1728341909
transform -1 0 10990 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2140_
timestamp 1728341909
transform -1 0 8410 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2142_
timestamp 1728341909
transform 1 0 1970 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2143_
timestamp 1728341909
transform -1 0 3010 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2145_
timestamp 1728341909
transform -1 0 6310 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2146_
timestamp 1728341909
transform 1 0 5610 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2148_
timestamp 1728341909
transform 1 0 9750 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2150_
timestamp 1728341909
transform -1 0 8590 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2151_
timestamp 1728341909
transform 1 0 8250 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__2153_
timestamp 1728341909
transform -1 0 9190 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2155_
timestamp 1728341909
transform 1 0 8090 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__2156_
timestamp 1728341909
transform -1 0 8370 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__2158_
timestamp 1728341909
transform 1 0 10410 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__2159_
timestamp 1728341909
transform 1 0 6110 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__2161_
timestamp 1728341909
transform 1 0 6670 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__2163_
timestamp 1728341909
transform -1 0 8430 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__2164_
timestamp 1728341909
transform 1 0 7190 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__2166_
timestamp 1728341909
transform -1 0 8230 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__2167_
timestamp 1728341909
transform -1 0 7930 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__2169_
timestamp 1728341909
transform 1 0 8230 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2171_
timestamp 1728341909
transform 1 0 8650 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2172_
timestamp 1728341909
transform -1 0 10510 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2174_
timestamp 1728341909
transform 1 0 4470 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2175_
timestamp 1728341909
transform -1 0 4030 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2177_
timestamp 1728341909
transform -1 0 6150 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2179_
timestamp 1728341909
transform 1 0 6450 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2180_
timestamp 1728341909
transform 1 0 7250 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2182_
timestamp 1728341909
transform -1 0 7250 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__2184_
timestamp 1728341909
transform 1 0 6550 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__2185_
timestamp 1728341909
transform -1 0 6690 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2187_
timestamp 1728341909
transform -1 0 9530 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__2188_
timestamp 1728341909
transform 1 0 9130 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__2190_
timestamp 1728341909
transform 1 0 8590 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__2192_
timestamp 1728341909
transform 1 0 7390 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2193_
timestamp 1728341909
transform 1 0 7610 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2195_
timestamp 1728341909
transform -1 0 8650 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__2196_
timestamp 1728341909
transform 1 0 8690 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__2198_
timestamp 1728341909
transform -1 0 7330 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__2200_
timestamp 1728341909
transform 1 0 9110 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__2201_
timestamp 1728341909
transform 1 0 8970 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2203_
timestamp 1728341909
transform 1 0 8490 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__2204_
timestamp 1728341909
transform -1 0 8490 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2206_
timestamp 1728341909
transform -1 0 8110 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2208_
timestamp 1728341909
transform -1 0 8370 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2209_
timestamp 1728341909
transform -1 0 7890 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2211_
timestamp 1728341909
transform -1 0 7290 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__2213_
timestamp 1728341909
transform -1 0 8070 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2214_
timestamp 1728341909
transform 1 0 8630 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2216_
timestamp 1728341909
transform 1 0 9310 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2217_
timestamp 1728341909
transform -1 0 9570 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2219_
timestamp 1728341909
transform -1 0 2330 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__2221_
timestamp 1728341909
transform 1 0 4190 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2222_
timestamp 1728341909
transform 1 0 4410 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2224_
timestamp 1728341909
transform -1 0 2910 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2225_
timestamp 1728341909
transform -1 0 5970 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2227_
timestamp 1728341909
transform -1 0 7070 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__2229_
timestamp 1728341909
transform 1 0 7870 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__2230_
timestamp 1728341909
transform -1 0 6270 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__2232_
timestamp 1728341909
transform 1 0 6930 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__2234_
timestamp 1728341909
transform 1 0 7410 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2235_
timestamp 1728341909
transform 1 0 9490 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2237_
timestamp 1728341909
transform 1 0 10030 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2238_
timestamp 1728341909
transform -1 0 9950 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2240_
timestamp 1728341909
transform 1 0 2770 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2242_
timestamp 1728341909
transform -1 0 4670 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2243_
timestamp 1728341909
transform 1 0 3450 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2245_
timestamp 1728341909
transform 1 0 7350 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2246_
timestamp 1728341909
transform 1 0 7370 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2248_
timestamp 1728341909
transform 1 0 3510 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2250_
timestamp 1728341909
transform 1 0 6750 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2251_
timestamp 1728341909
transform 1 0 7270 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2253_
timestamp 1728341909
transform 1 0 9430 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2254_
timestamp 1728341909
transform 1 0 5710 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2256_
timestamp 1728341909
transform 1 0 7210 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2258_
timestamp 1728341909
transform -1 0 3110 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__2259_
timestamp 1728341909
transform 1 0 3530 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2261_
timestamp 1728341909
transform -1 0 5710 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2263_
timestamp 1728341909
transform 1 0 4950 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2264_
timestamp 1728341909
transform -1 0 6250 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2266_
timestamp 1728341909
transform 1 0 7590 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__2267_
timestamp 1728341909
transform -1 0 5490 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__2269_
timestamp 1728341909
transform 1 0 5490 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__2271_
timestamp 1728341909
transform 1 0 6050 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__2272_
timestamp 1728341909
transform 1 0 5650 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__2274_
timestamp 1728341909
transform 1 0 5230 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__2275_
timestamp 1728341909
transform 1 0 5710 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__2277_
timestamp 1728341909
transform 1 0 7850 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__2279_
timestamp 1728341909
transform 1 0 6550 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__2280_
timestamp 1728341909
transform -1 0 6570 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2282_
timestamp 1728341909
transform 1 0 6610 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2283_
timestamp 1728341909
transform 1 0 7310 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2285_
timestamp 1728341909
transform 1 0 9710 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2287_
timestamp 1728341909
transform -1 0 1870 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2288_
timestamp 1728341909
transform -1 0 2310 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2290_
timestamp 1728341909
transform -1 0 1830 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2292_
timestamp 1728341909
transform 1 0 4170 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2293_
timestamp 1728341909
transform 1 0 4910 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2295_
timestamp 1728341909
transform -1 0 2310 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2296_
timestamp 1728341909
transform 1 0 3750 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2298_
timestamp 1728341909
transform 1 0 2050 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2300_
timestamp 1728341909
transform 1 0 3250 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2301_
timestamp 1728341909
transform -1 0 3710 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2303_
timestamp 1728341909
transform -1 0 5170 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2304_
timestamp 1728341909
transform 1 0 5410 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2306_
timestamp 1728341909
transform 1 0 2510 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2308_
timestamp 1728341909
transform -1 0 5670 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2309_
timestamp 1728341909
transform 1 0 4670 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2311_
timestamp 1728341909
transform -1 0 3830 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2313_
timestamp 1728341909
transform 1 0 5350 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2314_
timestamp 1728341909
transform 1 0 4530 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2316_
timestamp 1728341909
transform -1 0 9930 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2317_
timestamp 1728341909
transform 1 0 11230 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__2319_
timestamp 1728341909
transform -1 0 10550 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__2321_
timestamp 1728341909
transform 1 0 10650 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__2322_
timestamp 1728341909
transform 1 0 10550 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__2324_
timestamp 1728341909
transform 1 0 7010 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2325_
timestamp 1728341909
transform 1 0 9370 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__2327_
timestamp 1728341909
transform -1 0 9370 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__2329_
timestamp 1728341909
transform 1 0 9330 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2330_
timestamp 1728341909
transform -1 0 9090 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2332_
timestamp 1728341909
transform 1 0 9230 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2333_
timestamp 1728341909
transform 1 0 9490 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2335_
timestamp 1728341909
transform 1 0 5730 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2337_
timestamp 1728341909
transform -1 0 6030 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__2338_
timestamp 1728341909
transform -1 0 5970 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2340_
timestamp 1728341909
transform -1 0 9330 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2342_
timestamp 1728341909
transform 1 0 10190 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2343_
timestamp 1728341909
transform -1 0 9690 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2345_
timestamp 1728341909
transform -1 0 6970 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2346_
timestamp 1728341909
transform 1 0 6830 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2348_
timestamp 1728341909
transform 1 0 8170 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2350_
timestamp 1728341909
transform 1 0 7590 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2351_
timestamp 1728341909
transform -1 0 5290 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2353_
timestamp 1728341909
transform -1 0 4310 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2354_
timestamp 1728341909
transform 1 0 4790 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2356_
timestamp 1728341909
transform 1 0 5990 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2358_
timestamp 1728341909
transform 1 0 7030 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__2359_
timestamp 1728341909
transform 1 0 6390 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2361_
timestamp 1728341909
transform 1 0 7930 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__2362_
timestamp 1728341909
transform 1 0 7450 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__2364_
timestamp 1728341909
transform 1 0 8170 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__2366_
timestamp 1728341909
transform 1 0 7810 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2367_
timestamp 1728341909
transform 1 0 8090 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2369_
timestamp 1728341909
transform -1 0 10030 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2371_
timestamp 1728341909
transform -1 0 8850 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2372_
timestamp 1728341909
transform -1 0 8590 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2374_
timestamp 1728341909
transform 1 0 8170 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2375_
timestamp 1728341909
transform 1 0 6570 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2377_
timestamp 1728341909
transform -1 0 8790 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2379_
timestamp 1728341909
transform -1 0 6950 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2380_
timestamp 1728341909
transform -1 0 7090 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2382_
timestamp 1728341909
transform -1 0 8030 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2383_
timestamp 1728341909
transform 1 0 7750 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2385_
timestamp 1728341909
transform -1 0 7590 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2387_
timestamp 1728341909
transform -1 0 6470 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2388_
timestamp 1728341909
transform -1 0 9030 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2390_
timestamp 1728341909
transform -1 0 8350 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2392_
timestamp 1728341909
transform 1 0 8350 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2393_
timestamp 1728341909
transform 1 0 8310 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2395_
timestamp 1728341909
transform 1 0 8910 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2396_
timestamp 1728341909
transform 1 0 9190 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2398_
timestamp 1728341909
transform 1 0 8830 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2400_
timestamp 1728341909
transform 1 0 7450 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2401_
timestamp 1728341909
transform 1 0 8570 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2403_
timestamp 1728341909
transform -1 0 6710 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2404_
timestamp 1728341909
transform -1 0 7670 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2406_
timestamp 1728341909
transform 1 0 7170 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2408_
timestamp 1728341909
transform -1 0 6010 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2409_
timestamp 1728341909
transform 1 0 7090 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2411_
timestamp 1728341909
transform -1 0 6930 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2412_
timestamp 1728341909
transform -1 0 7590 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2414_
timestamp 1728341909
transform 1 0 6930 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2416_
timestamp 1728341909
transform 1 0 7870 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2417_
timestamp 1728341909
transform -1 0 9110 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2419_
timestamp 1728341909
transform 1 0 7150 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2421_
timestamp 1728341909
transform -1 0 9770 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__2422_
timestamp 1728341909
transform 1 0 8350 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__2424_
timestamp 1728341909
transform 1 0 8850 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__2425_
timestamp 1728341909
transform 1 0 3250 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2427_
timestamp 1728341909
transform 1 0 8910 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__2429_
timestamp 1728341909
transform 1 0 9530 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__2430_
timestamp 1728341909
transform 1 0 8890 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__2432_
timestamp 1728341909
transform 1 0 9570 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__2433_
timestamp 1728341909
transform -1 0 9990 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__2435_
timestamp 1728341909
transform 1 0 4530 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__2437_
timestamp 1728341909
transform 1 0 10970 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__2438_
timestamp 1728341909
transform -1 0 11030 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__2440_
timestamp 1728341909
transform 1 0 9130 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__2442_
timestamp 1728341909
transform -1 0 8350 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__2443_
timestamp 1728341909
transform 1 0 3910 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__2445_
timestamp 1728341909
transform -1 0 8690 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__2446_
timestamp 1728341909
transform 1 0 8330 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__2448_
timestamp 1728341909
transform 1 0 8570 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__2450_
timestamp 1728341909
transform -1 0 9050 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__2451_
timestamp 1728341909
transform 1 0 3910 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2453_
timestamp 1728341909
transform -1 0 6710 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__2454_
timestamp 1728341909
transform -1 0 6430 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__2456_
timestamp 1728341909
transform -1 0 8830 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__2458_
timestamp 1728341909
transform -1 0 6890 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__2459_
timestamp 1728341909
transform -1 0 3670 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__2461_
timestamp 1728341909
transform 1 0 7110 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__2462_
timestamp 1728341909
transform -1 0 7390 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__2464_
timestamp 1728341909
transform 1 0 4570 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__2466_
timestamp 1728341909
transform -1 0 3450 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2467_
timestamp 1728341909
transform 1 0 6270 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2469_
timestamp 1728341909
transform -1 0 6230 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__2471_
timestamp 1728341909
transform -1 0 8150 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__2472_
timestamp 1728341909
transform -1 0 6170 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__2474_
timestamp 1728341909
transform -1 0 5430 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__2475_
timestamp 1728341909
transform -1 0 7890 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__2477_
timestamp 1728341909
transform -1 0 5290 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2479_
timestamp 1728341909
transform -1 0 8110 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__2480_
timestamp 1728341909
transform 1 0 6010 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2482_
timestamp 1728341909
transform -1 0 2550 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__2483_
timestamp 1728341909
transform -1 0 4790 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__2485_
timestamp 1728341909
transform -1 0 7070 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__2487_
timestamp 1728341909
transform -1 0 5770 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2488_
timestamp 1728341909
transform 1 0 6530 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2490_
timestamp 1728341909
transform 1 0 7790 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2491_
timestamp 1728341909
transform -1 0 8030 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2493_
timestamp 1728341909
transform -1 0 5610 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__2495_
timestamp 1728341909
transform 1 0 6930 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__2496_
timestamp 1728341909
transform 1 0 7650 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__2498_
timestamp 1728341909
transform -1 0 8870 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__2500_
timestamp 1728341909
transform -1 0 7730 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__2501_
timestamp 1728341909
transform -1 0 6850 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__2503_
timestamp 1728341909
transform 1 0 11210 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__2504_
timestamp 1728341909
transform -1 0 4650 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__2506_
timestamp 1728341909
transform -1 0 6810 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__2508_
timestamp 1728341909
transform 1 0 5750 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__2509_
timestamp 1728341909
transform -1 0 8910 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__2511_
timestamp 1728341909
transform -1 0 7490 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__2512_
timestamp 1728341909
transform 1 0 7190 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__2514_
timestamp 1728341909
transform 1 0 7130 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__2516_
timestamp 1728341909
transform 1 0 8610 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__2517_
timestamp 1728341909
transform 1 0 10710 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__2519_
timestamp 1728341909
transform 1 0 10050 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__2521_
timestamp 1728341909
transform -1 0 8610 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__2522_
timestamp 1728341909
transform 1 0 6170 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__2524_
timestamp 1728341909
transform 1 0 8370 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__2525_
timestamp 1728341909
transform 1 0 6870 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__2527_
timestamp 1728341909
transform 1 0 8090 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__2529_
timestamp 1728341909
transform 1 0 7930 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__2530_
timestamp 1728341909
transform -1 0 7890 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__2532_
timestamp 1728341909
transform 1 0 7910 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__2533_
timestamp 1728341909
transform -1 0 5570 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__2535_
timestamp 1728341909
transform -1 0 7670 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__2537_
timestamp 1728341909
transform 1 0 7390 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__2538_
timestamp 1728341909
transform 1 0 8110 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__2540_
timestamp 1728341909
transform 1 0 5690 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__2541_
timestamp 1728341909
transform 1 0 6210 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__2543_
timestamp 1728341909
transform -1 0 6710 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__2545_
timestamp 1728341909
transform 1 0 6950 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__2546_
timestamp 1728341909
transform 1 0 6210 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__2548_
timestamp 1728341909
transform 1 0 7210 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__2550_
timestamp 1728341909
transform -1 0 7630 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__2551_
timestamp 1728341909
transform -1 0 6350 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__2553_
timestamp 1728341909
transform -1 0 5950 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__2554_
timestamp 1728341909
transform -1 0 5670 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__2556_
timestamp 1728341909
transform 1 0 5110 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__2558_
timestamp 1728341909
transform -1 0 6490 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__2559_
timestamp 1728341909
transform 1 0 6170 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__2561_
timestamp 1728341909
transform -1 0 5490 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__2562_
timestamp 1728341909
transform 1 0 5110 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__2564_
timestamp 1728341909
transform -1 0 4670 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__2566_
timestamp 1728341909
transform -1 0 5030 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2567_
timestamp 1728341909
transform 1 0 5230 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__2569_
timestamp 1728341909
transform -1 0 4250 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__2570_
timestamp 1728341909
transform 1 0 5270 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__2572_
timestamp 1728341909
transform -1 0 4510 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__2574_
timestamp 1728341909
transform 1 0 5470 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__2575_
timestamp 1728341909
transform -1 0 5030 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__2577_
timestamp 1728341909
transform 1 0 4950 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__2579_
timestamp 1728341909
transform 1 0 4750 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__2580_
timestamp 1728341909
transform 1 0 4790 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__2582_
timestamp 1728341909
transform -1 0 3370 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__2583_
timestamp 1728341909
transform 1 0 2310 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__2585_
timestamp 1728341909
transform -1 0 6430 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__2587_
timestamp 1728341909
transform -1 0 3530 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__2588_
timestamp 1728341909
transform -1 0 3050 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__2590_
timestamp 1728341909
transform 1 0 3670 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__2591_
timestamp 1728341909
transform -1 0 3150 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__2593_
timestamp 1728341909
transform -1 0 2750 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__2595_
timestamp 1728341909
transform -1 0 3850 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__2596_
timestamp 1728341909
transform 1 0 3450 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__2598_
timestamp 1728341909
transform -1 0 3270 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2600_
timestamp 1728341909
transform 1 0 2990 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__2601_
timestamp 1728341909
transform -1 0 2550 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2603_
timestamp 1728341909
transform -1 0 2410 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__2604_
timestamp 1728341909
transform 1 0 2550 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2606_
timestamp 1728341909
transform 1 0 2270 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2608_
timestamp 1728341909
transform -1 0 1150 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__2609_
timestamp 1728341909
transform 1 0 2110 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__2611_
timestamp 1728341909
transform -1 0 1330 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2612_
timestamp 1728341909
transform -1 0 1070 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2614_
timestamp 1728341909
transform -1 0 670 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__2616_
timestamp 1728341909
transform 1 0 1590 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__2617_
timestamp 1728341909
transform -1 0 1590 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2619_
timestamp 1728341909
transform 1 0 870 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__2620_
timestamp 1728341909
transform -1 0 1390 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__2622_
timestamp 1728341909
transform -1 0 1350 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__2624_
timestamp 1728341909
transform -1 0 630 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2625_
timestamp 1728341909
transform -1 0 2710 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2627_
timestamp 1728341909
transform 1 0 1470 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2629_
timestamp 1728341909
transform -1 0 3470 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__2630_
timestamp 1728341909
transform 1 0 4330 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__2632_
timestamp 1728341909
transform 1 0 10970 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__2633_
timestamp 1728341909
transform 1 0 3970 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__2635_
timestamp 1728341909
transform -1 0 2350 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__2637_
timestamp 1728341909
transform 1 0 4430 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2638_
timestamp 1728341909
transform 1 0 4930 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2640_
timestamp 1728341909
transform -1 0 9950 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__2641_
timestamp 1728341909
transform 1 0 10250 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__2643_
timestamp 1728341909
transform 1 0 10990 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__2645_
timestamp 1728341909
transform -1 0 9790 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__2646_
timestamp 1728341909
transform 1 0 10190 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__2648_
timestamp 1728341909
transform -1 0 4250 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__2650_
timestamp 1728341909
transform 1 0 9390 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__2651_
timestamp 1728341909
transform -1 0 5770 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__2653_
timestamp 1728341909
transform -1 0 7830 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__2654_
timestamp 1728341909
transform 1 0 4750 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__2656_
timestamp 1728341909
transform -1 0 6110 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__2658_
timestamp 1728341909
transform 1 0 6350 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__2659_
timestamp 1728341909
transform 1 0 7050 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__2661_
timestamp 1728341909
transform -1 0 4550 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__2662_
timestamp 1728341909
transform 1 0 4510 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__2664_
timestamp 1728341909
transform -1 0 6690 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2666_
timestamp 1728341909
transform 1 0 6930 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2667_
timestamp 1728341909
transform 1 0 7670 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2669_
timestamp 1728341909
transform 1 0 8070 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__2670_
timestamp 1728341909
transform -1 0 4290 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__2672_
timestamp 1728341909
transform 1 0 5310 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__2674_
timestamp 1728341909
transform -1 0 7490 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2675_
timestamp 1728341909
transform 1 0 7730 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2677_
timestamp 1728341909
transform 1 0 7850 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2679_
timestamp 1728341909
transform 1 0 4250 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__2680_
timestamp 1728341909
transform -1 0 4510 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__2682_
timestamp 1728341909
transform 1 0 6830 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__2683_
timestamp 1728341909
transform 1 0 4170 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2685_
timestamp 1728341909
transform 1 0 5550 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__2687_
timestamp 1728341909
transform 1 0 7430 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2688_
timestamp 1728341909
transform -1 0 7570 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__2690_
timestamp 1728341909
transform 1 0 6670 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2691_
timestamp 1728341909
transform 1 0 7170 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2693_
timestamp 1728341909
transform 1 0 5150 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2695_
timestamp 1728341909
transform 1 0 6730 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2696_
timestamp 1728341909
transform 1 0 6670 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__2698_
timestamp 1728341909
transform 1 0 6990 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2699_
timestamp 1728341909
transform -1 0 6430 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__2701_
timestamp 1728341909
transform -1 0 5570 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__2703_
timestamp 1728341909
transform -1 0 5670 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2704_
timestamp 1728341909
transform 1 0 5730 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2706_
timestamp 1728341909
transform -1 0 6250 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2708_
timestamp 1728341909
transform -1 0 2390 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__2709_
timestamp 1728341909
transform -1 0 5050 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__2711_
timestamp 1728341909
transform -1 0 5170 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__2712_
timestamp 1728341909
transform -1 0 5750 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__2714_
timestamp 1728341909
transform -1 0 6190 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2716_
timestamp 1728341909
transform -1 0 6750 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__2717_
timestamp 1728341909
transform 1 0 6690 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2719_
timestamp 1728341909
transform -1 0 6430 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2720_
timestamp 1728341909
transform 1 0 4730 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__2722_
timestamp 1728341909
transform 1 0 5250 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__2724_
timestamp 1728341909
transform 1 0 6230 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2725_
timestamp 1728341909
transform 1 0 6470 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2727_
timestamp 1728341909
transform 1 0 5930 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__2729_
timestamp 1728341909
transform -1 0 4270 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__2730_
timestamp 1728341909
transform -1 0 5310 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__2732_
timestamp 1728341909
transform -1 0 5730 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2733_
timestamp 1728341909
transform -1 0 5990 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2735_
timestamp 1728341909
transform 1 0 5510 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__2737_
timestamp 1728341909
transform 1 0 3830 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2738_
timestamp 1728341909
transform 1 0 4010 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__2740_
timestamp 1728341909
transform -1 0 3770 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__2741_
timestamp 1728341909
transform -1 0 4110 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2743_
timestamp 1728341909
transform 1 0 4990 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2745_
timestamp 1728341909
transform 1 0 5210 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2746_
timestamp 1728341909
transform 1 0 4710 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2748_
timestamp 1728341909
transform -1 0 5030 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__2749_
timestamp 1728341909
transform -1 0 5390 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__2751_
timestamp 1728341909
transform 1 0 4470 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2753_
timestamp 1728341909
transform -1 0 3510 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2754_
timestamp 1728341909
transform -1 0 3090 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2756_
timestamp 1728341909
transform -1 0 3730 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2758_
timestamp 1728341909
transform -1 0 3730 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2759_
timestamp 1728341909
transform -1 0 3610 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2761_
timestamp 1728341909
transform -1 0 3790 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2762_
timestamp 1728341909
transform -1 0 3550 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__2764_
timestamp 1728341909
transform 1 0 3390 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__2766_
timestamp 1728341909
transform 1 0 3790 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__2767_
timestamp 1728341909
transform -1 0 4490 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__2769_
timestamp 1728341909
transform 1 0 5230 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2770_
timestamp 1728341909
transform -1 0 4730 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2772_
timestamp 1728341909
transform -1 0 4990 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2774_
timestamp 1728341909
transform -1 0 2610 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__2775_
timestamp 1728341909
transform 1 0 3970 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2777_
timestamp 1728341909
transform 1 0 5230 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2778_
timestamp 1728341909
transform -1 0 4730 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2780_
timestamp 1728341909
transform 1 0 2830 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__2782_
timestamp 1728341909
transform -1 0 2850 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__2783_
timestamp 1728341909
transform 1 0 2550 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__2785_
timestamp 1728341909
transform -1 0 2330 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2787_
timestamp 1728341909
transform -1 0 3010 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2788_
timestamp 1728341909
transform -1 0 2510 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__2790_
timestamp 1728341909
transform 1 0 3290 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__2791_
timestamp 1728341909
transform -1 0 3030 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__2793_
timestamp 1728341909
transform -1 0 2350 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__2795_
timestamp 1728341909
transform 1 0 870 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2796_
timestamp 1728341909
transform 1 0 1810 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2798_
timestamp 1728341909
transform 1 0 1310 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2799_
timestamp 1728341909
transform -1 0 1590 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2801_
timestamp 1728341909
transform 1 0 1810 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2803_
timestamp 1728341909
transform 1 0 3370 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2804_
timestamp 1728341909
transform -1 0 530 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__2806_
timestamp 1728341909
transform -1 0 5490 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2808_
timestamp 1728341909
transform 1 0 4010 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2809_
timestamp 1728341909
transform -1 0 4470 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2811_
timestamp 1728341909
transform -1 0 4690 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2812_
timestamp 1728341909
transform 1 0 4310 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__2814_
timestamp 1728341909
transform 1 0 4190 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__2816_
timestamp 1728341909
transform 1 0 2570 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__2817_
timestamp 1728341909
transform -1 0 2850 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__2819_
timestamp 1728341909
transform 1 0 3250 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2820_
timestamp 1728341909
transform 1 0 3490 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2822_
timestamp 1728341909
transform -1 0 4830 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__2824_
timestamp 1728341909
transform 1 0 630 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__2825_
timestamp 1728341909
transform 1 0 610 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2827_
timestamp 1728341909
transform 1 0 1810 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__2828_
timestamp 1728341909
transform -1 0 2090 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__2830_
timestamp 1728341909
transform -1 0 1590 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__2832_
timestamp 1728341909
transform 1 0 2110 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2833_
timestamp 1728341909
transform -1 0 1130 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__2835_
timestamp 1728341909
transform 1 0 1190 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__2837_
timestamp 1728341909
transform 1 0 1730 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__2838_
timestamp 1728341909
transform -1 0 1610 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__2840_
timestamp 1728341909
transform 1 0 1330 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__2841_
timestamp 1728341909
transform 1 0 2130 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__2843_
timestamp 1728341909
transform -1 0 1890 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__2845_
timestamp 1728341909
transform -1 0 1590 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__2846_
timestamp 1728341909
transform 1 0 1370 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2848_
timestamp 1728341909
transform -1 0 1350 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__2849_
timestamp 1728341909
transform -1 0 1650 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2851_
timestamp 1728341909
transform -1 0 1110 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__2853_
timestamp 1728341909
transform -1 0 2370 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2854_
timestamp 1728341909
transform 1 0 850 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__2856_
timestamp 1728341909
transform -1 0 2050 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__2857_
timestamp 1728341909
transform -1 0 2450 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__2859_
timestamp 1728341909
transform -1 0 930 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2861_
timestamp 1728341909
transform -1 0 170 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__2862_
timestamp 1728341909
transform -1 0 1130 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__2864_
timestamp 1728341909
transform -1 0 410 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__2866_
timestamp 1728341909
transform 1 0 4550 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__2867_
timestamp 1728341909
transform 1 0 5650 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__2869_
timestamp 1728341909
transform -1 0 3310 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__2870_
timestamp 1728341909
transform -1 0 2370 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__2872_
timestamp 1728341909
transform -1 0 4670 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__2874_
timestamp 1728341909
transform -1 0 4210 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2875_
timestamp 1728341909
transform -1 0 1770 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2877_
timestamp 1728341909
transform -1 0 3570 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2878_
timestamp 1728341909
transform -1 0 4010 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__2880_
timestamp 1728341909
transform 1 0 1530 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__2882_
timestamp 1728341909
transform -1 0 2530 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__2883_
timestamp 1728341909
transform 1 0 4530 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__2885_
timestamp 1728341909
transform 1 0 3190 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2887_
timestamp 1728341909
transform 1 0 5210 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2888_
timestamp 1728341909
transform 1 0 3470 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2890_
timestamp 1728341909
transform -1 0 4470 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2891_
timestamp 1728341909
transform -1 0 4210 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__2893_
timestamp 1728341909
transform 1 0 3750 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2895_
timestamp 1728341909
transform 1 0 4530 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2896_
timestamp 1728341909
transform -1 0 3930 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2898_
timestamp 1728341909
transform 1 0 5250 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2899_
timestamp 1728341909
transform 1 0 5210 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2901_
timestamp 1728341909
transform -1 0 4950 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2903_
timestamp 1728341909
transform 1 0 2270 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2904_
timestamp 1728341909
transform 1 0 2530 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2906_
timestamp 1728341909
transform 1 0 1110 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2907_
timestamp 1728341909
transform 1 0 1310 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2909_
timestamp 1728341909
transform -1 0 1850 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2911_
timestamp 1728341909
transform -1 0 1630 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2912_
timestamp 1728341909
transform -1 0 2550 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2914_
timestamp 1728341909
transform 1 0 2310 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2916_
timestamp 1728341909
transform 1 0 1770 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2917_
timestamp 1728341909
transform -1 0 1850 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2919_
timestamp 1728341909
transform -1 0 2330 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2920_
timestamp 1728341909
transform -1 0 2050 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__2922_
timestamp 1728341909
transform -1 0 2030 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__2924_
timestamp 1728341909
transform -1 0 3030 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2925_
timestamp 1728341909
transform 1 0 3510 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2927_
timestamp 1728341909
transform -1 0 2530 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__2928_
timestamp 1728341909
transform 1 0 4670 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__2930_
timestamp 1728341909
transform -1 0 2790 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2932_
timestamp 1728341909
transform 1 0 3230 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2933_
timestamp 1728341909
transform -1 0 2790 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2935_
timestamp 1728341909
transform -1 0 1390 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2937_
timestamp 1728341909
transform 1 0 650 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2938_
timestamp 1728341909
transform 1 0 1810 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2940_
timestamp 1728341909
transform 1 0 3250 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2941_
timestamp 1728341909
transform 1 0 3250 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2943_
timestamp 1728341909
transform -1 0 3310 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2945_
timestamp 1728341909
transform 1 0 3250 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__2946_
timestamp 1728341909
transform 1 0 3690 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__2948_
timestamp 1728341909
transform -1 0 4270 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__2949_
timestamp 1728341909
transform 1 0 3230 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__2951_
timestamp 1728341909
transform -1 0 2790 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2953_
timestamp 1728341909
transform -1 0 2270 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__2954_
timestamp 1728341909
transform -1 0 2510 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__2956_
timestamp 1728341909
transform 1 0 3330 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__2957_
timestamp 1728341909
transform 1 0 3830 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__2959_
timestamp 1728341909
transform 1 0 3550 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__2961_
timestamp 1728341909
transform 1 0 2790 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2962_
timestamp 1728341909
transform 1 0 2530 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2964_
timestamp 1728341909
transform 1 0 2790 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2966_
timestamp 1728341909
transform 1 0 4190 0 1 1690
box -12 -8 32 252
use FILL  FILL_7__2967_
timestamp 1728341909
transform -1 0 4670 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2969_
timestamp 1728341909
transform -1 0 1410 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__2970_
timestamp 1728341909
transform -1 0 1590 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__2972_
timestamp 1728341909
transform -1 0 1350 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__2974_
timestamp 1728341909
transform -1 0 1850 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2975_
timestamp 1728341909
transform -1 0 2070 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2977_
timestamp 1728341909
transform -1 0 4510 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2978_
timestamp 1728341909
transform 1 0 4230 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2980_
timestamp 1728341909
transform -1 0 1090 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2982_
timestamp 1728341909
transform 1 0 2290 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__2983_
timestamp 1728341909
transform -1 0 610 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2985_
timestamp 1728341909
transform -1 0 170 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__2986_
timestamp 1728341909
transform -1 0 430 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2988_
timestamp 1728341909
transform -1 0 650 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2990_
timestamp 1728341909
transform 1 0 150 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__2991_
timestamp 1728341909
transform -1 0 430 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2993_
timestamp 1728341909
transform -1 0 1130 0 1 730
box -12 -8 32 252
use FILL  FILL_7__2995_
timestamp 1728341909
transform 1 0 670 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__2996_
timestamp 1728341909
transform -1 0 610 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__2998_
timestamp 1728341909
transform -1 0 170 0 1 250
box -12 -8 32 252
use FILL  FILL_7__2999_
timestamp 1728341909
transform -1 0 410 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__3001_
timestamp 1728341909
transform -1 0 170 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7__3003_
timestamp 1728341909
transform -1 0 170 0 1 730
box -12 -8 32 252
use FILL  FILL_7__3004_
timestamp 1728341909
transform -1 0 910 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__3006_
timestamp 1728341909
transform -1 0 170 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__3007_
timestamp 1728341909
transform 1 0 1870 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__3009_
timestamp 1728341909
transform -1 0 1390 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__3011_
timestamp 1728341909
transform -1 0 1150 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7__3012_
timestamp 1728341909
transform -1 0 1530 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__3014_
timestamp 1728341909
transform 1 0 1110 0 1 250
box -12 -8 32 252
use FILL  FILL_7__3016_
timestamp 1728341909
transform -1 0 1370 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__3017_
timestamp 1728341909
transform -1 0 1350 0 1 250
box -12 -8 32 252
use FILL  FILL_7__3019_
timestamp 1728341909
transform -1 0 1130 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7__3020_
timestamp 1728341909
transform -1 0 3770 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__3022_
timestamp 1728341909
transform 1 0 2870 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3024_
timestamp 1728341909
transform 1 0 3870 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__3025_
timestamp 1728341909
transform -1 0 4290 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__3027_
timestamp 1728341909
transform -1 0 3550 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__3028_
timestamp 1728341909
transform -1 0 4070 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3030_
timestamp 1728341909
transform 1 0 3550 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__3032_
timestamp 1728341909
transform -1 0 2630 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3033_
timestamp 1728341909
transform -1 0 2650 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__3035_
timestamp 1728341909
transform -1 0 3050 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__3036_
timestamp 1728341909
transform 1 0 3370 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__3038_
timestamp 1728341909
transform -1 0 3370 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3040_
timestamp 1728341909
transform 1 0 2250 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__3041_
timestamp 1728341909
transform 1 0 2790 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__3043_
timestamp 1728341909
transform 1 0 6390 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__3045_
timestamp 1728341909
transform 1 0 5830 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__3046_
timestamp 1728341909
transform 1 0 5550 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__3048_
timestamp 1728341909
transform 1 0 5230 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__3049_
timestamp 1728341909
transform 1 0 5930 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3051_
timestamp 1728341909
transform -1 0 6410 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__3053_
timestamp 1728341909
transform 1 0 6190 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__3054_
timestamp 1728341909
transform 1 0 5930 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__3056_
timestamp 1728341909
transform 1 0 4690 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__3057_
timestamp 1728341909
transform 1 0 4450 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__3059_
timestamp 1728341909
transform 1 0 4390 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__3061_
timestamp 1728341909
transform 1 0 4070 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__3062_
timestamp 1728341909
transform -1 0 4890 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__3064_
timestamp 1728341909
transform 1 0 6090 0 1 2170
box -12 -8 32 252
use FILL  FILL_7__3065_
timestamp 1728341909
transform 1 0 5870 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7__3067_
timestamp 1728341909
transform -1 0 6010 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__3069_
timestamp 1728341909
transform -1 0 6550 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__3070_
timestamp 1728341909
transform 1 0 6190 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3072_
timestamp 1728341909
transform 1 0 6670 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__3074_
timestamp 1728341909
transform 1 0 490 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__3075_
timestamp 1728341909
transform -1 0 650 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__3077_
timestamp 1728341909
transform 1 0 2090 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__3078_
timestamp 1728341909
transform -1 0 5590 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__3080_
timestamp 1728341909
transform 1 0 4330 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__3082_
timestamp 1728341909
transform -1 0 6970 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__3083_
timestamp 1728341909
transform 1 0 6130 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__3085_
timestamp 1728341909
transform -1 0 5090 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__3086_
timestamp 1728341909
transform 1 0 5570 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__3088_
timestamp 1728341909
transform -1 0 5710 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__3090_
timestamp 1728341909
transform 1 0 4850 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__3091_
timestamp 1728341909
transform -1 0 4810 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__3093_
timestamp 1728341909
transform -1 0 4070 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__3095_
timestamp 1728341909
transform 1 0 4810 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__3096_
timestamp 1728341909
transform 1 0 4790 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__3098_
timestamp 1728341909
transform -1 0 5130 0 1 2650
box -12 -8 32 252
use FILL  FILL_7__3099_
timestamp 1728341909
transform 1 0 5270 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7__3101_
timestamp 1728341909
transform 1 0 5210 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__3103_
timestamp 1728341909
transform 1 0 4950 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__3104_
timestamp 1728341909
transform -1 0 5090 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__3106_
timestamp 1728341909
transform 1 0 8590 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__3107_
timestamp 1728341909
transform 1 0 8350 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__3109_
timestamp 1728341909
transform -1 0 8650 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__3111_
timestamp 1728341909
transform 1 0 4590 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__3112_
timestamp 1728341909
transform 1 0 4830 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__3114_
timestamp 1728341909
transform 1 0 850 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__3115_
timestamp 1728341909
transform 1 0 4530 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__3117_
timestamp 1728341909
transform -1 0 410 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__3119_
timestamp 1728341909
transform -1 0 5010 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__3120_
timestamp 1728341909
transform 1 0 4510 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3122_
timestamp 1728341909
transform -1 0 4550 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__3124_
timestamp 1728341909
transform -1 0 4030 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3125_
timestamp 1728341909
transform -1 0 3770 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3127_
timestamp 1728341909
transform 1 0 4810 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__3128_
timestamp 1728341909
transform 1 0 4730 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__3130_
timestamp 1728341909
transform -1 0 1910 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3132_
timestamp 1728341909
transform 1 0 1130 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__3133_
timestamp 1728341909
transform 1 0 3990 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__3135_
timestamp 1728341909
transform 1 0 3310 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__3136_
timestamp 1728341909
transform 1 0 3790 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3138_
timestamp 1728341909
transform -1 0 4090 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__3140_
timestamp 1728341909
transform 1 0 890 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__3141_
timestamp 1728341909
transform -1 0 4070 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__3143_
timestamp 1728341909
transform -1 0 4270 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3145_
timestamp 1728341909
transform 1 0 3290 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3146_
timestamp 1728341909
transform -1 0 3370 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__3148_
timestamp 1728341909
transform -1 0 3570 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3149_
timestamp 1728341909
transform -1 0 3550 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__3151_
timestamp 1728341909
transform -1 0 2370 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__3153_
timestamp 1728341909
transform 1 0 4530 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3154_
timestamp 1728341909
transform -1 0 870 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__3156_
timestamp 1728341909
transform 1 0 3050 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3157_
timestamp 1728341909
transform -1 0 2830 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__3159_
timestamp 1728341909
transform 1 0 2590 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__3161_
timestamp 1728341909
transform -1 0 2750 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__3162_
timestamp 1728341909
transform -1 0 2530 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__3164_
timestamp 1728341909
transform 1 0 1330 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__3165_
timestamp 1728341909
transform -1 0 410 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__3167_
timestamp 1728341909
transform 1 0 2130 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3169_
timestamp 1728341909
transform -1 0 2370 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__3170_
timestamp 1728341909
transform 1 0 2110 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__3172_
timestamp 1728341909
transform 1 0 1970 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__3174_
timestamp 1728341909
transform -1 0 1870 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__3175_
timestamp 1728341909
transform -1 0 3110 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__3177_
timestamp 1728341909
transform 1 0 2350 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3178_
timestamp 1728341909
transform 1 0 2690 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3180_
timestamp 1728341909
transform 1 0 3290 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3182_
timestamp 1728341909
transform -1 0 3090 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__3183_
timestamp 1728341909
transform 1 0 2850 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__3185_
timestamp 1728341909
transform -1 0 2610 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__3186_
timestamp 1728341909
transform 1 0 2090 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__3188_
timestamp 1728341909
transform -1 0 170 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__3190_
timestamp 1728341909
transform -1 0 910 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3191_
timestamp 1728341909
transform -1 0 1170 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3193_
timestamp 1728341909
transform 1 0 1530 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__3194_
timestamp 1728341909
transform 1 0 3330 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__3196_
timestamp 1728341909
transform 1 0 2030 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__3198_
timestamp 1728341909
transform -1 0 2190 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3199_
timestamp 1728341909
transform -1 0 2450 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3201_
timestamp 1728341909
transform -1 0 1130 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__3203_
timestamp 1728341909
transform -1 0 1390 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3204_
timestamp 1728341909
transform -1 0 650 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3206_
timestamp 1728341909
transform 1 0 1150 0 -1 4090
box -12 -8 32 252
use FILL  FILL_7__3207_
timestamp 1728341909
transform -1 0 410 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__3209_
timestamp 1728341909
transform 1 0 390 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__3211_
timestamp 1728341909
transform -1 0 1650 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__3212_
timestamp 1728341909
transform -1 0 1390 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__3214_
timestamp 1728341909
transform 1 0 1410 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3215_
timestamp 1728341909
transform -1 0 1370 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__3217_
timestamp 1728341909
transform -1 0 410 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__3219_
timestamp 1728341909
transform -1 0 1690 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3220_
timestamp 1728341909
transform 1 0 1910 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3222_
timestamp 1728341909
transform -1 0 170 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3224_
timestamp 1728341909
transform 1 0 630 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__3225_
timestamp 1728341909
transform -1 0 410 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__3227_
timestamp 1728341909
transform -1 0 430 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__3228_
timestamp 1728341909
transform -1 0 170 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__3230_
timestamp 1728341909
transform 1 0 1810 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__3232_
timestamp 1728341909
transform -1 0 1870 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__3233_
timestamp 1728341909
transform 1 0 1170 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3235_
timestamp 1728341909
transform 1 0 1130 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__3236_
timestamp 1728341909
transform 1 0 1390 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__3238_
timestamp 1728341909
transform 1 0 2550 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7__3240_
timestamp 1728341909
transform -1 0 890 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__3241_
timestamp 1728341909
transform 1 0 9790 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__3243_
timestamp 1728341909
transform 1 0 9550 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__3244_
timestamp 1728341909
transform 1 0 8850 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__3246_
timestamp 1728341909
transform -1 0 9670 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__3248_
timestamp 1728341909
transform 1 0 10830 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__3249_
timestamp 1728341909
transform -1 0 9570 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__3251_
timestamp 1728341909
transform 1 0 9330 0 1 3130
box -12 -8 32 252
use FILL  FILL_7__3253_
timestamp 1728341909
transform -1 0 7970 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__3254_
timestamp 1728341909
transform -1 0 8230 0 1 3610
box -12 -8 32 252
use FILL  FILL_7__3256_
timestamp 1728341909
transform 1 0 8350 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3257_
timestamp 1728341909
transform 1 0 8110 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3259_
timestamp 1728341909
transform 1 0 9590 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__3261_
timestamp 1728341909
transform -1 0 10490 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__3262_
timestamp 1728341909
transform 1 0 10070 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__3264_
timestamp 1728341909
transform 1 0 9090 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7__3265_
timestamp 1728341909
transform -1 0 9830 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3267_
timestamp 1728341909
transform -1 0 9750 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__3269_
timestamp 1728341909
transform -1 0 10590 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__3270_
timestamp 1728341909
transform 1 0 10310 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3272_
timestamp 1728341909
transform 1 0 10350 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7__3273_
timestamp 1728341909
transform -1 0 10250 0 1 4570
box -12 -8 32 252
use FILL  FILL_7__3275_
timestamp 1728341909
transform 1 0 9670 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__3277_
timestamp 1728341909
transform -1 0 10750 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__3278_
timestamp 1728341909
transform 1 0 10210 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__3280_
timestamp 1728341909
transform 1 0 9330 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__3282_
timestamp 1728341909
transform -1 0 6970 0 1 4090
box -12 -8 32 252
use FILL  FILL_7__3283_
timestamp 1728341909
transform -1 0 6910 0 -1 5050
box -12 -8 32 252
use FILL  FILL_7__3285_
timestamp 1728341909
transform 1 0 7110 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3286_
timestamp 1728341909
transform -1 0 7370 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3288_
timestamp 1728341909
transform -1 0 6950 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3290_
timestamp 1728341909
transform 1 0 6630 0 1 5530
box -12 -8 32 252
use FILL  FILL_7__3291_
timestamp 1728341909
transform 1 0 7130 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__3293_
timestamp 1728341909
transform 1 0 7230 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__3294_
timestamp 1728341909
transform 1 0 6970 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__3296_
timestamp 1728341909
transform 1 0 5910 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__3298_
timestamp 1728341909
transform 1 0 5270 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__3299_
timestamp 1728341909
transform 1 0 5710 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3301_
timestamp 1728341909
transform 1 0 6970 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7__3303_
timestamp 1728341909
transform -1 0 3110 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__3304_
timestamp 1728341909
transform 1 0 2050 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__3306_
timestamp 1728341909
transform 1 0 3970 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__3307_
timestamp 1728341909
transform -1 0 4910 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__3309_
timestamp 1728341909
transform -1 0 170 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__3311_
timestamp 1728341909
transform -1 0 890 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__3312_
timestamp 1728341909
transform -1 0 390 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__3314_
timestamp 1728341909
transform -1 0 170 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__3315_
timestamp 1728341909
transform -1 0 170 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__3317_
timestamp 1728341909
transform -1 0 890 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__3450_
timestamp 1728341909
transform 1 0 3070 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__3451_
timestamp 1728341909
transform 1 0 3190 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__3453_
timestamp 1728341909
transform 1 0 3310 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__3454_
timestamp 1728341909
transform -1 0 3670 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__3456_
timestamp 1728341909
transform 1 0 9610 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__3458_
timestamp 1728341909
transform -1 0 10050 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3459_
timestamp 1728341909
transform 1 0 10490 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3461_
timestamp 1728341909
transform -1 0 10550 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__3463_
timestamp 1728341909
transform 1 0 10510 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7__3464_
timestamp 1728341909
transform -1 0 10310 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__3466_
timestamp 1728341909
transform -1 0 10290 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__3467_
timestamp 1728341909
transform 1 0 8350 0 1 6010
box -12 -8 32 252
use FILL  FILL_7__3469_
timestamp 1728341909
transform 1 0 8650 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3471_
timestamp 1728341909
transform 1 0 8730 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__3472_
timestamp 1728341909
transform 1 0 8970 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__3474_
timestamp 1728341909
transform -1 0 8910 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__3475_
timestamp 1728341909
transform -1 0 9030 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__3477_
timestamp 1728341909
transform 1 0 9270 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__3479_
timestamp 1728341909
transform 1 0 10630 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__3480_
timestamp 1728341909
transform -1 0 10190 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__3482_
timestamp 1728341909
transform -1 0 9850 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__3484_
timestamp 1728341909
transform 1 0 10970 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__3485_
timestamp 1728341909
transform 1 0 11250 0 1 6490
box -12 -8 32 252
use FILL  FILL_7__3487_
timestamp 1728341909
transform 1 0 10970 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3488_
timestamp 1728341909
transform 1 0 9610 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__3490_
timestamp 1728341909
transform -1 0 9770 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__3492_
timestamp 1728341909
transform 1 0 9990 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__3493_
timestamp 1728341909
transform 1 0 10250 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__3495_
timestamp 1728341909
transform -1 0 8890 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__3496_
timestamp 1728341909
transform 1 0 9510 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__3498_
timestamp 1728341909
transform 1 0 9890 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__3500_
timestamp 1728341909
transform -1 0 9570 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__3501_
timestamp 1728341909
transform -1 0 9810 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__3503_
timestamp 1728341909
transform 1 0 10130 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__3504_
timestamp 1728341909
transform -1 0 10090 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__3506_
timestamp 1728341909
transform 1 0 10850 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__3508_
timestamp 1728341909
transform -1 0 8590 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__3509_
timestamp 1728341909
transform 1 0 8510 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__3511_
timestamp 1728341909
transform -1 0 9050 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__3513_
timestamp 1728341909
transform -1 0 9070 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__3514_
timestamp 1728341909
transform -1 0 8830 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__3516_
timestamp 1728341909
transform 1 0 11070 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__3517_
timestamp 1728341909
transform -1 0 10390 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__3519_
timestamp 1728341909
transform 1 0 10950 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__3521_
timestamp 1728341909
transform 1 0 7570 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__3522_
timestamp 1728341909
transform -1 0 8090 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__3524_
timestamp 1728341909
transform 1 0 8610 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__3525_
timestamp 1728341909
transform 1 0 9030 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__3527_
timestamp 1728341909
transform -1 0 8370 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__3529_
timestamp 1728341909
transform 1 0 10110 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__3530_
timestamp 1728341909
transform 1 0 10210 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__3532_
timestamp 1728341909
transform 1 0 10390 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__3533_
timestamp 1728341909
transform -1 0 8310 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__3535_
timestamp 1728341909
transform -1 0 8130 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__3537_
timestamp 1728341909
transform 1 0 8450 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__3538_
timestamp 1728341909
transform -1 0 8730 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__3540_
timestamp 1728341909
transform 1 0 9850 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__3542_
timestamp 1728341909
transform -1 0 7590 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__3543_
timestamp 1728341909
transform -1 0 7850 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__3545_
timestamp 1728341909
transform 1 0 8930 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__3546_
timestamp 1728341909
transform -1 0 8370 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__3548_
timestamp 1728341909
transform -1 0 9050 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__3550_
timestamp 1728341909
transform 1 0 8990 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__3551_
timestamp 1728341909
transform 1 0 9270 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__3553_
timestamp 1728341909
transform 1 0 9150 0 -1 9850
box -12 -8 32 252
use FILL  FILL_7__3554_
timestamp 1728341909
transform 1 0 9070 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__3556_
timestamp 1728341909
transform 1 0 8550 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__3558_
timestamp 1728341909
transform -1 0 7850 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__3559_
timestamp 1728341909
transform 1 0 7810 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__3561_
timestamp 1728341909
transform -1 0 8070 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__3563_
timestamp 1728341909
transform -1 0 9050 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__3564_
timestamp 1728341909
transform 1 0 10150 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__3566_
timestamp 1728341909
transform 1 0 9990 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__3567_
timestamp 1728341909
transform 1 0 10070 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__3569_
timestamp 1728341909
transform 1 0 10290 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__3571_
timestamp 1728341909
transform -1 0 10730 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__3572_
timestamp 1728341909
transform -1 0 11230 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__3574_
timestamp 1728341909
transform 1 0 10850 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__3575_
timestamp 1728341909
transform 1 0 11250 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__3577_
timestamp 1728341909
transform -1 0 11270 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__3579_
timestamp 1728341909
transform -1 0 10570 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__3580_
timestamp 1728341909
transform -1 0 9270 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__3582_
timestamp 1728341909
transform 1 0 8810 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__3583_
timestamp 1728341909
transform -1 0 9130 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__3585_
timestamp 1728341909
transform -1 0 9610 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__3587_
timestamp 1728341909
transform -1 0 9330 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__3588_
timestamp 1728341909
transform 1 0 9350 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__3590_
timestamp 1728341909
transform -1 0 10330 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__3592_
timestamp 1728341909
transform 1 0 9830 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__3593_
timestamp 1728341909
transform -1 0 9610 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__3595_
timestamp 1728341909
transform 1 0 11010 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__3596_
timestamp 1728341909
transform -1 0 10970 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__3598_
timestamp 1728341909
transform 1 0 11250 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__3600_
timestamp 1728341909
transform 1 0 11090 0 -1 9370
box -12 -8 32 252
use FILL  FILL_7__3601_
timestamp 1728341909
transform 1 0 10270 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__3603_
timestamp 1728341909
transform 1 0 10570 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__3604_
timestamp 1728341909
transform 1 0 10790 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__3606_
timestamp 1728341909
transform 1 0 10750 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__3608_
timestamp 1728341909
transform -1 0 10290 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__3609_
timestamp 1728341909
transform 1 0 10790 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__3611_
timestamp 1728341909
transform 1 0 9410 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__3612_
timestamp 1728341909
transform 1 0 9670 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__3614_
timestamp 1728341909
transform -1 0 9930 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__3616_
timestamp 1728341909
transform -1 0 9110 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__3617_
timestamp 1728341909
transform -1 0 9370 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__3619_
timestamp 1728341909
transform 1 0 11010 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__3621_
timestamp 1728341909
transform -1 0 10530 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__3622_
timestamp 1728341909
transform 1 0 10770 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__3624_
timestamp 1728341909
transform 1 0 10790 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__3625_
timestamp 1728341909
transform 1 0 10890 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__3627_
timestamp 1728341909
transform -1 0 9770 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__3629_
timestamp 1728341909
transform 1 0 10730 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__3630_
timestamp 1728341909
transform 1 0 10530 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__3632_
timestamp 1728341909
transform -1 0 11030 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__3633_
timestamp 1728341909
transform 1 0 10990 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__3635_
timestamp 1728341909
transform -1 0 10530 0 1 10810
box -12 -8 32 252
use FILL  FILL_7__3637_
timestamp 1728341909
transform -1 0 10790 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__3638_
timestamp 1728341909
transform -1 0 10710 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__3640_
timestamp 1728341909
transform -1 0 11010 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__3642_
timestamp 1728341909
transform -1 0 11070 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__3643_
timestamp 1728341909
transform 1 0 10990 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__3645_
timestamp 1728341909
transform -1 0 10290 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__3646_
timestamp 1728341909
transform -1 0 11050 0 -1 8890
box -12 -8 32 252
use FILL  FILL_7__3648_
timestamp 1728341909
transform 1 0 11230 0 1 8410
box -12 -8 32 252
use FILL  FILL_7__3650_
timestamp 1728341909
transform 1 0 10430 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__3651_
timestamp 1728341909
transform 1 0 10530 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__3653_
timestamp 1728341909
transform 1 0 10710 0 -1 6970
box -12 -8 32 252
use FILL  FILL_7__3654_
timestamp 1728341909
transform 1 0 8510 0 1 9850
box -12 -8 32 252
use FILL  FILL_7__3656_
timestamp 1728341909
transform 1 0 8350 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__3658_
timestamp 1728341909
transform -1 0 8630 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__3659_
timestamp 1728341909
transform -1 0 8370 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7__3661_
timestamp 1728341909
transform -1 0 9350 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__3662_
timestamp 1728341909
transform -1 0 9590 0 1 10330
box -12 -8 32 252
use FILL  FILL_7__3664_
timestamp 1728341909
transform -1 0 9750 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__3666_
timestamp 1728341909
transform -1 0 8590 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__3667_
timestamp 1728341909
transform -1 0 9310 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7__3669_
timestamp 1728341909
transform -1 0 10270 0 1 9370
box -12 -8 32 252
use FILL  FILL_7__3671_
timestamp 1728341909
transform 1 0 8390 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__3672_
timestamp 1728341909
transform 1 0 8630 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__3674_
timestamp 1728341909
transform -1 0 10010 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__3675_
timestamp 1728341909
transform 1 0 10230 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__3677_
timestamp 1728341909
transform 1 0 9510 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__3691_
timestamp 1728341909
transform 1 0 7830 0 1 250
box -12 -8 32 252
use FILL  FILL_7__3692_
timestamp 1728341909
transform -1 0 8090 0 1 250
box -12 -8 32 252
use FILL  FILL_7__3694_
timestamp 1728341909
transform -1 0 170 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__3695_
timestamp 1728341909
transform 1 0 670 0 -1 10330
box -12 -8 32 252
use FILL  FILL_7__3697_
timestamp 1728341909
transform -1 0 170 0 -1 10810
box -12 -8 32 252
use FILL  FILL_7__3699_
timestamp 1728341909
transform 1 0 6230 0 1 1210
box -12 -8 32 252
use FILL  FILL_7__3700_
timestamp 1728341909
transform -1 0 6390 0 -1 730
box -12 -8 32 252
use FILL  FILL_7__3702_
timestamp 1728341909
transform -1 0 5350 0 1 5050
box -12 -8 32 252
use FILL  FILL_7__3703_
timestamp 1728341909
transform -1 0 3590 0 -1 250
box -12 -8 32 252
use FILL  FILL_7__3705_
timestamp 1728341909
transform -1 0 170 0 1 8890
box -12 -8 32 252
use FILL  FILL_7__3707_
timestamp 1728341909
transform 1 0 11230 0 1 6970
box -12 -8 32 252
use FILL  FILL_7__3708_
timestamp 1728341909
transform 1 0 11230 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7__3710_
timestamp 1728341909
transform 1 0 11010 0 1 7450
box -12 -8 32 252
use FILL  FILL_7__3712_
timestamp 1728341909
transform 1 0 11010 0 -1 8410
box -12 -8 32 252
use FILL  FILL_7__3713_
timestamp 1728341909
transform 1 0 11130 0 1 7930
box -12 -8 32 252
use FILL  FILL_7__3715_
timestamp 1728341909
transform 1 0 11230 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert0
timestamp 1728341909
transform 1 0 7870 0 1 10810
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert1
timestamp 1728341909
transform 1 0 9090 0 1 1690
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert3
timestamp 1728341909
transform 1 0 5770 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert4
timestamp 1728341909
transform 1 0 6870 0 1 1690
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert6
timestamp 1728341909
transform 1 0 7290 0 1 10330
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert8
timestamp 1728341909
transform -1 0 7650 0 -1 2170
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert9
timestamp 1728341909
transform 1 0 4570 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert11
timestamp 1728341909
transform -1 0 4890 0 1 2650
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert13
timestamp 1728341909
transform -1 0 5990 0 1 7450
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert14
timestamp 1728341909
transform 1 0 4630 0 1 2650
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert16
timestamp 1728341909
transform 1 0 2790 0 1 8410
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert17
timestamp 1728341909
transform 1 0 4290 0 1 6490
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert19
timestamp 1728341909
transform -1 0 430 0 1 8410
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert21
timestamp 1728341909
transform -1 0 7170 0 1 4570
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert22
timestamp 1728341909
transform -1 0 10550 0 1 4090
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert24
timestamp 1728341909
transform 1 0 8610 0 1 3130
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert25
timestamp 1728341909
transform -1 0 7170 0 1 3130
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert37
timestamp 1728341909
transform -1 0 1090 0 1 5530
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert38
timestamp 1728341909
transform 1 0 1370 0 1 4570
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert40
timestamp 1728341909
transform -1 0 2830 0 -1 6010
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert42
timestamp 1728341909
transform 1 0 8950 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert43
timestamp 1728341909
transform -1 0 8870 0 -1 3610
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert45
timestamp 1728341909
transform 1 0 3950 0 1 4090
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert46
timestamp 1728341909
transform 1 0 5310 0 1 4090
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert48
timestamp 1728341909
transform 1 0 5530 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert50
timestamp 1728341909
transform 1 0 8410 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert51
timestamp 1728341909
transform -1 0 10510 0 1 4570
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert53
timestamp 1728341909
transform -1 0 9630 0 -1 2650
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert54
timestamp 1728341909
transform -1 0 8470 0 -1 3130
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert56
timestamp 1728341909
transform 1 0 5110 0 -1 1210
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert58
timestamp 1728341909
transform 1 0 2030 0 1 1690
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert59
timestamp 1728341909
transform 1 0 4470 0 1 730
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert61
timestamp 1728341909
transform 1 0 10250 0 -1 7450
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert63
timestamp 1728341909
transform 1 0 9370 0 1 7450
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert64
timestamp 1728341909
transform 1 0 8710 0 1 1210
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert66
timestamp 1728341909
transform 1 0 5850 0 1 2650
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert67
timestamp 1728341909
transform 1 0 6690 0 1 5050
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert69
timestamp 1728341909
transform -1 0 6170 0 1 1690
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert71
timestamp 1728341909
transform 1 0 2550 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert72
timestamp 1728341909
transform 1 0 3990 0 1 1210
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert74
timestamp 1728341909
transform -1 0 3790 0 -1 1690
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert75
timestamp 1728341909
transform -1 0 870 0 1 2170
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert77
timestamp 1728341909
transform -1 0 8590 0 -1 5530
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert79
timestamp 1728341909
transform -1 0 9310 0 1 4570
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert80
timestamp 1728341909
transform 1 0 4290 0 -1 6490
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert82
timestamp 1728341909
transform 1 0 2290 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7_BUFX2_insert83
timestamp 1728341909
transform -1 0 2770 0 -1 7930
box -12 -8 32 252
use FILL  FILL_7_CLKBUF1_insert27
timestamp 1728341909
transform 1 0 3750 0 1 3130
box -12 -8 32 252
use FILL  FILL_7_CLKBUF1_insert29
timestamp 1728341909
transform 1 0 630 0 1 7930
box -12 -8 32 252
use FILL  FILL_7_CLKBUF1_insert30
timestamp 1728341909
transform 1 0 8310 0 1 5530
box -12 -8 32 252
use FILL  FILL_7_CLKBUF1_insert32
timestamp 1728341909
transform -1 0 3290 0 -1 4570
box -12 -8 32 252
use FILL  FILL_7_CLKBUF1_insert34
timestamp 1728341909
transform -1 0 170 0 -1 11290
box -12 -8 32 252
use FILL  FILL_7_CLKBUF1_insert35
timestamp 1728341909
transform -1 0 5590 0 1 5050
box -12 -8 32 252
<< labels >>
flabel metal1 s 11362 2 11422 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal3 s -24 10716 -16 10724 7 FreeSans 16 0 0 0 AB[15]
port 2 nsew
flabel metal3 s -24 10676 -16 10684 7 FreeSans 16 0 0 0 AB[14]
port 3 nsew
flabel metal3 s -24 10356 -16 10364 7 FreeSans 16 0 0 0 AB[13]
port 4 nsew
flabel metal3 s -24 10316 -16 10324 7 FreeSans 16 0 0 0 AB[12]
port 5 nsew
flabel metal3 s -24 10276 -16 10284 7 FreeSans 16 0 0 0 AB[11]
port 6 nsew
flabel metal3 s -24 10236 -16 10244 7 FreeSans 16 0 0 0 AB[10]
port 7 nsew
flabel metal3 s -24 10196 -16 10204 7 FreeSans 16 0 0 0 AB[9]
port 8 nsew
flabel metal3 s -24 8996 -16 9004 7 FreeSans 16 0 0 0 AB[8]
port 9 nsew
flabel metal2 s 3377 -23 3383 -17 7 FreeSans 16 270 0 0 AB[7]
port 10 nsew
flabel metal2 s 3617 -23 3623 -17 7 FreeSans 16 270 0 0 AB[6]
port 11 nsew
flabel metal2 s 5377 -23 5383 -17 7 FreeSans 16 270 0 0 AB[5]
port 12 nsew
flabel metal2 s 6357 -23 6363 -17 7 FreeSans 16 270 0 0 AB[4]
port 13 nsew
flabel metal2 s 6397 -23 6403 -17 7 FreeSans 16 270 0 0 AB[3]
port 14 nsew
flabel metal2 s 6437 -23 6443 -17 7 FreeSans 16 270 0 0 AB[2]
port 15 nsew
flabel metal2 s 8097 -23 8103 -17 7 FreeSans 16 270 0 0 AB[1]
port 16 nsew
flabel metal2 s 8137 -23 8143 -17 7 FreeSans 16 270 0 0 AB[0]
port 17 nsew
flabel metal2 s 8337 11337 8343 11343 3 FreeSans 16 90 0 0 DI[7]
port 18 nsew
flabel metal2 s 8157 11337 8163 11343 3 FreeSans 16 90 0 0 DI[6]
port 19 nsew
flabel metal2 s 7437 11337 7443 11343 3 FreeSans 16 90 0 0 DI[5]
port 20 nsew
flabel metal2 s 7177 11337 7183 11343 3 FreeSans 16 90 0 0 DI[4]
port 21 nsew
flabel metal2 s 7137 11337 7143 11343 3 FreeSans 16 90 0 0 DI[3]
port 22 nsew
flabel metal2 s 6977 11337 6983 11343 3 FreeSans 16 90 0 0 DI[2]
port 23 nsew
flabel metal2 s 6737 11337 6743 11343 3 FreeSans 16 90 0 0 DI[1]
port 24 nsew
flabel metal2 s 4377 11337 4383 11343 3 FreeSans 16 90 0 0 DI[0]
port 25 nsew
flabel metal3 s 11396 8356 11404 8364 3 FreeSans 16 0 0 0 DO[7]
port 26 nsew
flabel metal3 s 11396 8316 11404 8324 3 FreeSans 16 0 0 0 DO[6]
port 27 nsew
flabel metal3 s 11396 8276 11404 8284 3 FreeSans 16 0 0 0 DO[5]
port 28 nsew
flabel metal3 s 11396 7796 11404 7804 3 FreeSans 16 0 0 0 DO[4]
port 29 nsew
flabel metal3 s 11396 7576 11404 7584 3 FreeSans 16 0 0 0 DO[3]
port 30 nsew
flabel metal3 s 11396 7536 11404 7544 3 FreeSans 16 0 0 0 DO[2]
port 31 nsew
flabel metal3 s 11396 7316 11404 7324 3 FreeSans 16 0 0 0 DO[1]
port 32 nsew
flabel metal3 s 11396 7076 11404 7084 3 FreeSans 16 0 0 0 DO[0]
port 33 nsew
flabel metal2 s 3937 11337 3943 11343 3 FreeSans 16 90 0 0 IRQ
port 34 nsew
flabel metal3 s -24 5936 -16 5944 7 FreeSans 16 0 0 0 NMI
port 35 nsew
flabel metal2 s 4137 11337 4143 11343 3 FreeSans 16 90 0 0 RDY
port 36 nsew
flabel metal3 s 11396 5396 11404 5404 3 FreeSans 16 0 0 0 WE
port 37 nsew
flabel metal3 s -24 3256 -16 3264 7 FreeSans 16 0 0 0 clk
port 38 nsew
flabel metal3 s -24 4956 -16 4964 7 FreeSans 16 0 0 0 reset
port 39 nsew
<< properties >>
string FIXED_BBOX -40 -40 11400 11340
<< end >>
