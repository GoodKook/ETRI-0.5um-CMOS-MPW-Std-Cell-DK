magic
tech scmos
magscale 1 2
timestamp 1726561008
<< nwell >>
rect -12 154 152 272
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 50 14 54 54
rect 70 14 74 54
rect 80 14 84 54
rect 100 14 104 54
<< ptransistor >>
rect 20 166 24 246
rect 40 166 44 246
rect 50 166 54 246
rect 70 166 74 246
rect 80 166 84 246
rect 100 166 104 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 48 40 54
rect 24 14 26 48
rect 38 14 40 48
rect 44 14 50 54
rect 54 14 56 54
rect 68 14 70 54
rect 74 14 80 54
rect 84 48 100 54
rect 84 14 86 48
rect 98 14 100 48
rect 104 14 106 54
<< pdiffusion >>
rect 18 166 20 246
rect 24 180 26 246
rect 38 180 40 246
rect 24 166 40 180
rect 44 166 50 246
rect 54 166 56 246
rect 68 166 70 246
rect 74 166 80 246
rect 84 180 86 246
rect 98 180 100 246
rect 84 166 100 180
rect 104 166 106 246
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 48
rect 56 14 68 54
rect 86 14 98 48
rect 106 14 118 54
<< pdcontact >>
rect 6 166 18 246
rect 26 180 38 246
rect 56 166 68 246
rect 86 180 98 246
rect 106 166 118 246
<< psubstratepcontact >>
rect -6 -6 146 6
<< nsubstratencontact >>
rect -6 254 146 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 50 246 54 250
rect 70 246 74 250
rect 80 246 84 250
rect 100 246 104 250
rect 20 102 24 166
rect 40 160 44 166
rect 17 90 24 102
rect 20 54 24 90
rect 28 156 44 160
rect 28 62 32 156
rect 50 152 54 166
rect 70 154 74 166
rect 80 164 84 166
rect 100 164 104 166
rect 80 158 104 164
rect 50 148 56 152
rect 70 150 86 154
rect 52 114 56 148
rect 52 108 66 114
rect 82 110 86 150
rect 52 86 54 98
rect 28 58 44 62
rect 40 54 44 58
rect 50 54 54 86
rect 62 82 66 108
rect 62 78 74 82
rect 70 54 74 78
rect 100 74 104 158
rect 80 68 104 74
rect 80 54 84 68
rect 100 54 104 68
rect 20 10 24 14
rect 40 10 44 14
rect 50 10 54 14
rect 70 10 74 14
rect 80 10 84 14
rect 100 10 104 14
<< polycontact >>
rect 5 90 17 102
rect 32 128 44 140
rect 40 108 52 120
rect 40 86 52 98
rect 74 98 86 110
rect 104 116 116 128
<< metal1 >>
rect -6 266 146 268
rect -6 252 146 254
rect 26 246 38 252
rect 86 246 98 252
rect 18 166 36 172
rect 60 156 68 166
rect 100 166 106 174
rect 60 150 70 156
rect 64 136 70 150
rect 17 108 40 116
rect 58 116 74 122
rect 10 66 52 72
rect 58 78 65 116
rect 10 54 18 66
rect 58 64 63 78
rect 58 54 66 64
rect 100 54 118 60
rect 26 8 38 14
rect 86 8 98 14
rect -6 6 146 8
rect -6 -8 146 -6
<< m2contact >>
rect 22 152 36 166
rect 86 160 100 174
rect 43 140 57 142
rect 43 128 44 140
rect 44 128 57 140
rect 63 122 77 136
rect 3 102 17 116
rect 38 72 52 86
rect 103 102 117 116
rect 71 84 85 98
rect 63 64 77 78
rect 86 54 100 68
<< metal2 >>
rect 6 116 14 134
rect 28 92 34 152
rect 66 136 74 154
rect 51 112 57 128
rect 89 112 97 160
rect 51 104 97 112
rect 28 86 71 92
rect 28 84 38 86
rect 52 84 71 86
rect 91 68 97 104
rect 106 86 114 102
rect 66 46 74 64
<< m1p >>
rect -6 252 146 268
rect -6 -8 146 8
<< m2p >>
rect 66 138 74 154
rect 6 118 14 134
rect 106 86 114 100
rect 66 46 74 62
<< labels >>
rlabel metal1 -6 252 126 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -6 -8 126 8 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal2 10 130 10 130 1 A
port 1 n signal input
rlabel metal2 70 152 70 152 5 Y
port 3 n signal output
rlabel metal2 70 50 70 50 1 Y
port 3 n signal output
rlabel metal2 110 90 110 90 5 B
port 2 n signal input
<< properties >>
string FIXED_BBOX 0 0 140 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
