magic
tech scmos
magscale 1 3
timestamp 1569139307
<< checkpaint >>
rect -52 -52 192 88
<< pseudo_rpoly2 >>
rect 8 8 132 28
use poly2cont_CDNS_704676826059  poly2cont_CDNS_704676826059_0
timestamp 1569139307
transform 1 0 114 0 1 8
box 0 0 18 20
use poly2cont_CDNS_704676826059  poly2cont_CDNS_704676826059_1
timestamp 1569139307
transform 1 0 8 0 1 8
box 0 0 18 20
<< end >>
