magic
tech scmos
magscale 1 2
timestamp 1702306454
<< nwell >>
rect -13 154 73 272
<< ntransistor >>
rect 18 14 22 54
rect 38 14 42 54
<< ptransistor >>
rect 18 166 22 246
rect 38 166 42 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 14 24 54
rect 36 14 38 54
rect 42 14 44 54
<< pdiffusion >>
rect 4 245 18 246
rect 16 166 18 245
rect 22 166 24 246
rect 36 166 38 246
rect 42 166 44 246
<< ndcontact >>
rect 4 14 16 54
rect 24 14 36 54
rect 44 14 56 54
<< pdcontact >>
rect 4 166 16 245
rect 24 166 36 246
rect 44 166 56 246
<< psubstratepcontact >>
rect -6 -6 66 6
<< nsubstratencontact >>
rect -6 254 66 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 18 164 22 166
rect 38 164 42 166
rect 18 160 42 164
rect 18 117 22 160
rect 17 105 22 117
rect 18 62 22 105
rect 18 58 42 62
rect 18 54 22 58
rect 38 54 42 58
rect 18 10 22 14
rect 38 10 42 14
<< polycontact >>
rect 5 105 17 117
<< metal1 >>
rect -6 266 66 268
rect -6 252 66 254
rect 4 245 16 252
rect 44 246 56 252
rect 26 151 34 166
rect 26 143 54 151
rect 46 137 54 143
rect 3 123 17 137
rect 43 123 57 137
rect 5 117 17 123
rect 46 73 54 123
rect 26 65 54 73
rect 26 54 34 65
rect 4 8 16 14
rect 44 8 56 14
rect -6 6 66 8
rect -6 -8 66 -6
<< m1p >>
rect -6 252 66 268
rect 3 123 17 137
rect 43 123 57 137
rect -6 -8 66 8
<< labels >>
rlabel nsubstratencontact 30 260 30 260 0 vdd
port 3 nsew power bidirectional abutment
rlabel psubstratepcontact 30 0 30 0 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 10 127 10 127 0 A
port 1 nsew signal input
rlabel metal1 50 130 50 130 0 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 60 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
