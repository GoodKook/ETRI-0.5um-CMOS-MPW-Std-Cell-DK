magic
tech scmos
magscale 1 2
timestamp 1749781262
<< checkpaint >>
rect -48 809 340 834
rect -48 714 342 809
rect -40 142 342 714
rect 1316 553 7715 559
rect -40 54 468 142
rect -48 48 468 54
rect -48 40 480 48
rect -78 -66 480 40
rect -78 -140 468 -66
rect 90 -334 468 -140
rect 90 -664 584 -334
rect 164 -1140 584 -664
rect 164 -1382 542 -1140
rect 1002 -5146 7815 553
<< nwell >>
rect 153 174 172 188
<< metal1 >>
rect 0 0 26 754
rect 250 0 276 754
<< metal2 >>
rect 95 709 106 754
rect 141 715 176 729
rect 95 695 135 709
rect 165 689 176 715
rect 95 675 176 689
rect 95 619 106 675
rect 141 625 176 639
rect 95 605 135 619
rect 165 599 176 625
rect 95 585 176 599
rect 95 529 106 585
rect 141 535 176 549
rect 95 515 135 529
rect 165 509 176 535
rect 95 495 176 509
rect 95 439 106 495
rect 141 445 176 459
rect 95 425 135 439
rect 165 419 176 445
rect 95 405 176 419
rect 95 349 106 405
rect 141 355 176 369
rect 95 335 135 349
rect 165 329 176 355
rect 95 315 176 329
rect 95 259 106 315
rect 141 265 176 279
rect 95 245 135 259
rect 165 239 176 265
rect 95 225 176 239
rect 95 168 106 225
rect 153 174 176 188
rect 95 154 135 168
rect 165 148 176 174
rect 144 137 176 148
rect 144 116 155 137
rect 95 105 155 116
rect 95 77 106 105
rect 145 83 176 97
rect 95 63 135 77
rect 165 57 176 83
rect 146 43 176 57
rect 165 0 176 43
<< m2p >>
rect 95 695 106 754
rect 95 154 106 239
rect 95 105 155 116
rect 165 0 176 11
use NAND2X1  NAND2X1_8 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304996
transform 0 1 18 -1 0 100
box -12 -8 92 252
use NAND2X1  NAND2X1_9
timestamp 1728304996
transform 0 1 18 -1 0 191
box -12 -8 92 252
use NAND2X1  NAND2X1_10
timestamp 1728304996
transform 0 1 18 -1 0 282
box -12 -8 92 252
use NAND2X1  NAND2X1_11
timestamp 1728304996
transform 0 1 18 -1 0 372
box -12 -8 92 252
use NAND2X1  NAND2X1_12
timestamp 1728304996
transform 0 1 18 -1 0 462
box -12 -8 92 252
use NAND2X1  NAND2X1_13
timestamp 1728304996
transform 0 1 18 -1 0 552
box -12 -8 92 252
use NAND2X1  NAND2X1_14
timestamp 1728304996
transform 0 1 18 -1 0 642
box -12 -8 92 252
use NAND2X1  NAND2X1_15
timestamp 1728304996
transform 0 1 18 -1 0 732
box -12 -8 92 252
<< labels >>
rlabel metal1 250 728 276 754 0 vdd
port 1 nsew power bidirectional abutment
rlabel metal1 0 728 26 754 0 gnd
port 2 nsew ground bidirectional abutment
rlabel metal2 165 0 176 11 0 In
port 3 nsew signal input
rlabel metal2 95 105 155 116 0 Out1
port 4 nsew signal output
rlabel metal2 95 154 106 239 0 Out2
port 5 nsew signal output
rlabel metal2 95 695 106 754 0 Out3
port 6 nsew signal output
<< end >>
