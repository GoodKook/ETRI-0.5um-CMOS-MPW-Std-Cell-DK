** sch_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/DFFSR.sch
**.subckt DFFSR D R S CLK Q vdd gnd
*.ipin CLK
*.ipin D
*.opin Q
*.ipin S
*.ipin R
*.iopin vdd
*.iopin gnd
M1 net1 C_Bar net2 VDD pfet w=3u l=0.6u m=1
M2 net1 C net2 GND nfet w=3u l=0.6u m=1
M3 net5 C net2 VDD pfet w=3u l=0.6u m=1
M4 net5 C_Bar net2 GND nfet w=3u l=0.6u m=1
M6 net4 C_Bar net3 VDD pfet w=3u l=0.6u m=1
M5 net4 C net3 GND nfet w=3u l=0.6u m=1
M7 net4 C net6 VDD pfet w=3u l=0.6u m=1
M8 net4 C_Bar net6 GND nfet w=3u l=0.6u m=1
x1 CLK C_Bar vdd gnd INVX1
x2 C_Bar C vdd gnd INVX1
x4 S net2 net3 vdd gnd NAND2X1
x6 R net3 net1 vdd gnd NAND2X1
x7 R net4 net7 vdd gnd NAND2X1
x8 net7 S net6 vdd gnd NAND2X1
x3 D net5 vdd gnd INVX1
x5 net7 Q vdd gnd INVX1
**.ends

* expanding   symbol:  /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/INVX1.sym # of pins=4
** sym_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/INVX1.sym
** sch_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/INVX1.sch
.subckt INVX1 A Y vdd gnd
*.ipin A
*.opin Y
*.iopin vdd
*.iopin gnd
M1 Y A gnd GND nfet w=3u l=0.6u m=1
M2 Y A vdd VDD pfet w=6u l=0.6u m=1
.ends


* expanding   symbol:  /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/NAND2X1.sym # of pins=5
** sym_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/NAND2X1.sym
** sch_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/NAND2X1.sch
.subckt NAND2X1 A B Y vdd gnd
*.ipin A
*.ipin B
*.opin Y
*.iopin vdd
*.iopin gnd
M1 Y B net1 GND nfet w=6u l=0.6u m=1
M2 Y B vdd VDD pfet w=6u l=0.6u m=1
M3 net1 A gnd GND nfet w=6u l=0.6u m=1
M4 Y A vdd VDD pfet w=6u l=0.6u m=1
.ends

.end
