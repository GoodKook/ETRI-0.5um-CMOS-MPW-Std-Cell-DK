magic
tech scmos
magscale 1 3
timestamp 1725340527
<< checkpaint >>
rect -44 435 158 438
rect -44 432 170 435
rect -58 425 170 432
rect 278 425 454 435
rect -58 312 454 425
rect -58 116 470 312
rect -58 -36 459 116
rect -55 -38 459 -36
<< nwell >>
rect 35 300 375 375
rect 35 110 110 300
rect 300 110 375 300
rect 35 35 375 110
<< psubstratepdiff >>
rect 130 260 280 280
rect 130 150 150 260
rect 260 150 280 260
rect 130 130 280 150
<< nsubstratendiff >>
rect 45 345 365 365
rect 45 65 65 345
rect 195 195 215 215
rect 345 65 365 345
rect 45 45 365 65
<< genericcontact >>
rect 70 345 340 365
rect 45 75 65 340
rect 150 260 260 280
rect 130 150 150 260
rect 195 195 215 215
rect 260 150 280 260
rect 150 130 260 150
rect 345 70 365 340
rect 70 45 340 65
<< metal1 >>
rect 45 345 365 365
rect 45 65 65 345
rect 130 260 280 280
rect 130 150 150 260
rect 195 195 215 215
rect 260 150 280 260
rect 130 130 280 150
rect 345 65 365 345
rect 45 45 365 65
<< end >>
