magic
tech scmos
magscale 2 1
timestamp 1756367800
<< checkpaint >>
rect -39 402 403 450
rect -39 -40 451 402
<< metal1 >>
rect 1 290 407 362
rect 1 259 51 290
rect 57 278 70 290
rect 57 259 70 273
rect 76 259 82 290
rect 88 289 113 290
rect 124 289 148 290
rect 88 288 111 289
rect 126 288 148 289
rect 88 287 110 288
rect 128 287 148 288
rect 88 286 109 287
rect 88 284 108 286
rect 129 285 148 287
rect 170 285 174 290
rect 116 284 121 285
rect 88 280 107 284
rect 114 283 123 284
rect 114 281 124 283
rect 130 282 148 285
rect 131 281 148 282
rect 115 280 148 281
rect 88 278 108 280
rect 117 279 148 280
rect 121 278 148 279
rect 88 276 109 278
rect 125 277 148 278
rect 155 277 174 285
rect 127 276 148 277
rect 88 275 110 276
rect 128 275 148 276
rect 88 274 112 275
rect 129 274 148 275
rect 88 273 114 274
rect 130 273 148 274
rect 88 272 118 273
rect 88 271 121 272
rect 88 270 124 271
rect 88 269 108 270
rect 88 267 106 269
rect 113 267 125 270
rect 88 264 107 267
rect 114 266 124 267
rect 115 265 124 266
rect 117 264 121 265
rect 131 264 148 273
rect 168 272 174 277
rect 104 263 108 264
rect 130 263 148 264
rect 104 262 109 263
rect 129 262 148 263
rect 104 261 110 262
rect 128 261 148 262
rect 104 260 111 261
rect 127 260 148 261
rect 104 259 113 260
rect 125 259 148 260
rect 155 259 174 272
rect 181 259 186 290
rect 206 289 229 290
rect 208 288 229 289
rect 209 287 229 288
rect 210 285 229 287
rect 250 285 255 290
rect 261 285 267 290
rect 192 284 202 285
rect 192 282 204 284
rect 192 280 205 282
rect 192 278 204 280
rect 192 277 202 278
rect 211 277 229 285
rect 235 282 267 285
rect 235 277 255 282
rect 210 276 229 277
rect 209 275 229 276
rect 208 274 229 275
rect 207 273 229 274
rect 204 272 229 273
rect 248 272 255 277
rect 192 271 196 272
rect 205 271 229 272
rect 192 270 198 271
rect 206 270 229 271
rect 192 269 199 270
rect 207 269 229 270
rect 192 267 200 269
rect 208 268 229 269
rect 192 266 201 267
rect 209 266 229 268
rect 192 264 202 266
rect 210 265 229 266
rect 192 263 203 264
rect 211 263 229 265
rect 192 261 204 263
rect 212 261 229 263
rect 192 260 205 261
rect 213 260 229 261
rect 192 259 206 260
rect 214 259 229 260
rect 235 259 255 272
rect 261 259 267 282
rect 273 289 407 290
rect 273 288 284 289
rect 273 287 282 288
rect 273 286 280 287
rect 273 282 279 286
rect 285 283 407 289
rect 285 282 298 283
rect 305 282 325 283
rect 330 282 407 283
rect 273 277 276 282
rect 289 281 296 282
rect 307 281 316 282
rect 289 279 294 281
rect 309 279 316 281
rect 322 281 324 282
rect 322 280 323 281
rect 331 280 407 282
rect 289 278 293 279
rect 310 278 316 279
rect 330 278 407 280
rect 289 277 292 278
rect 300 277 303 278
rect 273 261 279 277
rect 285 276 292 277
rect 299 276 305 277
rect 285 266 291 276
rect 298 275 305 276
rect 311 275 316 278
rect 329 277 407 278
rect 325 276 407 277
rect 324 275 407 276
rect 298 274 306 275
rect 297 273 306 274
rect 312 269 316 275
rect 297 268 316 269
rect 298 266 316 268
rect 285 265 292 266
rect 299 265 305 266
rect 310 265 316 266
rect 286 264 288 265
rect 289 264 292 265
rect 300 264 304 265
rect 289 262 293 264
rect 311 263 316 265
rect 310 262 316 263
rect 290 261 294 262
rect 309 261 316 262
rect 273 260 280 261
rect 290 260 296 261
rect 308 260 316 261
rect 273 259 282 260
rect 289 259 297 260
rect 306 259 316 260
rect 323 259 407 275
rect 1 234 407 259
rect 1 228 66 234
rect 70 233 80 234
rect 84 233 85 234
rect 70 231 79 233
rect 83 231 85 233
rect 89 233 102 234
rect 89 232 96 233
rect 89 231 95 232
rect 97 231 101 233
rect 106 232 133 234
rect 105 231 132 232
rect 70 230 78 231
rect 82 230 94 231
rect 71 228 77 230
rect 82 229 93 230
rect 97 229 132 231
rect 137 230 144 234
rect 149 233 152 234
rect 148 231 152 233
rect 156 233 171 234
rect 178 233 218 234
rect 226 233 315 234
rect 322 233 407 234
rect 156 232 169 233
rect 180 232 217 233
rect 227 232 267 233
rect 268 232 313 233
rect 323 232 407 233
rect 1 223 67 228
rect 71 226 76 228
rect 81 227 84 229
rect 71 224 75 226
rect 80 225 84 227
rect 88 226 90 229
rect 99 228 101 229
rect 105 228 110 229
rect 117 228 132 229
rect 99 227 100 228
rect 105 227 108 228
rect 118 227 132 228
rect 98 226 100 227
rect 1 217 68 223
rect 72 222 74 224
rect 79 223 83 225
rect 88 224 92 226
rect 96 224 100 226
rect 72 220 73 222
rect 78 221 83 223
rect 77 220 83 221
rect 87 220 91 224
rect 95 223 100 224
rect 76 218 82 220
rect 87 219 90 220
rect 95 219 99 223
rect 104 222 107 227
rect 111 225 114 226
rect 111 224 115 225
rect 119 224 131 227
rect 136 226 143 230
rect 148 228 151 231
rect 156 230 168 232
rect 181 231 216 232
rect 228 231 265 232
rect 268 231 312 232
rect 324 231 407 232
rect 173 230 176 231
rect 181 230 215 231
rect 220 230 223 231
rect 229 230 264 231
rect 267 230 311 231
rect 156 229 167 230
rect 147 226 151 228
rect 155 226 167 229
rect 171 229 177 230
rect 182 229 215 230
rect 171 228 178 229
rect 182 228 191 229
rect 195 228 200 229
rect 172 227 192 228
rect 174 226 192 227
rect 196 226 199 228
rect 205 227 215 229
rect 219 228 225 230
rect 229 229 263 230
rect 267 229 310 230
rect 317 229 320 230
rect 325 229 407 231
rect 229 228 231 229
rect 220 227 231 228
rect 204 226 215 227
rect 222 226 231 227
rect 114 223 131 224
rect 147 223 150 226
rect 155 225 168 226
rect 176 225 192 226
rect 197 225 198 226
rect 203 225 215 226
rect 224 225 231 226
rect 235 227 241 229
rect 245 228 249 229
rect 256 228 261 229
rect 269 228 273 229
rect 279 228 286 229
rect 290 228 291 229
rect 296 228 299 229
rect 304 228 309 229
rect 315 228 321 229
rect 245 227 247 228
rect 257 227 260 228
rect 235 225 240 227
rect 244 226 247 227
rect 258 226 260 227
rect 269 227 272 228
rect 281 227 286 228
rect 297 227 298 228
rect 305 227 309 228
rect 314 227 322 228
rect 326 227 407 229
rect 269 226 271 227
rect 281 226 285 227
rect 244 225 246 226
rect 251 225 253 226
rect 259 225 262 226
rect 155 224 169 225
rect 178 224 193 225
rect 202 224 216 225
rect 226 224 232 225
rect 116 222 121 223
rect 128 222 131 223
rect 1 214 69 217
rect 75 216 82 218
rect 74 215 82 216
rect 86 215 90 219
rect 94 218 99 219
rect 103 221 108 222
rect 117 221 120 222
rect 103 220 110 221
rect 103 219 113 220
rect 118 219 120 221
rect 128 219 130 222
rect 135 220 142 222
rect 94 217 98 218
rect 103 217 105 219
rect 109 218 114 219
rect 110 217 113 218
rect 118 217 130 219
rect 134 219 142 220
rect 146 221 150 223
rect 154 223 170 224
rect 179 223 193 224
rect 201 223 218 224
rect 154 222 172 223
rect 154 221 174 222
rect 180 221 194 223
rect 200 222 220 223
rect 227 222 232 224
rect 199 221 222 222
rect 97 215 98 217
rect 74 214 81 215
rect 86 214 91 215
rect 96 214 98 215
rect 102 216 105 217
rect 118 216 129 217
rect 102 215 106 216
rect 117 215 129 216
rect 134 215 141 219
rect 146 217 149 221
rect 154 220 176 221
rect 154 219 165 220
rect 169 219 176 220
rect 153 218 165 219
rect 170 218 176 219
rect 180 219 193 221
rect 199 220 223 221
rect 180 218 192 219
rect 200 218 213 220
rect 217 218 224 220
rect 228 219 232 222
rect 236 223 239 225
rect 243 223 246 225
rect 250 224 255 225
rect 258 224 262 225
rect 253 223 262 224
rect 236 222 238 223
rect 242 222 246 223
rect 255 222 262 223
rect 266 224 270 226
rect 275 225 277 226
rect 236 219 237 222
rect 242 221 247 222
rect 241 220 249 221
rect 257 220 261 222
rect 266 221 269 224
rect 274 223 278 225
rect 273 222 279 223
rect 282 222 285 226
rect 291 225 293 226
rect 299 225 301 226
rect 290 224 293 225
rect 241 219 252 220
rect 228 218 233 219
rect 102 214 108 215
rect 115 214 129 215
rect 133 214 141 215
rect 145 216 149 217
rect 163 217 165 218
rect 171 217 175 218
rect 180 217 191 218
rect 163 216 166 217
rect 179 216 190 217
rect 195 216 197 217
rect 201 216 213 218
rect 218 217 222 218
rect 227 216 233 218
rect 240 217 244 219
rect 248 218 253 219
rect 258 218 261 220
rect 249 217 253 218
rect 145 214 148 216
rect 163 215 167 216
rect 178 215 189 216
rect 194 215 197 216
rect 202 215 214 216
rect 226 215 233 216
rect 239 215 245 217
rect 257 216 260 218
rect 265 217 269 221
rect 282 220 284 222
rect 289 221 293 224
rect 298 223 302 225
rect 273 218 284 220
rect 274 217 277 218
rect 267 216 270 217
rect 281 216 284 218
rect 288 220 293 221
rect 288 216 292 220
rect 297 219 301 223
rect 306 222 308 227
rect 313 225 407 227
rect 256 215 261 216
rect 163 214 169 215
rect 177 214 188 215
rect 193 214 198 215
rect 202 214 216 215
rect 224 214 233 215
rect 1 213 233 214
rect 238 214 247 215
rect 255 214 261 215
rect 267 215 271 216
rect 280 215 283 216
rect 267 214 272 215
rect 279 214 283 215
rect 287 215 292 216
rect 296 218 301 219
rect 305 218 308 222
rect 312 221 407 225
rect 312 220 320 221
rect 313 219 319 220
rect 314 218 318 219
rect 324 218 407 221
rect 287 214 291 215
rect 296 214 300 218
rect 305 217 309 218
rect 323 217 407 218
rect 304 216 310 217
rect 322 216 407 217
rect 304 215 311 216
rect 321 215 407 216
rect 304 214 312 215
rect 319 214 407 215
rect 238 213 407 214
rect 1 212 232 213
rect 1 209 229 212
rect 237 211 407 213
rect 236 210 407 211
rect 235 209 407 210
rect 1 149 407 209
rect 1 145 75 149
rect 81 147 87 149
rect 93 148 116 149
rect 123 148 131 149
rect 93 147 114 148
rect 125 147 131 148
rect 1 140 74 145
rect 81 144 86 147
rect 93 146 113 147
rect 93 145 112 146
rect 126 145 131 147
rect 135 146 147 149
rect 152 148 222 149
rect 151 147 222 148
rect 228 148 234 149
rect 151 146 221 147
rect 135 145 221 146
rect 93 144 111 145
rect 118 144 121 145
rect 1 135 73 140
rect 77 137 78 143
rect 81 142 85 144
rect 82 140 84 142
rect 82 138 83 140
rect 87 138 88 140
rect 92 139 95 144
rect 99 143 105 144
rect 109 143 111 144
rect 116 143 123 144
rect 99 141 104 143
rect 109 142 110 143
rect 99 139 103 141
rect 108 140 110 142
rect 115 142 123 143
rect 127 142 130 145
rect 134 144 221 145
rect 134 143 136 144
rect 141 143 146 144
rect 151 143 154 144
rect 158 143 159 144
rect 164 143 182 144
rect 188 143 195 144
rect 134 142 135 143
rect 115 141 130 142
rect 142 141 146 143
rect 92 138 96 139
rect 1 130 72 135
rect 76 131 78 137
rect 86 137 88 138
rect 86 136 87 137
rect 85 133 87 136
rect 84 132 87 133
rect 91 132 96 138
rect 100 137 102 139
rect 107 138 110 140
rect 100 135 101 137
rect 106 136 110 138
rect 105 134 110 136
rect 114 140 130 141
rect 136 140 138 141
rect 114 136 129 140
rect 134 138 138 140
rect 143 139 146 141
rect 150 142 154 143
rect 165 142 180 143
rect 190 142 195 143
rect 199 143 201 144
rect 206 143 221 144
rect 199 142 200 143
rect 207 142 221 143
rect 228 146 233 148
rect 240 147 259 149
rect 270 148 307 149
rect 312 148 407 149
rect 271 147 307 148
rect 228 143 232 146
rect 239 144 258 147
rect 272 146 307 147
rect 114 135 122 136
rect 126 135 129 136
rect 133 135 138 138
rect 114 134 121 135
rect 126 134 128 135
rect 133 134 137 135
rect 142 134 145 139
rect 150 138 153 142
rect 166 141 179 142
rect 159 140 161 141
rect 166 140 178 141
rect 184 140 186 141
rect 158 139 162 140
rect 167 139 178 140
rect 182 139 187 140
rect 191 139 195 142
rect 201 140 203 141
rect 200 139 204 140
rect 149 137 153 138
rect 157 137 163 139
rect 167 138 177 139
rect 104 132 110 134
rect 116 133 119 134
rect 125 132 128 134
rect 84 131 86 132
rect 1 129 71 130
rect 75 129 79 131
rect 83 129 86 131
rect 90 129 97 132
rect 103 131 111 132
rect 124 131 128 132
rect 103 130 112 131
rect 123 130 128 131
rect 132 130 137 134
rect 1 128 97 129
rect 102 129 114 130
rect 121 129 127 130
rect 132 129 136 130
rect 141 129 144 134
rect 149 133 152 137
rect 157 136 162 137
rect 167 136 168 138
rect 176 137 177 138
rect 182 137 188 139
rect 156 135 162 136
rect 157 134 162 135
rect 166 134 167 135
rect 175 134 177 137
rect 181 134 187 137
rect 192 136 194 139
rect 199 138 204 139
rect 208 138 220 142
rect 228 141 231 143
rect 239 142 241 144
rect 245 142 251 144
rect 256 143 258 144
rect 255 142 258 143
rect 262 144 267 145
rect 273 144 307 146
rect 311 144 407 148
rect 239 141 242 142
rect 199 137 203 138
rect 191 134 194 136
rect 198 134 203 137
rect 207 134 209 138
rect 217 137 220 138
rect 223 139 224 140
rect 228 139 230 141
rect 234 139 235 141
rect 217 135 219 137
rect 216 134 219 135
rect 223 134 225 139
rect 228 137 229 139
rect 233 137 234 139
rect 232 134 234 137
rect 238 136 242 141
rect 246 140 250 142
rect 255 141 257 142
rect 246 138 249 140
rect 254 139 257 141
rect 262 140 269 144
rect 273 143 279 144
rect 285 143 293 144
rect 301 143 306 144
rect 311 143 314 144
rect 319 143 407 144
rect 246 136 248 138
rect 253 137 257 139
rect 261 137 269 140
rect 274 142 278 143
rect 287 142 292 143
rect 302 142 306 143
rect 274 141 277 142
rect 287 141 291 142
rect 274 139 276 141
rect 281 140 283 141
rect 274 138 275 139
rect 280 138 284 140
rect 238 135 243 136
rect 246 135 247 136
rect 252 135 256 137
rect 261 135 268 137
rect 273 135 275 138
rect 279 137 285 138
rect 288 137 291 141
rect 295 140 298 141
rect 295 139 299 140
rect 303 139 306 142
rect 310 142 313 143
rect 318 142 407 143
rect 310 141 312 142
rect 317 141 407 142
rect 310 140 311 141
rect 316 140 407 141
rect 315 139 407 140
rect 297 138 305 139
rect 300 137 305 138
rect 314 137 407 139
rect 288 136 292 137
rect 301 136 305 137
rect 288 135 294 136
rect 157 133 161 134
rect 166 133 177 134
rect 182 133 186 134
rect 191 133 193 134
rect 198 133 202 134
rect 207 133 219 134
rect 148 132 152 133
rect 158 132 160 133
rect 148 129 151 132
rect 165 131 178 133
rect 183 132 185 133
rect 190 131 193 133
rect 164 130 179 131
rect 189 130 193 131
rect 102 128 151 129
rect 1 127 96 128
rect 101 127 151 128
rect 155 129 157 130
rect 162 129 180 130
rect 187 129 193 130
rect 197 129 202 133
rect 206 129 218 133
rect 222 129 225 134
rect 231 132 233 134
rect 230 130 233 132
rect 229 129 233 130
rect 237 129 243 135
rect 251 133 256 135
rect 260 134 267 135
rect 260 133 265 134
rect 272 133 275 135
rect 279 134 296 135
rect 302 134 305 136
rect 310 134 311 135
rect 315 134 407 137
rect 279 133 289 134
rect 293 133 298 134
rect 250 132 256 133
rect 271 132 275 133
rect 280 132 283 133
rect 250 131 255 132
rect 270 131 276 132
rect 287 131 289 133
rect 294 132 297 133
rect 302 132 304 134
rect 309 133 312 134
rect 249 129 255 131
rect 269 130 277 131
rect 286 130 290 131
rect 301 130 304 132
rect 267 129 278 130
rect 285 129 292 130
rect 299 129 304 130
rect 308 130 312 133
rect 316 130 407 134
rect 308 129 313 130
rect 317 129 407 130
rect 155 128 243 129
rect 155 127 242 128
rect 248 127 407 129
rect 1 124 93 127
rect 100 125 150 127
rect 155 126 239 127
rect 247 126 407 127
rect 98 124 150 125
rect 154 124 239 126
rect 246 125 407 126
rect 245 124 407 125
rect 1 111 407 124
rect 1 110 82 111
rect 88 110 95 111
rect 100 110 106 111
rect 111 110 117 111
rect 126 110 136 111
rect 141 110 162 111
rect 1 109 81 110
rect 89 109 94 110
rect 101 109 105 110
rect 112 109 117 110
rect 125 109 135 110
rect 142 109 162 110
rect 1 107 80 109
rect 84 107 86 109
rect 1 105 86 107
rect 90 108 93 109
rect 90 106 92 108
rect 96 107 98 109
rect 101 108 104 109
rect 108 108 109 109
rect 113 108 117 109
rect 90 105 91 106
rect 1 104 85 105
rect 1 103 84 104
rect 89 103 91 105
rect 95 104 98 107
rect 1 102 83 103
rect 88 102 91 103
rect 1 101 82 102
rect 87 101 91 102
rect 1 100 81 101
rect 86 100 91 101
rect 1 98 80 100
rect 85 99 91 100
rect 84 98 91 99
rect 94 101 98 104
rect 102 107 104 108
rect 107 107 110 108
rect 102 106 110 107
rect 102 105 109 106
rect 102 104 108 105
rect 113 104 116 108
rect 120 107 134 109
rect 138 108 139 109
rect 143 108 162 109
rect 165 108 174 111
rect 179 109 183 111
rect 188 110 206 111
rect 213 110 219 111
rect 188 109 205 110
rect 214 109 219 110
rect 222 109 232 111
rect 235 110 257 111
rect 235 109 256 110
rect 137 107 140 108
rect 119 106 140 107
rect 143 107 161 108
rect 143 106 146 107
rect 149 106 150 107
rect 153 106 155 107
rect 160 106 161 107
rect 165 106 173 108
rect 179 107 182 109
rect 188 108 204 109
rect 188 107 203 108
rect 208 107 211 108
rect 123 105 139 106
rect 143 105 145 106
rect 153 105 154 106
rect 124 104 137 105
rect 142 104 145 105
rect 152 104 154 105
rect 157 104 159 105
rect 164 104 173 106
rect 102 103 107 104
rect 112 103 115 104
rect 119 103 121 104
rect 101 102 106 103
rect 111 102 121 103
rect 125 103 137 104
rect 141 103 145 104
rect 150 103 153 104
rect 125 102 138 103
rect 101 101 105 102
rect 111 101 122 102
rect 94 99 97 101
rect 101 100 104 101
rect 110 100 114 101
rect 100 99 104 100
rect 109 99 114 100
rect 118 99 121 101
rect 125 100 139 102
rect 94 98 96 99
rect 100 98 103 99
rect 108 98 115 99
rect 118 98 120 99
rect 124 98 132 100
rect 135 99 139 100
rect 142 101 145 103
rect 149 102 153 103
rect 142 99 144 101
rect 148 99 152 102
rect 156 99 160 104
rect 164 101 172 104
rect 163 99 172 101
rect 175 99 176 106
rect 179 104 181 107
rect 179 102 180 104
rect 183 102 184 104
rect 187 102 190 107
rect 193 105 197 107
rect 201 106 202 107
rect 193 103 196 105
rect 200 104 202 106
rect 206 106 212 107
rect 215 106 218 109
rect 222 108 256 109
rect 221 107 256 108
rect 221 106 222 107
rect 227 106 231 107
rect 206 105 218 106
rect 205 104 218 105
rect 222 104 224 105
rect 182 100 183 102
rect 187 101 191 102
rect 194 101 195 103
rect 199 102 201 104
rect 198 101 201 102
rect 205 101 217 104
rect 221 102 224 104
rect 228 104 231 106
rect 234 104 237 107
rect 240 106 241 107
rect 245 106 256 107
rect 262 109 266 111
rect 262 107 265 109
rect 271 108 274 111
rect 284 110 287 111
rect 285 109 287 110
rect 286 108 287 109
rect 291 109 295 111
rect 299 109 304 111
rect 308 110 407 111
rect 246 105 256 106
rect 241 104 243 105
rect 228 103 230 104
rect 234 103 236 104
rect 136 98 138 99
rect 1 96 79 98
rect 89 97 92 98
rect 99 97 103 98
rect 112 97 115 98
rect 123 97 133 98
rect 141 97 144 99
rect 88 96 93 97
rect 98 96 102 97
rect 112 96 116 97
rect 122 96 134 97
rect 139 96 144 97
rect 147 97 153 99
rect 157 98 159 99
rect 163 97 171 99
rect 147 96 154 97
rect 162 96 171 97
rect 174 98 176 99
rect 174 96 177 98
rect 181 97 183 100
rect 180 96 182 97
rect 186 96 191 101
rect 198 100 202 101
rect 205 100 211 101
rect 197 99 202 100
rect 206 99 209 100
rect 214 99 217 101
rect 220 99 224 102
rect 227 99 230 103
rect 233 100 236 103
rect 240 102 244 104
rect 239 101 244 102
rect 196 98 202 99
rect 213 98 216 99
rect 220 98 223 99
rect 227 98 229 99
rect 233 98 235 100
rect 239 99 243 101
rect 247 100 255 105
rect 258 100 259 106
rect 262 105 264 107
rect 270 106 274 108
rect 277 107 282 108
rect 277 106 283 107
rect 262 103 263 105
rect 266 103 267 105
rect 270 103 273 106
rect 277 105 282 106
rect 286 105 288 108
rect 277 104 281 105
rect 285 103 288 105
rect 291 107 294 109
rect 299 107 303 109
rect 307 108 407 110
rect 291 105 293 107
rect 299 105 302 107
rect 306 106 407 108
rect 291 103 292 105
rect 296 104 297 105
rect 265 100 266 102
rect 247 99 254 100
rect 240 98 242 99
rect 246 98 254 99
rect 196 97 203 98
rect 212 97 216 98
rect 1 95 191 96
rect 195 96 204 97
rect 211 96 216 97
rect 219 96 223 98
rect 226 96 229 98
rect 232 96 235 98
rect 245 97 254 98
rect 195 95 235 96
rect 238 96 239 97
rect 244 96 254 97
rect 257 96 259 100
rect 264 98 266 100
rect 269 101 273 103
rect 284 102 288 103
rect 295 102 297 104
rect 300 103 301 105
rect 305 104 407 106
rect 304 102 407 104
rect 283 101 288 102
rect 263 96 265 98
rect 269 97 272 101
rect 276 99 288 101
rect 294 100 297 102
rect 303 100 407 102
rect 268 96 272 97
rect 275 96 288 99
rect 293 98 297 100
rect 302 98 407 100
rect 292 96 297 98
rect 301 96 407 98
rect 1 94 190 95
rect 1 92 188 94
rect 194 93 234 95
rect 238 93 407 96
rect 193 92 234 93
rect 237 92 407 93
rect 1 4 407 92
<< metal2 >>
rect 3 288 409 360
rect 3 257 53 288
rect 59 276 72 288
rect 59 257 72 271
rect 78 257 84 288
rect 90 287 115 288
rect 126 287 150 288
rect 90 286 113 287
rect 128 286 150 287
rect 90 285 112 286
rect 130 285 150 286
rect 90 284 111 285
rect 90 282 110 284
rect 131 283 150 285
rect 172 283 176 288
rect 118 282 123 283
rect 90 278 109 282
rect 116 281 125 282
rect 116 279 126 281
rect 132 280 150 283
rect 133 279 150 280
rect 117 278 150 279
rect 90 276 110 278
rect 119 277 150 278
rect 123 276 150 277
rect 90 274 111 276
rect 127 275 150 276
rect 157 275 176 283
rect 129 274 150 275
rect 90 273 112 274
rect 130 273 150 274
rect 90 272 114 273
rect 131 272 150 273
rect 90 271 116 272
rect 132 271 150 272
rect 90 270 120 271
rect 90 269 123 270
rect 90 268 126 269
rect 90 267 110 268
rect 90 265 108 267
rect 115 265 127 268
rect 90 262 109 265
rect 116 264 126 265
rect 117 263 126 264
rect 119 262 123 263
rect 133 262 150 271
rect 170 270 176 275
rect 106 261 110 262
rect 132 261 150 262
rect 106 260 111 261
rect 131 260 150 261
rect 106 259 112 260
rect 130 259 150 260
rect 106 258 113 259
rect 129 258 150 259
rect 106 257 115 258
rect 127 257 150 258
rect 157 257 176 270
rect 183 257 188 288
rect 208 287 231 288
rect 210 286 231 287
rect 211 285 231 286
rect 212 283 231 285
rect 252 283 257 288
rect 263 283 269 288
rect 194 282 204 283
rect 194 280 206 282
rect 194 278 207 280
rect 194 276 206 278
rect 194 275 204 276
rect 213 275 231 283
rect 237 280 269 283
rect 237 275 257 280
rect 212 274 231 275
rect 211 273 231 274
rect 210 272 231 273
rect 209 271 231 272
rect 206 270 231 271
rect 250 270 257 275
rect 194 269 198 270
rect 207 269 231 270
rect 194 268 200 269
rect 208 268 231 269
rect 194 267 201 268
rect 209 267 231 268
rect 194 265 202 267
rect 210 266 231 267
rect 194 264 203 265
rect 211 264 231 266
rect 194 262 204 264
rect 212 263 231 264
rect 194 261 205 262
rect 213 261 231 263
rect 194 259 206 261
rect 214 259 231 261
rect 194 258 207 259
rect 215 258 231 259
rect 194 257 208 258
rect 216 257 231 258
rect 237 257 257 270
rect 263 257 269 280
rect 275 287 409 288
rect 275 286 286 287
rect 275 285 284 286
rect 275 284 282 285
rect 275 280 281 284
rect 287 281 409 287
rect 287 280 300 281
rect 307 280 327 281
rect 332 280 409 281
rect 275 275 278 280
rect 291 279 298 280
rect 309 279 318 280
rect 291 277 296 279
rect 311 277 318 279
rect 324 279 326 280
rect 324 278 325 279
rect 333 278 409 280
rect 291 276 295 277
rect 312 276 318 277
rect 332 276 409 278
rect 291 275 294 276
rect 302 275 305 276
rect 275 259 281 275
rect 287 274 294 275
rect 301 274 307 275
rect 287 264 293 274
rect 300 273 307 274
rect 313 273 318 276
rect 331 275 409 276
rect 327 274 409 275
rect 326 273 409 274
rect 300 272 308 273
rect 299 271 308 272
rect 314 267 318 273
rect 299 266 318 267
rect 300 264 318 266
rect 287 263 294 264
rect 301 263 307 264
rect 312 263 318 264
rect 288 262 290 263
rect 291 262 294 263
rect 302 262 306 263
rect 291 260 295 262
rect 313 261 318 263
rect 312 260 318 261
rect 292 259 296 260
rect 311 259 318 260
rect 275 258 282 259
rect 292 258 298 259
rect 310 258 318 259
rect 275 257 284 258
rect 291 257 299 258
rect 308 257 318 258
rect 325 257 409 273
rect 3 232 409 257
rect 3 226 68 232
rect 72 231 82 232
rect 86 231 87 232
rect 72 229 81 231
rect 85 229 87 231
rect 91 231 104 232
rect 91 230 98 231
rect 91 229 97 230
rect 99 229 103 231
rect 108 230 135 232
rect 107 229 134 230
rect 72 228 80 229
rect 84 228 96 229
rect 73 226 79 228
rect 84 227 95 228
rect 99 227 134 229
rect 139 228 146 232
rect 151 231 154 232
rect 150 229 154 231
rect 158 231 173 232
rect 180 231 220 232
rect 228 231 317 232
rect 324 231 409 232
rect 158 230 171 231
rect 182 230 219 231
rect 229 230 269 231
rect 270 230 315 231
rect 325 230 409 231
rect 3 221 69 226
rect 73 224 78 226
rect 83 225 86 227
rect 73 222 77 224
rect 82 223 86 225
rect 90 224 92 227
rect 101 226 103 227
rect 107 226 112 227
rect 119 226 134 227
rect 101 225 102 226
rect 107 225 110 226
rect 120 225 134 226
rect 100 224 102 225
rect 3 215 70 221
rect 74 220 76 222
rect 81 221 85 223
rect 90 222 94 224
rect 98 222 102 224
rect 74 218 75 220
rect 80 219 85 221
rect 79 218 85 219
rect 89 218 93 222
rect 97 221 102 222
rect 78 216 84 218
rect 89 217 92 218
rect 97 217 101 221
rect 106 220 109 225
rect 113 223 116 224
rect 113 222 117 223
rect 121 222 133 225
rect 138 224 145 228
rect 150 226 153 229
rect 158 228 170 230
rect 183 229 218 230
rect 230 229 267 230
rect 270 229 314 230
rect 326 229 409 230
rect 175 228 178 229
rect 183 228 217 229
rect 222 228 225 229
rect 231 228 266 229
rect 269 228 313 229
rect 158 227 169 228
rect 149 224 153 226
rect 157 224 169 227
rect 173 227 179 228
rect 184 227 217 228
rect 173 226 180 227
rect 184 226 193 227
rect 197 226 202 227
rect 174 225 194 226
rect 176 224 194 225
rect 198 224 201 226
rect 207 225 217 227
rect 221 226 227 228
rect 231 227 265 228
rect 269 227 312 228
rect 319 227 322 228
rect 327 227 409 229
rect 231 226 233 227
rect 222 225 233 226
rect 206 224 217 225
rect 224 224 233 225
rect 116 221 133 222
rect 149 221 152 224
rect 157 223 170 224
rect 178 223 194 224
rect 199 223 200 224
rect 205 223 217 224
rect 226 223 233 224
rect 237 225 243 227
rect 247 226 251 227
rect 258 226 263 227
rect 271 226 275 227
rect 281 226 288 227
rect 292 226 293 227
rect 298 226 301 227
rect 306 226 311 227
rect 317 226 323 227
rect 247 225 249 226
rect 259 225 262 226
rect 237 223 242 225
rect 246 224 249 225
rect 260 224 262 225
rect 271 225 274 226
rect 283 225 288 226
rect 299 225 300 226
rect 307 225 311 226
rect 316 225 324 226
rect 328 225 409 227
rect 271 224 273 225
rect 283 224 287 225
rect 246 223 248 224
rect 253 223 255 224
rect 261 223 264 224
rect 157 222 171 223
rect 180 222 195 223
rect 204 222 218 223
rect 228 222 234 223
rect 118 220 123 221
rect 130 220 133 221
rect 3 212 71 215
rect 77 214 84 216
rect 76 213 84 214
rect 88 213 92 217
rect 96 216 101 217
rect 105 219 110 220
rect 119 219 122 220
rect 105 218 112 219
rect 105 217 115 218
rect 120 217 122 219
rect 130 217 132 220
rect 137 218 144 220
rect 96 215 100 216
rect 105 215 107 217
rect 111 216 116 217
rect 112 215 115 216
rect 120 215 132 217
rect 136 217 144 218
rect 148 219 152 221
rect 156 221 172 222
rect 181 221 195 222
rect 203 221 220 222
rect 156 220 174 221
rect 156 219 176 220
rect 182 219 196 221
rect 202 220 222 221
rect 229 220 234 222
rect 201 219 224 220
rect 99 213 100 215
rect 76 212 83 213
rect 88 212 93 213
rect 98 212 100 213
rect 104 214 107 215
rect 120 214 131 215
rect 104 213 108 214
rect 119 213 131 214
rect 136 213 143 217
rect 148 215 151 219
rect 156 218 178 219
rect 156 217 167 218
rect 171 217 178 218
rect 155 216 167 217
rect 172 216 178 217
rect 182 217 195 219
rect 201 218 225 219
rect 182 216 194 217
rect 202 216 215 218
rect 219 216 226 218
rect 230 217 234 220
rect 238 221 241 223
rect 245 221 248 223
rect 252 222 257 223
rect 260 222 264 223
rect 255 221 264 222
rect 238 220 240 221
rect 244 220 248 221
rect 257 220 264 221
rect 268 222 272 224
rect 277 223 279 224
rect 238 217 239 220
rect 244 219 249 220
rect 243 218 251 219
rect 259 218 263 220
rect 268 219 271 222
rect 276 221 280 223
rect 275 220 281 221
rect 284 220 287 224
rect 293 223 295 224
rect 301 223 303 224
rect 292 222 295 223
rect 243 217 254 218
rect 230 216 235 217
rect 104 212 110 213
rect 117 212 131 213
rect 135 212 143 213
rect 147 214 151 215
rect 165 215 167 216
rect 173 215 177 216
rect 182 215 193 216
rect 165 214 168 215
rect 181 214 192 215
rect 197 214 199 215
rect 203 214 215 216
rect 220 215 224 216
rect 229 214 235 216
rect 242 215 246 217
rect 250 216 255 217
rect 260 216 263 218
rect 251 215 255 216
rect 147 212 150 214
rect 165 213 169 214
rect 180 213 191 214
rect 196 213 199 214
rect 204 213 216 214
rect 228 213 235 214
rect 241 213 247 215
rect 259 214 262 216
rect 267 215 271 219
rect 284 218 286 220
rect 291 219 295 222
rect 300 221 304 223
rect 275 216 286 218
rect 276 215 279 216
rect 269 214 272 215
rect 283 214 286 216
rect 290 218 295 219
rect 290 214 294 218
rect 299 217 303 221
rect 308 220 310 225
rect 315 223 409 225
rect 258 213 263 214
rect 165 212 171 213
rect 179 212 190 213
rect 195 212 200 213
rect 204 212 218 213
rect 226 212 235 213
rect 3 211 235 212
rect 240 212 249 213
rect 257 212 263 213
rect 269 213 273 214
rect 282 213 285 214
rect 269 212 274 213
rect 281 212 285 213
rect 289 213 294 214
rect 298 216 303 217
rect 307 216 310 220
rect 314 219 409 223
rect 314 218 322 219
rect 315 217 321 218
rect 316 216 320 217
rect 326 216 409 219
rect 289 212 293 213
rect 298 212 302 216
rect 307 215 311 216
rect 325 215 409 216
rect 306 214 312 215
rect 324 214 409 215
rect 306 213 313 214
rect 323 213 409 214
rect 306 212 314 213
rect 321 212 409 213
rect 240 211 409 212
rect 3 210 234 211
rect 3 207 231 210
rect 239 209 409 211
rect 238 208 409 209
rect 237 207 409 208
rect 3 147 409 207
rect 3 143 77 147
rect 83 145 89 147
rect 95 146 118 147
rect 125 146 133 147
rect 95 145 116 146
rect 127 145 133 146
rect 3 138 76 143
rect 83 142 88 145
rect 95 144 115 145
rect 95 143 114 144
rect 128 143 133 145
rect 137 144 149 147
rect 154 146 224 147
rect 153 145 224 146
rect 230 146 236 147
rect 153 144 223 145
rect 137 143 223 144
rect 95 142 113 143
rect 120 142 123 143
rect 3 133 75 138
rect 79 135 80 141
rect 83 140 87 142
rect 84 138 86 140
rect 84 136 85 138
rect 89 136 90 138
rect 94 137 97 142
rect 101 141 107 142
rect 111 141 113 142
rect 118 141 125 142
rect 101 139 106 141
rect 111 140 112 141
rect 101 137 105 139
rect 110 138 112 140
rect 117 140 125 141
rect 129 140 132 143
rect 136 142 223 143
rect 136 141 138 142
rect 143 141 148 142
rect 153 141 156 142
rect 160 141 161 142
rect 166 141 184 142
rect 190 141 197 142
rect 136 140 137 141
rect 117 139 132 140
rect 144 139 148 141
rect 94 136 98 137
rect 3 128 74 133
rect 78 129 80 135
rect 88 135 90 136
rect 88 134 89 135
rect 87 131 89 134
rect 86 130 89 131
rect 93 130 98 136
rect 102 135 104 137
rect 109 136 112 138
rect 102 133 103 135
rect 108 134 112 136
rect 107 132 112 134
rect 116 138 132 139
rect 138 138 140 139
rect 116 134 131 138
rect 136 136 140 138
rect 145 137 148 139
rect 152 140 156 141
rect 167 140 182 141
rect 192 140 197 141
rect 201 141 203 142
rect 208 141 223 142
rect 201 140 202 141
rect 209 140 223 141
rect 230 144 235 146
rect 242 145 261 147
rect 272 146 309 147
rect 314 146 409 147
rect 273 145 309 146
rect 230 141 234 144
rect 241 142 260 145
rect 274 144 309 145
rect 116 133 124 134
rect 128 133 131 134
rect 135 133 140 136
rect 116 132 123 133
rect 128 132 130 133
rect 135 132 139 133
rect 144 132 147 137
rect 152 136 155 140
rect 168 139 181 140
rect 161 138 163 139
rect 168 138 180 139
rect 186 138 188 139
rect 160 137 164 138
rect 169 137 180 138
rect 184 137 189 138
rect 193 137 197 140
rect 203 138 205 139
rect 202 137 206 138
rect 151 135 155 136
rect 159 135 165 137
rect 169 136 179 137
rect 106 130 112 132
rect 118 131 121 132
rect 127 130 130 132
rect 86 129 88 130
rect 3 127 73 128
rect 77 127 81 129
rect 85 127 88 129
rect 92 127 99 130
rect 105 129 113 130
rect 126 129 130 130
rect 105 128 114 129
rect 125 128 130 129
rect 134 128 139 132
rect 3 126 99 127
rect 104 127 116 128
rect 123 127 129 128
rect 134 127 138 128
rect 143 127 146 132
rect 151 131 154 135
rect 159 134 164 135
rect 169 134 170 136
rect 178 135 179 136
rect 184 135 190 137
rect 158 133 164 134
rect 159 132 164 133
rect 168 132 169 133
rect 177 132 179 135
rect 183 132 189 135
rect 194 134 196 137
rect 201 136 206 137
rect 210 136 222 140
rect 230 139 233 141
rect 241 140 243 142
rect 247 140 253 142
rect 258 141 260 142
rect 257 140 260 141
rect 264 142 269 143
rect 275 142 309 144
rect 313 142 409 146
rect 241 139 244 140
rect 201 135 205 136
rect 193 132 196 134
rect 200 132 205 135
rect 209 132 211 136
rect 219 135 222 136
rect 225 137 226 138
rect 230 137 232 139
rect 236 137 237 139
rect 219 133 221 135
rect 218 132 221 133
rect 225 132 227 137
rect 230 135 231 137
rect 235 135 236 137
rect 234 132 236 135
rect 240 134 244 139
rect 248 138 252 140
rect 257 139 259 140
rect 248 136 251 138
rect 256 137 259 139
rect 264 138 271 142
rect 275 141 281 142
rect 287 141 295 142
rect 303 141 308 142
rect 313 141 316 142
rect 321 141 409 142
rect 248 134 250 136
rect 255 135 259 137
rect 263 135 271 138
rect 276 140 280 141
rect 289 140 294 141
rect 304 140 308 141
rect 276 139 279 140
rect 289 139 293 140
rect 276 137 278 139
rect 283 138 285 139
rect 276 136 277 137
rect 282 136 286 138
rect 240 133 245 134
rect 248 133 249 134
rect 254 133 258 135
rect 263 133 270 135
rect 275 133 277 136
rect 281 135 287 136
rect 290 135 293 139
rect 297 138 300 139
rect 297 137 301 138
rect 305 137 308 140
rect 312 140 315 141
rect 320 140 409 141
rect 312 139 314 140
rect 319 139 409 140
rect 312 138 313 139
rect 318 138 409 139
rect 317 137 409 138
rect 299 136 307 137
rect 302 135 307 136
rect 316 135 409 137
rect 290 134 294 135
rect 303 134 307 135
rect 290 133 296 134
rect 159 131 163 132
rect 168 131 179 132
rect 184 131 188 132
rect 193 131 195 132
rect 200 131 204 132
rect 209 131 221 132
rect 150 130 154 131
rect 160 130 162 131
rect 150 127 153 130
rect 167 129 180 131
rect 185 130 187 131
rect 192 129 195 131
rect 166 128 181 129
rect 191 128 195 129
rect 104 126 153 127
rect 3 125 98 126
rect 103 125 153 126
rect 157 127 159 128
rect 164 127 182 128
rect 189 127 195 128
rect 199 127 204 131
rect 208 127 220 131
rect 224 127 227 132
rect 233 130 235 132
rect 232 128 235 130
rect 231 127 235 128
rect 239 127 245 133
rect 253 131 258 133
rect 262 132 269 133
rect 262 131 267 132
rect 274 131 277 133
rect 281 132 298 133
rect 304 132 307 134
rect 312 132 313 133
rect 317 132 409 135
rect 281 131 291 132
rect 295 131 300 132
rect 252 130 258 131
rect 273 130 277 131
rect 282 130 285 131
rect 252 129 257 130
rect 272 129 278 130
rect 289 129 291 131
rect 296 130 299 131
rect 304 130 306 132
rect 311 131 314 132
rect 251 127 257 129
rect 271 128 279 129
rect 288 128 292 129
rect 303 128 306 130
rect 269 127 280 128
rect 287 127 294 128
rect 301 127 306 128
rect 310 128 314 131
rect 318 128 409 132
rect 310 127 315 128
rect 319 127 409 128
rect 157 126 245 127
rect 157 125 244 126
rect 250 125 409 127
rect 3 122 95 125
rect 102 123 152 125
rect 157 124 241 125
rect 249 124 409 125
rect 100 122 152 123
rect 156 122 241 124
rect 248 123 409 124
rect 247 122 409 123
rect 3 109 409 122
rect 3 108 84 109
rect 90 108 97 109
rect 102 108 108 109
rect 113 108 119 109
rect 128 108 138 109
rect 143 108 164 109
rect 3 107 83 108
rect 91 107 96 108
rect 103 107 107 108
rect 114 107 119 108
rect 127 107 137 108
rect 144 107 164 108
rect 3 105 82 107
rect 86 105 88 107
rect 3 103 88 105
rect 92 106 95 107
rect 92 104 94 106
rect 98 105 100 107
rect 103 106 106 107
rect 110 106 111 107
rect 115 106 119 107
rect 92 103 93 104
rect 3 102 87 103
rect 3 101 86 102
rect 91 101 93 103
rect 97 102 100 105
rect 3 100 85 101
rect 90 100 93 101
rect 3 99 84 100
rect 89 99 93 100
rect 3 98 83 99
rect 88 98 93 99
rect 3 96 82 98
rect 87 97 93 98
rect 86 96 93 97
rect 96 99 100 102
rect 104 105 106 106
rect 109 105 112 106
rect 104 104 112 105
rect 104 103 111 104
rect 104 102 110 103
rect 115 102 118 106
rect 122 105 136 107
rect 140 106 141 107
rect 145 106 164 107
rect 167 106 176 109
rect 181 107 185 109
rect 190 108 208 109
rect 215 108 221 109
rect 190 107 207 108
rect 216 107 221 108
rect 224 107 234 109
rect 237 108 259 109
rect 237 107 258 108
rect 139 105 142 106
rect 121 104 142 105
rect 145 105 163 106
rect 145 104 148 105
rect 151 104 152 105
rect 155 104 157 105
rect 162 104 163 105
rect 167 104 175 106
rect 181 105 184 107
rect 190 106 206 107
rect 190 105 205 106
rect 210 105 213 106
rect 125 103 141 104
rect 145 103 147 104
rect 155 103 156 104
rect 126 102 139 103
rect 144 102 147 103
rect 154 102 156 103
rect 159 102 161 103
rect 166 102 175 104
rect 104 101 109 102
rect 114 101 117 102
rect 121 101 123 102
rect 103 100 108 101
rect 113 100 123 101
rect 127 101 139 102
rect 143 101 147 102
rect 152 101 155 102
rect 127 100 140 101
rect 103 99 107 100
rect 113 99 124 100
rect 96 97 99 99
rect 103 98 106 99
rect 112 98 116 99
rect 102 97 106 98
rect 111 97 116 98
rect 120 97 123 99
rect 127 98 141 100
rect 96 96 98 97
rect 102 96 105 97
rect 110 96 117 97
rect 120 96 122 97
rect 126 96 134 98
rect 137 97 141 98
rect 144 99 147 101
rect 151 100 155 101
rect 144 97 146 99
rect 150 97 154 100
rect 158 97 162 102
rect 166 99 174 102
rect 165 97 174 99
rect 177 97 178 104
rect 181 102 183 105
rect 181 100 182 102
rect 185 100 186 102
rect 189 100 192 105
rect 195 103 199 105
rect 203 104 204 105
rect 195 101 198 103
rect 202 102 204 104
rect 208 104 214 105
rect 217 104 220 107
rect 224 106 258 107
rect 223 105 258 106
rect 223 104 224 105
rect 229 104 233 105
rect 208 103 220 104
rect 207 102 220 103
rect 224 102 226 103
rect 184 98 185 100
rect 189 99 193 100
rect 196 99 197 101
rect 201 100 203 102
rect 200 99 203 100
rect 207 99 219 102
rect 223 100 226 102
rect 230 102 233 104
rect 236 102 239 105
rect 242 104 243 105
rect 247 104 258 105
rect 264 107 268 109
rect 264 105 267 107
rect 273 106 276 109
rect 286 108 289 109
rect 287 107 289 108
rect 288 106 289 107
rect 293 107 297 109
rect 301 107 306 109
rect 310 108 409 109
rect 248 103 258 104
rect 243 102 245 103
rect 230 101 232 102
rect 236 101 238 102
rect 138 96 140 97
rect 3 94 81 96
rect 91 95 94 96
rect 101 95 105 96
rect 114 95 117 96
rect 125 95 135 96
rect 143 95 146 97
rect 90 94 95 95
rect 100 94 104 95
rect 114 94 118 95
rect 124 94 136 95
rect 141 94 146 95
rect 149 95 155 97
rect 159 96 161 97
rect 165 95 173 97
rect 149 94 156 95
rect 164 94 173 95
rect 176 96 178 97
rect 176 94 179 96
rect 183 95 185 98
rect 182 94 184 95
rect 188 94 193 99
rect 200 98 204 99
rect 207 98 213 99
rect 199 97 204 98
rect 208 97 211 98
rect 216 97 219 99
rect 222 97 226 100
rect 229 97 232 101
rect 235 98 238 101
rect 242 100 246 102
rect 241 99 246 100
rect 198 96 204 97
rect 215 96 218 97
rect 222 96 225 97
rect 229 96 231 97
rect 235 96 237 98
rect 241 97 245 99
rect 249 98 257 103
rect 260 98 261 104
rect 264 103 266 105
rect 272 104 276 106
rect 279 105 284 106
rect 279 104 285 105
rect 264 101 265 103
rect 268 101 269 103
rect 272 101 275 104
rect 279 103 284 104
rect 288 103 290 106
rect 279 102 283 103
rect 287 101 290 103
rect 293 105 296 107
rect 301 105 305 107
rect 309 106 409 108
rect 293 103 295 105
rect 301 103 304 105
rect 308 104 409 106
rect 293 101 294 103
rect 298 102 299 103
rect 267 98 268 100
rect 249 97 256 98
rect 242 96 244 97
rect 248 96 256 97
rect 198 95 205 96
rect 214 95 218 96
rect 3 93 193 94
rect 197 94 206 95
rect 213 94 218 95
rect 221 94 225 96
rect 228 94 231 96
rect 234 94 237 96
rect 247 95 256 96
rect 197 93 237 94
rect 240 94 241 95
rect 246 94 256 95
rect 259 94 261 98
rect 266 96 268 98
rect 271 99 275 101
rect 286 100 290 101
rect 297 100 299 102
rect 302 101 303 103
rect 307 102 409 104
rect 306 100 409 102
rect 285 99 290 100
rect 265 94 267 96
rect 271 95 274 99
rect 278 97 290 99
rect 296 98 299 100
rect 305 98 409 100
rect 270 94 274 95
rect 277 94 290 97
rect 295 96 299 98
rect 304 96 409 98
rect 294 94 299 96
rect 303 94 409 96
rect 3 92 192 93
rect 3 90 190 92
rect 196 91 236 93
rect 240 91 409 94
rect 195 90 236 91
rect 239 90 409 91
rect 3 2 409 90
<< metal3 >>
rect 5 286 411 358
rect 5 255 55 286
rect 61 274 74 286
rect 61 255 74 269
rect 80 255 86 286
rect 92 285 117 286
rect 128 285 152 286
rect 92 284 115 285
rect 130 284 152 285
rect 92 283 114 284
rect 132 283 152 284
rect 92 282 113 283
rect 92 280 112 282
rect 133 281 152 283
rect 174 281 178 286
rect 120 280 125 281
rect 92 276 111 280
rect 118 279 127 280
rect 118 277 128 279
rect 134 278 152 281
rect 135 277 152 278
rect 119 276 152 277
rect 92 274 112 276
rect 121 275 152 276
rect 125 274 152 275
rect 92 272 113 274
rect 129 273 152 274
rect 159 273 178 281
rect 131 272 152 273
rect 92 271 114 272
rect 132 271 152 272
rect 92 270 116 271
rect 133 270 152 271
rect 92 269 118 270
rect 134 269 152 270
rect 92 268 122 269
rect 92 267 125 268
rect 92 266 128 267
rect 92 265 112 266
rect 92 263 110 265
rect 117 263 129 266
rect 92 260 111 263
rect 118 262 128 263
rect 119 261 128 262
rect 121 260 125 261
rect 135 260 152 269
rect 172 268 178 273
rect 108 259 112 260
rect 134 259 152 260
rect 108 258 113 259
rect 133 258 152 259
rect 108 257 114 258
rect 132 257 152 258
rect 108 256 115 257
rect 131 256 152 257
rect 108 255 117 256
rect 129 255 152 256
rect 159 255 178 268
rect 185 255 190 286
rect 210 285 233 286
rect 212 284 233 285
rect 213 283 233 284
rect 214 281 233 283
rect 254 281 259 286
rect 265 281 271 286
rect 196 280 206 281
rect 196 278 208 280
rect 196 276 209 278
rect 196 274 208 276
rect 196 273 206 274
rect 215 273 233 281
rect 239 278 271 281
rect 239 273 259 278
rect 214 272 233 273
rect 213 271 233 272
rect 212 270 233 271
rect 211 269 233 270
rect 208 268 233 269
rect 252 268 259 273
rect 196 267 200 268
rect 209 267 233 268
rect 196 266 202 267
rect 210 266 233 267
rect 196 265 203 266
rect 211 265 233 266
rect 196 263 204 265
rect 212 264 233 265
rect 196 262 205 263
rect 213 262 233 264
rect 196 260 206 262
rect 214 261 233 262
rect 196 259 207 260
rect 215 259 233 261
rect 196 257 208 259
rect 216 257 233 259
rect 196 256 209 257
rect 217 256 233 257
rect 196 255 210 256
rect 218 255 233 256
rect 239 255 259 268
rect 265 255 271 278
rect 277 285 411 286
rect 277 284 288 285
rect 277 283 286 284
rect 277 282 284 283
rect 277 278 283 282
rect 289 279 411 285
rect 289 278 302 279
rect 309 278 329 279
rect 334 278 411 279
rect 277 273 280 278
rect 293 277 300 278
rect 311 277 320 278
rect 293 275 298 277
rect 313 275 320 277
rect 326 277 328 278
rect 326 276 327 277
rect 335 276 411 278
rect 293 274 297 275
rect 314 274 320 275
rect 334 274 411 276
rect 293 273 296 274
rect 304 273 307 274
rect 277 257 283 273
rect 289 272 296 273
rect 303 272 309 273
rect 289 262 295 272
rect 302 271 309 272
rect 315 271 320 274
rect 333 273 411 274
rect 329 272 411 273
rect 328 271 411 272
rect 302 270 310 271
rect 301 269 310 270
rect 316 265 320 271
rect 301 264 320 265
rect 302 262 320 264
rect 289 261 296 262
rect 303 261 309 262
rect 314 261 320 262
rect 290 260 292 261
rect 293 260 296 261
rect 304 260 308 261
rect 293 258 297 260
rect 315 259 320 261
rect 314 258 320 259
rect 294 257 298 258
rect 313 257 320 258
rect 277 256 284 257
rect 294 256 300 257
rect 312 256 320 257
rect 277 255 286 256
rect 293 255 301 256
rect 310 255 320 256
rect 327 255 411 271
rect 5 230 411 255
rect 5 224 70 230
rect 74 229 84 230
rect 88 229 89 230
rect 74 227 83 229
rect 87 227 89 229
rect 93 229 106 230
rect 93 228 100 229
rect 93 227 99 228
rect 101 227 105 229
rect 110 228 137 230
rect 109 227 136 228
rect 74 226 82 227
rect 86 226 98 227
rect 75 224 81 226
rect 86 225 97 226
rect 101 225 136 227
rect 141 226 148 230
rect 153 229 156 230
rect 152 227 156 229
rect 160 229 175 230
rect 182 229 222 230
rect 230 229 319 230
rect 326 229 411 230
rect 160 228 173 229
rect 184 228 221 229
rect 231 228 271 229
rect 272 228 317 229
rect 327 228 411 229
rect 5 219 71 224
rect 75 222 80 224
rect 85 223 88 225
rect 75 220 79 222
rect 84 221 88 223
rect 92 222 94 225
rect 103 224 105 225
rect 109 224 114 225
rect 121 224 136 225
rect 103 223 104 224
rect 109 223 112 224
rect 122 223 136 224
rect 102 222 104 223
rect 5 213 72 219
rect 76 218 78 220
rect 83 219 87 221
rect 92 220 96 222
rect 100 220 104 222
rect 76 216 77 218
rect 82 217 87 219
rect 81 216 87 217
rect 91 216 95 220
rect 99 219 104 220
rect 80 214 86 216
rect 91 215 94 216
rect 99 215 103 219
rect 108 218 111 223
rect 115 221 118 222
rect 115 220 119 221
rect 123 220 135 223
rect 140 222 147 226
rect 152 224 155 227
rect 160 226 172 228
rect 185 227 220 228
rect 232 227 269 228
rect 272 227 316 228
rect 328 227 411 228
rect 177 226 180 227
rect 185 226 219 227
rect 224 226 227 227
rect 233 226 268 227
rect 271 226 315 227
rect 160 225 171 226
rect 151 222 155 224
rect 159 222 171 225
rect 175 225 181 226
rect 186 225 219 226
rect 175 224 182 225
rect 186 224 195 225
rect 199 224 204 225
rect 176 223 196 224
rect 178 222 196 223
rect 200 222 203 224
rect 209 223 219 225
rect 223 224 229 226
rect 233 225 267 226
rect 271 225 314 226
rect 321 225 324 226
rect 329 225 411 227
rect 233 224 235 225
rect 224 223 235 224
rect 208 222 219 223
rect 226 222 235 223
rect 118 219 135 220
rect 151 219 154 222
rect 159 221 172 222
rect 180 221 196 222
rect 201 221 202 222
rect 207 221 219 222
rect 228 221 235 222
rect 239 223 245 225
rect 249 224 253 225
rect 260 224 265 225
rect 273 224 277 225
rect 283 224 290 225
rect 294 224 295 225
rect 300 224 303 225
rect 308 224 313 225
rect 319 224 325 225
rect 249 223 251 224
rect 261 223 264 224
rect 239 221 244 223
rect 248 222 251 223
rect 262 222 264 223
rect 273 223 276 224
rect 285 223 290 224
rect 301 223 302 224
rect 309 223 313 224
rect 318 223 326 224
rect 330 223 411 225
rect 273 222 275 223
rect 285 222 289 223
rect 248 221 250 222
rect 255 221 257 222
rect 263 221 266 222
rect 159 220 173 221
rect 182 220 197 221
rect 206 220 220 221
rect 230 220 236 221
rect 120 218 125 219
rect 132 218 135 219
rect 5 210 73 213
rect 79 212 86 214
rect 78 211 86 212
rect 90 211 94 215
rect 98 214 103 215
rect 107 217 112 218
rect 121 217 124 218
rect 107 216 114 217
rect 107 215 117 216
rect 122 215 124 217
rect 132 215 134 218
rect 139 216 146 218
rect 98 213 102 214
rect 107 213 109 215
rect 113 214 118 215
rect 114 213 117 214
rect 122 213 134 215
rect 138 215 146 216
rect 150 217 154 219
rect 158 219 174 220
rect 183 219 197 220
rect 205 219 222 220
rect 158 218 176 219
rect 158 217 178 218
rect 184 217 198 219
rect 204 218 224 219
rect 231 218 236 220
rect 203 217 226 218
rect 101 211 102 213
rect 78 210 85 211
rect 90 210 95 211
rect 100 210 102 211
rect 106 212 109 213
rect 122 212 133 213
rect 106 211 110 212
rect 121 211 133 212
rect 138 211 145 215
rect 150 213 153 217
rect 158 216 180 217
rect 158 215 169 216
rect 173 215 180 216
rect 157 214 169 215
rect 174 214 180 215
rect 184 215 197 217
rect 203 216 227 217
rect 184 214 196 215
rect 204 214 217 216
rect 221 214 228 216
rect 232 215 236 218
rect 240 219 243 221
rect 247 219 250 221
rect 254 220 259 221
rect 262 220 266 221
rect 257 219 266 220
rect 240 218 242 219
rect 246 218 250 219
rect 259 218 266 219
rect 270 220 274 222
rect 279 221 281 222
rect 240 215 241 218
rect 246 217 251 218
rect 245 216 253 217
rect 261 216 265 218
rect 270 217 273 220
rect 278 219 282 221
rect 277 218 283 219
rect 286 218 289 222
rect 295 221 297 222
rect 303 221 305 222
rect 294 220 297 221
rect 245 215 256 216
rect 232 214 237 215
rect 106 210 112 211
rect 119 210 133 211
rect 137 210 145 211
rect 149 212 153 213
rect 167 213 169 214
rect 175 213 179 214
rect 184 213 195 214
rect 167 212 170 213
rect 183 212 194 213
rect 199 212 201 213
rect 205 212 217 214
rect 222 213 226 214
rect 231 212 237 214
rect 244 213 248 215
rect 252 214 257 215
rect 262 214 265 216
rect 253 213 257 214
rect 149 210 152 212
rect 167 211 171 212
rect 182 211 193 212
rect 198 211 201 212
rect 206 211 218 212
rect 230 211 237 212
rect 243 211 249 213
rect 261 212 264 214
rect 269 213 273 217
rect 286 216 288 218
rect 293 217 297 220
rect 302 219 306 221
rect 277 214 288 216
rect 278 213 281 214
rect 271 212 274 213
rect 285 212 288 214
rect 292 216 297 217
rect 292 212 296 216
rect 301 215 305 219
rect 310 218 312 223
rect 317 221 411 223
rect 260 211 265 212
rect 167 210 173 211
rect 181 210 192 211
rect 197 210 202 211
rect 206 210 220 211
rect 228 210 237 211
rect 5 209 237 210
rect 242 210 251 211
rect 259 210 265 211
rect 271 211 275 212
rect 284 211 287 212
rect 271 210 276 211
rect 283 210 287 211
rect 291 211 296 212
rect 300 214 305 215
rect 309 214 312 218
rect 316 217 411 221
rect 316 216 324 217
rect 317 215 323 216
rect 318 214 322 215
rect 328 214 411 217
rect 291 210 295 211
rect 300 210 304 214
rect 309 213 313 214
rect 327 213 411 214
rect 308 212 314 213
rect 326 212 411 213
rect 308 211 315 212
rect 325 211 411 212
rect 308 210 316 211
rect 323 210 411 211
rect 242 209 411 210
rect 5 208 236 209
rect 5 205 233 208
rect 241 207 411 209
rect 240 206 411 207
rect 239 205 411 206
rect 5 145 411 205
rect 5 141 79 145
rect 85 143 91 145
rect 97 144 120 145
rect 127 144 135 145
rect 97 143 118 144
rect 129 143 135 144
rect 5 136 78 141
rect 85 140 90 143
rect 97 142 117 143
rect 97 141 116 142
rect 130 141 135 143
rect 139 142 151 145
rect 156 144 226 145
rect 155 143 226 144
rect 232 144 238 145
rect 155 142 225 143
rect 139 141 225 142
rect 97 140 115 141
rect 122 140 125 141
rect 5 131 77 136
rect 81 133 82 139
rect 85 138 89 140
rect 86 136 88 138
rect 86 134 87 136
rect 91 134 92 136
rect 96 135 99 140
rect 103 139 109 140
rect 113 139 115 140
rect 120 139 127 140
rect 103 137 108 139
rect 113 138 114 139
rect 103 135 107 137
rect 112 136 114 138
rect 119 138 127 139
rect 131 138 134 141
rect 138 140 225 141
rect 138 139 140 140
rect 145 139 150 140
rect 155 139 158 140
rect 162 139 163 140
rect 168 139 186 140
rect 192 139 199 140
rect 138 138 139 139
rect 119 137 134 138
rect 146 137 150 139
rect 96 134 100 135
rect 5 126 76 131
rect 80 127 82 133
rect 90 133 92 134
rect 90 132 91 133
rect 89 129 91 132
rect 88 128 91 129
rect 95 128 100 134
rect 104 133 106 135
rect 111 134 114 136
rect 104 131 105 133
rect 110 132 114 134
rect 109 130 114 132
rect 118 136 134 137
rect 140 136 142 137
rect 118 132 133 136
rect 138 134 142 136
rect 147 135 150 137
rect 154 138 158 139
rect 169 138 184 139
rect 194 138 199 139
rect 203 139 205 140
rect 210 139 225 140
rect 203 138 204 139
rect 211 138 225 139
rect 232 142 237 144
rect 244 143 263 145
rect 274 144 311 145
rect 316 144 411 145
rect 275 143 311 144
rect 232 139 236 142
rect 243 140 262 143
rect 276 142 311 143
rect 118 131 126 132
rect 130 131 133 132
rect 137 131 142 134
rect 118 130 125 131
rect 130 130 132 131
rect 137 130 141 131
rect 146 130 149 135
rect 154 134 157 138
rect 170 137 183 138
rect 163 136 165 137
rect 170 136 182 137
rect 188 136 190 137
rect 162 135 166 136
rect 171 135 182 136
rect 186 135 191 136
rect 195 135 199 138
rect 205 136 207 137
rect 204 135 208 136
rect 153 133 157 134
rect 161 133 167 135
rect 171 134 181 135
rect 108 128 114 130
rect 120 129 123 130
rect 129 128 132 130
rect 88 127 90 128
rect 5 125 75 126
rect 79 125 83 127
rect 87 125 90 127
rect 94 125 101 128
rect 107 127 115 128
rect 128 127 132 128
rect 107 126 116 127
rect 127 126 132 127
rect 136 126 141 130
rect 5 124 101 125
rect 106 125 118 126
rect 125 125 131 126
rect 136 125 140 126
rect 145 125 148 130
rect 153 129 156 133
rect 161 132 166 133
rect 171 132 172 134
rect 180 133 181 134
rect 186 133 192 135
rect 160 131 166 132
rect 161 130 166 131
rect 170 130 171 131
rect 179 130 181 133
rect 185 130 191 133
rect 196 132 198 135
rect 203 134 208 135
rect 212 134 224 138
rect 232 137 235 139
rect 243 138 245 140
rect 249 138 255 140
rect 260 139 262 140
rect 259 138 262 139
rect 266 140 271 141
rect 277 140 311 142
rect 315 140 411 144
rect 243 137 246 138
rect 203 133 207 134
rect 195 130 198 132
rect 202 130 207 133
rect 211 130 213 134
rect 221 133 224 134
rect 227 135 228 136
rect 232 135 234 137
rect 238 135 239 137
rect 221 131 223 133
rect 220 130 223 131
rect 227 130 229 135
rect 232 133 233 135
rect 237 133 238 135
rect 236 130 238 133
rect 242 132 246 137
rect 250 136 254 138
rect 259 137 261 138
rect 250 134 253 136
rect 258 135 261 137
rect 266 136 273 140
rect 277 139 283 140
rect 289 139 297 140
rect 305 139 310 140
rect 315 139 318 140
rect 323 139 411 140
rect 250 132 252 134
rect 257 133 261 135
rect 265 133 273 136
rect 278 138 282 139
rect 291 138 296 139
rect 306 138 310 139
rect 278 137 281 138
rect 291 137 295 138
rect 278 135 280 137
rect 285 136 287 137
rect 278 134 279 135
rect 284 134 288 136
rect 242 131 247 132
rect 250 131 251 132
rect 256 131 260 133
rect 265 131 272 133
rect 277 131 279 134
rect 283 133 289 134
rect 292 133 295 137
rect 299 136 302 137
rect 299 135 303 136
rect 307 135 310 138
rect 314 138 317 139
rect 322 138 411 139
rect 314 137 316 138
rect 321 137 411 138
rect 314 136 315 137
rect 320 136 411 137
rect 319 135 411 136
rect 301 134 309 135
rect 304 133 309 134
rect 318 133 411 135
rect 292 132 296 133
rect 305 132 309 133
rect 292 131 298 132
rect 161 129 165 130
rect 170 129 181 130
rect 186 129 190 130
rect 195 129 197 130
rect 202 129 206 130
rect 211 129 223 130
rect 152 128 156 129
rect 162 128 164 129
rect 152 125 155 128
rect 169 127 182 129
rect 187 128 189 129
rect 194 127 197 129
rect 168 126 183 127
rect 193 126 197 127
rect 106 124 155 125
rect 5 123 100 124
rect 105 123 155 124
rect 159 125 161 126
rect 166 125 184 126
rect 191 125 197 126
rect 201 125 206 129
rect 210 125 222 129
rect 226 125 229 130
rect 235 128 237 130
rect 234 126 237 128
rect 233 125 237 126
rect 241 125 247 131
rect 255 129 260 131
rect 264 130 271 131
rect 264 129 269 130
rect 276 129 279 131
rect 283 130 300 131
rect 306 130 309 132
rect 314 130 315 131
rect 319 130 411 133
rect 283 129 293 130
rect 297 129 302 130
rect 254 128 260 129
rect 275 128 279 129
rect 284 128 287 129
rect 254 127 259 128
rect 274 127 280 128
rect 291 127 293 129
rect 298 128 301 129
rect 306 128 308 130
rect 313 129 316 130
rect 253 125 259 127
rect 273 126 281 127
rect 290 126 294 127
rect 305 126 308 128
rect 271 125 282 126
rect 289 125 296 126
rect 303 125 308 126
rect 312 126 316 129
rect 320 126 411 130
rect 312 125 317 126
rect 321 125 411 126
rect 159 124 247 125
rect 159 123 246 124
rect 252 123 411 125
rect 5 120 97 123
rect 104 121 154 123
rect 159 122 243 123
rect 251 122 411 123
rect 102 120 154 121
rect 158 120 243 122
rect 250 121 411 122
rect 249 120 411 121
rect 5 107 411 120
rect 5 106 86 107
rect 92 106 99 107
rect 104 106 110 107
rect 115 106 121 107
rect 130 106 140 107
rect 145 106 166 107
rect 5 105 85 106
rect 93 105 98 106
rect 105 105 109 106
rect 116 105 121 106
rect 129 105 139 106
rect 146 105 166 106
rect 5 103 84 105
rect 88 103 90 105
rect 5 101 90 103
rect 94 104 97 105
rect 94 102 96 104
rect 100 103 102 105
rect 105 104 108 105
rect 112 104 113 105
rect 117 104 121 105
rect 94 101 95 102
rect 5 100 89 101
rect 5 99 88 100
rect 93 99 95 101
rect 99 100 102 103
rect 5 98 87 99
rect 92 98 95 99
rect 5 97 86 98
rect 91 97 95 98
rect 5 96 85 97
rect 90 96 95 97
rect 5 94 84 96
rect 89 95 95 96
rect 88 94 95 95
rect 98 97 102 100
rect 106 103 108 104
rect 111 103 114 104
rect 106 102 114 103
rect 106 101 113 102
rect 106 100 112 101
rect 117 100 120 104
rect 124 103 138 105
rect 142 104 143 105
rect 147 104 166 105
rect 169 104 178 107
rect 183 105 187 107
rect 192 106 210 107
rect 217 106 223 107
rect 192 105 209 106
rect 218 105 223 106
rect 226 105 236 107
rect 239 106 261 107
rect 239 105 260 106
rect 141 103 144 104
rect 123 102 144 103
rect 147 103 165 104
rect 147 102 150 103
rect 153 102 154 103
rect 157 102 159 103
rect 164 102 165 103
rect 169 102 177 104
rect 183 103 186 105
rect 192 104 208 105
rect 192 103 207 104
rect 212 103 215 104
rect 127 101 143 102
rect 147 101 149 102
rect 157 101 158 102
rect 128 100 141 101
rect 146 100 149 101
rect 156 100 158 101
rect 161 100 163 101
rect 168 100 177 102
rect 106 99 111 100
rect 116 99 119 100
rect 123 99 125 100
rect 105 98 110 99
rect 115 98 125 99
rect 129 99 141 100
rect 145 99 149 100
rect 154 99 157 100
rect 129 98 142 99
rect 105 97 109 98
rect 115 97 126 98
rect 98 95 101 97
rect 105 96 108 97
rect 114 96 118 97
rect 104 95 108 96
rect 113 95 118 96
rect 122 95 125 97
rect 129 96 143 98
rect 98 94 100 95
rect 104 94 107 95
rect 112 94 119 95
rect 122 94 124 95
rect 128 94 136 96
rect 139 95 143 96
rect 146 97 149 99
rect 153 98 157 99
rect 146 95 148 97
rect 152 95 156 98
rect 160 95 164 100
rect 168 97 176 100
rect 167 95 176 97
rect 179 95 180 102
rect 183 100 185 103
rect 183 98 184 100
rect 187 98 188 100
rect 191 98 194 103
rect 197 101 201 103
rect 205 102 206 103
rect 197 99 200 101
rect 204 100 206 102
rect 210 102 216 103
rect 219 102 222 105
rect 226 104 260 105
rect 225 103 260 104
rect 225 102 226 103
rect 231 102 235 103
rect 210 101 222 102
rect 209 100 222 101
rect 226 100 228 101
rect 186 96 187 98
rect 191 97 195 98
rect 198 97 199 99
rect 203 98 205 100
rect 202 97 205 98
rect 209 97 221 100
rect 225 98 228 100
rect 232 100 235 102
rect 238 100 241 103
rect 244 102 245 103
rect 249 102 260 103
rect 266 105 270 107
rect 266 103 269 105
rect 275 104 278 107
rect 288 106 291 107
rect 289 105 291 106
rect 290 104 291 105
rect 295 105 299 107
rect 303 105 308 107
rect 312 106 411 107
rect 250 101 260 102
rect 245 100 247 101
rect 232 99 234 100
rect 238 99 240 100
rect 140 94 142 95
rect 5 92 83 94
rect 93 93 96 94
rect 103 93 107 94
rect 116 93 119 94
rect 127 93 137 94
rect 145 93 148 95
rect 92 92 97 93
rect 102 92 106 93
rect 116 92 120 93
rect 126 92 138 93
rect 143 92 148 93
rect 151 93 157 95
rect 161 94 163 95
rect 167 93 175 95
rect 151 92 158 93
rect 166 92 175 93
rect 178 94 180 95
rect 178 92 181 94
rect 185 93 187 96
rect 184 92 186 93
rect 190 92 195 97
rect 202 96 206 97
rect 209 96 215 97
rect 201 95 206 96
rect 210 95 213 96
rect 218 95 221 97
rect 224 95 228 98
rect 231 95 234 99
rect 237 96 240 99
rect 244 98 248 100
rect 243 97 248 98
rect 200 94 206 95
rect 217 94 220 95
rect 224 94 227 95
rect 231 94 233 95
rect 237 94 239 96
rect 243 95 247 97
rect 251 96 259 101
rect 262 96 263 102
rect 266 101 268 103
rect 274 102 278 104
rect 281 103 286 104
rect 281 102 287 103
rect 266 99 267 101
rect 270 99 271 101
rect 274 99 277 102
rect 281 101 286 102
rect 290 101 292 104
rect 281 100 285 101
rect 289 99 292 101
rect 295 103 298 105
rect 303 103 307 105
rect 311 104 411 106
rect 295 101 297 103
rect 303 101 306 103
rect 310 102 411 104
rect 295 99 296 101
rect 300 100 301 101
rect 269 96 270 98
rect 251 95 258 96
rect 244 94 246 95
rect 250 94 258 95
rect 200 93 207 94
rect 216 93 220 94
rect 5 91 195 92
rect 199 92 208 93
rect 215 92 220 93
rect 223 92 227 94
rect 230 92 233 94
rect 236 92 239 94
rect 249 93 258 94
rect 199 91 239 92
rect 242 92 243 93
rect 248 92 258 93
rect 261 92 263 96
rect 268 94 270 96
rect 273 97 277 99
rect 288 98 292 99
rect 299 98 301 100
rect 304 99 305 101
rect 309 100 411 102
rect 308 98 411 100
rect 287 97 292 98
rect 267 92 269 94
rect 273 93 276 97
rect 280 95 292 97
rect 298 96 301 98
rect 307 96 411 98
rect 272 92 276 93
rect 279 92 292 95
rect 297 94 301 96
rect 306 94 411 96
rect 296 92 301 94
rect 305 92 411 94
rect 5 90 194 91
rect 5 88 192 90
rect 198 89 238 91
rect 242 89 411 92
rect 197 88 238 89
rect 241 88 411 89
rect 5 0 411 88
<< end >>
