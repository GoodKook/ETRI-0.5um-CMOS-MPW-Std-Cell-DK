magic
tech scmos
magscale 1 6
timestamp 1725342160
<< nwell >>
rect 0 0 176 260
<< ptransistor >>
rect 65 30 75 230
<< ndiffusion >>
rect 134 190 166 226
rect 134 178 144 190
rect 156 178 166 190
rect 134 134 166 178
rect 134 122 144 134
rect 156 122 166 134
rect 134 78 166 122
rect 134 66 144 78
rect 156 66 166 78
rect 134 30 166 66
<< pdiffusion >>
rect 28 220 65 230
rect 28 208 38 220
rect 50 208 65 220
rect 28 196 65 208
rect 28 184 38 196
rect 50 184 65 196
rect 28 172 65 184
rect 28 160 38 172
rect 50 160 65 172
rect 28 148 65 160
rect 28 136 38 148
rect 50 136 65 148
rect 28 124 65 136
rect 28 112 38 124
rect 50 112 65 124
rect 28 100 65 112
rect 28 88 38 100
rect 50 88 65 100
rect 28 76 65 88
rect 28 64 38 76
rect 50 64 65 76
rect 28 52 65 64
rect 28 40 38 52
rect 50 40 65 52
rect 28 30 65 40
rect 75 220 112 230
rect 75 208 90 220
rect 102 208 112 220
rect 75 196 112 208
rect 75 184 90 196
rect 102 184 112 196
rect 75 172 112 184
rect 75 160 90 172
rect 102 160 112 172
rect 75 148 112 160
rect 75 136 90 148
rect 102 136 112 148
rect 75 124 112 136
rect 75 112 90 124
rect 102 112 112 124
rect 75 100 112 112
rect 75 88 90 100
rect 102 88 112 100
rect 75 76 112 88
rect 75 64 90 76
rect 102 64 112 76
rect 75 52 112 64
rect 75 40 90 52
rect 102 40 112 52
rect 75 30 112 40
<< ndcontact >>
rect 144 178 156 190
rect 144 122 156 134
rect 144 66 156 78
<< pdcontact >>
rect 38 208 50 220
rect 38 184 50 196
rect 38 160 50 172
rect 38 136 50 148
rect 38 112 50 124
rect 38 88 50 100
rect 38 64 50 76
rect 38 40 50 52
rect 90 208 102 220
rect 90 184 102 196
rect 90 160 102 172
rect 90 136 102 148
rect 90 112 102 124
rect 90 88 102 100
rect 90 64 102 76
rect 90 40 102 52
<< polysilicon >>
rect 54 278 86 282
rect 54 254 58 278
rect 82 254 86 278
rect 54 250 86 254
rect 65 230 75 250
rect 65 20 75 30
<< polycontact >>
rect 58 254 82 278
<< metal1 >>
rect 52 278 88 284
rect 52 254 58 278
rect 82 254 88 278
rect 52 248 88 254
rect 26 220 62 232
rect 26 208 38 220
rect 50 208 62 220
rect 26 196 62 208
rect 26 184 38 196
rect 50 184 62 196
rect 26 172 62 184
rect 26 160 38 172
rect 50 160 62 172
rect 26 148 62 160
rect 26 136 38 148
rect 50 136 62 148
rect 26 124 62 136
rect 26 112 38 124
rect 50 112 62 124
rect 26 100 62 112
rect 26 88 38 100
rect 50 88 62 100
rect 26 76 62 88
rect 26 64 38 76
rect 50 64 62 76
rect 26 52 62 64
rect 26 40 38 52
rect 50 40 62 52
rect 26 28 62 40
rect 78 220 114 232
rect 78 208 90 220
rect 102 208 114 220
rect 78 196 114 208
rect 78 184 90 196
rect 102 184 114 196
rect 78 172 114 184
rect 78 160 90 172
rect 102 160 114 172
rect 78 148 114 160
rect 78 136 90 148
rect 102 136 114 148
rect 78 124 114 136
rect 78 112 90 124
rect 102 112 114 124
rect 78 100 114 112
rect 78 88 90 100
rect 102 88 114 100
rect 78 76 114 88
rect 78 64 90 76
rect 102 64 114 76
rect 78 52 114 64
rect 78 40 90 52
rect 102 40 114 52
rect 78 28 114 40
rect 132 190 168 228
rect 132 178 144 190
rect 156 178 168 190
rect 132 134 168 178
rect 132 122 144 134
rect 156 122 168 134
rect 132 78 168 122
rect 132 66 144 78
rect 156 66 168 78
rect 132 28 168 66
<< end >>
