magic
tech scmos
magscale 1 2
timestamp 1727267527
<< nwell >>
rect -12 154 92 272
<< ntransistor >>
rect 22 14 26 54
rect 32 14 36 54
<< ptransistor >>
rect 20 206 24 246
rect 40 206 44 246
<< ndiffusion >>
rect 20 14 22 54
rect 26 14 32 54
rect 36 14 42 54
<< pdiffusion >>
rect 18 206 20 246
rect 24 206 26 246
rect 38 206 40 246
rect 44 206 46 246
<< ndcontact >>
rect 8 14 20 54
rect 42 14 54 54
<< pdcontact >>
rect 6 206 18 246
rect 26 206 38 246
rect 46 206 58 246
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 254 86 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 20 123 24 206
rect 16 111 24 123
rect 18 80 24 111
rect 40 80 44 206
rect 18 74 26 80
rect 22 54 26 74
rect 32 74 44 80
rect 32 54 36 74
rect 22 10 26 14
rect 32 10 36 14
<< polycontact >>
rect 4 111 16 123
rect 44 111 56 123
<< metal1 >>
rect -6 266 86 268
rect -6 252 86 254
rect 6 246 18 252
rect 46 246 58 252
rect 26 117 34 206
rect 26 68 34 103
rect 26 62 54 68
rect 42 54 54 62
rect 8 8 20 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m2contact >>
rect 3 123 17 137
rect 43 123 57 137
rect 23 103 37 117
<< metal2 >>
rect 6 137 14 154
rect 46 137 54 154
rect 26 86 34 103
<< m1p >>
rect -6 252 86 268
rect -6 -8 86 8
<< m2p >>
rect 6 137 14 154
rect 46 137 54 154
rect 26 86 34 103
<< labels >>
rlabel metal1 -6 252 66 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -6 -8 66 8 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal2 30 91 30 91 1 Y
port 3 n signal output
rlabel metal2 10 151 10 151 1 A
port 1 n signal input
rlabel metal2 50 151 50 151 1 B
port 2 n signal input
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
