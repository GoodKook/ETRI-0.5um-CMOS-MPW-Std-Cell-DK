magic
tech scmos
magscale 1 2
timestamp 1740456754
<< nwell >>
rect -2 5664 5822 5782
rect 1235 5660 1271 5664
rect 3529 5396 3565 5400
rect -2 5184 5822 5396
rect 3529 4916 3565 4920
rect 4469 4916 4505 4920
rect -2 4704 5822 4916
rect 3775 4436 3811 4440
rect 5509 4436 5545 4440
rect -2 4342 5822 4436
rect -2 4224 5823 4342
rect 695 4220 731 4224
rect 4429 4220 4465 4224
rect 3695 3956 3731 3960
rect 4629 3956 4665 3960
rect -2 3744 5822 3956
rect 2009 3740 2045 3744
rect -2 3264 5822 3476
rect 2835 2996 2871 3000
rect 3349 2996 3385 3000
rect 3795 2996 3831 3000
rect -2 2784 5822 2996
rect 1535 2780 1571 2784
rect -2 2476 3982 2516
rect 4917 2476 5822 2516
rect -2 2344 5822 2476
rect -2 2304 2062 2344
rect 2518 2304 3882 2344
rect 4338 2304 5822 2344
rect 1035 2300 1071 2304
rect 5642 2296 5717 2304
rect -2 1996 2342 2036
rect 2798 1996 5822 2036
rect -2 1864 5822 1996
rect -2 1824 2182 1864
rect 2638 1824 5822 1864
rect 3222 1816 3297 1824
rect -2 1516 1762 1556
rect 2218 1516 3062 1556
rect 3518 1516 5822 1556
rect -2 1344 5822 1516
rect -2 864 5822 1076
rect 2655 860 2691 864
rect 5235 860 5271 864
rect 2215 596 2251 600
rect -2 384 5822 596
rect 1235 380 1271 384
rect 4962 376 5037 384
rect 5322 116 5397 124
rect -2 -2 5822 116
<< ntransistor >>
rect 85 5544 89 5584
rect 105 5544 109 5584
rect 125 5544 129 5584
rect 211 5544 215 5584
rect 231 5544 235 5584
rect 251 5544 255 5584
rect 392 5544 396 5564
rect 414 5544 418 5584
rect 422 5544 426 5584
rect 512 5544 516 5604
rect 520 5544 524 5604
rect 528 5544 532 5604
rect 665 5544 669 5584
rect 685 5544 689 5584
rect 705 5544 709 5584
rect 813 5544 817 5584
rect 823 5544 827 5584
rect 932 5544 936 5564
rect 954 5544 958 5584
rect 962 5544 966 5584
rect 1071 5544 1075 5564
rect 1091 5544 1095 5564
rect 1225 5544 1229 5584
rect 1245 5544 1249 5564
rect 1265 5544 1269 5564
rect 1375 5544 1379 5584
rect 1395 5544 1399 5584
rect 1405 5544 1409 5584
rect 1528 5544 1532 5604
rect 1536 5544 1540 5604
rect 1544 5544 1548 5604
rect 1672 5544 1676 5564
rect 1694 5544 1698 5584
rect 1702 5544 1706 5584
rect 1828 5544 1832 5604
rect 1836 5544 1840 5604
rect 1844 5544 1848 5604
rect 1931 5544 1935 5564
rect 2045 5544 2049 5584
rect 2065 5544 2069 5584
rect 2085 5544 2089 5584
rect 2171 5544 2175 5584
rect 2191 5544 2195 5584
rect 2211 5544 2215 5584
rect 2314 5544 2318 5584
rect 2322 5544 2326 5584
rect 2344 5544 2348 5564
rect 2473 5544 2477 5584
rect 2483 5544 2487 5584
rect 2608 5544 2612 5604
rect 2616 5544 2620 5604
rect 2624 5544 2628 5604
rect 2748 5544 2752 5604
rect 2756 5544 2760 5604
rect 2764 5544 2768 5604
rect 2853 5544 2857 5584
rect 2863 5544 2867 5584
rect 2985 5544 2989 5564
rect 3085 5544 3089 5584
rect 3105 5544 3109 5584
rect 3125 5544 3129 5584
rect 3255 5544 3259 5584
rect 3275 5544 3279 5584
rect 3285 5544 3289 5584
rect 3385 5544 3389 5564
rect 3405 5544 3409 5564
rect 3528 5544 3532 5604
rect 3536 5544 3540 5604
rect 3544 5544 3548 5604
rect 3665 5544 3669 5564
rect 3765 5544 3769 5564
rect 3851 5544 3855 5564
rect 3951 5544 3955 5584
rect 3971 5544 3975 5584
rect 3991 5544 3995 5584
rect 4091 5544 4095 5564
rect 4151 5544 4155 5584
rect 4173 5544 4177 5564
rect 4183 5544 4187 5564
rect 4203 5544 4207 5564
rect 4211 5544 4215 5564
rect 4257 5544 4261 5564
rect 4279 5544 4283 5564
rect 4289 5544 4293 5564
rect 4311 5544 4315 5564
rect 4321 5544 4325 5564
rect 4341 5544 4345 5584
rect 4465 5544 4469 5584
rect 4485 5544 4489 5584
rect 4505 5544 4509 5584
rect 4605 5544 4609 5584
rect 4625 5544 4629 5584
rect 4645 5544 4649 5584
rect 4665 5544 4669 5584
rect 4685 5544 4689 5584
rect 4705 5544 4709 5584
rect 4725 5544 4729 5584
rect 4745 5544 4749 5584
rect 4845 5544 4849 5564
rect 4945 5544 4949 5584
rect 4965 5544 4969 5584
rect 4985 5544 4989 5584
rect 5093 5544 5097 5584
rect 5103 5544 5107 5584
rect 5193 5544 5197 5584
rect 5203 5544 5207 5584
rect 5311 5544 5315 5584
rect 5331 5544 5335 5584
rect 5351 5544 5355 5584
rect 5451 5544 5455 5564
rect 5553 5544 5557 5584
rect 5563 5544 5567 5584
rect 5671 5544 5675 5564
rect 85 5476 89 5516
rect 105 5476 109 5516
rect 125 5476 129 5516
rect 268 5456 272 5516
rect 276 5456 280 5516
rect 284 5456 288 5516
rect 408 5456 412 5516
rect 416 5456 420 5516
rect 424 5456 428 5516
rect 548 5456 552 5516
rect 556 5456 560 5516
rect 564 5456 568 5516
rect 672 5456 676 5516
rect 680 5456 684 5516
rect 688 5456 692 5516
rect 811 5476 815 5516
rect 831 5476 835 5516
rect 851 5476 855 5516
rect 952 5456 956 5516
rect 960 5456 964 5516
rect 968 5456 972 5516
rect 1112 5496 1116 5516
rect 1134 5476 1138 5516
rect 1142 5476 1146 5516
rect 1232 5456 1236 5516
rect 1240 5456 1244 5516
rect 1248 5456 1252 5516
rect 1391 5496 1395 5516
rect 1411 5496 1415 5516
rect 1548 5456 1552 5516
rect 1556 5456 1560 5516
rect 1564 5456 1568 5516
rect 1651 5476 1655 5516
rect 1671 5476 1675 5516
rect 1691 5476 1695 5516
rect 1828 5456 1832 5516
rect 1836 5456 1840 5516
rect 1844 5456 1848 5516
rect 1968 5456 1972 5516
rect 1976 5456 1980 5516
rect 1984 5456 1988 5516
rect 2073 5476 2077 5516
rect 2083 5476 2087 5516
rect 2225 5496 2229 5516
rect 2335 5476 2339 5516
rect 2355 5476 2359 5516
rect 2365 5476 2369 5516
rect 2451 5476 2455 5516
rect 2471 5476 2475 5516
rect 2491 5476 2495 5516
rect 2648 5456 2652 5516
rect 2656 5456 2660 5516
rect 2664 5456 2668 5516
rect 2788 5456 2792 5516
rect 2796 5456 2800 5516
rect 2804 5456 2808 5516
rect 2891 5476 2895 5516
rect 2911 5476 2915 5516
rect 2931 5476 2935 5516
rect 3031 5496 3035 5516
rect 3133 5476 3137 5516
rect 3143 5476 3147 5516
rect 3272 5456 3276 5516
rect 3280 5456 3284 5516
rect 3288 5456 3292 5516
rect 3413 5476 3417 5516
rect 3423 5476 3427 5516
rect 3531 5496 3535 5516
rect 3551 5496 3555 5516
rect 3571 5476 3575 5516
rect 3708 5456 3712 5516
rect 3716 5456 3720 5516
rect 3724 5456 3728 5516
rect 3832 5496 3836 5516
rect 3854 5476 3858 5516
rect 3862 5476 3866 5516
rect 3953 5476 3957 5516
rect 3963 5476 3967 5516
rect 4085 5476 4089 5516
rect 4105 5476 4109 5516
rect 4125 5476 4129 5516
rect 4233 5476 4237 5516
rect 4243 5476 4247 5516
rect 4368 5456 4372 5516
rect 4376 5456 4380 5516
rect 4384 5456 4388 5516
rect 4494 5476 4498 5516
rect 4502 5476 4506 5516
rect 4524 5496 4528 5516
rect 4631 5496 4635 5516
rect 4731 5476 4735 5516
rect 4751 5476 4755 5516
rect 4771 5476 4775 5516
rect 4831 5476 4835 5516
rect 4853 5496 4857 5516
rect 4863 5496 4867 5516
rect 4883 5496 4887 5516
rect 4891 5496 4895 5516
rect 4937 5496 4941 5516
rect 4959 5496 4963 5516
rect 4969 5496 4973 5516
rect 4991 5496 4995 5516
rect 5001 5496 5005 5516
rect 5021 5476 5025 5516
rect 5111 5496 5115 5516
rect 5171 5476 5175 5516
rect 5193 5496 5197 5516
rect 5203 5496 5207 5516
rect 5223 5496 5227 5516
rect 5231 5496 5235 5516
rect 5277 5496 5281 5516
rect 5299 5496 5303 5516
rect 5309 5496 5313 5516
rect 5331 5496 5335 5516
rect 5341 5496 5345 5516
rect 5361 5476 5365 5516
rect 5451 5476 5455 5516
rect 5471 5476 5475 5516
rect 5491 5476 5495 5516
rect 5613 5476 5617 5516
rect 5623 5476 5627 5516
rect 5733 5476 5737 5516
rect 5743 5476 5747 5516
rect 108 5064 112 5124
rect 116 5064 120 5124
rect 124 5064 128 5124
rect 214 5064 218 5104
rect 222 5064 226 5104
rect 244 5064 248 5084
rect 351 5064 355 5084
rect 488 5064 492 5124
rect 496 5064 500 5124
rect 504 5064 508 5124
rect 594 5064 598 5104
rect 602 5064 606 5104
rect 624 5064 628 5084
rect 752 5064 756 5084
rect 774 5064 778 5104
rect 782 5064 786 5104
rect 872 5064 876 5124
rect 880 5064 884 5124
rect 888 5064 892 5124
rect 1048 5064 1052 5124
rect 1056 5064 1060 5124
rect 1064 5064 1068 5124
rect 1151 5064 1155 5084
rect 1288 5064 1292 5124
rect 1296 5064 1300 5124
rect 1304 5064 1308 5124
rect 1425 5064 1429 5104
rect 1445 5064 1449 5104
rect 1465 5064 1469 5104
rect 1565 5064 1569 5084
rect 1665 5064 1669 5104
rect 1685 5064 1689 5104
rect 1705 5064 1709 5104
rect 1885 5064 1889 5084
rect 1905 5064 1909 5084
rect 1925 5064 1929 5084
rect 2066 5064 2070 5104
rect 2074 5064 2078 5104
rect 2094 5064 2098 5104
rect 2102 5064 2106 5104
rect 2193 5064 2197 5104
rect 2203 5064 2207 5104
rect 2348 5064 2352 5124
rect 2356 5064 2360 5124
rect 2364 5064 2368 5124
rect 2472 5064 2476 5084
rect 2494 5064 2498 5104
rect 2502 5064 2506 5104
rect 2605 5064 2609 5084
rect 2705 5064 2709 5104
rect 2725 5064 2729 5104
rect 2745 5064 2749 5104
rect 2865 5064 2869 5104
rect 2885 5064 2889 5104
rect 2905 5064 2909 5104
rect 3015 5064 3019 5104
rect 3035 5064 3039 5104
rect 3045 5064 3049 5104
rect 3131 5064 3135 5084
rect 3151 5064 3155 5084
rect 3285 5064 3289 5084
rect 3385 5064 3389 5084
rect 3405 5064 3409 5084
rect 3525 5064 3529 5104
rect 3545 5064 3549 5104
rect 3565 5064 3569 5104
rect 3653 5064 3657 5104
rect 3663 5064 3667 5104
rect 3793 5064 3797 5104
rect 3803 5064 3807 5104
rect 3933 5064 3937 5104
rect 3943 5064 3947 5104
rect 4032 5064 4036 5124
rect 4040 5064 4044 5124
rect 4048 5064 4052 5124
rect 4185 5064 4189 5104
rect 4205 5064 4209 5104
rect 4225 5064 4229 5104
rect 4331 5064 4335 5104
rect 4351 5064 4355 5104
rect 4371 5064 4375 5104
rect 4471 5064 4475 5084
rect 4608 5064 4612 5124
rect 4616 5064 4620 5124
rect 4624 5064 4628 5124
rect 4714 5064 4718 5104
rect 4722 5064 4726 5104
rect 4744 5064 4748 5084
rect 4851 5064 4855 5084
rect 4871 5064 4875 5084
rect 4931 5064 4935 5104
rect 4953 5064 4957 5084
rect 4963 5064 4967 5084
rect 4983 5064 4987 5084
rect 4991 5064 4995 5084
rect 5037 5064 5041 5084
rect 5059 5064 5063 5084
rect 5069 5064 5073 5084
rect 5091 5064 5095 5084
rect 5101 5064 5105 5084
rect 5121 5064 5125 5104
rect 5211 5064 5215 5104
rect 5231 5064 5235 5104
rect 5251 5064 5255 5104
rect 5351 5064 5355 5084
rect 5451 5064 5455 5104
rect 5471 5064 5475 5104
rect 5491 5064 5495 5104
rect 5613 5064 5617 5104
rect 5623 5064 5627 5104
rect 5713 5064 5717 5104
rect 5723 5064 5727 5104
rect 85 4996 89 5036
rect 105 4996 109 5036
rect 125 4996 129 5036
rect 248 4976 252 5036
rect 256 4976 260 5036
rect 264 4976 268 5036
rect 352 4976 356 5036
rect 360 4976 364 5036
rect 368 4976 372 5036
rect 491 4996 495 5036
rect 511 4996 515 5036
rect 531 4996 535 5036
rect 653 4996 657 5036
rect 663 4996 667 5036
rect 765 4996 769 5036
rect 785 4996 789 5036
rect 805 4996 809 5036
rect 905 4996 909 5036
rect 925 4996 929 5036
rect 945 4996 949 5036
rect 1052 5016 1056 5036
rect 1074 4996 1078 5036
rect 1082 4996 1086 5036
rect 1185 4996 1189 5036
rect 1205 4996 1209 5036
rect 1225 4996 1229 5036
rect 1325 5016 1329 5036
rect 1433 4996 1437 5036
rect 1443 4996 1447 5036
rect 1588 4976 1592 5036
rect 1596 4976 1600 5036
rect 1604 4976 1608 5036
rect 1705 4996 1709 5036
rect 1725 4996 1729 5036
rect 1745 4996 1749 5036
rect 1834 4996 1838 5036
rect 1842 4996 1846 5036
rect 1864 5016 1868 5036
rect 1973 4996 1977 5036
rect 1983 4996 1987 5036
rect 2112 5016 2116 5036
rect 2134 4996 2138 5036
rect 2142 4996 2146 5036
rect 2265 5016 2269 5036
rect 2365 4996 2369 5036
rect 2385 4996 2389 5036
rect 2405 4996 2409 5036
rect 2528 4976 2532 5036
rect 2536 4976 2540 5036
rect 2544 4976 2548 5036
rect 2645 5016 2649 5036
rect 2773 4996 2777 5036
rect 2783 4996 2787 5036
rect 2871 5016 2875 5036
rect 2972 4976 2976 5036
rect 2980 4976 2984 5036
rect 2988 4976 2992 5036
rect 3125 4996 3129 5036
rect 3145 4996 3149 5036
rect 3165 4996 3169 5036
rect 3265 4996 3269 5036
rect 3285 4996 3289 5036
rect 3305 4996 3309 5036
rect 3412 5016 3416 5036
rect 3434 4996 3438 5036
rect 3442 4996 3446 5036
rect 3531 5016 3535 5036
rect 3551 5016 3555 5036
rect 3571 4996 3575 5036
rect 3685 5016 3689 5036
rect 3705 5016 3709 5036
rect 3828 4976 3832 5036
rect 3836 4976 3840 5036
rect 3844 4976 3848 5036
rect 3945 5016 3949 5036
rect 4032 4976 4036 5036
rect 4040 4976 4044 5036
rect 4048 4976 4052 5036
rect 4172 4976 4176 5036
rect 4180 4976 4184 5036
rect 4188 4976 4192 5036
rect 4335 4996 4339 5036
rect 4355 4996 4359 5036
rect 4365 4996 4369 5036
rect 4471 5016 4475 5036
rect 4491 5016 4495 5036
rect 4511 4996 4515 5036
rect 4611 5016 4615 5036
rect 4631 5016 4635 5036
rect 4745 4996 4749 5036
rect 4765 4996 4769 5036
rect 4785 4996 4789 5036
rect 4831 4996 4835 5036
rect 4853 5016 4857 5036
rect 4863 5016 4867 5036
rect 4883 5016 4887 5036
rect 4891 5016 4895 5036
rect 4937 5016 4941 5036
rect 4959 5016 4963 5036
rect 4969 5016 4973 5036
rect 4991 5016 4995 5036
rect 5001 5016 5005 5036
rect 5021 4996 5025 5036
rect 5111 4996 5115 5036
rect 5131 4996 5135 5036
rect 5151 4996 5155 5036
rect 5211 4996 5215 5036
rect 5233 5016 5237 5036
rect 5243 5016 5247 5036
rect 5263 5016 5267 5036
rect 5271 5016 5275 5036
rect 5317 5016 5321 5036
rect 5339 5016 5343 5036
rect 5349 5016 5353 5036
rect 5371 5016 5375 5036
rect 5381 5016 5385 5036
rect 5401 4996 5405 5036
rect 5513 4996 5517 5036
rect 5523 4996 5527 5036
rect 5613 4996 5617 5036
rect 5623 4996 5627 5036
rect 5753 4996 5757 5036
rect 5763 4996 5767 5036
rect 92 4584 96 4604
rect 114 4584 118 4624
rect 122 4584 126 4624
rect 248 4584 252 4644
rect 256 4584 260 4644
rect 264 4584 268 4644
rect 354 4584 358 4624
rect 362 4584 366 4624
rect 384 4584 388 4604
rect 493 4584 497 4624
rect 503 4584 507 4624
rect 648 4584 652 4644
rect 656 4584 660 4644
rect 664 4584 668 4644
rect 808 4584 812 4644
rect 816 4584 820 4644
rect 824 4584 828 4644
rect 911 4584 915 4604
rect 1011 4584 1015 4604
rect 1125 4584 1129 4604
rect 1225 4584 1229 4624
rect 1245 4584 1249 4624
rect 1265 4584 1269 4624
rect 1351 4584 1355 4624
rect 1371 4584 1375 4624
rect 1391 4584 1395 4624
rect 1491 4584 1495 4604
rect 1592 4584 1596 4644
rect 1600 4584 1604 4644
rect 1608 4584 1612 4644
rect 1745 4584 1749 4624
rect 1765 4584 1769 4624
rect 1785 4584 1789 4624
rect 1893 4584 1897 4624
rect 1903 4584 1907 4624
rect 1991 4584 1995 4624
rect 2011 4584 2015 4624
rect 2031 4584 2035 4624
rect 2168 4584 2172 4644
rect 2176 4584 2180 4644
rect 2184 4584 2188 4644
rect 2283 4584 2287 4624
rect 2305 4584 2309 4604
rect 2393 4584 2397 4624
rect 2403 4584 2407 4624
rect 2513 4584 2517 4624
rect 2523 4584 2527 4624
rect 2643 4584 2647 4624
rect 2665 4584 2669 4604
rect 2752 4584 2756 4644
rect 2760 4584 2764 4644
rect 2768 4584 2772 4644
rect 2905 4584 2909 4604
rect 2925 4584 2929 4604
rect 3031 4584 3035 4624
rect 3051 4584 3055 4624
rect 3071 4584 3075 4624
rect 3091 4584 3095 4624
rect 3213 4584 3217 4624
rect 3223 4584 3227 4624
rect 3348 4584 3352 4644
rect 3356 4584 3360 4644
rect 3364 4584 3368 4644
rect 3472 4584 3476 4604
rect 3494 4584 3498 4624
rect 3502 4584 3506 4624
rect 3628 4584 3632 4644
rect 3636 4584 3640 4644
rect 3644 4584 3648 4644
rect 3752 4584 3756 4604
rect 3774 4584 3778 4624
rect 3782 4584 3786 4624
rect 3872 4584 3876 4644
rect 3880 4584 3884 4644
rect 3888 4584 3892 4644
rect 4012 4584 4016 4644
rect 4020 4584 4024 4644
rect 4028 4584 4032 4644
rect 4151 4584 4155 4604
rect 4275 4584 4279 4624
rect 4295 4584 4299 4624
rect 4305 4584 4309 4624
rect 4448 4584 4452 4644
rect 4456 4584 4460 4644
rect 4464 4584 4468 4644
rect 4552 4584 4556 4644
rect 4560 4584 4564 4644
rect 4568 4584 4572 4644
rect 4691 4584 4695 4604
rect 4751 4584 4755 4624
rect 4773 4584 4777 4604
rect 4783 4584 4787 4604
rect 4803 4584 4807 4604
rect 4811 4584 4815 4604
rect 4857 4584 4861 4604
rect 4879 4584 4883 4604
rect 4889 4584 4893 4604
rect 4911 4584 4915 4604
rect 4921 4584 4925 4604
rect 4941 4584 4945 4624
rect 5031 4584 5035 4624
rect 5051 4584 5055 4624
rect 5071 4584 5075 4624
rect 5173 4584 5177 4624
rect 5183 4584 5187 4624
rect 5293 4584 5297 4624
rect 5303 4584 5307 4624
rect 5433 4584 5437 4624
rect 5443 4584 5447 4624
rect 5553 4584 5557 4624
rect 5563 4584 5567 4624
rect 5708 4584 5712 4644
rect 5716 4584 5720 4644
rect 5724 4584 5728 4644
rect 85 4516 89 4556
rect 105 4516 109 4556
rect 125 4516 129 4556
rect 248 4496 252 4556
rect 256 4496 260 4556
rect 264 4496 268 4556
rect 354 4516 358 4556
rect 362 4516 366 4556
rect 384 4536 388 4556
rect 525 4516 529 4556
rect 545 4516 549 4556
rect 565 4516 569 4556
rect 665 4516 669 4556
rect 685 4516 689 4556
rect 705 4516 709 4556
rect 791 4536 795 4556
rect 894 4516 898 4556
rect 902 4516 906 4556
rect 924 4536 928 4556
rect 1045 4536 1049 4556
rect 1168 4496 1172 4556
rect 1176 4496 1180 4556
rect 1184 4496 1188 4556
rect 1292 4536 1296 4556
rect 1314 4516 1318 4556
rect 1322 4516 1326 4556
rect 1425 4536 1429 4556
rect 1511 4516 1515 4556
rect 1531 4516 1535 4556
rect 1551 4516 1555 4556
rect 1673 4516 1677 4556
rect 1683 4516 1687 4556
rect 1808 4496 1812 4556
rect 1816 4496 1820 4556
rect 1824 4496 1828 4556
rect 1925 4536 1929 4556
rect 1945 4536 1949 4556
rect 2068 4496 2072 4556
rect 2076 4496 2080 4556
rect 2084 4496 2088 4556
rect 2228 4496 2232 4556
rect 2236 4496 2240 4556
rect 2244 4496 2248 4556
rect 2353 4516 2357 4556
rect 2363 4516 2367 4556
rect 2488 4496 2492 4556
rect 2496 4496 2500 4556
rect 2504 4496 2508 4556
rect 2592 4496 2596 4556
rect 2600 4496 2604 4556
rect 2608 4496 2612 4556
rect 2745 4536 2749 4556
rect 2845 4536 2849 4556
rect 2865 4536 2869 4556
rect 2988 4496 2992 4556
rect 2996 4496 3000 4556
rect 3004 4496 3008 4556
rect 3128 4496 3132 4556
rect 3136 4496 3140 4556
rect 3144 4496 3148 4556
rect 3231 4536 3235 4556
rect 3331 4516 3335 4556
rect 3351 4516 3355 4556
rect 3371 4516 3375 4556
rect 3495 4516 3499 4556
rect 3515 4516 3519 4556
rect 3525 4516 3529 4556
rect 3633 4516 3637 4556
rect 3643 4516 3647 4556
rect 3765 4516 3769 4556
rect 3785 4536 3789 4556
rect 3805 4536 3809 4556
rect 3893 4516 3897 4556
rect 3903 4516 3907 4556
rect 4023 4516 4027 4556
rect 4045 4536 4049 4556
rect 4131 4516 4135 4556
rect 4141 4516 4145 4556
rect 4161 4516 4165 4556
rect 4293 4516 4297 4556
rect 4303 4516 4307 4556
rect 4405 4516 4409 4556
rect 4425 4516 4429 4556
rect 4445 4516 4449 4556
rect 4533 4516 4537 4556
rect 4543 4516 4547 4556
rect 4673 4516 4677 4556
rect 4683 4516 4687 4556
rect 4771 4536 4775 4556
rect 4873 4516 4877 4556
rect 4883 4516 4887 4556
rect 4991 4516 4995 4556
rect 5011 4516 5015 4556
rect 5031 4516 5035 4556
rect 5091 4516 5095 4556
rect 5113 4536 5117 4556
rect 5123 4536 5127 4556
rect 5143 4536 5147 4556
rect 5151 4536 5155 4556
rect 5197 4536 5201 4556
rect 5219 4536 5223 4556
rect 5229 4536 5233 4556
rect 5251 4536 5255 4556
rect 5261 4536 5265 4556
rect 5281 4516 5285 4556
rect 5371 4516 5375 4556
rect 5391 4516 5395 4556
rect 5411 4516 5415 4556
rect 5511 4536 5515 4556
rect 5531 4536 5535 4556
rect 5551 4516 5555 4556
rect 5665 4516 5669 4556
rect 5685 4516 5689 4556
rect 5705 4516 5709 4556
rect 105 4104 109 4144
rect 125 4104 129 4144
rect 145 4104 149 4144
rect 245 4104 249 4144
rect 265 4104 269 4144
rect 285 4104 289 4144
rect 428 4104 432 4164
rect 436 4104 440 4164
rect 444 4104 448 4164
rect 568 4104 572 4164
rect 576 4104 580 4164
rect 584 4104 588 4164
rect 685 4104 689 4144
rect 705 4104 709 4124
rect 725 4104 729 4124
rect 825 4104 829 4144
rect 845 4104 849 4144
rect 865 4104 869 4144
rect 951 4104 955 4124
rect 1072 4104 1076 4124
rect 1094 4104 1098 4144
rect 1102 4104 1106 4144
rect 1248 4104 1252 4164
rect 1256 4104 1260 4164
rect 1264 4104 1268 4164
rect 1373 4104 1377 4144
rect 1383 4104 1387 4144
rect 1493 4104 1497 4144
rect 1503 4104 1507 4144
rect 1605 4104 1609 4124
rect 1625 4104 1629 4124
rect 1748 4104 1752 4164
rect 1756 4104 1760 4164
rect 1764 4104 1768 4164
rect 1888 4104 1892 4164
rect 1896 4104 1900 4164
rect 1904 4104 1908 4164
rect 1992 4104 1996 4164
rect 2000 4104 2004 4164
rect 2008 4104 2012 4164
rect 2132 4104 2136 4164
rect 2140 4104 2144 4164
rect 2148 4104 2152 4164
rect 2285 4104 2289 4124
rect 2305 4104 2309 4124
rect 2425 4104 2429 4144
rect 2445 4104 2449 4144
rect 2465 4104 2469 4144
rect 2608 4104 2612 4164
rect 2616 4104 2620 4164
rect 2624 4104 2628 4164
rect 2711 4104 2715 4124
rect 2832 4104 2836 4164
rect 2840 4104 2844 4164
rect 2848 4104 2852 4164
rect 2973 4104 2977 4144
rect 2983 4104 2987 4144
rect 3094 4104 3098 4144
rect 3102 4104 3106 4144
rect 3124 4104 3128 4124
rect 3234 4104 3238 4144
rect 3242 4104 3246 4144
rect 3264 4104 3268 4124
rect 3371 4104 3375 4144
rect 3391 4104 3395 4144
rect 3411 4104 3415 4144
rect 3531 4104 3535 4124
rect 3632 4104 3636 4164
rect 3640 4104 3644 4164
rect 3648 4104 3652 4164
rect 3772 4104 3776 4164
rect 3780 4104 3784 4164
rect 3788 4104 3792 4164
rect 3933 4104 3937 4144
rect 3943 4104 3947 4144
rect 4073 4104 4077 4144
rect 4083 4104 4087 4144
rect 4193 4104 4197 4144
rect 4203 4104 4207 4144
rect 4305 4104 4309 4144
rect 4325 4104 4329 4144
rect 4345 4104 4349 4144
rect 4431 4104 4435 4124
rect 4451 4104 4455 4124
rect 4471 4104 4475 4144
rect 4585 4104 4589 4144
rect 4605 4104 4609 4144
rect 4625 4104 4629 4144
rect 4731 4104 4735 4144
rect 4751 4104 4755 4144
rect 4771 4104 4775 4144
rect 4871 4104 4875 4124
rect 4891 4104 4895 4124
rect 4991 4104 4995 4124
rect 5114 4104 5118 4144
rect 5122 4104 5126 4144
rect 5144 4104 5148 4124
rect 5251 4104 5255 4144
rect 5271 4104 5275 4144
rect 5291 4104 5295 4144
rect 5391 4104 5395 4124
rect 5491 4104 5495 4144
rect 5511 4104 5515 4144
rect 5531 4104 5535 4144
rect 5595 4104 5599 4144
rect 5615 4104 5619 4124
rect 5625 4104 5629 4124
rect 5647 4104 5651 4124
rect 5657 4104 5661 4124
rect 5679 4104 5683 4124
rect 5725 4104 5729 4124
rect 5733 4104 5737 4124
rect 5753 4104 5757 4124
rect 5763 4104 5767 4124
rect 5785 4104 5789 4144
rect 85 4056 89 4076
rect 191 4036 195 4076
rect 211 4036 215 4076
rect 231 4036 235 4076
rect 345 4056 349 4076
rect 454 4036 458 4076
rect 462 4036 466 4076
rect 484 4056 488 4076
rect 605 4056 609 4076
rect 625 4056 629 4076
rect 745 4056 749 4076
rect 831 4036 835 4076
rect 851 4036 855 4076
rect 871 4036 875 4076
rect 971 4056 975 4076
rect 1072 4016 1076 4076
rect 1080 4016 1084 4076
rect 1088 4016 1092 4076
rect 1214 4036 1218 4076
rect 1222 4036 1226 4076
rect 1242 4036 1246 4076
rect 1250 4036 1254 4076
rect 1393 4036 1397 4076
rect 1403 4036 1407 4076
rect 1525 4056 1529 4076
rect 1625 4056 1629 4076
rect 1645 4056 1649 4076
rect 1745 4056 1749 4076
rect 1832 4016 1836 4076
rect 1840 4016 1844 4076
rect 1848 4016 1852 4076
rect 1985 4036 1989 4076
rect 2005 4036 2009 4076
rect 2025 4036 2029 4076
rect 2168 4016 2172 4076
rect 2176 4016 2180 4076
rect 2184 4016 2188 4076
rect 2272 4016 2276 4076
rect 2280 4016 2284 4076
rect 2288 4016 2292 4076
rect 2425 4036 2429 4076
rect 2445 4036 2449 4076
rect 2465 4036 2469 4076
rect 2573 4036 2577 4076
rect 2583 4036 2587 4076
rect 2673 4036 2677 4076
rect 2683 4036 2687 4076
rect 2792 4016 2796 4076
rect 2800 4016 2804 4076
rect 2808 4016 2812 4076
rect 2932 4016 2936 4076
rect 2940 4016 2944 4076
rect 2948 4016 2952 4076
rect 3085 4056 3089 4076
rect 3208 4016 3212 4076
rect 3216 4016 3220 4076
rect 3224 4016 3228 4076
rect 3325 4056 3329 4076
rect 3425 4036 3429 4076
rect 3445 4036 3449 4076
rect 3465 4036 3469 4076
rect 3553 4036 3557 4076
rect 3563 4036 3567 4076
rect 3685 4036 3689 4076
rect 3705 4056 3709 4076
rect 3725 4056 3729 4076
rect 3833 4036 3837 4076
rect 3843 4036 3847 4076
rect 3965 4036 3969 4076
rect 3985 4036 3989 4076
rect 4005 4036 4009 4076
rect 4112 4056 4116 4076
rect 4134 4036 4138 4076
rect 4142 4036 4146 4076
rect 4233 4036 4237 4076
rect 4243 4036 4247 4076
rect 4351 4036 4355 4076
rect 4371 4036 4375 4076
rect 4391 4036 4395 4076
rect 4491 4036 4495 4076
rect 4511 4036 4515 4076
rect 4531 4036 4535 4076
rect 4631 4056 4635 4076
rect 4651 4056 4655 4076
rect 4671 4036 4675 4076
rect 4793 4036 4797 4076
rect 4803 4036 4807 4076
rect 4892 4016 4896 4076
rect 4900 4016 4904 4076
rect 4908 4016 4912 4076
rect 5031 4056 5035 4076
rect 5145 4056 5149 4076
rect 5191 4036 5195 4076
rect 5213 4056 5217 4076
rect 5223 4056 5227 4076
rect 5243 4056 5247 4076
rect 5251 4056 5255 4076
rect 5297 4056 5301 4076
rect 5319 4056 5323 4076
rect 5329 4056 5333 4076
rect 5351 4056 5355 4076
rect 5361 4056 5365 4076
rect 5381 4036 5385 4076
rect 5431 4036 5435 4076
rect 5453 4056 5457 4076
rect 5463 4056 5467 4076
rect 5483 4056 5487 4076
rect 5491 4056 5495 4076
rect 5537 4056 5541 4076
rect 5559 4056 5563 4076
rect 5569 4056 5573 4076
rect 5591 4056 5595 4076
rect 5601 4056 5605 4076
rect 5621 4036 5625 4076
rect 5711 4036 5715 4076
rect 5731 4036 5735 4076
rect 5751 4036 5755 4076
rect 93 3624 97 3664
rect 103 3624 107 3664
rect 228 3624 232 3684
rect 236 3624 240 3684
rect 244 3624 248 3684
rect 405 3624 409 3644
rect 425 3624 429 3644
rect 445 3624 449 3644
rect 565 3624 569 3664
rect 585 3624 589 3664
rect 605 3624 609 3664
rect 713 3624 717 3664
rect 723 3624 727 3664
rect 811 3624 815 3664
rect 831 3624 835 3664
rect 851 3624 855 3664
rect 1006 3624 1010 3664
rect 1014 3624 1018 3664
rect 1034 3624 1038 3664
rect 1042 3624 1046 3664
rect 1133 3624 1137 3664
rect 1143 3624 1147 3664
rect 1252 3624 1256 3684
rect 1260 3624 1264 3684
rect 1268 3624 1272 3684
rect 1394 3624 1398 3664
rect 1402 3624 1406 3664
rect 1424 3624 1428 3644
rect 1531 3624 1535 3664
rect 1551 3624 1555 3664
rect 1571 3624 1575 3664
rect 1671 3624 1675 3644
rect 1793 3624 1797 3664
rect 1803 3624 1807 3664
rect 1893 3624 1897 3664
rect 1903 3624 1907 3664
rect 2011 3624 2015 3644
rect 2031 3624 2035 3644
rect 2051 3624 2055 3664
rect 2153 3624 2157 3664
rect 2163 3624 2167 3664
rect 2272 3624 2276 3684
rect 2280 3624 2284 3684
rect 2288 3624 2292 3684
rect 2425 3624 2429 3664
rect 2445 3624 2449 3664
rect 2465 3624 2469 3664
rect 2553 3624 2557 3664
rect 2563 3624 2567 3664
rect 2671 3624 2675 3664
rect 2691 3624 2695 3664
rect 2711 3624 2715 3664
rect 2825 3624 2829 3644
rect 2925 3624 2929 3664
rect 2945 3624 2949 3664
rect 2965 3624 2969 3664
rect 3053 3624 3057 3664
rect 3063 3624 3067 3664
rect 3213 3624 3217 3664
rect 3223 3624 3227 3664
rect 3325 3624 3329 3644
rect 3412 3624 3416 3684
rect 3420 3624 3424 3684
rect 3428 3624 3432 3684
rect 3551 3624 3555 3644
rect 3665 3624 3669 3644
rect 3685 3624 3689 3644
rect 3793 3624 3797 3664
rect 3803 3624 3807 3664
rect 3911 3624 3915 3644
rect 4025 3624 4029 3644
rect 4071 3624 4075 3664
rect 4093 3624 4097 3644
rect 4103 3624 4107 3644
rect 4123 3624 4127 3644
rect 4131 3624 4135 3644
rect 4177 3624 4181 3644
rect 4199 3624 4203 3644
rect 4209 3624 4213 3644
rect 4231 3624 4235 3644
rect 4241 3624 4245 3644
rect 4261 3624 4265 3664
rect 4365 3624 4369 3664
rect 4385 3624 4389 3664
rect 4405 3624 4409 3664
rect 4425 3624 4429 3664
rect 4513 3624 4517 3664
rect 4523 3624 4527 3664
rect 4631 3624 4635 3644
rect 4651 3624 4655 3644
rect 4751 3624 4755 3664
rect 4771 3624 4775 3664
rect 4791 3624 4795 3664
rect 4891 3624 4895 3664
rect 5033 3624 5037 3664
rect 5043 3624 5047 3664
rect 5131 3624 5135 3644
rect 5245 3624 5249 3664
rect 5265 3624 5269 3664
rect 5285 3624 5289 3664
rect 5305 3624 5309 3664
rect 5325 3624 5329 3664
rect 5345 3624 5349 3664
rect 5365 3624 5369 3664
rect 5385 3624 5389 3664
rect 5431 3624 5435 3664
rect 5453 3624 5457 3644
rect 5463 3624 5467 3644
rect 5483 3624 5487 3644
rect 5491 3624 5495 3644
rect 5537 3624 5541 3644
rect 5559 3624 5563 3644
rect 5569 3624 5573 3644
rect 5591 3624 5595 3644
rect 5601 3624 5605 3644
rect 5621 3624 5625 3664
rect 5733 3624 5737 3664
rect 5743 3624 5747 3664
rect 85 3556 89 3596
rect 105 3556 109 3596
rect 125 3556 129 3596
rect 214 3556 218 3596
rect 222 3556 226 3596
rect 244 3576 248 3596
rect 351 3576 355 3596
rect 451 3556 455 3596
rect 471 3556 475 3596
rect 491 3556 495 3596
rect 592 3536 596 3596
rect 600 3536 604 3596
rect 608 3536 612 3596
rect 773 3556 777 3596
rect 783 3556 787 3596
rect 893 3556 897 3596
rect 903 3556 907 3596
rect 991 3556 995 3596
rect 1011 3556 1015 3596
rect 1031 3556 1035 3596
rect 1168 3536 1172 3596
rect 1176 3536 1180 3596
rect 1184 3536 1188 3596
rect 1273 3556 1277 3596
rect 1283 3556 1287 3596
rect 1428 3536 1432 3596
rect 1436 3536 1440 3596
rect 1444 3536 1448 3596
rect 1531 3556 1535 3596
rect 1551 3556 1555 3596
rect 1571 3556 1575 3596
rect 1692 3576 1696 3596
rect 1714 3556 1718 3596
rect 1722 3556 1726 3596
rect 1848 3536 1852 3596
rect 1856 3536 1860 3596
rect 1864 3536 1868 3596
rect 1954 3556 1958 3596
rect 1962 3556 1966 3596
rect 1984 3576 1988 3596
rect 2105 3556 2109 3596
rect 2125 3556 2129 3596
rect 2145 3556 2149 3596
rect 2251 3556 2255 3596
rect 2271 3556 2275 3596
rect 2291 3556 2295 3596
rect 2412 3576 2416 3596
rect 2434 3556 2438 3596
rect 2442 3556 2446 3596
rect 2555 3556 2559 3596
rect 2575 3556 2579 3596
rect 2585 3556 2589 3596
rect 2673 3556 2677 3596
rect 2683 3556 2687 3596
rect 2805 3556 2809 3596
rect 2825 3556 2829 3596
rect 2845 3556 2849 3596
rect 2963 3556 2967 3596
rect 2985 3576 2989 3596
rect 3093 3556 3097 3596
rect 3103 3556 3107 3596
rect 3192 3536 3196 3596
rect 3200 3536 3204 3596
rect 3208 3536 3212 3596
rect 3368 3536 3372 3596
rect 3376 3536 3380 3596
rect 3384 3536 3388 3596
rect 3485 3556 3489 3596
rect 3505 3556 3509 3596
rect 3525 3556 3529 3596
rect 3625 3556 3629 3596
rect 3645 3556 3649 3596
rect 3665 3556 3669 3596
rect 3775 3556 3779 3596
rect 3795 3556 3799 3596
rect 3805 3556 3809 3596
rect 3891 3576 3895 3596
rect 3911 3576 3915 3596
rect 4045 3556 4049 3596
rect 4065 3556 4069 3596
rect 4085 3556 4089 3596
rect 4171 3576 4175 3596
rect 4271 3556 4275 3596
rect 4291 3556 4295 3596
rect 4311 3556 4315 3596
rect 4433 3556 4437 3596
rect 4443 3556 4447 3596
rect 4533 3556 4537 3596
rect 4543 3556 4547 3596
rect 4611 3556 4615 3596
rect 4633 3576 4637 3596
rect 4643 3576 4647 3596
rect 4663 3576 4667 3596
rect 4671 3576 4675 3596
rect 4717 3576 4721 3596
rect 4739 3576 4743 3596
rect 4749 3576 4753 3596
rect 4771 3576 4775 3596
rect 4781 3576 4785 3596
rect 4801 3556 4805 3596
rect 4913 3556 4917 3596
rect 4923 3556 4927 3596
rect 5025 3556 5029 3596
rect 5045 3556 5049 3596
rect 5065 3556 5069 3596
rect 5173 3556 5177 3596
rect 5183 3556 5187 3596
rect 5255 3556 5259 3596
rect 5275 3576 5279 3596
rect 5285 3576 5289 3596
rect 5307 3576 5311 3596
rect 5317 3576 5321 3596
rect 5339 3576 5343 3596
rect 5385 3576 5389 3596
rect 5393 3576 5397 3596
rect 5413 3576 5417 3596
rect 5423 3576 5427 3596
rect 5445 3556 5449 3596
rect 5553 3556 5557 3596
rect 5563 3556 5567 3596
rect 5651 3556 5655 3596
rect 5671 3556 5675 3596
rect 5691 3556 5695 3596
rect 85 3144 89 3164
rect 185 3144 189 3184
rect 205 3144 209 3184
rect 225 3144 229 3184
rect 325 3144 329 3164
rect 413 3144 417 3184
rect 423 3144 427 3184
rect 534 3144 538 3184
rect 542 3144 546 3184
rect 564 3144 568 3164
rect 671 3144 675 3184
rect 681 3144 685 3184
rect 701 3144 705 3184
rect 853 3144 857 3184
rect 863 3144 867 3184
rect 988 3144 992 3204
rect 996 3144 1000 3204
rect 1004 3144 1008 3204
rect 1128 3144 1132 3204
rect 1136 3144 1140 3204
rect 1144 3144 1148 3204
rect 1234 3144 1238 3184
rect 1242 3144 1246 3184
rect 1264 3144 1268 3164
rect 1385 3144 1389 3164
rect 1508 3144 1512 3204
rect 1516 3144 1520 3204
rect 1524 3144 1528 3204
rect 1648 3144 1652 3204
rect 1656 3144 1660 3204
rect 1664 3144 1668 3204
rect 1772 3144 1776 3164
rect 1794 3144 1798 3184
rect 1802 3144 1806 3184
rect 1933 3144 1937 3184
rect 1943 3144 1947 3184
rect 2052 3144 2056 3164
rect 2074 3144 2078 3184
rect 2082 3144 2086 3184
rect 2173 3144 2177 3184
rect 2183 3144 2187 3184
rect 2315 3144 2319 3184
rect 2335 3144 2339 3184
rect 2345 3144 2349 3184
rect 2433 3144 2437 3184
rect 2443 3144 2447 3184
rect 2565 3144 2569 3184
rect 2585 3144 2589 3184
rect 2605 3144 2609 3184
rect 2712 3144 2716 3164
rect 2734 3144 2738 3184
rect 2742 3144 2746 3184
rect 2832 3144 2836 3204
rect 2840 3144 2844 3204
rect 2848 3144 2852 3204
rect 2972 3144 2976 3204
rect 2980 3144 2984 3204
rect 2988 3144 2992 3204
rect 3133 3144 3137 3184
rect 3143 3144 3147 3184
rect 3273 3144 3277 3184
rect 3283 3144 3287 3184
rect 3371 3144 3375 3164
rect 3508 3144 3512 3204
rect 3516 3144 3520 3204
rect 3524 3144 3528 3204
rect 3614 3144 3618 3184
rect 3622 3144 3626 3184
rect 3644 3144 3648 3164
rect 3765 3144 3769 3184
rect 3785 3144 3789 3184
rect 3805 3144 3809 3184
rect 3891 3144 3895 3164
rect 3951 3144 3955 3184
rect 3973 3144 3977 3164
rect 3983 3144 3987 3164
rect 4003 3144 4007 3164
rect 4011 3144 4015 3164
rect 4057 3144 4061 3164
rect 4079 3144 4083 3164
rect 4089 3144 4093 3164
rect 4111 3144 4115 3164
rect 4121 3144 4125 3164
rect 4141 3144 4145 3184
rect 4231 3144 4235 3184
rect 4251 3144 4255 3184
rect 4271 3144 4275 3184
rect 4371 3144 4375 3184
rect 4391 3144 4395 3184
rect 4411 3144 4415 3184
rect 4471 3144 4475 3184
rect 4493 3144 4497 3164
rect 4503 3144 4507 3164
rect 4523 3144 4527 3164
rect 4531 3144 4535 3164
rect 4577 3144 4581 3164
rect 4599 3144 4603 3164
rect 4609 3144 4613 3164
rect 4631 3144 4635 3164
rect 4641 3144 4645 3164
rect 4661 3144 4665 3184
rect 4751 3144 4755 3184
rect 4771 3144 4775 3184
rect 4791 3144 4795 3184
rect 4913 3144 4917 3184
rect 4923 3144 4927 3184
rect 5025 3144 5029 3184
rect 5045 3144 5049 3184
rect 5065 3144 5069 3184
rect 5165 3144 5169 3164
rect 5273 3144 5277 3184
rect 5283 3144 5287 3184
rect 5371 3144 5375 3164
rect 5491 3144 5495 3184
rect 5511 3144 5515 3184
rect 5531 3144 5535 3184
rect 5673 3144 5677 3184
rect 5683 3144 5687 3184
rect 115 3076 119 3116
rect 135 3076 139 3116
rect 145 3076 149 3116
rect 252 3056 256 3116
rect 260 3056 264 3116
rect 268 3056 272 3116
rect 393 3076 397 3116
rect 403 3076 407 3116
rect 525 3076 529 3116
rect 545 3076 549 3116
rect 565 3076 569 3116
rect 651 3076 655 3116
rect 671 3076 675 3116
rect 691 3076 695 3116
rect 791 3076 795 3116
rect 811 3076 815 3116
rect 831 3076 835 3116
rect 931 3076 935 3116
rect 951 3076 955 3116
rect 971 3076 975 3116
rect 1093 3076 1097 3116
rect 1103 3076 1107 3116
rect 1225 3096 1229 3116
rect 1245 3096 1249 3116
rect 1331 3076 1335 3116
rect 1351 3076 1355 3116
rect 1371 3076 1375 3116
rect 1508 3056 1512 3116
rect 1516 3056 1520 3116
rect 1524 3056 1528 3116
rect 1652 3096 1656 3116
rect 1674 3076 1678 3116
rect 1682 3076 1686 3116
rect 1785 3076 1789 3116
rect 1805 3076 1809 3116
rect 1825 3076 1829 3116
rect 1911 3076 1915 3116
rect 1931 3076 1935 3116
rect 1951 3076 1955 3116
rect 2085 3076 2089 3116
rect 2105 3076 2109 3116
rect 2125 3076 2129 3116
rect 2225 3076 2229 3116
rect 2245 3076 2249 3116
rect 2265 3076 2269 3116
rect 2392 3096 2396 3116
rect 2414 3076 2418 3116
rect 2422 3076 2426 3116
rect 2532 3096 2536 3116
rect 2554 3076 2558 3116
rect 2562 3076 2566 3116
rect 2686 3076 2690 3116
rect 2694 3076 2698 3116
rect 2714 3076 2718 3116
rect 2722 3076 2726 3116
rect 2825 3076 2829 3116
rect 2845 3096 2849 3116
rect 2865 3096 2869 3116
rect 2951 3096 2955 3116
rect 2971 3096 2975 3116
rect 3093 3076 3097 3116
rect 3103 3076 3107 3116
rect 3235 3076 3239 3116
rect 3255 3076 3259 3116
rect 3265 3076 3269 3116
rect 3351 3096 3355 3116
rect 3371 3096 3375 3116
rect 3391 3076 3395 3116
rect 3505 3076 3509 3116
rect 3525 3076 3529 3116
rect 3545 3076 3549 3116
rect 3645 3076 3649 3116
rect 3665 3076 3669 3116
rect 3685 3076 3689 3116
rect 3785 3076 3789 3116
rect 3805 3096 3809 3116
rect 3825 3096 3829 3116
rect 3955 3076 3959 3116
rect 3975 3076 3979 3116
rect 3985 3076 3989 3116
rect 4071 3096 4075 3116
rect 4091 3096 4095 3116
rect 4192 3056 4196 3116
rect 4200 3056 4204 3116
rect 4208 3056 4212 3116
rect 4295 3076 4299 3116
rect 4315 3096 4319 3116
rect 4325 3096 4329 3116
rect 4347 3096 4351 3116
rect 4357 3096 4361 3116
rect 4379 3096 4383 3116
rect 4425 3096 4429 3116
rect 4433 3096 4437 3116
rect 4453 3096 4457 3116
rect 4463 3096 4467 3116
rect 4485 3076 4489 3116
rect 4591 3076 4595 3116
rect 4611 3076 4615 3116
rect 4631 3076 4635 3116
rect 4731 3076 4735 3116
rect 4751 3076 4755 3116
rect 4771 3076 4775 3116
rect 4893 3076 4897 3116
rect 4903 3076 4907 3116
rect 4993 3076 4997 3116
rect 5003 3076 5007 3116
rect 5075 3076 5079 3116
rect 5095 3096 5099 3116
rect 5105 3096 5109 3116
rect 5127 3096 5131 3116
rect 5137 3096 5141 3116
rect 5159 3096 5163 3116
rect 5205 3096 5209 3116
rect 5213 3096 5217 3116
rect 5233 3096 5237 3116
rect 5243 3096 5247 3116
rect 5265 3076 5269 3116
rect 5365 3076 5369 3116
rect 5385 3076 5389 3116
rect 5405 3076 5409 3116
rect 5425 3076 5429 3116
rect 5445 3076 5449 3116
rect 5465 3076 5469 3116
rect 5485 3076 5489 3116
rect 5505 3076 5509 3116
rect 5551 3076 5555 3116
rect 5573 3096 5577 3116
rect 5583 3096 5587 3116
rect 5603 3096 5607 3116
rect 5611 3096 5615 3116
rect 5657 3096 5661 3116
rect 5679 3096 5683 3116
rect 5689 3096 5693 3116
rect 5711 3096 5715 3116
rect 5721 3096 5725 3116
rect 5741 3076 5745 3116
rect 93 2664 97 2704
rect 103 2664 107 2704
rect 191 2664 195 2704
rect 211 2664 215 2704
rect 231 2664 235 2704
rect 345 2664 349 2684
rect 434 2664 438 2704
rect 442 2664 446 2704
rect 464 2664 468 2684
rect 593 2664 597 2704
rect 603 2664 607 2704
rect 691 2664 695 2704
rect 701 2664 705 2704
rect 721 2664 725 2704
rect 833 2664 837 2704
rect 843 2664 847 2704
rect 954 2664 958 2704
rect 962 2664 966 2704
rect 984 2664 988 2684
rect 1093 2664 1097 2704
rect 1103 2664 1107 2704
rect 1245 2664 1249 2704
rect 1265 2664 1269 2704
rect 1285 2664 1289 2704
rect 1371 2664 1375 2704
rect 1391 2664 1395 2704
rect 1411 2664 1415 2704
rect 1525 2664 1529 2704
rect 1545 2664 1549 2684
rect 1565 2664 1569 2684
rect 1651 2664 1655 2684
rect 1671 2664 1675 2684
rect 1795 2664 1799 2704
rect 1815 2664 1819 2704
rect 1825 2664 1829 2704
rect 1953 2664 1957 2704
rect 1963 2664 1967 2704
rect 2051 2664 2055 2704
rect 2071 2664 2075 2704
rect 2091 2664 2095 2704
rect 2215 2664 2219 2704
rect 2235 2664 2239 2704
rect 2245 2664 2249 2704
rect 2353 2664 2357 2704
rect 2363 2664 2367 2704
rect 2471 2664 2475 2684
rect 2491 2664 2495 2684
rect 2628 2664 2632 2724
rect 2636 2664 2640 2724
rect 2644 2664 2648 2724
rect 2755 2664 2759 2704
rect 2775 2664 2779 2704
rect 2785 2664 2789 2704
rect 2891 2664 2895 2704
rect 2911 2664 2915 2704
rect 2931 2664 2935 2704
rect 3068 2664 3072 2724
rect 3076 2664 3080 2724
rect 3084 2664 3088 2724
rect 3173 2664 3177 2704
rect 3183 2664 3187 2704
rect 3305 2664 3309 2704
rect 3325 2664 3329 2704
rect 3345 2664 3349 2704
rect 3455 2664 3459 2704
rect 3475 2664 3479 2704
rect 3485 2664 3489 2704
rect 3571 2664 3575 2684
rect 3591 2664 3595 2684
rect 3692 2664 3696 2724
rect 3700 2664 3704 2724
rect 3708 2664 3712 2724
rect 3833 2664 3837 2704
rect 3843 2664 3847 2704
rect 3965 2664 3969 2704
rect 4065 2664 4069 2704
rect 4085 2664 4089 2704
rect 4105 2664 4109 2704
rect 4193 2664 4197 2704
rect 4203 2664 4207 2704
rect 4311 2664 4315 2704
rect 4411 2664 4415 2684
rect 4471 2664 4475 2704
rect 4493 2664 4497 2684
rect 4503 2664 4507 2684
rect 4523 2664 4527 2684
rect 4531 2664 4535 2684
rect 4577 2664 4581 2684
rect 4599 2664 4603 2684
rect 4609 2664 4613 2684
rect 4631 2664 4635 2684
rect 4641 2664 4645 2684
rect 4661 2664 4665 2704
rect 4715 2664 4719 2704
rect 4735 2664 4739 2684
rect 4745 2664 4749 2684
rect 4767 2664 4771 2684
rect 4777 2664 4781 2684
rect 4799 2664 4803 2684
rect 4845 2664 4849 2684
rect 4853 2664 4857 2684
rect 4873 2664 4877 2684
rect 4883 2664 4887 2684
rect 4905 2664 4909 2704
rect 5011 2664 5015 2704
rect 5031 2664 5035 2704
rect 5051 2664 5055 2704
rect 5153 2664 5157 2704
rect 5163 2664 5167 2704
rect 5271 2664 5275 2704
rect 5291 2664 5295 2704
rect 5351 2664 5355 2704
rect 5373 2664 5377 2684
rect 5383 2664 5387 2684
rect 5403 2664 5407 2684
rect 5411 2664 5415 2684
rect 5457 2664 5461 2684
rect 5479 2664 5483 2684
rect 5489 2664 5493 2684
rect 5511 2664 5515 2684
rect 5521 2664 5525 2684
rect 5541 2664 5545 2704
rect 5631 2664 5635 2704
rect 5651 2664 5655 2704
rect 5671 2664 5675 2704
rect 85 2616 89 2636
rect 171 2616 175 2636
rect 292 2616 296 2636
rect 314 2596 318 2636
rect 322 2596 326 2636
rect 412 2576 416 2636
rect 420 2576 424 2636
rect 428 2576 432 2636
rect 551 2616 555 2636
rect 651 2616 655 2636
rect 671 2616 675 2636
rect 771 2596 775 2636
rect 791 2596 795 2636
rect 811 2596 815 2636
rect 934 2596 938 2636
rect 942 2596 946 2636
rect 964 2616 968 2636
rect 1085 2596 1089 2636
rect 1105 2596 1109 2636
rect 1125 2596 1129 2636
rect 1233 2596 1237 2636
rect 1243 2596 1247 2636
rect 1331 2596 1335 2636
rect 1341 2596 1345 2636
rect 1361 2596 1365 2636
rect 1508 2576 1512 2636
rect 1516 2576 1520 2636
rect 1524 2576 1528 2636
rect 1611 2616 1615 2636
rect 1711 2596 1715 2636
rect 1731 2596 1735 2636
rect 1751 2596 1755 2636
rect 1865 2596 1869 2636
rect 1885 2596 1889 2636
rect 1905 2596 1909 2636
rect 1991 2596 1995 2636
rect 2011 2596 2015 2636
rect 2031 2596 2035 2636
rect 2168 2576 2172 2636
rect 2176 2576 2180 2636
rect 2184 2576 2188 2636
rect 2292 2616 2296 2636
rect 2314 2596 2318 2636
rect 2322 2596 2326 2636
rect 2413 2596 2417 2636
rect 2423 2596 2427 2636
rect 2565 2596 2569 2636
rect 2585 2596 2589 2636
rect 2605 2596 2609 2636
rect 2691 2596 2695 2636
rect 2711 2596 2715 2636
rect 2731 2596 2735 2636
rect 2852 2616 2856 2636
rect 2874 2596 2878 2636
rect 2882 2596 2886 2636
rect 2985 2616 2989 2636
rect 3071 2596 3075 2636
rect 3091 2596 3095 2636
rect 3111 2596 3115 2636
rect 3233 2596 3237 2636
rect 3243 2596 3247 2636
rect 3388 2576 3392 2636
rect 3396 2576 3400 2636
rect 3404 2576 3408 2636
rect 3491 2596 3495 2636
rect 3501 2596 3505 2636
rect 3521 2596 3525 2636
rect 3633 2596 3637 2636
rect 3643 2596 3647 2636
rect 3754 2596 3758 2636
rect 3762 2596 3766 2636
rect 3782 2596 3786 2636
rect 3790 2596 3794 2636
rect 3911 2616 3915 2636
rect 3931 2616 3935 2636
rect 3999 2616 4003 2636
rect 4047 2596 4051 2636
rect 4059 2596 4063 2636
rect 4084 2596 4088 2636
rect 4096 2596 4100 2636
rect 4149 2616 4153 2636
rect 4169 2616 4173 2636
rect 4214 2616 4218 2636
rect 4234 2616 4238 2636
rect 4284 2616 4288 2636
rect 4304 2616 4308 2636
rect 4324 2616 4328 2636
rect 4374 2596 4378 2636
rect 4386 2596 4390 2636
rect 4410 2596 4414 2636
rect 4422 2596 4426 2636
rect 4474 2596 4478 2636
rect 4486 2596 4490 2636
rect 4510 2596 4514 2636
rect 4522 2596 4526 2636
rect 4572 2616 4576 2636
rect 4592 2616 4596 2636
rect 4612 2616 4616 2636
rect 4662 2616 4666 2636
rect 4682 2616 4686 2636
rect 4727 2616 4731 2636
rect 4747 2616 4751 2636
rect 4800 2596 4804 2636
rect 4812 2596 4816 2636
rect 4837 2596 4841 2636
rect 4849 2596 4853 2636
rect 4897 2616 4901 2636
rect 4955 2596 4959 2636
rect 4975 2616 4979 2636
rect 4985 2616 4989 2636
rect 5007 2616 5011 2636
rect 5017 2616 5021 2636
rect 5039 2616 5043 2636
rect 5085 2616 5089 2636
rect 5093 2616 5097 2636
rect 5113 2616 5117 2636
rect 5123 2616 5127 2636
rect 5145 2596 5149 2636
rect 5245 2596 5249 2636
rect 5265 2596 5269 2636
rect 5285 2596 5289 2636
rect 5305 2596 5309 2636
rect 5325 2596 5329 2636
rect 5345 2596 5349 2636
rect 5365 2596 5369 2636
rect 5385 2596 5389 2636
rect 5491 2596 5495 2636
rect 5511 2596 5515 2636
rect 5531 2596 5535 2636
rect 5551 2596 5555 2636
rect 5571 2596 5575 2636
rect 5591 2596 5595 2636
rect 5611 2596 5615 2636
rect 5631 2596 5635 2636
rect 5731 2596 5735 2636
rect 83 2184 87 2224
rect 105 2184 109 2204
rect 228 2184 232 2244
rect 236 2184 240 2244
rect 244 2184 248 2244
rect 333 2184 337 2224
rect 343 2184 347 2224
rect 451 2184 455 2224
rect 471 2184 475 2224
rect 491 2184 495 2224
rect 605 2184 609 2224
rect 625 2184 629 2224
rect 645 2184 649 2224
rect 788 2184 792 2244
rect 796 2184 800 2244
rect 804 2184 808 2244
rect 913 2184 917 2224
rect 923 2184 927 2224
rect 1025 2184 1029 2224
rect 1045 2184 1049 2204
rect 1065 2184 1069 2204
rect 1151 2184 1155 2224
rect 1288 2184 1292 2244
rect 1296 2184 1300 2244
rect 1304 2184 1308 2244
rect 1412 2184 1416 2204
rect 1434 2184 1438 2224
rect 1442 2184 1446 2224
rect 1565 2184 1569 2224
rect 1585 2184 1589 2224
rect 1605 2184 1609 2224
rect 1712 2184 1716 2204
rect 1734 2184 1738 2224
rect 1742 2184 1746 2224
rect 1868 2184 1872 2244
rect 1876 2184 1880 2244
rect 1884 2184 1888 2244
rect 2008 2184 2012 2244
rect 2016 2184 2020 2244
rect 2024 2184 2028 2244
rect 2079 2184 2083 2204
rect 2127 2184 2131 2224
rect 2139 2184 2143 2224
rect 2164 2184 2168 2224
rect 2176 2184 2180 2224
rect 2229 2184 2233 2204
rect 2249 2184 2253 2204
rect 2294 2184 2298 2204
rect 2314 2184 2318 2204
rect 2364 2184 2368 2204
rect 2384 2184 2388 2204
rect 2404 2184 2408 2204
rect 2454 2184 2458 2224
rect 2466 2184 2470 2224
rect 2490 2184 2494 2224
rect 2502 2184 2506 2224
rect 2603 2184 2607 2224
rect 2625 2184 2629 2204
rect 2731 2184 2735 2224
rect 2751 2184 2755 2224
rect 2771 2184 2775 2224
rect 2871 2184 2875 2224
rect 2891 2184 2895 2224
rect 2911 2184 2915 2224
rect 3033 2184 3037 2224
rect 3043 2184 3047 2224
rect 3153 2184 3157 2224
rect 3163 2184 3167 2224
rect 3292 2184 3296 2204
rect 3314 2184 3318 2224
rect 3322 2184 3326 2224
rect 3411 2184 3415 2204
rect 3431 2184 3435 2204
rect 3551 2184 3555 2224
rect 3571 2184 3575 2224
rect 3591 2184 3595 2224
rect 3693 2184 3697 2224
rect 3703 2184 3707 2224
rect 3811 2184 3815 2204
rect 3833 2184 3837 2224
rect 3899 2184 3903 2204
rect 3947 2184 3951 2224
rect 3959 2184 3963 2224
rect 3984 2184 3988 2224
rect 3996 2184 4000 2224
rect 4049 2184 4053 2204
rect 4069 2184 4073 2204
rect 4114 2184 4118 2204
rect 4134 2184 4138 2204
rect 4184 2184 4188 2204
rect 4204 2184 4208 2204
rect 4224 2184 4228 2204
rect 4274 2184 4278 2224
rect 4286 2184 4290 2224
rect 4310 2184 4314 2224
rect 4322 2184 4326 2224
rect 4411 2184 4415 2224
rect 4421 2184 4425 2224
rect 4441 2184 4445 2224
rect 4554 2184 4558 2224
rect 4562 2184 4566 2224
rect 4582 2184 4586 2224
rect 4590 2184 4594 2224
rect 4713 2184 4717 2224
rect 4723 2184 4727 2224
rect 4843 2184 4847 2224
rect 4865 2184 4869 2204
rect 4951 2184 4955 2204
rect 5054 2184 5058 2224
rect 5062 2184 5066 2224
rect 5082 2184 5086 2224
rect 5090 2184 5094 2224
rect 5213 2184 5217 2224
rect 5223 2184 5227 2224
rect 5331 2184 5335 2224
rect 5433 2184 5437 2224
rect 5443 2184 5447 2224
rect 5551 2184 5555 2204
rect 5651 2192 5655 2212
rect 5671 2192 5675 2232
rect 5681 2192 5685 2232
rect 5701 2192 5705 2232
rect 5711 2192 5715 2232
rect 103 2116 107 2156
rect 125 2136 129 2156
rect 268 2096 272 2156
rect 276 2096 280 2156
rect 284 2096 288 2156
rect 374 2116 378 2156
rect 382 2116 386 2156
rect 404 2136 408 2156
rect 525 2136 529 2156
rect 625 2116 629 2156
rect 645 2116 649 2156
rect 665 2116 669 2156
rect 772 2136 776 2156
rect 794 2116 798 2156
rect 802 2116 806 2156
rect 892 2096 896 2156
rect 900 2096 904 2156
rect 908 2096 912 2156
rect 1088 2096 1092 2156
rect 1096 2096 1100 2156
rect 1104 2096 1108 2156
rect 1205 2116 1209 2156
rect 1225 2116 1229 2156
rect 1245 2116 1249 2156
rect 1345 2116 1349 2156
rect 1365 2116 1369 2156
rect 1385 2116 1389 2156
rect 1492 2136 1496 2156
rect 1514 2116 1518 2156
rect 1522 2116 1526 2156
rect 1648 2096 1652 2156
rect 1656 2096 1660 2156
rect 1664 2096 1668 2156
rect 1751 2116 1755 2156
rect 1771 2116 1775 2156
rect 1791 2116 1795 2156
rect 1894 2116 1898 2156
rect 1902 2116 1906 2156
rect 1924 2136 1928 2156
rect 2105 2136 2109 2156
rect 2125 2136 2129 2156
rect 2145 2136 2149 2156
rect 2288 2096 2292 2156
rect 2296 2096 2300 2156
rect 2304 2096 2308 2156
rect 2359 2136 2363 2156
rect 2407 2116 2411 2156
rect 2419 2116 2423 2156
rect 2444 2116 2448 2156
rect 2456 2116 2460 2156
rect 2509 2136 2513 2156
rect 2529 2136 2533 2156
rect 2574 2136 2578 2156
rect 2594 2136 2598 2156
rect 2644 2136 2648 2156
rect 2664 2136 2668 2156
rect 2684 2136 2688 2156
rect 2734 2116 2738 2156
rect 2746 2116 2750 2156
rect 2770 2116 2774 2156
rect 2782 2116 2786 2156
rect 2871 2116 2875 2156
rect 2891 2116 2895 2156
rect 2911 2116 2915 2156
rect 3033 2116 3037 2156
rect 3043 2116 3047 2156
rect 3133 2116 3137 2156
rect 3143 2116 3147 2156
rect 3271 2136 3275 2156
rect 3291 2136 3295 2156
rect 3415 2116 3419 2156
rect 3435 2116 3439 2156
rect 3445 2116 3449 2156
rect 3534 2116 3538 2156
rect 3542 2116 3546 2156
rect 3564 2136 3568 2156
rect 3705 2116 3709 2156
rect 3812 2096 3816 2156
rect 3820 2096 3824 2156
rect 3828 2096 3832 2156
rect 3971 2116 3975 2156
rect 4115 2116 4119 2156
rect 4135 2116 4139 2156
rect 4145 2116 4149 2156
rect 4253 2116 4257 2156
rect 4263 2116 4267 2156
rect 4365 2116 4369 2156
rect 4385 2116 4389 2156
rect 4405 2116 4409 2156
rect 4491 2116 4495 2156
rect 4511 2116 4515 2156
rect 4531 2116 4535 2156
rect 4633 2116 4637 2156
rect 4643 2116 4647 2156
rect 4753 2116 4757 2156
rect 4763 2116 4767 2156
rect 4905 2116 4909 2156
rect 4925 2116 4929 2156
rect 4945 2116 4949 2156
rect 5045 2116 5049 2156
rect 5065 2116 5069 2156
rect 5085 2116 5089 2156
rect 5171 2136 5175 2156
rect 5271 2136 5275 2156
rect 5291 2136 5295 2156
rect 5393 2116 5397 2156
rect 5403 2116 5407 2156
rect 5511 2136 5515 2156
rect 5625 2136 5629 2156
rect 5711 2116 5715 2156
rect 5731 2116 5735 2156
rect 5751 2116 5755 2156
rect 108 1704 112 1764
rect 116 1704 120 1764
rect 124 1704 128 1764
rect 214 1704 218 1744
rect 222 1704 226 1744
rect 244 1704 248 1724
rect 365 1704 369 1744
rect 385 1704 389 1744
rect 405 1704 409 1744
rect 528 1704 532 1764
rect 536 1704 540 1764
rect 544 1704 548 1764
rect 665 1704 669 1724
rect 685 1704 689 1724
rect 774 1704 778 1744
rect 782 1704 786 1744
rect 804 1704 808 1724
rect 945 1704 949 1724
rect 1065 1704 1069 1744
rect 1085 1704 1089 1744
rect 1105 1704 1109 1744
rect 1205 1704 1209 1744
rect 1225 1704 1229 1744
rect 1245 1704 1249 1744
rect 1345 1704 1349 1724
rect 1445 1704 1449 1744
rect 1465 1704 1469 1744
rect 1485 1704 1489 1744
rect 1571 1704 1575 1744
rect 1591 1704 1595 1744
rect 1611 1704 1615 1744
rect 1725 1704 1729 1744
rect 1745 1704 1749 1744
rect 1765 1704 1769 1744
rect 1873 1704 1877 1744
rect 1883 1704 1887 1744
rect 1993 1704 1997 1744
rect 2003 1704 2007 1744
rect 2125 1704 2129 1744
rect 2145 1704 2149 1744
rect 2199 1704 2203 1724
rect 2247 1704 2251 1744
rect 2259 1704 2263 1744
rect 2284 1704 2288 1744
rect 2296 1704 2300 1744
rect 2349 1704 2353 1724
rect 2369 1704 2373 1724
rect 2414 1704 2418 1724
rect 2434 1704 2438 1724
rect 2484 1704 2488 1724
rect 2504 1704 2508 1724
rect 2524 1704 2528 1724
rect 2574 1704 2578 1744
rect 2586 1704 2590 1744
rect 2610 1704 2614 1744
rect 2622 1704 2626 1744
rect 2713 1704 2717 1744
rect 2723 1704 2727 1744
rect 2868 1704 2872 1764
rect 2876 1704 2880 1764
rect 2884 1704 2888 1764
rect 2985 1704 2989 1744
rect 3005 1704 3009 1744
rect 3025 1704 3029 1744
rect 3111 1704 3115 1724
rect 3131 1704 3135 1724
rect 3231 1712 3235 1732
rect 3251 1712 3255 1752
rect 3261 1712 3265 1752
rect 3281 1712 3285 1752
rect 3291 1712 3295 1752
rect 3405 1704 3409 1724
rect 3491 1704 3495 1744
rect 3511 1704 3515 1744
rect 3531 1704 3535 1744
rect 3551 1704 3555 1744
rect 3665 1704 3669 1744
rect 3685 1704 3689 1744
rect 3705 1704 3709 1744
rect 3825 1704 3829 1744
rect 3845 1704 3849 1744
rect 3865 1704 3869 1744
rect 3951 1704 3955 1744
rect 3971 1704 3975 1744
rect 3991 1704 3995 1744
rect 4113 1704 4117 1744
rect 4123 1704 4127 1744
rect 4246 1704 4250 1744
rect 4254 1704 4258 1744
rect 4274 1704 4278 1744
rect 4282 1704 4286 1744
rect 4393 1704 4397 1744
rect 4403 1704 4407 1744
rect 4491 1704 4495 1744
rect 4511 1704 4515 1744
rect 4531 1704 4535 1744
rect 4655 1704 4659 1744
rect 4675 1704 4679 1744
rect 4685 1704 4689 1744
rect 4785 1704 4789 1724
rect 4805 1704 4809 1724
rect 4913 1704 4917 1744
rect 4923 1704 4927 1744
rect 5046 1704 5050 1744
rect 5054 1704 5058 1744
rect 5074 1704 5078 1744
rect 5082 1704 5086 1744
rect 5185 1704 5189 1724
rect 5285 1704 5289 1724
rect 5305 1704 5309 1724
rect 5391 1704 5395 1744
rect 5411 1704 5415 1744
rect 5431 1704 5435 1744
rect 5545 1704 5549 1744
rect 5565 1704 5569 1744
rect 5585 1704 5589 1744
rect 5671 1704 5675 1744
rect 5691 1704 5695 1744
rect 92 1616 96 1676
rect 100 1616 104 1676
rect 108 1616 112 1676
rect 268 1616 272 1676
rect 276 1616 280 1676
rect 284 1616 288 1676
rect 374 1636 378 1676
rect 382 1636 386 1676
rect 404 1656 408 1676
rect 532 1656 536 1676
rect 554 1636 558 1676
rect 562 1636 566 1676
rect 653 1636 657 1676
rect 663 1636 667 1676
rect 771 1656 775 1676
rect 885 1636 889 1676
rect 905 1636 909 1676
rect 925 1636 929 1676
rect 1048 1616 1052 1676
rect 1056 1616 1060 1676
rect 1064 1616 1068 1676
rect 1173 1636 1177 1676
rect 1183 1636 1187 1676
rect 1291 1656 1295 1676
rect 1311 1656 1315 1676
rect 1423 1636 1427 1676
rect 1445 1656 1449 1676
rect 1565 1656 1569 1676
rect 1654 1636 1658 1676
rect 1662 1636 1666 1676
rect 1682 1636 1686 1676
rect 1690 1636 1694 1676
rect 1779 1656 1783 1676
rect 1827 1636 1831 1676
rect 1839 1636 1843 1676
rect 1864 1636 1868 1676
rect 1876 1636 1880 1676
rect 1929 1656 1933 1676
rect 1949 1656 1953 1676
rect 1994 1656 1998 1676
rect 2014 1656 2018 1676
rect 2064 1656 2068 1676
rect 2084 1656 2088 1676
rect 2104 1656 2108 1676
rect 2154 1636 2158 1676
rect 2166 1636 2170 1676
rect 2190 1636 2194 1676
rect 2202 1636 2206 1676
rect 2311 1636 2315 1676
rect 2331 1636 2335 1676
rect 2351 1636 2355 1676
rect 2453 1636 2457 1676
rect 2463 1636 2467 1676
rect 2585 1636 2589 1676
rect 2605 1636 2609 1676
rect 2625 1636 2629 1676
rect 2733 1636 2737 1676
rect 2743 1636 2747 1676
rect 2845 1636 2849 1676
rect 2865 1636 2869 1676
rect 2885 1636 2889 1676
rect 2985 1636 2989 1676
rect 3005 1636 3009 1676
rect 3025 1636 3029 1676
rect 3074 1636 3078 1676
rect 3086 1636 3090 1676
rect 3110 1636 3114 1676
rect 3122 1636 3126 1676
rect 3172 1656 3176 1676
rect 3192 1656 3196 1676
rect 3212 1656 3216 1676
rect 3262 1656 3266 1676
rect 3282 1656 3286 1676
rect 3327 1656 3331 1676
rect 3347 1656 3351 1676
rect 3400 1636 3404 1676
rect 3412 1636 3416 1676
rect 3437 1636 3441 1676
rect 3449 1636 3453 1676
rect 3497 1656 3501 1676
rect 3612 1656 3616 1676
rect 3634 1636 3638 1676
rect 3642 1636 3646 1676
rect 3731 1636 3735 1676
rect 3751 1636 3755 1676
rect 3771 1636 3775 1676
rect 3883 1636 3887 1676
rect 3905 1656 3909 1676
rect 4015 1636 4019 1676
rect 4035 1636 4039 1676
rect 4045 1636 4049 1676
rect 4133 1636 4137 1676
rect 4143 1636 4147 1676
rect 4286 1636 4290 1676
rect 4294 1636 4298 1676
rect 4314 1636 4318 1676
rect 4322 1636 4326 1676
rect 4446 1636 4450 1676
rect 4454 1636 4458 1676
rect 4474 1636 4478 1676
rect 4482 1636 4486 1676
rect 4594 1636 4598 1676
rect 4602 1636 4606 1676
rect 4622 1636 4626 1676
rect 4630 1636 4634 1676
rect 4753 1636 4757 1676
rect 4763 1636 4767 1676
rect 4871 1636 4875 1676
rect 4891 1636 4895 1676
rect 4911 1636 4915 1676
rect 5035 1636 5039 1676
rect 5055 1636 5059 1676
rect 5065 1636 5069 1676
rect 5172 1616 5176 1676
rect 5180 1616 5184 1676
rect 5188 1616 5192 1676
rect 5314 1636 5318 1676
rect 5322 1636 5326 1676
rect 5342 1636 5346 1676
rect 5350 1636 5354 1676
rect 5473 1636 5477 1676
rect 5483 1636 5487 1676
rect 5592 1616 5596 1676
rect 5600 1616 5604 1676
rect 5608 1616 5612 1676
rect 5765 1636 5769 1676
rect 108 1224 112 1284
rect 116 1224 120 1284
rect 124 1224 128 1284
rect 214 1224 218 1264
rect 222 1224 226 1264
rect 244 1224 248 1244
rect 388 1224 392 1284
rect 396 1224 400 1284
rect 404 1224 408 1284
rect 505 1224 509 1264
rect 525 1224 529 1264
rect 545 1224 549 1264
rect 645 1224 649 1264
rect 665 1224 669 1264
rect 685 1224 689 1264
rect 815 1224 819 1264
rect 835 1224 839 1264
rect 845 1224 849 1264
rect 933 1224 937 1264
rect 943 1224 947 1264
rect 1065 1224 1069 1244
rect 1152 1224 1156 1284
rect 1160 1224 1164 1284
rect 1168 1224 1172 1284
rect 1293 1224 1297 1264
rect 1303 1224 1307 1264
rect 1433 1224 1437 1264
rect 1443 1224 1447 1264
rect 1553 1224 1557 1264
rect 1563 1224 1567 1264
rect 1708 1224 1712 1284
rect 1716 1224 1720 1284
rect 1724 1224 1728 1284
rect 1813 1224 1817 1264
rect 1823 1224 1827 1264
rect 1968 1224 1972 1284
rect 1976 1224 1980 1284
rect 1984 1224 1988 1284
rect 2085 1224 2089 1244
rect 2228 1224 2232 1284
rect 2236 1224 2240 1284
rect 2244 1224 2248 1284
rect 2368 1224 2372 1284
rect 2376 1224 2380 1284
rect 2384 1224 2388 1284
rect 2471 1224 2475 1244
rect 2605 1224 2609 1264
rect 2625 1224 2629 1264
rect 2645 1224 2649 1264
rect 2734 1224 2738 1264
rect 2742 1224 2746 1264
rect 2764 1224 2768 1244
rect 2885 1224 2889 1264
rect 2905 1224 2909 1264
rect 2925 1224 2929 1264
rect 3025 1224 3029 1264
rect 3045 1224 3049 1264
rect 3065 1224 3069 1264
rect 3165 1224 3169 1264
rect 3185 1224 3189 1264
rect 3205 1224 3209 1264
rect 3305 1224 3309 1244
rect 3391 1224 3395 1244
rect 3503 1224 3507 1264
rect 3525 1224 3529 1244
rect 3652 1224 3656 1244
rect 3674 1224 3678 1264
rect 3682 1224 3686 1264
rect 3771 1224 3775 1264
rect 3791 1224 3795 1264
rect 3811 1224 3815 1264
rect 3925 1224 3929 1244
rect 4025 1224 4029 1264
rect 4045 1224 4049 1264
rect 4065 1224 4069 1264
rect 4165 1224 4169 1264
rect 4185 1224 4189 1264
rect 4205 1224 4209 1264
rect 4312 1224 4316 1244
rect 4334 1224 4338 1264
rect 4342 1224 4346 1264
rect 4445 1224 4449 1264
rect 4465 1224 4469 1264
rect 4485 1224 4489 1264
rect 4591 1224 4595 1264
rect 4611 1224 4615 1264
rect 4631 1224 4635 1264
rect 4733 1224 4737 1264
rect 4743 1224 4747 1264
rect 4851 1224 4855 1264
rect 4871 1224 4875 1264
rect 4891 1224 4895 1264
rect 4991 1224 4995 1244
rect 5011 1224 5015 1244
rect 5113 1224 5117 1264
rect 5123 1224 5127 1264
rect 5253 1224 5257 1264
rect 5263 1224 5267 1264
rect 5365 1224 5369 1264
rect 5385 1224 5389 1264
rect 5405 1224 5409 1264
rect 5491 1224 5495 1264
rect 5511 1224 5515 1264
rect 5531 1224 5535 1264
rect 5651 1224 5655 1264
rect 5671 1224 5675 1264
rect 5691 1224 5695 1264
rect 85 1176 89 1196
rect 174 1156 178 1196
rect 182 1156 186 1196
rect 204 1176 208 1196
rect 311 1156 315 1196
rect 331 1156 335 1196
rect 351 1156 355 1196
rect 451 1156 455 1196
rect 471 1156 475 1196
rect 491 1156 495 1196
rect 628 1136 632 1196
rect 636 1136 640 1196
rect 644 1136 648 1196
rect 731 1156 735 1196
rect 751 1156 755 1196
rect 771 1156 775 1196
rect 894 1156 898 1196
rect 902 1156 906 1196
rect 924 1176 928 1196
rect 1045 1156 1049 1196
rect 1065 1156 1069 1196
rect 1085 1156 1089 1196
rect 1185 1176 1189 1196
rect 1274 1156 1278 1196
rect 1282 1156 1286 1196
rect 1304 1176 1308 1196
rect 1425 1176 1429 1196
rect 1525 1176 1529 1196
rect 1545 1176 1549 1196
rect 1651 1176 1655 1196
rect 1788 1136 1792 1196
rect 1796 1136 1800 1196
rect 1804 1136 1808 1196
rect 1913 1156 1917 1196
rect 1923 1156 1927 1196
rect 2025 1156 2029 1196
rect 2045 1156 2049 1196
rect 2065 1156 2069 1196
rect 2188 1136 2192 1196
rect 2196 1136 2200 1196
rect 2204 1136 2208 1196
rect 2328 1136 2332 1196
rect 2336 1136 2340 1196
rect 2344 1136 2348 1196
rect 2445 1156 2449 1196
rect 2465 1156 2469 1196
rect 2485 1156 2489 1196
rect 2608 1136 2612 1196
rect 2616 1136 2620 1196
rect 2624 1136 2628 1196
rect 2731 1176 2735 1196
rect 2831 1176 2835 1196
rect 2851 1176 2855 1196
rect 2951 1176 2955 1196
rect 2971 1176 2975 1196
rect 3071 1156 3075 1196
rect 3081 1156 3085 1196
rect 3101 1156 3105 1196
rect 3225 1176 3229 1196
rect 3245 1176 3249 1196
rect 3365 1176 3369 1196
rect 3385 1176 3389 1196
rect 3485 1176 3489 1196
rect 3585 1156 3589 1196
rect 3605 1156 3609 1196
rect 3625 1156 3629 1196
rect 3725 1156 3729 1196
rect 3745 1156 3749 1196
rect 3765 1156 3769 1196
rect 3853 1156 3857 1196
rect 3863 1156 3867 1196
rect 3973 1156 3977 1196
rect 3983 1156 3987 1196
rect 4091 1176 4095 1196
rect 4111 1176 4115 1196
rect 4211 1176 4215 1196
rect 4332 1176 4336 1196
rect 4354 1156 4358 1196
rect 4362 1156 4366 1196
rect 4485 1156 4489 1196
rect 4505 1156 4509 1196
rect 4525 1156 4529 1196
rect 4632 1176 4636 1196
rect 4654 1156 4658 1196
rect 4662 1156 4666 1196
rect 4751 1156 4755 1196
rect 4771 1156 4775 1196
rect 4791 1156 4795 1196
rect 4891 1176 4895 1196
rect 4913 1156 4917 1196
rect 5011 1176 5015 1196
rect 5111 1176 5115 1196
rect 5233 1156 5237 1196
rect 5243 1156 5247 1196
rect 5365 1156 5369 1196
rect 5385 1156 5389 1196
rect 5405 1156 5409 1196
rect 5491 1176 5495 1196
rect 5511 1176 5515 1196
rect 5648 1136 5652 1196
rect 5656 1136 5660 1196
rect 5664 1136 5668 1196
rect 5765 1176 5769 1196
rect 108 744 112 804
rect 116 744 120 804
rect 124 744 128 804
rect 214 744 218 784
rect 222 744 226 784
rect 244 744 248 764
rect 388 744 392 804
rect 396 744 400 804
rect 404 744 408 804
rect 512 744 516 764
rect 534 744 538 784
rect 542 744 546 784
rect 668 744 672 804
rect 676 744 680 804
rect 684 744 688 804
rect 774 744 778 784
rect 782 744 786 784
rect 804 744 808 764
rect 925 744 929 784
rect 945 744 949 784
rect 965 744 969 784
rect 1088 744 1092 804
rect 1096 744 1100 804
rect 1104 744 1108 804
rect 1191 744 1195 784
rect 1211 744 1215 784
rect 1231 744 1235 784
rect 1368 744 1372 804
rect 1376 744 1380 804
rect 1384 744 1388 804
rect 1471 744 1475 764
rect 1573 744 1577 784
rect 1583 744 1587 784
rect 1748 744 1752 804
rect 1756 744 1760 804
rect 1764 744 1768 804
rect 1888 744 1892 804
rect 1896 744 1900 804
rect 1904 744 1908 804
rect 1992 744 1996 804
rect 2000 744 2004 804
rect 2008 744 2012 804
rect 2131 744 2135 784
rect 2151 744 2155 784
rect 2171 744 2175 784
rect 2271 744 2275 784
rect 2281 744 2285 784
rect 2301 744 2305 784
rect 2411 744 2415 764
rect 2533 744 2537 784
rect 2543 744 2547 784
rect 2645 744 2649 784
rect 2665 744 2669 764
rect 2685 744 2689 764
rect 2773 744 2777 784
rect 2783 744 2787 784
rect 2913 744 2917 784
rect 2923 744 2927 784
rect 3031 744 3035 764
rect 3145 744 3149 764
rect 3273 744 3277 784
rect 3283 744 3287 784
rect 3405 744 3409 764
rect 3425 744 3429 764
rect 3525 744 3529 764
rect 3545 744 3549 764
rect 3652 744 3656 764
rect 3674 744 3678 784
rect 3682 744 3686 784
rect 3785 744 3789 764
rect 3885 744 3889 784
rect 3905 744 3909 784
rect 3925 744 3929 784
rect 4013 744 4017 784
rect 4023 744 4027 784
rect 4145 744 4149 784
rect 4165 744 4169 784
rect 4185 744 4189 784
rect 4285 744 4289 784
rect 4305 744 4309 784
rect 4325 744 4329 784
rect 4431 744 4435 764
rect 4545 744 4549 784
rect 4565 744 4569 784
rect 4585 744 4589 784
rect 4674 744 4678 784
rect 4682 744 4686 784
rect 4704 744 4708 764
rect 4823 744 4827 784
rect 4845 744 4849 764
rect 4945 744 4949 784
rect 4965 744 4969 784
rect 4985 744 4989 784
rect 5074 744 5078 784
rect 5082 744 5086 784
rect 5104 744 5108 764
rect 5225 744 5229 784
rect 5245 744 5249 764
rect 5265 744 5269 764
rect 5385 744 5389 764
rect 5506 744 5510 784
rect 5514 744 5518 784
rect 5534 744 5538 784
rect 5542 744 5546 784
rect 5651 744 5655 784
rect 5671 744 5675 784
rect 5691 744 5695 784
rect 108 656 112 716
rect 116 656 120 716
rect 124 656 128 716
rect 252 696 256 716
rect 274 676 278 716
rect 282 676 286 716
rect 408 656 412 716
rect 416 656 420 716
rect 424 656 428 716
rect 525 676 529 716
rect 545 676 549 716
rect 565 676 569 716
rect 654 676 658 716
rect 662 676 666 716
rect 684 696 688 716
rect 793 676 797 716
rect 803 676 807 716
rect 945 676 949 716
rect 965 676 969 716
rect 985 676 989 716
rect 1108 656 1112 716
rect 1116 656 1120 716
rect 1124 656 1128 716
rect 1214 676 1218 716
rect 1222 676 1226 716
rect 1244 696 1248 716
rect 1372 696 1376 716
rect 1394 676 1398 716
rect 1402 676 1406 716
rect 1512 656 1516 716
rect 1520 656 1524 716
rect 1528 656 1532 716
rect 1665 676 1669 716
rect 1685 676 1689 716
rect 1705 676 1709 716
rect 1828 656 1832 716
rect 1836 656 1840 716
rect 1844 656 1848 716
rect 1934 676 1938 716
rect 1942 676 1946 716
rect 1964 696 1968 716
rect 2085 696 2089 716
rect 2105 696 2109 716
rect 2205 676 2209 716
rect 2225 696 2229 716
rect 2245 696 2249 716
rect 2331 676 2335 716
rect 2341 676 2345 716
rect 2361 676 2365 716
rect 2473 676 2477 716
rect 2483 676 2487 716
rect 2613 676 2617 716
rect 2623 676 2627 716
rect 2725 696 2729 716
rect 2745 696 2749 716
rect 2831 676 2835 716
rect 2851 676 2855 716
rect 2871 676 2875 716
rect 2993 676 2997 716
rect 3003 676 3007 716
rect 3094 676 3098 716
rect 3102 676 3106 716
rect 3124 696 3128 716
rect 3268 656 3272 716
rect 3276 656 3280 716
rect 3284 656 3288 716
rect 3373 676 3377 716
rect 3383 676 3387 716
rect 3505 676 3509 716
rect 3525 676 3529 716
rect 3545 676 3549 716
rect 3633 676 3637 716
rect 3643 676 3647 716
rect 3765 676 3769 716
rect 3785 676 3789 716
rect 3805 676 3809 716
rect 3891 676 3895 716
rect 3911 676 3915 716
rect 3931 676 3935 716
rect 4034 676 4038 716
rect 4042 676 4046 716
rect 4064 696 4068 716
rect 4191 676 4195 716
rect 4211 676 4215 716
rect 4231 676 4235 716
rect 4345 696 4349 716
rect 4452 696 4456 716
rect 4474 676 4478 716
rect 4482 676 4486 716
rect 4585 676 4589 716
rect 4605 676 4609 716
rect 4625 676 4629 716
rect 4725 676 4729 716
rect 4745 676 4749 716
rect 4765 676 4769 716
rect 4871 676 4875 716
rect 4891 676 4895 716
rect 4911 676 4915 716
rect 5011 696 5015 716
rect 5131 696 5135 716
rect 5153 676 5157 716
rect 5265 676 5269 716
rect 5285 676 5289 716
rect 5305 676 5309 716
rect 5391 676 5395 716
rect 5411 676 5415 716
rect 5431 676 5435 716
rect 5545 676 5549 716
rect 5565 676 5569 716
rect 5585 676 5589 716
rect 5671 696 5675 716
rect 5691 696 5695 716
rect 108 264 112 324
rect 116 264 120 324
rect 124 264 128 324
rect 225 264 229 304
rect 245 264 249 304
rect 265 264 269 304
rect 385 264 389 304
rect 405 264 409 304
rect 425 264 429 304
rect 548 264 552 324
rect 556 264 560 324
rect 564 264 568 324
rect 675 264 679 304
rect 695 264 699 304
rect 705 264 709 304
rect 828 264 832 324
rect 836 264 840 324
rect 844 264 848 324
rect 952 264 956 284
rect 974 264 978 304
rect 982 264 986 304
rect 1072 264 1076 324
rect 1080 264 1084 324
rect 1088 264 1092 324
rect 1225 264 1229 304
rect 1245 264 1249 284
rect 1265 264 1269 284
rect 1388 264 1392 324
rect 1396 264 1400 324
rect 1404 264 1408 324
rect 1525 264 1529 284
rect 1625 264 1629 304
rect 1645 264 1649 304
rect 1665 264 1669 304
rect 1775 264 1779 304
rect 1795 264 1799 304
rect 1805 264 1809 304
rect 1891 264 1895 284
rect 1911 264 1915 284
rect 2031 264 2035 284
rect 2145 264 2149 304
rect 2165 264 2169 304
rect 2185 264 2189 304
rect 2292 264 2296 284
rect 2314 264 2318 304
rect 2322 264 2326 304
rect 2425 264 2429 284
rect 2548 264 2552 324
rect 2556 264 2560 324
rect 2564 264 2568 324
rect 2651 264 2655 304
rect 2671 264 2675 304
rect 2691 264 2695 304
rect 2805 264 2809 284
rect 2905 264 2909 284
rect 2925 264 2929 284
rect 3011 264 3015 284
rect 3132 264 3136 284
rect 3154 264 3158 304
rect 3162 264 3166 304
rect 3274 264 3278 304
rect 3282 264 3286 304
rect 3304 264 3308 284
rect 3425 264 3429 284
rect 3531 264 3535 304
rect 3551 264 3555 304
rect 3571 264 3575 304
rect 3674 264 3678 304
rect 3682 264 3686 304
rect 3704 264 3708 284
rect 3848 264 3852 324
rect 3856 264 3860 324
rect 3864 264 3868 324
rect 3953 264 3957 304
rect 3963 264 3967 304
rect 4128 264 4132 324
rect 4136 264 4140 324
rect 4144 264 4148 324
rect 4245 264 4249 304
rect 4265 264 4269 304
rect 4285 264 4289 304
rect 4385 264 4389 284
rect 4493 264 4497 304
rect 4503 264 4507 304
rect 4605 264 4609 304
rect 4625 264 4629 304
rect 4645 264 4649 304
rect 4745 264 4749 284
rect 4845 264 4849 304
rect 4865 264 4869 304
rect 4885 264 4889 304
rect 4971 272 4975 292
rect 4991 272 4995 312
rect 5001 272 5005 312
rect 5021 272 5025 312
rect 5031 272 5035 312
rect 5145 264 5149 304
rect 5165 264 5169 304
rect 5185 264 5189 304
rect 5291 264 5295 304
rect 5311 264 5315 304
rect 5331 264 5335 304
rect 5472 264 5476 284
rect 5494 264 5498 304
rect 5502 264 5506 304
rect 5591 264 5595 304
rect 5611 264 5615 304
rect 5631 264 5635 304
rect 5733 264 5737 304
rect 5743 264 5747 304
rect 108 176 112 236
rect 116 176 120 236
rect 124 176 128 236
rect 214 196 218 236
rect 222 196 226 236
rect 244 216 248 236
rect 392 216 396 236
rect 414 196 418 236
rect 422 196 426 236
rect 525 196 529 236
rect 545 196 549 236
rect 565 196 569 236
rect 651 196 655 236
rect 671 196 675 236
rect 691 196 695 236
rect 828 176 832 236
rect 836 176 840 236
rect 844 176 848 236
rect 931 216 935 236
rect 1031 196 1035 236
rect 1051 196 1055 236
rect 1071 196 1075 236
rect 1174 196 1178 236
rect 1182 196 1186 236
rect 1204 216 1208 236
rect 1311 216 1315 236
rect 1331 216 1335 236
rect 1431 196 1435 236
rect 1441 196 1445 236
rect 1461 196 1465 236
rect 1585 216 1589 236
rect 1685 196 1689 236
rect 1705 196 1709 236
rect 1725 196 1729 236
rect 1833 196 1837 236
rect 1843 196 1847 236
rect 1932 176 1936 236
rect 1940 176 1944 236
rect 1948 176 1952 236
rect 2128 176 2132 236
rect 2136 176 2140 236
rect 2144 176 2148 236
rect 2231 216 2235 236
rect 2253 196 2257 236
rect 2373 196 2377 236
rect 2383 196 2387 236
rect 2471 196 2475 236
rect 2481 196 2485 236
rect 2501 196 2505 236
rect 2632 216 2636 236
rect 2654 196 2658 236
rect 2662 196 2666 236
rect 2775 196 2779 236
rect 2795 196 2799 236
rect 2805 196 2809 236
rect 2913 196 2917 236
rect 2923 196 2927 236
rect 3053 196 3057 236
rect 3063 196 3067 236
rect 3188 176 3192 236
rect 3196 176 3200 236
rect 3204 176 3208 236
rect 3305 216 3309 236
rect 3391 196 3395 236
rect 3411 196 3415 236
rect 3431 196 3435 236
rect 3545 216 3549 236
rect 3653 196 3657 236
rect 3663 196 3667 236
rect 3763 196 3767 236
rect 3785 216 3789 236
rect 3871 216 3875 236
rect 3893 196 3897 236
rect 4013 196 4017 236
rect 4023 196 4027 236
rect 4131 196 4135 236
rect 4141 196 4145 236
rect 4161 196 4165 236
rect 4305 216 4309 236
rect 4325 216 4329 236
rect 4413 196 4417 236
rect 4423 196 4427 236
rect 4568 176 4572 236
rect 4576 176 4580 236
rect 4584 176 4588 236
rect 4705 196 4709 236
rect 4725 196 4729 236
rect 4745 196 4749 236
rect 4833 196 4837 236
rect 4843 196 4847 236
rect 4965 196 4969 236
rect 4985 196 4989 236
rect 5005 196 5009 236
rect 5091 216 5095 236
rect 5111 216 5115 236
rect 5233 196 5237 236
rect 5243 196 5247 236
rect 5331 208 5335 228
rect 5351 188 5355 228
rect 5361 188 5365 228
rect 5381 188 5385 228
rect 5391 188 5395 228
rect 5491 216 5495 236
rect 5605 216 5609 236
rect 5693 196 5697 236
rect 5703 196 5707 236
<< ptransistor >>
rect 90 5716 94 5756
rect 112 5676 116 5756
rect 120 5676 124 5756
rect 216 5676 220 5756
rect 224 5676 228 5756
rect 246 5716 250 5756
rect 385 5676 389 5756
rect 405 5676 409 5756
rect 425 5676 429 5756
rect 511 5716 515 5756
rect 531 5716 535 5756
rect 551 5716 555 5756
rect 670 5716 674 5756
rect 692 5676 696 5756
rect 700 5676 704 5756
rect 805 5716 809 5756
rect 825 5716 829 5756
rect 925 5676 929 5756
rect 945 5676 949 5756
rect 965 5676 969 5756
rect 1071 5676 1075 5756
rect 1079 5676 1083 5756
rect 1235 5676 1239 5756
rect 1255 5676 1259 5756
rect 1265 5676 1269 5756
rect 1361 5676 1365 5756
rect 1383 5716 1387 5756
rect 1405 5716 1409 5756
rect 1505 5716 1509 5756
rect 1525 5716 1529 5756
rect 1545 5716 1549 5756
rect 1665 5676 1669 5756
rect 1685 5676 1689 5756
rect 1705 5676 1709 5756
rect 1805 5716 1809 5756
rect 1825 5716 1829 5756
rect 1845 5716 1849 5756
rect 1931 5716 1935 5756
rect 2050 5716 2054 5756
rect 2072 5676 2076 5756
rect 2080 5676 2084 5756
rect 2176 5676 2180 5756
rect 2184 5676 2188 5756
rect 2206 5716 2210 5756
rect 2311 5676 2315 5756
rect 2331 5676 2335 5756
rect 2351 5676 2355 5756
rect 2465 5716 2469 5756
rect 2485 5716 2489 5756
rect 2585 5716 2589 5756
rect 2605 5716 2609 5756
rect 2625 5716 2629 5756
rect 2725 5716 2729 5756
rect 2745 5716 2749 5756
rect 2765 5716 2769 5756
rect 2851 5716 2855 5756
rect 2871 5716 2875 5756
rect 2985 5716 2989 5756
rect 3090 5716 3094 5756
rect 3112 5676 3116 5756
rect 3120 5676 3124 5756
rect 3241 5676 3245 5756
rect 3263 5716 3267 5756
rect 3285 5716 3289 5756
rect 3397 5676 3401 5756
rect 3405 5676 3409 5756
rect 3505 5716 3509 5756
rect 3525 5716 3529 5756
rect 3545 5716 3549 5756
rect 3665 5716 3669 5756
rect 3765 5716 3769 5756
rect 3851 5716 3855 5756
rect 3956 5676 3960 5756
rect 3964 5676 3968 5756
rect 3986 5716 3990 5756
rect 4091 5716 4095 5756
rect 4151 5676 4155 5756
rect 4173 5736 4177 5756
rect 4181 5736 4185 5756
rect 4201 5716 4205 5756
rect 4209 5716 4213 5756
rect 4255 5716 4259 5756
rect 4275 5716 4279 5756
rect 4287 5716 4291 5756
rect 4307 5716 4311 5756
rect 4321 5716 4325 5756
rect 4341 5676 4345 5756
rect 4470 5716 4474 5756
rect 4492 5676 4496 5756
rect 4500 5676 4504 5756
rect 4605 5676 4609 5756
rect 4625 5676 4629 5756
rect 4645 5676 4649 5756
rect 4665 5676 4669 5756
rect 4685 5676 4689 5756
rect 4705 5676 4709 5756
rect 4725 5676 4729 5756
rect 4745 5676 4749 5756
rect 4845 5716 4849 5756
rect 4950 5716 4954 5756
rect 4972 5676 4976 5756
rect 4980 5676 4984 5756
rect 5085 5716 5089 5756
rect 5105 5716 5109 5756
rect 5191 5716 5195 5756
rect 5211 5716 5215 5756
rect 5316 5676 5320 5756
rect 5324 5676 5328 5756
rect 5346 5716 5350 5756
rect 5451 5716 5455 5756
rect 5551 5716 5555 5756
rect 5571 5716 5575 5756
rect 5671 5716 5675 5756
rect 90 5304 94 5344
rect 112 5304 116 5384
rect 120 5304 124 5384
rect 245 5304 249 5344
rect 265 5304 269 5344
rect 285 5304 289 5344
rect 385 5304 389 5344
rect 405 5304 409 5344
rect 425 5304 429 5344
rect 525 5304 529 5344
rect 545 5304 549 5344
rect 565 5304 569 5344
rect 671 5304 675 5344
rect 691 5304 695 5344
rect 711 5304 715 5344
rect 816 5304 820 5384
rect 824 5304 828 5384
rect 846 5304 850 5344
rect 951 5304 955 5344
rect 971 5304 975 5344
rect 991 5304 995 5344
rect 1105 5304 1109 5384
rect 1125 5304 1129 5384
rect 1145 5304 1149 5384
rect 1231 5304 1235 5344
rect 1251 5304 1255 5344
rect 1271 5304 1275 5344
rect 1391 5304 1395 5384
rect 1399 5304 1403 5384
rect 1525 5304 1529 5344
rect 1545 5304 1549 5344
rect 1565 5304 1569 5344
rect 1656 5304 1660 5384
rect 1664 5304 1668 5384
rect 1686 5304 1690 5344
rect 1805 5304 1809 5344
rect 1825 5304 1829 5344
rect 1845 5304 1849 5344
rect 1945 5304 1949 5344
rect 1965 5304 1969 5344
rect 1985 5304 1989 5344
rect 2071 5304 2075 5344
rect 2091 5304 2095 5344
rect 2225 5304 2229 5344
rect 2321 5304 2325 5384
rect 2343 5304 2347 5344
rect 2365 5304 2369 5344
rect 2456 5304 2460 5384
rect 2464 5304 2468 5384
rect 2486 5304 2490 5344
rect 2625 5304 2629 5344
rect 2645 5304 2649 5344
rect 2665 5304 2669 5344
rect 2765 5304 2769 5344
rect 2785 5304 2789 5344
rect 2805 5304 2809 5344
rect 2896 5304 2900 5384
rect 2904 5304 2908 5384
rect 2926 5304 2930 5344
rect 3031 5304 3035 5344
rect 3131 5304 3135 5344
rect 3151 5304 3155 5344
rect 3271 5304 3275 5344
rect 3291 5304 3295 5344
rect 3311 5304 3315 5344
rect 3411 5304 3415 5344
rect 3431 5304 3435 5344
rect 3531 5304 3535 5384
rect 3541 5304 3545 5384
rect 3561 5304 3565 5384
rect 3685 5304 3689 5344
rect 3705 5304 3709 5344
rect 3725 5304 3729 5344
rect 3825 5304 3829 5384
rect 3845 5304 3849 5384
rect 3865 5304 3869 5384
rect 3951 5304 3955 5344
rect 3971 5304 3975 5344
rect 4090 5304 4094 5344
rect 4112 5304 4116 5384
rect 4120 5304 4124 5384
rect 4225 5304 4229 5344
rect 4245 5304 4249 5344
rect 4345 5304 4349 5344
rect 4365 5304 4369 5344
rect 4385 5304 4389 5344
rect 4491 5304 4495 5384
rect 4511 5304 4515 5384
rect 4531 5304 4535 5384
rect 4631 5304 4635 5344
rect 4736 5304 4740 5384
rect 4744 5304 4748 5384
rect 4766 5304 4770 5344
rect 4831 5304 4835 5384
rect 4853 5304 4857 5324
rect 4861 5304 4865 5324
rect 4881 5304 4885 5344
rect 4889 5304 4893 5344
rect 4935 5304 4939 5344
rect 4955 5304 4959 5344
rect 4967 5304 4971 5344
rect 4987 5304 4991 5344
rect 5001 5304 5005 5344
rect 5021 5304 5025 5384
rect 5111 5304 5115 5344
rect 5171 5304 5175 5384
rect 5193 5304 5197 5324
rect 5201 5304 5205 5324
rect 5221 5304 5225 5344
rect 5229 5304 5233 5344
rect 5275 5304 5279 5344
rect 5295 5304 5299 5344
rect 5307 5304 5311 5344
rect 5327 5304 5331 5344
rect 5341 5304 5345 5344
rect 5361 5304 5365 5384
rect 5456 5304 5460 5384
rect 5464 5304 5468 5384
rect 5486 5304 5490 5344
rect 5611 5304 5615 5344
rect 5631 5304 5635 5344
rect 5731 5304 5735 5344
rect 5751 5304 5755 5344
rect 85 5236 89 5276
rect 105 5236 109 5276
rect 125 5236 129 5276
rect 211 5196 215 5276
rect 231 5196 235 5276
rect 251 5196 255 5276
rect 351 5236 355 5276
rect 465 5236 469 5276
rect 485 5236 489 5276
rect 505 5236 509 5276
rect 591 5196 595 5276
rect 611 5196 615 5276
rect 631 5196 635 5276
rect 745 5196 749 5276
rect 765 5196 769 5276
rect 785 5196 789 5276
rect 871 5236 875 5276
rect 891 5236 895 5276
rect 911 5236 915 5276
rect 1025 5236 1029 5276
rect 1045 5236 1049 5276
rect 1065 5236 1069 5276
rect 1151 5236 1155 5276
rect 1265 5236 1269 5276
rect 1285 5236 1289 5276
rect 1305 5236 1309 5276
rect 1430 5236 1434 5276
rect 1452 5196 1456 5276
rect 1460 5196 1464 5276
rect 1565 5236 1569 5276
rect 1670 5236 1674 5276
rect 1692 5196 1696 5276
rect 1700 5196 1704 5276
rect 1821 5208 1825 5268
rect 1841 5208 1845 5268
rect 1885 5216 1889 5276
rect 1905 5216 1909 5276
rect 1925 5216 1929 5276
rect 1945 5216 1949 5276
rect 2045 5196 2049 5276
rect 2065 5196 2069 5276
rect 2085 5196 2089 5276
rect 2105 5196 2109 5276
rect 2191 5236 2195 5276
rect 2211 5236 2215 5276
rect 2325 5236 2329 5276
rect 2345 5236 2349 5276
rect 2365 5236 2369 5276
rect 2465 5196 2469 5276
rect 2485 5196 2489 5276
rect 2505 5196 2509 5276
rect 2605 5236 2609 5276
rect 2710 5236 2714 5276
rect 2732 5196 2736 5276
rect 2740 5196 2744 5276
rect 2870 5236 2874 5276
rect 2892 5196 2896 5276
rect 2900 5196 2904 5276
rect 3001 5196 3005 5276
rect 3023 5236 3027 5276
rect 3045 5236 3049 5276
rect 3131 5196 3135 5276
rect 3139 5196 3143 5276
rect 3285 5236 3289 5276
rect 3397 5196 3401 5276
rect 3405 5196 3409 5276
rect 3530 5236 3534 5276
rect 3552 5196 3556 5276
rect 3560 5196 3564 5276
rect 3651 5236 3655 5276
rect 3671 5236 3675 5276
rect 3785 5236 3789 5276
rect 3805 5236 3809 5276
rect 3925 5236 3929 5276
rect 3945 5236 3949 5276
rect 4031 5236 4035 5276
rect 4051 5236 4055 5276
rect 4071 5236 4075 5276
rect 4190 5236 4194 5276
rect 4212 5196 4216 5276
rect 4220 5196 4224 5276
rect 4336 5196 4340 5276
rect 4344 5196 4348 5276
rect 4366 5236 4370 5276
rect 4471 5236 4475 5276
rect 4585 5236 4589 5276
rect 4605 5236 4609 5276
rect 4625 5236 4629 5276
rect 4711 5196 4715 5276
rect 4731 5196 4735 5276
rect 4751 5196 4755 5276
rect 4851 5196 4855 5276
rect 4859 5196 4863 5276
rect 4931 5196 4935 5276
rect 4953 5256 4957 5276
rect 4961 5256 4965 5276
rect 4981 5236 4985 5276
rect 4989 5236 4993 5276
rect 5035 5236 5039 5276
rect 5055 5236 5059 5276
rect 5067 5236 5071 5276
rect 5087 5236 5091 5276
rect 5101 5236 5105 5276
rect 5121 5196 5125 5276
rect 5216 5196 5220 5276
rect 5224 5196 5228 5276
rect 5246 5236 5250 5276
rect 5351 5236 5355 5276
rect 5456 5196 5460 5276
rect 5464 5196 5468 5276
rect 5486 5236 5490 5276
rect 5605 5236 5609 5276
rect 5625 5236 5629 5276
rect 5711 5236 5715 5276
rect 5731 5236 5735 5276
rect 90 4824 94 4864
rect 112 4824 116 4904
rect 120 4824 124 4904
rect 225 4824 229 4864
rect 245 4824 249 4864
rect 265 4824 269 4864
rect 351 4824 355 4864
rect 371 4824 375 4864
rect 391 4824 395 4864
rect 496 4824 500 4904
rect 504 4824 508 4904
rect 526 4824 530 4864
rect 645 4824 649 4864
rect 665 4824 669 4864
rect 770 4824 774 4864
rect 792 4824 796 4904
rect 800 4824 804 4904
rect 910 4824 914 4864
rect 932 4824 936 4904
rect 940 4824 944 4904
rect 1045 4824 1049 4904
rect 1065 4824 1069 4904
rect 1085 4824 1089 4904
rect 1190 4824 1194 4864
rect 1212 4824 1216 4904
rect 1220 4824 1224 4904
rect 1325 4824 1329 4864
rect 1425 4824 1429 4864
rect 1445 4824 1449 4864
rect 1565 4824 1569 4864
rect 1585 4824 1589 4864
rect 1605 4824 1609 4864
rect 1710 4824 1714 4864
rect 1732 4824 1736 4904
rect 1740 4824 1744 4904
rect 1831 4824 1835 4904
rect 1851 4824 1855 4904
rect 1871 4824 1875 4904
rect 1971 4824 1975 4864
rect 1991 4824 1995 4864
rect 2105 4824 2109 4904
rect 2125 4824 2129 4904
rect 2145 4824 2149 4904
rect 2265 4824 2269 4864
rect 2370 4824 2374 4864
rect 2392 4824 2396 4904
rect 2400 4824 2404 4904
rect 2505 4824 2509 4864
rect 2525 4824 2529 4864
rect 2545 4824 2549 4864
rect 2645 4824 2649 4864
rect 2765 4824 2769 4864
rect 2785 4824 2789 4864
rect 2871 4824 2875 4864
rect 2971 4824 2975 4864
rect 2991 4824 2995 4864
rect 3011 4824 3015 4864
rect 3130 4824 3134 4864
rect 3152 4824 3156 4904
rect 3160 4824 3164 4904
rect 3270 4824 3274 4864
rect 3292 4824 3296 4904
rect 3300 4824 3304 4904
rect 3405 4824 3409 4904
rect 3425 4824 3429 4904
rect 3445 4824 3449 4904
rect 3531 4824 3535 4904
rect 3541 4824 3545 4904
rect 3561 4824 3565 4904
rect 3697 4824 3701 4904
rect 3705 4824 3709 4904
rect 3805 4824 3809 4864
rect 3825 4824 3829 4864
rect 3845 4824 3849 4864
rect 3945 4824 3949 4864
rect 4031 4824 4035 4864
rect 4051 4824 4055 4864
rect 4071 4824 4075 4864
rect 4171 4824 4175 4864
rect 4191 4824 4195 4864
rect 4211 4824 4215 4864
rect 4321 4824 4325 4904
rect 4343 4824 4347 4864
rect 4365 4824 4369 4864
rect 4471 4824 4475 4904
rect 4481 4824 4485 4904
rect 4501 4824 4505 4904
rect 4611 4824 4615 4904
rect 4619 4824 4623 4904
rect 4750 4824 4754 4864
rect 4772 4824 4776 4904
rect 4780 4824 4784 4904
rect 4831 4824 4835 4904
rect 4853 4824 4857 4844
rect 4861 4824 4865 4844
rect 4881 4824 4885 4864
rect 4889 4824 4893 4864
rect 4935 4824 4939 4864
rect 4955 4824 4959 4864
rect 4967 4824 4971 4864
rect 4987 4824 4991 4864
rect 5001 4824 5005 4864
rect 5021 4824 5025 4904
rect 5116 4824 5120 4904
rect 5124 4824 5128 4904
rect 5146 4824 5150 4864
rect 5211 4824 5215 4904
rect 5233 4824 5237 4844
rect 5241 4824 5245 4844
rect 5261 4824 5265 4864
rect 5269 4824 5273 4864
rect 5315 4824 5319 4864
rect 5335 4824 5339 4864
rect 5347 4824 5351 4864
rect 5367 4824 5371 4864
rect 5381 4824 5385 4864
rect 5401 4824 5405 4904
rect 5505 4824 5509 4864
rect 5525 4824 5529 4864
rect 5611 4824 5615 4864
rect 5631 4824 5635 4864
rect 5751 4824 5755 4864
rect 5771 4824 5775 4864
rect 85 4716 89 4796
rect 105 4716 109 4796
rect 125 4716 129 4796
rect 225 4756 229 4796
rect 245 4756 249 4796
rect 265 4756 269 4796
rect 351 4716 355 4796
rect 371 4716 375 4796
rect 391 4716 395 4796
rect 491 4756 495 4796
rect 511 4756 515 4796
rect 625 4756 629 4796
rect 645 4756 649 4796
rect 665 4756 669 4796
rect 785 4756 789 4796
rect 805 4756 809 4796
rect 825 4756 829 4796
rect 911 4756 915 4796
rect 1011 4756 1015 4796
rect 1125 4756 1129 4796
rect 1230 4756 1234 4796
rect 1252 4716 1256 4796
rect 1260 4716 1264 4796
rect 1356 4716 1360 4796
rect 1364 4716 1368 4796
rect 1386 4756 1390 4796
rect 1491 4756 1495 4796
rect 1591 4756 1595 4796
rect 1611 4756 1615 4796
rect 1631 4756 1635 4796
rect 1750 4756 1754 4796
rect 1772 4716 1776 4796
rect 1780 4716 1784 4796
rect 1885 4756 1889 4796
rect 1905 4756 1909 4796
rect 1996 4716 2000 4796
rect 2004 4716 2008 4796
rect 2026 4756 2030 4796
rect 2145 4756 2149 4796
rect 2165 4756 2169 4796
rect 2185 4756 2189 4796
rect 2283 4716 2287 4796
rect 2305 4756 2309 4796
rect 2391 4756 2395 4796
rect 2411 4756 2415 4796
rect 2511 4756 2515 4796
rect 2531 4756 2535 4796
rect 2643 4716 2647 4796
rect 2665 4756 2669 4796
rect 2751 4756 2755 4796
rect 2771 4756 2775 4796
rect 2791 4756 2795 4796
rect 2917 4716 2921 4796
rect 2925 4716 2929 4796
rect 3031 4716 3035 4796
rect 3041 4716 3045 4796
rect 3071 4716 3075 4796
rect 3081 4716 3085 4796
rect 3205 4756 3209 4796
rect 3225 4756 3229 4796
rect 3325 4756 3329 4796
rect 3345 4756 3349 4796
rect 3365 4756 3369 4796
rect 3465 4716 3469 4796
rect 3485 4716 3489 4796
rect 3505 4716 3509 4796
rect 3605 4756 3609 4796
rect 3625 4756 3629 4796
rect 3645 4756 3649 4796
rect 3745 4716 3749 4796
rect 3765 4716 3769 4796
rect 3785 4716 3789 4796
rect 3871 4756 3875 4796
rect 3891 4756 3895 4796
rect 3911 4756 3915 4796
rect 4011 4756 4015 4796
rect 4031 4756 4035 4796
rect 4051 4756 4055 4796
rect 4151 4756 4155 4796
rect 4261 4716 4265 4796
rect 4283 4756 4287 4796
rect 4305 4756 4309 4796
rect 4425 4756 4429 4796
rect 4445 4756 4449 4796
rect 4465 4756 4469 4796
rect 4551 4756 4555 4796
rect 4571 4756 4575 4796
rect 4591 4756 4595 4796
rect 4691 4756 4695 4796
rect 4751 4716 4755 4796
rect 4773 4776 4777 4796
rect 4781 4776 4785 4796
rect 4801 4756 4805 4796
rect 4809 4756 4813 4796
rect 4855 4756 4859 4796
rect 4875 4756 4879 4796
rect 4887 4756 4891 4796
rect 4907 4756 4911 4796
rect 4921 4756 4925 4796
rect 4941 4716 4945 4796
rect 5036 4716 5040 4796
rect 5044 4716 5048 4796
rect 5066 4756 5070 4796
rect 5171 4756 5175 4796
rect 5191 4756 5195 4796
rect 5291 4756 5295 4796
rect 5311 4756 5315 4796
rect 5431 4756 5435 4796
rect 5451 4756 5455 4796
rect 5551 4756 5555 4796
rect 5571 4756 5575 4796
rect 5685 4756 5689 4796
rect 5705 4756 5709 4796
rect 5725 4756 5729 4796
rect 90 4344 94 4384
rect 112 4344 116 4424
rect 120 4344 124 4424
rect 225 4344 229 4384
rect 245 4344 249 4384
rect 265 4344 269 4384
rect 351 4344 355 4424
rect 371 4344 375 4424
rect 391 4344 395 4424
rect 530 4344 534 4384
rect 552 4344 556 4424
rect 560 4344 564 4424
rect 670 4344 674 4384
rect 692 4344 696 4424
rect 700 4344 704 4424
rect 791 4344 795 4384
rect 891 4344 895 4424
rect 911 4344 915 4424
rect 931 4344 935 4424
rect 1045 4344 1049 4384
rect 1145 4344 1149 4384
rect 1165 4344 1169 4384
rect 1185 4344 1189 4384
rect 1285 4344 1289 4424
rect 1305 4344 1309 4424
rect 1325 4344 1329 4424
rect 1425 4344 1429 4384
rect 1516 4344 1520 4424
rect 1524 4344 1528 4424
rect 1546 4344 1550 4384
rect 1665 4344 1669 4384
rect 1685 4344 1689 4384
rect 1785 4344 1789 4384
rect 1805 4344 1809 4384
rect 1825 4344 1829 4384
rect 1937 4344 1941 4424
rect 1945 4344 1949 4424
rect 2045 4344 2049 4384
rect 2065 4344 2069 4384
rect 2085 4344 2089 4384
rect 2205 4344 2209 4384
rect 2225 4344 2229 4384
rect 2245 4344 2249 4384
rect 2345 4344 2349 4384
rect 2365 4344 2369 4384
rect 2465 4344 2469 4384
rect 2485 4344 2489 4384
rect 2505 4344 2509 4384
rect 2591 4344 2595 4384
rect 2611 4344 2615 4384
rect 2631 4344 2635 4384
rect 2745 4344 2749 4384
rect 2857 4344 2861 4424
rect 2865 4344 2869 4424
rect 2965 4344 2969 4384
rect 2985 4344 2989 4384
rect 3005 4344 3009 4384
rect 3105 4344 3109 4384
rect 3125 4344 3129 4384
rect 3145 4344 3149 4384
rect 3231 4344 3235 4384
rect 3336 4344 3340 4424
rect 3344 4344 3348 4424
rect 3366 4344 3370 4384
rect 3481 4344 3485 4424
rect 3503 4344 3507 4384
rect 3525 4344 3529 4384
rect 3631 4344 3635 4384
rect 3651 4344 3655 4384
rect 3775 4344 3779 4424
rect 3795 4344 3799 4424
rect 3805 4344 3809 4424
rect 3891 4344 3895 4384
rect 3911 4344 3915 4384
rect 4023 4344 4027 4424
rect 4045 4344 4049 4384
rect 4131 4344 4135 4384
rect 4153 4344 4157 4384
rect 4175 4344 4179 4424
rect 4285 4344 4289 4384
rect 4305 4344 4309 4384
rect 4410 4344 4414 4384
rect 4432 4344 4436 4424
rect 4440 4344 4444 4424
rect 4531 4344 4535 4384
rect 4551 4344 4555 4384
rect 4665 4344 4669 4384
rect 4685 4344 4689 4384
rect 4771 4344 4775 4384
rect 4871 4344 4875 4384
rect 4891 4344 4895 4384
rect 4996 4344 5000 4424
rect 5004 4344 5008 4424
rect 5026 4344 5030 4384
rect 5091 4344 5095 4424
rect 5113 4344 5117 4364
rect 5121 4344 5125 4364
rect 5141 4344 5145 4384
rect 5149 4344 5153 4384
rect 5195 4344 5199 4384
rect 5215 4344 5219 4384
rect 5227 4344 5231 4384
rect 5247 4344 5251 4384
rect 5261 4344 5265 4384
rect 5281 4344 5285 4424
rect 5376 4344 5380 4424
rect 5384 4344 5388 4424
rect 5406 4344 5410 4384
rect 5511 4344 5515 4424
rect 5521 4344 5525 4424
rect 5541 4344 5545 4424
rect 5670 4344 5674 4384
rect 5692 4344 5696 4424
rect 5700 4344 5704 4424
rect 110 4276 114 4316
rect 132 4236 136 4316
rect 140 4236 144 4316
rect 250 4276 254 4316
rect 272 4236 276 4316
rect 280 4236 284 4316
rect 405 4276 409 4316
rect 425 4276 429 4316
rect 445 4276 449 4316
rect 545 4276 549 4316
rect 565 4276 569 4316
rect 585 4276 589 4316
rect 695 4236 699 4316
rect 715 4236 719 4316
rect 725 4236 729 4316
rect 830 4276 834 4316
rect 852 4236 856 4316
rect 860 4236 864 4316
rect 951 4276 955 4316
rect 1065 4236 1069 4316
rect 1085 4236 1089 4316
rect 1105 4236 1109 4316
rect 1225 4276 1229 4316
rect 1245 4276 1249 4316
rect 1265 4276 1269 4316
rect 1365 4276 1369 4316
rect 1385 4276 1389 4316
rect 1485 4276 1489 4316
rect 1505 4276 1509 4316
rect 1617 4236 1621 4316
rect 1625 4236 1629 4316
rect 1725 4276 1729 4316
rect 1745 4276 1749 4316
rect 1765 4276 1769 4316
rect 1865 4276 1869 4316
rect 1885 4276 1889 4316
rect 1905 4276 1909 4316
rect 1991 4276 1995 4316
rect 2011 4276 2015 4316
rect 2031 4276 2035 4316
rect 2131 4276 2135 4316
rect 2151 4276 2155 4316
rect 2171 4276 2175 4316
rect 2297 4236 2301 4316
rect 2305 4236 2309 4316
rect 2430 4276 2434 4316
rect 2452 4236 2456 4316
rect 2460 4236 2464 4316
rect 2585 4276 2589 4316
rect 2605 4276 2609 4316
rect 2625 4276 2629 4316
rect 2711 4276 2715 4316
rect 2831 4276 2835 4316
rect 2851 4276 2855 4316
rect 2871 4276 2875 4316
rect 2971 4276 2975 4316
rect 2991 4276 2995 4316
rect 3091 4236 3095 4316
rect 3111 4236 3115 4316
rect 3131 4236 3135 4316
rect 3231 4236 3235 4316
rect 3251 4236 3255 4316
rect 3271 4236 3275 4316
rect 3376 4236 3380 4316
rect 3384 4236 3388 4316
rect 3406 4276 3410 4316
rect 3531 4276 3535 4316
rect 3631 4276 3635 4316
rect 3651 4276 3655 4316
rect 3671 4276 3675 4316
rect 3771 4276 3775 4316
rect 3791 4276 3795 4316
rect 3811 4276 3815 4316
rect 3925 4276 3929 4316
rect 3945 4276 3949 4316
rect 4065 4276 4069 4316
rect 4085 4276 4089 4316
rect 4185 4276 4189 4316
rect 4205 4276 4209 4316
rect 4310 4276 4314 4316
rect 4332 4236 4336 4316
rect 4340 4236 4344 4316
rect 4431 4236 4435 4316
rect 4441 4236 4445 4316
rect 4461 4236 4465 4316
rect 4590 4276 4594 4316
rect 4612 4236 4616 4316
rect 4620 4236 4624 4316
rect 4736 4236 4740 4316
rect 4744 4236 4748 4316
rect 4766 4276 4770 4316
rect 4871 4236 4875 4316
rect 4879 4236 4883 4316
rect 4991 4276 4995 4316
rect 5111 4236 5115 4316
rect 5131 4236 5135 4316
rect 5151 4236 5155 4316
rect 5256 4236 5260 4316
rect 5264 4236 5268 4316
rect 5286 4276 5290 4316
rect 5391 4276 5395 4316
rect 5496 4236 5500 4316
rect 5504 4236 5508 4316
rect 5526 4276 5530 4316
rect 5595 4236 5599 4316
rect 5615 4276 5619 4316
rect 5629 4276 5633 4316
rect 5649 4276 5653 4316
rect 5661 4276 5665 4316
rect 5681 4276 5685 4316
rect 5727 4276 5731 4316
rect 5735 4276 5739 4316
rect 5755 4296 5759 4316
rect 5763 4296 5767 4316
rect 5785 4236 5789 4316
rect 85 3864 89 3904
rect 196 3864 200 3944
rect 204 3864 208 3944
rect 226 3864 230 3904
rect 345 3864 349 3904
rect 451 3864 455 3944
rect 471 3864 475 3944
rect 491 3864 495 3944
rect 617 3864 621 3944
rect 625 3864 629 3944
rect 745 3864 749 3904
rect 836 3864 840 3944
rect 844 3864 848 3944
rect 866 3864 870 3904
rect 971 3864 975 3904
rect 1071 3864 1075 3904
rect 1091 3864 1095 3904
rect 1111 3864 1115 3904
rect 1211 3864 1215 3944
rect 1231 3864 1235 3944
rect 1251 3864 1255 3944
rect 1271 3864 1275 3944
rect 1391 3864 1395 3904
rect 1411 3864 1415 3904
rect 1525 3864 1529 3904
rect 1637 3864 1641 3944
rect 1645 3864 1649 3944
rect 1745 3864 1749 3904
rect 1831 3864 1835 3904
rect 1851 3864 1855 3904
rect 1871 3864 1875 3904
rect 1990 3864 1994 3904
rect 2012 3864 2016 3944
rect 2020 3864 2024 3944
rect 2145 3864 2149 3904
rect 2165 3864 2169 3904
rect 2185 3864 2189 3904
rect 2271 3864 2275 3904
rect 2291 3864 2295 3904
rect 2311 3864 2315 3904
rect 2430 3864 2434 3904
rect 2452 3864 2456 3944
rect 2460 3864 2464 3944
rect 2565 3864 2569 3904
rect 2585 3864 2589 3904
rect 2671 3864 2675 3904
rect 2691 3864 2695 3904
rect 2791 3864 2795 3904
rect 2811 3864 2815 3904
rect 2831 3864 2835 3904
rect 2931 3864 2935 3904
rect 2951 3864 2955 3904
rect 2971 3864 2975 3904
rect 3085 3864 3089 3904
rect 3185 3864 3189 3904
rect 3205 3864 3209 3904
rect 3225 3864 3229 3904
rect 3325 3864 3329 3904
rect 3430 3864 3434 3904
rect 3452 3864 3456 3944
rect 3460 3864 3464 3944
rect 3551 3864 3555 3904
rect 3571 3864 3575 3904
rect 3695 3864 3699 3944
rect 3715 3864 3719 3944
rect 3725 3864 3729 3944
rect 3831 3864 3835 3904
rect 3851 3864 3855 3904
rect 3970 3864 3974 3904
rect 3992 3864 3996 3944
rect 4000 3864 4004 3944
rect 4105 3864 4109 3944
rect 4125 3864 4129 3944
rect 4145 3864 4149 3944
rect 4231 3864 4235 3904
rect 4251 3864 4255 3904
rect 4356 3864 4360 3944
rect 4364 3864 4368 3944
rect 4386 3864 4390 3904
rect 4496 3864 4500 3944
rect 4504 3864 4508 3944
rect 4526 3864 4530 3904
rect 4631 3864 4635 3944
rect 4641 3864 4645 3944
rect 4661 3864 4665 3944
rect 4785 3864 4789 3904
rect 4805 3864 4809 3904
rect 4891 3864 4895 3904
rect 4911 3864 4915 3904
rect 4931 3864 4935 3904
rect 5031 3864 5035 3904
rect 5145 3864 5149 3904
rect 5191 3864 5195 3944
rect 5213 3864 5217 3884
rect 5221 3864 5225 3884
rect 5241 3864 5245 3904
rect 5249 3864 5253 3904
rect 5295 3864 5299 3904
rect 5315 3864 5319 3904
rect 5327 3864 5331 3904
rect 5347 3864 5351 3904
rect 5361 3864 5365 3904
rect 5381 3864 5385 3944
rect 5431 3864 5435 3944
rect 5453 3864 5457 3884
rect 5461 3864 5465 3884
rect 5481 3864 5485 3904
rect 5489 3864 5493 3904
rect 5535 3864 5539 3904
rect 5555 3864 5559 3904
rect 5567 3864 5571 3904
rect 5587 3864 5591 3904
rect 5601 3864 5605 3904
rect 5621 3864 5625 3944
rect 5716 3864 5720 3944
rect 5724 3864 5728 3944
rect 5746 3864 5750 3904
rect 85 3796 89 3836
rect 105 3796 109 3836
rect 205 3796 209 3836
rect 225 3796 229 3836
rect 245 3796 249 3836
rect 341 3768 345 3828
rect 361 3768 365 3828
rect 405 3776 409 3836
rect 425 3776 429 3836
rect 445 3776 449 3836
rect 465 3776 469 3836
rect 570 3796 574 3836
rect 592 3756 596 3836
rect 600 3756 604 3836
rect 705 3796 709 3836
rect 725 3796 729 3836
rect 816 3756 820 3836
rect 824 3756 828 3836
rect 846 3796 850 3836
rect 985 3756 989 3836
rect 1005 3756 1009 3836
rect 1025 3756 1029 3836
rect 1045 3756 1049 3836
rect 1131 3796 1135 3836
rect 1151 3796 1155 3836
rect 1251 3796 1255 3836
rect 1271 3796 1275 3836
rect 1291 3796 1295 3836
rect 1391 3756 1395 3836
rect 1411 3756 1415 3836
rect 1431 3756 1435 3836
rect 1536 3756 1540 3836
rect 1544 3756 1548 3836
rect 1566 3796 1570 3836
rect 1671 3796 1675 3836
rect 1785 3796 1789 3836
rect 1805 3796 1809 3836
rect 1891 3796 1895 3836
rect 1911 3796 1915 3836
rect 2011 3756 2015 3836
rect 2021 3756 2025 3836
rect 2041 3756 2045 3836
rect 2151 3796 2155 3836
rect 2171 3796 2175 3836
rect 2271 3796 2275 3836
rect 2291 3796 2295 3836
rect 2311 3796 2315 3836
rect 2430 3796 2434 3836
rect 2452 3756 2456 3836
rect 2460 3756 2464 3836
rect 2551 3796 2555 3836
rect 2571 3796 2575 3836
rect 2676 3756 2680 3836
rect 2684 3756 2688 3836
rect 2706 3796 2710 3836
rect 2825 3796 2829 3836
rect 2930 3796 2934 3836
rect 2952 3756 2956 3836
rect 2960 3756 2964 3836
rect 3051 3796 3055 3836
rect 3071 3796 3075 3836
rect 3205 3796 3209 3836
rect 3225 3796 3229 3836
rect 3325 3796 3329 3836
rect 3411 3796 3415 3836
rect 3431 3796 3435 3836
rect 3451 3796 3455 3836
rect 3551 3796 3555 3836
rect 3677 3756 3681 3836
rect 3685 3756 3689 3836
rect 3791 3796 3795 3836
rect 3811 3796 3815 3836
rect 3911 3796 3915 3836
rect 4025 3796 4029 3836
rect 4071 3756 4075 3836
rect 4093 3816 4097 3836
rect 4101 3816 4105 3836
rect 4121 3796 4125 3836
rect 4129 3796 4133 3836
rect 4175 3796 4179 3836
rect 4195 3796 4199 3836
rect 4207 3796 4211 3836
rect 4227 3796 4231 3836
rect 4241 3796 4245 3836
rect 4261 3756 4265 3836
rect 4375 3756 4379 3836
rect 4385 3756 4389 3836
rect 4415 3756 4419 3836
rect 4425 3756 4429 3836
rect 4511 3796 4515 3836
rect 4531 3796 4535 3836
rect 4631 3756 4635 3836
rect 4639 3756 4643 3836
rect 4756 3756 4760 3836
rect 4764 3756 4768 3836
rect 4786 3796 4790 3836
rect 4891 3756 4895 3836
rect 5025 3796 5029 3836
rect 5045 3796 5049 3836
rect 5131 3796 5135 3836
rect 5245 3756 5249 3836
rect 5265 3756 5269 3836
rect 5285 3756 5289 3836
rect 5305 3756 5309 3836
rect 5325 3756 5329 3836
rect 5345 3756 5349 3836
rect 5365 3756 5369 3836
rect 5385 3756 5389 3836
rect 5431 3756 5435 3836
rect 5453 3816 5457 3836
rect 5461 3816 5465 3836
rect 5481 3796 5485 3836
rect 5489 3796 5493 3836
rect 5535 3796 5539 3836
rect 5555 3796 5559 3836
rect 5567 3796 5571 3836
rect 5587 3796 5591 3836
rect 5601 3796 5605 3836
rect 5621 3756 5625 3836
rect 5725 3796 5729 3836
rect 5745 3796 5749 3836
rect 90 3384 94 3424
rect 112 3384 116 3464
rect 120 3384 124 3464
rect 211 3384 215 3464
rect 231 3384 235 3464
rect 251 3384 255 3464
rect 351 3384 355 3424
rect 456 3384 460 3464
rect 464 3384 468 3464
rect 486 3384 490 3424
rect 591 3384 595 3424
rect 611 3384 615 3424
rect 631 3384 635 3424
rect 765 3384 769 3424
rect 785 3384 789 3424
rect 885 3384 889 3424
rect 905 3384 909 3424
rect 996 3384 1000 3464
rect 1004 3384 1008 3464
rect 1026 3384 1030 3424
rect 1145 3384 1149 3424
rect 1165 3384 1169 3424
rect 1185 3384 1189 3424
rect 1271 3384 1275 3424
rect 1291 3384 1295 3424
rect 1405 3384 1409 3424
rect 1425 3384 1429 3424
rect 1445 3384 1449 3424
rect 1536 3384 1540 3464
rect 1544 3384 1548 3464
rect 1566 3384 1570 3424
rect 1685 3384 1689 3464
rect 1705 3384 1709 3464
rect 1725 3384 1729 3464
rect 1825 3384 1829 3424
rect 1845 3384 1849 3424
rect 1865 3384 1869 3424
rect 1951 3384 1955 3464
rect 1971 3384 1975 3464
rect 1991 3384 1995 3464
rect 2110 3384 2114 3424
rect 2132 3384 2136 3464
rect 2140 3384 2144 3464
rect 2256 3384 2260 3464
rect 2264 3384 2268 3464
rect 2286 3384 2290 3424
rect 2405 3384 2409 3464
rect 2425 3384 2429 3464
rect 2445 3384 2449 3464
rect 2541 3384 2545 3464
rect 2563 3384 2567 3424
rect 2585 3384 2589 3424
rect 2671 3384 2675 3424
rect 2691 3384 2695 3424
rect 2810 3384 2814 3424
rect 2832 3384 2836 3464
rect 2840 3384 2844 3464
rect 2963 3384 2967 3464
rect 2985 3384 2989 3424
rect 3085 3384 3089 3424
rect 3105 3384 3109 3424
rect 3191 3384 3195 3424
rect 3211 3384 3215 3424
rect 3231 3384 3235 3424
rect 3345 3384 3349 3424
rect 3365 3384 3369 3424
rect 3385 3384 3389 3424
rect 3490 3384 3494 3424
rect 3512 3384 3516 3464
rect 3520 3384 3524 3464
rect 3630 3384 3634 3424
rect 3652 3384 3656 3464
rect 3660 3384 3664 3464
rect 3761 3384 3765 3464
rect 3783 3384 3787 3424
rect 3805 3384 3809 3424
rect 3891 3384 3895 3464
rect 3899 3384 3903 3464
rect 4050 3384 4054 3424
rect 4072 3384 4076 3464
rect 4080 3384 4084 3464
rect 4171 3384 4175 3424
rect 4276 3384 4280 3464
rect 4284 3384 4288 3464
rect 4306 3384 4310 3424
rect 4425 3384 4429 3424
rect 4445 3384 4449 3424
rect 4531 3384 4535 3424
rect 4551 3384 4555 3424
rect 4611 3384 4615 3464
rect 4633 3384 4637 3404
rect 4641 3384 4645 3404
rect 4661 3384 4665 3424
rect 4669 3384 4673 3424
rect 4715 3384 4719 3424
rect 4735 3384 4739 3424
rect 4747 3384 4751 3424
rect 4767 3384 4771 3424
rect 4781 3384 4785 3424
rect 4801 3384 4805 3464
rect 4905 3384 4909 3424
rect 4925 3384 4929 3424
rect 5030 3384 5034 3424
rect 5052 3384 5056 3464
rect 5060 3384 5064 3464
rect 5171 3384 5175 3424
rect 5191 3384 5195 3424
rect 5255 3384 5259 3464
rect 5275 3384 5279 3424
rect 5289 3384 5293 3424
rect 5309 3384 5313 3424
rect 5321 3384 5325 3424
rect 5341 3384 5345 3424
rect 5387 3384 5391 3424
rect 5395 3384 5399 3424
rect 5415 3384 5419 3404
rect 5423 3384 5427 3404
rect 5445 3384 5449 3464
rect 5545 3384 5549 3424
rect 5565 3384 5569 3424
rect 5656 3384 5660 3464
rect 5664 3384 5668 3464
rect 5686 3384 5690 3424
rect 85 3316 89 3356
rect 190 3316 194 3356
rect 212 3276 216 3356
rect 220 3276 224 3356
rect 325 3316 329 3356
rect 411 3316 415 3356
rect 431 3316 435 3356
rect 531 3276 535 3356
rect 551 3276 555 3356
rect 571 3276 575 3356
rect 671 3316 675 3356
rect 693 3316 697 3356
rect 715 3276 719 3356
rect 845 3316 849 3356
rect 865 3316 869 3356
rect 965 3316 969 3356
rect 985 3316 989 3356
rect 1005 3316 1009 3356
rect 1105 3316 1109 3356
rect 1125 3316 1129 3356
rect 1145 3316 1149 3356
rect 1231 3276 1235 3356
rect 1251 3276 1255 3356
rect 1271 3276 1275 3356
rect 1385 3316 1389 3356
rect 1485 3316 1489 3356
rect 1505 3316 1509 3356
rect 1525 3316 1529 3356
rect 1625 3316 1629 3356
rect 1645 3316 1649 3356
rect 1665 3316 1669 3356
rect 1765 3276 1769 3356
rect 1785 3276 1789 3356
rect 1805 3276 1809 3356
rect 1925 3316 1929 3356
rect 1945 3316 1949 3356
rect 2045 3276 2049 3356
rect 2065 3276 2069 3356
rect 2085 3276 2089 3356
rect 2171 3316 2175 3356
rect 2191 3316 2195 3356
rect 2301 3276 2305 3356
rect 2323 3316 2327 3356
rect 2345 3316 2349 3356
rect 2431 3316 2435 3356
rect 2451 3316 2455 3356
rect 2570 3316 2574 3356
rect 2592 3276 2596 3356
rect 2600 3276 2604 3356
rect 2705 3276 2709 3356
rect 2725 3276 2729 3356
rect 2745 3276 2749 3356
rect 2831 3316 2835 3356
rect 2851 3316 2855 3356
rect 2871 3316 2875 3356
rect 2971 3316 2975 3356
rect 2991 3316 2995 3356
rect 3011 3316 3015 3356
rect 3125 3316 3129 3356
rect 3145 3316 3149 3356
rect 3265 3316 3269 3356
rect 3285 3316 3289 3356
rect 3371 3316 3375 3356
rect 3485 3316 3489 3356
rect 3505 3316 3509 3356
rect 3525 3316 3529 3356
rect 3611 3276 3615 3356
rect 3631 3276 3635 3356
rect 3651 3276 3655 3356
rect 3770 3316 3774 3356
rect 3792 3276 3796 3356
rect 3800 3276 3804 3356
rect 3891 3316 3895 3356
rect 3951 3276 3955 3356
rect 3973 3336 3977 3356
rect 3981 3336 3985 3356
rect 4001 3316 4005 3356
rect 4009 3316 4013 3356
rect 4055 3316 4059 3356
rect 4075 3316 4079 3356
rect 4087 3316 4091 3356
rect 4107 3316 4111 3356
rect 4121 3316 4125 3356
rect 4141 3276 4145 3356
rect 4236 3276 4240 3356
rect 4244 3276 4248 3356
rect 4266 3316 4270 3356
rect 4376 3276 4380 3356
rect 4384 3276 4388 3356
rect 4406 3316 4410 3356
rect 4471 3276 4475 3356
rect 4493 3336 4497 3356
rect 4501 3336 4505 3356
rect 4521 3316 4525 3356
rect 4529 3316 4533 3356
rect 4575 3316 4579 3356
rect 4595 3316 4599 3356
rect 4607 3316 4611 3356
rect 4627 3316 4631 3356
rect 4641 3316 4645 3356
rect 4661 3276 4665 3356
rect 4756 3276 4760 3356
rect 4764 3276 4768 3356
rect 4786 3316 4790 3356
rect 4905 3316 4909 3356
rect 4925 3316 4929 3356
rect 5030 3316 5034 3356
rect 5052 3276 5056 3356
rect 5060 3276 5064 3356
rect 5165 3316 5169 3356
rect 5265 3316 5269 3356
rect 5285 3316 5289 3356
rect 5371 3316 5375 3356
rect 5496 3276 5500 3356
rect 5504 3276 5508 3356
rect 5526 3316 5530 3356
rect 5665 3316 5669 3356
rect 5685 3316 5689 3356
rect 101 2904 105 2984
rect 123 2904 127 2944
rect 145 2904 149 2944
rect 251 2904 255 2944
rect 271 2904 275 2944
rect 291 2904 295 2944
rect 391 2904 395 2944
rect 411 2904 415 2944
rect 530 2904 534 2944
rect 552 2904 556 2984
rect 560 2904 564 2984
rect 656 2904 660 2984
rect 664 2904 668 2984
rect 686 2904 690 2944
rect 796 2904 800 2984
rect 804 2904 808 2984
rect 826 2904 830 2944
rect 936 2904 940 2984
rect 944 2904 948 2984
rect 966 2904 970 2944
rect 1085 2904 1089 2944
rect 1105 2904 1109 2944
rect 1237 2904 1241 2984
rect 1245 2904 1249 2984
rect 1336 2904 1340 2984
rect 1344 2904 1348 2984
rect 1366 2904 1370 2944
rect 1485 2904 1489 2944
rect 1505 2904 1509 2944
rect 1525 2904 1529 2944
rect 1645 2904 1649 2984
rect 1665 2904 1669 2984
rect 1685 2904 1689 2984
rect 1790 2904 1794 2944
rect 1812 2904 1816 2984
rect 1820 2904 1824 2984
rect 1916 2904 1920 2984
rect 1924 2904 1928 2984
rect 1946 2904 1950 2944
rect 2090 2904 2094 2944
rect 2112 2904 2116 2984
rect 2120 2904 2124 2984
rect 2230 2904 2234 2944
rect 2252 2904 2256 2984
rect 2260 2904 2264 2984
rect 2385 2904 2389 2984
rect 2405 2904 2409 2984
rect 2425 2904 2429 2984
rect 2525 2904 2529 2984
rect 2545 2904 2549 2984
rect 2565 2904 2569 2984
rect 2665 2904 2669 2984
rect 2685 2904 2689 2984
rect 2705 2904 2709 2984
rect 2725 2904 2729 2984
rect 2835 2904 2839 2984
rect 2855 2904 2859 2984
rect 2865 2904 2869 2984
rect 2951 2904 2955 2984
rect 2959 2904 2963 2984
rect 3091 2904 3095 2944
rect 3111 2904 3115 2944
rect 3221 2904 3225 2984
rect 3243 2904 3247 2944
rect 3265 2904 3269 2944
rect 3351 2904 3355 2984
rect 3361 2904 3365 2984
rect 3381 2904 3385 2984
rect 3510 2904 3514 2944
rect 3532 2904 3536 2984
rect 3540 2904 3544 2984
rect 3650 2904 3654 2944
rect 3672 2904 3676 2984
rect 3680 2904 3684 2984
rect 3795 2904 3799 2984
rect 3815 2904 3819 2984
rect 3825 2904 3829 2984
rect 3941 2904 3945 2984
rect 3963 2904 3967 2944
rect 3985 2904 3989 2944
rect 4071 2904 4075 2984
rect 4079 2904 4083 2984
rect 4191 2904 4195 2944
rect 4211 2904 4215 2944
rect 4231 2904 4235 2944
rect 4295 2904 4299 2984
rect 4315 2904 4319 2944
rect 4329 2904 4333 2944
rect 4349 2904 4353 2944
rect 4361 2904 4365 2944
rect 4381 2904 4385 2944
rect 4427 2904 4431 2944
rect 4435 2904 4439 2944
rect 4455 2904 4459 2924
rect 4463 2904 4467 2924
rect 4485 2904 4489 2984
rect 4596 2904 4600 2984
rect 4604 2904 4608 2984
rect 4626 2904 4630 2944
rect 4736 2904 4740 2984
rect 4744 2904 4748 2984
rect 4766 2904 4770 2944
rect 4885 2904 4889 2944
rect 4905 2904 4909 2944
rect 4991 2904 4995 2944
rect 5011 2904 5015 2944
rect 5075 2904 5079 2984
rect 5095 2904 5099 2944
rect 5109 2904 5113 2944
rect 5129 2904 5133 2944
rect 5141 2904 5145 2944
rect 5161 2904 5165 2944
rect 5207 2904 5211 2944
rect 5215 2904 5219 2944
rect 5235 2904 5239 2924
rect 5243 2904 5247 2924
rect 5265 2904 5269 2984
rect 5365 2904 5369 2984
rect 5385 2904 5389 2984
rect 5405 2904 5409 2984
rect 5425 2904 5429 2984
rect 5445 2904 5449 2984
rect 5465 2904 5469 2984
rect 5485 2904 5489 2984
rect 5505 2904 5509 2984
rect 5551 2904 5555 2984
rect 5573 2904 5577 2924
rect 5581 2904 5585 2924
rect 5601 2904 5605 2944
rect 5609 2904 5613 2944
rect 5655 2904 5659 2944
rect 5675 2904 5679 2944
rect 5687 2904 5691 2944
rect 5707 2904 5711 2944
rect 5721 2904 5725 2944
rect 5741 2904 5745 2984
rect 85 2836 89 2876
rect 105 2836 109 2876
rect 196 2796 200 2876
rect 204 2796 208 2876
rect 226 2836 230 2876
rect 345 2836 349 2876
rect 431 2796 435 2876
rect 451 2796 455 2876
rect 471 2796 475 2876
rect 585 2836 589 2876
rect 605 2836 609 2876
rect 691 2836 695 2876
rect 713 2836 717 2876
rect 735 2796 739 2876
rect 831 2836 835 2876
rect 851 2836 855 2876
rect 951 2796 955 2876
rect 971 2796 975 2876
rect 991 2796 995 2876
rect 1091 2836 1095 2876
rect 1111 2836 1115 2876
rect 1250 2836 1254 2876
rect 1272 2796 1276 2876
rect 1280 2796 1284 2876
rect 1376 2796 1380 2876
rect 1384 2796 1388 2876
rect 1406 2836 1410 2876
rect 1535 2796 1539 2876
rect 1555 2796 1559 2876
rect 1565 2796 1569 2876
rect 1651 2796 1655 2876
rect 1659 2796 1663 2876
rect 1781 2796 1785 2876
rect 1803 2836 1807 2876
rect 1825 2836 1829 2876
rect 1945 2836 1949 2876
rect 1965 2836 1969 2876
rect 2056 2796 2060 2876
rect 2064 2796 2068 2876
rect 2086 2836 2090 2876
rect 2201 2796 2205 2876
rect 2223 2836 2227 2876
rect 2245 2836 2249 2876
rect 2345 2836 2349 2876
rect 2365 2836 2369 2876
rect 2471 2796 2475 2876
rect 2479 2796 2483 2876
rect 2605 2836 2609 2876
rect 2625 2836 2629 2876
rect 2645 2836 2649 2876
rect 2741 2796 2745 2876
rect 2763 2836 2767 2876
rect 2785 2836 2789 2876
rect 2896 2796 2900 2876
rect 2904 2796 2908 2876
rect 2926 2836 2930 2876
rect 3045 2836 3049 2876
rect 3065 2836 3069 2876
rect 3085 2836 3089 2876
rect 3171 2836 3175 2876
rect 3191 2836 3195 2876
rect 3310 2836 3314 2876
rect 3332 2796 3336 2876
rect 3340 2796 3344 2876
rect 3441 2796 3445 2876
rect 3463 2836 3467 2876
rect 3485 2836 3489 2876
rect 3571 2796 3575 2876
rect 3579 2796 3583 2876
rect 3691 2836 3695 2876
rect 3711 2836 3715 2876
rect 3731 2836 3735 2876
rect 3831 2836 3835 2876
rect 3851 2836 3855 2876
rect 3965 2796 3969 2876
rect 4070 2836 4074 2876
rect 4092 2796 4096 2876
rect 4100 2796 4104 2876
rect 4191 2836 4195 2876
rect 4211 2836 4215 2876
rect 4311 2796 4315 2876
rect 4411 2836 4415 2876
rect 4471 2796 4475 2876
rect 4493 2856 4497 2876
rect 4501 2856 4505 2876
rect 4521 2836 4525 2876
rect 4529 2836 4533 2876
rect 4575 2836 4579 2876
rect 4595 2836 4599 2876
rect 4607 2836 4611 2876
rect 4627 2836 4631 2876
rect 4641 2836 4645 2876
rect 4661 2796 4665 2876
rect 4715 2796 4719 2876
rect 4735 2836 4739 2876
rect 4749 2836 4753 2876
rect 4769 2836 4773 2876
rect 4781 2836 4785 2876
rect 4801 2836 4805 2876
rect 4847 2836 4851 2876
rect 4855 2836 4859 2876
rect 4875 2856 4879 2876
rect 4883 2856 4887 2876
rect 4905 2796 4909 2876
rect 5016 2796 5020 2876
rect 5024 2796 5028 2876
rect 5046 2836 5050 2876
rect 5151 2836 5155 2876
rect 5171 2836 5175 2876
rect 5271 2796 5275 2876
rect 5291 2796 5295 2876
rect 5351 2796 5355 2876
rect 5373 2856 5377 2876
rect 5381 2856 5385 2876
rect 5401 2836 5405 2876
rect 5409 2836 5413 2876
rect 5455 2836 5459 2876
rect 5475 2836 5479 2876
rect 5487 2836 5491 2876
rect 5507 2836 5511 2876
rect 5521 2836 5525 2876
rect 5541 2796 5545 2876
rect 5636 2796 5640 2876
rect 5644 2796 5648 2876
rect 5666 2836 5670 2876
rect 85 2424 89 2464
rect 171 2424 175 2464
rect 285 2424 289 2504
rect 305 2424 309 2504
rect 325 2424 329 2504
rect 411 2424 415 2464
rect 431 2424 435 2464
rect 451 2424 455 2464
rect 551 2424 555 2464
rect 651 2424 655 2504
rect 659 2424 663 2504
rect 776 2424 780 2504
rect 784 2424 788 2504
rect 806 2424 810 2464
rect 931 2424 935 2504
rect 951 2424 955 2504
rect 971 2424 975 2504
rect 1090 2424 1094 2464
rect 1112 2424 1116 2504
rect 1120 2424 1124 2504
rect 1225 2424 1229 2464
rect 1245 2424 1249 2464
rect 1331 2424 1335 2464
rect 1353 2424 1357 2464
rect 1375 2424 1379 2504
rect 1485 2424 1489 2464
rect 1505 2424 1509 2464
rect 1525 2424 1529 2464
rect 1611 2424 1615 2464
rect 1716 2424 1720 2504
rect 1724 2424 1728 2504
rect 1746 2424 1750 2464
rect 1870 2424 1874 2464
rect 1892 2424 1896 2504
rect 1900 2424 1904 2504
rect 1996 2424 2000 2504
rect 2004 2424 2008 2504
rect 2026 2424 2030 2464
rect 2145 2424 2149 2464
rect 2165 2424 2169 2464
rect 2185 2424 2189 2464
rect 2285 2424 2289 2504
rect 2305 2424 2309 2504
rect 2325 2424 2329 2504
rect 2411 2424 2415 2464
rect 2431 2424 2435 2464
rect 2570 2424 2574 2464
rect 2592 2424 2596 2504
rect 2600 2424 2604 2504
rect 2696 2424 2700 2504
rect 2704 2424 2708 2504
rect 2726 2424 2730 2464
rect 2845 2424 2849 2504
rect 2865 2424 2869 2504
rect 2885 2424 2889 2504
rect 2985 2424 2989 2464
rect 3076 2424 3080 2504
rect 3084 2424 3088 2504
rect 3106 2424 3110 2464
rect 3231 2424 3235 2464
rect 3251 2424 3255 2464
rect 3365 2424 3369 2464
rect 3385 2424 3389 2464
rect 3405 2424 3409 2464
rect 3491 2424 3495 2464
rect 3513 2424 3517 2464
rect 3535 2424 3539 2504
rect 3631 2424 3635 2464
rect 3651 2424 3655 2464
rect 3751 2424 3755 2504
rect 3771 2424 3775 2504
rect 3791 2424 3795 2504
rect 3811 2424 3815 2504
rect 3911 2424 3915 2504
rect 3919 2424 3923 2504
rect 3999 2424 4003 2464
rect 4044 2424 4048 2464
rect 4064 2424 4068 2464
rect 4084 2424 4088 2464
rect 4104 2424 4108 2464
rect 4149 2424 4153 2444
rect 4169 2424 4173 2444
rect 4214 2424 4218 2464
rect 4234 2424 4238 2464
rect 4279 2424 4283 2464
rect 4299 2424 4303 2444
rect 4319 2424 4323 2444
rect 4364 2424 4368 2464
rect 4384 2424 4388 2464
rect 4404 2424 4408 2464
rect 4424 2424 4428 2464
rect 4472 2424 4476 2464
rect 4492 2424 4496 2464
rect 4512 2424 4516 2464
rect 4532 2424 4536 2464
rect 4577 2424 4581 2444
rect 4597 2424 4601 2444
rect 4617 2424 4621 2464
rect 4662 2424 4666 2464
rect 4682 2424 4686 2464
rect 4727 2424 4731 2444
rect 4747 2424 4751 2444
rect 4792 2424 4796 2464
rect 4812 2424 4816 2464
rect 4832 2424 4836 2464
rect 4852 2424 4856 2464
rect 4897 2424 4901 2464
rect 4955 2424 4959 2504
rect 4975 2424 4979 2464
rect 4989 2424 4993 2464
rect 5009 2424 5013 2464
rect 5021 2424 5025 2464
rect 5041 2424 5045 2464
rect 5087 2424 5091 2464
rect 5095 2424 5099 2464
rect 5115 2424 5119 2444
rect 5123 2424 5127 2444
rect 5145 2424 5149 2504
rect 5245 2424 5249 2504
rect 5265 2424 5269 2504
rect 5285 2424 5289 2504
rect 5305 2424 5309 2504
rect 5325 2424 5329 2504
rect 5345 2424 5349 2504
rect 5365 2424 5369 2504
rect 5385 2424 5389 2504
rect 5491 2424 5495 2504
rect 5511 2424 5515 2504
rect 5531 2424 5535 2504
rect 5551 2424 5555 2504
rect 5571 2424 5575 2504
rect 5591 2424 5595 2504
rect 5611 2424 5615 2504
rect 5631 2424 5635 2504
rect 5731 2424 5735 2504
rect 83 2316 87 2396
rect 105 2356 109 2396
rect 205 2356 209 2396
rect 225 2356 229 2396
rect 245 2356 249 2396
rect 331 2356 335 2396
rect 351 2356 355 2396
rect 456 2316 460 2396
rect 464 2316 468 2396
rect 486 2356 490 2396
rect 610 2356 614 2396
rect 632 2316 636 2396
rect 640 2316 644 2396
rect 765 2356 769 2396
rect 785 2356 789 2396
rect 805 2356 809 2396
rect 905 2356 909 2396
rect 925 2356 929 2396
rect 1035 2316 1039 2396
rect 1055 2316 1059 2396
rect 1065 2316 1069 2396
rect 1151 2316 1155 2396
rect 1265 2356 1269 2396
rect 1285 2356 1289 2396
rect 1305 2356 1309 2396
rect 1405 2316 1409 2396
rect 1425 2316 1429 2396
rect 1445 2316 1449 2396
rect 1570 2356 1574 2396
rect 1592 2316 1596 2396
rect 1600 2316 1604 2396
rect 1705 2316 1709 2396
rect 1725 2316 1729 2396
rect 1745 2316 1749 2396
rect 1845 2356 1849 2396
rect 1865 2356 1869 2396
rect 1885 2356 1889 2396
rect 1985 2356 1989 2396
rect 2005 2356 2009 2396
rect 2025 2356 2029 2396
rect 2079 2356 2083 2396
rect 2124 2356 2128 2396
rect 2144 2356 2148 2396
rect 2164 2356 2168 2396
rect 2184 2356 2188 2396
rect 2229 2376 2233 2396
rect 2249 2376 2253 2396
rect 2294 2356 2298 2396
rect 2314 2356 2318 2396
rect 2359 2356 2363 2396
rect 2379 2376 2383 2396
rect 2399 2376 2403 2396
rect 2444 2356 2448 2396
rect 2464 2356 2468 2396
rect 2484 2356 2488 2396
rect 2504 2356 2508 2396
rect 2603 2316 2607 2396
rect 2625 2356 2629 2396
rect 2736 2316 2740 2396
rect 2744 2316 2748 2396
rect 2766 2356 2770 2396
rect 2876 2316 2880 2396
rect 2884 2316 2888 2396
rect 2906 2356 2910 2396
rect 3025 2356 3029 2396
rect 3045 2356 3049 2396
rect 3151 2356 3155 2396
rect 3171 2356 3175 2396
rect 3285 2316 3289 2396
rect 3305 2316 3309 2396
rect 3325 2316 3329 2396
rect 3411 2316 3415 2396
rect 3419 2316 3423 2396
rect 3556 2316 3560 2396
rect 3564 2316 3568 2396
rect 3586 2356 3590 2396
rect 3691 2356 3695 2396
rect 3711 2356 3715 2396
rect 3811 2356 3815 2396
rect 3833 2316 3837 2396
rect 3899 2356 3903 2396
rect 3944 2356 3948 2396
rect 3964 2356 3968 2396
rect 3984 2356 3988 2396
rect 4004 2356 4008 2396
rect 4049 2376 4053 2396
rect 4069 2376 4073 2396
rect 4114 2356 4118 2396
rect 4134 2356 4138 2396
rect 4179 2356 4183 2396
rect 4199 2376 4203 2396
rect 4219 2376 4223 2396
rect 4264 2356 4268 2396
rect 4284 2356 4288 2396
rect 4304 2356 4308 2396
rect 4324 2356 4328 2396
rect 4411 2356 4415 2396
rect 4433 2356 4437 2396
rect 4455 2316 4459 2396
rect 4551 2316 4555 2396
rect 4571 2316 4575 2396
rect 4591 2316 4595 2396
rect 4611 2316 4615 2396
rect 4711 2356 4715 2396
rect 4731 2356 4735 2396
rect 4843 2316 4847 2396
rect 4865 2356 4869 2396
rect 4951 2356 4955 2396
rect 5051 2316 5055 2396
rect 5071 2316 5075 2396
rect 5091 2316 5095 2396
rect 5111 2316 5115 2396
rect 5211 2356 5215 2396
rect 5231 2356 5235 2396
rect 5331 2316 5335 2396
rect 5431 2356 5435 2396
rect 5451 2356 5455 2396
rect 5551 2356 5555 2396
rect 5651 2348 5655 2388
rect 5671 2308 5675 2388
rect 5681 2308 5685 2388
rect 5701 2316 5705 2396
rect 5711 2316 5715 2396
rect 103 1944 107 2024
rect 125 1944 129 1984
rect 245 1944 249 1984
rect 265 1944 269 1984
rect 285 1944 289 1984
rect 371 1944 375 2024
rect 391 1944 395 2024
rect 411 1944 415 2024
rect 525 1944 529 1984
rect 630 1944 634 1984
rect 652 1944 656 2024
rect 660 1944 664 2024
rect 765 1944 769 2024
rect 785 1944 789 2024
rect 805 1944 809 2024
rect 891 1944 895 1984
rect 911 1944 915 1984
rect 931 1944 935 1984
rect 1065 1944 1069 1984
rect 1085 1944 1089 1984
rect 1105 1944 1109 1984
rect 1210 1944 1214 1984
rect 1232 1944 1236 2024
rect 1240 1944 1244 2024
rect 1350 1944 1354 1984
rect 1372 1944 1376 2024
rect 1380 1944 1384 2024
rect 1485 1944 1489 2024
rect 1505 1944 1509 2024
rect 1525 1944 1529 2024
rect 1625 1944 1629 1984
rect 1645 1944 1649 1984
rect 1665 1944 1669 1984
rect 1756 1944 1760 2024
rect 1764 1944 1768 2024
rect 1786 1944 1790 1984
rect 1891 1944 1895 2024
rect 1911 1944 1915 2024
rect 1931 1944 1935 2024
rect 2041 1952 2045 2012
rect 2061 1952 2065 2012
rect 2105 1944 2109 2004
rect 2125 1944 2129 2004
rect 2145 1944 2149 2004
rect 2165 1944 2169 2004
rect 2265 1944 2269 1984
rect 2285 1944 2289 1984
rect 2305 1944 2309 1984
rect 2359 1944 2363 1984
rect 2404 1944 2408 1984
rect 2424 1944 2428 1984
rect 2444 1944 2448 1984
rect 2464 1944 2468 1984
rect 2509 1944 2513 1964
rect 2529 1944 2533 1964
rect 2574 1944 2578 1984
rect 2594 1944 2598 1984
rect 2639 1944 2643 1984
rect 2659 1944 2663 1964
rect 2679 1944 2683 1964
rect 2724 1944 2728 1984
rect 2744 1944 2748 1984
rect 2764 1944 2768 1984
rect 2784 1944 2788 1984
rect 2876 1944 2880 2024
rect 2884 1944 2888 2024
rect 2906 1944 2910 1984
rect 3025 1944 3029 1984
rect 3045 1944 3049 1984
rect 3131 1944 3135 1984
rect 3151 1944 3155 1984
rect 3271 1944 3275 2024
rect 3279 1944 3283 2024
rect 3401 1944 3405 2024
rect 3423 1944 3427 1984
rect 3445 1944 3449 1984
rect 3531 1944 3535 2024
rect 3551 1944 3555 2024
rect 3571 1944 3575 2024
rect 3705 1944 3709 2024
rect 3811 1944 3815 1984
rect 3831 1944 3835 1984
rect 3851 1944 3855 1984
rect 3971 1944 3975 2024
rect 4101 1944 4105 2024
rect 4123 1944 4127 1984
rect 4145 1944 4149 1984
rect 4245 1944 4249 1984
rect 4265 1944 4269 1984
rect 4370 1944 4374 1984
rect 4392 1944 4396 2024
rect 4400 1944 4404 2024
rect 4496 1944 4500 2024
rect 4504 1944 4508 2024
rect 4526 1944 4530 1984
rect 4631 1944 4635 1984
rect 4651 1944 4655 1984
rect 4751 1944 4755 1984
rect 4771 1944 4775 1984
rect 4910 1944 4914 1984
rect 4932 1944 4936 2024
rect 4940 1944 4944 2024
rect 5050 1944 5054 1984
rect 5072 1944 5076 2024
rect 5080 1944 5084 2024
rect 5171 1944 5175 1984
rect 5271 1944 5275 2024
rect 5279 1944 5283 2024
rect 5391 1944 5395 1984
rect 5411 1944 5415 1984
rect 5511 1944 5515 1984
rect 5625 1944 5629 1984
rect 5716 1944 5720 2024
rect 5724 1944 5728 2024
rect 5746 1944 5750 1984
rect 85 1876 89 1916
rect 105 1876 109 1916
rect 125 1876 129 1916
rect 211 1836 215 1916
rect 231 1836 235 1916
rect 251 1836 255 1916
rect 370 1876 374 1916
rect 392 1836 396 1916
rect 400 1836 404 1916
rect 505 1876 509 1916
rect 525 1876 529 1916
rect 545 1876 549 1916
rect 677 1836 681 1916
rect 685 1836 689 1916
rect 771 1836 775 1916
rect 791 1836 795 1916
rect 811 1836 815 1916
rect 945 1876 949 1916
rect 1070 1876 1074 1916
rect 1092 1836 1096 1916
rect 1100 1836 1104 1916
rect 1210 1876 1214 1916
rect 1232 1836 1236 1916
rect 1240 1836 1244 1916
rect 1345 1876 1349 1916
rect 1450 1876 1454 1916
rect 1472 1836 1476 1916
rect 1480 1836 1484 1916
rect 1576 1836 1580 1916
rect 1584 1836 1588 1916
rect 1606 1876 1610 1916
rect 1730 1876 1734 1916
rect 1752 1836 1756 1916
rect 1760 1836 1764 1916
rect 1865 1876 1869 1916
rect 1885 1876 1889 1916
rect 1985 1876 1989 1916
rect 2005 1876 2009 1916
rect 2125 1836 2129 1916
rect 2145 1836 2149 1916
rect 2199 1876 2203 1916
rect 2244 1876 2248 1916
rect 2264 1876 2268 1916
rect 2284 1876 2288 1916
rect 2304 1876 2308 1916
rect 2349 1896 2353 1916
rect 2369 1896 2373 1916
rect 2414 1876 2418 1916
rect 2434 1876 2438 1916
rect 2479 1876 2483 1916
rect 2499 1896 2503 1916
rect 2519 1896 2523 1916
rect 2564 1876 2568 1916
rect 2584 1876 2588 1916
rect 2604 1876 2608 1916
rect 2624 1876 2628 1916
rect 2711 1876 2715 1916
rect 2731 1876 2735 1916
rect 2845 1876 2849 1916
rect 2865 1876 2869 1916
rect 2885 1876 2889 1916
rect 2990 1876 2994 1916
rect 3012 1836 3016 1916
rect 3020 1836 3024 1916
rect 3111 1836 3115 1916
rect 3119 1836 3123 1916
rect 3231 1868 3235 1908
rect 3251 1828 3255 1908
rect 3261 1828 3265 1908
rect 3281 1836 3285 1916
rect 3291 1836 3295 1916
rect 3405 1876 3409 1916
rect 3491 1836 3495 1916
rect 3501 1836 3505 1916
rect 3531 1836 3535 1916
rect 3541 1836 3545 1916
rect 3670 1876 3674 1916
rect 3692 1836 3696 1916
rect 3700 1836 3704 1916
rect 3830 1876 3834 1916
rect 3852 1836 3856 1916
rect 3860 1836 3864 1916
rect 3956 1836 3960 1916
rect 3964 1836 3968 1916
rect 3986 1876 3990 1916
rect 4105 1876 4109 1916
rect 4125 1876 4129 1916
rect 4225 1836 4229 1916
rect 4245 1836 4249 1916
rect 4265 1836 4269 1916
rect 4285 1836 4289 1916
rect 4385 1876 4389 1916
rect 4405 1876 4409 1916
rect 4496 1836 4500 1916
rect 4504 1836 4508 1916
rect 4526 1876 4530 1916
rect 4641 1836 4645 1916
rect 4663 1876 4667 1916
rect 4685 1876 4689 1916
rect 4797 1836 4801 1916
rect 4805 1836 4809 1916
rect 4905 1876 4909 1916
rect 4925 1876 4929 1916
rect 5025 1836 5029 1916
rect 5045 1836 5049 1916
rect 5065 1836 5069 1916
rect 5085 1836 5089 1916
rect 5185 1876 5189 1916
rect 5297 1836 5301 1916
rect 5305 1836 5309 1916
rect 5396 1836 5400 1916
rect 5404 1836 5408 1916
rect 5426 1876 5430 1916
rect 5550 1876 5554 1916
rect 5572 1836 5576 1916
rect 5580 1836 5584 1916
rect 5671 1836 5675 1916
rect 5691 1836 5695 1916
rect 91 1464 95 1504
rect 111 1464 115 1504
rect 131 1464 135 1504
rect 245 1464 249 1504
rect 265 1464 269 1504
rect 285 1464 289 1504
rect 371 1464 375 1544
rect 391 1464 395 1544
rect 411 1464 415 1544
rect 525 1464 529 1544
rect 545 1464 549 1544
rect 565 1464 569 1544
rect 651 1464 655 1504
rect 671 1464 675 1504
rect 771 1464 775 1504
rect 890 1464 894 1504
rect 912 1464 916 1544
rect 920 1464 924 1544
rect 1025 1464 1029 1504
rect 1045 1464 1049 1504
rect 1065 1464 1069 1504
rect 1165 1464 1169 1504
rect 1185 1464 1189 1504
rect 1291 1464 1295 1544
rect 1299 1464 1303 1544
rect 1423 1464 1427 1544
rect 1445 1464 1449 1504
rect 1565 1464 1569 1504
rect 1651 1464 1655 1544
rect 1671 1464 1675 1544
rect 1691 1464 1695 1544
rect 1711 1464 1715 1544
rect 1779 1464 1783 1504
rect 1824 1464 1828 1504
rect 1844 1464 1848 1504
rect 1864 1464 1868 1504
rect 1884 1464 1888 1504
rect 1929 1464 1933 1484
rect 1949 1464 1953 1484
rect 1994 1464 1998 1504
rect 2014 1464 2018 1504
rect 2059 1464 2063 1504
rect 2079 1464 2083 1484
rect 2099 1464 2103 1484
rect 2144 1464 2148 1504
rect 2164 1464 2168 1504
rect 2184 1464 2188 1504
rect 2204 1464 2208 1504
rect 2316 1464 2320 1544
rect 2324 1464 2328 1544
rect 2346 1464 2350 1504
rect 2451 1464 2455 1504
rect 2471 1464 2475 1504
rect 2590 1464 2594 1504
rect 2612 1464 2616 1544
rect 2620 1464 2624 1544
rect 2725 1464 2729 1504
rect 2745 1464 2749 1504
rect 2850 1464 2854 1504
rect 2872 1464 2876 1544
rect 2880 1464 2884 1544
rect 2990 1464 2994 1504
rect 3012 1464 3016 1544
rect 3020 1464 3024 1544
rect 3072 1464 3076 1504
rect 3092 1464 3096 1504
rect 3112 1464 3116 1504
rect 3132 1464 3136 1504
rect 3177 1464 3181 1484
rect 3197 1464 3201 1484
rect 3217 1464 3221 1504
rect 3262 1464 3266 1504
rect 3282 1464 3286 1504
rect 3327 1464 3331 1484
rect 3347 1464 3351 1484
rect 3392 1464 3396 1504
rect 3412 1464 3416 1504
rect 3432 1464 3436 1504
rect 3452 1464 3456 1504
rect 3497 1464 3501 1504
rect 3605 1464 3609 1544
rect 3625 1464 3629 1544
rect 3645 1464 3649 1544
rect 3736 1464 3740 1544
rect 3744 1464 3748 1544
rect 3766 1464 3770 1504
rect 3883 1464 3887 1544
rect 3905 1464 3909 1504
rect 4001 1464 4005 1544
rect 4023 1464 4027 1504
rect 4045 1464 4049 1504
rect 4131 1464 4135 1504
rect 4151 1464 4155 1504
rect 4265 1464 4269 1544
rect 4285 1464 4289 1544
rect 4305 1464 4309 1544
rect 4325 1464 4329 1544
rect 4425 1464 4429 1544
rect 4445 1464 4449 1544
rect 4465 1464 4469 1544
rect 4485 1464 4489 1544
rect 4591 1464 4595 1544
rect 4611 1464 4615 1544
rect 4631 1464 4635 1544
rect 4651 1464 4655 1544
rect 4751 1464 4755 1504
rect 4771 1464 4775 1504
rect 4876 1464 4880 1544
rect 4884 1464 4888 1544
rect 4906 1464 4910 1504
rect 5021 1464 5025 1544
rect 5043 1464 5047 1504
rect 5065 1464 5069 1504
rect 5171 1464 5175 1504
rect 5191 1464 5195 1504
rect 5211 1464 5215 1504
rect 5311 1464 5315 1544
rect 5331 1464 5335 1544
rect 5351 1464 5355 1544
rect 5371 1464 5375 1544
rect 5471 1464 5475 1504
rect 5491 1464 5495 1504
rect 5591 1464 5595 1504
rect 5611 1464 5615 1504
rect 5631 1464 5635 1504
rect 5765 1464 5769 1544
rect 85 1396 89 1436
rect 105 1396 109 1436
rect 125 1396 129 1436
rect 211 1356 215 1436
rect 231 1356 235 1436
rect 251 1356 255 1436
rect 365 1396 369 1436
rect 385 1396 389 1436
rect 405 1396 409 1436
rect 510 1396 514 1436
rect 532 1356 536 1436
rect 540 1356 544 1436
rect 650 1396 654 1436
rect 672 1356 676 1436
rect 680 1356 684 1436
rect 801 1356 805 1436
rect 823 1396 827 1436
rect 845 1396 849 1436
rect 931 1396 935 1436
rect 951 1396 955 1436
rect 1065 1396 1069 1436
rect 1151 1396 1155 1436
rect 1171 1396 1175 1436
rect 1191 1396 1195 1436
rect 1291 1396 1295 1436
rect 1311 1396 1315 1436
rect 1425 1396 1429 1436
rect 1445 1396 1449 1436
rect 1545 1396 1549 1436
rect 1565 1396 1569 1436
rect 1685 1396 1689 1436
rect 1705 1396 1709 1436
rect 1725 1396 1729 1436
rect 1811 1396 1815 1436
rect 1831 1396 1835 1436
rect 1945 1396 1949 1436
rect 1965 1396 1969 1436
rect 1985 1396 1989 1436
rect 2085 1396 2089 1436
rect 2205 1396 2209 1436
rect 2225 1396 2229 1436
rect 2245 1396 2249 1436
rect 2345 1396 2349 1436
rect 2365 1396 2369 1436
rect 2385 1396 2389 1436
rect 2471 1396 2475 1436
rect 2610 1396 2614 1436
rect 2632 1356 2636 1436
rect 2640 1356 2644 1436
rect 2731 1356 2735 1436
rect 2751 1356 2755 1436
rect 2771 1356 2775 1436
rect 2890 1396 2894 1436
rect 2912 1356 2916 1436
rect 2920 1356 2924 1436
rect 3030 1396 3034 1436
rect 3052 1356 3056 1436
rect 3060 1356 3064 1436
rect 3170 1396 3174 1436
rect 3192 1356 3196 1436
rect 3200 1356 3204 1436
rect 3305 1396 3309 1436
rect 3391 1396 3395 1436
rect 3503 1356 3507 1436
rect 3525 1396 3529 1436
rect 3645 1356 3649 1436
rect 3665 1356 3669 1436
rect 3685 1356 3689 1436
rect 3776 1356 3780 1436
rect 3784 1356 3788 1436
rect 3806 1396 3810 1436
rect 3925 1396 3929 1436
rect 4030 1396 4034 1436
rect 4052 1356 4056 1436
rect 4060 1356 4064 1436
rect 4170 1396 4174 1436
rect 4192 1356 4196 1436
rect 4200 1356 4204 1436
rect 4305 1356 4309 1436
rect 4325 1356 4329 1436
rect 4345 1356 4349 1436
rect 4450 1396 4454 1436
rect 4472 1356 4476 1436
rect 4480 1356 4484 1436
rect 4596 1356 4600 1436
rect 4604 1356 4608 1436
rect 4626 1396 4630 1436
rect 4731 1396 4735 1436
rect 4751 1396 4755 1436
rect 4856 1356 4860 1436
rect 4864 1356 4868 1436
rect 4886 1396 4890 1436
rect 4991 1356 4995 1436
rect 4999 1356 5003 1436
rect 5111 1396 5115 1436
rect 5131 1396 5135 1436
rect 5245 1396 5249 1436
rect 5265 1396 5269 1436
rect 5370 1396 5374 1436
rect 5392 1356 5396 1436
rect 5400 1356 5404 1436
rect 5496 1356 5500 1436
rect 5504 1356 5508 1436
rect 5526 1396 5530 1436
rect 5656 1356 5660 1436
rect 5664 1356 5668 1436
rect 5686 1396 5690 1436
rect 85 984 89 1024
rect 171 984 175 1064
rect 191 984 195 1064
rect 211 984 215 1064
rect 316 984 320 1064
rect 324 984 328 1064
rect 346 984 350 1024
rect 456 984 460 1064
rect 464 984 468 1064
rect 486 984 490 1024
rect 605 984 609 1024
rect 625 984 629 1024
rect 645 984 649 1024
rect 736 984 740 1064
rect 744 984 748 1064
rect 766 984 770 1024
rect 891 984 895 1064
rect 911 984 915 1064
rect 931 984 935 1064
rect 1050 984 1054 1024
rect 1072 984 1076 1064
rect 1080 984 1084 1064
rect 1185 984 1189 1024
rect 1271 984 1275 1064
rect 1291 984 1295 1064
rect 1311 984 1315 1064
rect 1425 984 1429 1024
rect 1537 984 1541 1064
rect 1545 984 1549 1064
rect 1651 984 1655 1024
rect 1765 984 1769 1024
rect 1785 984 1789 1024
rect 1805 984 1809 1024
rect 1905 984 1909 1024
rect 1925 984 1929 1024
rect 2030 984 2034 1024
rect 2052 984 2056 1064
rect 2060 984 2064 1064
rect 2165 984 2169 1024
rect 2185 984 2189 1024
rect 2205 984 2209 1024
rect 2305 984 2309 1024
rect 2325 984 2329 1024
rect 2345 984 2349 1024
rect 2450 984 2454 1024
rect 2472 984 2476 1064
rect 2480 984 2484 1064
rect 2585 984 2589 1024
rect 2605 984 2609 1024
rect 2625 984 2629 1024
rect 2731 984 2735 1024
rect 2831 984 2835 1064
rect 2839 984 2843 1064
rect 2951 984 2955 1064
rect 2959 984 2963 1064
rect 3071 984 3075 1024
rect 3093 984 3097 1024
rect 3115 984 3119 1064
rect 3237 984 3241 1064
rect 3245 984 3249 1064
rect 3377 984 3381 1064
rect 3385 984 3389 1064
rect 3485 984 3489 1024
rect 3590 984 3594 1024
rect 3612 984 3616 1064
rect 3620 984 3624 1064
rect 3730 984 3734 1024
rect 3752 984 3756 1064
rect 3760 984 3764 1064
rect 3851 984 3855 1024
rect 3871 984 3875 1024
rect 3971 984 3975 1024
rect 3991 984 3995 1024
rect 4091 984 4095 1064
rect 4099 984 4103 1064
rect 4211 984 4215 1024
rect 4325 984 4329 1064
rect 4345 984 4349 1064
rect 4365 984 4369 1064
rect 4490 984 4494 1024
rect 4512 984 4516 1064
rect 4520 984 4524 1064
rect 4625 984 4629 1064
rect 4645 984 4649 1064
rect 4665 984 4669 1064
rect 4756 984 4760 1064
rect 4764 984 4768 1064
rect 4786 984 4790 1024
rect 4891 984 4895 1024
rect 4913 984 4917 1064
rect 5011 984 5015 1024
rect 5111 984 5115 1024
rect 5225 984 5229 1024
rect 5245 984 5249 1024
rect 5370 984 5374 1024
rect 5392 984 5396 1064
rect 5400 984 5404 1064
rect 5491 984 5495 1064
rect 5499 984 5503 1064
rect 5625 984 5629 1024
rect 5645 984 5649 1024
rect 5665 984 5669 1024
rect 5765 984 5769 1024
rect 85 916 89 956
rect 105 916 109 956
rect 125 916 129 956
rect 211 876 215 956
rect 231 876 235 956
rect 251 876 255 956
rect 365 916 369 956
rect 385 916 389 956
rect 405 916 409 956
rect 505 876 509 956
rect 525 876 529 956
rect 545 876 549 956
rect 645 916 649 956
rect 665 916 669 956
rect 685 916 689 956
rect 771 876 775 956
rect 791 876 795 956
rect 811 876 815 956
rect 930 916 934 956
rect 952 876 956 956
rect 960 876 964 956
rect 1065 916 1069 956
rect 1085 916 1089 956
rect 1105 916 1109 956
rect 1196 876 1200 956
rect 1204 876 1208 956
rect 1226 916 1230 956
rect 1345 916 1349 956
rect 1365 916 1369 956
rect 1385 916 1389 956
rect 1471 916 1475 956
rect 1571 916 1575 956
rect 1591 916 1595 956
rect 1725 916 1729 956
rect 1745 916 1749 956
rect 1765 916 1769 956
rect 1865 916 1869 956
rect 1885 916 1889 956
rect 1905 916 1909 956
rect 1991 916 1995 956
rect 2011 916 2015 956
rect 2031 916 2035 956
rect 2136 876 2140 956
rect 2144 876 2148 956
rect 2166 916 2170 956
rect 2271 916 2275 956
rect 2293 916 2297 956
rect 2315 876 2319 956
rect 2411 916 2415 956
rect 2525 916 2529 956
rect 2545 916 2549 956
rect 2655 876 2659 956
rect 2675 876 2679 956
rect 2685 876 2689 956
rect 2771 916 2775 956
rect 2791 916 2795 956
rect 2905 916 2909 956
rect 2925 916 2929 956
rect 3031 916 3035 956
rect 3145 916 3149 956
rect 3265 916 3269 956
rect 3285 916 3289 956
rect 3417 876 3421 956
rect 3425 876 3429 956
rect 3537 876 3541 956
rect 3545 876 3549 956
rect 3645 876 3649 956
rect 3665 876 3669 956
rect 3685 876 3689 956
rect 3785 916 3789 956
rect 3890 916 3894 956
rect 3912 876 3916 956
rect 3920 876 3924 956
rect 4011 916 4015 956
rect 4031 916 4035 956
rect 4150 916 4154 956
rect 4172 876 4176 956
rect 4180 876 4184 956
rect 4290 916 4294 956
rect 4312 876 4316 956
rect 4320 876 4324 956
rect 4431 916 4435 956
rect 4550 916 4554 956
rect 4572 876 4576 956
rect 4580 876 4584 956
rect 4671 876 4675 956
rect 4691 876 4695 956
rect 4711 876 4715 956
rect 4823 876 4827 956
rect 4845 916 4849 956
rect 4950 916 4954 956
rect 4972 876 4976 956
rect 4980 876 4984 956
rect 5071 876 5075 956
rect 5091 876 5095 956
rect 5111 876 5115 956
rect 5235 876 5239 956
rect 5255 876 5259 956
rect 5265 876 5269 956
rect 5385 916 5389 956
rect 5485 876 5489 956
rect 5505 876 5509 956
rect 5525 876 5529 956
rect 5545 876 5549 956
rect 5656 876 5660 956
rect 5664 876 5668 956
rect 5686 916 5690 956
rect 85 504 89 544
rect 105 504 109 544
rect 125 504 129 544
rect 245 504 249 584
rect 265 504 269 584
rect 285 504 289 584
rect 385 504 389 544
rect 405 504 409 544
rect 425 504 429 544
rect 530 504 534 544
rect 552 504 556 584
rect 560 504 564 584
rect 651 504 655 584
rect 671 504 675 584
rect 691 504 695 584
rect 791 504 795 544
rect 811 504 815 544
rect 950 504 954 544
rect 972 504 976 584
rect 980 504 984 584
rect 1085 504 1089 544
rect 1105 504 1109 544
rect 1125 504 1129 544
rect 1211 504 1215 584
rect 1231 504 1235 584
rect 1251 504 1255 584
rect 1365 504 1369 584
rect 1385 504 1389 584
rect 1405 504 1409 584
rect 1511 504 1515 544
rect 1531 504 1535 544
rect 1551 504 1555 544
rect 1670 504 1674 544
rect 1692 504 1696 584
rect 1700 504 1704 584
rect 1805 504 1809 544
rect 1825 504 1829 544
rect 1845 504 1849 544
rect 1931 504 1935 584
rect 1951 504 1955 584
rect 1971 504 1975 584
rect 2097 504 2101 584
rect 2105 504 2109 584
rect 2215 504 2219 584
rect 2235 504 2239 584
rect 2245 504 2249 584
rect 2331 504 2335 544
rect 2353 504 2357 544
rect 2375 504 2379 584
rect 2471 504 2475 544
rect 2491 504 2495 544
rect 2605 504 2609 544
rect 2625 504 2629 544
rect 2737 504 2741 584
rect 2745 504 2749 584
rect 2836 504 2840 584
rect 2844 504 2848 584
rect 2866 504 2870 544
rect 2985 504 2989 544
rect 3005 504 3009 544
rect 3091 504 3095 584
rect 3111 504 3115 584
rect 3131 504 3135 584
rect 3245 504 3249 544
rect 3265 504 3269 544
rect 3285 504 3289 544
rect 3371 504 3375 544
rect 3391 504 3395 544
rect 3510 504 3514 544
rect 3532 504 3536 584
rect 3540 504 3544 584
rect 3631 504 3635 544
rect 3651 504 3655 544
rect 3770 504 3774 544
rect 3792 504 3796 584
rect 3800 504 3804 584
rect 3896 504 3900 584
rect 3904 504 3908 584
rect 3926 504 3930 544
rect 4031 504 4035 584
rect 4051 504 4055 584
rect 4071 504 4075 584
rect 4196 504 4200 584
rect 4204 504 4208 584
rect 4226 504 4230 544
rect 4345 504 4349 544
rect 4445 504 4449 584
rect 4465 504 4469 584
rect 4485 504 4489 584
rect 4590 504 4594 544
rect 4612 504 4616 584
rect 4620 504 4624 584
rect 4730 504 4734 544
rect 4752 504 4756 584
rect 4760 504 4764 584
rect 4876 504 4880 584
rect 4884 504 4888 584
rect 4906 504 4910 544
rect 5011 504 5015 544
rect 5131 504 5135 544
rect 5153 504 5157 584
rect 5270 504 5274 544
rect 5292 504 5296 584
rect 5300 504 5304 584
rect 5396 504 5400 584
rect 5404 504 5408 584
rect 5426 504 5430 544
rect 5550 504 5554 544
rect 5572 504 5576 584
rect 5580 504 5584 584
rect 5671 504 5675 584
rect 5679 504 5683 584
rect 85 436 89 476
rect 105 436 109 476
rect 125 436 129 476
rect 230 436 234 476
rect 252 396 256 476
rect 260 396 264 476
rect 390 436 394 476
rect 412 396 416 476
rect 420 396 424 476
rect 525 436 529 476
rect 545 436 549 476
rect 565 436 569 476
rect 661 396 665 476
rect 683 436 687 476
rect 705 436 709 476
rect 805 436 809 476
rect 825 436 829 476
rect 845 436 849 476
rect 945 396 949 476
rect 965 396 969 476
rect 985 396 989 476
rect 1071 436 1075 476
rect 1091 436 1095 476
rect 1111 436 1115 476
rect 1235 396 1239 476
rect 1255 396 1259 476
rect 1265 396 1269 476
rect 1365 436 1369 476
rect 1385 436 1389 476
rect 1405 436 1409 476
rect 1525 436 1529 476
rect 1630 436 1634 476
rect 1652 396 1656 476
rect 1660 396 1664 476
rect 1761 396 1765 476
rect 1783 436 1787 476
rect 1805 436 1809 476
rect 1891 396 1895 476
rect 1899 396 1903 476
rect 2031 436 2035 476
rect 2150 436 2154 476
rect 2172 396 2176 476
rect 2180 396 2184 476
rect 2285 396 2289 476
rect 2305 396 2309 476
rect 2325 396 2329 476
rect 2425 436 2429 476
rect 2525 436 2529 476
rect 2545 436 2549 476
rect 2565 436 2569 476
rect 2656 396 2660 476
rect 2664 396 2668 476
rect 2686 436 2690 476
rect 2805 436 2809 476
rect 2917 396 2921 476
rect 2925 396 2929 476
rect 3011 436 3015 476
rect 3125 396 3129 476
rect 3145 396 3149 476
rect 3165 396 3169 476
rect 3271 396 3275 476
rect 3291 396 3295 476
rect 3311 396 3315 476
rect 3425 436 3429 476
rect 3536 396 3540 476
rect 3544 396 3548 476
rect 3566 436 3570 476
rect 3671 396 3675 476
rect 3691 396 3695 476
rect 3711 396 3715 476
rect 3825 436 3829 476
rect 3845 436 3849 476
rect 3865 436 3869 476
rect 3951 436 3955 476
rect 3971 436 3975 476
rect 4105 436 4109 476
rect 4125 436 4129 476
rect 4145 436 4149 476
rect 4250 436 4254 476
rect 4272 396 4276 476
rect 4280 396 4284 476
rect 4385 436 4389 476
rect 4485 436 4489 476
rect 4505 436 4509 476
rect 4610 436 4614 476
rect 4632 396 4636 476
rect 4640 396 4644 476
rect 4745 436 4749 476
rect 4850 436 4854 476
rect 4872 396 4876 476
rect 4880 396 4884 476
rect 4971 428 4975 468
rect 4991 388 4995 468
rect 5001 388 5005 468
rect 5021 396 5025 476
rect 5031 396 5035 476
rect 5150 436 5154 476
rect 5172 396 5176 476
rect 5180 396 5184 476
rect 5296 396 5300 476
rect 5304 396 5308 476
rect 5326 436 5330 476
rect 5465 396 5469 476
rect 5485 396 5489 476
rect 5505 396 5509 476
rect 5596 396 5600 476
rect 5604 396 5608 476
rect 5626 436 5630 476
rect 5731 436 5735 476
rect 5751 436 5755 476
rect 85 24 89 64
rect 105 24 109 64
rect 125 24 129 64
rect 211 24 215 104
rect 231 24 235 104
rect 251 24 255 104
rect 385 24 389 104
rect 405 24 409 104
rect 425 24 429 104
rect 530 24 534 64
rect 552 24 556 104
rect 560 24 564 104
rect 656 24 660 104
rect 664 24 668 104
rect 686 24 690 64
rect 805 24 809 64
rect 825 24 829 64
rect 845 24 849 64
rect 931 24 935 64
rect 1036 24 1040 104
rect 1044 24 1048 104
rect 1066 24 1070 64
rect 1171 24 1175 104
rect 1191 24 1195 104
rect 1211 24 1215 104
rect 1311 24 1315 104
rect 1319 24 1323 104
rect 1431 24 1435 64
rect 1453 24 1457 64
rect 1475 24 1479 104
rect 1585 24 1589 64
rect 1690 24 1694 64
rect 1712 24 1716 104
rect 1720 24 1724 104
rect 1825 24 1829 64
rect 1845 24 1849 64
rect 1931 24 1935 64
rect 1951 24 1955 64
rect 1971 24 1975 64
rect 2105 24 2109 64
rect 2125 24 2129 64
rect 2145 24 2149 64
rect 2231 24 2235 64
rect 2253 24 2257 104
rect 2365 24 2369 64
rect 2385 24 2389 64
rect 2471 24 2475 64
rect 2493 24 2497 64
rect 2515 24 2519 104
rect 2625 24 2629 104
rect 2645 24 2649 104
rect 2665 24 2669 104
rect 2761 24 2765 104
rect 2783 24 2787 64
rect 2805 24 2809 64
rect 2911 24 2915 64
rect 2931 24 2935 64
rect 3045 24 3049 64
rect 3065 24 3069 64
rect 3165 24 3169 64
rect 3185 24 3189 64
rect 3205 24 3209 64
rect 3305 24 3309 64
rect 3396 24 3400 104
rect 3404 24 3408 104
rect 3426 24 3430 64
rect 3545 24 3549 64
rect 3645 24 3649 64
rect 3665 24 3669 64
rect 3763 24 3767 104
rect 3785 24 3789 64
rect 3871 24 3875 64
rect 3893 24 3897 104
rect 4005 24 4009 64
rect 4025 24 4029 64
rect 4131 24 4135 64
rect 4153 24 4157 64
rect 4175 24 4179 104
rect 4317 24 4321 104
rect 4325 24 4329 104
rect 4411 24 4415 64
rect 4431 24 4435 64
rect 4545 24 4549 64
rect 4565 24 4569 64
rect 4585 24 4589 64
rect 4710 24 4714 64
rect 4732 24 4736 104
rect 4740 24 4744 104
rect 4831 24 4835 64
rect 4851 24 4855 64
rect 4970 24 4974 64
rect 4992 24 4996 104
rect 5000 24 5004 104
rect 5091 24 5095 104
rect 5099 24 5103 104
rect 5225 24 5229 64
rect 5245 24 5249 64
rect 5331 32 5335 72
rect 5351 32 5355 112
rect 5361 32 5365 112
rect 5381 24 5385 104
rect 5391 24 5395 104
rect 5491 24 5495 64
rect 5605 24 5609 64
rect 5691 24 5695 64
rect 5711 24 5715 64
<< ndiffusion >>
rect 83 5544 85 5584
rect 89 5544 91 5584
rect 103 5544 105 5584
rect 109 5572 125 5584
rect 109 5544 111 5572
rect 123 5544 125 5572
rect 129 5544 131 5584
rect 209 5544 211 5584
rect 215 5572 231 5584
rect 215 5544 217 5572
rect 229 5544 231 5572
rect 235 5544 237 5584
rect 249 5544 251 5584
rect 255 5544 257 5584
rect 390 5544 392 5564
rect 396 5544 400 5564
rect 412 5544 414 5584
rect 418 5544 422 5584
rect 426 5544 428 5584
rect 510 5544 512 5604
rect 516 5544 520 5604
rect 524 5544 528 5604
rect 532 5602 546 5604
rect 532 5544 534 5602
rect 663 5544 665 5584
rect 669 5544 671 5584
rect 683 5544 685 5584
rect 689 5572 705 5584
rect 689 5544 691 5572
rect 703 5544 705 5572
rect 709 5544 711 5584
rect 811 5544 813 5584
rect 817 5544 823 5584
rect 827 5544 829 5584
rect 930 5544 932 5564
rect 936 5544 940 5564
rect 952 5544 954 5584
rect 958 5544 962 5584
rect 966 5544 968 5584
rect 1069 5544 1071 5564
rect 1075 5544 1077 5564
rect 1089 5544 1091 5564
rect 1095 5544 1097 5564
rect 1223 5544 1225 5584
rect 1229 5564 1241 5584
rect 1514 5602 1528 5604
rect 1229 5544 1231 5564
rect 1243 5544 1245 5564
rect 1249 5544 1251 5564
rect 1263 5544 1265 5564
rect 1269 5544 1271 5564
rect 1373 5544 1375 5584
rect 1379 5544 1381 5584
rect 1393 5544 1395 5584
rect 1399 5544 1405 5584
rect 1409 5544 1411 5584
rect 1526 5544 1528 5602
rect 1532 5544 1536 5604
rect 1540 5544 1544 5604
rect 1548 5544 1550 5604
rect 1814 5602 1828 5604
rect 1670 5544 1672 5564
rect 1676 5544 1680 5564
rect 1692 5544 1694 5584
rect 1698 5544 1702 5584
rect 1706 5544 1708 5584
rect 1826 5544 1828 5602
rect 1832 5544 1836 5604
rect 1840 5544 1844 5604
rect 1848 5544 1850 5604
rect 1929 5544 1931 5564
rect 1935 5544 1937 5564
rect 2043 5544 2045 5584
rect 2049 5544 2051 5584
rect 2063 5544 2065 5584
rect 2069 5572 2085 5584
rect 2069 5544 2071 5572
rect 2083 5544 2085 5572
rect 2089 5544 2091 5584
rect 2169 5544 2171 5584
rect 2175 5572 2191 5584
rect 2175 5544 2177 5572
rect 2189 5544 2191 5572
rect 2195 5544 2197 5584
rect 2209 5544 2211 5584
rect 2215 5544 2217 5584
rect 2312 5544 2314 5584
rect 2318 5544 2322 5584
rect 2326 5544 2328 5584
rect 2594 5602 2608 5604
rect 2340 5544 2344 5564
rect 2348 5544 2350 5564
rect 2471 5544 2473 5584
rect 2477 5544 2483 5584
rect 2487 5544 2489 5584
rect 2606 5544 2608 5602
rect 2612 5544 2616 5604
rect 2620 5544 2624 5604
rect 2628 5544 2630 5604
rect 2734 5602 2748 5604
rect 2746 5544 2748 5602
rect 2752 5544 2756 5604
rect 2760 5544 2764 5604
rect 2768 5544 2770 5604
rect 2851 5544 2853 5584
rect 2857 5544 2863 5584
rect 2867 5544 2869 5584
rect 2983 5544 2985 5564
rect 2989 5544 2991 5564
rect 3083 5544 3085 5584
rect 3089 5544 3091 5584
rect 3103 5544 3105 5584
rect 3109 5572 3125 5584
rect 3109 5544 3111 5572
rect 3123 5544 3125 5572
rect 3129 5544 3131 5584
rect 3253 5544 3255 5584
rect 3259 5544 3261 5584
rect 3273 5544 3275 5584
rect 3279 5544 3285 5584
rect 3289 5544 3291 5584
rect 3514 5602 3528 5604
rect 3383 5544 3385 5564
rect 3389 5544 3391 5564
rect 3403 5544 3405 5564
rect 3409 5544 3411 5564
rect 3526 5544 3528 5602
rect 3532 5544 3536 5604
rect 3540 5544 3544 5604
rect 3548 5544 3550 5604
rect 3663 5544 3665 5564
rect 3669 5544 3671 5564
rect 3763 5544 3765 5564
rect 3769 5544 3771 5564
rect 3849 5544 3851 5564
rect 3855 5544 3857 5564
rect 3949 5544 3951 5584
rect 3955 5572 3971 5584
rect 3955 5544 3957 5572
rect 3969 5544 3971 5572
rect 3975 5544 3977 5584
rect 3989 5544 3991 5584
rect 3995 5544 3997 5584
rect 4089 5544 4091 5564
rect 4095 5544 4097 5564
rect 4149 5544 4151 5584
rect 4155 5564 4168 5584
rect 4331 5564 4341 5584
rect 4155 5544 4159 5564
rect 4171 5544 4173 5564
rect 4177 5544 4183 5564
rect 4187 5544 4189 5564
rect 4201 5544 4203 5564
rect 4207 5544 4211 5564
rect 4215 5544 4217 5564
rect 4255 5544 4257 5564
rect 4261 5544 4265 5564
rect 4277 5544 4279 5564
rect 4283 5544 4289 5564
rect 4293 5544 4295 5564
rect 4307 5544 4311 5564
rect 4315 5544 4321 5564
rect 4325 5544 4327 5564
rect 4339 5544 4341 5564
rect 4345 5544 4347 5584
rect 4463 5544 4465 5584
rect 4469 5544 4471 5584
rect 4483 5544 4485 5584
rect 4489 5572 4505 5584
rect 4489 5544 4491 5572
rect 4503 5544 4505 5572
rect 4509 5544 4511 5584
rect 4603 5544 4605 5584
rect 4609 5544 4611 5584
rect 4623 5544 4625 5584
rect 4629 5544 4631 5584
rect 4643 5544 4645 5584
rect 4649 5544 4651 5584
rect 4663 5544 4665 5584
rect 4669 5544 4671 5584
rect 4683 5544 4685 5584
rect 4689 5544 4691 5584
rect 4703 5544 4705 5584
rect 4709 5544 4711 5584
rect 4723 5544 4725 5584
rect 4729 5544 4731 5584
rect 4743 5544 4745 5584
rect 4749 5544 4751 5584
rect 4843 5544 4845 5564
rect 4849 5544 4851 5564
rect 4943 5544 4945 5584
rect 4949 5544 4951 5584
rect 4963 5544 4965 5584
rect 4969 5572 4985 5584
rect 4969 5544 4971 5572
rect 4983 5544 4985 5572
rect 4989 5544 4991 5584
rect 5091 5544 5093 5584
rect 5097 5544 5103 5584
rect 5107 5544 5109 5584
rect 5191 5544 5193 5584
rect 5197 5544 5203 5584
rect 5207 5544 5209 5584
rect 5309 5544 5311 5584
rect 5315 5572 5331 5584
rect 5315 5544 5317 5572
rect 5329 5544 5331 5572
rect 5335 5544 5337 5584
rect 5349 5544 5351 5584
rect 5355 5544 5357 5584
rect 5449 5544 5451 5564
rect 5455 5544 5457 5564
rect 5551 5544 5553 5584
rect 5557 5544 5563 5584
rect 5567 5544 5569 5584
rect 5669 5544 5671 5564
rect 5675 5544 5677 5564
rect 83 5476 85 5516
rect 89 5476 91 5516
rect 103 5476 105 5516
rect 109 5488 111 5516
rect 123 5488 125 5516
rect 109 5476 125 5488
rect 129 5476 131 5516
rect 266 5458 268 5516
rect 254 5456 268 5458
rect 272 5456 276 5516
rect 280 5456 284 5516
rect 288 5456 290 5516
rect 406 5458 408 5516
rect 394 5456 408 5458
rect 412 5456 416 5516
rect 420 5456 424 5516
rect 428 5456 430 5516
rect 546 5458 548 5516
rect 534 5456 548 5458
rect 552 5456 556 5516
rect 560 5456 564 5516
rect 568 5456 570 5516
rect 670 5456 672 5516
rect 676 5456 680 5516
rect 684 5456 688 5516
rect 692 5458 694 5516
rect 809 5476 811 5516
rect 815 5488 817 5516
rect 829 5488 831 5516
rect 815 5476 831 5488
rect 835 5476 837 5516
rect 849 5476 851 5516
rect 855 5476 857 5516
rect 692 5456 706 5458
rect 950 5456 952 5516
rect 956 5456 960 5516
rect 964 5456 968 5516
rect 972 5458 974 5516
rect 1110 5496 1112 5516
rect 1116 5496 1120 5516
rect 972 5456 986 5458
rect 1132 5476 1134 5516
rect 1138 5476 1142 5516
rect 1146 5476 1148 5516
rect 1230 5456 1232 5516
rect 1236 5456 1240 5516
rect 1244 5456 1248 5516
rect 1252 5458 1254 5516
rect 1389 5496 1391 5516
rect 1395 5496 1397 5516
rect 1409 5496 1411 5516
rect 1415 5496 1417 5516
rect 1252 5456 1266 5458
rect 1546 5458 1548 5516
rect 1534 5456 1548 5458
rect 1552 5456 1556 5516
rect 1560 5456 1564 5516
rect 1568 5456 1570 5516
rect 1649 5476 1651 5516
rect 1655 5488 1657 5516
rect 1669 5488 1671 5516
rect 1655 5476 1671 5488
rect 1675 5476 1677 5516
rect 1689 5476 1691 5516
rect 1695 5476 1697 5516
rect 1826 5458 1828 5516
rect 1814 5456 1828 5458
rect 1832 5456 1836 5516
rect 1840 5456 1844 5516
rect 1848 5456 1850 5516
rect 1966 5458 1968 5516
rect 1954 5456 1968 5458
rect 1972 5456 1976 5516
rect 1980 5456 1984 5516
rect 1988 5456 1990 5516
rect 2071 5476 2073 5516
rect 2077 5476 2083 5516
rect 2087 5476 2089 5516
rect 2223 5496 2225 5516
rect 2229 5496 2231 5516
rect 2333 5476 2335 5516
rect 2339 5476 2341 5516
rect 2353 5476 2355 5516
rect 2359 5476 2365 5516
rect 2369 5476 2371 5516
rect 2449 5476 2451 5516
rect 2455 5488 2457 5516
rect 2469 5488 2471 5516
rect 2455 5476 2471 5488
rect 2475 5476 2477 5516
rect 2489 5476 2491 5516
rect 2495 5476 2497 5516
rect 2646 5458 2648 5516
rect 2634 5456 2648 5458
rect 2652 5456 2656 5516
rect 2660 5456 2664 5516
rect 2668 5456 2670 5516
rect 2786 5458 2788 5516
rect 2774 5456 2788 5458
rect 2792 5456 2796 5516
rect 2800 5456 2804 5516
rect 2808 5456 2810 5516
rect 2889 5476 2891 5516
rect 2895 5488 2897 5516
rect 2909 5488 2911 5516
rect 2895 5476 2911 5488
rect 2915 5476 2917 5516
rect 2929 5476 2931 5516
rect 2935 5476 2937 5516
rect 3029 5496 3031 5516
rect 3035 5496 3037 5516
rect 3131 5476 3133 5516
rect 3137 5476 3143 5516
rect 3147 5476 3149 5516
rect 3270 5456 3272 5516
rect 3276 5456 3280 5516
rect 3284 5456 3288 5516
rect 3292 5458 3294 5516
rect 3411 5476 3413 5516
rect 3417 5476 3423 5516
rect 3427 5476 3429 5516
rect 3529 5496 3531 5516
rect 3535 5496 3537 5516
rect 3549 5496 3551 5516
rect 3555 5496 3557 5516
rect 3569 5496 3571 5516
rect 3292 5456 3306 5458
rect 3559 5476 3571 5496
rect 3575 5476 3577 5516
rect 3706 5458 3708 5516
rect 3694 5456 3708 5458
rect 3712 5456 3716 5516
rect 3720 5456 3724 5516
rect 3728 5456 3730 5516
rect 3830 5496 3832 5516
rect 3836 5496 3840 5516
rect 3852 5476 3854 5516
rect 3858 5476 3862 5516
rect 3866 5476 3868 5516
rect 3951 5476 3953 5516
rect 3957 5476 3963 5516
rect 3967 5476 3969 5516
rect 4083 5476 4085 5516
rect 4089 5476 4091 5516
rect 4103 5476 4105 5516
rect 4109 5488 4111 5516
rect 4123 5488 4125 5516
rect 4109 5476 4125 5488
rect 4129 5476 4131 5516
rect 4231 5476 4233 5516
rect 4237 5476 4243 5516
rect 4247 5476 4249 5516
rect 4366 5458 4368 5516
rect 4354 5456 4368 5458
rect 4372 5456 4376 5516
rect 4380 5456 4384 5516
rect 4388 5456 4390 5516
rect 4492 5476 4494 5516
rect 4498 5476 4502 5516
rect 4506 5476 4508 5516
rect 4520 5496 4524 5516
rect 4528 5496 4530 5516
rect 4629 5496 4631 5516
rect 4635 5496 4637 5516
rect 4729 5476 4731 5516
rect 4735 5488 4737 5516
rect 4749 5488 4751 5516
rect 4735 5476 4751 5488
rect 4755 5476 4757 5516
rect 4769 5476 4771 5516
rect 4775 5476 4777 5516
rect 4829 5476 4831 5516
rect 4835 5496 4839 5516
rect 4851 5496 4853 5516
rect 4857 5496 4863 5516
rect 4867 5496 4869 5516
rect 4881 5496 4883 5516
rect 4887 5496 4891 5516
rect 4895 5496 4897 5516
rect 4935 5496 4937 5516
rect 4941 5496 4945 5516
rect 4957 5496 4959 5516
rect 4963 5496 4969 5516
rect 4973 5496 4975 5516
rect 4987 5496 4991 5516
rect 4995 5496 5001 5516
rect 5005 5496 5007 5516
rect 5019 5496 5021 5516
rect 4835 5476 4848 5496
rect 5011 5476 5021 5496
rect 5025 5476 5027 5516
rect 5109 5496 5111 5516
rect 5115 5496 5117 5516
rect 5169 5476 5171 5516
rect 5175 5496 5179 5516
rect 5191 5496 5193 5516
rect 5197 5496 5203 5516
rect 5207 5496 5209 5516
rect 5221 5496 5223 5516
rect 5227 5496 5231 5516
rect 5235 5496 5237 5516
rect 5275 5496 5277 5516
rect 5281 5496 5285 5516
rect 5297 5496 5299 5516
rect 5303 5496 5309 5516
rect 5313 5496 5315 5516
rect 5327 5496 5331 5516
rect 5335 5496 5341 5516
rect 5345 5496 5347 5516
rect 5359 5496 5361 5516
rect 5175 5476 5188 5496
rect 5351 5476 5361 5496
rect 5365 5476 5367 5516
rect 5449 5476 5451 5516
rect 5455 5488 5457 5516
rect 5469 5488 5471 5516
rect 5455 5476 5471 5488
rect 5475 5476 5477 5516
rect 5489 5476 5491 5516
rect 5495 5476 5497 5516
rect 5611 5476 5613 5516
rect 5617 5476 5623 5516
rect 5627 5476 5629 5516
rect 5731 5476 5733 5516
rect 5737 5476 5743 5516
rect 5747 5476 5749 5516
rect 94 5122 108 5124
rect 106 5064 108 5122
rect 112 5064 116 5124
rect 120 5064 124 5124
rect 128 5064 130 5124
rect 212 5064 214 5104
rect 218 5064 222 5104
rect 226 5064 228 5104
rect 474 5122 488 5124
rect 240 5064 244 5084
rect 248 5064 250 5084
rect 349 5064 351 5084
rect 355 5064 357 5084
rect 486 5064 488 5122
rect 492 5064 496 5124
rect 500 5064 504 5124
rect 508 5064 510 5124
rect 592 5064 594 5104
rect 598 5064 602 5104
rect 606 5064 608 5104
rect 620 5064 624 5084
rect 628 5064 630 5084
rect 750 5064 752 5084
rect 756 5064 760 5084
rect 772 5064 774 5104
rect 778 5064 782 5104
rect 786 5064 788 5104
rect 870 5064 872 5124
rect 876 5064 880 5124
rect 884 5064 888 5124
rect 892 5122 906 5124
rect 892 5064 894 5122
rect 1034 5122 1048 5124
rect 1046 5064 1048 5122
rect 1052 5064 1056 5124
rect 1060 5064 1064 5124
rect 1068 5064 1070 5124
rect 1274 5122 1288 5124
rect 1149 5064 1151 5084
rect 1155 5064 1157 5084
rect 1286 5064 1288 5122
rect 1292 5064 1296 5124
rect 1300 5064 1304 5124
rect 1308 5064 1310 5124
rect 1423 5064 1425 5104
rect 1429 5064 1431 5104
rect 1443 5064 1445 5104
rect 1449 5092 1465 5104
rect 1449 5064 1451 5092
rect 1463 5064 1465 5092
rect 1469 5064 1471 5104
rect 1563 5064 1565 5084
rect 1569 5064 1571 5084
rect 1663 5064 1665 5104
rect 1669 5064 1671 5104
rect 1683 5064 1685 5104
rect 1689 5092 1705 5104
rect 1689 5064 1691 5092
rect 1703 5064 1705 5092
rect 1709 5064 1711 5104
rect 2334 5122 2348 5124
rect 1883 5064 1885 5084
rect 1889 5064 1891 5084
rect 1903 5064 1905 5084
rect 1909 5064 1911 5084
rect 1923 5064 1925 5084
rect 1929 5064 1931 5084
rect 2064 5064 2066 5104
rect 2070 5064 2074 5104
rect 2078 5064 2080 5104
rect 2092 5064 2094 5104
rect 2098 5064 2102 5104
rect 2106 5064 2108 5104
rect 2191 5064 2193 5104
rect 2197 5064 2203 5104
rect 2207 5064 2209 5104
rect 2346 5064 2348 5122
rect 2352 5064 2356 5124
rect 2360 5064 2364 5124
rect 2368 5064 2370 5124
rect 2470 5064 2472 5084
rect 2476 5064 2480 5084
rect 2492 5064 2494 5104
rect 2498 5064 2502 5104
rect 2506 5064 2508 5104
rect 2603 5064 2605 5084
rect 2609 5064 2611 5084
rect 2703 5064 2705 5104
rect 2709 5064 2711 5104
rect 2723 5064 2725 5104
rect 2729 5092 2745 5104
rect 2729 5064 2731 5092
rect 2743 5064 2745 5092
rect 2749 5064 2751 5104
rect 2863 5064 2865 5104
rect 2869 5064 2871 5104
rect 2883 5064 2885 5104
rect 2889 5092 2905 5104
rect 2889 5064 2891 5092
rect 2903 5064 2905 5092
rect 2909 5064 2911 5104
rect 3013 5064 3015 5104
rect 3019 5064 3021 5104
rect 3033 5064 3035 5104
rect 3039 5064 3045 5104
rect 3049 5064 3051 5104
rect 3129 5064 3131 5084
rect 3135 5064 3137 5084
rect 3149 5064 3151 5084
rect 3155 5064 3157 5084
rect 3283 5064 3285 5084
rect 3289 5064 3291 5084
rect 3383 5064 3385 5084
rect 3389 5064 3391 5084
rect 3403 5064 3405 5084
rect 3409 5064 3411 5084
rect 3523 5064 3525 5104
rect 3529 5064 3531 5104
rect 3543 5064 3545 5104
rect 3549 5092 3565 5104
rect 3549 5064 3551 5092
rect 3563 5064 3565 5092
rect 3569 5064 3571 5104
rect 3651 5064 3653 5104
rect 3657 5064 3663 5104
rect 3667 5064 3669 5104
rect 3791 5064 3793 5104
rect 3797 5064 3803 5104
rect 3807 5064 3809 5104
rect 3931 5064 3933 5104
rect 3937 5064 3943 5104
rect 3947 5064 3949 5104
rect 4030 5064 4032 5124
rect 4036 5064 4040 5124
rect 4044 5064 4048 5124
rect 4052 5122 4066 5124
rect 4052 5064 4054 5122
rect 4183 5064 4185 5104
rect 4189 5064 4191 5104
rect 4203 5064 4205 5104
rect 4209 5092 4225 5104
rect 4209 5064 4211 5092
rect 4223 5064 4225 5092
rect 4229 5064 4231 5104
rect 4329 5064 4331 5104
rect 4335 5092 4351 5104
rect 4335 5064 4337 5092
rect 4349 5064 4351 5092
rect 4355 5064 4357 5104
rect 4369 5064 4371 5104
rect 4375 5064 4377 5104
rect 4594 5122 4608 5124
rect 4469 5064 4471 5084
rect 4475 5064 4477 5084
rect 4606 5064 4608 5122
rect 4612 5064 4616 5124
rect 4620 5064 4624 5124
rect 4628 5064 4630 5124
rect 4712 5064 4714 5104
rect 4718 5064 4722 5104
rect 4726 5064 4728 5104
rect 4740 5064 4744 5084
rect 4748 5064 4750 5084
rect 4849 5064 4851 5084
rect 4855 5064 4857 5084
rect 4869 5064 4871 5084
rect 4875 5064 4877 5084
rect 4929 5064 4931 5104
rect 4935 5084 4948 5104
rect 5111 5084 5121 5104
rect 4935 5064 4939 5084
rect 4951 5064 4953 5084
rect 4957 5064 4963 5084
rect 4967 5064 4969 5084
rect 4981 5064 4983 5084
rect 4987 5064 4991 5084
rect 4995 5064 4997 5084
rect 5035 5064 5037 5084
rect 5041 5064 5045 5084
rect 5057 5064 5059 5084
rect 5063 5064 5069 5084
rect 5073 5064 5075 5084
rect 5087 5064 5091 5084
rect 5095 5064 5101 5084
rect 5105 5064 5107 5084
rect 5119 5064 5121 5084
rect 5125 5064 5127 5104
rect 5209 5064 5211 5104
rect 5215 5092 5231 5104
rect 5215 5064 5217 5092
rect 5229 5064 5231 5092
rect 5235 5064 5237 5104
rect 5249 5064 5251 5104
rect 5255 5064 5257 5104
rect 5349 5064 5351 5084
rect 5355 5064 5357 5084
rect 5449 5064 5451 5104
rect 5455 5092 5471 5104
rect 5455 5064 5457 5092
rect 5469 5064 5471 5092
rect 5475 5064 5477 5104
rect 5489 5064 5491 5104
rect 5495 5064 5497 5104
rect 5611 5064 5613 5104
rect 5617 5064 5623 5104
rect 5627 5064 5629 5104
rect 5711 5064 5713 5104
rect 5717 5064 5723 5104
rect 5727 5064 5729 5104
rect 83 4996 85 5036
rect 89 4996 91 5036
rect 103 4996 105 5036
rect 109 5008 111 5036
rect 123 5008 125 5036
rect 109 4996 125 5008
rect 129 4996 131 5036
rect 246 4978 248 5036
rect 234 4976 248 4978
rect 252 4976 256 5036
rect 260 4976 264 5036
rect 268 4976 270 5036
rect 350 4976 352 5036
rect 356 4976 360 5036
rect 364 4976 368 5036
rect 372 4978 374 5036
rect 489 4996 491 5036
rect 495 5008 497 5036
rect 509 5008 511 5036
rect 495 4996 511 5008
rect 515 4996 517 5036
rect 529 4996 531 5036
rect 535 4996 537 5036
rect 651 4996 653 5036
rect 657 4996 663 5036
rect 667 4996 669 5036
rect 763 4996 765 5036
rect 769 4996 771 5036
rect 783 4996 785 5036
rect 789 5008 791 5036
rect 803 5008 805 5036
rect 789 4996 805 5008
rect 809 4996 811 5036
rect 903 4996 905 5036
rect 909 4996 911 5036
rect 923 4996 925 5036
rect 929 5008 931 5036
rect 943 5008 945 5036
rect 929 4996 945 5008
rect 949 4996 951 5036
rect 1050 5016 1052 5036
rect 1056 5016 1060 5036
rect 372 4976 386 4978
rect 1072 4996 1074 5036
rect 1078 4996 1082 5036
rect 1086 4996 1088 5036
rect 1183 4996 1185 5036
rect 1189 4996 1191 5036
rect 1203 4996 1205 5036
rect 1209 5008 1211 5036
rect 1223 5008 1225 5036
rect 1209 4996 1225 5008
rect 1229 4996 1231 5036
rect 1323 5016 1325 5036
rect 1329 5016 1331 5036
rect 1431 4996 1433 5036
rect 1437 4996 1443 5036
rect 1447 4996 1449 5036
rect 1586 4978 1588 5036
rect 1574 4976 1588 4978
rect 1592 4976 1596 5036
rect 1600 4976 1604 5036
rect 1608 4976 1610 5036
rect 1703 4996 1705 5036
rect 1709 4996 1711 5036
rect 1723 4996 1725 5036
rect 1729 5008 1731 5036
rect 1743 5008 1745 5036
rect 1729 4996 1745 5008
rect 1749 4996 1751 5036
rect 1832 4996 1834 5036
rect 1838 4996 1842 5036
rect 1846 4996 1848 5036
rect 1860 5016 1864 5036
rect 1868 5016 1870 5036
rect 1971 4996 1973 5036
rect 1977 4996 1983 5036
rect 1987 4996 1989 5036
rect 2110 5016 2112 5036
rect 2116 5016 2120 5036
rect 2132 4996 2134 5036
rect 2138 4996 2142 5036
rect 2146 4996 2148 5036
rect 2263 5016 2265 5036
rect 2269 5016 2271 5036
rect 2363 4996 2365 5036
rect 2369 4996 2371 5036
rect 2383 4996 2385 5036
rect 2389 5008 2391 5036
rect 2403 5008 2405 5036
rect 2389 4996 2405 5008
rect 2409 4996 2411 5036
rect 2526 4978 2528 5036
rect 2514 4976 2528 4978
rect 2532 4976 2536 5036
rect 2540 4976 2544 5036
rect 2548 4976 2550 5036
rect 2643 5016 2645 5036
rect 2649 5016 2651 5036
rect 2771 4996 2773 5036
rect 2777 4996 2783 5036
rect 2787 4996 2789 5036
rect 2869 5016 2871 5036
rect 2875 5016 2877 5036
rect 2970 4976 2972 5036
rect 2976 4976 2980 5036
rect 2984 4976 2988 5036
rect 2992 4978 2994 5036
rect 3123 4996 3125 5036
rect 3129 4996 3131 5036
rect 3143 4996 3145 5036
rect 3149 5008 3151 5036
rect 3163 5008 3165 5036
rect 3149 4996 3165 5008
rect 3169 4996 3171 5036
rect 3263 4996 3265 5036
rect 3269 4996 3271 5036
rect 3283 4996 3285 5036
rect 3289 5008 3291 5036
rect 3303 5008 3305 5036
rect 3289 4996 3305 5008
rect 3309 4996 3311 5036
rect 3410 5016 3412 5036
rect 3416 5016 3420 5036
rect 2992 4976 3006 4978
rect 3432 4996 3434 5036
rect 3438 4996 3442 5036
rect 3446 4996 3448 5036
rect 3529 5016 3531 5036
rect 3535 5016 3537 5036
rect 3549 5016 3551 5036
rect 3555 5016 3557 5036
rect 3569 5016 3571 5036
rect 3559 4996 3571 5016
rect 3575 4996 3577 5036
rect 3683 5016 3685 5036
rect 3689 5016 3691 5036
rect 3703 5016 3705 5036
rect 3709 5016 3711 5036
rect 3826 4978 3828 5036
rect 3814 4976 3828 4978
rect 3832 4976 3836 5036
rect 3840 4976 3844 5036
rect 3848 4976 3850 5036
rect 3943 5016 3945 5036
rect 3949 5016 3951 5036
rect 4030 4976 4032 5036
rect 4036 4976 4040 5036
rect 4044 4976 4048 5036
rect 4052 4978 4054 5036
rect 4052 4976 4066 4978
rect 4170 4976 4172 5036
rect 4176 4976 4180 5036
rect 4184 4976 4188 5036
rect 4192 4978 4194 5036
rect 4333 4996 4335 5036
rect 4339 4996 4341 5036
rect 4353 4996 4355 5036
rect 4359 4996 4365 5036
rect 4369 4996 4371 5036
rect 4469 5016 4471 5036
rect 4475 5016 4477 5036
rect 4489 5016 4491 5036
rect 4495 5016 4497 5036
rect 4509 5016 4511 5036
rect 4192 4976 4206 4978
rect 4499 4996 4511 5016
rect 4515 4996 4517 5036
rect 4609 5016 4611 5036
rect 4615 5016 4617 5036
rect 4629 5016 4631 5036
rect 4635 5016 4637 5036
rect 4743 4996 4745 5036
rect 4749 4996 4751 5036
rect 4763 4996 4765 5036
rect 4769 5008 4771 5036
rect 4783 5008 4785 5036
rect 4769 4996 4785 5008
rect 4789 4996 4791 5036
rect 4829 4996 4831 5036
rect 4835 5016 4839 5036
rect 4851 5016 4853 5036
rect 4857 5016 4863 5036
rect 4867 5016 4869 5036
rect 4881 5016 4883 5036
rect 4887 5016 4891 5036
rect 4895 5016 4897 5036
rect 4935 5016 4937 5036
rect 4941 5016 4945 5036
rect 4957 5016 4959 5036
rect 4963 5016 4969 5036
rect 4973 5016 4975 5036
rect 4987 5016 4991 5036
rect 4995 5016 5001 5036
rect 5005 5016 5007 5036
rect 5019 5016 5021 5036
rect 4835 4996 4848 5016
rect 5011 4996 5021 5016
rect 5025 4996 5027 5036
rect 5109 4996 5111 5036
rect 5115 5008 5117 5036
rect 5129 5008 5131 5036
rect 5115 4996 5131 5008
rect 5135 4996 5137 5036
rect 5149 4996 5151 5036
rect 5155 4996 5157 5036
rect 5209 4996 5211 5036
rect 5215 5016 5219 5036
rect 5231 5016 5233 5036
rect 5237 5016 5243 5036
rect 5247 5016 5249 5036
rect 5261 5016 5263 5036
rect 5267 5016 5271 5036
rect 5275 5016 5277 5036
rect 5315 5016 5317 5036
rect 5321 5016 5325 5036
rect 5337 5016 5339 5036
rect 5343 5016 5349 5036
rect 5353 5016 5355 5036
rect 5367 5016 5371 5036
rect 5375 5016 5381 5036
rect 5385 5016 5387 5036
rect 5399 5016 5401 5036
rect 5215 4996 5228 5016
rect 5391 4996 5401 5016
rect 5405 4996 5407 5036
rect 5511 4996 5513 5036
rect 5517 4996 5523 5036
rect 5527 4996 5529 5036
rect 5611 4996 5613 5036
rect 5617 4996 5623 5036
rect 5627 4996 5629 5036
rect 5751 4996 5753 5036
rect 5757 4996 5763 5036
rect 5767 4996 5769 5036
rect 234 4642 248 4644
rect 90 4584 92 4604
rect 96 4584 100 4604
rect 112 4584 114 4624
rect 118 4584 122 4624
rect 126 4584 128 4624
rect 246 4584 248 4642
rect 252 4584 256 4644
rect 260 4584 264 4644
rect 268 4584 270 4644
rect 352 4584 354 4624
rect 358 4584 362 4624
rect 366 4584 368 4624
rect 634 4642 648 4644
rect 380 4584 384 4604
rect 388 4584 390 4604
rect 491 4584 493 4624
rect 497 4584 503 4624
rect 507 4584 509 4624
rect 646 4584 648 4642
rect 652 4584 656 4644
rect 660 4584 664 4644
rect 668 4584 670 4644
rect 794 4642 808 4644
rect 806 4584 808 4642
rect 812 4584 816 4644
rect 820 4584 824 4644
rect 828 4584 830 4644
rect 909 4584 911 4604
rect 915 4584 917 4604
rect 1009 4584 1011 4604
rect 1015 4584 1017 4604
rect 1123 4584 1125 4604
rect 1129 4584 1131 4604
rect 1223 4584 1225 4624
rect 1229 4584 1231 4624
rect 1243 4584 1245 4624
rect 1249 4612 1265 4624
rect 1249 4584 1251 4612
rect 1263 4584 1265 4612
rect 1269 4584 1271 4624
rect 1349 4584 1351 4624
rect 1355 4612 1371 4624
rect 1355 4584 1357 4612
rect 1369 4584 1371 4612
rect 1375 4584 1377 4624
rect 1389 4584 1391 4624
rect 1395 4584 1397 4624
rect 1489 4584 1491 4604
rect 1495 4584 1497 4604
rect 1590 4584 1592 4644
rect 1596 4584 1600 4644
rect 1604 4584 1608 4644
rect 1612 4642 1626 4644
rect 1612 4584 1614 4642
rect 2154 4642 2168 4644
rect 1743 4584 1745 4624
rect 1749 4584 1751 4624
rect 1763 4584 1765 4624
rect 1769 4612 1785 4624
rect 1769 4584 1771 4612
rect 1783 4584 1785 4612
rect 1789 4584 1791 4624
rect 1891 4584 1893 4624
rect 1897 4584 1903 4624
rect 1907 4584 1909 4624
rect 1989 4584 1991 4624
rect 1995 4612 2011 4624
rect 1995 4584 1997 4612
rect 2009 4584 2011 4612
rect 2015 4584 2017 4624
rect 2029 4584 2031 4624
rect 2035 4584 2037 4624
rect 2166 4584 2168 4642
rect 2172 4584 2176 4644
rect 2180 4584 2184 4644
rect 2188 4584 2190 4644
rect 2281 4584 2283 4624
rect 2287 4584 2289 4624
rect 2301 4584 2305 4604
rect 2309 4584 2311 4604
rect 2391 4584 2393 4624
rect 2397 4584 2403 4624
rect 2407 4584 2409 4624
rect 2511 4584 2513 4624
rect 2517 4584 2523 4624
rect 2527 4584 2529 4624
rect 2641 4584 2643 4624
rect 2647 4584 2649 4624
rect 2661 4584 2665 4604
rect 2669 4584 2671 4604
rect 2750 4584 2752 4644
rect 2756 4584 2760 4644
rect 2764 4584 2768 4644
rect 2772 4642 2786 4644
rect 2772 4584 2774 4642
rect 3334 4642 3348 4644
rect 2903 4584 2905 4604
rect 2909 4584 2911 4604
rect 2923 4584 2925 4604
rect 2929 4584 2931 4604
rect 3029 4584 3031 4624
rect 3035 4614 3051 4624
rect 3035 4584 3037 4614
rect 3049 4584 3051 4614
rect 3055 4584 3057 4624
rect 3069 4584 3071 4624
rect 3075 4596 3077 4624
rect 3089 4596 3091 4624
rect 3075 4584 3091 4596
rect 3095 4584 3097 4624
rect 3211 4584 3213 4624
rect 3217 4584 3223 4624
rect 3227 4584 3229 4624
rect 3346 4584 3348 4642
rect 3352 4584 3356 4644
rect 3360 4584 3364 4644
rect 3368 4584 3370 4644
rect 3614 4642 3628 4644
rect 3470 4584 3472 4604
rect 3476 4584 3480 4604
rect 3492 4584 3494 4624
rect 3498 4584 3502 4624
rect 3506 4584 3508 4624
rect 3626 4584 3628 4642
rect 3632 4584 3636 4644
rect 3640 4584 3644 4644
rect 3648 4584 3650 4644
rect 3750 4584 3752 4604
rect 3756 4584 3760 4604
rect 3772 4584 3774 4624
rect 3778 4584 3782 4624
rect 3786 4584 3788 4624
rect 3870 4584 3872 4644
rect 3876 4584 3880 4644
rect 3884 4584 3888 4644
rect 3892 4642 3906 4644
rect 3892 4584 3894 4642
rect 4010 4584 4012 4644
rect 4016 4584 4020 4644
rect 4024 4584 4028 4644
rect 4032 4642 4046 4644
rect 4032 4584 4034 4642
rect 4434 4642 4448 4644
rect 4149 4584 4151 4604
rect 4155 4584 4157 4604
rect 4273 4584 4275 4624
rect 4279 4584 4281 4624
rect 4293 4584 4295 4624
rect 4299 4584 4305 4624
rect 4309 4584 4311 4624
rect 4446 4584 4448 4642
rect 4452 4584 4456 4644
rect 4460 4584 4464 4644
rect 4468 4584 4470 4644
rect 4550 4584 4552 4644
rect 4556 4584 4560 4644
rect 4564 4584 4568 4644
rect 4572 4642 4586 4644
rect 4572 4584 4574 4642
rect 4689 4584 4691 4604
rect 4695 4584 4697 4604
rect 4749 4584 4751 4624
rect 4755 4604 4768 4624
rect 5694 4642 5708 4644
rect 4931 4604 4941 4624
rect 4755 4584 4759 4604
rect 4771 4584 4773 4604
rect 4777 4584 4783 4604
rect 4787 4584 4789 4604
rect 4801 4584 4803 4604
rect 4807 4584 4811 4604
rect 4815 4584 4817 4604
rect 4855 4584 4857 4604
rect 4861 4584 4865 4604
rect 4877 4584 4879 4604
rect 4883 4584 4889 4604
rect 4893 4584 4895 4604
rect 4907 4584 4911 4604
rect 4915 4584 4921 4604
rect 4925 4584 4927 4604
rect 4939 4584 4941 4604
rect 4945 4584 4947 4624
rect 5029 4584 5031 4624
rect 5035 4612 5051 4624
rect 5035 4584 5037 4612
rect 5049 4584 5051 4612
rect 5055 4584 5057 4624
rect 5069 4584 5071 4624
rect 5075 4584 5077 4624
rect 5171 4584 5173 4624
rect 5177 4584 5183 4624
rect 5187 4584 5189 4624
rect 5291 4584 5293 4624
rect 5297 4584 5303 4624
rect 5307 4584 5309 4624
rect 5431 4584 5433 4624
rect 5437 4584 5443 4624
rect 5447 4584 5449 4624
rect 5551 4584 5553 4624
rect 5557 4584 5563 4624
rect 5567 4584 5569 4624
rect 5706 4584 5708 4642
rect 5712 4584 5716 4644
rect 5720 4584 5724 4644
rect 5728 4584 5730 4644
rect 83 4516 85 4556
rect 89 4516 91 4556
rect 103 4516 105 4556
rect 109 4528 111 4556
rect 123 4528 125 4556
rect 109 4516 125 4528
rect 129 4516 131 4556
rect 246 4498 248 4556
rect 234 4496 248 4498
rect 252 4496 256 4556
rect 260 4496 264 4556
rect 268 4496 270 4556
rect 352 4516 354 4556
rect 358 4516 362 4556
rect 366 4516 368 4556
rect 380 4536 384 4556
rect 388 4536 390 4556
rect 523 4516 525 4556
rect 529 4516 531 4556
rect 543 4516 545 4556
rect 549 4528 551 4556
rect 563 4528 565 4556
rect 549 4516 565 4528
rect 569 4516 571 4556
rect 663 4516 665 4556
rect 669 4516 671 4556
rect 683 4516 685 4556
rect 689 4528 691 4556
rect 703 4528 705 4556
rect 689 4516 705 4528
rect 709 4516 711 4556
rect 789 4536 791 4556
rect 795 4536 797 4556
rect 892 4516 894 4556
rect 898 4516 902 4556
rect 906 4516 908 4556
rect 920 4536 924 4556
rect 928 4536 930 4556
rect 1043 4536 1045 4556
rect 1049 4536 1051 4556
rect 1166 4498 1168 4556
rect 1154 4496 1168 4498
rect 1172 4496 1176 4556
rect 1180 4496 1184 4556
rect 1188 4496 1190 4556
rect 1290 4536 1292 4556
rect 1296 4536 1300 4556
rect 1312 4516 1314 4556
rect 1318 4516 1322 4556
rect 1326 4516 1328 4556
rect 1423 4536 1425 4556
rect 1429 4536 1431 4556
rect 1509 4516 1511 4556
rect 1515 4528 1517 4556
rect 1529 4528 1531 4556
rect 1515 4516 1531 4528
rect 1535 4516 1537 4556
rect 1549 4516 1551 4556
rect 1555 4516 1557 4556
rect 1671 4516 1673 4556
rect 1677 4516 1683 4556
rect 1687 4516 1689 4556
rect 1806 4498 1808 4556
rect 1794 4496 1808 4498
rect 1812 4496 1816 4556
rect 1820 4496 1824 4556
rect 1828 4496 1830 4556
rect 1923 4536 1925 4556
rect 1929 4536 1931 4556
rect 1943 4536 1945 4556
rect 1949 4536 1951 4556
rect 2066 4498 2068 4556
rect 2054 4496 2068 4498
rect 2072 4496 2076 4556
rect 2080 4496 2084 4556
rect 2088 4496 2090 4556
rect 2226 4498 2228 4556
rect 2214 4496 2228 4498
rect 2232 4496 2236 4556
rect 2240 4496 2244 4556
rect 2248 4496 2250 4556
rect 2351 4516 2353 4556
rect 2357 4516 2363 4556
rect 2367 4516 2369 4556
rect 2486 4498 2488 4556
rect 2474 4496 2488 4498
rect 2492 4496 2496 4556
rect 2500 4496 2504 4556
rect 2508 4496 2510 4556
rect 2590 4496 2592 4556
rect 2596 4496 2600 4556
rect 2604 4496 2608 4556
rect 2612 4498 2614 4556
rect 2743 4536 2745 4556
rect 2749 4536 2751 4556
rect 2843 4536 2845 4556
rect 2849 4536 2851 4556
rect 2863 4536 2865 4556
rect 2869 4536 2871 4556
rect 2612 4496 2626 4498
rect 2986 4498 2988 4556
rect 2974 4496 2988 4498
rect 2992 4496 2996 4556
rect 3000 4496 3004 4556
rect 3008 4496 3010 4556
rect 3126 4498 3128 4556
rect 3114 4496 3128 4498
rect 3132 4496 3136 4556
rect 3140 4496 3144 4556
rect 3148 4496 3150 4556
rect 3229 4536 3231 4556
rect 3235 4536 3237 4556
rect 3329 4516 3331 4556
rect 3335 4528 3337 4556
rect 3349 4528 3351 4556
rect 3335 4516 3351 4528
rect 3355 4516 3357 4556
rect 3369 4516 3371 4556
rect 3375 4516 3377 4556
rect 3493 4516 3495 4556
rect 3499 4516 3501 4556
rect 3513 4516 3515 4556
rect 3519 4516 3525 4556
rect 3529 4516 3531 4556
rect 3631 4516 3633 4556
rect 3637 4516 3643 4556
rect 3647 4516 3649 4556
rect 3763 4516 3765 4556
rect 3769 4536 3771 4556
rect 3783 4536 3785 4556
rect 3789 4536 3791 4556
rect 3803 4536 3805 4556
rect 3809 4536 3811 4556
rect 3769 4516 3781 4536
rect 3891 4516 3893 4556
rect 3897 4516 3903 4556
rect 3907 4516 3909 4556
rect 4021 4516 4023 4556
rect 4027 4516 4029 4556
rect 4041 4536 4045 4556
rect 4049 4536 4051 4556
rect 4129 4516 4131 4556
rect 4135 4516 4141 4556
rect 4145 4516 4147 4556
rect 4159 4516 4161 4556
rect 4165 4516 4167 4556
rect 4291 4516 4293 4556
rect 4297 4516 4303 4556
rect 4307 4516 4309 4556
rect 4403 4516 4405 4556
rect 4409 4516 4411 4556
rect 4423 4516 4425 4556
rect 4429 4528 4431 4556
rect 4443 4528 4445 4556
rect 4429 4516 4445 4528
rect 4449 4516 4451 4556
rect 4531 4516 4533 4556
rect 4537 4516 4543 4556
rect 4547 4516 4549 4556
rect 4671 4516 4673 4556
rect 4677 4516 4683 4556
rect 4687 4516 4689 4556
rect 4769 4536 4771 4556
rect 4775 4536 4777 4556
rect 4871 4516 4873 4556
rect 4877 4516 4883 4556
rect 4887 4516 4889 4556
rect 4989 4516 4991 4556
rect 4995 4528 4997 4556
rect 5009 4528 5011 4556
rect 4995 4516 5011 4528
rect 5015 4516 5017 4556
rect 5029 4516 5031 4556
rect 5035 4516 5037 4556
rect 5089 4516 5091 4556
rect 5095 4536 5099 4556
rect 5111 4536 5113 4556
rect 5117 4536 5123 4556
rect 5127 4536 5129 4556
rect 5141 4536 5143 4556
rect 5147 4536 5151 4556
rect 5155 4536 5157 4556
rect 5195 4536 5197 4556
rect 5201 4536 5205 4556
rect 5217 4536 5219 4556
rect 5223 4536 5229 4556
rect 5233 4536 5235 4556
rect 5247 4536 5251 4556
rect 5255 4536 5261 4556
rect 5265 4536 5267 4556
rect 5279 4536 5281 4556
rect 5095 4516 5108 4536
rect 5271 4516 5281 4536
rect 5285 4516 5287 4556
rect 5369 4516 5371 4556
rect 5375 4528 5377 4556
rect 5389 4528 5391 4556
rect 5375 4516 5391 4528
rect 5395 4516 5397 4556
rect 5409 4516 5411 4556
rect 5415 4516 5417 4556
rect 5509 4536 5511 4556
rect 5515 4536 5517 4556
rect 5529 4536 5531 4556
rect 5535 4536 5537 4556
rect 5549 4536 5551 4556
rect 5539 4516 5551 4536
rect 5555 4516 5557 4556
rect 5663 4516 5665 4556
rect 5669 4516 5671 4556
rect 5683 4516 5685 4556
rect 5689 4528 5691 4556
rect 5703 4528 5705 4556
rect 5689 4516 5705 4528
rect 5709 4516 5711 4556
rect 414 4162 428 4164
rect 103 4104 105 4144
rect 109 4104 111 4144
rect 123 4104 125 4144
rect 129 4132 145 4144
rect 129 4104 131 4132
rect 143 4104 145 4132
rect 149 4104 151 4144
rect 243 4104 245 4144
rect 249 4104 251 4144
rect 263 4104 265 4144
rect 269 4132 285 4144
rect 269 4104 271 4132
rect 283 4104 285 4132
rect 289 4104 291 4144
rect 426 4104 428 4162
rect 432 4104 436 4164
rect 440 4104 444 4164
rect 448 4104 450 4164
rect 554 4162 568 4164
rect 566 4104 568 4162
rect 572 4104 576 4164
rect 580 4104 584 4164
rect 588 4104 590 4164
rect 683 4104 685 4144
rect 689 4124 701 4144
rect 689 4104 691 4124
rect 703 4104 705 4124
rect 709 4104 711 4124
rect 723 4104 725 4124
rect 729 4104 731 4124
rect 823 4104 825 4144
rect 829 4104 831 4144
rect 843 4104 845 4144
rect 849 4132 865 4144
rect 849 4104 851 4132
rect 863 4104 865 4132
rect 869 4104 871 4144
rect 1234 4162 1248 4164
rect 949 4104 951 4124
rect 955 4104 957 4124
rect 1070 4104 1072 4124
rect 1076 4104 1080 4124
rect 1092 4104 1094 4144
rect 1098 4104 1102 4144
rect 1106 4104 1108 4144
rect 1246 4104 1248 4162
rect 1252 4104 1256 4164
rect 1260 4104 1264 4164
rect 1268 4104 1270 4164
rect 1371 4104 1373 4144
rect 1377 4104 1383 4144
rect 1387 4104 1389 4144
rect 1491 4104 1493 4144
rect 1497 4104 1503 4144
rect 1507 4104 1509 4144
rect 1734 4162 1748 4164
rect 1603 4104 1605 4124
rect 1609 4104 1611 4124
rect 1623 4104 1625 4124
rect 1629 4104 1631 4124
rect 1746 4104 1748 4162
rect 1752 4104 1756 4164
rect 1760 4104 1764 4164
rect 1768 4104 1770 4164
rect 1874 4162 1888 4164
rect 1886 4104 1888 4162
rect 1892 4104 1896 4164
rect 1900 4104 1904 4164
rect 1908 4104 1910 4164
rect 1990 4104 1992 4164
rect 1996 4104 2000 4164
rect 2004 4104 2008 4164
rect 2012 4162 2026 4164
rect 2012 4104 2014 4162
rect 2130 4104 2132 4164
rect 2136 4104 2140 4164
rect 2144 4104 2148 4164
rect 2152 4162 2166 4164
rect 2152 4104 2154 4162
rect 2594 4162 2608 4164
rect 2283 4104 2285 4124
rect 2289 4104 2291 4124
rect 2303 4104 2305 4124
rect 2309 4104 2311 4124
rect 2423 4104 2425 4144
rect 2429 4104 2431 4144
rect 2443 4104 2445 4144
rect 2449 4132 2465 4144
rect 2449 4104 2451 4132
rect 2463 4104 2465 4132
rect 2469 4104 2471 4144
rect 2606 4104 2608 4162
rect 2612 4104 2616 4164
rect 2620 4104 2624 4164
rect 2628 4104 2630 4164
rect 2709 4104 2711 4124
rect 2715 4104 2717 4124
rect 2830 4104 2832 4164
rect 2836 4104 2840 4164
rect 2844 4104 2848 4164
rect 2852 4162 2866 4164
rect 2852 4104 2854 4162
rect 2971 4104 2973 4144
rect 2977 4104 2983 4144
rect 2987 4104 2989 4144
rect 3092 4104 3094 4144
rect 3098 4104 3102 4144
rect 3106 4104 3108 4144
rect 3120 4104 3124 4124
rect 3128 4104 3130 4124
rect 3232 4104 3234 4144
rect 3238 4104 3242 4144
rect 3246 4104 3248 4144
rect 3260 4104 3264 4124
rect 3268 4104 3270 4124
rect 3369 4104 3371 4144
rect 3375 4132 3391 4144
rect 3375 4104 3377 4132
rect 3389 4104 3391 4132
rect 3395 4104 3397 4144
rect 3409 4104 3411 4144
rect 3415 4104 3417 4144
rect 3529 4104 3531 4124
rect 3535 4104 3537 4124
rect 3630 4104 3632 4164
rect 3636 4104 3640 4164
rect 3644 4104 3648 4164
rect 3652 4162 3666 4164
rect 3652 4104 3654 4162
rect 3770 4104 3772 4164
rect 3776 4104 3780 4164
rect 3784 4104 3788 4164
rect 3792 4162 3806 4164
rect 3792 4104 3794 4162
rect 3931 4104 3933 4144
rect 3937 4104 3943 4144
rect 3947 4104 3949 4144
rect 4071 4104 4073 4144
rect 4077 4104 4083 4144
rect 4087 4104 4089 4144
rect 4191 4104 4193 4144
rect 4197 4104 4203 4144
rect 4207 4104 4209 4144
rect 4303 4104 4305 4144
rect 4309 4104 4311 4144
rect 4323 4104 4325 4144
rect 4329 4132 4345 4144
rect 4329 4104 4331 4132
rect 4343 4104 4345 4132
rect 4349 4104 4351 4144
rect 4459 4124 4471 4144
rect 4429 4104 4431 4124
rect 4435 4104 4437 4124
rect 4449 4104 4451 4124
rect 4455 4104 4457 4124
rect 4469 4104 4471 4124
rect 4475 4104 4477 4144
rect 4583 4104 4585 4144
rect 4589 4104 4591 4144
rect 4603 4104 4605 4144
rect 4609 4132 4625 4144
rect 4609 4104 4611 4132
rect 4623 4104 4625 4132
rect 4629 4104 4631 4144
rect 4729 4104 4731 4144
rect 4735 4132 4751 4144
rect 4735 4104 4737 4132
rect 4749 4104 4751 4132
rect 4755 4104 4757 4144
rect 4769 4104 4771 4144
rect 4775 4104 4777 4144
rect 4869 4104 4871 4124
rect 4875 4104 4877 4124
rect 4889 4104 4891 4124
rect 4895 4104 4897 4124
rect 4989 4104 4991 4124
rect 4995 4104 4997 4124
rect 5112 4104 5114 4144
rect 5118 4104 5122 4144
rect 5126 4104 5128 4144
rect 5140 4104 5144 4124
rect 5148 4104 5150 4124
rect 5249 4104 5251 4144
rect 5255 4132 5271 4144
rect 5255 4104 5257 4132
rect 5269 4104 5271 4132
rect 5275 4104 5277 4144
rect 5289 4104 5291 4144
rect 5295 4104 5297 4144
rect 5389 4104 5391 4124
rect 5395 4104 5397 4124
rect 5489 4104 5491 4144
rect 5495 4132 5511 4144
rect 5495 4104 5497 4132
rect 5509 4104 5511 4132
rect 5515 4104 5517 4144
rect 5529 4104 5531 4144
rect 5535 4104 5537 4144
rect 5593 4104 5595 4144
rect 5599 4124 5609 4144
rect 5772 4124 5785 4144
rect 5599 4104 5601 4124
rect 5613 4104 5615 4124
rect 5619 4104 5625 4124
rect 5629 4104 5633 4124
rect 5645 4104 5647 4124
rect 5651 4104 5657 4124
rect 5661 4104 5663 4124
rect 5675 4104 5679 4124
rect 5683 4104 5685 4124
rect 5723 4104 5725 4124
rect 5729 4104 5733 4124
rect 5737 4104 5739 4124
rect 5751 4104 5753 4124
rect 5757 4104 5763 4124
rect 5767 4104 5769 4124
rect 5781 4104 5785 4124
rect 5789 4104 5791 4144
rect 83 4056 85 4076
rect 89 4056 91 4076
rect 189 4036 191 4076
rect 195 4048 197 4076
rect 209 4048 211 4076
rect 195 4036 211 4048
rect 215 4036 217 4076
rect 229 4036 231 4076
rect 235 4036 237 4076
rect 343 4056 345 4076
rect 349 4056 351 4076
rect 452 4036 454 4076
rect 458 4036 462 4076
rect 466 4036 468 4076
rect 480 4056 484 4076
rect 488 4056 490 4076
rect 603 4056 605 4076
rect 609 4056 611 4076
rect 623 4056 625 4076
rect 629 4056 631 4076
rect 743 4056 745 4076
rect 749 4056 751 4076
rect 829 4036 831 4076
rect 835 4048 837 4076
rect 849 4048 851 4076
rect 835 4036 851 4048
rect 855 4036 857 4076
rect 869 4036 871 4076
rect 875 4036 877 4076
rect 969 4056 971 4076
rect 975 4056 977 4076
rect 1070 4016 1072 4076
rect 1076 4016 1080 4076
rect 1084 4016 1088 4076
rect 1092 4018 1094 4076
rect 1212 4036 1214 4076
rect 1218 4036 1222 4076
rect 1226 4036 1228 4076
rect 1240 4036 1242 4076
rect 1246 4036 1250 4076
rect 1254 4036 1256 4076
rect 1391 4036 1393 4076
rect 1397 4036 1403 4076
rect 1407 4036 1409 4076
rect 1523 4056 1525 4076
rect 1529 4056 1531 4076
rect 1623 4056 1625 4076
rect 1629 4056 1631 4076
rect 1643 4056 1645 4076
rect 1649 4056 1651 4076
rect 1743 4056 1745 4076
rect 1749 4056 1751 4076
rect 1092 4016 1106 4018
rect 1830 4016 1832 4076
rect 1836 4016 1840 4076
rect 1844 4016 1848 4076
rect 1852 4018 1854 4076
rect 1983 4036 1985 4076
rect 1989 4036 1991 4076
rect 2003 4036 2005 4076
rect 2009 4048 2011 4076
rect 2023 4048 2025 4076
rect 2009 4036 2025 4048
rect 2029 4036 2031 4076
rect 1852 4016 1866 4018
rect 2166 4018 2168 4076
rect 2154 4016 2168 4018
rect 2172 4016 2176 4076
rect 2180 4016 2184 4076
rect 2188 4016 2190 4076
rect 2270 4016 2272 4076
rect 2276 4016 2280 4076
rect 2284 4016 2288 4076
rect 2292 4018 2294 4076
rect 2423 4036 2425 4076
rect 2429 4036 2431 4076
rect 2443 4036 2445 4076
rect 2449 4048 2451 4076
rect 2463 4048 2465 4076
rect 2449 4036 2465 4048
rect 2469 4036 2471 4076
rect 2571 4036 2573 4076
rect 2577 4036 2583 4076
rect 2587 4036 2589 4076
rect 2671 4036 2673 4076
rect 2677 4036 2683 4076
rect 2687 4036 2689 4076
rect 2292 4016 2306 4018
rect 2790 4016 2792 4076
rect 2796 4016 2800 4076
rect 2804 4016 2808 4076
rect 2812 4018 2814 4076
rect 2812 4016 2826 4018
rect 2930 4016 2932 4076
rect 2936 4016 2940 4076
rect 2944 4016 2948 4076
rect 2952 4018 2954 4076
rect 3083 4056 3085 4076
rect 3089 4056 3091 4076
rect 2952 4016 2966 4018
rect 3206 4018 3208 4076
rect 3194 4016 3208 4018
rect 3212 4016 3216 4076
rect 3220 4016 3224 4076
rect 3228 4016 3230 4076
rect 3323 4056 3325 4076
rect 3329 4056 3331 4076
rect 3423 4036 3425 4076
rect 3429 4036 3431 4076
rect 3443 4036 3445 4076
rect 3449 4048 3451 4076
rect 3463 4048 3465 4076
rect 3449 4036 3465 4048
rect 3469 4036 3471 4076
rect 3551 4036 3553 4076
rect 3557 4036 3563 4076
rect 3567 4036 3569 4076
rect 3683 4036 3685 4076
rect 3689 4056 3691 4076
rect 3703 4056 3705 4076
rect 3709 4056 3711 4076
rect 3723 4056 3725 4076
rect 3729 4056 3731 4076
rect 3689 4036 3701 4056
rect 3831 4036 3833 4076
rect 3837 4036 3843 4076
rect 3847 4036 3849 4076
rect 3963 4036 3965 4076
rect 3969 4036 3971 4076
rect 3983 4036 3985 4076
rect 3989 4048 3991 4076
rect 4003 4048 4005 4076
rect 3989 4036 4005 4048
rect 4009 4036 4011 4076
rect 4110 4056 4112 4076
rect 4116 4056 4120 4076
rect 4132 4036 4134 4076
rect 4138 4036 4142 4076
rect 4146 4036 4148 4076
rect 4231 4036 4233 4076
rect 4237 4036 4243 4076
rect 4247 4036 4249 4076
rect 4349 4036 4351 4076
rect 4355 4048 4357 4076
rect 4369 4048 4371 4076
rect 4355 4036 4371 4048
rect 4375 4036 4377 4076
rect 4389 4036 4391 4076
rect 4395 4036 4397 4076
rect 4489 4036 4491 4076
rect 4495 4048 4497 4076
rect 4509 4048 4511 4076
rect 4495 4036 4511 4048
rect 4515 4036 4517 4076
rect 4529 4036 4531 4076
rect 4535 4036 4537 4076
rect 4629 4056 4631 4076
rect 4635 4056 4637 4076
rect 4649 4056 4651 4076
rect 4655 4056 4657 4076
rect 4669 4056 4671 4076
rect 4659 4036 4671 4056
rect 4675 4036 4677 4076
rect 4791 4036 4793 4076
rect 4797 4036 4803 4076
rect 4807 4036 4809 4076
rect 4890 4016 4892 4076
rect 4896 4016 4900 4076
rect 4904 4016 4908 4076
rect 4912 4018 4914 4076
rect 5029 4056 5031 4076
rect 5035 4056 5037 4076
rect 5143 4056 5145 4076
rect 5149 4056 5151 4076
rect 4912 4016 4926 4018
rect 5189 4036 5191 4076
rect 5195 4056 5199 4076
rect 5211 4056 5213 4076
rect 5217 4056 5223 4076
rect 5227 4056 5229 4076
rect 5241 4056 5243 4076
rect 5247 4056 5251 4076
rect 5255 4056 5257 4076
rect 5295 4056 5297 4076
rect 5301 4056 5305 4076
rect 5317 4056 5319 4076
rect 5323 4056 5329 4076
rect 5333 4056 5335 4076
rect 5347 4056 5351 4076
rect 5355 4056 5361 4076
rect 5365 4056 5367 4076
rect 5379 4056 5381 4076
rect 5195 4036 5208 4056
rect 5371 4036 5381 4056
rect 5385 4036 5387 4076
rect 5429 4036 5431 4076
rect 5435 4056 5439 4076
rect 5451 4056 5453 4076
rect 5457 4056 5463 4076
rect 5467 4056 5469 4076
rect 5481 4056 5483 4076
rect 5487 4056 5491 4076
rect 5495 4056 5497 4076
rect 5535 4056 5537 4076
rect 5541 4056 5545 4076
rect 5557 4056 5559 4076
rect 5563 4056 5569 4076
rect 5573 4056 5575 4076
rect 5587 4056 5591 4076
rect 5595 4056 5601 4076
rect 5605 4056 5607 4076
rect 5619 4056 5621 4076
rect 5435 4036 5448 4056
rect 5611 4036 5621 4056
rect 5625 4036 5627 4076
rect 5709 4036 5711 4076
rect 5715 4048 5717 4076
rect 5729 4048 5731 4076
rect 5715 4036 5731 4048
rect 5735 4036 5737 4076
rect 5749 4036 5751 4076
rect 5755 4036 5757 4076
rect 214 3682 228 3684
rect 91 3624 93 3664
rect 97 3624 103 3664
rect 107 3624 109 3664
rect 226 3624 228 3682
rect 232 3624 236 3684
rect 240 3624 244 3684
rect 248 3624 250 3684
rect 403 3624 405 3644
rect 409 3624 411 3644
rect 423 3624 425 3644
rect 429 3624 431 3644
rect 443 3624 445 3644
rect 449 3624 451 3644
rect 563 3624 565 3664
rect 569 3624 571 3664
rect 583 3624 585 3664
rect 589 3652 605 3664
rect 589 3624 591 3652
rect 603 3624 605 3652
rect 609 3624 611 3664
rect 711 3624 713 3664
rect 717 3624 723 3664
rect 727 3624 729 3664
rect 809 3624 811 3664
rect 815 3652 831 3664
rect 815 3624 817 3652
rect 829 3624 831 3652
rect 835 3624 837 3664
rect 849 3624 851 3664
rect 855 3624 857 3664
rect 1004 3624 1006 3664
rect 1010 3624 1014 3664
rect 1018 3624 1020 3664
rect 1032 3624 1034 3664
rect 1038 3624 1042 3664
rect 1046 3624 1048 3664
rect 1131 3624 1133 3664
rect 1137 3624 1143 3664
rect 1147 3624 1149 3664
rect 1250 3624 1252 3684
rect 1256 3624 1260 3684
rect 1264 3624 1268 3684
rect 1272 3682 1286 3684
rect 1272 3624 1274 3682
rect 1392 3624 1394 3664
rect 1398 3624 1402 3664
rect 1406 3624 1408 3664
rect 1420 3624 1424 3644
rect 1428 3624 1430 3644
rect 1529 3624 1531 3664
rect 1535 3652 1551 3664
rect 1535 3624 1537 3652
rect 1549 3624 1551 3652
rect 1555 3624 1557 3664
rect 1569 3624 1571 3664
rect 1575 3624 1577 3664
rect 1669 3624 1671 3644
rect 1675 3624 1677 3644
rect 1791 3624 1793 3664
rect 1797 3624 1803 3664
rect 1807 3624 1809 3664
rect 1891 3624 1893 3664
rect 1897 3624 1903 3664
rect 1907 3624 1909 3664
rect 2039 3644 2051 3664
rect 2009 3624 2011 3644
rect 2015 3624 2017 3644
rect 2029 3624 2031 3644
rect 2035 3624 2037 3644
rect 2049 3624 2051 3644
rect 2055 3624 2057 3664
rect 2151 3624 2153 3664
rect 2157 3624 2163 3664
rect 2167 3624 2169 3664
rect 2270 3624 2272 3684
rect 2276 3624 2280 3684
rect 2284 3624 2288 3684
rect 2292 3682 2306 3684
rect 2292 3624 2294 3682
rect 2423 3624 2425 3664
rect 2429 3624 2431 3664
rect 2443 3624 2445 3664
rect 2449 3652 2465 3664
rect 2449 3624 2451 3652
rect 2463 3624 2465 3652
rect 2469 3624 2471 3664
rect 2551 3624 2553 3664
rect 2557 3624 2563 3664
rect 2567 3624 2569 3664
rect 2669 3624 2671 3664
rect 2675 3652 2691 3664
rect 2675 3624 2677 3652
rect 2689 3624 2691 3652
rect 2695 3624 2697 3664
rect 2709 3624 2711 3664
rect 2715 3624 2717 3664
rect 2823 3624 2825 3644
rect 2829 3624 2831 3644
rect 2923 3624 2925 3664
rect 2929 3624 2931 3664
rect 2943 3624 2945 3664
rect 2949 3652 2965 3664
rect 2949 3624 2951 3652
rect 2963 3624 2965 3652
rect 2969 3624 2971 3664
rect 3051 3624 3053 3664
rect 3057 3624 3063 3664
rect 3067 3624 3069 3664
rect 3211 3624 3213 3664
rect 3217 3624 3223 3664
rect 3227 3624 3229 3664
rect 3323 3624 3325 3644
rect 3329 3624 3331 3644
rect 3410 3624 3412 3684
rect 3416 3624 3420 3684
rect 3424 3624 3428 3684
rect 3432 3682 3446 3684
rect 3432 3624 3434 3682
rect 3549 3624 3551 3644
rect 3555 3624 3557 3644
rect 3663 3624 3665 3644
rect 3669 3624 3671 3644
rect 3683 3624 3685 3644
rect 3689 3624 3691 3644
rect 3791 3624 3793 3664
rect 3797 3624 3803 3664
rect 3807 3624 3809 3664
rect 3909 3624 3911 3644
rect 3915 3624 3917 3644
rect 4023 3624 4025 3644
rect 4029 3624 4031 3644
rect 4069 3624 4071 3664
rect 4075 3644 4088 3664
rect 4251 3644 4261 3664
rect 4075 3624 4079 3644
rect 4091 3624 4093 3644
rect 4097 3624 4103 3644
rect 4107 3624 4109 3644
rect 4121 3624 4123 3644
rect 4127 3624 4131 3644
rect 4135 3624 4137 3644
rect 4175 3624 4177 3644
rect 4181 3624 4185 3644
rect 4197 3624 4199 3644
rect 4203 3624 4209 3644
rect 4213 3624 4215 3644
rect 4227 3624 4231 3644
rect 4235 3624 4241 3644
rect 4245 3624 4247 3644
rect 4259 3624 4261 3644
rect 4265 3624 4267 3664
rect 4363 3624 4365 3664
rect 4369 3636 4371 3664
rect 4383 3636 4385 3664
rect 4369 3624 4385 3636
rect 4389 3624 4391 3664
rect 4403 3624 4405 3664
rect 4409 3654 4425 3664
rect 4409 3624 4411 3654
rect 4423 3624 4425 3654
rect 4429 3624 4431 3664
rect 4511 3624 4513 3664
rect 4517 3624 4523 3664
rect 4527 3624 4529 3664
rect 4629 3624 4631 3644
rect 4635 3624 4637 3644
rect 4649 3624 4651 3644
rect 4655 3624 4657 3644
rect 4749 3624 4751 3664
rect 4755 3652 4771 3664
rect 4755 3624 4757 3652
rect 4769 3624 4771 3652
rect 4775 3624 4777 3664
rect 4789 3624 4791 3664
rect 4795 3624 4797 3664
rect 4889 3624 4891 3664
rect 4895 3624 4897 3664
rect 5031 3624 5033 3664
rect 5037 3624 5043 3664
rect 5047 3624 5049 3664
rect 5129 3624 5131 3644
rect 5135 3624 5137 3644
rect 5243 3624 5245 3664
rect 5249 3624 5251 3664
rect 5263 3624 5265 3664
rect 5269 3624 5271 3664
rect 5283 3624 5285 3664
rect 5289 3624 5291 3664
rect 5303 3624 5305 3664
rect 5309 3624 5311 3664
rect 5323 3624 5325 3664
rect 5329 3624 5331 3664
rect 5343 3624 5345 3664
rect 5349 3624 5351 3664
rect 5363 3624 5365 3664
rect 5369 3624 5371 3664
rect 5383 3624 5385 3664
rect 5389 3624 5391 3664
rect 5429 3624 5431 3664
rect 5435 3644 5448 3664
rect 5611 3644 5621 3664
rect 5435 3624 5439 3644
rect 5451 3624 5453 3644
rect 5457 3624 5463 3644
rect 5467 3624 5469 3644
rect 5481 3624 5483 3644
rect 5487 3624 5491 3644
rect 5495 3624 5497 3644
rect 5535 3624 5537 3644
rect 5541 3624 5545 3644
rect 5557 3624 5559 3644
rect 5563 3624 5569 3644
rect 5573 3624 5575 3644
rect 5587 3624 5591 3644
rect 5595 3624 5601 3644
rect 5605 3624 5607 3644
rect 5619 3624 5621 3644
rect 5625 3624 5627 3664
rect 5731 3624 5733 3664
rect 5737 3624 5743 3664
rect 5747 3624 5749 3664
rect 83 3556 85 3596
rect 89 3556 91 3596
rect 103 3556 105 3596
rect 109 3568 111 3596
rect 123 3568 125 3596
rect 109 3556 125 3568
rect 129 3556 131 3596
rect 212 3556 214 3596
rect 218 3556 222 3596
rect 226 3556 228 3596
rect 240 3576 244 3596
rect 248 3576 250 3596
rect 349 3576 351 3596
rect 355 3576 357 3596
rect 449 3556 451 3596
rect 455 3568 457 3596
rect 469 3568 471 3596
rect 455 3556 471 3568
rect 475 3556 477 3596
rect 489 3556 491 3596
rect 495 3556 497 3596
rect 590 3536 592 3596
rect 596 3536 600 3596
rect 604 3536 608 3596
rect 612 3538 614 3596
rect 771 3556 773 3596
rect 777 3556 783 3596
rect 787 3556 789 3596
rect 891 3556 893 3596
rect 897 3556 903 3596
rect 907 3556 909 3596
rect 989 3556 991 3596
rect 995 3568 997 3596
rect 1009 3568 1011 3596
rect 995 3556 1011 3568
rect 1015 3556 1017 3596
rect 1029 3556 1031 3596
rect 1035 3556 1037 3596
rect 612 3536 626 3538
rect 1166 3538 1168 3596
rect 1154 3536 1168 3538
rect 1172 3536 1176 3596
rect 1180 3536 1184 3596
rect 1188 3536 1190 3596
rect 1271 3556 1273 3596
rect 1277 3556 1283 3596
rect 1287 3556 1289 3596
rect 1426 3538 1428 3596
rect 1414 3536 1428 3538
rect 1432 3536 1436 3596
rect 1440 3536 1444 3596
rect 1448 3536 1450 3596
rect 1529 3556 1531 3596
rect 1535 3568 1537 3596
rect 1549 3568 1551 3596
rect 1535 3556 1551 3568
rect 1555 3556 1557 3596
rect 1569 3556 1571 3596
rect 1575 3556 1577 3596
rect 1690 3576 1692 3596
rect 1696 3576 1700 3596
rect 1712 3556 1714 3596
rect 1718 3556 1722 3596
rect 1726 3556 1728 3596
rect 1846 3538 1848 3596
rect 1834 3536 1848 3538
rect 1852 3536 1856 3596
rect 1860 3536 1864 3596
rect 1868 3536 1870 3596
rect 1952 3556 1954 3596
rect 1958 3556 1962 3596
rect 1966 3556 1968 3596
rect 1980 3576 1984 3596
rect 1988 3576 1990 3596
rect 2103 3556 2105 3596
rect 2109 3556 2111 3596
rect 2123 3556 2125 3596
rect 2129 3568 2131 3596
rect 2143 3568 2145 3596
rect 2129 3556 2145 3568
rect 2149 3556 2151 3596
rect 2249 3556 2251 3596
rect 2255 3568 2257 3596
rect 2269 3568 2271 3596
rect 2255 3556 2271 3568
rect 2275 3556 2277 3596
rect 2289 3556 2291 3596
rect 2295 3556 2297 3596
rect 2410 3576 2412 3596
rect 2416 3576 2420 3596
rect 2432 3556 2434 3596
rect 2438 3556 2442 3596
rect 2446 3556 2448 3596
rect 2553 3556 2555 3596
rect 2559 3556 2561 3596
rect 2573 3556 2575 3596
rect 2579 3556 2585 3596
rect 2589 3556 2591 3596
rect 2671 3556 2673 3596
rect 2677 3556 2683 3596
rect 2687 3556 2689 3596
rect 2803 3556 2805 3596
rect 2809 3556 2811 3596
rect 2823 3556 2825 3596
rect 2829 3568 2831 3596
rect 2843 3568 2845 3596
rect 2829 3556 2845 3568
rect 2849 3556 2851 3596
rect 2961 3556 2963 3596
rect 2967 3556 2969 3596
rect 2981 3576 2985 3596
rect 2989 3576 2991 3596
rect 3091 3556 3093 3596
rect 3097 3556 3103 3596
rect 3107 3556 3109 3596
rect 3190 3536 3192 3596
rect 3196 3536 3200 3596
rect 3204 3536 3208 3596
rect 3212 3538 3214 3596
rect 3212 3536 3226 3538
rect 3366 3538 3368 3596
rect 3354 3536 3368 3538
rect 3372 3536 3376 3596
rect 3380 3536 3384 3596
rect 3388 3536 3390 3596
rect 3483 3556 3485 3596
rect 3489 3556 3491 3596
rect 3503 3556 3505 3596
rect 3509 3568 3511 3596
rect 3523 3568 3525 3596
rect 3509 3556 3525 3568
rect 3529 3556 3531 3596
rect 3623 3556 3625 3596
rect 3629 3556 3631 3596
rect 3643 3556 3645 3596
rect 3649 3568 3651 3596
rect 3663 3568 3665 3596
rect 3649 3556 3665 3568
rect 3669 3556 3671 3596
rect 3773 3556 3775 3596
rect 3779 3556 3781 3596
rect 3793 3556 3795 3596
rect 3799 3556 3805 3596
rect 3809 3556 3811 3596
rect 3889 3576 3891 3596
rect 3895 3576 3897 3596
rect 3909 3576 3911 3596
rect 3915 3576 3917 3596
rect 4043 3556 4045 3596
rect 4049 3556 4051 3596
rect 4063 3556 4065 3596
rect 4069 3568 4071 3596
rect 4083 3568 4085 3596
rect 4069 3556 4085 3568
rect 4089 3556 4091 3596
rect 4169 3576 4171 3596
rect 4175 3576 4177 3596
rect 4269 3556 4271 3596
rect 4275 3568 4277 3596
rect 4289 3568 4291 3596
rect 4275 3556 4291 3568
rect 4295 3556 4297 3596
rect 4309 3556 4311 3596
rect 4315 3556 4317 3596
rect 4431 3556 4433 3596
rect 4437 3556 4443 3596
rect 4447 3556 4449 3596
rect 4531 3556 4533 3596
rect 4537 3556 4543 3596
rect 4547 3556 4549 3596
rect 4609 3556 4611 3596
rect 4615 3576 4619 3596
rect 4631 3576 4633 3596
rect 4637 3576 4643 3596
rect 4647 3576 4649 3596
rect 4661 3576 4663 3596
rect 4667 3576 4671 3596
rect 4675 3576 4677 3596
rect 4715 3576 4717 3596
rect 4721 3576 4725 3596
rect 4737 3576 4739 3596
rect 4743 3576 4749 3596
rect 4753 3576 4755 3596
rect 4767 3576 4771 3596
rect 4775 3576 4781 3596
rect 4785 3576 4787 3596
rect 4799 3576 4801 3596
rect 4615 3556 4628 3576
rect 4791 3556 4801 3576
rect 4805 3556 4807 3596
rect 4911 3556 4913 3596
rect 4917 3556 4923 3596
rect 4927 3556 4929 3596
rect 5023 3556 5025 3596
rect 5029 3556 5031 3596
rect 5043 3556 5045 3596
rect 5049 3568 5051 3596
rect 5063 3568 5065 3596
rect 5049 3556 5065 3568
rect 5069 3556 5071 3596
rect 5171 3556 5173 3596
rect 5177 3556 5183 3596
rect 5187 3556 5189 3596
rect 5253 3556 5255 3596
rect 5259 3576 5261 3596
rect 5273 3576 5275 3596
rect 5279 3576 5285 3596
rect 5289 3576 5293 3596
rect 5305 3576 5307 3596
rect 5311 3576 5317 3596
rect 5321 3576 5323 3596
rect 5335 3576 5339 3596
rect 5343 3576 5345 3596
rect 5383 3576 5385 3596
rect 5389 3576 5393 3596
rect 5397 3576 5399 3596
rect 5411 3576 5413 3596
rect 5417 3576 5423 3596
rect 5427 3576 5429 3596
rect 5441 3576 5445 3596
rect 5259 3556 5269 3576
rect 5432 3556 5445 3576
rect 5449 3556 5451 3596
rect 5551 3556 5553 3596
rect 5557 3556 5563 3596
rect 5567 3556 5569 3596
rect 5649 3556 5651 3596
rect 5655 3568 5657 3596
rect 5669 3568 5671 3596
rect 5655 3556 5671 3568
rect 5675 3556 5677 3596
rect 5689 3556 5691 3596
rect 5695 3556 5697 3596
rect 83 3144 85 3164
rect 89 3144 91 3164
rect 183 3144 185 3184
rect 189 3144 191 3184
rect 203 3144 205 3184
rect 209 3172 225 3184
rect 209 3144 211 3172
rect 223 3144 225 3172
rect 229 3144 231 3184
rect 323 3144 325 3164
rect 329 3144 331 3164
rect 411 3144 413 3184
rect 417 3144 423 3184
rect 427 3144 429 3184
rect 532 3144 534 3184
rect 538 3144 542 3184
rect 546 3144 548 3184
rect 974 3202 988 3204
rect 560 3144 564 3164
rect 568 3144 570 3164
rect 669 3144 671 3184
rect 675 3144 681 3184
rect 685 3144 687 3184
rect 699 3144 701 3184
rect 705 3144 707 3184
rect 851 3144 853 3184
rect 857 3144 863 3184
rect 867 3144 869 3184
rect 986 3144 988 3202
rect 992 3144 996 3204
rect 1000 3144 1004 3204
rect 1008 3144 1010 3204
rect 1114 3202 1128 3204
rect 1126 3144 1128 3202
rect 1132 3144 1136 3204
rect 1140 3144 1144 3204
rect 1148 3144 1150 3204
rect 1232 3144 1234 3184
rect 1238 3144 1242 3184
rect 1246 3144 1248 3184
rect 1494 3202 1508 3204
rect 1260 3144 1264 3164
rect 1268 3144 1270 3164
rect 1383 3144 1385 3164
rect 1389 3144 1391 3164
rect 1506 3144 1508 3202
rect 1512 3144 1516 3204
rect 1520 3144 1524 3204
rect 1528 3144 1530 3204
rect 1634 3202 1648 3204
rect 1646 3144 1648 3202
rect 1652 3144 1656 3204
rect 1660 3144 1664 3204
rect 1668 3144 1670 3204
rect 1770 3144 1772 3164
rect 1776 3144 1780 3164
rect 1792 3144 1794 3184
rect 1798 3144 1802 3184
rect 1806 3144 1808 3184
rect 1931 3144 1933 3184
rect 1937 3144 1943 3184
rect 1947 3144 1949 3184
rect 2050 3144 2052 3164
rect 2056 3144 2060 3164
rect 2072 3144 2074 3184
rect 2078 3144 2082 3184
rect 2086 3144 2088 3184
rect 2171 3144 2173 3184
rect 2177 3144 2183 3184
rect 2187 3144 2189 3184
rect 2313 3144 2315 3184
rect 2319 3144 2321 3184
rect 2333 3144 2335 3184
rect 2339 3144 2345 3184
rect 2349 3144 2351 3184
rect 2431 3144 2433 3184
rect 2437 3144 2443 3184
rect 2447 3144 2449 3184
rect 2563 3144 2565 3184
rect 2569 3144 2571 3184
rect 2583 3144 2585 3184
rect 2589 3172 2605 3184
rect 2589 3144 2591 3172
rect 2603 3144 2605 3172
rect 2609 3144 2611 3184
rect 2710 3144 2712 3164
rect 2716 3144 2720 3164
rect 2732 3144 2734 3184
rect 2738 3144 2742 3184
rect 2746 3144 2748 3184
rect 2830 3144 2832 3204
rect 2836 3144 2840 3204
rect 2844 3144 2848 3204
rect 2852 3202 2866 3204
rect 2852 3144 2854 3202
rect 2970 3144 2972 3204
rect 2976 3144 2980 3204
rect 2984 3144 2988 3204
rect 2992 3202 3006 3204
rect 2992 3144 2994 3202
rect 3131 3144 3133 3184
rect 3137 3144 3143 3184
rect 3147 3144 3149 3184
rect 3271 3144 3273 3184
rect 3277 3144 3283 3184
rect 3287 3144 3289 3184
rect 3494 3202 3508 3204
rect 3369 3144 3371 3164
rect 3375 3144 3377 3164
rect 3506 3144 3508 3202
rect 3512 3144 3516 3204
rect 3520 3144 3524 3204
rect 3528 3144 3530 3204
rect 3612 3144 3614 3184
rect 3618 3144 3622 3184
rect 3626 3144 3628 3184
rect 3640 3144 3644 3164
rect 3648 3144 3650 3164
rect 3763 3144 3765 3184
rect 3769 3144 3771 3184
rect 3783 3144 3785 3184
rect 3789 3172 3805 3184
rect 3789 3144 3791 3172
rect 3803 3144 3805 3172
rect 3809 3144 3811 3184
rect 3889 3144 3891 3164
rect 3895 3144 3897 3164
rect 3949 3144 3951 3184
rect 3955 3164 3968 3184
rect 4131 3164 4141 3184
rect 3955 3144 3959 3164
rect 3971 3144 3973 3164
rect 3977 3144 3983 3164
rect 3987 3144 3989 3164
rect 4001 3144 4003 3164
rect 4007 3144 4011 3164
rect 4015 3144 4017 3164
rect 4055 3144 4057 3164
rect 4061 3144 4065 3164
rect 4077 3144 4079 3164
rect 4083 3144 4089 3164
rect 4093 3144 4095 3164
rect 4107 3144 4111 3164
rect 4115 3144 4121 3164
rect 4125 3144 4127 3164
rect 4139 3144 4141 3164
rect 4145 3144 4147 3184
rect 4229 3144 4231 3184
rect 4235 3172 4251 3184
rect 4235 3144 4237 3172
rect 4249 3144 4251 3172
rect 4255 3144 4257 3184
rect 4269 3144 4271 3184
rect 4275 3144 4277 3184
rect 4369 3144 4371 3184
rect 4375 3172 4391 3184
rect 4375 3144 4377 3172
rect 4389 3144 4391 3172
rect 4395 3144 4397 3184
rect 4409 3144 4411 3184
rect 4415 3144 4417 3184
rect 4469 3144 4471 3184
rect 4475 3164 4488 3184
rect 4651 3164 4661 3184
rect 4475 3144 4479 3164
rect 4491 3144 4493 3164
rect 4497 3144 4503 3164
rect 4507 3144 4509 3164
rect 4521 3144 4523 3164
rect 4527 3144 4531 3164
rect 4535 3144 4537 3164
rect 4575 3144 4577 3164
rect 4581 3144 4585 3164
rect 4597 3144 4599 3164
rect 4603 3144 4609 3164
rect 4613 3144 4615 3164
rect 4627 3144 4631 3164
rect 4635 3144 4641 3164
rect 4645 3144 4647 3164
rect 4659 3144 4661 3164
rect 4665 3144 4667 3184
rect 4749 3144 4751 3184
rect 4755 3172 4771 3184
rect 4755 3144 4757 3172
rect 4769 3144 4771 3172
rect 4775 3144 4777 3184
rect 4789 3144 4791 3184
rect 4795 3144 4797 3184
rect 4911 3144 4913 3184
rect 4917 3144 4923 3184
rect 4927 3144 4929 3184
rect 5023 3144 5025 3184
rect 5029 3144 5031 3184
rect 5043 3144 5045 3184
rect 5049 3172 5065 3184
rect 5049 3144 5051 3172
rect 5063 3144 5065 3172
rect 5069 3144 5071 3184
rect 5163 3144 5165 3164
rect 5169 3144 5171 3164
rect 5271 3144 5273 3184
rect 5277 3144 5283 3184
rect 5287 3144 5289 3184
rect 5369 3144 5371 3164
rect 5375 3144 5377 3164
rect 5489 3144 5491 3184
rect 5495 3172 5511 3184
rect 5495 3144 5497 3172
rect 5509 3144 5511 3172
rect 5515 3144 5517 3184
rect 5529 3144 5531 3184
rect 5535 3144 5537 3184
rect 5671 3144 5673 3184
rect 5677 3144 5683 3184
rect 5687 3144 5689 3184
rect 113 3076 115 3116
rect 119 3076 121 3116
rect 133 3076 135 3116
rect 139 3076 145 3116
rect 149 3076 151 3116
rect 250 3056 252 3116
rect 256 3056 260 3116
rect 264 3056 268 3116
rect 272 3058 274 3116
rect 391 3076 393 3116
rect 397 3076 403 3116
rect 407 3076 409 3116
rect 523 3076 525 3116
rect 529 3076 531 3116
rect 543 3076 545 3116
rect 549 3088 551 3116
rect 563 3088 565 3116
rect 549 3076 565 3088
rect 569 3076 571 3116
rect 649 3076 651 3116
rect 655 3088 657 3116
rect 669 3088 671 3116
rect 655 3076 671 3088
rect 675 3076 677 3116
rect 689 3076 691 3116
rect 695 3076 697 3116
rect 789 3076 791 3116
rect 795 3088 797 3116
rect 809 3088 811 3116
rect 795 3076 811 3088
rect 815 3076 817 3116
rect 829 3076 831 3116
rect 835 3076 837 3116
rect 929 3076 931 3116
rect 935 3088 937 3116
rect 949 3088 951 3116
rect 935 3076 951 3088
rect 955 3076 957 3116
rect 969 3076 971 3116
rect 975 3076 977 3116
rect 1091 3076 1093 3116
rect 1097 3076 1103 3116
rect 1107 3076 1109 3116
rect 1223 3096 1225 3116
rect 1229 3096 1231 3116
rect 1243 3096 1245 3116
rect 1249 3096 1251 3116
rect 272 3056 286 3058
rect 1329 3076 1331 3116
rect 1335 3088 1337 3116
rect 1349 3088 1351 3116
rect 1335 3076 1351 3088
rect 1355 3076 1357 3116
rect 1369 3076 1371 3116
rect 1375 3076 1377 3116
rect 1506 3058 1508 3116
rect 1494 3056 1508 3058
rect 1512 3056 1516 3116
rect 1520 3056 1524 3116
rect 1528 3056 1530 3116
rect 1650 3096 1652 3116
rect 1656 3096 1660 3116
rect 1672 3076 1674 3116
rect 1678 3076 1682 3116
rect 1686 3076 1688 3116
rect 1783 3076 1785 3116
rect 1789 3076 1791 3116
rect 1803 3076 1805 3116
rect 1809 3088 1811 3116
rect 1823 3088 1825 3116
rect 1809 3076 1825 3088
rect 1829 3076 1831 3116
rect 1909 3076 1911 3116
rect 1915 3088 1917 3116
rect 1929 3088 1931 3116
rect 1915 3076 1931 3088
rect 1935 3076 1937 3116
rect 1949 3076 1951 3116
rect 1955 3076 1957 3116
rect 2083 3076 2085 3116
rect 2089 3076 2091 3116
rect 2103 3076 2105 3116
rect 2109 3088 2111 3116
rect 2123 3088 2125 3116
rect 2109 3076 2125 3088
rect 2129 3076 2131 3116
rect 2223 3076 2225 3116
rect 2229 3076 2231 3116
rect 2243 3076 2245 3116
rect 2249 3088 2251 3116
rect 2263 3088 2265 3116
rect 2249 3076 2265 3088
rect 2269 3076 2271 3116
rect 2390 3096 2392 3116
rect 2396 3096 2400 3116
rect 2412 3076 2414 3116
rect 2418 3076 2422 3116
rect 2426 3076 2428 3116
rect 2530 3096 2532 3116
rect 2536 3096 2540 3116
rect 2552 3076 2554 3116
rect 2558 3076 2562 3116
rect 2566 3076 2568 3116
rect 2684 3076 2686 3116
rect 2690 3076 2694 3116
rect 2698 3076 2700 3116
rect 2712 3076 2714 3116
rect 2718 3076 2722 3116
rect 2726 3076 2728 3116
rect 2823 3076 2825 3116
rect 2829 3096 2831 3116
rect 2843 3096 2845 3116
rect 2849 3096 2851 3116
rect 2863 3096 2865 3116
rect 2869 3096 2871 3116
rect 2949 3096 2951 3116
rect 2955 3096 2957 3116
rect 2969 3096 2971 3116
rect 2975 3096 2977 3116
rect 2829 3076 2841 3096
rect 3091 3076 3093 3116
rect 3097 3076 3103 3116
rect 3107 3076 3109 3116
rect 3233 3076 3235 3116
rect 3239 3076 3241 3116
rect 3253 3076 3255 3116
rect 3259 3076 3265 3116
rect 3269 3076 3271 3116
rect 3349 3096 3351 3116
rect 3355 3096 3357 3116
rect 3369 3096 3371 3116
rect 3375 3096 3377 3116
rect 3389 3096 3391 3116
rect 3379 3076 3391 3096
rect 3395 3076 3397 3116
rect 3503 3076 3505 3116
rect 3509 3076 3511 3116
rect 3523 3076 3525 3116
rect 3529 3088 3531 3116
rect 3543 3088 3545 3116
rect 3529 3076 3545 3088
rect 3549 3076 3551 3116
rect 3643 3076 3645 3116
rect 3649 3076 3651 3116
rect 3663 3076 3665 3116
rect 3669 3088 3671 3116
rect 3683 3088 3685 3116
rect 3669 3076 3685 3088
rect 3689 3076 3691 3116
rect 3783 3076 3785 3116
rect 3789 3096 3791 3116
rect 3803 3096 3805 3116
rect 3809 3096 3811 3116
rect 3823 3096 3825 3116
rect 3829 3096 3831 3116
rect 3789 3076 3801 3096
rect 3953 3076 3955 3116
rect 3959 3076 3961 3116
rect 3973 3076 3975 3116
rect 3979 3076 3985 3116
rect 3989 3076 3991 3116
rect 4069 3096 4071 3116
rect 4075 3096 4077 3116
rect 4089 3096 4091 3116
rect 4095 3096 4097 3116
rect 4190 3056 4192 3116
rect 4196 3056 4200 3116
rect 4204 3056 4208 3116
rect 4212 3058 4214 3116
rect 4293 3076 4295 3116
rect 4299 3096 4301 3116
rect 4313 3096 4315 3116
rect 4319 3096 4325 3116
rect 4329 3096 4333 3116
rect 4345 3096 4347 3116
rect 4351 3096 4357 3116
rect 4361 3096 4363 3116
rect 4375 3096 4379 3116
rect 4383 3096 4385 3116
rect 4423 3096 4425 3116
rect 4429 3096 4433 3116
rect 4437 3096 4439 3116
rect 4451 3096 4453 3116
rect 4457 3096 4463 3116
rect 4467 3096 4469 3116
rect 4481 3096 4485 3116
rect 4299 3076 4309 3096
rect 4212 3056 4226 3058
rect 4472 3076 4485 3096
rect 4489 3076 4491 3116
rect 4589 3076 4591 3116
rect 4595 3088 4597 3116
rect 4609 3088 4611 3116
rect 4595 3076 4611 3088
rect 4615 3076 4617 3116
rect 4629 3076 4631 3116
rect 4635 3076 4637 3116
rect 4729 3076 4731 3116
rect 4735 3088 4737 3116
rect 4749 3088 4751 3116
rect 4735 3076 4751 3088
rect 4755 3076 4757 3116
rect 4769 3076 4771 3116
rect 4775 3076 4777 3116
rect 4891 3076 4893 3116
rect 4897 3076 4903 3116
rect 4907 3076 4909 3116
rect 4991 3076 4993 3116
rect 4997 3076 5003 3116
rect 5007 3076 5009 3116
rect 5073 3076 5075 3116
rect 5079 3096 5081 3116
rect 5093 3096 5095 3116
rect 5099 3096 5105 3116
rect 5109 3096 5113 3116
rect 5125 3096 5127 3116
rect 5131 3096 5137 3116
rect 5141 3096 5143 3116
rect 5155 3096 5159 3116
rect 5163 3096 5165 3116
rect 5203 3096 5205 3116
rect 5209 3096 5213 3116
rect 5217 3096 5219 3116
rect 5231 3096 5233 3116
rect 5237 3096 5243 3116
rect 5247 3096 5249 3116
rect 5261 3096 5265 3116
rect 5079 3076 5089 3096
rect 5252 3076 5265 3096
rect 5269 3076 5271 3116
rect 5363 3076 5365 3116
rect 5369 3076 5371 3116
rect 5383 3076 5385 3116
rect 5389 3076 5391 3116
rect 5403 3076 5405 3116
rect 5409 3076 5411 3116
rect 5423 3076 5425 3116
rect 5429 3076 5431 3116
rect 5443 3076 5445 3116
rect 5449 3076 5451 3116
rect 5463 3076 5465 3116
rect 5469 3076 5471 3116
rect 5483 3076 5485 3116
rect 5489 3076 5491 3116
rect 5503 3076 5505 3116
rect 5509 3076 5511 3116
rect 5549 3076 5551 3116
rect 5555 3096 5559 3116
rect 5571 3096 5573 3116
rect 5577 3096 5583 3116
rect 5587 3096 5589 3116
rect 5601 3096 5603 3116
rect 5607 3096 5611 3116
rect 5615 3096 5617 3116
rect 5655 3096 5657 3116
rect 5661 3096 5665 3116
rect 5677 3096 5679 3116
rect 5683 3096 5689 3116
rect 5693 3096 5695 3116
rect 5707 3096 5711 3116
rect 5715 3096 5721 3116
rect 5725 3096 5727 3116
rect 5739 3096 5741 3116
rect 5555 3076 5568 3096
rect 5731 3076 5741 3096
rect 5745 3076 5747 3116
rect 91 2664 93 2704
rect 97 2664 103 2704
rect 107 2664 109 2704
rect 189 2664 191 2704
rect 195 2692 211 2704
rect 195 2664 197 2692
rect 209 2664 211 2692
rect 215 2664 217 2704
rect 229 2664 231 2704
rect 235 2664 237 2704
rect 343 2664 345 2684
rect 349 2664 351 2684
rect 432 2664 434 2704
rect 438 2664 442 2704
rect 446 2664 448 2704
rect 460 2664 464 2684
rect 468 2664 470 2684
rect 591 2664 593 2704
rect 597 2664 603 2704
rect 607 2664 609 2704
rect 689 2664 691 2704
rect 695 2664 701 2704
rect 705 2664 707 2704
rect 719 2664 721 2704
rect 725 2664 727 2704
rect 831 2664 833 2704
rect 837 2664 843 2704
rect 847 2664 849 2704
rect 952 2664 954 2704
rect 958 2664 962 2704
rect 966 2664 968 2704
rect 980 2664 984 2684
rect 988 2664 990 2684
rect 1091 2664 1093 2704
rect 1097 2664 1103 2704
rect 1107 2664 1109 2704
rect 1243 2664 1245 2704
rect 1249 2664 1251 2704
rect 1263 2664 1265 2704
rect 1269 2692 1285 2704
rect 1269 2664 1271 2692
rect 1283 2664 1285 2692
rect 1289 2664 1291 2704
rect 1369 2664 1371 2704
rect 1375 2692 1391 2704
rect 1375 2664 1377 2692
rect 1389 2664 1391 2692
rect 1395 2664 1397 2704
rect 1409 2664 1411 2704
rect 1415 2664 1417 2704
rect 1523 2664 1525 2704
rect 1529 2684 1541 2704
rect 1529 2664 1531 2684
rect 1543 2664 1545 2684
rect 1549 2664 1551 2684
rect 1563 2664 1565 2684
rect 1569 2664 1571 2684
rect 1649 2664 1651 2684
rect 1655 2664 1657 2684
rect 1669 2664 1671 2684
rect 1675 2664 1677 2684
rect 1793 2664 1795 2704
rect 1799 2664 1801 2704
rect 1813 2664 1815 2704
rect 1819 2664 1825 2704
rect 1829 2664 1831 2704
rect 1951 2664 1953 2704
rect 1957 2664 1963 2704
rect 1967 2664 1969 2704
rect 2049 2664 2051 2704
rect 2055 2692 2071 2704
rect 2055 2664 2057 2692
rect 2069 2664 2071 2692
rect 2075 2664 2077 2704
rect 2089 2664 2091 2704
rect 2095 2664 2097 2704
rect 2213 2664 2215 2704
rect 2219 2664 2221 2704
rect 2233 2664 2235 2704
rect 2239 2664 2245 2704
rect 2249 2664 2251 2704
rect 2351 2664 2353 2704
rect 2357 2664 2363 2704
rect 2367 2664 2369 2704
rect 2614 2722 2628 2724
rect 2469 2664 2471 2684
rect 2475 2664 2477 2684
rect 2489 2664 2491 2684
rect 2495 2664 2497 2684
rect 2626 2664 2628 2722
rect 2632 2664 2636 2724
rect 2640 2664 2644 2724
rect 2648 2664 2650 2724
rect 3054 2722 3068 2724
rect 2753 2664 2755 2704
rect 2759 2664 2761 2704
rect 2773 2664 2775 2704
rect 2779 2664 2785 2704
rect 2789 2664 2791 2704
rect 2889 2664 2891 2704
rect 2895 2692 2911 2704
rect 2895 2664 2897 2692
rect 2909 2664 2911 2692
rect 2915 2664 2917 2704
rect 2929 2664 2931 2704
rect 2935 2664 2937 2704
rect 3066 2664 3068 2722
rect 3072 2664 3076 2724
rect 3080 2664 3084 2724
rect 3088 2664 3090 2724
rect 3171 2664 3173 2704
rect 3177 2664 3183 2704
rect 3187 2664 3189 2704
rect 3303 2664 3305 2704
rect 3309 2664 3311 2704
rect 3323 2664 3325 2704
rect 3329 2692 3345 2704
rect 3329 2664 3331 2692
rect 3343 2664 3345 2692
rect 3349 2664 3351 2704
rect 3453 2664 3455 2704
rect 3459 2664 3461 2704
rect 3473 2664 3475 2704
rect 3479 2664 3485 2704
rect 3489 2664 3491 2704
rect 3569 2664 3571 2684
rect 3575 2664 3577 2684
rect 3589 2664 3591 2684
rect 3595 2664 3597 2684
rect 3690 2664 3692 2724
rect 3696 2664 3700 2724
rect 3704 2664 3708 2724
rect 3712 2722 3726 2724
rect 3712 2664 3714 2722
rect 3831 2664 3833 2704
rect 3837 2664 3843 2704
rect 3847 2664 3849 2704
rect 3963 2664 3965 2704
rect 3969 2664 3971 2704
rect 4063 2664 4065 2704
rect 4069 2664 4071 2704
rect 4083 2664 4085 2704
rect 4089 2692 4105 2704
rect 4089 2664 4091 2692
rect 4103 2664 4105 2692
rect 4109 2664 4111 2704
rect 4191 2664 4193 2704
rect 4197 2664 4203 2704
rect 4207 2664 4209 2704
rect 4309 2664 4311 2704
rect 4315 2664 4317 2704
rect 4409 2664 4411 2684
rect 4415 2664 4417 2684
rect 4469 2664 4471 2704
rect 4475 2684 4488 2704
rect 4651 2684 4661 2704
rect 4475 2664 4479 2684
rect 4491 2664 4493 2684
rect 4497 2664 4503 2684
rect 4507 2664 4509 2684
rect 4521 2664 4523 2684
rect 4527 2664 4531 2684
rect 4535 2664 4537 2684
rect 4575 2664 4577 2684
rect 4581 2664 4585 2684
rect 4597 2664 4599 2684
rect 4603 2664 4609 2684
rect 4613 2664 4615 2684
rect 4627 2664 4631 2684
rect 4635 2664 4641 2684
rect 4645 2664 4647 2684
rect 4659 2664 4661 2684
rect 4665 2664 4667 2704
rect 4713 2664 4715 2704
rect 4719 2684 4729 2704
rect 4892 2684 4905 2704
rect 4719 2664 4721 2684
rect 4733 2664 4735 2684
rect 4739 2664 4745 2684
rect 4749 2664 4753 2684
rect 4765 2664 4767 2684
rect 4771 2664 4777 2684
rect 4781 2664 4783 2684
rect 4795 2664 4799 2684
rect 4803 2664 4805 2684
rect 4843 2664 4845 2684
rect 4849 2664 4853 2684
rect 4857 2664 4859 2684
rect 4871 2664 4873 2684
rect 4877 2664 4883 2684
rect 4887 2664 4889 2684
rect 4901 2664 4905 2684
rect 4909 2664 4911 2704
rect 5009 2664 5011 2704
rect 5015 2692 5031 2704
rect 5015 2664 5017 2692
rect 5029 2664 5031 2692
rect 5035 2664 5037 2704
rect 5049 2664 5051 2704
rect 5055 2664 5057 2704
rect 5151 2664 5153 2704
rect 5157 2664 5163 2704
rect 5167 2664 5169 2704
rect 5269 2664 5271 2704
rect 5275 2664 5277 2704
rect 5289 2664 5291 2704
rect 5295 2664 5297 2704
rect 5349 2664 5351 2704
rect 5355 2684 5368 2704
rect 5531 2684 5541 2704
rect 5355 2664 5359 2684
rect 5371 2664 5373 2684
rect 5377 2664 5383 2684
rect 5387 2664 5389 2684
rect 5401 2664 5403 2684
rect 5407 2664 5411 2684
rect 5415 2664 5417 2684
rect 5455 2664 5457 2684
rect 5461 2664 5465 2684
rect 5477 2664 5479 2684
rect 5483 2664 5489 2684
rect 5493 2664 5495 2684
rect 5507 2664 5511 2684
rect 5515 2664 5521 2684
rect 5525 2664 5527 2684
rect 5539 2664 5541 2684
rect 5545 2664 5547 2704
rect 5629 2664 5631 2704
rect 5635 2692 5651 2704
rect 5635 2664 5637 2692
rect 5649 2664 5651 2692
rect 5655 2664 5657 2704
rect 5669 2664 5671 2704
rect 5675 2664 5677 2704
rect 83 2616 85 2636
rect 89 2616 91 2636
rect 169 2616 171 2636
rect 175 2616 177 2636
rect 290 2616 292 2636
rect 296 2616 300 2636
rect 312 2596 314 2636
rect 318 2596 322 2636
rect 326 2596 328 2636
rect 410 2576 412 2636
rect 416 2576 420 2636
rect 424 2576 428 2636
rect 432 2578 434 2636
rect 549 2616 551 2636
rect 555 2616 557 2636
rect 649 2616 651 2636
rect 655 2616 657 2636
rect 669 2616 671 2636
rect 675 2616 677 2636
rect 432 2576 446 2578
rect 769 2596 771 2636
rect 775 2608 777 2636
rect 789 2608 791 2636
rect 775 2596 791 2608
rect 795 2596 797 2636
rect 809 2596 811 2636
rect 815 2596 817 2636
rect 932 2596 934 2636
rect 938 2596 942 2636
rect 946 2596 948 2636
rect 960 2616 964 2636
rect 968 2616 970 2636
rect 1083 2596 1085 2636
rect 1089 2596 1091 2636
rect 1103 2596 1105 2636
rect 1109 2608 1111 2636
rect 1123 2608 1125 2636
rect 1109 2596 1125 2608
rect 1129 2596 1131 2636
rect 1231 2596 1233 2636
rect 1237 2596 1243 2636
rect 1247 2596 1249 2636
rect 1329 2596 1331 2636
rect 1335 2596 1341 2636
rect 1345 2596 1347 2636
rect 1359 2596 1361 2636
rect 1365 2596 1367 2636
rect 1506 2578 1508 2636
rect 1494 2576 1508 2578
rect 1512 2576 1516 2636
rect 1520 2576 1524 2636
rect 1528 2576 1530 2636
rect 1609 2616 1611 2636
rect 1615 2616 1617 2636
rect 1709 2596 1711 2636
rect 1715 2608 1717 2636
rect 1729 2608 1731 2636
rect 1715 2596 1731 2608
rect 1735 2596 1737 2636
rect 1749 2596 1751 2636
rect 1755 2596 1757 2636
rect 1863 2596 1865 2636
rect 1869 2596 1871 2636
rect 1883 2596 1885 2636
rect 1889 2608 1891 2636
rect 1903 2608 1905 2636
rect 1889 2596 1905 2608
rect 1909 2596 1911 2636
rect 1989 2596 1991 2636
rect 1995 2608 1997 2636
rect 2009 2608 2011 2636
rect 1995 2596 2011 2608
rect 2015 2596 2017 2636
rect 2029 2596 2031 2636
rect 2035 2596 2037 2636
rect 2166 2578 2168 2636
rect 2154 2576 2168 2578
rect 2172 2576 2176 2636
rect 2180 2576 2184 2636
rect 2188 2576 2190 2636
rect 2290 2616 2292 2636
rect 2296 2616 2300 2636
rect 2312 2596 2314 2636
rect 2318 2596 2322 2636
rect 2326 2596 2328 2636
rect 2411 2596 2413 2636
rect 2417 2596 2423 2636
rect 2427 2596 2429 2636
rect 2563 2596 2565 2636
rect 2569 2596 2571 2636
rect 2583 2596 2585 2636
rect 2589 2608 2591 2636
rect 2603 2608 2605 2636
rect 2589 2596 2605 2608
rect 2609 2596 2611 2636
rect 2689 2596 2691 2636
rect 2695 2608 2697 2636
rect 2709 2608 2711 2636
rect 2695 2596 2711 2608
rect 2715 2596 2717 2636
rect 2729 2596 2731 2636
rect 2735 2596 2737 2636
rect 2850 2616 2852 2636
rect 2856 2616 2860 2636
rect 2872 2596 2874 2636
rect 2878 2596 2882 2636
rect 2886 2596 2888 2636
rect 2983 2616 2985 2636
rect 2989 2616 2991 2636
rect 3069 2596 3071 2636
rect 3075 2608 3077 2636
rect 3089 2608 3091 2636
rect 3075 2596 3091 2608
rect 3095 2596 3097 2636
rect 3109 2596 3111 2636
rect 3115 2596 3117 2636
rect 3231 2596 3233 2636
rect 3237 2596 3243 2636
rect 3247 2596 3249 2636
rect 3386 2578 3388 2636
rect 3374 2576 3388 2578
rect 3392 2576 3396 2636
rect 3400 2576 3404 2636
rect 3408 2576 3410 2636
rect 3489 2596 3491 2636
rect 3495 2596 3501 2636
rect 3505 2596 3507 2636
rect 3519 2596 3521 2636
rect 3525 2596 3527 2636
rect 3631 2596 3633 2636
rect 3637 2596 3643 2636
rect 3647 2596 3649 2636
rect 3752 2596 3754 2636
rect 3758 2596 3762 2636
rect 3766 2596 3768 2636
rect 3780 2596 3782 2636
rect 3786 2596 3790 2636
rect 3794 2596 3796 2636
rect 3909 2616 3911 2636
rect 3915 2616 3917 2636
rect 3929 2616 3931 2636
rect 3935 2616 3937 2636
rect 3997 2616 3999 2636
rect 4003 2616 4005 2636
rect 4043 2596 4047 2636
rect 4051 2596 4059 2636
rect 4063 2596 4067 2636
rect 4079 2596 4084 2636
rect 4088 2596 4096 2636
rect 4100 2596 4104 2636
rect 4147 2616 4149 2636
rect 4153 2616 4155 2636
rect 4167 2616 4169 2636
rect 4173 2616 4175 2636
rect 4212 2616 4214 2636
rect 4218 2616 4220 2636
rect 4232 2616 4234 2636
rect 4238 2616 4240 2636
rect 4282 2616 4284 2636
rect 4288 2616 4290 2636
rect 4302 2616 4304 2636
rect 4308 2616 4310 2636
rect 4322 2616 4324 2636
rect 4328 2616 4330 2636
rect 4370 2596 4374 2636
rect 4378 2596 4386 2636
rect 4390 2596 4394 2636
rect 4406 2596 4410 2636
rect 4414 2596 4422 2636
rect 4426 2596 4430 2636
rect 4470 2596 4474 2636
rect 4478 2596 4486 2636
rect 4490 2596 4494 2636
rect 4506 2596 4510 2636
rect 4514 2596 4522 2636
rect 4526 2596 4530 2636
rect 4570 2616 4572 2636
rect 4576 2616 4578 2636
rect 4590 2616 4592 2636
rect 4596 2616 4598 2636
rect 4610 2616 4612 2636
rect 4616 2616 4618 2636
rect 4660 2616 4662 2636
rect 4666 2616 4668 2636
rect 4680 2616 4682 2636
rect 4686 2616 4688 2636
rect 4725 2616 4727 2636
rect 4731 2616 4733 2636
rect 4745 2616 4747 2636
rect 4751 2616 4753 2636
rect 4796 2596 4800 2636
rect 4804 2596 4812 2636
rect 4816 2596 4821 2636
rect 4833 2596 4837 2636
rect 4841 2596 4849 2636
rect 4853 2596 4857 2636
rect 4895 2616 4897 2636
rect 4901 2616 4903 2636
rect 4953 2596 4955 2636
rect 4959 2616 4961 2636
rect 4973 2616 4975 2636
rect 4979 2616 4985 2636
rect 4989 2616 4993 2636
rect 5005 2616 5007 2636
rect 5011 2616 5017 2636
rect 5021 2616 5023 2636
rect 5035 2616 5039 2636
rect 5043 2616 5045 2636
rect 5083 2616 5085 2636
rect 5089 2616 5093 2636
rect 5097 2616 5099 2636
rect 5111 2616 5113 2636
rect 5117 2616 5123 2636
rect 5127 2616 5129 2636
rect 5141 2616 5145 2636
rect 4959 2596 4969 2616
rect 5132 2596 5145 2616
rect 5149 2596 5151 2636
rect 5243 2596 5245 2636
rect 5249 2596 5251 2636
rect 5263 2596 5265 2636
rect 5269 2596 5271 2636
rect 5283 2596 5285 2636
rect 5289 2596 5291 2636
rect 5303 2596 5305 2636
rect 5309 2596 5311 2636
rect 5323 2596 5325 2636
rect 5329 2596 5331 2636
rect 5343 2596 5345 2636
rect 5349 2596 5351 2636
rect 5363 2596 5365 2636
rect 5369 2596 5371 2636
rect 5383 2596 5385 2636
rect 5389 2596 5391 2636
rect 5489 2596 5491 2636
rect 5495 2596 5497 2636
rect 5509 2596 5511 2636
rect 5515 2596 5517 2636
rect 5529 2596 5531 2636
rect 5535 2596 5537 2636
rect 5549 2596 5551 2636
rect 5555 2596 5557 2636
rect 5569 2596 5571 2636
rect 5575 2596 5577 2636
rect 5589 2596 5591 2636
rect 5595 2596 5597 2636
rect 5609 2596 5611 2636
rect 5615 2596 5617 2636
rect 5629 2596 5631 2636
rect 5635 2596 5637 2636
rect 5729 2596 5731 2636
rect 5735 2596 5737 2636
rect 81 2184 83 2224
rect 87 2184 89 2224
rect 214 2242 228 2244
rect 101 2184 105 2204
rect 109 2184 111 2204
rect 226 2184 228 2242
rect 232 2184 236 2244
rect 240 2184 244 2244
rect 248 2184 250 2244
rect 774 2242 788 2244
rect 331 2184 333 2224
rect 337 2184 343 2224
rect 347 2184 349 2224
rect 449 2184 451 2224
rect 455 2212 471 2224
rect 455 2184 457 2212
rect 469 2184 471 2212
rect 475 2184 477 2224
rect 489 2184 491 2224
rect 495 2184 497 2224
rect 603 2184 605 2224
rect 609 2184 611 2224
rect 623 2184 625 2224
rect 629 2212 645 2224
rect 629 2184 631 2212
rect 643 2184 645 2212
rect 649 2184 651 2224
rect 786 2184 788 2242
rect 792 2184 796 2244
rect 800 2184 804 2244
rect 808 2184 810 2244
rect 911 2184 913 2224
rect 917 2184 923 2224
rect 927 2184 929 2224
rect 1023 2184 1025 2224
rect 1029 2204 1041 2224
rect 1274 2242 1288 2244
rect 1029 2184 1031 2204
rect 1043 2184 1045 2204
rect 1049 2184 1051 2204
rect 1063 2184 1065 2204
rect 1069 2184 1071 2204
rect 1149 2184 1151 2224
rect 1155 2184 1157 2224
rect 1286 2184 1288 2242
rect 1292 2184 1296 2244
rect 1300 2184 1304 2244
rect 1308 2184 1310 2244
rect 1410 2184 1412 2204
rect 1416 2184 1420 2204
rect 1432 2184 1434 2224
rect 1438 2184 1442 2224
rect 1446 2184 1448 2224
rect 1563 2184 1565 2224
rect 1569 2184 1571 2224
rect 1583 2184 1585 2224
rect 1589 2212 1605 2224
rect 1589 2184 1591 2212
rect 1603 2184 1605 2212
rect 1609 2184 1611 2224
rect 1854 2242 1868 2244
rect 1710 2184 1712 2204
rect 1716 2184 1720 2204
rect 1732 2184 1734 2224
rect 1738 2184 1742 2224
rect 1746 2184 1748 2224
rect 1866 2184 1868 2242
rect 1872 2184 1876 2244
rect 1880 2184 1884 2244
rect 1888 2184 1890 2244
rect 1994 2242 2008 2244
rect 2006 2184 2008 2242
rect 2012 2184 2016 2244
rect 2020 2184 2024 2244
rect 2028 2184 2030 2244
rect 2077 2184 2079 2204
rect 2083 2184 2085 2204
rect 2123 2184 2127 2224
rect 2131 2184 2139 2224
rect 2143 2184 2147 2224
rect 2159 2184 2164 2224
rect 2168 2184 2176 2224
rect 2180 2184 2184 2224
rect 2227 2184 2229 2204
rect 2233 2184 2235 2204
rect 2247 2184 2249 2204
rect 2253 2184 2255 2204
rect 2292 2184 2294 2204
rect 2298 2184 2300 2204
rect 2312 2184 2314 2204
rect 2318 2184 2320 2204
rect 2362 2184 2364 2204
rect 2368 2184 2370 2204
rect 2382 2184 2384 2204
rect 2388 2184 2390 2204
rect 2402 2184 2404 2204
rect 2408 2184 2410 2204
rect 2450 2184 2454 2224
rect 2458 2184 2466 2224
rect 2470 2184 2474 2224
rect 2486 2184 2490 2224
rect 2494 2184 2502 2224
rect 2506 2184 2510 2224
rect 2601 2184 2603 2224
rect 2607 2184 2609 2224
rect 2621 2184 2625 2204
rect 2629 2184 2631 2204
rect 2729 2184 2731 2224
rect 2735 2212 2751 2224
rect 2735 2184 2737 2212
rect 2749 2184 2751 2212
rect 2755 2184 2757 2224
rect 2769 2184 2771 2224
rect 2775 2184 2777 2224
rect 2869 2184 2871 2224
rect 2875 2212 2891 2224
rect 2875 2184 2877 2212
rect 2889 2184 2891 2212
rect 2895 2184 2897 2224
rect 2909 2184 2911 2224
rect 2915 2184 2917 2224
rect 3031 2184 3033 2224
rect 3037 2184 3043 2224
rect 3047 2184 3049 2224
rect 3151 2184 3153 2224
rect 3157 2184 3163 2224
rect 3167 2184 3169 2224
rect 3290 2184 3292 2204
rect 3296 2184 3300 2204
rect 3312 2184 3314 2224
rect 3318 2184 3322 2224
rect 3326 2184 3328 2224
rect 3409 2184 3411 2204
rect 3415 2184 3417 2204
rect 3429 2184 3431 2204
rect 3435 2184 3437 2204
rect 3549 2184 3551 2224
rect 3555 2212 3571 2224
rect 3555 2184 3557 2212
rect 3569 2184 3571 2212
rect 3575 2184 3577 2224
rect 3589 2184 3591 2224
rect 3595 2184 3597 2224
rect 3691 2184 3693 2224
rect 3697 2184 3703 2224
rect 3707 2184 3709 2224
rect 3809 2184 3811 2204
rect 3815 2184 3819 2204
rect 3831 2184 3833 2224
rect 3837 2184 3839 2224
rect 3897 2184 3899 2204
rect 3903 2184 3905 2204
rect 3943 2184 3947 2224
rect 3951 2184 3959 2224
rect 3963 2184 3967 2224
rect 3979 2184 3984 2224
rect 3988 2184 3996 2224
rect 4000 2184 4004 2224
rect 4047 2184 4049 2204
rect 4053 2184 4055 2204
rect 4067 2184 4069 2204
rect 4073 2184 4075 2204
rect 4112 2184 4114 2204
rect 4118 2184 4120 2204
rect 4132 2184 4134 2204
rect 4138 2184 4140 2204
rect 4182 2184 4184 2204
rect 4188 2184 4190 2204
rect 4202 2184 4204 2204
rect 4208 2184 4210 2204
rect 4222 2184 4224 2204
rect 4228 2184 4230 2204
rect 4270 2184 4274 2224
rect 4278 2184 4286 2224
rect 4290 2184 4294 2224
rect 4306 2184 4310 2224
rect 4314 2184 4322 2224
rect 4326 2184 4330 2224
rect 4409 2184 4411 2224
rect 4415 2184 4421 2224
rect 4425 2184 4427 2224
rect 4439 2184 4441 2224
rect 4445 2184 4447 2224
rect 4552 2184 4554 2224
rect 4558 2184 4562 2224
rect 4566 2184 4568 2224
rect 4580 2184 4582 2224
rect 4586 2184 4590 2224
rect 4594 2184 4596 2224
rect 4711 2184 4713 2224
rect 4717 2184 4723 2224
rect 4727 2184 4729 2224
rect 4841 2184 4843 2224
rect 4847 2184 4849 2224
rect 4861 2184 4865 2204
rect 4869 2184 4871 2204
rect 4949 2184 4951 2204
rect 4955 2184 4957 2204
rect 5052 2184 5054 2224
rect 5058 2184 5062 2224
rect 5066 2184 5068 2224
rect 5080 2184 5082 2224
rect 5086 2184 5090 2224
rect 5094 2184 5096 2224
rect 5211 2184 5213 2224
rect 5217 2184 5223 2224
rect 5227 2184 5229 2224
rect 5329 2184 5331 2224
rect 5335 2184 5337 2224
rect 5431 2184 5433 2224
rect 5437 2184 5443 2224
rect 5447 2184 5449 2224
rect 5659 2212 5671 2232
rect 5549 2184 5551 2204
rect 5555 2184 5557 2204
rect 5649 2192 5651 2212
rect 5655 2192 5657 2212
rect 5669 2192 5671 2212
rect 5675 2192 5681 2232
rect 5685 2224 5701 2232
rect 5685 2192 5687 2224
rect 5699 2192 5701 2224
rect 5705 2192 5711 2232
rect 5715 2192 5717 2232
rect 101 2116 103 2156
rect 107 2116 109 2156
rect 121 2136 125 2156
rect 129 2136 131 2156
rect 266 2098 268 2156
rect 254 2096 268 2098
rect 272 2096 276 2156
rect 280 2096 284 2156
rect 288 2096 290 2156
rect 372 2116 374 2156
rect 378 2116 382 2156
rect 386 2116 388 2156
rect 400 2136 404 2156
rect 408 2136 410 2156
rect 523 2136 525 2156
rect 529 2136 531 2156
rect 623 2116 625 2156
rect 629 2116 631 2156
rect 643 2116 645 2156
rect 649 2128 651 2156
rect 663 2128 665 2156
rect 649 2116 665 2128
rect 669 2116 671 2156
rect 770 2136 772 2156
rect 776 2136 780 2156
rect 792 2116 794 2156
rect 798 2116 802 2156
rect 806 2116 808 2156
rect 890 2096 892 2156
rect 896 2096 900 2156
rect 904 2096 908 2156
rect 912 2098 914 2156
rect 912 2096 926 2098
rect 1086 2098 1088 2156
rect 1074 2096 1088 2098
rect 1092 2096 1096 2156
rect 1100 2096 1104 2156
rect 1108 2096 1110 2156
rect 1203 2116 1205 2156
rect 1209 2116 1211 2156
rect 1223 2116 1225 2156
rect 1229 2128 1231 2156
rect 1243 2128 1245 2156
rect 1229 2116 1245 2128
rect 1249 2116 1251 2156
rect 1343 2116 1345 2156
rect 1349 2116 1351 2156
rect 1363 2116 1365 2156
rect 1369 2128 1371 2156
rect 1383 2128 1385 2156
rect 1369 2116 1385 2128
rect 1389 2116 1391 2156
rect 1490 2136 1492 2156
rect 1496 2136 1500 2156
rect 1512 2116 1514 2156
rect 1518 2116 1522 2156
rect 1526 2116 1528 2156
rect 1646 2098 1648 2156
rect 1634 2096 1648 2098
rect 1652 2096 1656 2156
rect 1660 2096 1664 2156
rect 1668 2096 1670 2156
rect 1749 2116 1751 2156
rect 1755 2128 1757 2156
rect 1769 2128 1771 2156
rect 1755 2116 1771 2128
rect 1775 2116 1777 2156
rect 1789 2116 1791 2156
rect 1795 2116 1797 2156
rect 1892 2116 1894 2156
rect 1898 2116 1902 2156
rect 1906 2116 1908 2156
rect 1920 2136 1924 2156
rect 1928 2136 1930 2156
rect 2103 2136 2105 2156
rect 2109 2136 2111 2156
rect 2123 2136 2125 2156
rect 2129 2136 2131 2156
rect 2143 2136 2145 2156
rect 2149 2136 2151 2156
rect 2286 2098 2288 2156
rect 2274 2096 2288 2098
rect 2292 2096 2296 2156
rect 2300 2096 2304 2156
rect 2308 2096 2310 2156
rect 2357 2136 2359 2156
rect 2363 2136 2365 2156
rect 2403 2116 2407 2156
rect 2411 2116 2419 2156
rect 2423 2116 2427 2156
rect 2439 2116 2444 2156
rect 2448 2116 2456 2156
rect 2460 2116 2464 2156
rect 2507 2136 2509 2156
rect 2513 2136 2515 2156
rect 2527 2136 2529 2156
rect 2533 2136 2535 2156
rect 2572 2136 2574 2156
rect 2578 2136 2580 2156
rect 2592 2136 2594 2156
rect 2598 2136 2600 2156
rect 2642 2136 2644 2156
rect 2648 2136 2650 2156
rect 2662 2136 2664 2156
rect 2668 2136 2670 2156
rect 2682 2136 2684 2156
rect 2688 2136 2690 2156
rect 2730 2116 2734 2156
rect 2738 2116 2746 2156
rect 2750 2116 2754 2156
rect 2766 2116 2770 2156
rect 2774 2116 2782 2156
rect 2786 2116 2790 2156
rect 2869 2116 2871 2156
rect 2875 2128 2877 2156
rect 2889 2128 2891 2156
rect 2875 2116 2891 2128
rect 2895 2116 2897 2156
rect 2909 2116 2911 2156
rect 2915 2116 2917 2156
rect 3031 2116 3033 2156
rect 3037 2116 3043 2156
rect 3047 2116 3049 2156
rect 3131 2116 3133 2156
rect 3137 2116 3143 2156
rect 3147 2116 3149 2156
rect 3269 2136 3271 2156
rect 3275 2136 3277 2156
rect 3289 2136 3291 2156
rect 3295 2136 3297 2156
rect 3413 2116 3415 2156
rect 3419 2116 3421 2156
rect 3433 2116 3435 2156
rect 3439 2116 3445 2156
rect 3449 2116 3451 2156
rect 3532 2116 3534 2156
rect 3538 2116 3542 2156
rect 3546 2116 3548 2156
rect 3560 2136 3564 2156
rect 3568 2136 3570 2156
rect 3703 2116 3705 2156
rect 3709 2116 3711 2156
rect 3810 2096 3812 2156
rect 3816 2096 3820 2156
rect 3824 2096 3828 2156
rect 3832 2098 3834 2156
rect 3969 2116 3971 2156
rect 3975 2116 3977 2156
rect 4113 2116 4115 2156
rect 4119 2116 4121 2156
rect 4133 2116 4135 2156
rect 4139 2116 4145 2156
rect 4149 2116 4151 2156
rect 4251 2116 4253 2156
rect 4257 2116 4263 2156
rect 4267 2116 4269 2156
rect 4363 2116 4365 2156
rect 4369 2116 4371 2156
rect 4383 2116 4385 2156
rect 4389 2128 4391 2156
rect 4403 2128 4405 2156
rect 4389 2116 4405 2128
rect 4409 2116 4411 2156
rect 4489 2116 4491 2156
rect 4495 2128 4497 2156
rect 4509 2128 4511 2156
rect 4495 2116 4511 2128
rect 4515 2116 4517 2156
rect 4529 2116 4531 2156
rect 4535 2116 4537 2156
rect 4631 2116 4633 2156
rect 4637 2116 4643 2156
rect 4647 2116 4649 2156
rect 4751 2116 4753 2156
rect 4757 2116 4763 2156
rect 4767 2116 4769 2156
rect 4903 2116 4905 2156
rect 4909 2116 4911 2156
rect 4923 2116 4925 2156
rect 4929 2128 4931 2156
rect 4943 2128 4945 2156
rect 4929 2116 4945 2128
rect 4949 2116 4951 2156
rect 5043 2116 5045 2156
rect 5049 2116 5051 2156
rect 5063 2116 5065 2156
rect 5069 2128 5071 2156
rect 5083 2128 5085 2156
rect 5069 2116 5085 2128
rect 5089 2116 5091 2156
rect 5169 2136 5171 2156
rect 5175 2136 5177 2156
rect 5269 2136 5271 2156
rect 5275 2136 5277 2156
rect 5289 2136 5291 2156
rect 5295 2136 5297 2156
rect 3832 2096 3846 2098
rect 5391 2116 5393 2156
rect 5397 2116 5403 2156
rect 5407 2116 5409 2156
rect 5509 2136 5511 2156
rect 5515 2136 5517 2156
rect 5623 2136 5625 2156
rect 5629 2136 5631 2156
rect 5709 2116 5711 2156
rect 5715 2128 5717 2156
rect 5729 2128 5731 2156
rect 5715 2116 5731 2128
rect 5735 2116 5737 2156
rect 5749 2116 5751 2156
rect 5755 2116 5757 2156
rect 94 1762 108 1764
rect 106 1704 108 1762
rect 112 1704 116 1764
rect 120 1704 124 1764
rect 128 1704 130 1764
rect 212 1704 214 1744
rect 218 1704 222 1744
rect 226 1704 228 1744
rect 514 1762 528 1764
rect 240 1704 244 1724
rect 248 1704 250 1724
rect 363 1704 365 1744
rect 369 1704 371 1744
rect 383 1704 385 1744
rect 389 1732 405 1744
rect 389 1704 391 1732
rect 403 1704 405 1732
rect 409 1704 411 1744
rect 526 1704 528 1762
rect 532 1704 536 1764
rect 540 1704 544 1764
rect 548 1704 550 1764
rect 663 1704 665 1724
rect 669 1704 671 1724
rect 683 1704 685 1724
rect 689 1704 691 1724
rect 772 1704 774 1744
rect 778 1704 782 1744
rect 786 1704 788 1744
rect 800 1704 804 1724
rect 808 1704 810 1724
rect 943 1704 945 1724
rect 949 1704 951 1724
rect 1063 1704 1065 1744
rect 1069 1704 1071 1744
rect 1083 1704 1085 1744
rect 1089 1732 1105 1744
rect 1089 1704 1091 1732
rect 1103 1704 1105 1732
rect 1109 1704 1111 1744
rect 1203 1704 1205 1744
rect 1209 1704 1211 1744
rect 1223 1704 1225 1744
rect 1229 1732 1245 1744
rect 1229 1704 1231 1732
rect 1243 1704 1245 1732
rect 1249 1704 1251 1744
rect 1343 1704 1345 1724
rect 1349 1704 1351 1724
rect 1443 1704 1445 1744
rect 1449 1704 1451 1744
rect 1463 1704 1465 1744
rect 1469 1732 1485 1744
rect 1469 1704 1471 1732
rect 1483 1704 1485 1732
rect 1489 1704 1491 1744
rect 1569 1704 1571 1744
rect 1575 1732 1591 1744
rect 1575 1704 1577 1732
rect 1589 1704 1591 1732
rect 1595 1704 1597 1744
rect 1609 1704 1611 1744
rect 1615 1704 1617 1744
rect 1723 1704 1725 1744
rect 1729 1704 1731 1744
rect 1743 1704 1745 1744
rect 1749 1732 1765 1744
rect 1749 1704 1751 1732
rect 1763 1704 1765 1732
rect 1769 1704 1771 1744
rect 1871 1704 1873 1744
rect 1877 1704 1883 1744
rect 1887 1704 1889 1744
rect 1991 1704 1993 1744
rect 1997 1704 2003 1744
rect 2007 1704 2009 1744
rect 2123 1704 2125 1744
rect 2129 1704 2131 1744
rect 2143 1704 2145 1744
rect 2149 1704 2151 1744
rect 2197 1704 2199 1724
rect 2203 1704 2205 1724
rect 2243 1704 2247 1744
rect 2251 1704 2259 1744
rect 2263 1704 2267 1744
rect 2279 1704 2284 1744
rect 2288 1704 2296 1744
rect 2300 1704 2304 1744
rect 2854 1762 2868 1764
rect 2347 1704 2349 1724
rect 2353 1704 2355 1724
rect 2367 1704 2369 1724
rect 2373 1704 2375 1724
rect 2412 1704 2414 1724
rect 2418 1704 2420 1724
rect 2432 1704 2434 1724
rect 2438 1704 2440 1724
rect 2482 1704 2484 1724
rect 2488 1704 2490 1724
rect 2502 1704 2504 1724
rect 2508 1704 2510 1724
rect 2522 1704 2524 1724
rect 2528 1704 2530 1724
rect 2570 1704 2574 1744
rect 2578 1704 2586 1744
rect 2590 1704 2594 1744
rect 2606 1704 2610 1744
rect 2614 1704 2622 1744
rect 2626 1704 2630 1744
rect 2711 1704 2713 1744
rect 2717 1704 2723 1744
rect 2727 1704 2729 1744
rect 2866 1704 2868 1762
rect 2872 1704 2876 1764
rect 2880 1704 2884 1764
rect 2888 1704 2890 1764
rect 2983 1704 2985 1744
rect 2989 1704 2991 1744
rect 3003 1704 3005 1744
rect 3009 1732 3025 1744
rect 3009 1704 3011 1732
rect 3023 1704 3025 1732
rect 3029 1704 3031 1744
rect 3239 1732 3251 1752
rect 3109 1704 3111 1724
rect 3115 1704 3117 1724
rect 3129 1704 3131 1724
rect 3135 1704 3137 1724
rect 3229 1712 3231 1732
rect 3235 1712 3237 1732
rect 3249 1712 3251 1732
rect 3255 1712 3261 1752
rect 3265 1744 3281 1752
rect 3265 1712 3267 1744
rect 3279 1712 3281 1744
rect 3285 1712 3291 1752
rect 3295 1712 3297 1752
rect 3403 1704 3405 1724
rect 3409 1704 3411 1724
rect 3489 1704 3491 1744
rect 3495 1734 3511 1744
rect 3495 1704 3497 1734
rect 3509 1704 3511 1734
rect 3515 1704 3517 1744
rect 3529 1704 3531 1744
rect 3535 1716 3537 1744
rect 3549 1716 3551 1744
rect 3535 1704 3551 1716
rect 3555 1704 3557 1744
rect 3663 1704 3665 1744
rect 3669 1704 3671 1744
rect 3683 1704 3685 1744
rect 3689 1732 3705 1744
rect 3689 1704 3691 1732
rect 3703 1704 3705 1732
rect 3709 1704 3711 1744
rect 3823 1704 3825 1744
rect 3829 1704 3831 1744
rect 3843 1704 3845 1744
rect 3849 1732 3865 1744
rect 3849 1704 3851 1732
rect 3863 1704 3865 1732
rect 3869 1704 3871 1744
rect 3949 1704 3951 1744
rect 3955 1732 3971 1744
rect 3955 1704 3957 1732
rect 3969 1704 3971 1732
rect 3975 1704 3977 1744
rect 3989 1704 3991 1744
rect 3995 1704 3997 1744
rect 4111 1704 4113 1744
rect 4117 1704 4123 1744
rect 4127 1704 4129 1744
rect 4244 1704 4246 1744
rect 4250 1704 4254 1744
rect 4258 1704 4260 1744
rect 4272 1704 4274 1744
rect 4278 1704 4282 1744
rect 4286 1704 4288 1744
rect 4391 1704 4393 1744
rect 4397 1704 4403 1744
rect 4407 1704 4409 1744
rect 4489 1704 4491 1744
rect 4495 1732 4511 1744
rect 4495 1704 4497 1732
rect 4509 1704 4511 1732
rect 4515 1704 4517 1744
rect 4529 1704 4531 1744
rect 4535 1704 4537 1744
rect 4653 1704 4655 1744
rect 4659 1704 4661 1744
rect 4673 1704 4675 1744
rect 4679 1704 4685 1744
rect 4689 1704 4691 1744
rect 4783 1704 4785 1724
rect 4789 1704 4791 1724
rect 4803 1704 4805 1724
rect 4809 1704 4811 1724
rect 4911 1704 4913 1744
rect 4917 1704 4923 1744
rect 4927 1704 4929 1744
rect 5044 1704 5046 1744
rect 5050 1704 5054 1744
rect 5058 1704 5060 1744
rect 5072 1704 5074 1744
rect 5078 1704 5082 1744
rect 5086 1704 5088 1744
rect 5183 1704 5185 1724
rect 5189 1704 5191 1724
rect 5283 1704 5285 1724
rect 5289 1704 5291 1724
rect 5303 1704 5305 1724
rect 5309 1704 5311 1724
rect 5389 1704 5391 1744
rect 5395 1732 5411 1744
rect 5395 1704 5397 1732
rect 5409 1704 5411 1732
rect 5415 1704 5417 1744
rect 5429 1704 5431 1744
rect 5435 1704 5437 1744
rect 5543 1704 5545 1744
rect 5549 1704 5551 1744
rect 5563 1704 5565 1744
rect 5569 1732 5585 1744
rect 5569 1704 5571 1732
rect 5583 1704 5585 1732
rect 5589 1704 5591 1744
rect 5669 1704 5671 1744
rect 5675 1704 5677 1744
rect 5689 1704 5691 1744
rect 5695 1704 5697 1744
rect 90 1616 92 1676
rect 96 1616 100 1676
rect 104 1616 108 1676
rect 112 1618 114 1676
rect 112 1616 126 1618
rect 266 1618 268 1676
rect 254 1616 268 1618
rect 272 1616 276 1676
rect 280 1616 284 1676
rect 288 1616 290 1676
rect 372 1636 374 1676
rect 378 1636 382 1676
rect 386 1636 388 1676
rect 400 1656 404 1676
rect 408 1656 410 1676
rect 530 1656 532 1676
rect 536 1656 540 1676
rect 552 1636 554 1676
rect 558 1636 562 1676
rect 566 1636 568 1676
rect 651 1636 653 1676
rect 657 1636 663 1676
rect 667 1636 669 1676
rect 769 1656 771 1676
rect 775 1656 777 1676
rect 883 1636 885 1676
rect 889 1636 891 1676
rect 903 1636 905 1676
rect 909 1648 911 1676
rect 923 1648 925 1676
rect 909 1636 925 1648
rect 929 1636 931 1676
rect 1046 1618 1048 1676
rect 1034 1616 1048 1618
rect 1052 1616 1056 1676
rect 1060 1616 1064 1676
rect 1068 1616 1070 1676
rect 1171 1636 1173 1676
rect 1177 1636 1183 1676
rect 1187 1636 1189 1676
rect 1289 1656 1291 1676
rect 1295 1656 1297 1676
rect 1309 1656 1311 1676
rect 1315 1656 1317 1676
rect 1421 1636 1423 1676
rect 1427 1636 1429 1676
rect 1441 1656 1445 1676
rect 1449 1656 1451 1676
rect 1563 1656 1565 1676
rect 1569 1656 1571 1676
rect 1652 1636 1654 1676
rect 1658 1636 1662 1676
rect 1666 1636 1668 1676
rect 1680 1636 1682 1676
rect 1686 1636 1690 1676
rect 1694 1636 1696 1676
rect 1777 1656 1779 1676
rect 1783 1656 1785 1676
rect 1823 1636 1827 1676
rect 1831 1636 1839 1676
rect 1843 1636 1847 1676
rect 1859 1636 1864 1676
rect 1868 1636 1876 1676
rect 1880 1636 1884 1676
rect 1927 1656 1929 1676
rect 1933 1656 1935 1676
rect 1947 1656 1949 1676
rect 1953 1656 1955 1676
rect 1992 1656 1994 1676
rect 1998 1656 2000 1676
rect 2012 1656 2014 1676
rect 2018 1656 2020 1676
rect 2062 1656 2064 1676
rect 2068 1656 2070 1676
rect 2082 1656 2084 1676
rect 2088 1656 2090 1676
rect 2102 1656 2104 1676
rect 2108 1656 2110 1676
rect 2150 1636 2154 1676
rect 2158 1636 2166 1676
rect 2170 1636 2174 1676
rect 2186 1636 2190 1676
rect 2194 1636 2202 1676
rect 2206 1636 2210 1676
rect 2309 1636 2311 1676
rect 2315 1648 2317 1676
rect 2329 1648 2331 1676
rect 2315 1636 2331 1648
rect 2335 1636 2337 1676
rect 2349 1636 2351 1676
rect 2355 1636 2357 1676
rect 2451 1636 2453 1676
rect 2457 1636 2463 1676
rect 2467 1636 2469 1676
rect 2583 1636 2585 1676
rect 2589 1636 2591 1676
rect 2603 1636 2605 1676
rect 2609 1648 2611 1676
rect 2623 1648 2625 1676
rect 2609 1636 2625 1648
rect 2629 1636 2631 1676
rect 2731 1636 2733 1676
rect 2737 1636 2743 1676
rect 2747 1636 2749 1676
rect 2843 1636 2845 1676
rect 2849 1636 2851 1676
rect 2863 1636 2865 1676
rect 2869 1648 2871 1676
rect 2883 1648 2885 1676
rect 2869 1636 2885 1648
rect 2889 1636 2891 1676
rect 2983 1636 2985 1676
rect 2989 1636 2991 1676
rect 3003 1636 3005 1676
rect 3009 1648 3011 1676
rect 3023 1648 3025 1676
rect 3009 1636 3025 1648
rect 3029 1636 3031 1676
rect 3070 1636 3074 1676
rect 3078 1636 3086 1676
rect 3090 1636 3094 1676
rect 3106 1636 3110 1676
rect 3114 1636 3122 1676
rect 3126 1636 3130 1676
rect 3170 1656 3172 1676
rect 3176 1656 3178 1676
rect 3190 1656 3192 1676
rect 3196 1656 3198 1676
rect 3210 1656 3212 1676
rect 3216 1656 3218 1676
rect 3260 1656 3262 1676
rect 3266 1656 3268 1676
rect 3280 1656 3282 1676
rect 3286 1656 3288 1676
rect 3325 1656 3327 1676
rect 3331 1656 3333 1676
rect 3345 1656 3347 1676
rect 3351 1656 3353 1676
rect 3396 1636 3400 1676
rect 3404 1636 3412 1676
rect 3416 1636 3421 1676
rect 3433 1636 3437 1676
rect 3441 1636 3449 1676
rect 3453 1636 3457 1676
rect 3495 1656 3497 1676
rect 3501 1656 3503 1676
rect 3610 1656 3612 1676
rect 3616 1656 3620 1676
rect 3632 1636 3634 1676
rect 3638 1636 3642 1676
rect 3646 1636 3648 1676
rect 3729 1636 3731 1676
rect 3735 1648 3737 1676
rect 3749 1648 3751 1676
rect 3735 1636 3751 1648
rect 3755 1636 3757 1676
rect 3769 1636 3771 1676
rect 3775 1636 3777 1676
rect 3881 1636 3883 1676
rect 3887 1636 3889 1676
rect 3901 1656 3905 1676
rect 3909 1656 3911 1676
rect 4013 1636 4015 1676
rect 4019 1636 4021 1676
rect 4033 1636 4035 1676
rect 4039 1636 4045 1676
rect 4049 1636 4051 1676
rect 4131 1636 4133 1676
rect 4137 1636 4143 1676
rect 4147 1636 4149 1676
rect 4284 1636 4286 1676
rect 4290 1636 4294 1676
rect 4298 1636 4300 1676
rect 4312 1636 4314 1676
rect 4318 1636 4322 1676
rect 4326 1636 4328 1676
rect 4444 1636 4446 1676
rect 4450 1636 4454 1676
rect 4458 1636 4460 1676
rect 4472 1636 4474 1676
rect 4478 1636 4482 1676
rect 4486 1636 4488 1676
rect 4592 1636 4594 1676
rect 4598 1636 4602 1676
rect 4606 1636 4608 1676
rect 4620 1636 4622 1676
rect 4626 1636 4630 1676
rect 4634 1636 4636 1676
rect 4751 1636 4753 1676
rect 4757 1636 4763 1676
rect 4767 1636 4769 1676
rect 4869 1636 4871 1676
rect 4875 1648 4877 1676
rect 4889 1648 4891 1676
rect 4875 1636 4891 1648
rect 4895 1636 4897 1676
rect 4909 1636 4911 1676
rect 4915 1636 4917 1676
rect 5033 1636 5035 1676
rect 5039 1636 5041 1676
rect 5053 1636 5055 1676
rect 5059 1636 5065 1676
rect 5069 1636 5071 1676
rect 5170 1616 5172 1676
rect 5176 1616 5180 1676
rect 5184 1616 5188 1676
rect 5192 1618 5194 1676
rect 5312 1636 5314 1676
rect 5318 1636 5322 1676
rect 5326 1636 5328 1676
rect 5340 1636 5342 1676
rect 5346 1636 5350 1676
rect 5354 1636 5356 1676
rect 5471 1636 5473 1676
rect 5477 1636 5483 1676
rect 5487 1636 5489 1676
rect 5192 1616 5206 1618
rect 5590 1616 5592 1676
rect 5596 1616 5600 1676
rect 5604 1616 5608 1676
rect 5612 1618 5614 1676
rect 5763 1636 5765 1676
rect 5769 1636 5771 1676
rect 5612 1616 5626 1618
rect 94 1282 108 1284
rect 106 1224 108 1282
rect 112 1224 116 1284
rect 120 1224 124 1284
rect 128 1224 130 1284
rect 212 1224 214 1264
rect 218 1224 222 1264
rect 226 1224 228 1264
rect 374 1282 388 1284
rect 240 1224 244 1244
rect 248 1224 250 1244
rect 386 1224 388 1282
rect 392 1224 396 1284
rect 400 1224 404 1284
rect 408 1224 410 1284
rect 503 1224 505 1264
rect 509 1224 511 1264
rect 523 1224 525 1264
rect 529 1252 545 1264
rect 529 1224 531 1252
rect 543 1224 545 1252
rect 549 1224 551 1264
rect 643 1224 645 1264
rect 649 1224 651 1264
rect 663 1224 665 1264
rect 669 1252 685 1264
rect 669 1224 671 1252
rect 683 1224 685 1252
rect 689 1224 691 1264
rect 813 1224 815 1264
rect 819 1224 821 1264
rect 833 1224 835 1264
rect 839 1224 845 1264
rect 849 1224 851 1264
rect 931 1224 933 1264
rect 937 1224 943 1264
rect 947 1224 949 1264
rect 1063 1224 1065 1244
rect 1069 1224 1071 1244
rect 1150 1224 1152 1284
rect 1156 1224 1160 1284
rect 1164 1224 1168 1284
rect 1172 1282 1186 1284
rect 1172 1224 1174 1282
rect 1694 1282 1708 1284
rect 1291 1224 1293 1264
rect 1297 1224 1303 1264
rect 1307 1224 1309 1264
rect 1431 1224 1433 1264
rect 1437 1224 1443 1264
rect 1447 1224 1449 1264
rect 1551 1224 1553 1264
rect 1557 1224 1563 1264
rect 1567 1224 1569 1264
rect 1706 1224 1708 1282
rect 1712 1224 1716 1284
rect 1720 1224 1724 1284
rect 1728 1224 1730 1284
rect 1954 1282 1968 1284
rect 1811 1224 1813 1264
rect 1817 1224 1823 1264
rect 1827 1224 1829 1264
rect 1966 1224 1968 1282
rect 1972 1224 1976 1284
rect 1980 1224 1984 1284
rect 1988 1224 1990 1284
rect 2214 1282 2228 1284
rect 2083 1224 2085 1244
rect 2089 1224 2091 1244
rect 2226 1224 2228 1282
rect 2232 1224 2236 1284
rect 2240 1224 2244 1284
rect 2248 1224 2250 1284
rect 2354 1282 2368 1284
rect 2366 1224 2368 1282
rect 2372 1224 2376 1284
rect 2380 1224 2384 1284
rect 2388 1224 2390 1284
rect 2469 1224 2471 1244
rect 2475 1224 2477 1244
rect 2603 1224 2605 1264
rect 2609 1224 2611 1264
rect 2623 1224 2625 1264
rect 2629 1252 2645 1264
rect 2629 1224 2631 1252
rect 2643 1224 2645 1252
rect 2649 1224 2651 1264
rect 2732 1224 2734 1264
rect 2738 1224 2742 1264
rect 2746 1224 2748 1264
rect 2760 1224 2764 1244
rect 2768 1224 2770 1244
rect 2883 1224 2885 1264
rect 2889 1224 2891 1264
rect 2903 1224 2905 1264
rect 2909 1252 2925 1264
rect 2909 1224 2911 1252
rect 2923 1224 2925 1252
rect 2929 1224 2931 1264
rect 3023 1224 3025 1264
rect 3029 1224 3031 1264
rect 3043 1224 3045 1264
rect 3049 1252 3065 1264
rect 3049 1224 3051 1252
rect 3063 1224 3065 1252
rect 3069 1224 3071 1264
rect 3163 1224 3165 1264
rect 3169 1224 3171 1264
rect 3183 1224 3185 1264
rect 3189 1252 3205 1264
rect 3189 1224 3191 1252
rect 3203 1224 3205 1252
rect 3209 1224 3211 1264
rect 3303 1224 3305 1244
rect 3309 1224 3311 1244
rect 3389 1224 3391 1244
rect 3395 1224 3397 1244
rect 3501 1224 3503 1264
rect 3507 1224 3509 1264
rect 3521 1224 3525 1244
rect 3529 1224 3531 1244
rect 3650 1224 3652 1244
rect 3656 1224 3660 1244
rect 3672 1224 3674 1264
rect 3678 1224 3682 1264
rect 3686 1224 3688 1264
rect 3769 1224 3771 1264
rect 3775 1252 3791 1264
rect 3775 1224 3777 1252
rect 3789 1224 3791 1252
rect 3795 1224 3797 1264
rect 3809 1224 3811 1264
rect 3815 1224 3817 1264
rect 3923 1224 3925 1244
rect 3929 1224 3931 1244
rect 4023 1224 4025 1264
rect 4029 1224 4031 1264
rect 4043 1224 4045 1264
rect 4049 1252 4065 1264
rect 4049 1224 4051 1252
rect 4063 1224 4065 1252
rect 4069 1224 4071 1264
rect 4163 1224 4165 1264
rect 4169 1224 4171 1264
rect 4183 1224 4185 1264
rect 4189 1252 4205 1264
rect 4189 1224 4191 1252
rect 4203 1224 4205 1252
rect 4209 1224 4211 1264
rect 4310 1224 4312 1244
rect 4316 1224 4320 1244
rect 4332 1224 4334 1264
rect 4338 1224 4342 1264
rect 4346 1224 4348 1264
rect 4443 1224 4445 1264
rect 4449 1224 4451 1264
rect 4463 1224 4465 1264
rect 4469 1252 4485 1264
rect 4469 1224 4471 1252
rect 4483 1224 4485 1252
rect 4489 1224 4491 1264
rect 4589 1224 4591 1264
rect 4595 1252 4611 1264
rect 4595 1224 4597 1252
rect 4609 1224 4611 1252
rect 4615 1224 4617 1264
rect 4629 1224 4631 1264
rect 4635 1224 4637 1264
rect 4731 1224 4733 1264
rect 4737 1224 4743 1264
rect 4747 1224 4749 1264
rect 4849 1224 4851 1264
rect 4855 1252 4871 1264
rect 4855 1224 4857 1252
rect 4869 1224 4871 1252
rect 4875 1224 4877 1264
rect 4889 1224 4891 1264
rect 4895 1224 4897 1264
rect 4989 1224 4991 1244
rect 4995 1224 4997 1244
rect 5009 1224 5011 1244
rect 5015 1224 5017 1244
rect 5111 1224 5113 1264
rect 5117 1224 5123 1264
rect 5127 1224 5129 1264
rect 5251 1224 5253 1264
rect 5257 1224 5263 1264
rect 5267 1224 5269 1264
rect 5363 1224 5365 1264
rect 5369 1224 5371 1264
rect 5383 1224 5385 1264
rect 5389 1252 5405 1264
rect 5389 1224 5391 1252
rect 5403 1224 5405 1252
rect 5409 1224 5411 1264
rect 5489 1224 5491 1264
rect 5495 1252 5511 1264
rect 5495 1224 5497 1252
rect 5509 1224 5511 1252
rect 5515 1224 5517 1264
rect 5529 1224 5531 1264
rect 5535 1224 5537 1264
rect 5649 1224 5651 1264
rect 5655 1252 5671 1264
rect 5655 1224 5657 1252
rect 5669 1224 5671 1252
rect 5675 1224 5677 1264
rect 5689 1224 5691 1264
rect 5695 1224 5697 1264
rect 83 1176 85 1196
rect 89 1176 91 1196
rect 172 1156 174 1196
rect 178 1156 182 1196
rect 186 1156 188 1196
rect 200 1176 204 1196
rect 208 1176 210 1196
rect 309 1156 311 1196
rect 315 1168 317 1196
rect 329 1168 331 1196
rect 315 1156 331 1168
rect 335 1156 337 1196
rect 349 1156 351 1196
rect 355 1156 357 1196
rect 449 1156 451 1196
rect 455 1168 457 1196
rect 469 1168 471 1196
rect 455 1156 471 1168
rect 475 1156 477 1196
rect 489 1156 491 1196
rect 495 1156 497 1196
rect 626 1138 628 1196
rect 614 1136 628 1138
rect 632 1136 636 1196
rect 640 1136 644 1196
rect 648 1136 650 1196
rect 729 1156 731 1196
rect 735 1168 737 1196
rect 749 1168 751 1196
rect 735 1156 751 1168
rect 755 1156 757 1196
rect 769 1156 771 1196
rect 775 1156 777 1196
rect 892 1156 894 1196
rect 898 1156 902 1196
rect 906 1156 908 1196
rect 920 1176 924 1196
rect 928 1176 930 1196
rect 1043 1156 1045 1196
rect 1049 1156 1051 1196
rect 1063 1156 1065 1196
rect 1069 1168 1071 1196
rect 1083 1168 1085 1196
rect 1069 1156 1085 1168
rect 1089 1156 1091 1196
rect 1183 1176 1185 1196
rect 1189 1176 1191 1196
rect 1272 1156 1274 1196
rect 1278 1156 1282 1196
rect 1286 1156 1288 1196
rect 1300 1176 1304 1196
rect 1308 1176 1310 1196
rect 1423 1176 1425 1196
rect 1429 1176 1431 1196
rect 1523 1176 1525 1196
rect 1529 1176 1531 1196
rect 1543 1176 1545 1196
rect 1549 1176 1551 1196
rect 1649 1176 1651 1196
rect 1655 1176 1657 1196
rect 1786 1138 1788 1196
rect 1774 1136 1788 1138
rect 1792 1136 1796 1196
rect 1800 1136 1804 1196
rect 1808 1136 1810 1196
rect 1911 1156 1913 1196
rect 1917 1156 1923 1196
rect 1927 1156 1929 1196
rect 2023 1156 2025 1196
rect 2029 1156 2031 1196
rect 2043 1156 2045 1196
rect 2049 1168 2051 1196
rect 2063 1168 2065 1196
rect 2049 1156 2065 1168
rect 2069 1156 2071 1196
rect 2186 1138 2188 1196
rect 2174 1136 2188 1138
rect 2192 1136 2196 1196
rect 2200 1136 2204 1196
rect 2208 1136 2210 1196
rect 2326 1138 2328 1196
rect 2314 1136 2328 1138
rect 2332 1136 2336 1196
rect 2340 1136 2344 1196
rect 2348 1136 2350 1196
rect 2443 1156 2445 1196
rect 2449 1156 2451 1196
rect 2463 1156 2465 1196
rect 2469 1168 2471 1196
rect 2483 1168 2485 1196
rect 2469 1156 2485 1168
rect 2489 1156 2491 1196
rect 2606 1138 2608 1196
rect 2594 1136 2608 1138
rect 2612 1136 2616 1196
rect 2620 1136 2624 1196
rect 2628 1136 2630 1196
rect 2729 1176 2731 1196
rect 2735 1176 2737 1196
rect 2829 1176 2831 1196
rect 2835 1176 2837 1196
rect 2849 1176 2851 1196
rect 2855 1176 2857 1196
rect 2949 1176 2951 1196
rect 2955 1176 2957 1196
rect 2969 1176 2971 1196
rect 2975 1176 2977 1196
rect 3069 1156 3071 1196
rect 3075 1156 3081 1196
rect 3085 1156 3087 1196
rect 3099 1156 3101 1196
rect 3105 1156 3107 1196
rect 3223 1176 3225 1196
rect 3229 1176 3231 1196
rect 3243 1176 3245 1196
rect 3249 1176 3251 1196
rect 3363 1176 3365 1196
rect 3369 1176 3371 1196
rect 3383 1176 3385 1196
rect 3389 1176 3391 1196
rect 3483 1176 3485 1196
rect 3489 1176 3491 1196
rect 3583 1156 3585 1196
rect 3589 1156 3591 1196
rect 3603 1156 3605 1196
rect 3609 1168 3611 1196
rect 3623 1168 3625 1196
rect 3609 1156 3625 1168
rect 3629 1156 3631 1196
rect 3723 1156 3725 1196
rect 3729 1156 3731 1196
rect 3743 1156 3745 1196
rect 3749 1168 3751 1196
rect 3763 1168 3765 1196
rect 3749 1156 3765 1168
rect 3769 1156 3771 1196
rect 3851 1156 3853 1196
rect 3857 1156 3863 1196
rect 3867 1156 3869 1196
rect 3971 1156 3973 1196
rect 3977 1156 3983 1196
rect 3987 1156 3989 1196
rect 4089 1176 4091 1196
rect 4095 1176 4097 1196
rect 4109 1176 4111 1196
rect 4115 1176 4117 1196
rect 4209 1176 4211 1196
rect 4215 1176 4217 1196
rect 4330 1176 4332 1196
rect 4336 1176 4340 1196
rect 4352 1156 4354 1196
rect 4358 1156 4362 1196
rect 4366 1156 4368 1196
rect 4483 1156 4485 1196
rect 4489 1156 4491 1196
rect 4503 1156 4505 1196
rect 4509 1168 4511 1196
rect 4523 1168 4525 1196
rect 4509 1156 4525 1168
rect 4529 1156 4531 1196
rect 4630 1176 4632 1196
rect 4636 1176 4640 1196
rect 4652 1156 4654 1196
rect 4658 1156 4662 1196
rect 4666 1156 4668 1196
rect 4749 1156 4751 1196
rect 4755 1168 4757 1196
rect 4769 1168 4771 1196
rect 4755 1156 4771 1168
rect 4775 1156 4777 1196
rect 4789 1156 4791 1196
rect 4795 1156 4797 1196
rect 4889 1176 4891 1196
rect 4895 1176 4899 1196
rect 4911 1156 4913 1196
rect 4917 1156 4919 1196
rect 5009 1176 5011 1196
rect 5015 1176 5017 1196
rect 5109 1176 5111 1196
rect 5115 1176 5117 1196
rect 5231 1156 5233 1196
rect 5237 1156 5243 1196
rect 5247 1156 5249 1196
rect 5363 1156 5365 1196
rect 5369 1156 5371 1196
rect 5383 1156 5385 1196
rect 5389 1168 5391 1196
rect 5403 1168 5405 1196
rect 5389 1156 5405 1168
rect 5409 1156 5411 1196
rect 5489 1176 5491 1196
rect 5495 1176 5497 1196
rect 5509 1176 5511 1196
rect 5515 1176 5517 1196
rect 5646 1138 5648 1196
rect 5634 1136 5648 1138
rect 5652 1136 5656 1196
rect 5660 1136 5664 1196
rect 5668 1136 5670 1196
rect 5763 1176 5765 1196
rect 5769 1176 5771 1196
rect 94 802 108 804
rect 106 744 108 802
rect 112 744 116 804
rect 120 744 124 804
rect 128 744 130 804
rect 212 744 214 784
rect 218 744 222 784
rect 226 744 228 784
rect 374 802 388 804
rect 240 744 244 764
rect 248 744 250 764
rect 386 744 388 802
rect 392 744 396 804
rect 400 744 404 804
rect 408 744 410 804
rect 654 802 668 804
rect 510 744 512 764
rect 516 744 520 764
rect 532 744 534 784
rect 538 744 542 784
rect 546 744 548 784
rect 666 744 668 802
rect 672 744 676 804
rect 680 744 684 804
rect 688 744 690 804
rect 772 744 774 784
rect 778 744 782 784
rect 786 744 788 784
rect 1074 802 1088 804
rect 800 744 804 764
rect 808 744 810 764
rect 923 744 925 784
rect 929 744 931 784
rect 943 744 945 784
rect 949 772 965 784
rect 949 744 951 772
rect 963 744 965 772
rect 969 744 971 784
rect 1086 744 1088 802
rect 1092 744 1096 804
rect 1100 744 1104 804
rect 1108 744 1110 804
rect 1354 802 1368 804
rect 1189 744 1191 784
rect 1195 772 1211 784
rect 1195 744 1197 772
rect 1209 744 1211 772
rect 1215 744 1217 784
rect 1229 744 1231 784
rect 1235 744 1237 784
rect 1366 744 1368 802
rect 1372 744 1376 804
rect 1380 744 1384 804
rect 1388 744 1390 804
rect 1734 802 1748 804
rect 1469 744 1471 764
rect 1475 744 1477 764
rect 1571 744 1573 784
rect 1577 744 1583 784
rect 1587 744 1589 784
rect 1746 744 1748 802
rect 1752 744 1756 804
rect 1760 744 1764 804
rect 1768 744 1770 804
rect 1874 802 1888 804
rect 1886 744 1888 802
rect 1892 744 1896 804
rect 1900 744 1904 804
rect 1908 744 1910 804
rect 1990 744 1992 804
rect 1996 744 2000 804
rect 2004 744 2008 804
rect 2012 802 2026 804
rect 2012 744 2014 802
rect 2129 744 2131 784
rect 2135 772 2151 784
rect 2135 744 2137 772
rect 2149 744 2151 772
rect 2155 744 2157 784
rect 2169 744 2171 784
rect 2175 744 2177 784
rect 2269 744 2271 784
rect 2275 744 2281 784
rect 2285 744 2287 784
rect 2299 744 2301 784
rect 2305 744 2307 784
rect 2409 744 2411 764
rect 2415 744 2417 764
rect 2531 744 2533 784
rect 2537 744 2543 784
rect 2547 744 2549 784
rect 2643 744 2645 784
rect 2649 764 2661 784
rect 2649 744 2651 764
rect 2663 744 2665 764
rect 2669 744 2671 764
rect 2683 744 2685 764
rect 2689 744 2691 764
rect 2771 744 2773 784
rect 2777 744 2783 784
rect 2787 744 2789 784
rect 2911 744 2913 784
rect 2917 744 2923 784
rect 2927 744 2929 784
rect 3029 744 3031 764
rect 3035 744 3037 764
rect 3143 744 3145 764
rect 3149 744 3151 764
rect 3271 744 3273 784
rect 3277 744 3283 784
rect 3287 744 3289 784
rect 3403 744 3405 764
rect 3409 744 3411 764
rect 3423 744 3425 764
rect 3429 744 3431 764
rect 3523 744 3525 764
rect 3529 744 3531 764
rect 3543 744 3545 764
rect 3549 744 3551 764
rect 3650 744 3652 764
rect 3656 744 3660 764
rect 3672 744 3674 784
rect 3678 744 3682 784
rect 3686 744 3688 784
rect 3783 744 3785 764
rect 3789 744 3791 764
rect 3883 744 3885 784
rect 3889 744 3891 784
rect 3903 744 3905 784
rect 3909 772 3925 784
rect 3909 744 3911 772
rect 3923 744 3925 772
rect 3929 744 3931 784
rect 4011 744 4013 784
rect 4017 744 4023 784
rect 4027 744 4029 784
rect 4143 744 4145 784
rect 4149 744 4151 784
rect 4163 744 4165 784
rect 4169 772 4185 784
rect 4169 744 4171 772
rect 4183 744 4185 772
rect 4189 744 4191 784
rect 4283 744 4285 784
rect 4289 744 4291 784
rect 4303 744 4305 784
rect 4309 772 4325 784
rect 4309 744 4311 772
rect 4323 744 4325 772
rect 4329 744 4331 784
rect 4429 744 4431 764
rect 4435 744 4437 764
rect 4543 744 4545 784
rect 4549 744 4551 784
rect 4563 744 4565 784
rect 4569 772 4585 784
rect 4569 744 4571 772
rect 4583 744 4585 772
rect 4589 744 4591 784
rect 4672 744 4674 784
rect 4678 744 4682 784
rect 4686 744 4688 784
rect 4700 744 4704 764
rect 4708 744 4710 764
rect 4821 744 4823 784
rect 4827 744 4829 784
rect 4841 744 4845 764
rect 4849 744 4851 764
rect 4943 744 4945 784
rect 4949 744 4951 784
rect 4963 744 4965 784
rect 4969 772 4985 784
rect 4969 744 4971 772
rect 4983 744 4985 772
rect 4989 744 4991 784
rect 5072 744 5074 784
rect 5078 744 5082 784
rect 5086 744 5088 784
rect 5100 744 5104 764
rect 5108 744 5110 764
rect 5223 744 5225 784
rect 5229 764 5241 784
rect 5229 744 5231 764
rect 5243 744 5245 764
rect 5249 744 5251 764
rect 5263 744 5265 764
rect 5269 744 5271 764
rect 5383 744 5385 764
rect 5389 744 5391 764
rect 5504 744 5506 784
rect 5510 744 5514 784
rect 5518 744 5520 784
rect 5532 744 5534 784
rect 5538 744 5542 784
rect 5546 744 5548 784
rect 5649 744 5651 784
rect 5655 772 5671 784
rect 5655 744 5657 772
rect 5669 744 5671 772
rect 5675 744 5677 784
rect 5689 744 5691 784
rect 5695 744 5697 784
rect 106 658 108 716
rect 94 656 108 658
rect 112 656 116 716
rect 120 656 124 716
rect 128 656 130 716
rect 250 696 252 716
rect 256 696 260 716
rect 272 676 274 716
rect 278 676 282 716
rect 286 676 288 716
rect 406 658 408 716
rect 394 656 408 658
rect 412 656 416 716
rect 420 656 424 716
rect 428 656 430 716
rect 523 676 525 716
rect 529 676 531 716
rect 543 676 545 716
rect 549 688 551 716
rect 563 688 565 716
rect 549 676 565 688
rect 569 676 571 716
rect 652 676 654 716
rect 658 676 662 716
rect 666 676 668 716
rect 680 696 684 716
rect 688 696 690 716
rect 791 676 793 716
rect 797 676 803 716
rect 807 676 809 716
rect 943 676 945 716
rect 949 676 951 716
rect 963 676 965 716
rect 969 688 971 716
rect 983 688 985 716
rect 969 676 985 688
rect 989 676 991 716
rect 1106 658 1108 716
rect 1094 656 1108 658
rect 1112 656 1116 716
rect 1120 656 1124 716
rect 1128 656 1130 716
rect 1212 676 1214 716
rect 1218 676 1222 716
rect 1226 676 1228 716
rect 1240 696 1244 716
rect 1248 696 1250 716
rect 1370 696 1372 716
rect 1376 696 1380 716
rect 1392 676 1394 716
rect 1398 676 1402 716
rect 1406 676 1408 716
rect 1510 656 1512 716
rect 1516 656 1520 716
rect 1524 656 1528 716
rect 1532 658 1534 716
rect 1663 676 1665 716
rect 1669 676 1671 716
rect 1683 676 1685 716
rect 1689 688 1691 716
rect 1703 688 1705 716
rect 1689 676 1705 688
rect 1709 676 1711 716
rect 1532 656 1546 658
rect 1826 658 1828 716
rect 1814 656 1828 658
rect 1832 656 1836 716
rect 1840 656 1844 716
rect 1848 656 1850 716
rect 1932 676 1934 716
rect 1938 676 1942 716
rect 1946 676 1948 716
rect 1960 696 1964 716
rect 1968 696 1970 716
rect 2083 696 2085 716
rect 2089 696 2091 716
rect 2103 696 2105 716
rect 2109 696 2111 716
rect 2203 676 2205 716
rect 2209 696 2211 716
rect 2223 696 2225 716
rect 2229 696 2231 716
rect 2243 696 2245 716
rect 2249 696 2251 716
rect 2209 676 2221 696
rect 2329 676 2331 716
rect 2335 676 2341 716
rect 2345 676 2347 716
rect 2359 676 2361 716
rect 2365 676 2367 716
rect 2471 676 2473 716
rect 2477 676 2483 716
rect 2487 676 2489 716
rect 2611 676 2613 716
rect 2617 676 2623 716
rect 2627 676 2629 716
rect 2723 696 2725 716
rect 2729 696 2731 716
rect 2743 696 2745 716
rect 2749 696 2751 716
rect 2829 676 2831 716
rect 2835 688 2837 716
rect 2849 688 2851 716
rect 2835 676 2851 688
rect 2855 676 2857 716
rect 2869 676 2871 716
rect 2875 676 2877 716
rect 2991 676 2993 716
rect 2997 676 3003 716
rect 3007 676 3009 716
rect 3092 676 3094 716
rect 3098 676 3102 716
rect 3106 676 3108 716
rect 3120 696 3124 716
rect 3128 696 3130 716
rect 3266 658 3268 716
rect 3254 656 3268 658
rect 3272 656 3276 716
rect 3280 656 3284 716
rect 3288 656 3290 716
rect 3371 676 3373 716
rect 3377 676 3383 716
rect 3387 676 3389 716
rect 3503 676 3505 716
rect 3509 676 3511 716
rect 3523 676 3525 716
rect 3529 688 3531 716
rect 3543 688 3545 716
rect 3529 676 3545 688
rect 3549 676 3551 716
rect 3631 676 3633 716
rect 3637 676 3643 716
rect 3647 676 3649 716
rect 3763 676 3765 716
rect 3769 676 3771 716
rect 3783 676 3785 716
rect 3789 688 3791 716
rect 3803 688 3805 716
rect 3789 676 3805 688
rect 3809 676 3811 716
rect 3889 676 3891 716
rect 3895 688 3897 716
rect 3909 688 3911 716
rect 3895 676 3911 688
rect 3915 676 3917 716
rect 3929 676 3931 716
rect 3935 676 3937 716
rect 4032 676 4034 716
rect 4038 676 4042 716
rect 4046 676 4048 716
rect 4060 696 4064 716
rect 4068 696 4070 716
rect 4189 676 4191 716
rect 4195 688 4197 716
rect 4209 688 4211 716
rect 4195 676 4211 688
rect 4215 676 4217 716
rect 4229 676 4231 716
rect 4235 676 4237 716
rect 4343 696 4345 716
rect 4349 696 4351 716
rect 4450 696 4452 716
rect 4456 696 4460 716
rect 4472 676 4474 716
rect 4478 676 4482 716
rect 4486 676 4488 716
rect 4583 676 4585 716
rect 4589 676 4591 716
rect 4603 676 4605 716
rect 4609 688 4611 716
rect 4623 688 4625 716
rect 4609 676 4625 688
rect 4629 676 4631 716
rect 4723 676 4725 716
rect 4729 676 4731 716
rect 4743 676 4745 716
rect 4749 688 4751 716
rect 4763 688 4765 716
rect 4749 676 4765 688
rect 4769 676 4771 716
rect 4869 676 4871 716
rect 4875 688 4877 716
rect 4889 688 4891 716
rect 4875 676 4891 688
rect 4895 676 4897 716
rect 4909 676 4911 716
rect 4915 676 4917 716
rect 5009 696 5011 716
rect 5015 696 5017 716
rect 5129 696 5131 716
rect 5135 696 5139 716
rect 5151 676 5153 716
rect 5157 676 5159 716
rect 5263 676 5265 716
rect 5269 676 5271 716
rect 5283 676 5285 716
rect 5289 688 5291 716
rect 5303 688 5305 716
rect 5289 676 5305 688
rect 5309 676 5311 716
rect 5389 676 5391 716
rect 5395 688 5397 716
rect 5409 688 5411 716
rect 5395 676 5411 688
rect 5415 676 5417 716
rect 5429 676 5431 716
rect 5435 676 5437 716
rect 5543 676 5545 716
rect 5549 676 5551 716
rect 5563 676 5565 716
rect 5569 688 5571 716
rect 5583 688 5585 716
rect 5569 676 5585 688
rect 5589 676 5591 716
rect 5669 696 5671 716
rect 5675 696 5677 716
rect 5689 696 5691 716
rect 5695 696 5697 716
rect 94 322 108 324
rect 106 264 108 322
rect 112 264 116 324
rect 120 264 124 324
rect 128 264 130 324
rect 534 322 548 324
rect 223 264 225 304
rect 229 264 231 304
rect 243 264 245 304
rect 249 292 265 304
rect 249 264 251 292
rect 263 264 265 292
rect 269 264 271 304
rect 383 264 385 304
rect 389 264 391 304
rect 403 264 405 304
rect 409 292 425 304
rect 409 264 411 292
rect 423 264 425 292
rect 429 264 431 304
rect 546 264 548 322
rect 552 264 556 324
rect 560 264 564 324
rect 568 264 570 324
rect 814 322 828 324
rect 673 264 675 304
rect 679 264 681 304
rect 693 264 695 304
rect 699 264 705 304
rect 709 264 711 304
rect 826 264 828 322
rect 832 264 836 324
rect 840 264 844 324
rect 848 264 850 324
rect 950 264 952 284
rect 956 264 960 284
rect 972 264 974 304
rect 978 264 982 304
rect 986 264 988 304
rect 1070 264 1072 324
rect 1076 264 1080 324
rect 1084 264 1088 324
rect 1092 322 1106 324
rect 1092 264 1094 322
rect 1223 264 1225 304
rect 1229 284 1241 304
rect 1374 322 1388 324
rect 1229 264 1231 284
rect 1243 264 1245 284
rect 1249 264 1251 284
rect 1263 264 1265 284
rect 1269 264 1271 284
rect 1386 264 1388 322
rect 1392 264 1396 324
rect 1400 264 1404 324
rect 1408 264 1410 324
rect 1523 264 1525 284
rect 1529 264 1531 284
rect 1623 264 1625 304
rect 1629 264 1631 304
rect 1643 264 1645 304
rect 1649 292 1665 304
rect 1649 264 1651 292
rect 1663 264 1665 292
rect 1669 264 1671 304
rect 1773 264 1775 304
rect 1779 264 1781 304
rect 1793 264 1795 304
rect 1799 264 1805 304
rect 1809 264 1811 304
rect 1889 264 1891 284
rect 1895 264 1897 284
rect 1909 264 1911 284
rect 1915 264 1917 284
rect 2029 264 2031 284
rect 2035 264 2037 284
rect 2143 264 2145 304
rect 2149 264 2151 304
rect 2163 264 2165 304
rect 2169 292 2185 304
rect 2169 264 2171 292
rect 2183 264 2185 292
rect 2189 264 2191 304
rect 2290 264 2292 284
rect 2296 264 2300 284
rect 2312 264 2314 304
rect 2318 264 2322 304
rect 2326 264 2328 304
rect 2534 322 2548 324
rect 2423 264 2425 284
rect 2429 264 2431 284
rect 2546 264 2548 322
rect 2552 264 2556 324
rect 2560 264 2564 324
rect 2568 264 2570 324
rect 2649 264 2651 304
rect 2655 292 2671 304
rect 2655 264 2657 292
rect 2669 264 2671 292
rect 2675 264 2677 304
rect 2689 264 2691 304
rect 2695 264 2697 304
rect 2803 264 2805 284
rect 2809 264 2811 284
rect 2903 264 2905 284
rect 2909 264 2911 284
rect 2923 264 2925 284
rect 2929 264 2931 284
rect 3009 264 3011 284
rect 3015 264 3017 284
rect 3130 264 3132 284
rect 3136 264 3140 284
rect 3152 264 3154 304
rect 3158 264 3162 304
rect 3166 264 3168 304
rect 3272 264 3274 304
rect 3278 264 3282 304
rect 3286 264 3288 304
rect 3300 264 3304 284
rect 3308 264 3310 284
rect 3423 264 3425 284
rect 3429 264 3431 284
rect 3529 264 3531 304
rect 3535 292 3551 304
rect 3535 264 3537 292
rect 3549 264 3551 292
rect 3555 264 3557 304
rect 3569 264 3571 304
rect 3575 264 3577 304
rect 3672 264 3674 304
rect 3678 264 3682 304
rect 3686 264 3688 304
rect 3834 322 3848 324
rect 3700 264 3704 284
rect 3708 264 3710 284
rect 3846 264 3848 322
rect 3852 264 3856 324
rect 3860 264 3864 324
rect 3868 264 3870 324
rect 4114 322 4128 324
rect 3951 264 3953 304
rect 3957 264 3963 304
rect 3967 264 3969 304
rect 4126 264 4128 322
rect 4132 264 4136 324
rect 4140 264 4144 324
rect 4148 264 4150 324
rect 4243 264 4245 304
rect 4249 264 4251 304
rect 4263 264 4265 304
rect 4269 292 4285 304
rect 4269 264 4271 292
rect 4283 264 4285 292
rect 4289 264 4291 304
rect 4383 264 4385 284
rect 4389 264 4391 284
rect 4491 264 4493 304
rect 4497 264 4503 304
rect 4507 264 4509 304
rect 4603 264 4605 304
rect 4609 264 4611 304
rect 4623 264 4625 304
rect 4629 292 4645 304
rect 4629 264 4631 292
rect 4643 264 4645 292
rect 4649 264 4651 304
rect 4743 264 4745 284
rect 4749 264 4751 284
rect 4843 264 4845 304
rect 4849 264 4851 304
rect 4863 264 4865 304
rect 4869 292 4885 304
rect 4869 264 4871 292
rect 4883 264 4885 292
rect 4889 264 4891 304
rect 4979 292 4991 312
rect 4969 272 4971 292
rect 4975 272 4977 292
rect 4989 272 4991 292
rect 4995 272 5001 312
rect 5005 304 5021 312
rect 5005 272 5007 304
rect 5019 272 5021 304
rect 5025 272 5031 312
rect 5035 272 5037 312
rect 5143 264 5145 304
rect 5149 264 5151 304
rect 5163 264 5165 304
rect 5169 292 5185 304
rect 5169 264 5171 292
rect 5183 264 5185 292
rect 5189 264 5191 304
rect 5289 264 5291 304
rect 5295 292 5311 304
rect 5295 264 5297 292
rect 5309 264 5311 292
rect 5315 264 5317 304
rect 5329 264 5331 304
rect 5335 264 5337 304
rect 5470 264 5472 284
rect 5476 264 5480 284
rect 5492 264 5494 304
rect 5498 264 5502 304
rect 5506 264 5508 304
rect 5589 264 5591 304
rect 5595 292 5611 304
rect 5595 264 5597 292
rect 5609 264 5611 292
rect 5615 264 5617 304
rect 5629 264 5631 304
rect 5635 264 5637 304
rect 5731 264 5733 304
rect 5737 264 5743 304
rect 5747 264 5749 304
rect 106 178 108 236
rect 94 176 108 178
rect 112 176 116 236
rect 120 176 124 236
rect 128 176 130 236
rect 212 196 214 236
rect 218 196 222 236
rect 226 196 228 236
rect 240 216 244 236
rect 248 216 250 236
rect 390 216 392 236
rect 396 216 400 236
rect 412 196 414 236
rect 418 196 422 236
rect 426 196 428 236
rect 523 196 525 236
rect 529 196 531 236
rect 543 196 545 236
rect 549 208 551 236
rect 563 208 565 236
rect 549 196 565 208
rect 569 196 571 236
rect 649 196 651 236
rect 655 208 657 236
rect 669 208 671 236
rect 655 196 671 208
rect 675 196 677 236
rect 689 196 691 236
rect 695 196 697 236
rect 826 178 828 236
rect 814 176 828 178
rect 832 176 836 236
rect 840 176 844 236
rect 848 176 850 236
rect 929 216 931 236
rect 935 216 937 236
rect 1029 196 1031 236
rect 1035 208 1037 236
rect 1049 208 1051 236
rect 1035 196 1051 208
rect 1055 196 1057 236
rect 1069 196 1071 236
rect 1075 196 1077 236
rect 1172 196 1174 236
rect 1178 196 1182 236
rect 1186 196 1188 236
rect 1200 216 1204 236
rect 1208 216 1210 236
rect 1309 216 1311 236
rect 1315 216 1317 236
rect 1329 216 1331 236
rect 1335 216 1337 236
rect 1429 196 1431 236
rect 1435 196 1441 236
rect 1445 196 1447 236
rect 1459 196 1461 236
rect 1465 196 1467 236
rect 1583 216 1585 236
rect 1589 216 1591 236
rect 1683 196 1685 236
rect 1689 196 1691 236
rect 1703 196 1705 236
rect 1709 208 1711 236
rect 1723 208 1725 236
rect 1709 196 1725 208
rect 1729 196 1731 236
rect 1831 196 1833 236
rect 1837 196 1843 236
rect 1847 196 1849 236
rect 1930 176 1932 236
rect 1936 176 1940 236
rect 1944 176 1948 236
rect 1952 178 1954 236
rect 1952 176 1966 178
rect 2126 178 2128 236
rect 2114 176 2128 178
rect 2132 176 2136 236
rect 2140 176 2144 236
rect 2148 176 2150 236
rect 2229 216 2231 236
rect 2235 216 2239 236
rect 2251 196 2253 236
rect 2257 196 2259 236
rect 2371 196 2373 236
rect 2377 196 2383 236
rect 2387 196 2389 236
rect 2469 196 2471 236
rect 2475 196 2481 236
rect 2485 196 2487 236
rect 2499 196 2501 236
rect 2505 196 2507 236
rect 2630 216 2632 236
rect 2636 216 2640 236
rect 2652 196 2654 236
rect 2658 196 2662 236
rect 2666 196 2668 236
rect 2773 196 2775 236
rect 2779 196 2781 236
rect 2793 196 2795 236
rect 2799 196 2805 236
rect 2809 196 2811 236
rect 2911 196 2913 236
rect 2917 196 2923 236
rect 2927 196 2929 236
rect 3051 196 3053 236
rect 3057 196 3063 236
rect 3067 196 3069 236
rect 3186 178 3188 236
rect 3174 176 3188 178
rect 3192 176 3196 236
rect 3200 176 3204 236
rect 3208 176 3210 236
rect 3303 216 3305 236
rect 3309 216 3311 236
rect 3389 196 3391 236
rect 3395 208 3397 236
rect 3409 208 3411 236
rect 3395 196 3411 208
rect 3415 196 3417 236
rect 3429 196 3431 236
rect 3435 196 3437 236
rect 3543 216 3545 236
rect 3549 216 3551 236
rect 3651 196 3653 236
rect 3657 196 3663 236
rect 3667 196 3669 236
rect 3761 196 3763 236
rect 3767 196 3769 236
rect 3781 216 3785 236
rect 3789 216 3791 236
rect 3869 216 3871 236
rect 3875 216 3879 236
rect 3891 196 3893 236
rect 3897 196 3899 236
rect 4011 196 4013 236
rect 4017 196 4023 236
rect 4027 196 4029 236
rect 4129 196 4131 236
rect 4135 196 4141 236
rect 4145 196 4147 236
rect 4159 196 4161 236
rect 4165 196 4167 236
rect 4303 216 4305 236
rect 4309 216 4311 236
rect 4323 216 4325 236
rect 4329 216 4331 236
rect 4411 196 4413 236
rect 4417 196 4423 236
rect 4427 196 4429 236
rect 4566 178 4568 236
rect 4554 176 4568 178
rect 4572 176 4576 236
rect 4580 176 4584 236
rect 4588 176 4590 236
rect 4703 196 4705 236
rect 4709 196 4711 236
rect 4723 196 4725 236
rect 4729 208 4731 236
rect 4743 208 4745 236
rect 4729 196 4745 208
rect 4749 196 4751 236
rect 4831 196 4833 236
rect 4837 196 4843 236
rect 4847 196 4849 236
rect 4963 196 4965 236
rect 4969 196 4971 236
rect 4983 196 4985 236
rect 4989 208 4991 236
rect 5003 208 5005 236
rect 4989 196 5005 208
rect 5009 196 5011 236
rect 5089 216 5091 236
rect 5095 216 5097 236
rect 5109 216 5111 236
rect 5115 216 5117 236
rect 5231 196 5233 236
rect 5237 196 5243 236
rect 5247 196 5249 236
rect 5329 208 5331 228
rect 5335 208 5337 228
rect 5349 208 5351 228
rect 5339 188 5351 208
rect 5355 188 5361 228
rect 5365 196 5367 228
rect 5379 196 5381 228
rect 5365 188 5381 196
rect 5385 188 5391 228
rect 5395 188 5397 228
rect 5489 216 5491 236
rect 5495 216 5497 236
rect 5603 216 5605 236
rect 5609 216 5611 236
rect 5691 196 5693 236
rect 5697 196 5703 236
rect 5707 196 5709 236
<< pdiffusion >>
rect 88 5716 90 5756
rect 94 5716 98 5756
rect 110 5676 112 5756
rect 116 5676 120 5756
rect 124 5676 126 5756
rect 214 5676 216 5756
rect 220 5676 224 5756
rect 228 5676 230 5756
rect 242 5716 246 5756
rect 250 5716 252 5756
rect 383 5676 385 5756
rect 389 5676 391 5756
rect 403 5676 405 5756
rect 409 5688 411 5756
rect 423 5688 425 5756
rect 409 5676 425 5688
rect 429 5684 431 5756
rect 509 5716 511 5756
rect 515 5716 517 5756
rect 529 5716 531 5756
rect 535 5720 537 5756
rect 549 5720 551 5756
rect 535 5716 551 5720
rect 555 5716 557 5756
rect 668 5716 670 5756
rect 674 5716 678 5756
rect 429 5676 443 5684
rect 690 5676 692 5756
rect 696 5676 700 5756
rect 704 5676 706 5756
rect 803 5716 805 5756
rect 809 5716 811 5756
rect 823 5716 825 5756
rect 829 5716 831 5756
rect 923 5676 925 5756
rect 929 5676 931 5756
rect 943 5676 945 5756
rect 949 5688 951 5756
rect 963 5688 965 5756
rect 949 5676 965 5688
rect 969 5684 971 5756
rect 969 5676 983 5684
rect 1069 5676 1071 5756
rect 1075 5676 1079 5756
rect 1083 5676 1085 5756
rect 1233 5677 1235 5756
rect 1221 5676 1235 5677
rect 1239 5677 1241 5756
rect 1253 5677 1255 5756
rect 1239 5676 1255 5677
rect 1259 5676 1265 5756
rect 1269 5676 1271 5756
rect 1359 5676 1361 5756
rect 1365 5676 1367 5756
rect 1379 5716 1383 5756
rect 1387 5716 1391 5756
rect 1403 5716 1405 5756
rect 1409 5716 1411 5756
rect 1503 5716 1505 5756
rect 1509 5720 1511 5756
rect 1523 5720 1525 5756
rect 1509 5716 1525 5720
rect 1529 5716 1531 5756
rect 1543 5716 1545 5756
rect 1549 5716 1551 5756
rect 1663 5676 1665 5756
rect 1669 5676 1671 5756
rect 1683 5676 1685 5756
rect 1689 5688 1691 5756
rect 1703 5688 1705 5756
rect 1689 5676 1705 5688
rect 1709 5684 1711 5756
rect 1803 5716 1805 5756
rect 1809 5720 1811 5756
rect 1823 5720 1825 5756
rect 1809 5716 1825 5720
rect 1829 5716 1831 5756
rect 1843 5716 1845 5756
rect 1849 5716 1851 5756
rect 1929 5716 1931 5756
rect 1935 5716 1937 5756
rect 2048 5716 2050 5756
rect 2054 5716 2058 5756
rect 1709 5676 1723 5684
rect 2070 5676 2072 5756
rect 2076 5676 2080 5756
rect 2084 5676 2086 5756
rect 2174 5676 2176 5756
rect 2180 5676 2184 5756
rect 2188 5676 2190 5756
rect 2202 5716 2206 5756
rect 2210 5716 2212 5756
rect 2309 5684 2311 5756
rect 2297 5676 2311 5684
rect 2315 5688 2317 5756
rect 2329 5688 2331 5756
rect 2315 5676 2331 5688
rect 2335 5676 2337 5756
rect 2349 5676 2351 5756
rect 2355 5676 2357 5756
rect 2463 5716 2465 5756
rect 2469 5716 2471 5756
rect 2483 5716 2485 5756
rect 2489 5716 2491 5756
rect 2583 5716 2585 5756
rect 2589 5720 2591 5756
rect 2603 5720 2605 5756
rect 2589 5716 2605 5720
rect 2609 5716 2611 5756
rect 2623 5716 2625 5756
rect 2629 5716 2631 5756
rect 2723 5716 2725 5756
rect 2729 5720 2731 5756
rect 2743 5720 2745 5756
rect 2729 5716 2745 5720
rect 2749 5716 2751 5756
rect 2763 5716 2765 5756
rect 2769 5716 2771 5756
rect 2849 5716 2851 5756
rect 2855 5716 2857 5756
rect 2869 5716 2871 5756
rect 2875 5716 2877 5756
rect 2983 5716 2985 5756
rect 2989 5716 2991 5756
rect 3088 5716 3090 5756
rect 3094 5716 3098 5756
rect 3110 5676 3112 5756
rect 3116 5676 3120 5756
rect 3124 5676 3126 5756
rect 3239 5676 3241 5756
rect 3245 5676 3247 5756
rect 3259 5716 3263 5756
rect 3267 5716 3271 5756
rect 3283 5716 3285 5756
rect 3289 5716 3291 5756
rect 3395 5676 3397 5756
rect 3401 5676 3405 5756
rect 3409 5676 3411 5756
rect 3503 5716 3505 5756
rect 3509 5720 3511 5756
rect 3523 5720 3525 5756
rect 3509 5716 3525 5720
rect 3529 5716 3531 5756
rect 3543 5716 3545 5756
rect 3549 5716 3551 5756
rect 3663 5716 3665 5756
rect 3669 5716 3671 5756
rect 3763 5716 3765 5756
rect 3769 5716 3771 5756
rect 3849 5716 3851 5756
rect 3855 5716 3857 5756
rect 3954 5676 3956 5756
rect 3960 5676 3964 5756
rect 3968 5676 3970 5756
rect 3982 5716 3986 5756
rect 3990 5716 3992 5756
rect 4089 5716 4091 5756
rect 4095 5716 4097 5756
rect 4149 5676 4151 5756
rect 4155 5736 4157 5756
rect 4169 5736 4173 5756
rect 4177 5736 4181 5756
rect 4185 5736 4187 5756
rect 4199 5736 4201 5756
rect 4155 5676 4164 5736
rect 4190 5716 4201 5736
rect 4205 5716 4209 5756
rect 4213 5716 4215 5756
rect 4253 5716 4255 5756
rect 4259 5716 4261 5756
rect 4273 5716 4275 5756
rect 4279 5716 4287 5756
rect 4291 5716 4293 5756
rect 4305 5716 4307 5756
rect 4311 5716 4321 5756
rect 4325 5716 4327 5756
rect 4339 5716 4341 5756
rect 4332 5676 4341 5716
rect 4345 5676 4347 5756
rect 4468 5716 4470 5756
rect 4474 5716 4478 5756
rect 4490 5676 4492 5756
rect 4496 5676 4500 5756
rect 4504 5676 4506 5756
rect 4603 5676 4605 5756
rect 4609 5676 4611 5756
rect 4623 5676 4625 5756
rect 4629 5676 4631 5756
rect 4643 5676 4645 5756
rect 4649 5676 4651 5756
rect 4663 5676 4665 5756
rect 4669 5676 4671 5756
rect 4683 5676 4685 5756
rect 4689 5676 4691 5756
rect 4703 5676 4705 5756
rect 4709 5676 4711 5756
rect 4723 5676 4725 5756
rect 4729 5676 4731 5756
rect 4743 5676 4745 5756
rect 4749 5676 4751 5756
rect 4843 5716 4845 5756
rect 4849 5716 4851 5756
rect 4948 5716 4950 5756
rect 4954 5716 4958 5756
rect 4970 5676 4972 5756
rect 4976 5676 4980 5756
rect 4984 5676 4986 5756
rect 5083 5716 5085 5756
rect 5089 5716 5091 5756
rect 5103 5716 5105 5756
rect 5109 5716 5111 5756
rect 5189 5716 5191 5756
rect 5195 5716 5197 5756
rect 5209 5716 5211 5756
rect 5215 5716 5217 5756
rect 5314 5676 5316 5756
rect 5320 5676 5324 5756
rect 5328 5676 5330 5756
rect 5342 5716 5346 5756
rect 5350 5716 5352 5756
rect 5449 5716 5451 5756
rect 5455 5716 5457 5756
rect 5549 5716 5551 5756
rect 5555 5716 5557 5756
rect 5569 5716 5571 5756
rect 5575 5716 5577 5756
rect 5669 5716 5671 5756
rect 5675 5716 5677 5756
rect 88 5304 90 5344
rect 94 5304 98 5344
rect 110 5304 112 5384
rect 116 5304 120 5384
rect 124 5304 126 5384
rect 243 5304 245 5344
rect 249 5340 265 5344
rect 249 5304 251 5340
rect 263 5304 265 5340
rect 269 5304 271 5344
rect 283 5304 285 5344
rect 289 5304 291 5344
rect 383 5304 385 5344
rect 389 5340 405 5344
rect 389 5304 391 5340
rect 403 5304 405 5340
rect 409 5304 411 5344
rect 423 5304 425 5344
rect 429 5304 431 5344
rect 523 5304 525 5344
rect 529 5340 545 5344
rect 529 5304 531 5340
rect 543 5304 545 5340
rect 549 5304 551 5344
rect 563 5304 565 5344
rect 569 5304 571 5344
rect 669 5304 671 5344
rect 675 5304 677 5344
rect 689 5304 691 5344
rect 695 5340 711 5344
rect 695 5304 697 5340
rect 709 5304 711 5340
rect 715 5304 717 5344
rect 814 5304 816 5384
rect 820 5304 824 5384
rect 828 5304 830 5384
rect 842 5304 846 5344
rect 850 5304 852 5344
rect 949 5304 951 5344
rect 955 5304 957 5344
rect 969 5304 971 5344
rect 975 5340 991 5344
rect 975 5304 977 5340
rect 989 5304 991 5340
rect 995 5304 997 5344
rect 1103 5304 1105 5384
rect 1109 5304 1111 5384
rect 1123 5304 1125 5384
rect 1129 5372 1145 5384
rect 1129 5304 1131 5372
rect 1143 5304 1145 5372
rect 1149 5376 1163 5384
rect 1149 5304 1151 5376
rect 1229 5304 1231 5344
rect 1235 5304 1237 5344
rect 1249 5304 1251 5344
rect 1255 5340 1271 5344
rect 1255 5304 1257 5340
rect 1269 5304 1271 5340
rect 1275 5304 1277 5344
rect 1389 5304 1391 5384
rect 1395 5304 1399 5384
rect 1403 5304 1405 5384
rect 1523 5304 1525 5344
rect 1529 5340 1545 5344
rect 1529 5304 1531 5340
rect 1543 5304 1545 5340
rect 1549 5304 1551 5344
rect 1563 5304 1565 5344
rect 1569 5304 1571 5344
rect 1654 5304 1656 5384
rect 1660 5304 1664 5384
rect 1668 5304 1670 5384
rect 1682 5304 1686 5344
rect 1690 5304 1692 5344
rect 1803 5304 1805 5344
rect 1809 5340 1825 5344
rect 1809 5304 1811 5340
rect 1823 5304 1825 5340
rect 1829 5304 1831 5344
rect 1843 5304 1845 5344
rect 1849 5304 1851 5344
rect 1943 5304 1945 5344
rect 1949 5340 1965 5344
rect 1949 5304 1951 5340
rect 1963 5304 1965 5340
rect 1969 5304 1971 5344
rect 1983 5304 1985 5344
rect 1989 5304 1991 5344
rect 2069 5304 2071 5344
rect 2075 5304 2077 5344
rect 2089 5304 2091 5344
rect 2095 5304 2097 5344
rect 2223 5304 2225 5344
rect 2229 5304 2231 5344
rect 2319 5304 2321 5384
rect 2325 5304 2327 5384
rect 2339 5304 2343 5344
rect 2347 5304 2351 5344
rect 2363 5304 2365 5344
rect 2369 5304 2371 5344
rect 2454 5304 2456 5384
rect 2460 5304 2464 5384
rect 2468 5304 2470 5384
rect 2482 5304 2486 5344
rect 2490 5304 2492 5344
rect 2623 5304 2625 5344
rect 2629 5340 2645 5344
rect 2629 5304 2631 5340
rect 2643 5304 2645 5340
rect 2649 5304 2651 5344
rect 2663 5304 2665 5344
rect 2669 5304 2671 5344
rect 2763 5304 2765 5344
rect 2769 5340 2785 5344
rect 2769 5304 2771 5340
rect 2783 5304 2785 5340
rect 2789 5304 2791 5344
rect 2803 5304 2805 5344
rect 2809 5304 2811 5344
rect 2894 5304 2896 5384
rect 2900 5304 2904 5384
rect 2908 5304 2910 5384
rect 2922 5304 2926 5344
rect 2930 5304 2932 5344
rect 3029 5304 3031 5344
rect 3035 5304 3037 5344
rect 3129 5304 3131 5344
rect 3135 5304 3137 5344
rect 3149 5304 3151 5344
rect 3155 5304 3157 5344
rect 3269 5304 3271 5344
rect 3275 5304 3277 5344
rect 3289 5304 3291 5344
rect 3295 5340 3311 5344
rect 3295 5304 3297 5340
rect 3309 5304 3311 5340
rect 3315 5304 3317 5344
rect 3409 5304 3411 5344
rect 3415 5304 3417 5344
rect 3429 5304 3431 5344
rect 3435 5304 3437 5344
rect 3529 5304 3531 5384
rect 3535 5304 3541 5384
rect 3545 5383 3561 5384
rect 3545 5304 3547 5383
rect 3559 5304 3561 5383
rect 3565 5383 3579 5384
rect 3565 5304 3567 5383
rect 3683 5304 3685 5344
rect 3689 5340 3705 5344
rect 3689 5304 3691 5340
rect 3703 5304 3705 5340
rect 3709 5304 3711 5344
rect 3723 5304 3725 5344
rect 3729 5304 3731 5344
rect 3823 5304 3825 5384
rect 3829 5304 3831 5384
rect 3843 5304 3845 5384
rect 3849 5372 3865 5384
rect 3849 5304 3851 5372
rect 3863 5304 3865 5372
rect 3869 5376 3883 5384
rect 3869 5304 3871 5376
rect 3949 5304 3951 5344
rect 3955 5304 3957 5344
rect 3969 5304 3971 5344
rect 3975 5304 3977 5344
rect 4088 5304 4090 5344
rect 4094 5304 4098 5344
rect 4110 5304 4112 5384
rect 4116 5304 4120 5384
rect 4124 5304 4126 5384
rect 4477 5376 4491 5384
rect 4223 5304 4225 5344
rect 4229 5304 4231 5344
rect 4243 5304 4245 5344
rect 4249 5304 4251 5344
rect 4343 5304 4345 5344
rect 4349 5340 4365 5344
rect 4349 5304 4351 5340
rect 4363 5304 4365 5340
rect 4369 5304 4371 5344
rect 4383 5304 4385 5344
rect 4389 5304 4391 5344
rect 4489 5304 4491 5376
rect 4495 5372 4511 5384
rect 4495 5304 4497 5372
rect 4509 5304 4511 5372
rect 4515 5304 4517 5384
rect 4529 5304 4531 5384
rect 4535 5304 4537 5384
rect 4629 5304 4631 5344
rect 4635 5304 4637 5344
rect 4734 5304 4736 5384
rect 4740 5304 4744 5384
rect 4748 5304 4750 5384
rect 4762 5304 4766 5344
rect 4770 5304 4772 5344
rect 4829 5304 4831 5384
rect 4835 5324 4844 5384
rect 5012 5344 5021 5384
rect 4870 5324 4881 5344
rect 4835 5304 4837 5324
rect 4849 5304 4853 5324
rect 4857 5304 4861 5324
rect 4865 5304 4867 5324
rect 4879 5304 4881 5324
rect 4885 5304 4889 5344
rect 4893 5304 4895 5344
rect 4933 5304 4935 5344
rect 4939 5304 4941 5344
rect 4953 5304 4955 5344
rect 4959 5304 4967 5344
rect 4971 5304 4973 5344
rect 4985 5304 4987 5344
rect 4991 5304 5001 5344
rect 5005 5304 5007 5344
rect 5019 5304 5021 5344
rect 5025 5304 5027 5384
rect 5109 5304 5111 5344
rect 5115 5304 5117 5344
rect 5169 5304 5171 5384
rect 5175 5324 5184 5384
rect 5352 5344 5361 5384
rect 5210 5324 5221 5344
rect 5175 5304 5177 5324
rect 5189 5304 5193 5324
rect 5197 5304 5201 5324
rect 5205 5304 5207 5324
rect 5219 5304 5221 5324
rect 5225 5304 5229 5344
rect 5233 5304 5235 5344
rect 5273 5304 5275 5344
rect 5279 5304 5281 5344
rect 5293 5304 5295 5344
rect 5299 5304 5307 5344
rect 5311 5304 5313 5344
rect 5325 5304 5327 5344
rect 5331 5304 5341 5344
rect 5345 5304 5347 5344
rect 5359 5304 5361 5344
rect 5365 5304 5367 5384
rect 5454 5304 5456 5384
rect 5460 5304 5464 5384
rect 5468 5304 5470 5384
rect 5482 5304 5486 5344
rect 5490 5304 5492 5344
rect 5609 5304 5611 5344
rect 5615 5304 5617 5344
rect 5629 5304 5631 5344
rect 5635 5304 5637 5344
rect 5729 5304 5731 5344
rect 5735 5304 5737 5344
rect 5749 5304 5751 5344
rect 5755 5304 5757 5344
rect 83 5236 85 5276
rect 89 5240 91 5276
rect 103 5240 105 5276
rect 89 5236 105 5240
rect 109 5236 111 5276
rect 123 5236 125 5276
rect 129 5236 131 5276
rect 209 5204 211 5276
rect 197 5196 211 5204
rect 215 5208 217 5276
rect 229 5208 231 5276
rect 215 5196 231 5208
rect 235 5196 237 5276
rect 249 5196 251 5276
rect 255 5196 257 5276
rect 349 5236 351 5276
rect 355 5236 357 5276
rect 463 5236 465 5276
rect 469 5240 471 5276
rect 483 5240 485 5276
rect 469 5236 485 5240
rect 489 5236 491 5276
rect 503 5236 505 5276
rect 509 5236 511 5276
rect 589 5204 591 5276
rect 577 5196 591 5204
rect 595 5208 597 5276
rect 609 5208 611 5276
rect 595 5196 611 5208
rect 615 5196 617 5276
rect 629 5196 631 5276
rect 635 5196 637 5276
rect 743 5196 745 5276
rect 749 5196 751 5276
rect 763 5196 765 5276
rect 769 5208 771 5276
rect 783 5208 785 5276
rect 769 5196 785 5208
rect 789 5204 791 5276
rect 869 5236 871 5276
rect 875 5236 877 5276
rect 889 5236 891 5276
rect 895 5240 897 5276
rect 909 5240 911 5276
rect 895 5236 911 5240
rect 915 5236 917 5276
rect 1023 5236 1025 5276
rect 1029 5240 1031 5276
rect 1043 5240 1045 5276
rect 1029 5236 1045 5240
rect 1049 5236 1051 5276
rect 1063 5236 1065 5276
rect 1069 5236 1071 5276
rect 1149 5236 1151 5276
rect 1155 5236 1157 5276
rect 1263 5236 1265 5276
rect 1269 5240 1271 5276
rect 1283 5240 1285 5276
rect 1269 5236 1285 5240
rect 1289 5236 1291 5276
rect 1303 5236 1305 5276
rect 1309 5236 1311 5276
rect 1428 5236 1430 5276
rect 1434 5236 1438 5276
rect 789 5196 803 5204
rect 1450 5196 1452 5276
rect 1456 5196 1460 5276
rect 1464 5196 1466 5276
rect 1563 5236 1565 5276
rect 1569 5236 1571 5276
rect 1668 5236 1670 5276
rect 1674 5236 1678 5276
rect 1690 5196 1692 5276
rect 1696 5196 1700 5276
rect 1704 5196 1706 5276
rect 1819 5208 1821 5268
rect 1825 5264 1841 5268
rect 1825 5212 1827 5264
rect 1839 5212 1841 5264
rect 1825 5208 1841 5212
rect 1845 5208 1847 5268
rect 1883 5218 1885 5276
rect 1871 5216 1885 5218
rect 1889 5264 1905 5276
rect 1889 5216 1891 5264
rect 1903 5216 1905 5264
rect 1909 5216 1911 5276
rect 1923 5216 1925 5276
rect 1929 5216 1931 5276
rect 1943 5216 1945 5276
rect 1949 5216 1951 5276
rect 2043 5196 2045 5276
rect 2049 5264 2065 5276
rect 2049 5196 2051 5264
rect 2063 5196 2065 5264
rect 2069 5198 2071 5276
rect 2083 5198 2085 5276
rect 2069 5196 2085 5198
rect 2089 5210 2091 5276
rect 2103 5210 2105 5276
rect 2089 5196 2105 5210
rect 2109 5198 2111 5276
rect 2189 5236 2191 5276
rect 2195 5236 2197 5276
rect 2209 5236 2211 5276
rect 2215 5236 2217 5276
rect 2323 5236 2325 5276
rect 2329 5240 2331 5276
rect 2343 5240 2345 5276
rect 2329 5236 2345 5240
rect 2349 5236 2351 5276
rect 2363 5236 2365 5276
rect 2369 5236 2371 5276
rect 2109 5196 2123 5198
rect 2463 5196 2465 5276
rect 2469 5196 2471 5276
rect 2483 5196 2485 5276
rect 2489 5208 2491 5276
rect 2503 5208 2505 5276
rect 2489 5196 2505 5208
rect 2509 5204 2511 5276
rect 2603 5236 2605 5276
rect 2609 5236 2611 5276
rect 2708 5236 2710 5276
rect 2714 5236 2718 5276
rect 2509 5196 2523 5204
rect 2730 5196 2732 5276
rect 2736 5196 2740 5276
rect 2744 5196 2746 5276
rect 2868 5236 2870 5276
rect 2874 5236 2878 5276
rect 2890 5196 2892 5276
rect 2896 5196 2900 5276
rect 2904 5196 2906 5276
rect 2999 5196 3001 5276
rect 3005 5196 3007 5276
rect 3019 5236 3023 5276
rect 3027 5236 3031 5276
rect 3043 5236 3045 5276
rect 3049 5236 3051 5276
rect 3129 5196 3131 5276
rect 3135 5196 3139 5276
rect 3143 5196 3145 5276
rect 3283 5236 3285 5276
rect 3289 5236 3291 5276
rect 3395 5196 3397 5276
rect 3401 5196 3405 5276
rect 3409 5196 3411 5276
rect 3528 5236 3530 5276
rect 3534 5236 3538 5276
rect 3550 5196 3552 5276
rect 3556 5196 3560 5276
rect 3564 5196 3566 5276
rect 3649 5236 3651 5276
rect 3655 5236 3657 5276
rect 3669 5236 3671 5276
rect 3675 5236 3677 5276
rect 3783 5236 3785 5276
rect 3789 5236 3791 5276
rect 3803 5236 3805 5276
rect 3809 5236 3811 5276
rect 3923 5236 3925 5276
rect 3929 5236 3931 5276
rect 3943 5236 3945 5276
rect 3949 5236 3951 5276
rect 4029 5236 4031 5276
rect 4035 5236 4037 5276
rect 4049 5236 4051 5276
rect 4055 5240 4057 5276
rect 4069 5240 4071 5276
rect 4055 5236 4071 5240
rect 4075 5236 4077 5276
rect 4188 5236 4190 5276
rect 4194 5236 4198 5276
rect 4210 5196 4212 5276
rect 4216 5196 4220 5276
rect 4224 5196 4226 5276
rect 4334 5196 4336 5276
rect 4340 5196 4344 5276
rect 4348 5196 4350 5276
rect 4362 5236 4366 5276
rect 4370 5236 4372 5276
rect 4469 5236 4471 5276
rect 4475 5236 4477 5276
rect 4583 5236 4585 5276
rect 4589 5240 4591 5276
rect 4603 5240 4605 5276
rect 4589 5236 4605 5240
rect 4609 5236 4611 5276
rect 4623 5236 4625 5276
rect 4629 5236 4631 5276
rect 4709 5204 4711 5276
rect 4697 5196 4711 5204
rect 4715 5208 4717 5276
rect 4729 5208 4731 5276
rect 4715 5196 4731 5208
rect 4735 5196 4737 5276
rect 4749 5196 4751 5276
rect 4755 5196 4757 5276
rect 4849 5196 4851 5276
rect 4855 5196 4859 5276
rect 4863 5196 4865 5276
rect 4929 5196 4931 5276
rect 4935 5256 4937 5276
rect 4949 5256 4953 5276
rect 4957 5256 4961 5276
rect 4965 5256 4967 5276
rect 4979 5256 4981 5276
rect 4935 5196 4944 5256
rect 4970 5236 4981 5256
rect 4985 5236 4989 5276
rect 4993 5236 4995 5276
rect 5033 5236 5035 5276
rect 5039 5236 5041 5276
rect 5053 5236 5055 5276
rect 5059 5236 5067 5276
rect 5071 5236 5073 5276
rect 5085 5236 5087 5276
rect 5091 5236 5101 5276
rect 5105 5236 5107 5276
rect 5119 5236 5121 5276
rect 5112 5196 5121 5236
rect 5125 5196 5127 5276
rect 5214 5196 5216 5276
rect 5220 5196 5224 5276
rect 5228 5196 5230 5276
rect 5242 5236 5246 5276
rect 5250 5236 5252 5276
rect 5349 5236 5351 5276
rect 5355 5236 5357 5276
rect 5454 5196 5456 5276
rect 5460 5196 5464 5276
rect 5468 5196 5470 5276
rect 5482 5236 5486 5276
rect 5490 5236 5492 5276
rect 5603 5236 5605 5276
rect 5609 5236 5611 5276
rect 5623 5236 5625 5276
rect 5629 5236 5631 5276
rect 5709 5236 5711 5276
rect 5715 5236 5717 5276
rect 5729 5236 5731 5276
rect 5735 5236 5737 5276
rect 88 4824 90 4864
rect 94 4824 98 4864
rect 110 4824 112 4904
rect 116 4824 120 4904
rect 124 4824 126 4904
rect 223 4824 225 4864
rect 229 4860 245 4864
rect 229 4824 231 4860
rect 243 4824 245 4860
rect 249 4824 251 4864
rect 263 4824 265 4864
rect 269 4824 271 4864
rect 349 4824 351 4864
rect 355 4824 357 4864
rect 369 4824 371 4864
rect 375 4860 391 4864
rect 375 4824 377 4860
rect 389 4824 391 4860
rect 395 4824 397 4864
rect 494 4824 496 4904
rect 500 4824 504 4904
rect 508 4824 510 4904
rect 522 4824 526 4864
rect 530 4824 532 4864
rect 643 4824 645 4864
rect 649 4824 651 4864
rect 663 4824 665 4864
rect 669 4824 671 4864
rect 768 4824 770 4864
rect 774 4824 778 4864
rect 790 4824 792 4904
rect 796 4824 800 4904
rect 804 4824 806 4904
rect 908 4824 910 4864
rect 914 4824 918 4864
rect 930 4824 932 4904
rect 936 4824 940 4904
rect 944 4824 946 4904
rect 1043 4824 1045 4904
rect 1049 4824 1051 4904
rect 1063 4824 1065 4904
rect 1069 4892 1085 4904
rect 1069 4824 1071 4892
rect 1083 4824 1085 4892
rect 1089 4896 1103 4904
rect 1089 4824 1091 4896
rect 1188 4824 1190 4864
rect 1194 4824 1198 4864
rect 1210 4824 1212 4904
rect 1216 4824 1220 4904
rect 1224 4824 1226 4904
rect 1323 4824 1325 4864
rect 1329 4824 1331 4864
rect 1423 4824 1425 4864
rect 1429 4824 1431 4864
rect 1443 4824 1445 4864
rect 1449 4824 1451 4864
rect 1563 4824 1565 4864
rect 1569 4860 1585 4864
rect 1569 4824 1571 4860
rect 1583 4824 1585 4860
rect 1589 4824 1591 4864
rect 1603 4824 1605 4864
rect 1609 4824 1611 4864
rect 1708 4824 1710 4864
rect 1714 4824 1718 4864
rect 1730 4824 1732 4904
rect 1736 4824 1740 4904
rect 1744 4824 1746 4904
rect 1817 4896 1831 4904
rect 1829 4824 1831 4896
rect 1835 4892 1851 4904
rect 1835 4824 1837 4892
rect 1849 4824 1851 4892
rect 1855 4824 1857 4904
rect 1869 4824 1871 4904
rect 1875 4824 1877 4904
rect 1969 4824 1971 4864
rect 1975 4824 1977 4864
rect 1989 4824 1991 4864
rect 1995 4824 1997 4864
rect 2103 4824 2105 4904
rect 2109 4824 2111 4904
rect 2123 4824 2125 4904
rect 2129 4892 2145 4904
rect 2129 4824 2131 4892
rect 2143 4824 2145 4892
rect 2149 4896 2163 4904
rect 2149 4824 2151 4896
rect 2263 4824 2265 4864
rect 2269 4824 2271 4864
rect 2368 4824 2370 4864
rect 2374 4824 2378 4864
rect 2390 4824 2392 4904
rect 2396 4824 2400 4904
rect 2404 4824 2406 4904
rect 2503 4824 2505 4864
rect 2509 4860 2525 4864
rect 2509 4824 2511 4860
rect 2523 4824 2525 4860
rect 2529 4824 2531 4864
rect 2543 4824 2545 4864
rect 2549 4824 2551 4864
rect 2643 4824 2645 4864
rect 2649 4824 2651 4864
rect 2763 4824 2765 4864
rect 2769 4824 2771 4864
rect 2783 4824 2785 4864
rect 2789 4824 2791 4864
rect 2869 4824 2871 4864
rect 2875 4824 2877 4864
rect 2969 4824 2971 4864
rect 2975 4824 2977 4864
rect 2989 4824 2991 4864
rect 2995 4860 3011 4864
rect 2995 4824 2997 4860
rect 3009 4824 3011 4860
rect 3015 4824 3017 4864
rect 3128 4824 3130 4864
rect 3134 4824 3138 4864
rect 3150 4824 3152 4904
rect 3156 4824 3160 4904
rect 3164 4824 3166 4904
rect 3268 4824 3270 4864
rect 3274 4824 3278 4864
rect 3290 4824 3292 4904
rect 3296 4824 3300 4904
rect 3304 4824 3306 4904
rect 3403 4824 3405 4904
rect 3409 4824 3411 4904
rect 3423 4824 3425 4904
rect 3429 4892 3445 4904
rect 3429 4824 3431 4892
rect 3443 4824 3445 4892
rect 3449 4896 3463 4904
rect 3449 4824 3451 4896
rect 3529 4824 3531 4904
rect 3535 4824 3541 4904
rect 3545 4903 3561 4904
rect 3545 4824 3547 4903
rect 3559 4824 3561 4903
rect 3565 4903 3579 4904
rect 3565 4824 3567 4903
rect 3695 4824 3697 4904
rect 3701 4824 3705 4904
rect 3709 4824 3711 4904
rect 3803 4824 3805 4864
rect 3809 4860 3825 4864
rect 3809 4824 3811 4860
rect 3823 4824 3825 4860
rect 3829 4824 3831 4864
rect 3843 4824 3845 4864
rect 3849 4824 3851 4864
rect 3943 4824 3945 4864
rect 3949 4824 3951 4864
rect 4029 4824 4031 4864
rect 4035 4824 4037 4864
rect 4049 4824 4051 4864
rect 4055 4860 4071 4864
rect 4055 4824 4057 4860
rect 4069 4824 4071 4860
rect 4075 4824 4077 4864
rect 4169 4824 4171 4864
rect 4175 4824 4177 4864
rect 4189 4824 4191 4864
rect 4195 4860 4211 4864
rect 4195 4824 4197 4860
rect 4209 4824 4211 4860
rect 4215 4824 4217 4864
rect 4319 4824 4321 4904
rect 4325 4824 4327 4904
rect 4339 4824 4343 4864
rect 4347 4824 4351 4864
rect 4363 4824 4365 4864
rect 4369 4824 4371 4864
rect 4469 4824 4471 4904
rect 4475 4824 4481 4904
rect 4485 4903 4501 4904
rect 4485 4824 4487 4903
rect 4499 4824 4501 4903
rect 4505 4903 4519 4904
rect 4505 4824 4507 4903
rect 4609 4824 4611 4904
rect 4615 4824 4619 4904
rect 4623 4824 4625 4904
rect 4748 4824 4750 4864
rect 4754 4824 4758 4864
rect 4770 4824 4772 4904
rect 4776 4824 4780 4904
rect 4784 4824 4786 4904
rect 4829 4824 4831 4904
rect 4835 4844 4844 4904
rect 5012 4864 5021 4904
rect 4870 4844 4881 4864
rect 4835 4824 4837 4844
rect 4849 4824 4853 4844
rect 4857 4824 4861 4844
rect 4865 4824 4867 4844
rect 4879 4824 4881 4844
rect 4885 4824 4889 4864
rect 4893 4824 4895 4864
rect 4933 4824 4935 4864
rect 4939 4824 4941 4864
rect 4953 4824 4955 4864
rect 4959 4824 4967 4864
rect 4971 4824 4973 4864
rect 4985 4824 4987 4864
rect 4991 4824 5001 4864
rect 5005 4824 5007 4864
rect 5019 4824 5021 4864
rect 5025 4824 5027 4904
rect 5114 4824 5116 4904
rect 5120 4824 5124 4904
rect 5128 4824 5130 4904
rect 5142 4824 5146 4864
rect 5150 4824 5152 4864
rect 5209 4824 5211 4904
rect 5215 4844 5224 4904
rect 5392 4864 5401 4904
rect 5250 4844 5261 4864
rect 5215 4824 5217 4844
rect 5229 4824 5233 4844
rect 5237 4824 5241 4844
rect 5245 4824 5247 4844
rect 5259 4824 5261 4844
rect 5265 4824 5269 4864
rect 5273 4824 5275 4864
rect 5313 4824 5315 4864
rect 5319 4824 5321 4864
rect 5333 4824 5335 4864
rect 5339 4824 5347 4864
rect 5351 4824 5353 4864
rect 5365 4824 5367 4864
rect 5371 4824 5381 4864
rect 5385 4824 5387 4864
rect 5399 4824 5401 4864
rect 5405 4824 5407 4904
rect 5503 4824 5505 4864
rect 5509 4824 5511 4864
rect 5523 4824 5525 4864
rect 5529 4824 5531 4864
rect 5609 4824 5611 4864
rect 5615 4824 5617 4864
rect 5629 4824 5631 4864
rect 5635 4824 5637 4864
rect 5749 4824 5751 4864
rect 5755 4824 5757 4864
rect 5769 4824 5771 4864
rect 5775 4824 5777 4864
rect 83 4716 85 4796
rect 89 4716 91 4796
rect 103 4716 105 4796
rect 109 4728 111 4796
rect 123 4728 125 4796
rect 109 4716 125 4728
rect 129 4724 131 4796
rect 223 4756 225 4796
rect 229 4760 231 4796
rect 243 4760 245 4796
rect 229 4756 245 4760
rect 249 4756 251 4796
rect 263 4756 265 4796
rect 269 4756 271 4796
rect 129 4716 143 4724
rect 349 4724 351 4796
rect 337 4716 351 4724
rect 355 4728 357 4796
rect 369 4728 371 4796
rect 355 4716 371 4728
rect 375 4716 377 4796
rect 389 4716 391 4796
rect 395 4716 397 4796
rect 489 4756 491 4796
rect 495 4756 497 4796
rect 509 4756 511 4796
rect 515 4756 517 4796
rect 623 4756 625 4796
rect 629 4760 631 4796
rect 643 4760 645 4796
rect 629 4756 645 4760
rect 649 4756 651 4796
rect 663 4756 665 4796
rect 669 4756 671 4796
rect 783 4756 785 4796
rect 789 4760 791 4796
rect 803 4760 805 4796
rect 789 4756 805 4760
rect 809 4756 811 4796
rect 823 4756 825 4796
rect 829 4756 831 4796
rect 909 4756 911 4796
rect 915 4756 917 4796
rect 1009 4756 1011 4796
rect 1015 4756 1017 4796
rect 1123 4756 1125 4796
rect 1129 4756 1131 4796
rect 1228 4756 1230 4796
rect 1234 4756 1238 4796
rect 1250 4716 1252 4796
rect 1256 4716 1260 4796
rect 1264 4716 1266 4796
rect 1354 4716 1356 4796
rect 1360 4716 1364 4796
rect 1368 4716 1370 4796
rect 1382 4756 1386 4796
rect 1390 4756 1392 4796
rect 1489 4756 1491 4796
rect 1495 4756 1497 4796
rect 1589 4756 1591 4796
rect 1595 4756 1597 4796
rect 1609 4756 1611 4796
rect 1615 4760 1617 4796
rect 1629 4760 1631 4796
rect 1615 4756 1631 4760
rect 1635 4756 1637 4796
rect 1748 4756 1750 4796
rect 1754 4756 1758 4796
rect 1770 4716 1772 4796
rect 1776 4716 1780 4796
rect 1784 4716 1786 4796
rect 1883 4756 1885 4796
rect 1889 4756 1891 4796
rect 1903 4756 1905 4796
rect 1909 4756 1911 4796
rect 1994 4716 1996 4796
rect 2000 4716 2004 4796
rect 2008 4716 2010 4796
rect 2022 4756 2026 4796
rect 2030 4756 2032 4796
rect 2143 4756 2145 4796
rect 2149 4760 2151 4796
rect 2163 4760 2165 4796
rect 2149 4756 2165 4760
rect 2169 4756 2171 4796
rect 2183 4756 2185 4796
rect 2189 4756 2191 4796
rect 2281 4716 2283 4796
rect 2287 4716 2289 4796
rect 2301 4756 2305 4796
rect 2309 4756 2311 4796
rect 2389 4756 2391 4796
rect 2395 4756 2397 4796
rect 2409 4756 2411 4796
rect 2415 4756 2417 4796
rect 2509 4756 2511 4796
rect 2515 4756 2517 4796
rect 2529 4756 2531 4796
rect 2535 4756 2537 4796
rect 2641 4716 2643 4796
rect 2647 4716 2649 4796
rect 2661 4756 2665 4796
rect 2669 4756 2671 4796
rect 2749 4756 2751 4796
rect 2755 4756 2757 4796
rect 2769 4756 2771 4796
rect 2775 4760 2777 4796
rect 2789 4760 2791 4796
rect 2775 4756 2791 4760
rect 2795 4756 2797 4796
rect 2915 4716 2917 4796
rect 2921 4716 2925 4796
rect 2929 4716 2931 4796
rect 3029 4716 3031 4796
rect 3035 4716 3041 4796
rect 3045 4716 3047 4796
rect 3069 4716 3071 4796
rect 3075 4716 3081 4796
rect 3085 4716 3087 4796
rect 3203 4756 3205 4796
rect 3209 4756 3211 4796
rect 3223 4756 3225 4796
rect 3229 4756 3231 4796
rect 3323 4756 3325 4796
rect 3329 4760 3331 4796
rect 3343 4760 3345 4796
rect 3329 4756 3345 4760
rect 3349 4756 3351 4796
rect 3363 4756 3365 4796
rect 3369 4756 3371 4796
rect 3463 4716 3465 4796
rect 3469 4716 3471 4796
rect 3483 4716 3485 4796
rect 3489 4728 3491 4796
rect 3503 4728 3505 4796
rect 3489 4716 3505 4728
rect 3509 4724 3511 4796
rect 3603 4756 3605 4796
rect 3609 4760 3611 4796
rect 3623 4760 3625 4796
rect 3609 4756 3625 4760
rect 3629 4756 3631 4796
rect 3643 4756 3645 4796
rect 3649 4756 3651 4796
rect 3509 4716 3523 4724
rect 3743 4716 3745 4796
rect 3749 4716 3751 4796
rect 3763 4716 3765 4796
rect 3769 4728 3771 4796
rect 3783 4728 3785 4796
rect 3769 4716 3785 4728
rect 3789 4724 3791 4796
rect 3869 4756 3871 4796
rect 3875 4756 3877 4796
rect 3889 4756 3891 4796
rect 3895 4760 3897 4796
rect 3909 4760 3911 4796
rect 3895 4756 3911 4760
rect 3915 4756 3917 4796
rect 4009 4756 4011 4796
rect 4015 4756 4017 4796
rect 4029 4756 4031 4796
rect 4035 4760 4037 4796
rect 4049 4760 4051 4796
rect 4035 4756 4051 4760
rect 4055 4756 4057 4796
rect 4149 4756 4151 4796
rect 4155 4756 4157 4796
rect 3789 4716 3803 4724
rect 4259 4716 4261 4796
rect 4265 4716 4267 4796
rect 4279 4756 4283 4796
rect 4287 4756 4291 4796
rect 4303 4756 4305 4796
rect 4309 4756 4311 4796
rect 4423 4756 4425 4796
rect 4429 4760 4431 4796
rect 4443 4760 4445 4796
rect 4429 4756 4445 4760
rect 4449 4756 4451 4796
rect 4463 4756 4465 4796
rect 4469 4756 4471 4796
rect 4549 4756 4551 4796
rect 4555 4756 4557 4796
rect 4569 4756 4571 4796
rect 4575 4760 4577 4796
rect 4589 4760 4591 4796
rect 4575 4756 4591 4760
rect 4595 4756 4597 4796
rect 4689 4756 4691 4796
rect 4695 4756 4697 4796
rect 4749 4716 4751 4796
rect 4755 4776 4757 4796
rect 4769 4776 4773 4796
rect 4777 4776 4781 4796
rect 4785 4776 4787 4796
rect 4799 4776 4801 4796
rect 4755 4716 4764 4776
rect 4790 4756 4801 4776
rect 4805 4756 4809 4796
rect 4813 4756 4815 4796
rect 4853 4756 4855 4796
rect 4859 4756 4861 4796
rect 4873 4756 4875 4796
rect 4879 4756 4887 4796
rect 4891 4756 4893 4796
rect 4905 4756 4907 4796
rect 4911 4756 4921 4796
rect 4925 4756 4927 4796
rect 4939 4756 4941 4796
rect 4932 4716 4941 4756
rect 4945 4716 4947 4796
rect 5034 4716 5036 4796
rect 5040 4716 5044 4796
rect 5048 4716 5050 4796
rect 5062 4756 5066 4796
rect 5070 4756 5072 4796
rect 5169 4756 5171 4796
rect 5175 4756 5177 4796
rect 5189 4756 5191 4796
rect 5195 4756 5197 4796
rect 5289 4756 5291 4796
rect 5295 4756 5297 4796
rect 5309 4756 5311 4796
rect 5315 4756 5317 4796
rect 5429 4756 5431 4796
rect 5435 4756 5437 4796
rect 5449 4756 5451 4796
rect 5455 4756 5457 4796
rect 5549 4756 5551 4796
rect 5555 4756 5557 4796
rect 5569 4756 5571 4796
rect 5575 4756 5577 4796
rect 5683 4756 5685 4796
rect 5689 4760 5691 4796
rect 5703 4760 5705 4796
rect 5689 4756 5705 4760
rect 5709 4756 5711 4796
rect 5723 4756 5725 4796
rect 5729 4756 5731 4796
rect 88 4344 90 4384
rect 94 4344 98 4384
rect 110 4344 112 4424
rect 116 4344 120 4424
rect 124 4344 126 4424
rect 337 4416 351 4424
rect 223 4344 225 4384
rect 229 4380 245 4384
rect 229 4344 231 4380
rect 243 4344 245 4380
rect 249 4344 251 4384
rect 263 4344 265 4384
rect 269 4344 271 4384
rect 349 4344 351 4416
rect 355 4412 371 4424
rect 355 4344 357 4412
rect 369 4344 371 4412
rect 375 4344 377 4424
rect 389 4344 391 4424
rect 395 4344 397 4424
rect 528 4344 530 4384
rect 534 4344 538 4384
rect 550 4344 552 4424
rect 556 4344 560 4424
rect 564 4344 566 4424
rect 668 4344 670 4384
rect 674 4344 678 4384
rect 690 4344 692 4424
rect 696 4344 700 4424
rect 704 4344 706 4424
rect 877 4416 891 4424
rect 789 4344 791 4384
rect 795 4344 797 4384
rect 889 4344 891 4416
rect 895 4412 911 4424
rect 895 4344 897 4412
rect 909 4344 911 4412
rect 915 4344 917 4424
rect 929 4344 931 4424
rect 935 4344 937 4424
rect 1043 4344 1045 4384
rect 1049 4344 1051 4384
rect 1143 4344 1145 4384
rect 1149 4380 1165 4384
rect 1149 4344 1151 4380
rect 1163 4344 1165 4380
rect 1169 4344 1171 4384
rect 1183 4344 1185 4384
rect 1189 4344 1191 4384
rect 1283 4344 1285 4424
rect 1289 4344 1291 4424
rect 1303 4344 1305 4424
rect 1309 4412 1325 4424
rect 1309 4344 1311 4412
rect 1323 4344 1325 4412
rect 1329 4416 1343 4424
rect 1329 4344 1331 4416
rect 1423 4344 1425 4384
rect 1429 4344 1431 4384
rect 1514 4344 1516 4424
rect 1520 4344 1524 4424
rect 1528 4344 1530 4424
rect 1542 4344 1546 4384
rect 1550 4344 1552 4384
rect 1663 4344 1665 4384
rect 1669 4344 1671 4384
rect 1683 4344 1685 4384
rect 1689 4344 1691 4384
rect 1783 4344 1785 4384
rect 1789 4380 1805 4384
rect 1789 4344 1791 4380
rect 1803 4344 1805 4380
rect 1809 4344 1811 4384
rect 1823 4344 1825 4384
rect 1829 4344 1831 4384
rect 1935 4344 1937 4424
rect 1941 4344 1945 4424
rect 1949 4344 1951 4424
rect 2043 4344 2045 4384
rect 2049 4380 2065 4384
rect 2049 4344 2051 4380
rect 2063 4344 2065 4380
rect 2069 4344 2071 4384
rect 2083 4344 2085 4384
rect 2089 4344 2091 4384
rect 2203 4344 2205 4384
rect 2209 4380 2225 4384
rect 2209 4344 2211 4380
rect 2223 4344 2225 4380
rect 2229 4344 2231 4384
rect 2243 4344 2245 4384
rect 2249 4344 2251 4384
rect 2343 4344 2345 4384
rect 2349 4344 2351 4384
rect 2363 4344 2365 4384
rect 2369 4344 2371 4384
rect 2463 4344 2465 4384
rect 2469 4380 2485 4384
rect 2469 4344 2471 4380
rect 2483 4344 2485 4380
rect 2489 4344 2491 4384
rect 2503 4344 2505 4384
rect 2509 4344 2511 4384
rect 2589 4344 2591 4384
rect 2595 4344 2597 4384
rect 2609 4344 2611 4384
rect 2615 4380 2631 4384
rect 2615 4344 2617 4380
rect 2629 4344 2631 4380
rect 2635 4344 2637 4384
rect 2743 4344 2745 4384
rect 2749 4344 2751 4384
rect 2855 4344 2857 4424
rect 2861 4344 2865 4424
rect 2869 4344 2871 4424
rect 2963 4344 2965 4384
rect 2969 4380 2985 4384
rect 2969 4344 2971 4380
rect 2983 4344 2985 4380
rect 2989 4344 2991 4384
rect 3003 4344 3005 4384
rect 3009 4344 3011 4384
rect 3103 4344 3105 4384
rect 3109 4380 3125 4384
rect 3109 4344 3111 4380
rect 3123 4344 3125 4380
rect 3129 4344 3131 4384
rect 3143 4344 3145 4384
rect 3149 4344 3151 4384
rect 3229 4344 3231 4384
rect 3235 4344 3237 4384
rect 3334 4344 3336 4424
rect 3340 4344 3344 4424
rect 3348 4344 3350 4424
rect 3362 4344 3366 4384
rect 3370 4344 3372 4384
rect 3479 4344 3481 4424
rect 3485 4344 3487 4424
rect 3761 4423 3775 4424
rect 3499 4344 3503 4384
rect 3507 4344 3511 4384
rect 3523 4344 3525 4384
rect 3529 4344 3531 4384
rect 3629 4344 3631 4384
rect 3635 4344 3637 4384
rect 3649 4344 3651 4384
rect 3655 4344 3657 4384
rect 3773 4344 3775 4423
rect 3779 4423 3795 4424
rect 3779 4344 3781 4423
rect 3793 4344 3795 4423
rect 3799 4344 3805 4424
rect 3809 4344 3811 4424
rect 3889 4344 3891 4384
rect 3895 4344 3897 4384
rect 3909 4344 3911 4384
rect 3915 4344 3917 4384
rect 4021 4344 4023 4424
rect 4027 4344 4029 4424
rect 4041 4344 4045 4384
rect 4049 4344 4051 4384
rect 4129 4344 4131 4384
rect 4135 4344 4137 4384
rect 4149 4344 4153 4384
rect 4157 4344 4161 4384
rect 4173 4344 4175 4424
rect 4179 4344 4181 4424
rect 4283 4344 4285 4384
rect 4289 4344 4291 4384
rect 4303 4344 4305 4384
rect 4309 4344 4311 4384
rect 4408 4344 4410 4384
rect 4414 4344 4418 4384
rect 4430 4344 4432 4424
rect 4436 4344 4440 4424
rect 4444 4344 4446 4424
rect 4529 4344 4531 4384
rect 4535 4344 4537 4384
rect 4549 4344 4551 4384
rect 4555 4344 4557 4384
rect 4663 4344 4665 4384
rect 4669 4344 4671 4384
rect 4683 4344 4685 4384
rect 4689 4344 4691 4384
rect 4769 4344 4771 4384
rect 4775 4344 4777 4384
rect 4869 4344 4871 4384
rect 4875 4344 4877 4384
rect 4889 4344 4891 4384
rect 4895 4344 4897 4384
rect 4994 4344 4996 4424
rect 5000 4344 5004 4424
rect 5008 4344 5010 4424
rect 5022 4344 5026 4384
rect 5030 4344 5032 4384
rect 5089 4344 5091 4424
rect 5095 4364 5104 4424
rect 5272 4384 5281 4424
rect 5130 4364 5141 4384
rect 5095 4344 5097 4364
rect 5109 4344 5113 4364
rect 5117 4344 5121 4364
rect 5125 4344 5127 4364
rect 5139 4344 5141 4364
rect 5145 4344 5149 4384
rect 5153 4344 5155 4384
rect 5193 4344 5195 4384
rect 5199 4344 5201 4384
rect 5213 4344 5215 4384
rect 5219 4344 5227 4384
rect 5231 4344 5233 4384
rect 5245 4344 5247 4384
rect 5251 4344 5261 4384
rect 5265 4344 5267 4384
rect 5279 4344 5281 4384
rect 5285 4344 5287 4424
rect 5374 4344 5376 4424
rect 5380 4344 5384 4424
rect 5388 4344 5390 4424
rect 5402 4344 5406 4384
rect 5410 4344 5412 4384
rect 5509 4344 5511 4424
rect 5515 4344 5521 4424
rect 5525 4423 5541 4424
rect 5525 4344 5527 4423
rect 5539 4344 5541 4423
rect 5545 4423 5559 4424
rect 5545 4344 5547 4423
rect 5668 4344 5670 4384
rect 5674 4344 5678 4384
rect 5690 4344 5692 4424
rect 5696 4344 5700 4424
rect 5704 4344 5706 4424
rect 108 4276 110 4316
rect 114 4276 118 4316
rect 130 4236 132 4316
rect 136 4236 140 4316
rect 144 4236 146 4316
rect 248 4276 250 4316
rect 254 4276 258 4316
rect 270 4236 272 4316
rect 276 4236 280 4316
rect 284 4236 286 4316
rect 403 4276 405 4316
rect 409 4280 411 4316
rect 423 4280 425 4316
rect 409 4276 425 4280
rect 429 4276 431 4316
rect 443 4276 445 4316
rect 449 4276 451 4316
rect 543 4276 545 4316
rect 549 4280 551 4316
rect 563 4280 565 4316
rect 549 4276 565 4280
rect 569 4276 571 4316
rect 583 4276 585 4316
rect 589 4276 591 4316
rect 693 4237 695 4316
rect 681 4236 695 4237
rect 699 4237 701 4316
rect 713 4237 715 4316
rect 699 4236 715 4237
rect 719 4236 725 4316
rect 729 4236 731 4316
rect 828 4276 830 4316
rect 834 4276 838 4316
rect 850 4236 852 4316
rect 856 4236 860 4316
rect 864 4236 866 4316
rect 949 4276 951 4316
rect 955 4276 957 4316
rect 1063 4236 1065 4316
rect 1069 4236 1071 4316
rect 1083 4236 1085 4316
rect 1089 4248 1091 4316
rect 1103 4248 1105 4316
rect 1089 4236 1105 4248
rect 1109 4244 1111 4316
rect 1223 4276 1225 4316
rect 1229 4280 1231 4316
rect 1243 4280 1245 4316
rect 1229 4276 1245 4280
rect 1249 4276 1251 4316
rect 1263 4276 1265 4316
rect 1269 4276 1271 4316
rect 1363 4276 1365 4316
rect 1369 4276 1371 4316
rect 1383 4276 1385 4316
rect 1389 4276 1391 4316
rect 1483 4276 1485 4316
rect 1489 4276 1491 4316
rect 1503 4276 1505 4316
rect 1509 4276 1511 4316
rect 1109 4236 1123 4244
rect 1615 4236 1617 4316
rect 1621 4236 1625 4316
rect 1629 4236 1631 4316
rect 1723 4276 1725 4316
rect 1729 4280 1731 4316
rect 1743 4280 1745 4316
rect 1729 4276 1745 4280
rect 1749 4276 1751 4316
rect 1763 4276 1765 4316
rect 1769 4276 1771 4316
rect 1863 4276 1865 4316
rect 1869 4280 1871 4316
rect 1883 4280 1885 4316
rect 1869 4276 1885 4280
rect 1889 4276 1891 4316
rect 1903 4276 1905 4316
rect 1909 4276 1911 4316
rect 1989 4276 1991 4316
rect 1995 4276 1997 4316
rect 2009 4276 2011 4316
rect 2015 4280 2017 4316
rect 2029 4280 2031 4316
rect 2015 4276 2031 4280
rect 2035 4276 2037 4316
rect 2129 4276 2131 4316
rect 2135 4276 2137 4316
rect 2149 4276 2151 4316
rect 2155 4280 2157 4316
rect 2169 4280 2171 4316
rect 2155 4276 2171 4280
rect 2175 4276 2177 4316
rect 2295 4236 2297 4316
rect 2301 4236 2305 4316
rect 2309 4236 2311 4316
rect 2428 4276 2430 4316
rect 2434 4276 2438 4316
rect 2450 4236 2452 4316
rect 2456 4236 2460 4316
rect 2464 4236 2466 4316
rect 2583 4276 2585 4316
rect 2589 4280 2591 4316
rect 2603 4280 2605 4316
rect 2589 4276 2605 4280
rect 2609 4276 2611 4316
rect 2623 4276 2625 4316
rect 2629 4276 2631 4316
rect 2709 4276 2711 4316
rect 2715 4276 2717 4316
rect 2829 4276 2831 4316
rect 2835 4276 2837 4316
rect 2849 4276 2851 4316
rect 2855 4280 2857 4316
rect 2869 4280 2871 4316
rect 2855 4276 2871 4280
rect 2875 4276 2877 4316
rect 2969 4276 2971 4316
rect 2975 4276 2977 4316
rect 2989 4276 2991 4316
rect 2995 4276 2997 4316
rect 3089 4244 3091 4316
rect 3077 4236 3091 4244
rect 3095 4248 3097 4316
rect 3109 4248 3111 4316
rect 3095 4236 3111 4248
rect 3115 4236 3117 4316
rect 3129 4236 3131 4316
rect 3135 4236 3137 4316
rect 3229 4244 3231 4316
rect 3217 4236 3231 4244
rect 3235 4248 3237 4316
rect 3249 4248 3251 4316
rect 3235 4236 3251 4248
rect 3255 4236 3257 4316
rect 3269 4236 3271 4316
rect 3275 4236 3277 4316
rect 3374 4236 3376 4316
rect 3380 4236 3384 4316
rect 3388 4236 3390 4316
rect 3402 4276 3406 4316
rect 3410 4276 3412 4316
rect 3529 4276 3531 4316
rect 3535 4276 3537 4316
rect 3629 4276 3631 4316
rect 3635 4276 3637 4316
rect 3649 4276 3651 4316
rect 3655 4280 3657 4316
rect 3669 4280 3671 4316
rect 3655 4276 3671 4280
rect 3675 4276 3677 4316
rect 3769 4276 3771 4316
rect 3775 4276 3777 4316
rect 3789 4276 3791 4316
rect 3795 4280 3797 4316
rect 3809 4280 3811 4316
rect 3795 4276 3811 4280
rect 3815 4276 3817 4316
rect 3923 4276 3925 4316
rect 3929 4276 3931 4316
rect 3943 4276 3945 4316
rect 3949 4276 3951 4316
rect 4063 4276 4065 4316
rect 4069 4276 4071 4316
rect 4083 4276 4085 4316
rect 4089 4276 4091 4316
rect 4183 4276 4185 4316
rect 4189 4276 4191 4316
rect 4203 4276 4205 4316
rect 4209 4276 4211 4316
rect 4308 4276 4310 4316
rect 4314 4276 4318 4316
rect 4330 4236 4332 4316
rect 4336 4236 4340 4316
rect 4344 4236 4346 4316
rect 4429 4236 4431 4316
rect 4435 4236 4441 4316
rect 4445 4237 4447 4316
rect 4459 4237 4461 4316
rect 4445 4236 4461 4237
rect 4465 4237 4467 4316
rect 4588 4276 4590 4316
rect 4594 4276 4598 4316
rect 4465 4236 4479 4237
rect 4610 4236 4612 4316
rect 4616 4236 4620 4316
rect 4624 4236 4626 4316
rect 4734 4236 4736 4316
rect 4740 4236 4744 4316
rect 4748 4236 4750 4316
rect 4762 4276 4766 4316
rect 4770 4276 4772 4316
rect 4869 4236 4871 4316
rect 4875 4236 4879 4316
rect 4883 4236 4885 4316
rect 4989 4276 4991 4316
rect 4995 4276 4997 4316
rect 5109 4244 5111 4316
rect 5097 4236 5111 4244
rect 5115 4248 5117 4316
rect 5129 4248 5131 4316
rect 5115 4236 5131 4248
rect 5135 4236 5137 4316
rect 5149 4236 5151 4316
rect 5155 4236 5157 4316
rect 5254 4236 5256 4316
rect 5260 4236 5264 4316
rect 5268 4236 5270 4316
rect 5282 4276 5286 4316
rect 5290 4276 5292 4316
rect 5389 4276 5391 4316
rect 5395 4276 5397 4316
rect 5494 4236 5496 4316
rect 5500 4236 5504 4316
rect 5508 4236 5510 4316
rect 5522 4276 5526 4316
rect 5530 4276 5532 4316
rect 5593 4236 5595 4316
rect 5599 4276 5601 4316
rect 5613 4276 5615 4316
rect 5619 4276 5629 4316
rect 5633 4276 5635 4316
rect 5647 4276 5649 4316
rect 5653 4276 5661 4316
rect 5665 4276 5667 4316
rect 5679 4276 5681 4316
rect 5685 4276 5687 4316
rect 5725 4276 5727 4316
rect 5731 4276 5735 4316
rect 5739 4296 5741 4316
rect 5753 4296 5755 4316
rect 5759 4296 5763 4316
rect 5767 4296 5771 4316
rect 5783 4296 5785 4316
rect 5739 4276 5750 4296
rect 5599 4236 5608 4276
rect 5776 4236 5785 4296
rect 5789 4236 5791 4316
rect 83 3864 85 3904
rect 89 3864 91 3904
rect 194 3864 196 3944
rect 200 3864 204 3944
rect 208 3864 210 3944
rect 437 3936 451 3944
rect 222 3864 226 3904
rect 230 3864 232 3904
rect 343 3864 345 3904
rect 349 3864 351 3904
rect 449 3864 451 3936
rect 455 3932 471 3944
rect 455 3864 457 3932
rect 469 3864 471 3932
rect 475 3864 477 3944
rect 489 3864 491 3944
rect 495 3864 497 3944
rect 615 3864 617 3944
rect 621 3864 625 3944
rect 629 3864 631 3944
rect 743 3864 745 3904
rect 749 3864 751 3904
rect 834 3864 836 3944
rect 840 3864 844 3944
rect 848 3864 850 3944
rect 1197 3942 1211 3944
rect 862 3864 866 3904
rect 870 3864 872 3904
rect 969 3864 971 3904
rect 975 3864 977 3904
rect 1069 3864 1071 3904
rect 1075 3864 1077 3904
rect 1089 3864 1091 3904
rect 1095 3900 1111 3904
rect 1095 3864 1097 3900
rect 1109 3864 1111 3900
rect 1115 3864 1117 3904
rect 1209 3864 1211 3942
rect 1215 3930 1231 3944
rect 1215 3864 1217 3930
rect 1229 3864 1231 3930
rect 1235 3942 1251 3944
rect 1235 3864 1237 3942
rect 1249 3864 1251 3942
rect 1255 3876 1257 3944
rect 1269 3876 1271 3944
rect 1255 3864 1271 3876
rect 1275 3864 1277 3944
rect 1389 3864 1391 3904
rect 1395 3864 1397 3904
rect 1409 3864 1411 3904
rect 1415 3864 1417 3904
rect 1523 3864 1525 3904
rect 1529 3864 1531 3904
rect 1635 3864 1637 3944
rect 1641 3864 1645 3944
rect 1649 3864 1651 3944
rect 1743 3864 1745 3904
rect 1749 3864 1751 3904
rect 1829 3864 1831 3904
rect 1835 3864 1837 3904
rect 1849 3864 1851 3904
rect 1855 3900 1871 3904
rect 1855 3864 1857 3900
rect 1869 3864 1871 3900
rect 1875 3864 1877 3904
rect 1988 3864 1990 3904
rect 1994 3864 1998 3904
rect 2010 3864 2012 3944
rect 2016 3864 2020 3944
rect 2024 3864 2026 3944
rect 2143 3864 2145 3904
rect 2149 3900 2165 3904
rect 2149 3864 2151 3900
rect 2163 3864 2165 3900
rect 2169 3864 2171 3904
rect 2183 3864 2185 3904
rect 2189 3864 2191 3904
rect 2269 3864 2271 3904
rect 2275 3864 2277 3904
rect 2289 3864 2291 3904
rect 2295 3900 2311 3904
rect 2295 3864 2297 3900
rect 2309 3864 2311 3900
rect 2315 3864 2317 3904
rect 2428 3864 2430 3904
rect 2434 3864 2438 3904
rect 2450 3864 2452 3944
rect 2456 3864 2460 3944
rect 2464 3864 2466 3944
rect 2563 3864 2565 3904
rect 2569 3864 2571 3904
rect 2583 3864 2585 3904
rect 2589 3864 2591 3904
rect 2669 3864 2671 3904
rect 2675 3864 2677 3904
rect 2689 3864 2691 3904
rect 2695 3864 2697 3904
rect 2789 3864 2791 3904
rect 2795 3864 2797 3904
rect 2809 3864 2811 3904
rect 2815 3900 2831 3904
rect 2815 3864 2817 3900
rect 2829 3864 2831 3900
rect 2835 3864 2837 3904
rect 2929 3864 2931 3904
rect 2935 3864 2937 3904
rect 2949 3864 2951 3904
rect 2955 3900 2971 3904
rect 2955 3864 2957 3900
rect 2969 3864 2971 3900
rect 2975 3864 2977 3904
rect 3083 3864 3085 3904
rect 3089 3864 3091 3904
rect 3183 3864 3185 3904
rect 3189 3900 3205 3904
rect 3189 3864 3191 3900
rect 3203 3864 3205 3900
rect 3209 3864 3211 3904
rect 3223 3864 3225 3904
rect 3229 3864 3231 3904
rect 3323 3864 3325 3904
rect 3329 3864 3331 3904
rect 3428 3864 3430 3904
rect 3434 3864 3438 3904
rect 3450 3864 3452 3944
rect 3456 3864 3460 3944
rect 3464 3864 3466 3944
rect 3681 3943 3695 3944
rect 3549 3864 3551 3904
rect 3555 3864 3557 3904
rect 3569 3864 3571 3904
rect 3575 3864 3577 3904
rect 3693 3864 3695 3943
rect 3699 3943 3715 3944
rect 3699 3864 3701 3943
rect 3713 3864 3715 3943
rect 3719 3864 3725 3944
rect 3729 3864 3731 3944
rect 3829 3864 3831 3904
rect 3835 3864 3837 3904
rect 3849 3864 3851 3904
rect 3855 3864 3857 3904
rect 3968 3864 3970 3904
rect 3974 3864 3978 3904
rect 3990 3864 3992 3944
rect 3996 3864 4000 3944
rect 4004 3864 4006 3944
rect 4103 3864 4105 3944
rect 4109 3864 4111 3944
rect 4123 3864 4125 3944
rect 4129 3932 4145 3944
rect 4129 3864 4131 3932
rect 4143 3864 4145 3932
rect 4149 3936 4163 3944
rect 4149 3864 4151 3936
rect 4229 3864 4231 3904
rect 4235 3864 4237 3904
rect 4249 3864 4251 3904
rect 4255 3864 4257 3904
rect 4354 3864 4356 3944
rect 4360 3864 4364 3944
rect 4368 3864 4370 3944
rect 4382 3864 4386 3904
rect 4390 3864 4392 3904
rect 4494 3864 4496 3944
rect 4500 3864 4504 3944
rect 4508 3864 4510 3944
rect 4522 3864 4526 3904
rect 4530 3864 4532 3904
rect 4629 3864 4631 3944
rect 4635 3864 4641 3944
rect 4645 3943 4661 3944
rect 4645 3864 4647 3943
rect 4659 3864 4661 3943
rect 4665 3943 4679 3944
rect 4665 3864 4667 3943
rect 4783 3864 4785 3904
rect 4789 3864 4791 3904
rect 4803 3864 4805 3904
rect 4809 3864 4811 3904
rect 4889 3864 4891 3904
rect 4895 3864 4897 3904
rect 4909 3864 4911 3904
rect 4915 3900 4931 3904
rect 4915 3864 4917 3900
rect 4929 3864 4931 3900
rect 4935 3864 4937 3904
rect 5029 3864 5031 3904
rect 5035 3864 5037 3904
rect 5143 3864 5145 3904
rect 5149 3864 5151 3904
rect 5189 3864 5191 3944
rect 5195 3884 5204 3944
rect 5372 3904 5381 3944
rect 5230 3884 5241 3904
rect 5195 3864 5197 3884
rect 5209 3864 5213 3884
rect 5217 3864 5221 3884
rect 5225 3864 5227 3884
rect 5239 3864 5241 3884
rect 5245 3864 5249 3904
rect 5253 3864 5255 3904
rect 5293 3864 5295 3904
rect 5299 3864 5301 3904
rect 5313 3864 5315 3904
rect 5319 3864 5327 3904
rect 5331 3864 5333 3904
rect 5345 3864 5347 3904
rect 5351 3864 5361 3904
rect 5365 3864 5367 3904
rect 5379 3864 5381 3904
rect 5385 3864 5387 3944
rect 5429 3864 5431 3944
rect 5435 3884 5444 3944
rect 5612 3904 5621 3944
rect 5470 3884 5481 3904
rect 5435 3864 5437 3884
rect 5449 3864 5453 3884
rect 5457 3864 5461 3884
rect 5465 3864 5467 3884
rect 5479 3864 5481 3884
rect 5485 3864 5489 3904
rect 5493 3864 5495 3904
rect 5533 3864 5535 3904
rect 5539 3864 5541 3904
rect 5553 3864 5555 3904
rect 5559 3864 5567 3904
rect 5571 3864 5573 3904
rect 5585 3864 5587 3904
rect 5591 3864 5601 3904
rect 5605 3864 5607 3904
rect 5619 3864 5621 3904
rect 5625 3864 5627 3944
rect 5714 3864 5716 3944
rect 5720 3864 5724 3944
rect 5728 3864 5730 3944
rect 5742 3864 5746 3904
rect 5750 3864 5752 3904
rect 83 3796 85 3836
rect 89 3796 91 3836
rect 103 3796 105 3836
rect 109 3796 111 3836
rect 203 3796 205 3836
rect 209 3800 211 3836
rect 223 3800 225 3836
rect 209 3796 225 3800
rect 229 3796 231 3836
rect 243 3796 245 3836
rect 249 3796 251 3836
rect 339 3768 341 3828
rect 345 3824 361 3828
rect 345 3772 347 3824
rect 359 3772 361 3824
rect 345 3768 361 3772
rect 365 3768 367 3828
rect 403 3778 405 3836
rect 391 3776 405 3778
rect 409 3824 425 3836
rect 409 3776 411 3824
rect 423 3776 425 3824
rect 429 3776 431 3836
rect 443 3776 445 3836
rect 449 3776 451 3836
rect 463 3776 465 3836
rect 469 3776 471 3836
rect 568 3796 570 3836
rect 574 3796 578 3836
rect 590 3756 592 3836
rect 596 3756 600 3836
rect 604 3756 606 3836
rect 703 3796 705 3836
rect 709 3796 711 3836
rect 723 3796 725 3836
rect 729 3796 731 3836
rect 814 3756 816 3836
rect 820 3756 824 3836
rect 828 3756 830 3836
rect 842 3796 846 3836
rect 850 3796 852 3836
rect 983 3756 985 3836
rect 989 3824 1005 3836
rect 989 3756 991 3824
rect 1003 3756 1005 3824
rect 1009 3758 1011 3836
rect 1023 3758 1025 3836
rect 1009 3756 1025 3758
rect 1029 3770 1031 3836
rect 1043 3770 1045 3836
rect 1029 3756 1045 3770
rect 1049 3758 1051 3836
rect 1129 3796 1131 3836
rect 1135 3796 1137 3836
rect 1149 3796 1151 3836
rect 1155 3796 1157 3836
rect 1249 3796 1251 3836
rect 1255 3796 1257 3836
rect 1269 3796 1271 3836
rect 1275 3800 1277 3836
rect 1289 3800 1291 3836
rect 1275 3796 1291 3800
rect 1295 3796 1297 3836
rect 1049 3756 1063 3758
rect 1389 3764 1391 3836
rect 1377 3756 1391 3764
rect 1395 3768 1397 3836
rect 1409 3768 1411 3836
rect 1395 3756 1411 3768
rect 1415 3756 1417 3836
rect 1429 3756 1431 3836
rect 1435 3756 1437 3836
rect 1534 3756 1536 3836
rect 1540 3756 1544 3836
rect 1548 3756 1550 3836
rect 1562 3796 1566 3836
rect 1570 3796 1572 3836
rect 1669 3796 1671 3836
rect 1675 3796 1677 3836
rect 1783 3796 1785 3836
rect 1789 3796 1791 3836
rect 1803 3796 1805 3836
rect 1809 3796 1811 3836
rect 1889 3796 1891 3836
rect 1895 3796 1897 3836
rect 1909 3796 1911 3836
rect 1915 3796 1917 3836
rect 2009 3756 2011 3836
rect 2015 3756 2021 3836
rect 2025 3757 2027 3836
rect 2039 3757 2041 3836
rect 2025 3756 2041 3757
rect 2045 3757 2047 3836
rect 2149 3796 2151 3836
rect 2155 3796 2157 3836
rect 2169 3796 2171 3836
rect 2175 3796 2177 3836
rect 2269 3796 2271 3836
rect 2275 3796 2277 3836
rect 2289 3796 2291 3836
rect 2295 3800 2297 3836
rect 2309 3800 2311 3836
rect 2295 3796 2311 3800
rect 2315 3796 2317 3836
rect 2428 3796 2430 3836
rect 2434 3796 2438 3836
rect 2045 3756 2059 3757
rect 2450 3756 2452 3836
rect 2456 3756 2460 3836
rect 2464 3756 2466 3836
rect 2549 3796 2551 3836
rect 2555 3796 2557 3836
rect 2569 3796 2571 3836
rect 2575 3796 2577 3836
rect 2674 3756 2676 3836
rect 2680 3756 2684 3836
rect 2688 3756 2690 3836
rect 2702 3796 2706 3836
rect 2710 3796 2712 3836
rect 2823 3796 2825 3836
rect 2829 3796 2831 3836
rect 2928 3796 2930 3836
rect 2934 3796 2938 3836
rect 2950 3756 2952 3836
rect 2956 3756 2960 3836
rect 2964 3756 2966 3836
rect 3049 3796 3051 3836
rect 3055 3796 3057 3836
rect 3069 3796 3071 3836
rect 3075 3796 3077 3836
rect 3203 3796 3205 3836
rect 3209 3796 3211 3836
rect 3223 3796 3225 3836
rect 3229 3796 3231 3836
rect 3323 3796 3325 3836
rect 3329 3796 3331 3836
rect 3409 3796 3411 3836
rect 3415 3796 3417 3836
rect 3429 3796 3431 3836
rect 3435 3800 3437 3836
rect 3449 3800 3451 3836
rect 3435 3796 3451 3800
rect 3455 3796 3457 3836
rect 3549 3796 3551 3836
rect 3555 3796 3557 3836
rect 3675 3756 3677 3836
rect 3681 3756 3685 3836
rect 3689 3756 3691 3836
rect 3789 3796 3791 3836
rect 3795 3796 3797 3836
rect 3809 3796 3811 3836
rect 3815 3796 3817 3836
rect 3909 3796 3911 3836
rect 3915 3796 3917 3836
rect 4023 3796 4025 3836
rect 4029 3796 4031 3836
rect 4069 3756 4071 3836
rect 4075 3816 4077 3836
rect 4089 3816 4093 3836
rect 4097 3816 4101 3836
rect 4105 3816 4107 3836
rect 4119 3816 4121 3836
rect 4075 3756 4084 3816
rect 4110 3796 4121 3816
rect 4125 3796 4129 3836
rect 4133 3796 4135 3836
rect 4173 3796 4175 3836
rect 4179 3796 4181 3836
rect 4193 3796 4195 3836
rect 4199 3796 4207 3836
rect 4211 3796 4213 3836
rect 4225 3796 4227 3836
rect 4231 3796 4241 3836
rect 4245 3796 4247 3836
rect 4259 3796 4261 3836
rect 4252 3756 4261 3796
rect 4265 3756 4267 3836
rect 4373 3756 4375 3836
rect 4379 3756 4385 3836
rect 4389 3756 4391 3836
rect 4413 3756 4415 3836
rect 4419 3756 4425 3836
rect 4429 3756 4431 3836
rect 4509 3796 4511 3836
rect 4515 3796 4517 3836
rect 4529 3796 4531 3836
rect 4535 3796 4537 3836
rect 4629 3756 4631 3836
rect 4635 3756 4639 3836
rect 4643 3756 4645 3836
rect 4754 3756 4756 3836
rect 4760 3756 4764 3836
rect 4768 3756 4770 3836
rect 4782 3796 4786 3836
rect 4790 3796 4792 3836
rect 4889 3756 4891 3836
rect 4895 3756 4897 3836
rect 5023 3796 5025 3836
rect 5029 3796 5031 3836
rect 5043 3796 5045 3836
rect 5049 3796 5051 3836
rect 5129 3796 5131 3836
rect 5135 3796 5137 3836
rect 5243 3756 5245 3836
rect 5249 3756 5251 3836
rect 5263 3756 5265 3836
rect 5269 3756 5271 3836
rect 5283 3756 5285 3836
rect 5289 3756 5291 3836
rect 5303 3756 5305 3836
rect 5309 3756 5311 3836
rect 5323 3756 5325 3836
rect 5329 3756 5331 3836
rect 5343 3756 5345 3836
rect 5349 3756 5351 3836
rect 5363 3756 5365 3836
rect 5369 3756 5371 3836
rect 5383 3756 5385 3836
rect 5389 3756 5391 3836
rect 5429 3756 5431 3836
rect 5435 3816 5437 3836
rect 5449 3816 5453 3836
rect 5457 3816 5461 3836
rect 5465 3816 5467 3836
rect 5479 3816 5481 3836
rect 5435 3756 5444 3816
rect 5470 3796 5481 3816
rect 5485 3796 5489 3836
rect 5493 3796 5495 3836
rect 5533 3796 5535 3836
rect 5539 3796 5541 3836
rect 5553 3796 5555 3836
rect 5559 3796 5567 3836
rect 5571 3796 5573 3836
rect 5585 3796 5587 3836
rect 5591 3796 5601 3836
rect 5605 3796 5607 3836
rect 5619 3796 5621 3836
rect 5612 3756 5621 3796
rect 5625 3756 5627 3836
rect 5723 3796 5725 3836
rect 5729 3796 5731 3836
rect 5743 3796 5745 3836
rect 5749 3796 5751 3836
rect 88 3384 90 3424
rect 94 3384 98 3424
rect 110 3384 112 3464
rect 116 3384 120 3464
rect 124 3384 126 3464
rect 197 3456 211 3464
rect 209 3384 211 3456
rect 215 3452 231 3464
rect 215 3384 217 3452
rect 229 3384 231 3452
rect 235 3384 237 3464
rect 249 3384 251 3464
rect 255 3384 257 3464
rect 349 3384 351 3424
rect 355 3384 357 3424
rect 454 3384 456 3464
rect 460 3384 464 3464
rect 468 3384 470 3464
rect 482 3384 486 3424
rect 490 3384 492 3424
rect 589 3384 591 3424
rect 595 3384 597 3424
rect 609 3384 611 3424
rect 615 3420 631 3424
rect 615 3384 617 3420
rect 629 3384 631 3420
rect 635 3384 637 3424
rect 763 3384 765 3424
rect 769 3384 771 3424
rect 783 3384 785 3424
rect 789 3384 791 3424
rect 883 3384 885 3424
rect 889 3384 891 3424
rect 903 3384 905 3424
rect 909 3384 911 3424
rect 994 3384 996 3464
rect 1000 3384 1004 3464
rect 1008 3384 1010 3464
rect 1022 3384 1026 3424
rect 1030 3384 1032 3424
rect 1143 3384 1145 3424
rect 1149 3420 1165 3424
rect 1149 3384 1151 3420
rect 1163 3384 1165 3420
rect 1169 3384 1171 3424
rect 1183 3384 1185 3424
rect 1189 3384 1191 3424
rect 1269 3384 1271 3424
rect 1275 3384 1277 3424
rect 1289 3384 1291 3424
rect 1295 3384 1297 3424
rect 1403 3384 1405 3424
rect 1409 3420 1425 3424
rect 1409 3384 1411 3420
rect 1423 3384 1425 3420
rect 1429 3384 1431 3424
rect 1443 3384 1445 3424
rect 1449 3384 1451 3424
rect 1534 3384 1536 3464
rect 1540 3384 1544 3464
rect 1548 3384 1550 3464
rect 1562 3384 1566 3424
rect 1570 3384 1572 3424
rect 1683 3384 1685 3464
rect 1689 3384 1691 3464
rect 1703 3384 1705 3464
rect 1709 3452 1725 3464
rect 1709 3384 1711 3452
rect 1723 3384 1725 3452
rect 1729 3456 1743 3464
rect 1729 3384 1731 3456
rect 1937 3456 1951 3464
rect 1823 3384 1825 3424
rect 1829 3420 1845 3424
rect 1829 3384 1831 3420
rect 1843 3384 1845 3420
rect 1849 3384 1851 3424
rect 1863 3384 1865 3424
rect 1869 3384 1871 3424
rect 1949 3384 1951 3456
rect 1955 3452 1971 3464
rect 1955 3384 1957 3452
rect 1969 3384 1971 3452
rect 1975 3384 1977 3464
rect 1989 3384 1991 3464
rect 1995 3384 1997 3464
rect 2108 3384 2110 3424
rect 2114 3384 2118 3424
rect 2130 3384 2132 3464
rect 2136 3384 2140 3464
rect 2144 3384 2146 3464
rect 2254 3384 2256 3464
rect 2260 3384 2264 3464
rect 2268 3384 2270 3464
rect 2282 3384 2286 3424
rect 2290 3384 2292 3424
rect 2403 3384 2405 3464
rect 2409 3384 2411 3464
rect 2423 3384 2425 3464
rect 2429 3452 2445 3464
rect 2429 3384 2431 3452
rect 2443 3384 2445 3452
rect 2449 3456 2463 3464
rect 2449 3384 2451 3456
rect 2539 3384 2541 3464
rect 2545 3384 2547 3464
rect 2559 3384 2563 3424
rect 2567 3384 2571 3424
rect 2583 3384 2585 3424
rect 2589 3384 2591 3424
rect 2669 3384 2671 3424
rect 2675 3384 2677 3424
rect 2689 3384 2691 3424
rect 2695 3384 2697 3424
rect 2808 3384 2810 3424
rect 2814 3384 2818 3424
rect 2830 3384 2832 3464
rect 2836 3384 2840 3464
rect 2844 3384 2846 3464
rect 2961 3384 2963 3464
rect 2967 3384 2969 3464
rect 2981 3384 2985 3424
rect 2989 3384 2991 3424
rect 3083 3384 3085 3424
rect 3089 3384 3091 3424
rect 3103 3384 3105 3424
rect 3109 3384 3111 3424
rect 3189 3384 3191 3424
rect 3195 3384 3197 3424
rect 3209 3384 3211 3424
rect 3215 3420 3231 3424
rect 3215 3384 3217 3420
rect 3229 3384 3231 3420
rect 3235 3384 3237 3424
rect 3343 3384 3345 3424
rect 3349 3420 3365 3424
rect 3349 3384 3351 3420
rect 3363 3384 3365 3420
rect 3369 3384 3371 3424
rect 3383 3384 3385 3424
rect 3389 3384 3391 3424
rect 3488 3384 3490 3424
rect 3494 3384 3498 3424
rect 3510 3384 3512 3464
rect 3516 3384 3520 3464
rect 3524 3384 3526 3464
rect 3628 3384 3630 3424
rect 3634 3384 3638 3424
rect 3650 3384 3652 3464
rect 3656 3384 3660 3464
rect 3664 3384 3666 3464
rect 3759 3384 3761 3464
rect 3765 3384 3767 3464
rect 3779 3384 3783 3424
rect 3787 3384 3791 3424
rect 3803 3384 3805 3424
rect 3809 3384 3811 3424
rect 3889 3384 3891 3464
rect 3895 3384 3899 3464
rect 3903 3384 3905 3464
rect 4048 3384 4050 3424
rect 4054 3384 4058 3424
rect 4070 3384 4072 3464
rect 4076 3384 4080 3464
rect 4084 3384 4086 3464
rect 4169 3384 4171 3424
rect 4175 3384 4177 3424
rect 4274 3384 4276 3464
rect 4280 3384 4284 3464
rect 4288 3384 4290 3464
rect 4302 3384 4306 3424
rect 4310 3384 4312 3424
rect 4423 3384 4425 3424
rect 4429 3384 4431 3424
rect 4443 3384 4445 3424
rect 4449 3384 4451 3424
rect 4529 3384 4531 3424
rect 4535 3384 4537 3424
rect 4549 3384 4551 3424
rect 4555 3384 4557 3424
rect 4609 3384 4611 3464
rect 4615 3404 4624 3464
rect 4792 3424 4801 3464
rect 4650 3404 4661 3424
rect 4615 3384 4617 3404
rect 4629 3384 4633 3404
rect 4637 3384 4641 3404
rect 4645 3384 4647 3404
rect 4659 3384 4661 3404
rect 4665 3384 4669 3424
rect 4673 3384 4675 3424
rect 4713 3384 4715 3424
rect 4719 3384 4721 3424
rect 4733 3384 4735 3424
rect 4739 3384 4747 3424
rect 4751 3384 4753 3424
rect 4765 3384 4767 3424
rect 4771 3384 4781 3424
rect 4785 3384 4787 3424
rect 4799 3384 4801 3424
rect 4805 3384 4807 3464
rect 4903 3384 4905 3424
rect 4909 3384 4911 3424
rect 4923 3384 4925 3424
rect 4929 3384 4931 3424
rect 5028 3384 5030 3424
rect 5034 3384 5038 3424
rect 5050 3384 5052 3464
rect 5056 3384 5060 3464
rect 5064 3384 5066 3464
rect 5169 3384 5171 3424
rect 5175 3384 5177 3424
rect 5189 3384 5191 3424
rect 5195 3384 5197 3424
rect 5253 3384 5255 3464
rect 5259 3424 5268 3464
rect 5259 3384 5261 3424
rect 5273 3384 5275 3424
rect 5279 3384 5289 3424
rect 5293 3384 5295 3424
rect 5307 3384 5309 3424
rect 5313 3384 5321 3424
rect 5325 3384 5327 3424
rect 5339 3384 5341 3424
rect 5345 3384 5347 3424
rect 5385 3384 5387 3424
rect 5391 3384 5395 3424
rect 5399 3404 5410 3424
rect 5436 3404 5445 3464
rect 5399 3384 5401 3404
rect 5413 3384 5415 3404
rect 5419 3384 5423 3404
rect 5427 3384 5431 3404
rect 5443 3384 5445 3404
rect 5449 3384 5451 3464
rect 5543 3384 5545 3424
rect 5549 3384 5551 3424
rect 5563 3384 5565 3424
rect 5569 3384 5571 3424
rect 5654 3384 5656 3464
rect 5660 3384 5664 3464
rect 5668 3384 5670 3464
rect 5682 3384 5686 3424
rect 5690 3384 5692 3424
rect 83 3316 85 3356
rect 89 3316 91 3356
rect 188 3316 190 3356
rect 194 3316 198 3356
rect 210 3276 212 3356
rect 216 3276 220 3356
rect 224 3276 226 3356
rect 323 3316 325 3356
rect 329 3316 331 3356
rect 409 3316 411 3356
rect 415 3316 417 3356
rect 429 3316 431 3356
rect 435 3316 437 3356
rect 529 3284 531 3356
rect 517 3276 531 3284
rect 535 3288 537 3356
rect 549 3288 551 3356
rect 535 3276 551 3288
rect 555 3276 557 3356
rect 569 3276 571 3356
rect 575 3276 577 3356
rect 669 3316 671 3356
rect 675 3316 677 3356
rect 689 3316 693 3356
rect 697 3316 701 3356
rect 713 3276 715 3356
rect 719 3276 721 3356
rect 843 3316 845 3356
rect 849 3316 851 3356
rect 863 3316 865 3356
rect 869 3316 871 3356
rect 963 3316 965 3356
rect 969 3320 971 3356
rect 983 3320 985 3356
rect 969 3316 985 3320
rect 989 3316 991 3356
rect 1003 3316 1005 3356
rect 1009 3316 1011 3356
rect 1103 3316 1105 3356
rect 1109 3320 1111 3356
rect 1123 3320 1125 3356
rect 1109 3316 1125 3320
rect 1129 3316 1131 3356
rect 1143 3316 1145 3356
rect 1149 3316 1151 3356
rect 1229 3284 1231 3356
rect 1217 3276 1231 3284
rect 1235 3288 1237 3356
rect 1249 3288 1251 3356
rect 1235 3276 1251 3288
rect 1255 3276 1257 3356
rect 1269 3276 1271 3356
rect 1275 3276 1277 3356
rect 1383 3316 1385 3356
rect 1389 3316 1391 3356
rect 1483 3316 1485 3356
rect 1489 3320 1491 3356
rect 1503 3320 1505 3356
rect 1489 3316 1505 3320
rect 1509 3316 1511 3356
rect 1523 3316 1525 3356
rect 1529 3316 1531 3356
rect 1623 3316 1625 3356
rect 1629 3320 1631 3356
rect 1643 3320 1645 3356
rect 1629 3316 1645 3320
rect 1649 3316 1651 3356
rect 1663 3316 1665 3356
rect 1669 3316 1671 3356
rect 1763 3276 1765 3356
rect 1769 3276 1771 3356
rect 1783 3276 1785 3356
rect 1789 3288 1791 3356
rect 1803 3288 1805 3356
rect 1789 3276 1805 3288
rect 1809 3284 1811 3356
rect 1923 3316 1925 3356
rect 1929 3316 1931 3356
rect 1943 3316 1945 3356
rect 1949 3316 1951 3356
rect 1809 3276 1823 3284
rect 2043 3276 2045 3356
rect 2049 3276 2051 3356
rect 2063 3276 2065 3356
rect 2069 3288 2071 3356
rect 2083 3288 2085 3356
rect 2069 3276 2085 3288
rect 2089 3284 2091 3356
rect 2169 3316 2171 3356
rect 2175 3316 2177 3356
rect 2189 3316 2191 3356
rect 2195 3316 2197 3356
rect 2089 3276 2103 3284
rect 2299 3276 2301 3356
rect 2305 3276 2307 3356
rect 2319 3316 2323 3356
rect 2327 3316 2331 3356
rect 2343 3316 2345 3356
rect 2349 3316 2351 3356
rect 2429 3316 2431 3356
rect 2435 3316 2437 3356
rect 2449 3316 2451 3356
rect 2455 3316 2457 3356
rect 2568 3316 2570 3356
rect 2574 3316 2578 3356
rect 2590 3276 2592 3356
rect 2596 3276 2600 3356
rect 2604 3276 2606 3356
rect 2703 3276 2705 3356
rect 2709 3276 2711 3356
rect 2723 3276 2725 3356
rect 2729 3288 2731 3356
rect 2743 3288 2745 3356
rect 2729 3276 2745 3288
rect 2749 3284 2751 3356
rect 2829 3316 2831 3356
rect 2835 3316 2837 3356
rect 2849 3316 2851 3356
rect 2855 3320 2857 3356
rect 2869 3320 2871 3356
rect 2855 3316 2871 3320
rect 2875 3316 2877 3356
rect 2969 3316 2971 3356
rect 2975 3316 2977 3356
rect 2989 3316 2991 3356
rect 2995 3320 2997 3356
rect 3009 3320 3011 3356
rect 2995 3316 3011 3320
rect 3015 3316 3017 3356
rect 3123 3316 3125 3356
rect 3129 3316 3131 3356
rect 3143 3316 3145 3356
rect 3149 3316 3151 3356
rect 3263 3316 3265 3356
rect 3269 3316 3271 3356
rect 3283 3316 3285 3356
rect 3289 3316 3291 3356
rect 3369 3316 3371 3356
rect 3375 3316 3377 3356
rect 3483 3316 3485 3356
rect 3489 3320 3491 3356
rect 3503 3320 3505 3356
rect 3489 3316 3505 3320
rect 3509 3316 3511 3356
rect 3523 3316 3525 3356
rect 3529 3316 3531 3356
rect 2749 3276 2763 3284
rect 3609 3284 3611 3356
rect 3597 3276 3611 3284
rect 3615 3288 3617 3356
rect 3629 3288 3631 3356
rect 3615 3276 3631 3288
rect 3635 3276 3637 3356
rect 3649 3276 3651 3356
rect 3655 3276 3657 3356
rect 3768 3316 3770 3356
rect 3774 3316 3778 3356
rect 3790 3276 3792 3356
rect 3796 3276 3800 3356
rect 3804 3276 3806 3356
rect 3889 3316 3891 3356
rect 3895 3316 3897 3356
rect 3949 3276 3951 3356
rect 3955 3336 3957 3356
rect 3969 3336 3973 3356
rect 3977 3336 3981 3356
rect 3985 3336 3987 3356
rect 3999 3336 4001 3356
rect 3955 3276 3964 3336
rect 3990 3316 4001 3336
rect 4005 3316 4009 3356
rect 4013 3316 4015 3356
rect 4053 3316 4055 3356
rect 4059 3316 4061 3356
rect 4073 3316 4075 3356
rect 4079 3316 4087 3356
rect 4091 3316 4093 3356
rect 4105 3316 4107 3356
rect 4111 3316 4121 3356
rect 4125 3316 4127 3356
rect 4139 3316 4141 3356
rect 4132 3276 4141 3316
rect 4145 3276 4147 3356
rect 4234 3276 4236 3356
rect 4240 3276 4244 3356
rect 4248 3276 4250 3356
rect 4262 3316 4266 3356
rect 4270 3316 4272 3356
rect 4374 3276 4376 3356
rect 4380 3276 4384 3356
rect 4388 3276 4390 3356
rect 4402 3316 4406 3356
rect 4410 3316 4412 3356
rect 4469 3276 4471 3356
rect 4475 3336 4477 3356
rect 4489 3336 4493 3356
rect 4497 3336 4501 3356
rect 4505 3336 4507 3356
rect 4519 3336 4521 3356
rect 4475 3276 4484 3336
rect 4510 3316 4521 3336
rect 4525 3316 4529 3356
rect 4533 3316 4535 3356
rect 4573 3316 4575 3356
rect 4579 3316 4581 3356
rect 4593 3316 4595 3356
rect 4599 3316 4607 3356
rect 4611 3316 4613 3356
rect 4625 3316 4627 3356
rect 4631 3316 4641 3356
rect 4645 3316 4647 3356
rect 4659 3316 4661 3356
rect 4652 3276 4661 3316
rect 4665 3276 4667 3356
rect 4754 3276 4756 3356
rect 4760 3276 4764 3356
rect 4768 3276 4770 3356
rect 4782 3316 4786 3356
rect 4790 3316 4792 3356
rect 4903 3316 4905 3356
rect 4909 3316 4911 3356
rect 4923 3316 4925 3356
rect 4929 3316 4931 3356
rect 5028 3316 5030 3356
rect 5034 3316 5038 3356
rect 5050 3276 5052 3356
rect 5056 3276 5060 3356
rect 5064 3276 5066 3356
rect 5163 3316 5165 3356
rect 5169 3316 5171 3356
rect 5263 3316 5265 3356
rect 5269 3316 5271 3356
rect 5283 3316 5285 3356
rect 5289 3316 5291 3356
rect 5369 3316 5371 3356
rect 5375 3316 5377 3356
rect 5494 3276 5496 3356
rect 5500 3276 5504 3356
rect 5508 3276 5510 3356
rect 5522 3316 5526 3356
rect 5530 3316 5532 3356
rect 5663 3316 5665 3356
rect 5669 3316 5671 3356
rect 5683 3316 5685 3356
rect 5689 3316 5691 3356
rect 99 2904 101 2984
rect 105 2904 107 2984
rect 119 2904 123 2944
rect 127 2904 131 2944
rect 143 2904 145 2944
rect 149 2904 151 2944
rect 249 2904 251 2944
rect 255 2904 257 2944
rect 269 2904 271 2944
rect 275 2940 291 2944
rect 275 2904 277 2940
rect 289 2904 291 2940
rect 295 2904 297 2944
rect 389 2904 391 2944
rect 395 2904 397 2944
rect 409 2904 411 2944
rect 415 2904 417 2944
rect 528 2904 530 2944
rect 534 2904 538 2944
rect 550 2904 552 2984
rect 556 2904 560 2984
rect 564 2904 566 2984
rect 654 2904 656 2984
rect 660 2904 664 2984
rect 668 2904 670 2984
rect 682 2904 686 2944
rect 690 2904 692 2944
rect 794 2904 796 2984
rect 800 2904 804 2984
rect 808 2904 810 2984
rect 822 2904 826 2944
rect 830 2904 832 2944
rect 934 2904 936 2984
rect 940 2904 944 2984
rect 948 2904 950 2984
rect 962 2904 966 2944
rect 970 2904 972 2944
rect 1083 2904 1085 2944
rect 1089 2904 1091 2944
rect 1103 2904 1105 2944
rect 1109 2904 1111 2944
rect 1235 2904 1237 2984
rect 1241 2904 1245 2984
rect 1249 2904 1251 2984
rect 1334 2904 1336 2984
rect 1340 2904 1344 2984
rect 1348 2904 1350 2984
rect 1362 2904 1366 2944
rect 1370 2904 1372 2944
rect 1483 2904 1485 2944
rect 1489 2940 1505 2944
rect 1489 2904 1491 2940
rect 1503 2904 1505 2940
rect 1509 2904 1511 2944
rect 1523 2904 1525 2944
rect 1529 2904 1531 2944
rect 1643 2904 1645 2984
rect 1649 2904 1651 2984
rect 1663 2904 1665 2984
rect 1669 2972 1685 2984
rect 1669 2904 1671 2972
rect 1683 2904 1685 2972
rect 1689 2976 1703 2984
rect 1689 2904 1691 2976
rect 1788 2904 1790 2944
rect 1794 2904 1798 2944
rect 1810 2904 1812 2984
rect 1816 2904 1820 2984
rect 1824 2904 1826 2984
rect 1914 2904 1916 2984
rect 1920 2904 1924 2984
rect 1928 2904 1930 2984
rect 1942 2904 1946 2944
rect 1950 2904 1952 2944
rect 2088 2904 2090 2944
rect 2094 2904 2098 2944
rect 2110 2904 2112 2984
rect 2116 2904 2120 2984
rect 2124 2904 2126 2984
rect 2228 2904 2230 2944
rect 2234 2904 2238 2944
rect 2250 2904 2252 2984
rect 2256 2904 2260 2984
rect 2264 2904 2266 2984
rect 2383 2904 2385 2984
rect 2389 2904 2391 2984
rect 2403 2904 2405 2984
rect 2409 2972 2425 2984
rect 2409 2904 2411 2972
rect 2423 2904 2425 2972
rect 2429 2976 2443 2984
rect 2429 2904 2431 2976
rect 2523 2904 2525 2984
rect 2529 2904 2531 2984
rect 2543 2904 2545 2984
rect 2549 2972 2565 2984
rect 2549 2904 2551 2972
rect 2563 2904 2565 2972
rect 2569 2976 2583 2984
rect 2569 2904 2571 2976
rect 2663 2904 2665 2984
rect 2669 2916 2671 2984
rect 2683 2916 2685 2984
rect 2669 2904 2685 2916
rect 2689 2982 2705 2984
rect 2689 2904 2691 2982
rect 2703 2904 2705 2982
rect 2709 2970 2725 2984
rect 2709 2904 2711 2970
rect 2723 2904 2725 2970
rect 2729 2982 2743 2984
rect 2729 2904 2731 2982
rect 2821 2983 2835 2984
rect 2833 2904 2835 2983
rect 2839 2983 2855 2984
rect 2839 2904 2841 2983
rect 2853 2904 2855 2983
rect 2859 2904 2865 2984
rect 2869 2904 2871 2984
rect 2949 2904 2951 2984
rect 2955 2904 2959 2984
rect 2963 2904 2965 2984
rect 3089 2904 3091 2944
rect 3095 2904 3097 2944
rect 3109 2904 3111 2944
rect 3115 2904 3117 2944
rect 3219 2904 3221 2984
rect 3225 2904 3227 2984
rect 3239 2904 3243 2944
rect 3247 2904 3251 2944
rect 3263 2904 3265 2944
rect 3269 2904 3271 2944
rect 3349 2904 3351 2984
rect 3355 2904 3361 2984
rect 3365 2983 3381 2984
rect 3365 2904 3367 2983
rect 3379 2904 3381 2983
rect 3385 2983 3399 2984
rect 3385 2904 3387 2983
rect 3508 2904 3510 2944
rect 3514 2904 3518 2944
rect 3530 2904 3532 2984
rect 3536 2904 3540 2984
rect 3544 2904 3546 2984
rect 3648 2904 3650 2944
rect 3654 2904 3658 2944
rect 3670 2904 3672 2984
rect 3676 2904 3680 2984
rect 3684 2904 3686 2984
rect 3781 2983 3795 2984
rect 3793 2904 3795 2983
rect 3799 2983 3815 2984
rect 3799 2904 3801 2983
rect 3813 2904 3815 2983
rect 3819 2904 3825 2984
rect 3829 2904 3831 2984
rect 3939 2904 3941 2984
rect 3945 2904 3947 2984
rect 3959 2904 3963 2944
rect 3967 2904 3971 2944
rect 3983 2904 3985 2944
rect 3989 2904 3991 2944
rect 4069 2904 4071 2984
rect 4075 2904 4079 2984
rect 4083 2904 4085 2984
rect 4189 2904 4191 2944
rect 4195 2904 4197 2944
rect 4209 2904 4211 2944
rect 4215 2940 4231 2944
rect 4215 2904 4217 2940
rect 4229 2904 4231 2940
rect 4235 2904 4237 2944
rect 4293 2904 4295 2984
rect 4299 2944 4308 2984
rect 4299 2904 4301 2944
rect 4313 2904 4315 2944
rect 4319 2904 4329 2944
rect 4333 2904 4335 2944
rect 4347 2904 4349 2944
rect 4353 2904 4361 2944
rect 4365 2904 4367 2944
rect 4379 2904 4381 2944
rect 4385 2904 4387 2944
rect 4425 2904 4427 2944
rect 4431 2904 4435 2944
rect 4439 2924 4450 2944
rect 4476 2924 4485 2984
rect 4439 2904 4441 2924
rect 4453 2904 4455 2924
rect 4459 2904 4463 2924
rect 4467 2904 4471 2924
rect 4483 2904 4485 2924
rect 4489 2904 4491 2984
rect 4594 2904 4596 2984
rect 4600 2904 4604 2984
rect 4608 2904 4610 2984
rect 4622 2904 4626 2944
rect 4630 2904 4632 2944
rect 4734 2904 4736 2984
rect 4740 2904 4744 2984
rect 4748 2904 4750 2984
rect 4762 2904 4766 2944
rect 4770 2904 4772 2944
rect 4883 2904 4885 2944
rect 4889 2904 4891 2944
rect 4903 2904 4905 2944
rect 4909 2904 4911 2944
rect 4989 2904 4991 2944
rect 4995 2904 4997 2944
rect 5009 2904 5011 2944
rect 5015 2904 5017 2944
rect 5073 2904 5075 2984
rect 5079 2944 5088 2984
rect 5079 2904 5081 2944
rect 5093 2904 5095 2944
rect 5099 2904 5109 2944
rect 5113 2904 5115 2944
rect 5127 2904 5129 2944
rect 5133 2904 5141 2944
rect 5145 2904 5147 2944
rect 5159 2904 5161 2944
rect 5165 2904 5167 2944
rect 5205 2904 5207 2944
rect 5211 2904 5215 2944
rect 5219 2924 5230 2944
rect 5256 2924 5265 2984
rect 5219 2904 5221 2924
rect 5233 2904 5235 2924
rect 5239 2904 5243 2924
rect 5247 2904 5251 2924
rect 5263 2904 5265 2924
rect 5269 2904 5271 2984
rect 5363 2904 5365 2984
rect 5369 2904 5371 2984
rect 5383 2904 5385 2984
rect 5389 2904 5391 2984
rect 5403 2904 5405 2984
rect 5409 2904 5411 2984
rect 5423 2904 5425 2984
rect 5429 2904 5431 2984
rect 5443 2904 5445 2984
rect 5449 2904 5451 2984
rect 5463 2904 5465 2984
rect 5469 2904 5471 2984
rect 5483 2904 5485 2984
rect 5489 2904 5491 2984
rect 5503 2904 5505 2984
rect 5509 2904 5511 2984
rect 5549 2904 5551 2984
rect 5555 2924 5564 2984
rect 5732 2944 5741 2984
rect 5590 2924 5601 2944
rect 5555 2904 5557 2924
rect 5569 2904 5573 2924
rect 5577 2904 5581 2924
rect 5585 2904 5587 2924
rect 5599 2904 5601 2924
rect 5605 2904 5609 2944
rect 5613 2904 5615 2944
rect 5653 2904 5655 2944
rect 5659 2904 5661 2944
rect 5673 2904 5675 2944
rect 5679 2904 5687 2944
rect 5691 2904 5693 2944
rect 5705 2904 5707 2944
rect 5711 2904 5721 2944
rect 5725 2904 5727 2944
rect 5739 2904 5741 2944
rect 5745 2904 5747 2984
rect 83 2836 85 2876
rect 89 2836 91 2876
rect 103 2836 105 2876
rect 109 2836 111 2876
rect 194 2796 196 2876
rect 200 2796 204 2876
rect 208 2796 210 2876
rect 222 2836 226 2876
rect 230 2836 232 2876
rect 343 2836 345 2876
rect 349 2836 351 2876
rect 429 2804 431 2876
rect 417 2796 431 2804
rect 435 2808 437 2876
rect 449 2808 451 2876
rect 435 2796 451 2808
rect 455 2796 457 2876
rect 469 2796 471 2876
rect 475 2796 477 2876
rect 583 2836 585 2876
rect 589 2836 591 2876
rect 603 2836 605 2876
rect 609 2836 611 2876
rect 689 2836 691 2876
rect 695 2836 697 2876
rect 709 2836 713 2876
rect 717 2836 721 2876
rect 733 2796 735 2876
rect 739 2796 741 2876
rect 829 2836 831 2876
rect 835 2836 837 2876
rect 849 2836 851 2876
rect 855 2836 857 2876
rect 949 2804 951 2876
rect 937 2796 951 2804
rect 955 2808 957 2876
rect 969 2808 971 2876
rect 955 2796 971 2808
rect 975 2796 977 2876
rect 989 2796 991 2876
rect 995 2796 997 2876
rect 1089 2836 1091 2876
rect 1095 2836 1097 2876
rect 1109 2836 1111 2876
rect 1115 2836 1117 2876
rect 1248 2836 1250 2876
rect 1254 2836 1258 2876
rect 1270 2796 1272 2876
rect 1276 2796 1280 2876
rect 1284 2796 1286 2876
rect 1374 2796 1376 2876
rect 1380 2796 1384 2876
rect 1388 2796 1390 2876
rect 1402 2836 1406 2876
rect 1410 2836 1412 2876
rect 1533 2797 1535 2876
rect 1521 2796 1535 2797
rect 1539 2797 1541 2876
rect 1553 2797 1555 2876
rect 1539 2796 1555 2797
rect 1559 2796 1565 2876
rect 1569 2796 1571 2876
rect 1649 2796 1651 2876
rect 1655 2796 1659 2876
rect 1663 2796 1665 2876
rect 1779 2796 1781 2876
rect 1785 2796 1787 2876
rect 1799 2836 1803 2876
rect 1807 2836 1811 2876
rect 1823 2836 1825 2876
rect 1829 2836 1831 2876
rect 1943 2836 1945 2876
rect 1949 2836 1951 2876
rect 1963 2836 1965 2876
rect 1969 2836 1971 2876
rect 2054 2796 2056 2876
rect 2060 2796 2064 2876
rect 2068 2796 2070 2876
rect 2082 2836 2086 2876
rect 2090 2836 2092 2876
rect 2199 2796 2201 2876
rect 2205 2796 2207 2876
rect 2219 2836 2223 2876
rect 2227 2836 2231 2876
rect 2243 2836 2245 2876
rect 2249 2836 2251 2876
rect 2343 2836 2345 2876
rect 2349 2836 2351 2876
rect 2363 2836 2365 2876
rect 2369 2836 2371 2876
rect 2469 2796 2471 2876
rect 2475 2796 2479 2876
rect 2483 2796 2485 2876
rect 2603 2836 2605 2876
rect 2609 2840 2611 2876
rect 2623 2840 2625 2876
rect 2609 2836 2625 2840
rect 2629 2836 2631 2876
rect 2643 2836 2645 2876
rect 2649 2836 2651 2876
rect 2739 2796 2741 2876
rect 2745 2796 2747 2876
rect 2759 2836 2763 2876
rect 2767 2836 2771 2876
rect 2783 2836 2785 2876
rect 2789 2836 2791 2876
rect 2894 2796 2896 2876
rect 2900 2796 2904 2876
rect 2908 2796 2910 2876
rect 2922 2836 2926 2876
rect 2930 2836 2932 2876
rect 3043 2836 3045 2876
rect 3049 2840 3051 2876
rect 3063 2840 3065 2876
rect 3049 2836 3065 2840
rect 3069 2836 3071 2876
rect 3083 2836 3085 2876
rect 3089 2836 3091 2876
rect 3169 2836 3171 2876
rect 3175 2836 3177 2876
rect 3189 2836 3191 2876
rect 3195 2836 3197 2876
rect 3308 2836 3310 2876
rect 3314 2836 3318 2876
rect 3330 2796 3332 2876
rect 3336 2796 3340 2876
rect 3344 2796 3346 2876
rect 3439 2796 3441 2876
rect 3445 2796 3447 2876
rect 3459 2836 3463 2876
rect 3467 2836 3471 2876
rect 3483 2836 3485 2876
rect 3489 2836 3491 2876
rect 3569 2796 3571 2876
rect 3575 2796 3579 2876
rect 3583 2796 3585 2876
rect 3689 2836 3691 2876
rect 3695 2836 3697 2876
rect 3709 2836 3711 2876
rect 3715 2840 3717 2876
rect 3729 2840 3731 2876
rect 3715 2836 3731 2840
rect 3735 2836 3737 2876
rect 3829 2836 3831 2876
rect 3835 2836 3837 2876
rect 3849 2836 3851 2876
rect 3855 2836 3857 2876
rect 3963 2796 3965 2876
rect 3969 2796 3971 2876
rect 4068 2836 4070 2876
rect 4074 2836 4078 2876
rect 4090 2796 4092 2876
rect 4096 2796 4100 2876
rect 4104 2796 4106 2876
rect 4189 2836 4191 2876
rect 4195 2836 4197 2876
rect 4209 2836 4211 2876
rect 4215 2836 4217 2876
rect 4309 2796 4311 2876
rect 4315 2796 4317 2876
rect 4409 2836 4411 2876
rect 4415 2836 4417 2876
rect 4469 2796 4471 2876
rect 4475 2856 4477 2876
rect 4489 2856 4493 2876
rect 4497 2856 4501 2876
rect 4505 2856 4507 2876
rect 4519 2856 4521 2876
rect 4475 2796 4484 2856
rect 4510 2836 4521 2856
rect 4525 2836 4529 2876
rect 4533 2836 4535 2876
rect 4573 2836 4575 2876
rect 4579 2836 4581 2876
rect 4593 2836 4595 2876
rect 4599 2836 4607 2876
rect 4611 2836 4613 2876
rect 4625 2836 4627 2876
rect 4631 2836 4641 2876
rect 4645 2836 4647 2876
rect 4659 2836 4661 2876
rect 4652 2796 4661 2836
rect 4665 2796 4667 2876
rect 4713 2796 4715 2876
rect 4719 2836 4721 2876
rect 4733 2836 4735 2876
rect 4739 2836 4749 2876
rect 4753 2836 4755 2876
rect 4767 2836 4769 2876
rect 4773 2836 4781 2876
rect 4785 2836 4787 2876
rect 4799 2836 4801 2876
rect 4805 2836 4807 2876
rect 4845 2836 4847 2876
rect 4851 2836 4855 2876
rect 4859 2856 4861 2876
rect 4873 2856 4875 2876
rect 4879 2856 4883 2876
rect 4887 2856 4891 2876
rect 4903 2856 4905 2876
rect 4859 2836 4870 2856
rect 4719 2796 4728 2836
rect 4896 2796 4905 2856
rect 4909 2796 4911 2876
rect 5014 2796 5016 2876
rect 5020 2796 5024 2876
rect 5028 2796 5030 2876
rect 5042 2836 5046 2876
rect 5050 2836 5052 2876
rect 5149 2836 5151 2876
rect 5155 2836 5157 2876
rect 5169 2836 5171 2876
rect 5175 2836 5177 2876
rect 5257 2874 5271 2876
rect 5269 2796 5271 2874
rect 5275 2796 5277 2876
rect 5289 2796 5291 2876
rect 5295 2796 5297 2876
rect 5349 2796 5351 2876
rect 5355 2856 5357 2876
rect 5369 2856 5373 2876
rect 5377 2856 5381 2876
rect 5385 2856 5387 2876
rect 5399 2856 5401 2876
rect 5355 2796 5364 2856
rect 5390 2836 5401 2856
rect 5405 2836 5409 2876
rect 5413 2836 5415 2876
rect 5453 2836 5455 2876
rect 5459 2836 5461 2876
rect 5473 2836 5475 2876
rect 5479 2836 5487 2876
rect 5491 2836 5493 2876
rect 5505 2836 5507 2876
rect 5511 2836 5521 2876
rect 5525 2836 5527 2876
rect 5539 2836 5541 2876
rect 5532 2796 5541 2836
rect 5545 2796 5547 2876
rect 5634 2796 5636 2876
rect 5640 2796 5644 2876
rect 5648 2796 5650 2876
rect 5662 2836 5666 2876
rect 5670 2836 5672 2876
rect 83 2424 85 2464
rect 89 2424 91 2464
rect 169 2424 171 2464
rect 175 2424 177 2464
rect 283 2424 285 2504
rect 289 2424 291 2504
rect 303 2424 305 2504
rect 309 2492 325 2504
rect 309 2424 311 2492
rect 323 2424 325 2492
rect 329 2496 343 2504
rect 329 2424 331 2496
rect 409 2424 411 2464
rect 415 2424 417 2464
rect 429 2424 431 2464
rect 435 2460 451 2464
rect 435 2424 437 2460
rect 449 2424 451 2460
rect 455 2424 457 2464
rect 549 2424 551 2464
rect 555 2424 557 2464
rect 649 2424 651 2504
rect 655 2424 659 2504
rect 663 2424 665 2504
rect 774 2424 776 2504
rect 780 2424 784 2504
rect 788 2424 790 2504
rect 917 2496 931 2504
rect 802 2424 806 2464
rect 810 2424 812 2464
rect 929 2424 931 2496
rect 935 2492 951 2504
rect 935 2424 937 2492
rect 949 2424 951 2492
rect 955 2424 957 2504
rect 969 2424 971 2504
rect 975 2424 977 2504
rect 1088 2424 1090 2464
rect 1094 2424 1098 2464
rect 1110 2424 1112 2504
rect 1116 2424 1120 2504
rect 1124 2424 1126 2504
rect 1223 2424 1225 2464
rect 1229 2424 1231 2464
rect 1243 2424 1245 2464
rect 1249 2424 1251 2464
rect 1329 2424 1331 2464
rect 1335 2424 1337 2464
rect 1349 2424 1353 2464
rect 1357 2424 1361 2464
rect 1373 2424 1375 2504
rect 1379 2424 1381 2504
rect 1483 2424 1485 2464
rect 1489 2460 1505 2464
rect 1489 2424 1491 2460
rect 1503 2424 1505 2460
rect 1509 2424 1511 2464
rect 1523 2424 1525 2464
rect 1529 2424 1531 2464
rect 1609 2424 1611 2464
rect 1615 2424 1617 2464
rect 1714 2424 1716 2504
rect 1720 2424 1724 2504
rect 1728 2424 1730 2504
rect 1742 2424 1746 2464
rect 1750 2424 1752 2464
rect 1868 2424 1870 2464
rect 1874 2424 1878 2464
rect 1890 2424 1892 2504
rect 1896 2424 1900 2504
rect 1904 2424 1906 2504
rect 1994 2424 1996 2504
rect 2000 2424 2004 2504
rect 2008 2424 2010 2504
rect 2022 2424 2026 2464
rect 2030 2424 2032 2464
rect 2143 2424 2145 2464
rect 2149 2460 2165 2464
rect 2149 2424 2151 2460
rect 2163 2424 2165 2460
rect 2169 2424 2171 2464
rect 2183 2424 2185 2464
rect 2189 2424 2191 2464
rect 2283 2424 2285 2504
rect 2289 2424 2291 2504
rect 2303 2424 2305 2504
rect 2309 2492 2325 2504
rect 2309 2424 2311 2492
rect 2323 2424 2325 2492
rect 2329 2496 2343 2504
rect 2329 2424 2331 2496
rect 2409 2424 2411 2464
rect 2415 2424 2417 2464
rect 2429 2424 2431 2464
rect 2435 2424 2437 2464
rect 2568 2424 2570 2464
rect 2574 2424 2578 2464
rect 2590 2424 2592 2504
rect 2596 2424 2600 2504
rect 2604 2424 2606 2504
rect 2694 2424 2696 2504
rect 2700 2424 2704 2504
rect 2708 2424 2710 2504
rect 2722 2424 2726 2464
rect 2730 2424 2732 2464
rect 2843 2424 2845 2504
rect 2849 2424 2851 2504
rect 2863 2424 2865 2504
rect 2869 2492 2885 2504
rect 2869 2424 2871 2492
rect 2883 2424 2885 2492
rect 2889 2496 2903 2504
rect 2889 2424 2891 2496
rect 2983 2424 2985 2464
rect 2989 2424 2991 2464
rect 3074 2424 3076 2504
rect 3080 2424 3084 2504
rect 3088 2424 3090 2504
rect 3102 2424 3106 2464
rect 3110 2424 3112 2464
rect 3229 2424 3231 2464
rect 3235 2424 3237 2464
rect 3249 2424 3251 2464
rect 3255 2424 3257 2464
rect 3363 2424 3365 2464
rect 3369 2460 3385 2464
rect 3369 2424 3371 2460
rect 3383 2424 3385 2460
rect 3389 2424 3391 2464
rect 3403 2424 3405 2464
rect 3409 2424 3411 2464
rect 3489 2424 3491 2464
rect 3495 2424 3497 2464
rect 3509 2424 3513 2464
rect 3517 2424 3521 2464
rect 3533 2424 3535 2504
rect 3539 2424 3541 2504
rect 3737 2502 3751 2504
rect 3629 2424 3631 2464
rect 3635 2424 3637 2464
rect 3649 2424 3651 2464
rect 3655 2424 3657 2464
rect 3749 2424 3751 2502
rect 3755 2490 3771 2504
rect 3755 2424 3757 2490
rect 3769 2424 3771 2490
rect 3775 2502 3791 2504
rect 3775 2424 3777 2502
rect 3789 2424 3791 2502
rect 3795 2436 3797 2504
rect 3809 2436 3811 2504
rect 3795 2424 3811 2436
rect 3815 2424 3817 2504
rect 3909 2424 3911 2504
rect 3915 2424 3919 2504
rect 3923 2424 3925 2504
rect 3997 2424 3999 2464
rect 4003 2424 4005 2464
rect 4042 2424 4044 2464
rect 4048 2424 4050 2464
rect 4062 2424 4064 2464
rect 4068 2424 4070 2464
rect 4082 2424 4084 2464
rect 4088 2424 4090 2464
rect 4102 2424 4104 2464
rect 4108 2424 4110 2464
rect 4147 2424 4149 2444
rect 4153 2424 4155 2444
rect 4167 2424 4169 2444
rect 4173 2424 4175 2444
rect 4212 2424 4214 2464
rect 4218 2424 4220 2464
rect 4232 2424 4234 2464
rect 4238 2424 4240 2464
rect 4277 2424 4279 2464
rect 4283 2444 4295 2464
rect 4350 2447 4364 2464
rect 4283 2424 4285 2444
rect 4297 2424 4299 2444
rect 4303 2424 4305 2444
rect 4317 2424 4319 2444
rect 4323 2424 4325 2444
rect 4362 2424 4364 2447
rect 4368 2424 4370 2464
rect 4382 2424 4384 2464
rect 4388 2424 4390 2464
rect 4402 2424 4404 2464
rect 4408 2424 4410 2464
rect 4422 2424 4424 2464
rect 4428 2424 4430 2464
rect 4470 2424 4472 2464
rect 4476 2424 4478 2464
rect 4490 2424 4492 2464
rect 4496 2424 4498 2464
rect 4510 2424 4512 2464
rect 4516 2424 4518 2464
rect 4530 2424 4532 2464
rect 4536 2447 4550 2464
rect 4536 2424 4538 2447
rect 4605 2444 4617 2464
rect 4575 2424 4577 2444
rect 4581 2424 4583 2444
rect 4595 2424 4597 2444
rect 4601 2424 4603 2444
rect 4615 2424 4617 2444
rect 4621 2424 4623 2464
rect 4660 2424 4662 2464
rect 4666 2424 4668 2464
rect 4680 2424 4682 2464
rect 4686 2424 4688 2464
rect 4725 2424 4727 2444
rect 4731 2424 4733 2444
rect 4745 2424 4747 2444
rect 4751 2424 4753 2444
rect 4790 2424 4792 2464
rect 4796 2424 4798 2464
rect 4810 2424 4812 2464
rect 4816 2424 4818 2464
rect 4830 2424 4832 2464
rect 4836 2424 4838 2464
rect 4850 2424 4852 2464
rect 4856 2424 4858 2464
rect 4895 2424 4897 2464
rect 4901 2424 4903 2464
rect 4953 2424 4955 2504
rect 4959 2464 4968 2504
rect 4959 2424 4961 2464
rect 4973 2424 4975 2464
rect 4979 2424 4989 2464
rect 4993 2424 4995 2464
rect 5007 2424 5009 2464
rect 5013 2424 5021 2464
rect 5025 2424 5027 2464
rect 5039 2424 5041 2464
rect 5045 2424 5047 2464
rect 5085 2424 5087 2464
rect 5091 2424 5095 2464
rect 5099 2444 5110 2464
rect 5136 2444 5145 2504
rect 5099 2424 5101 2444
rect 5113 2424 5115 2444
rect 5119 2424 5123 2444
rect 5127 2424 5131 2444
rect 5143 2424 5145 2444
rect 5149 2424 5151 2504
rect 5243 2424 5245 2504
rect 5249 2424 5251 2504
rect 5263 2424 5265 2504
rect 5269 2424 5271 2504
rect 5283 2424 5285 2504
rect 5289 2424 5291 2504
rect 5303 2424 5305 2504
rect 5309 2424 5311 2504
rect 5323 2424 5325 2504
rect 5329 2424 5331 2504
rect 5343 2424 5345 2504
rect 5349 2424 5351 2504
rect 5363 2424 5365 2504
rect 5369 2424 5371 2504
rect 5383 2424 5385 2504
rect 5389 2424 5391 2504
rect 5489 2424 5491 2504
rect 5495 2424 5497 2504
rect 5509 2424 5511 2504
rect 5515 2424 5517 2504
rect 5529 2424 5531 2504
rect 5535 2424 5537 2504
rect 5549 2424 5551 2504
rect 5555 2424 5557 2504
rect 5569 2424 5571 2504
rect 5575 2424 5577 2504
rect 5589 2424 5591 2504
rect 5595 2424 5597 2504
rect 5609 2424 5611 2504
rect 5615 2424 5617 2504
rect 5629 2424 5631 2504
rect 5635 2424 5637 2504
rect 5729 2424 5731 2504
rect 5735 2424 5737 2504
rect 81 2316 83 2396
rect 87 2316 89 2396
rect 101 2356 105 2396
rect 109 2356 111 2396
rect 203 2356 205 2396
rect 209 2360 211 2396
rect 223 2360 225 2396
rect 209 2356 225 2360
rect 229 2356 231 2396
rect 243 2356 245 2396
rect 249 2356 251 2396
rect 329 2356 331 2396
rect 335 2356 337 2396
rect 349 2356 351 2396
rect 355 2356 357 2396
rect 454 2316 456 2396
rect 460 2316 464 2396
rect 468 2316 470 2396
rect 482 2356 486 2396
rect 490 2356 492 2396
rect 608 2356 610 2396
rect 614 2356 618 2396
rect 630 2316 632 2396
rect 636 2316 640 2396
rect 644 2316 646 2396
rect 763 2356 765 2396
rect 769 2360 771 2396
rect 783 2360 785 2396
rect 769 2356 785 2360
rect 789 2356 791 2396
rect 803 2356 805 2396
rect 809 2356 811 2396
rect 903 2356 905 2396
rect 909 2356 911 2396
rect 923 2356 925 2396
rect 929 2356 931 2396
rect 1033 2317 1035 2396
rect 1021 2316 1035 2317
rect 1039 2317 1041 2396
rect 1053 2317 1055 2396
rect 1039 2316 1055 2317
rect 1059 2316 1065 2396
rect 1069 2316 1071 2396
rect 1149 2316 1151 2396
rect 1155 2316 1157 2396
rect 1263 2356 1265 2396
rect 1269 2360 1271 2396
rect 1283 2360 1285 2396
rect 1269 2356 1285 2360
rect 1289 2356 1291 2396
rect 1303 2356 1305 2396
rect 1309 2356 1311 2396
rect 1403 2316 1405 2396
rect 1409 2316 1411 2396
rect 1423 2316 1425 2396
rect 1429 2328 1431 2396
rect 1443 2328 1445 2396
rect 1429 2316 1445 2328
rect 1449 2324 1451 2396
rect 1568 2356 1570 2396
rect 1574 2356 1578 2396
rect 1449 2316 1463 2324
rect 1590 2316 1592 2396
rect 1596 2316 1600 2396
rect 1604 2316 1606 2396
rect 1703 2316 1705 2396
rect 1709 2316 1711 2396
rect 1723 2316 1725 2396
rect 1729 2328 1731 2396
rect 1743 2328 1745 2396
rect 1729 2316 1745 2328
rect 1749 2324 1751 2396
rect 1843 2356 1845 2396
rect 1849 2360 1851 2396
rect 1863 2360 1865 2396
rect 1849 2356 1865 2360
rect 1869 2356 1871 2396
rect 1883 2356 1885 2396
rect 1889 2356 1891 2396
rect 1983 2356 1985 2396
rect 1989 2360 1991 2396
rect 2003 2360 2005 2396
rect 1989 2356 2005 2360
rect 2009 2356 2011 2396
rect 2023 2356 2025 2396
rect 2029 2356 2031 2396
rect 2077 2356 2079 2396
rect 2083 2356 2085 2396
rect 2122 2356 2124 2396
rect 2128 2356 2130 2396
rect 2142 2356 2144 2396
rect 2148 2356 2150 2396
rect 2162 2356 2164 2396
rect 2168 2356 2170 2396
rect 2182 2356 2184 2396
rect 2188 2356 2190 2396
rect 2227 2376 2229 2396
rect 2233 2376 2235 2396
rect 2247 2376 2249 2396
rect 2253 2376 2255 2396
rect 1749 2316 1763 2324
rect 2292 2356 2294 2396
rect 2298 2356 2300 2396
rect 2312 2356 2314 2396
rect 2318 2356 2320 2396
rect 2357 2356 2359 2396
rect 2363 2376 2365 2396
rect 2377 2376 2379 2396
rect 2383 2376 2385 2396
rect 2397 2376 2399 2396
rect 2403 2376 2405 2396
rect 2363 2356 2375 2376
rect 2442 2373 2444 2396
rect 2430 2356 2444 2373
rect 2448 2356 2450 2396
rect 2462 2356 2464 2396
rect 2468 2356 2470 2396
rect 2482 2356 2484 2396
rect 2488 2356 2490 2396
rect 2502 2356 2504 2396
rect 2508 2356 2510 2396
rect 2601 2316 2603 2396
rect 2607 2316 2609 2396
rect 2621 2356 2625 2396
rect 2629 2356 2631 2396
rect 2734 2316 2736 2396
rect 2740 2316 2744 2396
rect 2748 2316 2750 2396
rect 2762 2356 2766 2396
rect 2770 2356 2772 2396
rect 2874 2316 2876 2396
rect 2880 2316 2884 2396
rect 2888 2316 2890 2396
rect 2902 2356 2906 2396
rect 2910 2356 2912 2396
rect 3023 2356 3025 2396
rect 3029 2356 3031 2396
rect 3043 2356 3045 2396
rect 3049 2356 3051 2396
rect 3149 2356 3151 2396
rect 3155 2356 3157 2396
rect 3169 2356 3171 2396
rect 3175 2356 3177 2396
rect 3283 2316 3285 2396
rect 3289 2316 3291 2396
rect 3303 2316 3305 2396
rect 3309 2328 3311 2396
rect 3323 2328 3325 2396
rect 3309 2316 3325 2328
rect 3329 2324 3331 2396
rect 3329 2316 3343 2324
rect 3409 2316 3411 2396
rect 3415 2316 3419 2396
rect 3423 2316 3425 2396
rect 3554 2316 3556 2396
rect 3560 2316 3564 2396
rect 3568 2316 3570 2396
rect 3582 2356 3586 2396
rect 3590 2356 3592 2396
rect 3689 2356 3691 2396
rect 3695 2356 3697 2396
rect 3709 2356 3711 2396
rect 3715 2356 3717 2396
rect 3809 2356 3811 2396
rect 3815 2356 3819 2396
rect 3831 2316 3833 2396
rect 3837 2316 3839 2396
rect 3897 2356 3899 2396
rect 3903 2356 3905 2396
rect 3942 2356 3944 2396
rect 3948 2356 3950 2396
rect 3962 2356 3964 2396
rect 3968 2356 3970 2396
rect 3982 2356 3984 2396
rect 3988 2356 3990 2396
rect 4002 2356 4004 2396
rect 4008 2356 4010 2396
rect 4047 2376 4049 2396
rect 4053 2376 4055 2396
rect 4067 2376 4069 2396
rect 4073 2376 4075 2396
rect 4112 2356 4114 2396
rect 4118 2356 4120 2396
rect 4132 2356 4134 2396
rect 4138 2356 4140 2396
rect 4177 2356 4179 2396
rect 4183 2376 4185 2396
rect 4197 2376 4199 2396
rect 4203 2376 4205 2396
rect 4217 2376 4219 2396
rect 4223 2376 4225 2396
rect 4183 2356 4195 2376
rect 4262 2373 4264 2396
rect 4250 2356 4264 2373
rect 4268 2356 4270 2396
rect 4282 2356 4284 2396
rect 4288 2356 4290 2396
rect 4302 2356 4304 2396
rect 4308 2356 4310 2396
rect 4322 2356 4324 2396
rect 4328 2356 4330 2396
rect 4409 2356 4411 2396
rect 4415 2356 4417 2396
rect 4429 2356 4433 2396
rect 4437 2356 4441 2396
rect 4453 2316 4455 2396
rect 4459 2316 4461 2396
rect 4549 2318 4551 2396
rect 4537 2316 4551 2318
rect 4555 2330 4557 2396
rect 4569 2330 4571 2396
rect 4555 2316 4571 2330
rect 4575 2318 4577 2396
rect 4589 2318 4591 2396
rect 4575 2316 4591 2318
rect 4595 2384 4611 2396
rect 4595 2316 4597 2384
rect 4609 2316 4611 2384
rect 4615 2316 4617 2396
rect 4709 2356 4711 2396
rect 4715 2356 4717 2396
rect 4729 2356 4731 2396
rect 4735 2356 4737 2396
rect 4841 2316 4843 2396
rect 4847 2316 4849 2396
rect 4861 2356 4865 2396
rect 4869 2356 4871 2396
rect 4949 2356 4951 2396
rect 4955 2356 4957 2396
rect 5049 2318 5051 2396
rect 5037 2316 5051 2318
rect 5055 2330 5057 2396
rect 5069 2330 5071 2396
rect 5055 2316 5071 2330
rect 5075 2318 5077 2396
rect 5089 2318 5091 2396
rect 5075 2316 5091 2318
rect 5095 2384 5111 2396
rect 5095 2316 5097 2384
rect 5109 2316 5111 2384
rect 5115 2316 5117 2396
rect 5209 2356 5211 2396
rect 5215 2356 5217 2396
rect 5229 2356 5231 2396
rect 5235 2356 5237 2396
rect 5329 2316 5331 2396
rect 5335 2316 5337 2396
rect 5429 2356 5431 2396
rect 5435 2356 5437 2396
rect 5449 2356 5451 2396
rect 5455 2356 5457 2396
rect 5549 2356 5551 2396
rect 5555 2356 5557 2396
rect 5692 2388 5701 2396
rect 5649 2348 5651 2388
rect 5655 2348 5657 2388
rect 5669 2348 5671 2388
rect 5661 2308 5671 2348
rect 5675 2308 5681 2388
rect 5685 2324 5687 2388
rect 5699 2324 5701 2388
rect 5685 2316 5701 2324
rect 5705 2316 5711 2396
rect 5715 2316 5717 2396
rect 5685 2308 5693 2316
rect 101 1944 103 2024
rect 107 1944 109 2024
rect 357 2016 371 2024
rect 121 1944 125 1984
rect 129 1944 131 1984
rect 243 1944 245 1984
rect 249 1980 265 1984
rect 249 1944 251 1980
rect 263 1944 265 1980
rect 269 1944 271 1984
rect 283 1944 285 1984
rect 289 1944 291 1984
rect 369 1944 371 2016
rect 375 2012 391 2024
rect 375 1944 377 2012
rect 389 1944 391 2012
rect 395 1944 397 2024
rect 409 1944 411 2024
rect 415 1944 417 2024
rect 523 1944 525 1984
rect 529 1944 531 1984
rect 628 1944 630 1984
rect 634 1944 638 1984
rect 650 1944 652 2024
rect 656 1944 660 2024
rect 664 1944 666 2024
rect 763 1944 765 2024
rect 769 1944 771 2024
rect 783 1944 785 2024
rect 789 2012 805 2024
rect 789 1944 791 2012
rect 803 1944 805 2012
rect 809 2016 823 2024
rect 809 1944 811 2016
rect 889 1944 891 1984
rect 895 1944 897 1984
rect 909 1944 911 1984
rect 915 1980 931 1984
rect 915 1944 917 1980
rect 929 1944 931 1980
rect 935 1944 937 1984
rect 1063 1944 1065 1984
rect 1069 1980 1085 1984
rect 1069 1944 1071 1980
rect 1083 1944 1085 1980
rect 1089 1944 1091 1984
rect 1103 1944 1105 1984
rect 1109 1944 1111 1984
rect 1208 1944 1210 1984
rect 1214 1944 1218 1984
rect 1230 1944 1232 2024
rect 1236 1944 1240 2024
rect 1244 1944 1246 2024
rect 1348 1944 1350 1984
rect 1354 1944 1358 1984
rect 1370 1944 1372 2024
rect 1376 1944 1380 2024
rect 1384 1944 1386 2024
rect 1483 1944 1485 2024
rect 1489 1944 1491 2024
rect 1503 1944 1505 2024
rect 1509 2012 1525 2024
rect 1509 1944 1511 2012
rect 1523 1944 1525 2012
rect 1529 2016 1543 2024
rect 1529 1944 1531 2016
rect 1623 1944 1625 1984
rect 1629 1980 1645 1984
rect 1629 1944 1631 1980
rect 1643 1944 1645 1980
rect 1649 1944 1651 1984
rect 1663 1944 1665 1984
rect 1669 1944 1671 1984
rect 1754 1944 1756 2024
rect 1760 1944 1764 2024
rect 1768 1944 1770 2024
rect 1877 2016 1891 2024
rect 1782 1944 1786 1984
rect 1790 1944 1792 1984
rect 1889 1944 1891 2016
rect 1895 2012 1911 2024
rect 1895 1944 1897 2012
rect 1909 1944 1911 2012
rect 1915 1944 1917 2024
rect 1929 1944 1931 2024
rect 1935 1944 1937 2024
rect 2039 1952 2041 2012
rect 2045 2008 2061 2012
rect 2045 1956 2047 2008
rect 2059 1956 2061 2008
rect 2045 1952 2061 1956
rect 2065 1952 2067 2012
rect 2091 2002 2105 2004
rect 2103 1944 2105 2002
rect 2109 1956 2111 2004
rect 2123 1956 2125 2004
rect 2109 1944 2125 1956
rect 2129 1944 2131 2004
rect 2143 1944 2145 2004
rect 2149 1944 2151 2004
rect 2163 1944 2165 2004
rect 2169 1944 2171 2004
rect 2263 1944 2265 1984
rect 2269 1980 2285 1984
rect 2269 1944 2271 1980
rect 2283 1944 2285 1980
rect 2289 1944 2291 1984
rect 2303 1944 2305 1984
rect 2309 1944 2311 1984
rect 2357 1944 2359 1984
rect 2363 1944 2365 1984
rect 2402 1944 2404 1984
rect 2408 1944 2410 1984
rect 2422 1944 2424 1984
rect 2428 1944 2430 1984
rect 2442 1944 2444 1984
rect 2448 1944 2450 1984
rect 2462 1944 2464 1984
rect 2468 1944 2470 1984
rect 2507 1944 2509 1964
rect 2513 1944 2515 1964
rect 2527 1944 2529 1964
rect 2533 1944 2535 1964
rect 2572 1944 2574 1984
rect 2578 1944 2580 1984
rect 2592 1944 2594 1984
rect 2598 1944 2600 1984
rect 2637 1944 2639 1984
rect 2643 1964 2655 1984
rect 2710 1967 2724 1984
rect 2643 1944 2645 1964
rect 2657 1944 2659 1964
rect 2663 1944 2665 1964
rect 2677 1944 2679 1964
rect 2683 1944 2685 1964
rect 2722 1944 2724 1967
rect 2728 1944 2730 1984
rect 2742 1944 2744 1984
rect 2748 1944 2750 1984
rect 2762 1944 2764 1984
rect 2768 1944 2770 1984
rect 2782 1944 2784 1984
rect 2788 1944 2790 1984
rect 2874 1944 2876 2024
rect 2880 1944 2884 2024
rect 2888 1944 2890 2024
rect 2902 1944 2906 1984
rect 2910 1944 2912 1984
rect 3023 1944 3025 1984
rect 3029 1944 3031 1984
rect 3043 1944 3045 1984
rect 3049 1944 3051 1984
rect 3129 1944 3131 1984
rect 3135 1944 3137 1984
rect 3149 1944 3151 1984
rect 3155 1944 3157 1984
rect 3269 1944 3271 2024
rect 3275 1944 3279 2024
rect 3283 1944 3285 2024
rect 3399 1944 3401 2024
rect 3405 1944 3407 2024
rect 3517 2016 3531 2024
rect 3419 1944 3423 1984
rect 3427 1944 3431 1984
rect 3443 1944 3445 1984
rect 3449 1944 3451 1984
rect 3529 1944 3531 2016
rect 3535 2012 3551 2024
rect 3535 1944 3537 2012
rect 3549 1944 3551 2012
rect 3555 1944 3557 2024
rect 3569 1944 3571 2024
rect 3575 1944 3577 2024
rect 3703 1944 3705 2024
rect 3709 1944 3711 2024
rect 3809 1944 3811 1984
rect 3815 1944 3817 1984
rect 3829 1944 3831 1984
rect 3835 1980 3851 1984
rect 3835 1944 3837 1980
rect 3849 1944 3851 1980
rect 3855 1944 3857 1984
rect 3969 1944 3971 2024
rect 3975 1944 3977 2024
rect 4099 1944 4101 2024
rect 4105 1944 4107 2024
rect 4119 1944 4123 1984
rect 4127 1944 4131 1984
rect 4143 1944 4145 1984
rect 4149 1944 4151 1984
rect 4243 1944 4245 1984
rect 4249 1944 4251 1984
rect 4263 1944 4265 1984
rect 4269 1944 4271 1984
rect 4368 1944 4370 1984
rect 4374 1944 4378 1984
rect 4390 1944 4392 2024
rect 4396 1944 4400 2024
rect 4404 1944 4406 2024
rect 4494 1944 4496 2024
rect 4500 1944 4504 2024
rect 4508 1944 4510 2024
rect 4522 1944 4526 1984
rect 4530 1944 4532 1984
rect 4629 1944 4631 1984
rect 4635 1944 4637 1984
rect 4649 1944 4651 1984
rect 4655 1944 4657 1984
rect 4749 1944 4751 1984
rect 4755 1944 4757 1984
rect 4769 1944 4771 1984
rect 4775 1944 4777 1984
rect 4908 1944 4910 1984
rect 4914 1944 4918 1984
rect 4930 1944 4932 2024
rect 4936 1944 4940 2024
rect 4944 1944 4946 2024
rect 5048 1944 5050 1984
rect 5054 1944 5058 1984
rect 5070 1944 5072 2024
rect 5076 1944 5080 2024
rect 5084 1944 5086 2024
rect 5169 1944 5171 1984
rect 5175 1944 5177 1984
rect 5269 1944 5271 2024
rect 5275 1944 5279 2024
rect 5283 1944 5285 2024
rect 5389 1944 5391 1984
rect 5395 1944 5397 1984
rect 5409 1944 5411 1984
rect 5415 1944 5417 1984
rect 5509 1944 5511 1984
rect 5515 1944 5517 1984
rect 5623 1944 5625 1984
rect 5629 1944 5631 1984
rect 5714 1944 5716 2024
rect 5720 1944 5724 2024
rect 5728 1944 5730 2024
rect 5742 1944 5746 1984
rect 5750 1944 5752 1984
rect 83 1876 85 1916
rect 89 1880 91 1916
rect 103 1880 105 1916
rect 89 1876 105 1880
rect 109 1876 111 1916
rect 123 1876 125 1916
rect 129 1876 131 1916
rect 209 1844 211 1916
rect 197 1836 211 1844
rect 215 1848 217 1916
rect 229 1848 231 1916
rect 215 1836 231 1848
rect 235 1836 237 1916
rect 249 1836 251 1916
rect 255 1836 257 1916
rect 368 1876 370 1916
rect 374 1876 378 1916
rect 390 1836 392 1916
rect 396 1836 400 1916
rect 404 1836 406 1916
rect 503 1876 505 1916
rect 509 1880 511 1916
rect 523 1880 525 1916
rect 509 1876 525 1880
rect 529 1876 531 1916
rect 543 1876 545 1916
rect 549 1876 551 1916
rect 675 1836 677 1916
rect 681 1836 685 1916
rect 689 1836 691 1916
rect 769 1844 771 1916
rect 757 1836 771 1844
rect 775 1848 777 1916
rect 789 1848 791 1916
rect 775 1836 791 1848
rect 795 1836 797 1916
rect 809 1836 811 1916
rect 815 1836 817 1916
rect 943 1876 945 1916
rect 949 1876 951 1916
rect 1068 1876 1070 1916
rect 1074 1876 1078 1916
rect 1090 1836 1092 1916
rect 1096 1836 1100 1916
rect 1104 1836 1106 1916
rect 1208 1876 1210 1916
rect 1214 1876 1218 1916
rect 1230 1836 1232 1916
rect 1236 1836 1240 1916
rect 1244 1836 1246 1916
rect 1343 1876 1345 1916
rect 1349 1876 1351 1916
rect 1448 1876 1450 1916
rect 1454 1876 1458 1916
rect 1470 1836 1472 1916
rect 1476 1836 1480 1916
rect 1484 1836 1486 1916
rect 1574 1836 1576 1916
rect 1580 1836 1584 1916
rect 1588 1836 1590 1916
rect 1602 1876 1606 1916
rect 1610 1876 1612 1916
rect 1728 1876 1730 1916
rect 1734 1876 1738 1916
rect 1750 1836 1752 1916
rect 1756 1836 1760 1916
rect 1764 1836 1766 1916
rect 1863 1876 1865 1916
rect 1869 1876 1871 1916
rect 1883 1876 1885 1916
rect 1889 1876 1891 1916
rect 1983 1876 1985 1916
rect 1989 1876 1991 1916
rect 2003 1876 2005 1916
rect 2009 1876 2011 1916
rect 2123 1836 2125 1916
rect 2129 1836 2131 1916
rect 2143 1836 2145 1916
rect 2149 1914 2163 1916
rect 2149 1836 2151 1914
rect 2197 1876 2199 1916
rect 2203 1876 2205 1916
rect 2242 1876 2244 1916
rect 2248 1876 2250 1916
rect 2262 1876 2264 1916
rect 2268 1876 2270 1916
rect 2282 1876 2284 1916
rect 2288 1876 2290 1916
rect 2302 1876 2304 1916
rect 2308 1876 2310 1916
rect 2347 1896 2349 1916
rect 2353 1896 2355 1916
rect 2367 1896 2369 1916
rect 2373 1896 2375 1916
rect 2412 1876 2414 1916
rect 2418 1876 2420 1916
rect 2432 1876 2434 1916
rect 2438 1876 2440 1916
rect 2477 1876 2479 1916
rect 2483 1896 2485 1916
rect 2497 1896 2499 1916
rect 2503 1896 2505 1916
rect 2517 1896 2519 1916
rect 2523 1896 2525 1916
rect 2483 1876 2495 1896
rect 2562 1893 2564 1916
rect 2550 1876 2564 1893
rect 2568 1876 2570 1916
rect 2582 1876 2584 1916
rect 2588 1876 2590 1916
rect 2602 1876 2604 1916
rect 2608 1876 2610 1916
rect 2622 1876 2624 1916
rect 2628 1876 2630 1916
rect 2709 1876 2711 1916
rect 2715 1876 2717 1916
rect 2729 1876 2731 1916
rect 2735 1876 2737 1916
rect 2843 1876 2845 1916
rect 2849 1880 2851 1916
rect 2863 1880 2865 1916
rect 2849 1876 2865 1880
rect 2869 1876 2871 1916
rect 2883 1876 2885 1916
rect 2889 1876 2891 1916
rect 2988 1876 2990 1916
rect 2994 1876 2998 1916
rect 3010 1836 3012 1916
rect 3016 1836 3020 1916
rect 3024 1836 3026 1916
rect 3109 1836 3111 1916
rect 3115 1836 3119 1916
rect 3123 1836 3125 1916
rect 3272 1908 3281 1916
rect 3229 1868 3231 1908
rect 3235 1868 3237 1908
rect 3249 1868 3251 1908
rect 3241 1828 3251 1868
rect 3255 1828 3261 1908
rect 3265 1844 3267 1908
rect 3279 1844 3281 1908
rect 3265 1836 3281 1844
rect 3285 1836 3291 1916
rect 3295 1836 3297 1916
rect 3403 1876 3405 1916
rect 3409 1876 3411 1916
rect 3265 1828 3273 1836
rect 3489 1836 3491 1916
rect 3495 1836 3501 1916
rect 3505 1836 3507 1916
rect 3529 1836 3531 1916
rect 3535 1836 3541 1916
rect 3545 1836 3547 1916
rect 3668 1876 3670 1916
rect 3674 1876 3678 1916
rect 3690 1836 3692 1916
rect 3696 1836 3700 1916
rect 3704 1836 3706 1916
rect 3828 1876 3830 1916
rect 3834 1876 3838 1916
rect 3850 1836 3852 1916
rect 3856 1836 3860 1916
rect 3864 1836 3866 1916
rect 3954 1836 3956 1916
rect 3960 1836 3964 1916
rect 3968 1836 3970 1916
rect 3982 1876 3986 1916
rect 3990 1876 3992 1916
rect 4103 1876 4105 1916
rect 4109 1876 4111 1916
rect 4123 1876 4125 1916
rect 4129 1876 4131 1916
rect 4223 1836 4225 1916
rect 4229 1904 4245 1916
rect 4229 1836 4231 1904
rect 4243 1836 4245 1904
rect 4249 1838 4251 1916
rect 4263 1838 4265 1916
rect 4249 1836 4265 1838
rect 4269 1850 4271 1916
rect 4283 1850 4285 1916
rect 4269 1836 4285 1850
rect 4289 1838 4291 1916
rect 4383 1876 4385 1916
rect 4389 1876 4391 1916
rect 4403 1876 4405 1916
rect 4409 1876 4411 1916
rect 4289 1836 4303 1838
rect 4494 1836 4496 1916
rect 4500 1836 4504 1916
rect 4508 1836 4510 1916
rect 4522 1876 4526 1916
rect 4530 1876 4532 1916
rect 4639 1836 4641 1916
rect 4645 1836 4647 1916
rect 4659 1876 4663 1916
rect 4667 1876 4671 1916
rect 4683 1876 4685 1916
rect 4689 1876 4691 1916
rect 4795 1836 4797 1916
rect 4801 1836 4805 1916
rect 4809 1836 4811 1916
rect 4903 1876 4905 1916
rect 4909 1876 4911 1916
rect 4923 1876 4925 1916
rect 4929 1876 4931 1916
rect 5023 1836 5025 1916
rect 5029 1904 5045 1916
rect 5029 1836 5031 1904
rect 5043 1836 5045 1904
rect 5049 1838 5051 1916
rect 5063 1838 5065 1916
rect 5049 1836 5065 1838
rect 5069 1850 5071 1916
rect 5083 1850 5085 1916
rect 5069 1836 5085 1850
rect 5089 1838 5091 1916
rect 5183 1876 5185 1916
rect 5189 1876 5191 1916
rect 5089 1836 5103 1838
rect 5295 1836 5297 1916
rect 5301 1836 5305 1916
rect 5309 1836 5311 1916
rect 5394 1836 5396 1916
rect 5400 1836 5404 1916
rect 5408 1836 5410 1916
rect 5422 1876 5426 1916
rect 5430 1876 5432 1916
rect 5548 1876 5550 1916
rect 5554 1876 5558 1916
rect 5570 1836 5572 1916
rect 5576 1836 5580 1916
rect 5584 1836 5586 1916
rect 5657 1914 5671 1916
rect 5669 1836 5671 1914
rect 5675 1836 5677 1916
rect 5689 1836 5691 1916
rect 5695 1836 5697 1916
rect 357 1536 371 1544
rect 89 1464 91 1504
rect 95 1464 97 1504
rect 109 1464 111 1504
rect 115 1500 131 1504
rect 115 1464 117 1500
rect 129 1464 131 1500
rect 135 1464 137 1504
rect 243 1464 245 1504
rect 249 1500 265 1504
rect 249 1464 251 1500
rect 263 1464 265 1500
rect 269 1464 271 1504
rect 283 1464 285 1504
rect 289 1464 291 1504
rect 369 1464 371 1536
rect 375 1532 391 1544
rect 375 1464 377 1532
rect 389 1464 391 1532
rect 395 1464 397 1544
rect 409 1464 411 1544
rect 415 1464 417 1544
rect 523 1464 525 1544
rect 529 1464 531 1544
rect 543 1464 545 1544
rect 549 1532 565 1544
rect 549 1464 551 1532
rect 563 1464 565 1532
rect 569 1536 583 1544
rect 569 1464 571 1536
rect 649 1464 651 1504
rect 655 1464 657 1504
rect 669 1464 671 1504
rect 675 1464 677 1504
rect 769 1464 771 1504
rect 775 1464 777 1504
rect 888 1464 890 1504
rect 894 1464 898 1504
rect 910 1464 912 1544
rect 916 1464 920 1544
rect 924 1464 926 1544
rect 1023 1464 1025 1504
rect 1029 1500 1045 1504
rect 1029 1464 1031 1500
rect 1043 1464 1045 1500
rect 1049 1464 1051 1504
rect 1063 1464 1065 1504
rect 1069 1464 1071 1504
rect 1163 1464 1165 1504
rect 1169 1464 1171 1504
rect 1183 1464 1185 1504
rect 1189 1464 1191 1504
rect 1289 1464 1291 1544
rect 1295 1464 1299 1544
rect 1303 1464 1305 1544
rect 1421 1464 1423 1544
rect 1427 1464 1429 1544
rect 1637 1542 1651 1544
rect 1441 1464 1445 1504
rect 1449 1464 1451 1504
rect 1563 1464 1565 1504
rect 1569 1464 1571 1504
rect 1649 1464 1651 1542
rect 1655 1530 1671 1544
rect 1655 1464 1657 1530
rect 1669 1464 1671 1530
rect 1675 1542 1691 1544
rect 1675 1464 1677 1542
rect 1689 1464 1691 1542
rect 1695 1476 1697 1544
rect 1709 1476 1711 1544
rect 1695 1464 1711 1476
rect 1715 1464 1717 1544
rect 1777 1464 1779 1504
rect 1783 1464 1785 1504
rect 1822 1464 1824 1504
rect 1828 1464 1830 1504
rect 1842 1464 1844 1504
rect 1848 1464 1850 1504
rect 1862 1464 1864 1504
rect 1868 1464 1870 1504
rect 1882 1464 1884 1504
rect 1888 1464 1890 1504
rect 1927 1464 1929 1484
rect 1933 1464 1935 1484
rect 1947 1464 1949 1484
rect 1953 1464 1955 1484
rect 1992 1464 1994 1504
rect 1998 1464 2000 1504
rect 2012 1464 2014 1504
rect 2018 1464 2020 1504
rect 2057 1464 2059 1504
rect 2063 1484 2075 1504
rect 2130 1487 2144 1504
rect 2063 1464 2065 1484
rect 2077 1464 2079 1484
rect 2083 1464 2085 1484
rect 2097 1464 2099 1484
rect 2103 1464 2105 1484
rect 2142 1464 2144 1487
rect 2148 1464 2150 1504
rect 2162 1464 2164 1504
rect 2168 1464 2170 1504
rect 2182 1464 2184 1504
rect 2188 1464 2190 1504
rect 2202 1464 2204 1504
rect 2208 1464 2210 1504
rect 2314 1464 2316 1544
rect 2320 1464 2324 1544
rect 2328 1464 2330 1544
rect 2342 1464 2346 1504
rect 2350 1464 2352 1504
rect 2449 1464 2451 1504
rect 2455 1464 2457 1504
rect 2469 1464 2471 1504
rect 2475 1464 2477 1504
rect 2588 1464 2590 1504
rect 2594 1464 2598 1504
rect 2610 1464 2612 1544
rect 2616 1464 2620 1544
rect 2624 1464 2626 1544
rect 2723 1464 2725 1504
rect 2729 1464 2731 1504
rect 2743 1464 2745 1504
rect 2749 1464 2751 1504
rect 2848 1464 2850 1504
rect 2854 1464 2858 1504
rect 2870 1464 2872 1544
rect 2876 1464 2880 1544
rect 2884 1464 2886 1544
rect 2988 1464 2990 1504
rect 2994 1464 2998 1504
rect 3010 1464 3012 1544
rect 3016 1464 3020 1544
rect 3024 1464 3026 1544
rect 3070 1464 3072 1504
rect 3076 1464 3078 1504
rect 3090 1464 3092 1504
rect 3096 1464 3098 1504
rect 3110 1464 3112 1504
rect 3116 1464 3118 1504
rect 3130 1464 3132 1504
rect 3136 1487 3150 1504
rect 3136 1464 3138 1487
rect 3205 1484 3217 1504
rect 3175 1464 3177 1484
rect 3181 1464 3183 1484
rect 3195 1464 3197 1484
rect 3201 1464 3203 1484
rect 3215 1464 3217 1484
rect 3221 1464 3223 1504
rect 3260 1464 3262 1504
rect 3266 1464 3268 1504
rect 3280 1464 3282 1504
rect 3286 1464 3288 1504
rect 3325 1464 3327 1484
rect 3331 1464 3333 1484
rect 3345 1464 3347 1484
rect 3351 1464 3353 1484
rect 3390 1464 3392 1504
rect 3396 1464 3398 1504
rect 3410 1464 3412 1504
rect 3416 1464 3418 1504
rect 3430 1464 3432 1504
rect 3436 1464 3438 1504
rect 3450 1464 3452 1504
rect 3456 1464 3458 1504
rect 3495 1464 3497 1504
rect 3501 1464 3503 1504
rect 3603 1464 3605 1544
rect 3609 1464 3611 1544
rect 3623 1464 3625 1544
rect 3629 1532 3645 1544
rect 3629 1464 3631 1532
rect 3643 1464 3645 1532
rect 3649 1536 3663 1544
rect 3649 1464 3651 1536
rect 3734 1464 3736 1544
rect 3740 1464 3744 1544
rect 3748 1464 3750 1544
rect 3762 1464 3766 1504
rect 3770 1464 3772 1504
rect 3881 1464 3883 1544
rect 3887 1464 3889 1544
rect 3901 1464 3905 1504
rect 3909 1464 3911 1504
rect 3999 1464 4001 1544
rect 4005 1464 4007 1544
rect 4019 1464 4023 1504
rect 4027 1464 4031 1504
rect 4043 1464 4045 1504
rect 4049 1464 4051 1504
rect 4129 1464 4131 1504
rect 4135 1464 4137 1504
rect 4149 1464 4151 1504
rect 4155 1464 4157 1504
rect 4263 1464 4265 1544
rect 4269 1476 4271 1544
rect 4283 1476 4285 1544
rect 4269 1464 4285 1476
rect 4289 1542 4305 1544
rect 4289 1464 4291 1542
rect 4303 1464 4305 1542
rect 4309 1530 4325 1544
rect 4309 1464 4311 1530
rect 4323 1464 4325 1530
rect 4329 1542 4343 1544
rect 4329 1464 4331 1542
rect 4423 1464 4425 1544
rect 4429 1476 4431 1544
rect 4443 1476 4445 1544
rect 4429 1464 4445 1476
rect 4449 1542 4465 1544
rect 4449 1464 4451 1542
rect 4463 1464 4465 1542
rect 4469 1530 4485 1544
rect 4469 1464 4471 1530
rect 4483 1464 4485 1530
rect 4489 1542 4503 1544
rect 4489 1464 4491 1542
rect 4577 1542 4591 1544
rect 4589 1464 4591 1542
rect 4595 1530 4611 1544
rect 4595 1464 4597 1530
rect 4609 1464 4611 1530
rect 4615 1542 4631 1544
rect 4615 1464 4617 1542
rect 4629 1464 4631 1542
rect 4635 1476 4637 1544
rect 4649 1476 4651 1544
rect 4635 1464 4651 1476
rect 4655 1464 4657 1544
rect 4749 1464 4751 1504
rect 4755 1464 4757 1504
rect 4769 1464 4771 1504
rect 4775 1464 4777 1504
rect 4874 1464 4876 1544
rect 4880 1464 4884 1544
rect 4888 1464 4890 1544
rect 4902 1464 4906 1504
rect 4910 1464 4912 1504
rect 5019 1464 5021 1544
rect 5025 1464 5027 1544
rect 5297 1542 5311 1544
rect 5039 1464 5043 1504
rect 5047 1464 5051 1504
rect 5063 1464 5065 1504
rect 5069 1464 5071 1504
rect 5169 1464 5171 1504
rect 5175 1464 5177 1504
rect 5189 1464 5191 1504
rect 5195 1500 5211 1504
rect 5195 1464 5197 1500
rect 5209 1464 5211 1500
rect 5215 1464 5217 1504
rect 5309 1464 5311 1542
rect 5315 1530 5331 1544
rect 5315 1464 5317 1530
rect 5329 1464 5331 1530
rect 5335 1542 5351 1544
rect 5335 1464 5337 1542
rect 5349 1464 5351 1542
rect 5355 1476 5357 1544
rect 5369 1476 5371 1544
rect 5355 1464 5371 1476
rect 5375 1464 5377 1544
rect 5469 1464 5471 1504
rect 5475 1464 5477 1504
rect 5489 1464 5491 1504
rect 5495 1464 5497 1504
rect 5589 1464 5591 1504
rect 5595 1464 5597 1504
rect 5609 1464 5611 1504
rect 5615 1500 5631 1504
rect 5615 1464 5617 1500
rect 5629 1464 5631 1500
rect 5635 1464 5637 1504
rect 5763 1464 5765 1544
rect 5769 1464 5771 1544
rect 83 1396 85 1436
rect 89 1400 91 1436
rect 103 1400 105 1436
rect 89 1396 105 1400
rect 109 1396 111 1436
rect 123 1396 125 1436
rect 129 1396 131 1436
rect 209 1364 211 1436
rect 197 1356 211 1364
rect 215 1368 217 1436
rect 229 1368 231 1436
rect 215 1356 231 1368
rect 235 1356 237 1436
rect 249 1356 251 1436
rect 255 1356 257 1436
rect 363 1396 365 1436
rect 369 1400 371 1436
rect 383 1400 385 1436
rect 369 1396 385 1400
rect 389 1396 391 1436
rect 403 1396 405 1436
rect 409 1396 411 1436
rect 508 1396 510 1436
rect 514 1396 518 1436
rect 530 1356 532 1436
rect 536 1356 540 1436
rect 544 1356 546 1436
rect 648 1396 650 1436
rect 654 1396 658 1436
rect 670 1356 672 1436
rect 676 1356 680 1436
rect 684 1356 686 1436
rect 799 1356 801 1436
rect 805 1356 807 1436
rect 819 1396 823 1436
rect 827 1396 831 1436
rect 843 1396 845 1436
rect 849 1396 851 1436
rect 929 1396 931 1436
rect 935 1396 937 1436
rect 949 1396 951 1436
rect 955 1396 957 1436
rect 1063 1396 1065 1436
rect 1069 1396 1071 1436
rect 1149 1396 1151 1436
rect 1155 1396 1157 1436
rect 1169 1396 1171 1436
rect 1175 1400 1177 1436
rect 1189 1400 1191 1436
rect 1175 1396 1191 1400
rect 1195 1396 1197 1436
rect 1289 1396 1291 1436
rect 1295 1396 1297 1436
rect 1309 1396 1311 1436
rect 1315 1396 1317 1436
rect 1423 1396 1425 1436
rect 1429 1396 1431 1436
rect 1443 1396 1445 1436
rect 1449 1396 1451 1436
rect 1543 1396 1545 1436
rect 1549 1396 1551 1436
rect 1563 1396 1565 1436
rect 1569 1396 1571 1436
rect 1683 1396 1685 1436
rect 1689 1400 1691 1436
rect 1703 1400 1705 1436
rect 1689 1396 1705 1400
rect 1709 1396 1711 1436
rect 1723 1396 1725 1436
rect 1729 1396 1731 1436
rect 1809 1396 1811 1436
rect 1815 1396 1817 1436
rect 1829 1396 1831 1436
rect 1835 1396 1837 1436
rect 1943 1396 1945 1436
rect 1949 1400 1951 1436
rect 1963 1400 1965 1436
rect 1949 1396 1965 1400
rect 1969 1396 1971 1436
rect 1983 1396 1985 1436
rect 1989 1396 1991 1436
rect 2083 1396 2085 1436
rect 2089 1396 2091 1436
rect 2203 1396 2205 1436
rect 2209 1400 2211 1436
rect 2223 1400 2225 1436
rect 2209 1396 2225 1400
rect 2229 1396 2231 1436
rect 2243 1396 2245 1436
rect 2249 1396 2251 1436
rect 2343 1396 2345 1436
rect 2349 1400 2351 1436
rect 2363 1400 2365 1436
rect 2349 1396 2365 1400
rect 2369 1396 2371 1436
rect 2383 1396 2385 1436
rect 2389 1396 2391 1436
rect 2469 1396 2471 1436
rect 2475 1396 2477 1436
rect 2608 1396 2610 1436
rect 2614 1396 2618 1436
rect 2630 1356 2632 1436
rect 2636 1356 2640 1436
rect 2644 1356 2646 1436
rect 2729 1364 2731 1436
rect 2717 1356 2731 1364
rect 2735 1368 2737 1436
rect 2749 1368 2751 1436
rect 2735 1356 2751 1368
rect 2755 1356 2757 1436
rect 2769 1356 2771 1436
rect 2775 1356 2777 1436
rect 2888 1396 2890 1436
rect 2894 1396 2898 1436
rect 2910 1356 2912 1436
rect 2916 1356 2920 1436
rect 2924 1356 2926 1436
rect 3028 1396 3030 1436
rect 3034 1396 3038 1436
rect 3050 1356 3052 1436
rect 3056 1356 3060 1436
rect 3064 1356 3066 1436
rect 3168 1396 3170 1436
rect 3174 1396 3178 1436
rect 3190 1356 3192 1436
rect 3196 1356 3200 1436
rect 3204 1356 3206 1436
rect 3303 1396 3305 1436
rect 3309 1396 3311 1436
rect 3389 1396 3391 1436
rect 3395 1396 3397 1436
rect 3501 1356 3503 1436
rect 3507 1356 3509 1436
rect 3521 1396 3525 1436
rect 3529 1396 3531 1436
rect 3643 1356 3645 1436
rect 3649 1356 3651 1436
rect 3663 1356 3665 1436
rect 3669 1368 3671 1436
rect 3683 1368 3685 1436
rect 3669 1356 3685 1368
rect 3689 1364 3691 1436
rect 3689 1356 3703 1364
rect 3774 1356 3776 1436
rect 3780 1356 3784 1436
rect 3788 1356 3790 1436
rect 3802 1396 3806 1436
rect 3810 1396 3812 1436
rect 3923 1396 3925 1436
rect 3929 1396 3931 1436
rect 4028 1396 4030 1436
rect 4034 1396 4038 1436
rect 4050 1356 4052 1436
rect 4056 1356 4060 1436
rect 4064 1356 4066 1436
rect 4168 1396 4170 1436
rect 4174 1396 4178 1436
rect 4190 1356 4192 1436
rect 4196 1356 4200 1436
rect 4204 1356 4206 1436
rect 4303 1356 4305 1436
rect 4309 1356 4311 1436
rect 4323 1356 4325 1436
rect 4329 1368 4331 1436
rect 4343 1368 4345 1436
rect 4329 1356 4345 1368
rect 4349 1364 4351 1436
rect 4448 1396 4450 1436
rect 4454 1396 4458 1436
rect 4349 1356 4363 1364
rect 4470 1356 4472 1436
rect 4476 1356 4480 1436
rect 4484 1356 4486 1436
rect 4594 1356 4596 1436
rect 4600 1356 4604 1436
rect 4608 1356 4610 1436
rect 4622 1396 4626 1436
rect 4630 1396 4632 1436
rect 4729 1396 4731 1436
rect 4735 1396 4737 1436
rect 4749 1396 4751 1436
rect 4755 1396 4757 1436
rect 4854 1356 4856 1436
rect 4860 1356 4864 1436
rect 4868 1356 4870 1436
rect 4882 1396 4886 1436
rect 4890 1396 4892 1436
rect 4989 1356 4991 1436
rect 4995 1356 4999 1436
rect 5003 1356 5005 1436
rect 5109 1396 5111 1436
rect 5115 1396 5117 1436
rect 5129 1396 5131 1436
rect 5135 1396 5137 1436
rect 5243 1396 5245 1436
rect 5249 1396 5251 1436
rect 5263 1396 5265 1436
rect 5269 1396 5271 1436
rect 5368 1396 5370 1436
rect 5374 1396 5378 1436
rect 5390 1356 5392 1436
rect 5396 1356 5400 1436
rect 5404 1356 5406 1436
rect 5494 1356 5496 1436
rect 5500 1356 5504 1436
rect 5508 1356 5510 1436
rect 5522 1396 5526 1436
rect 5530 1396 5532 1436
rect 5654 1356 5656 1436
rect 5660 1356 5664 1436
rect 5668 1356 5670 1436
rect 5682 1396 5686 1436
rect 5690 1396 5692 1436
rect 157 1056 171 1064
rect 83 984 85 1024
rect 89 984 91 1024
rect 169 984 171 1056
rect 175 1052 191 1064
rect 175 984 177 1052
rect 189 984 191 1052
rect 195 984 197 1064
rect 209 984 211 1064
rect 215 984 217 1064
rect 314 984 316 1064
rect 320 984 324 1064
rect 328 984 330 1064
rect 342 984 346 1024
rect 350 984 352 1024
rect 454 984 456 1064
rect 460 984 464 1064
rect 468 984 470 1064
rect 482 984 486 1024
rect 490 984 492 1024
rect 603 984 605 1024
rect 609 1020 625 1024
rect 609 984 611 1020
rect 623 984 625 1020
rect 629 984 631 1024
rect 643 984 645 1024
rect 649 984 651 1024
rect 734 984 736 1064
rect 740 984 744 1064
rect 748 984 750 1064
rect 877 1056 891 1064
rect 762 984 766 1024
rect 770 984 772 1024
rect 889 984 891 1056
rect 895 1052 911 1064
rect 895 984 897 1052
rect 909 984 911 1052
rect 915 984 917 1064
rect 929 984 931 1064
rect 935 984 937 1064
rect 1048 984 1050 1024
rect 1054 984 1058 1024
rect 1070 984 1072 1064
rect 1076 984 1080 1064
rect 1084 984 1086 1064
rect 1257 1056 1271 1064
rect 1183 984 1185 1024
rect 1189 984 1191 1024
rect 1269 984 1271 1056
rect 1275 1052 1291 1064
rect 1275 984 1277 1052
rect 1289 984 1291 1052
rect 1295 984 1297 1064
rect 1309 984 1311 1064
rect 1315 984 1317 1064
rect 1423 984 1425 1024
rect 1429 984 1431 1024
rect 1535 984 1537 1064
rect 1541 984 1545 1064
rect 1549 984 1551 1064
rect 1649 984 1651 1024
rect 1655 984 1657 1024
rect 1763 984 1765 1024
rect 1769 1020 1785 1024
rect 1769 984 1771 1020
rect 1783 984 1785 1020
rect 1789 984 1791 1024
rect 1803 984 1805 1024
rect 1809 984 1811 1024
rect 1903 984 1905 1024
rect 1909 984 1911 1024
rect 1923 984 1925 1024
rect 1929 984 1931 1024
rect 2028 984 2030 1024
rect 2034 984 2038 1024
rect 2050 984 2052 1064
rect 2056 984 2060 1064
rect 2064 984 2066 1064
rect 2163 984 2165 1024
rect 2169 1020 2185 1024
rect 2169 984 2171 1020
rect 2183 984 2185 1020
rect 2189 984 2191 1024
rect 2203 984 2205 1024
rect 2209 984 2211 1024
rect 2303 984 2305 1024
rect 2309 1020 2325 1024
rect 2309 984 2311 1020
rect 2323 984 2325 1020
rect 2329 984 2331 1024
rect 2343 984 2345 1024
rect 2349 984 2351 1024
rect 2448 984 2450 1024
rect 2454 984 2458 1024
rect 2470 984 2472 1064
rect 2476 984 2480 1064
rect 2484 984 2486 1064
rect 2583 984 2585 1024
rect 2589 1020 2605 1024
rect 2589 984 2591 1020
rect 2603 984 2605 1020
rect 2609 984 2611 1024
rect 2623 984 2625 1024
rect 2629 984 2631 1024
rect 2729 984 2731 1024
rect 2735 984 2737 1024
rect 2829 984 2831 1064
rect 2835 984 2839 1064
rect 2843 984 2845 1064
rect 2949 984 2951 1064
rect 2955 984 2959 1064
rect 2963 984 2965 1064
rect 3069 984 3071 1024
rect 3075 984 3077 1024
rect 3089 984 3093 1024
rect 3097 984 3101 1024
rect 3113 984 3115 1064
rect 3119 984 3121 1064
rect 3235 984 3237 1064
rect 3241 984 3245 1064
rect 3249 984 3251 1064
rect 3375 984 3377 1064
rect 3381 984 3385 1064
rect 3389 984 3391 1064
rect 3483 984 3485 1024
rect 3489 984 3491 1024
rect 3588 984 3590 1024
rect 3594 984 3598 1024
rect 3610 984 3612 1064
rect 3616 984 3620 1064
rect 3624 984 3626 1064
rect 3728 984 3730 1024
rect 3734 984 3738 1024
rect 3750 984 3752 1064
rect 3756 984 3760 1064
rect 3764 984 3766 1064
rect 3849 984 3851 1024
rect 3855 984 3857 1024
rect 3869 984 3871 1024
rect 3875 984 3877 1024
rect 3969 984 3971 1024
rect 3975 984 3977 1024
rect 3989 984 3991 1024
rect 3995 984 3997 1024
rect 4089 984 4091 1064
rect 4095 984 4099 1064
rect 4103 984 4105 1064
rect 4209 984 4211 1024
rect 4215 984 4217 1024
rect 4323 984 4325 1064
rect 4329 984 4331 1064
rect 4343 984 4345 1064
rect 4349 1052 4365 1064
rect 4349 984 4351 1052
rect 4363 984 4365 1052
rect 4369 1056 4383 1064
rect 4369 984 4371 1056
rect 4488 984 4490 1024
rect 4494 984 4498 1024
rect 4510 984 4512 1064
rect 4516 984 4520 1064
rect 4524 984 4526 1064
rect 4623 984 4625 1064
rect 4629 984 4631 1064
rect 4643 984 4645 1064
rect 4649 1052 4665 1064
rect 4649 984 4651 1052
rect 4663 984 4665 1052
rect 4669 1056 4683 1064
rect 4669 984 4671 1056
rect 4754 984 4756 1064
rect 4760 984 4764 1064
rect 4768 984 4770 1064
rect 4782 984 4786 1024
rect 4790 984 4792 1024
rect 4889 984 4891 1024
rect 4895 984 4899 1024
rect 4911 984 4913 1064
rect 4917 984 4919 1064
rect 5009 984 5011 1024
rect 5015 984 5017 1024
rect 5109 984 5111 1024
rect 5115 984 5117 1024
rect 5223 984 5225 1024
rect 5229 984 5231 1024
rect 5243 984 5245 1024
rect 5249 984 5251 1024
rect 5368 984 5370 1024
rect 5374 984 5378 1024
rect 5390 984 5392 1064
rect 5396 984 5400 1064
rect 5404 984 5406 1064
rect 5489 984 5491 1064
rect 5495 984 5499 1064
rect 5503 984 5505 1064
rect 5623 984 5625 1024
rect 5629 1020 5645 1024
rect 5629 984 5631 1020
rect 5643 984 5645 1020
rect 5649 984 5651 1024
rect 5663 984 5665 1024
rect 5669 984 5671 1024
rect 5763 984 5765 1024
rect 5769 984 5771 1024
rect 83 916 85 956
rect 89 920 91 956
rect 103 920 105 956
rect 89 916 105 920
rect 109 916 111 956
rect 123 916 125 956
rect 129 916 131 956
rect 209 884 211 956
rect 197 876 211 884
rect 215 888 217 956
rect 229 888 231 956
rect 215 876 231 888
rect 235 876 237 956
rect 249 876 251 956
rect 255 876 257 956
rect 363 916 365 956
rect 369 920 371 956
rect 383 920 385 956
rect 369 916 385 920
rect 389 916 391 956
rect 403 916 405 956
rect 409 916 411 956
rect 503 876 505 956
rect 509 876 511 956
rect 523 876 525 956
rect 529 888 531 956
rect 543 888 545 956
rect 529 876 545 888
rect 549 884 551 956
rect 643 916 645 956
rect 649 920 651 956
rect 663 920 665 956
rect 649 916 665 920
rect 669 916 671 956
rect 683 916 685 956
rect 689 916 691 956
rect 549 876 563 884
rect 769 884 771 956
rect 757 876 771 884
rect 775 888 777 956
rect 789 888 791 956
rect 775 876 791 888
rect 795 876 797 956
rect 809 876 811 956
rect 815 876 817 956
rect 928 916 930 956
rect 934 916 938 956
rect 950 876 952 956
rect 956 876 960 956
rect 964 876 966 956
rect 1063 916 1065 956
rect 1069 920 1071 956
rect 1083 920 1085 956
rect 1069 916 1085 920
rect 1089 916 1091 956
rect 1103 916 1105 956
rect 1109 916 1111 956
rect 1194 876 1196 956
rect 1200 876 1204 956
rect 1208 876 1210 956
rect 1222 916 1226 956
rect 1230 916 1232 956
rect 1343 916 1345 956
rect 1349 920 1351 956
rect 1363 920 1365 956
rect 1349 916 1365 920
rect 1369 916 1371 956
rect 1383 916 1385 956
rect 1389 916 1391 956
rect 1469 916 1471 956
rect 1475 916 1477 956
rect 1569 916 1571 956
rect 1575 916 1577 956
rect 1589 916 1591 956
rect 1595 916 1597 956
rect 1723 916 1725 956
rect 1729 920 1731 956
rect 1743 920 1745 956
rect 1729 916 1745 920
rect 1749 916 1751 956
rect 1763 916 1765 956
rect 1769 916 1771 956
rect 1863 916 1865 956
rect 1869 920 1871 956
rect 1883 920 1885 956
rect 1869 916 1885 920
rect 1889 916 1891 956
rect 1903 916 1905 956
rect 1909 916 1911 956
rect 1989 916 1991 956
rect 1995 916 1997 956
rect 2009 916 2011 956
rect 2015 920 2017 956
rect 2029 920 2031 956
rect 2015 916 2031 920
rect 2035 916 2037 956
rect 2134 876 2136 956
rect 2140 876 2144 956
rect 2148 876 2150 956
rect 2162 916 2166 956
rect 2170 916 2172 956
rect 2269 916 2271 956
rect 2275 916 2277 956
rect 2289 916 2293 956
rect 2297 916 2301 956
rect 2313 876 2315 956
rect 2319 876 2321 956
rect 2409 916 2411 956
rect 2415 916 2417 956
rect 2523 916 2525 956
rect 2529 916 2531 956
rect 2543 916 2545 956
rect 2549 916 2551 956
rect 2653 877 2655 956
rect 2641 876 2655 877
rect 2659 877 2661 956
rect 2673 877 2675 956
rect 2659 876 2675 877
rect 2679 876 2685 956
rect 2689 876 2691 956
rect 2769 916 2771 956
rect 2775 916 2777 956
rect 2789 916 2791 956
rect 2795 916 2797 956
rect 2903 916 2905 956
rect 2909 916 2911 956
rect 2923 916 2925 956
rect 2929 916 2931 956
rect 3029 916 3031 956
rect 3035 916 3037 956
rect 3143 916 3145 956
rect 3149 916 3151 956
rect 3263 916 3265 956
rect 3269 916 3271 956
rect 3283 916 3285 956
rect 3289 916 3291 956
rect 3415 876 3417 956
rect 3421 876 3425 956
rect 3429 876 3431 956
rect 3535 876 3537 956
rect 3541 876 3545 956
rect 3549 876 3551 956
rect 3643 876 3645 956
rect 3649 876 3651 956
rect 3663 876 3665 956
rect 3669 888 3671 956
rect 3683 888 3685 956
rect 3669 876 3685 888
rect 3689 884 3691 956
rect 3783 916 3785 956
rect 3789 916 3791 956
rect 3888 916 3890 956
rect 3894 916 3898 956
rect 3689 876 3703 884
rect 3910 876 3912 956
rect 3916 876 3920 956
rect 3924 876 3926 956
rect 4009 916 4011 956
rect 4015 916 4017 956
rect 4029 916 4031 956
rect 4035 916 4037 956
rect 4148 916 4150 956
rect 4154 916 4158 956
rect 4170 876 4172 956
rect 4176 876 4180 956
rect 4184 876 4186 956
rect 4288 916 4290 956
rect 4294 916 4298 956
rect 4310 876 4312 956
rect 4316 876 4320 956
rect 4324 876 4326 956
rect 4429 916 4431 956
rect 4435 916 4437 956
rect 4548 916 4550 956
rect 4554 916 4558 956
rect 4570 876 4572 956
rect 4576 876 4580 956
rect 4584 876 4586 956
rect 4669 884 4671 956
rect 4657 876 4671 884
rect 4675 888 4677 956
rect 4689 888 4691 956
rect 4675 876 4691 888
rect 4695 876 4697 956
rect 4709 876 4711 956
rect 4715 876 4717 956
rect 4821 876 4823 956
rect 4827 876 4829 956
rect 4841 916 4845 956
rect 4849 916 4851 956
rect 4948 916 4950 956
rect 4954 916 4958 956
rect 4970 876 4972 956
rect 4976 876 4980 956
rect 4984 876 4986 956
rect 5069 884 5071 956
rect 5057 876 5071 884
rect 5075 888 5077 956
rect 5089 888 5091 956
rect 5075 876 5091 888
rect 5095 876 5097 956
rect 5109 876 5111 956
rect 5115 876 5117 956
rect 5233 877 5235 956
rect 5221 876 5235 877
rect 5239 877 5241 956
rect 5253 877 5255 956
rect 5239 876 5255 877
rect 5259 876 5265 956
rect 5269 876 5271 956
rect 5383 916 5385 956
rect 5389 916 5391 956
rect 5483 876 5485 956
rect 5489 944 5505 956
rect 5489 876 5491 944
rect 5503 876 5505 944
rect 5509 878 5511 956
rect 5523 878 5525 956
rect 5509 876 5525 878
rect 5529 890 5531 956
rect 5543 890 5545 956
rect 5529 876 5545 890
rect 5549 878 5551 956
rect 5549 876 5563 878
rect 5654 876 5656 956
rect 5660 876 5664 956
rect 5668 876 5670 956
rect 5682 916 5686 956
rect 5690 916 5692 956
rect 83 504 85 544
rect 89 540 105 544
rect 89 504 91 540
rect 103 504 105 540
rect 109 504 111 544
rect 123 504 125 544
rect 129 504 131 544
rect 243 504 245 584
rect 249 504 251 584
rect 263 504 265 584
rect 269 572 285 584
rect 269 504 271 572
rect 283 504 285 572
rect 289 576 303 584
rect 289 504 291 576
rect 383 504 385 544
rect 389 540 405 544
rect 389 504 391 540
rect 403 504 405 540
rect 409 504 411 544
rect 423 504 425 544
rect 429 504 431 544
rect 528 504 530 544
rect 534 504 538 544
rect 550 504 552 584
rect 556 504 560 584
rect 564 504 566 584
rect 637 576 651 584
rect 649 504 651 576
rect 655 572 671 584
rect 655 504 657 572
rect 669 504 671 572
rect 675 504 677 584
rect 689 504 691 584
rect 695 504 697 584
rect 789 504 791 544
rect 795 504 797 544
rect 809 504 811 544
rect 815 504 817 544
rect 948 504 950 544
rect 954 504 958 544
rect 970 504 972 584
rect 976 504 980 584
rect 984 504 986 584
rect 1197 576 1211 584
rect 1083 504 1085 544
rect 1089 540 1105 544
rect 1089 504 1091 540
rect 1103 504 1105 540
rect 1109 504 1111 544
rect 1123 504 1125 544
rect 1129 504 1131 544
rect 1209 504 1211 576
rect 1215 572 1231 584
rect 1215 504 1217 572
rect 1229 504 1231 572
rect 1235 504 1237 584
rect 1249 504 1251 584
rect 1255 504 1257 584
rect 1363 504 1365 584
rect 1369 504 1371 584
rect 1383 504 1385 584
rect 1389 572 1405 584
rect 1389 504 1391 572
rect 1403 504 1405 572
rect 1409 576 1423 584
rect 1409 504 1411 576
rect 1509 504 1511 544
rect 1515 504 1517 544
rect 1529 504 1531 544
rect 1535 540 1551 544
rect 1535 504 1537 540
rect 1549 504 1551 540
rect 1555 504 1557 544
rect 1668 504 1670 544
rect 1674 504 1678 544
rect 1690 504 1692 584
rect 1696 504 1700 584
rect 1704 504 1706 584
rect 1917 576 1931 584
rect 1803 504 1805 544
rect 1809 540 1825 544
rect 1809 504 1811 540
rect 1823 504 1825 540
rect 1829 504 1831 544
rect 1843 504 1845 544
rect 1849 504 1851 544
rect 1929 504 1931 576
rect 1935 572 1951 584
rect 1935 504 1937 572
rect 1949 504 1951 572
rect 1955 504 1957 584
rect 1969 504 1971 584
rect 1975 504 1977 584
rect 2095 504 2097 584
rect 2101 504 2105 584
rect 2109 504 2111 584
rect 2201 583 2215 584
rect 2213 504 2215 583
rect 2219 583 2235 584
rect 2219 504 2221 583
rect 2233 504 2235 583
rect 2239 504 2245 584
rect 2249 504 2251 584
rect 2329 504 2331 544
rect 2335 504 2337 544
rect 2349 504 2353 544
rect 2357 504 2361 544
rect 2373 504 2375 584
rect 2379 504 2381 584
rect 2469 504 2471 544
rect 2475 504 2477 544
rect 2489 504 2491 544
rect 2495 504 2497 544
rect 2603 504 2605 544
rect 2609 504 2611 544
rect 2623 504 2625 544
rect 2629 504 2631 544
rect 2735 504 2737 584
rect 2741 504 2745 584
rect 2749 504 2751 584
rect 2834 504 2836 584
rect 2840 504 2844 584
rect 2848 504 2850 584
rect 3077 576 3091 584
rect 2862 504 2866 544
rect 2870 504 2872 544
rect 2983 504 2985 544
rect 2989 504 2991 544
rect 3003 504 3005 544
rect 3009 504 3011 544
rect 3089 504 3091 576
rect 3095 572 3111 584
rect 3095 504 3097 572
rect 3109 504 3111 572
rect 3115 504 3117 584
rect 3129 504 3131 584
rect 3135 504 3137 584
rect 3243 504 3245 544
rect 3249 540 3265 544
rect 3249 504 3251 540
rect 3263 504 3265 540
rect 3269 504 3271 544
rect 3283 504 3285 544
rect 3289 504 3291 544
rect 3369 504 3371 544
rect 3375 504 3377 544
rect 3389 504 3391 544
rect 3395 504 3397 544
rect 3508 504 3510 544
rect 3514 504 3518 544
rect 3530 504 3532 584
rect 3536 504 3540 584
rect 3544 504 3546 584
rect 3629 504 3631 544
rect 3635 504 3637 544
rect 3649 504 3651 544
rect 3655 504 3657 544
rect 3768 504 3770 544
rect 3774 504 3778 544
rect 3790 504 3792 584
rect 3796 504 3800 584
rect 3804 504 3806 584
rect 3894 504 3896 584
rect 3900 504 3904 584
rect 3908 504 3910 584
rect 4017 576 4031 584
rect 3922 504 3926 544
rect 3930 504 3932 544
rect 4029 504 4031 576
rect 4035 572 4051 584
rect 4035 504 4037 572
rect 4049 504 4051 572
rect 4055 504 4057 584
rect 4069 504 4071 584
rect 4075 504 4077 584
rect 4194 504 4196 584
rect 4200 504 4204 584
rect 4208 504 4210 584
rect 4222 504 4226 544
rect 4230 504 4232 544
rect 4343 504 4345 544
rect 4349 504 4351 544
rect 4443 504 4445 584
rect 4449 504 4451 584
rect 4463 504 4465 584
rect 4469 572 4485 584
rect 4469 504 4471 572
rect 4483 504 4485 572
rect 4489 576 4503 584
rect 4489 504 4491 576
rect 4588 504 4590 544
rect 4594 504 4598 544
rect 4610 504 4612 584
rect 4616 504 4620 584
rect 4624 504 4626 584
rect 4728 504 4730 544
rect 4734 504 4738 544
rect 4750 504 4752 584
rect 4756 504 4760 584
rect 4764 504 4766 584
rect 4874 504 4876 584
rect 4880 504 4884 584
rect 4888 504 4890 584
rect 4902 504 4906 544
rect 4910 504 4912 544
rect 5009 504 5011 544
rect 5015 504 5017 544
rect 5129 504 5131 544
rect 5135 504 5139 544
rect 5151 504 5153 584
rect 5157 504 5159 584
rect 5268 504 5270 544
rect 5274 504 5278 544
rect 5290 504 5292 584
rect 5296 504 5300 584
rect 5304 504 5306 584
rect 5394 504 5396 584
rect 5400 504 5404 584
rect 5408 504 5410 584
rect 5422 504 5426 544
rect 5430 504 5432 544
rect 5548 504 5550 544
rect 5554 504 5558 544
rect 5570 504 5572 584
rect 5576 504 5580 584
rect 5584 504 5586 584
rect 5669 504 5671 584
rect 5675 504 5679 584
rect 5683 504 5685 584
rect 83 436 85 476
rect 89 440 91 476
rect 103 440 105 476
rect 89 436 105 440
rect 109 436 111 476
rect 123 436 125 476
rect 129 436 131 476
rect 228 436 230 476
rect 234 436 238 476
rect 250 396 252 476
rect 256 396 260 476
rect 264 396 266 476
rect 388 436 390 476
rect 394 436 398 476
rect 410 396 412 476
rect 416 396 420 476
rect 424 396 426 476
rect 523 436 525 476
rect 529 440 531 476
rect 543 440 545 476
rect 529 436 545 440
rect 549 436 551 476
rect 563 436 565 476
rect 569 436 571 476
rect 659 396 661 476
rect 665 396 667 476
rect 679 436 683 476
rect 687 436 691 476
rect 703 436 705 476
rect 709 436 711 476
rect 803 436 805 476
rect 809 440 811 476
rect 823 440 825 476
rect 809 436 825 440
rect 829 436 831 476
rect 843 436 845 476
rect 849 436 851 476
rect 943 396 945 476
rect 949 396 951 476
rect 963 396 965 476
rect 969 408 971 476
rect 983 408 985 476
rect 969 396 985 408
rect 989 404 991 476
rect 1069 436 1071 476
rect 1075 436 1077 476
rect 1089 436 1091 476
rect 1095 440 1097 476
rect 1109 440 1111 476
rect 1095 436 1111 440
rect 1115 436 1117 476
rect 989 396 1003 404
rect 1233 397 1235 476
rect 1221 396 1235 397
rect 1239 397 1241 476
rect 1253 397 1255 476
rect 1239 396 1255 397
rect 1259 396 1265 476
rect 1269 396 1271 476
rect 1363 436 1365 476
rect 1369 440 1371 476
rect 1383 440 1385 476
rect 1369 436 1385 440
rect 1389 436 1391 476
rect 1403 436 1405 476
rect 1409 436 1411 476
rect 1523 436 1525 476
rect 1529 436 1531 476
rect 1628 436 1630 476
rect 1634 436 1638 476
rect 1650 396 1652 476
rect 1656 396 1660 476
rect 1664 396 1666 476
rect 1759 396 1761 476
rect 1765 396 1767 476
rect 1779 436 1783 476
rect 1787 436 1791 476
rect 1803 436 1805 476
rect 1809 436 1811 476
rect 1889 396 1891 476
rect 1895 396 1899 476
rect 1903 396 1905 476
rect 2029 436 2031 476
rect 2035 436 2037 476
rect 2148 436 2150 476
rect 2154 436 2158 476
rect 2170 396 2172 476
rect 2176 396 2180 476
rect 2184 396 2186 476
rect 2283 396 2285 476
rect 2289 396 2291 476
rect 2303 396 2305 476
rect 2309 408 2311 476
rect 2323 408 2325 476
rect 2309 396 2325 408
rect 2329 404 2331 476
rect 2423 436 2425 476
rect 2429 436 2431 476
rect 2523 436 2525 476
rect 2529 440 2531 476
rect 2543 440 2545 476
rect 2529 436 2545 440
rect 2549 436 2551 476
rect 2563 436 2565 476
rect 2569 436 2571 476
rect 2329 396 2343 404
rect 2654 396 2656 476
rect 2660 396 2664 476
rect 2668 396 2670 476
rect 2682 436 2686 476
rect 2690 436 2692 476
rect 2803 436 2805 476
rect 2809 436 2811 476
rect 2915 396 2917 476
rect 2921 396 2925 476
rect 2929 396 2931 476
rect 3009 436 3011 476
rect 3015 436 3017 476
rect 3123 396 3125 476
rect 3129 396 3131 476
rect 3143 396 3145 476
rect 3149 408 3151 476
rect 3163 408 3165 476
rect 3149 396 3165 408
rect 3169 404 3171 476
rect 3169 396 3183 404
rect 3269 404 3271 476
rect 3257 396 3271 404
rect 3275 408 3277 476
rect 3289 408 3291 476
rect 3275 396 3291 408
rect 3295 396 3297 476
rect 3309 396 3311 476
rect 3315 396 3317 476
rect 3423 436 3425 476
rect 3429 436 3431 476
rect 3534 396 3536 476
rect 3540 396 3544 476
rect 3548 396 3550 476
rect 3562 436 3566 476
rect 3570 436 3572 476
rect 3669 404 3671 476
rect 3657 396 3671 404
rect 3675 408 3677 476
rect 3689 408 3691 476
rect 3675 396 3691 408
rect 3695 396 3697 476
rect 3709 396 3711 476
rect 3715 396 3717 476
rect 3823 436 3825 476
rect 3829 440 3831 476
rect 3843 440 3845 476
rect 3829 436 3845 440
rect 3849 436 3851 476
rect 3863 436 3865 476
rect 3869 436 3871 476
rect 3949 436 3951 476
rect 3955 436 3957 476
rect 3969 436 3971 476
rect 3975 436 3977 476
rect 4103 436 4105 476
rect 4109 440 4111 476
rect 4123 440 4125 476
rect 4109 436 4125 440
rect 4129 436 4131 476
rect 4143 436 4145 476
rect 4149 436 4151 476
rect 4248 436 4250 476
rect 4254 436 4258 476
rect 4270 396 4272 476
rect 4276 396 4280 476
rect 4284 396 4286 476
rect 4383 436 4385 476
rect 4389 436 4391 476
rect 4483 436 4485 476
rect 4489 436 4491 476
rect 4503 436 4505 476
rect 4509 436 4511 476
rect 4608 436 4610 476
rect 4614 436 4618 476
rect 4630 396 4632 476
rect 4636 396 4640 476
rect 4644 396 4646 476
rect 4743 436 4745 476
rect 4749 436 4751 476
rect 4848 436 4850 476
rect 4854 436 4858 476
rect 4870 396 4872 476
rect 4876 396 4880 476
rect 4884 396 4886 476
rect 5012 468 5021 476
rect 4969 428 4971 468
rect 4975 428 4977 468
rect 4989 428 4991 468
rect 4981 388 4991 428
rect 4995 388 5001 468
rect 5005 404 5007 468
rect 5019 404 5021 468
rect 5005 396 5021 404
rect 5025 396 5031 476
rect 5035 396 5037 476
rect 5148 436 5150 476
rect 5154 436 5158 476
rect 5005 388 5013 396
rect 5170 396 5172 476
rect 5176 396 5180 476
rect 5184 396 5186 476
rect 5294 396 5296 476
rect 5300 396 5304 476
rect 5308 396 5310 476
rect 5322 436 5326 476
rect 5330 436 5332 476
rect 5463 396 5465 476
rect 5469 396 5471 476
rect 5483 396 5485 476
rect 5489 408 5491 476
rect 5503 408 5505 476
rect 5489 396 5505 408
rect 5509 404 5511 476
rect 5509 396 5523 404
rect 5594 396 5596 476
rect 5600 396 5604 476
rect 5608 396 5610 476
rect 5622 436 5626 476
rect 5630 436 5632 476
rect 5729 436 5731 476
rect 5735 436 5737 476
rect 5749 436 5751 476
rect 5755 436 5757 476
rect 197 96 211 104
rect 83 24 85 64
rect 89 60 105 64
rect 89 24 91 60
rect 103 24 105 60
rect 109 24 111 64
rect 123 24 125 64
rect 129 24 131 64
rect 209 24 211 96
rect 215 92 231 104
rect 215 24 217 92
rect 229 24 231 92
rect 235 24 237 104
rect 249 24 251 104
rect 255 24 257 104
rect 383 24 385 104
rect 389 24 391 104
rect 403 24 405 104
rect 409 92 425 104
rect 409 24 411 92
rect 423 24 425 92
rect 429 96 443 104
rect 429 24 431 96
rect 528 24 530 64
rect 534 24 538 64
rect 550 24 552 104
rect 556 24 560 104
rect 564 24 566 104
rect 654 24 656 104
rect 660 24 664 104
rect 668 24 670 104
rect 682 24 686 64
rect 690 24 692 64
rect 803 24 805 64
rect 809 60 825 64
rect 809 24 811 60
rect 823 24 825 60
rect 829 24 831 64
rect 843 24 845 64
rect 849 24 851 64
rect 929 24 931 64
rect 935 24 937 64
rect 1034 24 1036 104
rect 1040 24 1044 104
rect 1048 24 1050 104
rect 1157 96 1171 104
rect 1062 24 1066 64
rect 1070 24 1072 64
rect 1169 24 1171 96
rect 1175 92 1191 104
rect 1175 24 1177 92
rect 1189 24 1191 92
rect 1195 24 1197 104
rect 1209 24 1211 104
rect 1215 24 1217 104
rect 1309 24 1311 104
rect 1315 24 1319 104
rect 1323 24 1325 104
rect 1429 24 1431 64
rect 1435 24 1437 64
rect 1449 24 1453 64
rect 1457 24 1461 64
rect 1473 24 1475 104
rect 1479 24 1481 104
rect 1583 24 1585 64
rect 1589 24 1591 64
rect 1688 24 1690 64
rect 1694 24 1698 64
rect 1710 24 1712 104
rect 1716 24 1720 104
rect 1724 24 1726 104
rect 1823 24 1825 64
rect 1829 24 1831 64
rect 1843 24 1845 64
rect 1849 24 1851 64
rect 1929 24 1931 64
rect 1935 24 1937 64
rect 1949 24 1951 64
rect 1955 60 1971 64
rect 1955 24 1957 60
rect 1969 24 1971 60
rect 1975 24 1977 64
rect 2103 24 2105 64
rect 2109 60 2125 64
rect 2109 24 2111 60
rect 2123 24 2125 60
rect 2129 24 2131 64
rect 2143 24 2145 64
rect 2149 24 2151 64
rect 2229 24 2231 64
rect 2235 24 2239 64
rect 2251 24 2253 104
rect 2257 24 2259 104
rect 2363 24 2365 64
rect 2369 24 2371 64
rect 2383 24 2385 64
rect 2389 24 2391 64
rect 2469 24 2471 64
rect 2475 24 2477 64
rect 2489 24 2493 64
rect 2497 24 2501 64
rect 2513 24 2515 104
rect 2519 24 2521 104
rect 2623 24 2625 104
rect 2629 24 2631 104
rect 2643 24 2645 104
rect 2649 92 2665 104
rect 2649 24 2651 92
rect 2663 24 2665 92
rect 2669 96 2683 104
rect 2669 24 2671 96
rect 2759 24 2761 104
rect 2765 24 2767 104
rect 2779 24 2783 64
rect 2787 24 2791 64
rect 2803 24 2805 64
rect 2809 24 2811 64
rect 2909 24 2911 64
rect 2915 24 2917 64
rect 2929 24 2931 64
rect 2935 24 2937 64
rect 3043 24 3045 64
rect 3049 24 3051 64
rect 3063 24 3065 64
rect 3069 24 3071 64
rect 3163 24 3165 64
rect 3169 60 3185 64
rect 3169 24 3171 60
rect 3183 24 3185 60
rect 3189 24 3191 64
rect 3203 24 3205 64
rect 3209 24 3211 64
rect 3303 24 3305 64
rect 3309 24 3311 64
rect 3394 24 3396 104
rect 3400 24 3404 104
rect 3408 24 3410 104
rect 3422 24 3426 64
rect 3430 24 3432 64
rect 3543 24 3545 64
rect 3549 24 3551 64
rect 3643 24 3645 64
rect 3649 24 3651 64
rect 3663 24 3665 64
rect 3669 24 3671 64
rect 3761 24 3763 104
rect 3767 24 3769 104
rect 3781 24 3785 64
rect 3789 24 3791 64
rect 3869 24 3871 64
rect 3875 24 3879 64
rect 3891 24 3893 104
rect 3897 24 3899 104
rect 4003 24 4005 64
rect 4009 24 4011 64
rect 4023 24 4025 64
rect 4029 24 4031 64
rect 4129 24 4131 64
rect 4135 24 4137 64
rect 4149 24 4153 64
rect 4157 24 4161 64
rect 4173 24 4175 104
rect 4179 24 4181 104
rect 4315 24 4317 104
rect 4321 24 4325 104
rect 4329 24 4331 104
rect 4409 24 4411 64
rect 4415 24 4417 64
rect 4429 24 4431 64
rect 4435 24 4437 64
rect 4543 24 4545 64
rect 4549 60 4565 64
rect 4549 24 4551 60
rect 4563 24 4565 60
rect 4569 24 4571 64
rect 4583 24 4585 64
rect 4589 24 4591 64
rect 4708 24 4710 64
rect 4714 24 4718 64
rect 4730 24 4732 104
rect 4736 24 4740 104
rect 4744 24 4746 104
rect 4829 24 4831 64
rect 4835 24 4837 64
rect 4849 24 4851 64
rect 4855 24 4857 64
rect 4968 24 4970 64
rect 4974 24 4978 64
rect 4990 24 4992 104
rect 4996 24 5000 104
rect 5004 24 5006 104
rect 5089 24 5091 104
rect 5095 24 5099 104
rect 5103 24 5105 104
rect 5341 72 5351 112
rect 5223 24 5225 64
rect 5229 24 5231 64
rect 5243 24 5245 64
rect 5249 24 5251 64
rect 5329 32 5331 72
rect 5335 32 5337 72
rect 5349 32 5351 72
rect 5355 32 5361 112
rect 5365 104 5373 112
rect 5365 96 5381 104
rect 5365 32 5367 96
rect 5379 32 5381 96
rect 5372 24 5381 32
rect 5385 24 5391 104
rect 5395 24 5397 104
rect 5489 24 5491 64
rect 5495 24 5497 64
rect 5603 24 5605 64
rect 5609 24 5611 64
rect 5689 24 5691 64
rect 5695 24 5697 64
rect 5709 24 5711 64
rect 5715 24 5717 64
<< ndcontact >>
rect 71 5544 83 5584
rect 91 5544 103 5584
rect 111 5544 123 5572
rect 131 5544 143 5584
rect 197 5544 209 5584
rect 217 5544 229 5572
rect 237 5544 249 5584
rect 257 5544 269 5584
rect 378 5544 390 5564
rect 400 5544 412 5584
rect 428 5544 440 5584
rect 498 5544 510 5604
rect 534 5544 546 5602
rect 651 5544 663 5584
rect 671 5544 683 5584
rect 691 5544 703 5572
rect 711 5544 723 5584
rect 799 5544 811 5584
rect 829 5544 841 5584
rect 918 5544 930 5564
rect 940 5544 952 5584
rect 968 5544 980 5584
rect 1057 5544 1069 5564
rect 1077 5544 1089 5564
rect 1097 5544 1109 5564
rect 1211 5544 1223 5584
rect 1231 5544 1243 5564
rect 1251 5544 1263 5564
rect 1271 5544 1283 5564
rect 1361 5544 1373 5584
rect 1381 5544 1393 5584
rect 1411 5544 1423 5584
rect 1514 5544 1526 5602
rect 1550 5544 1562 5604
rect 1658 5544 1670 5564
rect 1680 5544 1692 5584
rect 1708 5544 1720 5584
rect 1814 5544 1826 5602
rect 1850 5544 1862 5604
rect 1917 5544 1929 5564
rect 1937 5544 1949 5564
rect 2031 5544 2043 5584
rect 2051 5544 2063 5584
rect 2071 5544 2083 5572
rect 2091 5544 2103 5584
rect 2157 5544 2169 5584
rect 2177 5544 2189 5572
rect 2197 5544 2209 5584
rect 2217 5544 2229 5584
rect 2300 5544 2312 5584
rect 2328 5544 2340 5584
rect 2350 5544 2362 5564
rect 2459 5544 2471 5584
rect 2489 5544 2501 5584
rect 2594 5544 2606 5602
rect 2630 5544 2642 5604
rect 2734 5544 2746 5602
rect 2770 5544 2782 5604
rect 2839 5544 2851 5584
rect 2869 5544 2881 5584
rect 2971 5544 2983 5564
rect 2991 5544 3003 5564
rect 3071 5544 3083 5584
rect 3091 5544 3103 5584
rect 3111 5544 3123 5572
rect 3131 5544 3143 5584
rect 3241 5544 3253 5584
rect 3261 5544 3273 5584
rect 3291 5544 3303 5584
rect 3371 5544 3383 5564
rect 3391 5544 3403 5564
rect 3411 5544 3423 5564
rect 3514 5544 3526 5602
rect 3550 5544 3562 5604
rect 3651 5544 3663 5564
rect 3671 5544 3683 5564
rect 3751 5544 3763 5564
rect 3771 5544 3783 5564
rect 3837 5544 3849 5564
rect 3857 5544 3869 5564
rect 3937 5544 3949 5584
rect 3957 5544 3969 5572
rect 3977 5544 3989 5584
rect 3997 5544 4009 5584
rect 4077 5544 4089 5564
rect 4097 5544 4109 5564
rect 4137 5544 4149 5584
rect 4159 5544 4171 5564
rect 4189 5544 4201 5564
rect 4217 5544 4229 5564
rect 4243 5544 4255 5564
rect 4265 5544 4277 5564
rect 4295 5544 4307 5564
rect 4327 5544 4339 5564
rect 4347 5544 4359 5584
rect 4451 5544 4463 5584
rect 4471 5544 4483 5584
rect 4491 5544 4503 5572
rect 4511 5544 4523 5584
rect 4591 5544 4603 5584
rect 4611 5544 4623 5584
rect 4631 5544 4643 5584
rect 4651 5544 4663 5584
rect 4671 5544 4683 5584
rect 4691 5544 4703 5584
rect 4711 5544 4723 5584
rect 4731 5544 4743 5584
rect 4751 5544 4763 5584
rect 4831 5544 4843 5564
rect 4851 5544 4863 5564
rect 4931 5544 4943 5584
rect 4951 5544 4963 5584
rect 4971 5544 4983 5572
rect 4991 5544 5003 5584
rect 5079 5544 5091 5584
rect 5109 5544 5121 5584
rect 5179 5544 5191 5584
rect 5209 5544 5221 5584
rect 5297 5544 5309 5584
rect 5317 5544 5329 5572
rect 5337 5544 5349 5584
rect 5357 5544 5369 5584
rect 5437 5544 5449 5564
rect 5457 5544 5469 5564
rect 5539 5544 5551 5584
rect 5569 5544 5581 5584
rect 5657 5544 5669 5564
rect 5677 5544 5689 5564
rect 71 5476 83 5516
rect 91 5476 103 5516
rect 111 5488 123 5516
rect 131 5476 143 5516
rect 254 5458 266 5516
rect 290 5456 302 5516
rect 394 5458 406 5516
rect 430 5456 442 5516
rect 534 5458 546 5516
rect 570 5456 582 5516
rect 658 5456 670 5516
rect 694 5458 706 5516
rect 797 5476 809 5516
rect 817 5488 829 5516
rect 837 5476 849 5516
rect 857 5476 869 5516
rect 938 5456 950 5516
rect 974 5458 986 5516
rect 1098 5496 1110 5516
rect 1120 5476 1132 5516
rect 1148 5476 1160 5516
rect 1218 5456 1230 5516
rect 1254 5458 1266 5516
rect 1377 5496 1389 5516
rect 1397 5496 1409 5516
rect 1417 5496 1429 5516
rect 1534 5458 1546 5516
rect 1570 5456 1582 5516
rect 1637 5476 1649 5516
rect 1657 5488 1669 5516
rect 1677 5476 1689 5516
rect 1697 5476 1709 5516
rect 1814 5458 1826 5516
rect 1850 5456 1862 5516
rect 1954 5458 1966 5516
rect 1990 5456 2002 5516
rect 2059 5476 2071 5516
rect 2089 5476 2101 5516
rect 2211 5496 2223 5516
rect 2231 5496 2243 5516
rect 2321 5476 2333 5516
rect 2341 5476 2353 5516
rect 2371 5476 2383 5516
rect 2437 5476 2449 5516
rect 2457 5488 2469 5516
rect 2477 5476 2489 5516
rect 2497 5476 2509 5516
rect 2634 5458 2646 5516
rect 2670 5456 2682 5516
rect 2774 5458 2786 5516
rect 2810 5456 2822 5516
rect 2877 5476 2889 5516
rect 2897 5488 2909 5516
rect 2917 5476 2929 5516
rect 2937 5476 2949 5516
rect 3017 5496 3029 5516
rect 3037 5496 3049 5516
rect 3119 5476 3131 5516
rect 3149 5476 3161 5516
rect 3258 5456 3270 5516
rect 3294 5458 3306 5516
rect 3399 5476 3411 5516
rect 3429 5476 3441 5516
rect 3517 5496 3529 5516
rect 3537 5496 3549 5516
rect 3557 5496 3569 5516
rect 3577 5476 3589 5516
rect 3694 5458 3706 5516
rect 3730 5456 3742 5516
rect 3818 5496 3830 5516
rect 3840 5476 3852 5516
rect 3868 5476 3880 5516
rect 3939 5476 3951 5516
rect 3969 5476 3981 5516
rect 4071 5476 4083 5516
rect 4091 5476 4103 5516
rect 4111 5488 4123 5516
rect 4131 5476 4143 5516
rect 4219 5476 4231 5516
rect 4249 5476 4261 5516
rect 4354 5458 4366 5516
rect 4390 5456 4402 5516
rect 4480 5476 4492 5516
rect 4508 5476 4520 5516
rect 4530 5496 4542 5516
rect 4617 5496 4629 5516
rect 4637 5496 4649 5516
rect 4717 5476 4729 5516
rect 4737 5488 4749 5516
rect 4757 5476 4769 5516
rect 4777 5476 4789 5516
rect 4817 5476 4829 5516
rect 4839 5496 4851 5516
rect 4869 5496 4881 5516
rect 4897 5496 4909 5516
rect 4923 5496 4935 5516
rect 4945 5496 4957 5516
rect 4975 5496 4987 5516
rect 5007 5496 5019 5516
rect 5027 5476 5039 5516
rect 5097 5496 5109 5516
rect 5117 5496 5129 5516
rect 5157 5476 5169 5516
rect 5179 5496 5191 5516
rect 5209 5496 5221 5516
rect 5237 5496 5249 5516
rect 5263 5496 5275 5516
rect 5285 5496 5297 5516
rect 5315 5496 5327 5516
rect 5347 5496 5359 5516
rect 5367 5476 5379 5516
rect 5437 5476 5449 5516
rect 5457 5488 5469 5516
rect 5477 5476 5489 5516
rect 5497 5476 5509 5516
rect 5599 5476 5611 5516
rect 5629 5476 5641 5516
rect 5719 5476 5731 5516
rect 5749 5476 5761 5516
rect 94 5064 106 5122
rect 130 5064 142 5124
rect 200 5064 212 5104
rect 228 5064 240 5104
rect 250 5064 262 5084
rect 337 5064 349 5084
rect 357 5064 369 5084
rect 474 5064 486 5122
rect 510 5064 522 5124
rect 580 5064 592 5104
rect 608 5064 620 5104
rect 630 5064 642 5084
rect 738 5064 750 5084
rect 760 5064 772 5104
rect 788 5064 800 5104
rect 858 5064 870 5124
rect 894 5064 906 5122
rect 1034 5064 1046 5122
rect 1070 5064 1082 5124
rect 1137 5064 1149 5084
rect 1157 5064 1169 5084
rect 1274 5064 1286 5122
rect 1310 5064 1322 5124
rect 1411 5064 1423 5104
rect 1431 5064 1443 5104
rect 1451 5064 1463 5092
rect 1471 5064 1483 5104
rect 1551 5064 1563 5084
rect 1571 5064 1583 5084
rect 1651 5064 1663 5104
rect 1671 5064 1683 5104
rect 1691 5064 1703 5092
rect 1711 5064 1723 5104
rect 1871 5064 1883 5084
rect 1891 5064 1903 5084
rect 1911 5064 1923 5084
rect 1931 5064 1945 5084
rect 2052 5064 2064 5104
rect 2080 5064 2092 5104
rect 2108 5064 2120 5104
rect 2179 5064 2191 5104
rect 2209 5064 2221 5104
rect 2334 5064 2346 5122
rect 2370 5064 2382 5124
rect 2458 5064 2470 5084
rect 2480 5064 2492 5104
rect 2508 5064 2520 5104
rect 2591 5064 2603 5084
rect 2611 5064 2623 5084
rect 2691 5064 2703 5104
rect 2711 5064 2723 5104
rect 2731 5064 2743 5092
rect 2751 5064 2763 5104
rect 2851 5064 2863 5104
rect 2871 5064 2883 5104
rect 2891 5064 2903 5092
rect 2911 5064 2923 5104
rect 3001 5064 3013 5104
rect 3021 5064 3033 5104
rect 3051 5064 3063 5104
rect 3117 5064 3129 5084
rect 3137 5064 3149 5084
rect 3157 5064 3169 5084
rect 3271 5064 3283 5084
rect 3291 5064 3303 5084
rect 3371 5064 3383 5084
rect 3391 5064 3403 5084
rect 3411 5064 3423 5084
rect 3511 5064 3523 5104
rect 3531 5064 3543 5104
rect 3551 5064 3563 5092
rect 3571 5064 3583 5104
rect 3639 5064 3651 5104
rect 3669 5064 3681 5104
rect 3779 5064 3791 5104
rect 3809 5064 3821 5104
rect 3919 5064 3931 5104
rect 3949 5064 3961 5104
rect 4018 5064 4030 5124
rect 4054 5064 4066 5122
rect 4171 5064 4183 5104
rect 4191 5064 4203 5104
rect 4211 5064 4223 5092
rect 4231 5064 4243 5104
rect 4317 5064 4329 5104
rect 4337 5064 4349 5092
rect 4357 5064 4369 5104
rect 4377 5064 4389 5104
rect 4457 5064 4469 5084
rect 4477 5064 4489 5084
rect 4594 5064 4606 5122
rect 4630 5064 4642 5124
rect 4700 5064 4712 5104
rect 4728 5064 4740 5104
rect 4750 5064 4762 5084
rect 4837 5064 4849 5084
rect 4857 5064 4869 5084
rect 4877 5064 4889 5084
rect 4917 5064 4929 5104
rect 4939 5064 4951 5084
rect 4969 5064 4981 5084
rect 4997 5064 5009 5084
rect 5023 5064 5035 5084
rect 5045 5064 5057 5084
rect 5075 5064 5087 5084
rect 5107 5064 5119 5084
rect 5127 5064 5139 5104
rect 5197 5064 5209 5104
rect 5217 5064 5229 5092
rect 5237 5064 5249 5104
rect 5257 5064 5269 5104
rect 5337 5064 5349 5084
rect 5357 5064 5369 5084
rect 5437 5064 5449 5104
rect 5457 5064 5469 5092
rect 5477 5064 5489 5104
rect 5497 5064 5509 5104
rect 5599 5064 5611 5104
rect 5629 5064 5641 5104
rect 5699 5064 5711 5104
rect 5729 5064 5741 5104
rect 71 4996 83 5036
rect 91 4996 103 5036
rect 111 5008 123 5036
rect 131 4996 143 5036
rect 234 4978 246 5036
rect 270 4976 282 5036
rect 338 4976 350 5036
rect 374 4978 386 5036
rect 477 4996 489 5036
rect 497 5008 509 5036
rect 517 4996 529 5036
rect 537 4996 549 5036
rect 639 4996 651 5036
rect 669 4996 681 5036
rect 751 4996 763 5036
rect 771 4996 783 5036
rect 791 5008 803 5036
rect 811 4996 823 5036
rect 891 4996 903 5036
rect 911 4996 923 5036
rect 931 5008 943 5036
rect 951 4996 963 5036
rect 1038 5016 1050 5036
rect 1060 4996 1072 5036
rect 1088 4996 1100 5036
rect 1171 4996 1183 5036
rect 1191 4996 1203 5036
rect 1211 5008 1223 5036
rect 1231 4996 1243 5036
rect 1311 5016 1323 5036
rect 1331 5016 1343 5036
rect 1419 4996 1431 5036
rect 1449 4996 1461 5036
rect 1574 4978 1586 5036
rect 1610 4976 1622 5036
rect 1691 4996 1703 5036
rect 1711 4996 1723 5036
rect 1731 5008 1743 5036
rect 1751 4996 1763 5036
rect 1820 4996 1832 5036
rect 1848 4996 1860 5036
rect 1870 5016 1882 5036
rect 1959 4996 1971 5036
rect 1989 4996 2001 5036
rect 2098 5016 2110 5036
rect 2120 4996 2132 5036
rect 2148 4996 2160 5036
rect 2251 5016 2263 5036
rect 2271 5016 2283 5036
rect 2351 4996 2363 5036
rect 2371 4996 2383 5036
rect 2391 5008 2403 5036
rect 2411 4996 2423 5036
rect 2514 4978 2526 5036
rect 2550 4976 2562 5036
rect 2631 5016 2643 5036
rect 2651 5016 2663 5036
rect 2759 4996 2771 5036
rect 2789 4996 2801 5036
rect 2857 5016 2869 5036
rect 2877 5016 2889 5036
rect 2958 4976 2970 5036
rect 2994 4978 3006 5036
rect 3111 4996 3123 5036
rect 3131 4996 3143 5036
rect 3151 5008 3163 5036
rect 3171 4996 3183 5036
rect 3251 4996 3263 5036
rect 3271 4996 3283 5036
rect 3291 5008 3303 5036
rect 3311 4996 3323 5036
rect 3398 5016 3410 5036
rect 3420 4996 3432 5036
rect 3448 4996 3460 5036
rect 3517 5016 3529 5036
rect 3537 5016 3549 5036
rect 3557 5016 3569 5036
rect 3577 4996 3589 5036
rect 3671 5016 3683 5036
rect 3691 5016 3703 5036
rect 3711 5016 3723 5036
rect 3814 4978 3826 5036
rect 3850 4976 3862 5036
rect 3931 5016 3943 5036
rect 3951 5016 3963 5036
rect 4018 4976 4030 5036
rect 4054 4978 4066 5036
rect 4158 4976 4170 5036
rect 4194 4978 4206 5036
rect 4321 4996 4333 5036
rect 4341 4996 4353 5036
rect 4371 4996 4383 5036
rect 4457 5016 4469 5036
rect 4477 5016 4489 5036
rect 4497 5016 4509 5036
rect 4517 4996 4529 5036
rect 4597 5016 4609 5036
rect 4617 5016 4629 5036
rect 4637 5016 4649 5036
rect 4731 4996 4743 5036
rect 4751 4996 4763 5036
rect 4771 5008 4783 5036
rect 4791 4996 4803 5036
rect 4817 4996 4829 5036
rect 4839 5016 4851 5036
rect 4869 5016 4881 5036
rect 4897 5016 4909 5036
rect 4923 5016 4935 5036
rect 4945 5016 4957 5036
rect 4975 5016 4987 5036
rect 5007 5016 5019 5036
rect 5027 4996 5039 5036
rect 5097 4996 5109 5036
rect 5117 5008 5129 5036
rect 5137 4996 5149 5036
rect 5157 4996 5169 5036
rect 5197 4996 5209 5036
rect 5219 5016 5231 5036
rect 5249 5016 5261 5036
rect 5277 5016 5289 5036
rect 5303 5016 5315 5036
rect 5325 5016 5337 5036
rect 5355 5016 5367 5036
rect 5387 5016 5399 5036
rect 5407 4996 5419 5036
rect 5499 4996 5511 5036
rect 5529 4996 5541 5036
rect 5599 4996 5611 5036
rect 5629 4996 5641 5036
rect 5739 4996 5751 5036
rect 5769 4996 5781 5036
rect 78 4584 90 4604
rect 100 4584 112 4624
rect 128 4584 140 4624
rect 234 4584 246 4642
rect 270 4584 282 4644
rect 340 4584 352 4624
rect 368 4584 380 4624
rect 390 4584 402 4604
rect 479 4584 491 4624
rect 509 4584 521 4624
rect 634 4584 646 4642
rect 670 4584 682 4644
rect 794 4584 806 4642
rect 830 4584 842 4644
rect 897 4584 909 4604
rect 917 4584 929 4604
rect 997 4584 1009 4604
rect 1017 4584 1029 4604
rect 1111 4584 1123 4604
rect 1131 4584 1143 4604
rect 1211 4584 1223 4624
rect 1231 4584 1243 4624
rect 1251 4584 1263 4612
rect 1271 4584 1283 4624
rect 1337 4584 1349 4624
rect 1357 4584 1369 4612
rect 1377 4584 1389 4624
rect 1397 4584 1409 4624
rect 1477 4584 1489 4604
rect 1497 4584 1509 4604
rect 1578 4584 1590 4644
rect 1614 4584 1626 4642
rect 1731 4584 1743 4624
rect 1751 4584 1763 4624
rect 1771 4584 1783 4612
rect 1791 4584 1803 4624
rect 1879 4584 1891 4624
rect 1909 4584 1921 4624
rect 1977 4584 1989 4624
rect 1997 4584 2009 4612
rect 2017 4584 2029 4624
rect 2037 4584 2049 4624
rect 2154 4584 2166 4642
rect 2190 4584 2202 4644
rect 2269 4584 2281 4624
rect 2289 4584 2301 4624
rect 2311 4584 2323 4604
rect 2379 4584 2391 4624
rect 2409 4584 2421 4624
rect 2499 4584 2511 4624
rect 2529 4584 2541 4624
rect 2629 4584 2641 4624
rect 2649 4584 2661 4624
rect 2671 4584 2683 4604
rect 2738 4584 2750 4644
rect 2774 4584 2786 4642
rect 2891 4584 2903 4604
rect 2911 4584 2923 4604
rect 2931 4584 2943 4604
rect 3017 4584 3029 4624
rect 3037 4584 3049 4614
rect 3057 4584 3069 4624
rect 3077 4596 3089 4624
rect 3097 4584 3109 4624
rect 3199 4584 3211 4624
rect 3229 4584 3241 4624
rect 3334 4584 3346 4642
rect 3370 4584 3382 4644
rect 3458 4584 3470 4604
rect 3480 4584 3492 4624
rect 3508 4584 3520 4624
rect 3614 4584 3626 4642
rect 3650 4584 3662 4644
rect 3738 4584 3750 4604
rect 3760 4584 3772 4624
rect 3788 4584 3800 4624
rect 3858 4584 3870 4644
rect 3894 4584 3906 4642
rect 3998 4584 4010 4644
rect 4034 4584 4046 4642
rect 4137 4584 4149 4604
rect 4157 4584 4169 4604
rect 4261 4584 4273 4624
rect 4281 4584 4293 4624
rect 4311 4584 4323 4624
rect 4434 4584 4446 4642
rect 4470 4584 4482 4644
rect 4538 4584 4550 4644
rect 4574 4584 4586 4642
rect 4677 4584 4689 4604
rect 4697 4584 4709 4604
rect 4737 4584 4749 4624
rect 4759 4584 4771 4604
rect 4789 4584 4801 4604
rect 4817 4584 4829 4604
rect 4843 4584 4855 4604
rect 4865 4584 4877 4604
rect 4895 4584 4907 4604
rect 4927 4584 4939 4604
rect 4947 4584 4959 4624
rect 5017 4584 5029 4624
rect 5037 4584 5049 4612
rect 5057 4584 5069 4624
rect 5077 4584 5089 4624
rect 5159 4584 5171 4624
rect 5189 4584 5201 4624
rect 5279 4584 5291 4624
rect 5309 4584 5321 4624
rect 5419 4584 5431 4624
rect 5449 4584 5461 4624
rect 5539 4584 5551 4624
rect 5569 4584 5581 4624
rect 5694 4584 5706 4642
rect 5730 4584 5742 4644
rect 71 4516 83 4556
rect 91 4516 103 4556
rect 111 4528 123 4556
rect 131 4516 143 4556
rect 234 4498 246 4556
rect 270 4496 282 4556
rect 340 4516 352 4556
rect 368 4516 380 4556
rect 390 4536 402 4556
rect 511 4516 523 4556
rect 531 4516 543 4556
rect 551 4528 563 4556
rect 571 4516 583 4556
rect 651 4516 663 4556
rect 671 4516 683 4556
rect 691 4528 703 4556
rect 711 4516 723 4556
rect 777 4536 789 4556
rect 797 4536 809 4556
rect 880 4516 892 4556
rect 908 4516 920 4556
rect 930 4536 942 4556
rect 1031 4536 1043 4556
rect 1051 4536 1063 4556
rect 1154 4498 1166 4556
rect 1190 4496 1202 4556
rect 1278 4536 1290 4556
rect 1300 4516 1312 4556
rect 1328 4516 1340 4556
rect 1411 4536 1423 4556
rect 1431 4536 1443 4556
rect 1497 4516 1509 4556
rect 1517 4528 1529 4556
rect 1537 4516 1549 4556
rect 1557 4516 1569 4556
rect 1659 4516 1671 4556
rect 1689 4516 1701 4556
rect 1794 4498 1806 4556
rect 1830 4496 1842 4556
rect 1911 4536 1923 4556
rect 1931 4536 1943 4556
rect 1951 4536 1963 4556
rect 2054 4498 2066 4556
rect 2090 4496 2102 4556
rect 2214 4498 2226 4556
rect 2250 4496 2262 4556
rect 2339 4516 2351 4556
rect 2369 4516 2381 4556
rect 2474 4498 2486 4556
rect 2510 4496 2522 4556
rect 2578 4496 2590 4556
rect 2614 4498 2626 4556
rect 2731 4536 2743 4556
rect 2751 4536 2763 4556
rect 2831 4536 2843 4556
rect 2851 4536 2863 4556
rect 2871 4536 2883 4556
rect 2974 4498 2986 4556
rect 3010 4496 3022 4556
rect 3114 4498 3126 4556
rect 3150 4496 3162 4556
rect 3217 4536 3229 4556
rect 3237 4536 3249 4556
rect 3317 4516 3329 4556
rect 3337 4528 3349 4556
rect 3357 4516 3369 4556
rect 3377 4516 3389 4556
rect 3481 4516 3493 4556
rect 3501 4516 3513 4556
rect 3531 4516 3543 4556
rect 3619 4516 3631 4556
rect 3649 4516 3661 4556
rect 3751 4516 3763 4556
rect 3771 4536 3783 4556
rect 3791 4536 3803 4556
rect 3811 4536 3823 4556
rect 3879 4516 3891 4556
rect 3909 4516 3921 4556
rect 4009 4516 4021 4556
rect 4029 4516 4041 4556
rect 4051 4536 4063 4556
rect 4117 4516 4129 4556
rect 4147 4516 4159 4556
rect 4167 4516 4179 4556
rect 4279 4516 4291 4556
rect 4309 4516 4321 4556
rect 4391 4516 4403 4556
rect 4411 4516 4423 4556
rect 4431 4528 4443 4556
rect 4451 4516 4463 4556
rect 4519 4516 4531 4556
rect 4549 4516 4561 4556
rect 4659 4516 4671 4556
rect 4689 4516 4701 4556
rect 4757 4536 4769 4556
rect 4777 4536 4789 4556
rect 4859 4516 4871 4556
rect 4889 4516 4901 4556
rect 4977 4516 4989 4556
rect 4997 4528 5009 4556
rect 5017 4516 5029 4556
rect 5037 4516 5049 4556
rect 5077 4516 5089 4556
rect 5099 4536 5111 4556
rect 5129 4536 5141 4556
rect 5157 4536 5169 4556
rect 5183 4536 5195 4556
rect 5205 4536 5217 4556
rect 5235 4536 5247 4556
rect 5267 4536 5279 4556
rect 5287 4516 5299 4556
rect 5357 4516 5369 4556
rect 5377 4528 5389 4556
rect 5397 4516 5409 4556
rect 5417 4516 5429 4556
rect 5497 4536 5509 4556
rect 5517 4536 5529 4556
rect 5537 4536 5549 4556
rect 5557 4516 5569 4556
rect 5651 4516 5663 4556
rect 5671 4516 5683 4556
rect 5691 4528 5703 4556
rect 5711 4516 5723 4556
rect 91 4104 103 4144
rect 111 4104 123 4144
rect 131 4104 143 4132
rect 151 4104 163 4144
rect 231 4104 243 4144
rect 251 4104 263 4144
rect 271 4104 283 4132
rect 291 4104 303 4144
rect 414 4104 426 4162
rect 450 4104 462 4164
rect 554 4104 566 4162
rect 590 4104 602 4164
rect 671 4104 683 4144
rect 691 4104 703 4124
rect 711 4104 723 4124
rect 731 4104 743 4124
rect 811 4104 823 4144
rect 831 4104 843 4144
rect 851 4104 863 4132
rect 871 4104 883 4144
rect 937 4104 949 4124
rect 957 4104 969 4124
rect 1058 4104 1070 4124
rect 1080 4104 1092 4144
rect 1108 4104 1120 4144
rect 1234 4104 1246 4162
rect 1270 4104 1282 4164
rect 1359 4104 1371 4144
rect 1389 4104 1401 4144
rect 1479 4104 1491 4144
rect 1509 4104 1521 4144
rect 1591 4104 1603 4124
rect 1611 4104 1623 4124
rect 1631 4104 1643 4124
rect 1734 4104 1746 4162
rect 1770 4104 1782 4164
rect 1874 4104 1886 4162
rect 1910 4104 1922 4164
rect 1978 4104 1990 4164
rect 2014 4104 2026 4162
rect 2118 4104 2130 4164
rect 2154 4104 2166 4162
rect 2271 4104 2283 4124
rect 2291 4104 2303 4124
rect 2311 4104 2323 4124
rect 2411 4104 2423 4144
rect 2431 4104 2443 4144
rect 2451 4104 2463 4132
rect 2471 4104 2483 4144
rect 2594 4104 2606 4162
rect 2630 4104 2642 4164
rect 2697 4104 2709 4124
rect 2717 4104 2729 4124
rect 2818 4104 2830 4164
rect 2854 4104 2866 4162
rect 2959 4104 2971 4144
rect 2989 4104 3001 4144
rect 3080 4104 3092 4144
rect 3108 4104 3120 4144
rect 3130 4104 3142 4124
rect 3220 4104 3232 4144
rect 3248 4104 3260 4144
rect 3270 4104 3282 4124
rect 3357 4104 3369 4144
rect 3377 4104 3389 4132
rect 3397 4104 3409 4144
rect 3417 4104 3429 4144
rect 3517 4104 3529 4124
rect 3537 4104 3549 4124
rect 3618 4104 3630 4164
rect 3654 4104 3666 4162
rect 3758 4104 3770 4164
rect 3794 4104 3806 4162
rect 3919 4104 3931 4144
rect 3949 4104 3961 4144
rect 4059 4104 4071 4144
rect 4089 4104 4101 4144
rect 4179 4104 4191 4144
rect 4209 4104 4221 4144
rect 4291 4104 4303 4144
rect 4311 4104 4323 4144
rect 4331 4104 4343 4132
rect 4351 4104 4363 4144
rect 4417 4104 4429 4124
rect 4437 4104 4449 4124
rect 4457 4104 4469 4124
rect 4477 4104 4489 4144
rect 4571 4104 4583 4144
rect 4591 4104 4603 4144
rect 4611 4104 4623 4132
rect 4631 4104 4643 4144
rect 4717 4104 4729 4144
rect 4737 4104 4749 4132
rect 4757 4104 4769 4144
rect 4777 4104 4789 4144
rect 4857 4104 4869 4124
rect 4877 4104 4889 4124
rect 4897 4104 4909 4124
rect 4977 4104 4989 4124
rect 4997 4104 5009 4124
rect 5100 4104 5112 4144
rect 5128 4104 5140 4144
rect 5150 4104 5162 4124
rect 5237 4104 5249 4144
rect 5257 4104 5269 4132
rect 5277 4104 5289 4144
rect 5297 4104 5309 4144
rect 5377 4104 5389 4124
rect 5397 4104 5409 4124
rect 5477 4104 5489 4144
rect 5497 4104 5509 4132
rect 5517 4104 5529 4144
rect 5537 4104 5549 4144
rect 5581 4104 5593 4144
rect 5601 4104 5613 4124
rect 5633 4104 5645 4124
rect 5663 4104 5675 4124
rect 5685 4104 5697 4124
rect 5711 4104 5723 4124
rect 5739 4104 5751 4124
rect 5769 4104 5781 4124
rect 5791 4104 5803 4144
rect 71 4056 83 4076
rect 91 4056 103 4076
rect 177 4036 189 4076
rect 197 4048 209 4076
rect 217 4036 229 4076
rect 237 4036 249 4076
rect 331 4056 343 4076
rect 351 4056 363 4076
rect 440 4036 452 4076
rect 468 4036 480 4076
rect 490 4056 502 4076
rect 591 4056 603 4076
rect 611 4056 623 4076
rect 631 4056 643 4076
rect 731 4056 743 4076
rect 751 4056 763 4076
rect 817 4036 829 4076
rect 837 4048 849 4076
rect 857 4036 869 4076
rect 877 4036 889 4076
rect 957 4056 969 4076
rect 977 4056 989 4076
rect 1058 4016 1070 4076
rect 1094 4018 1106 4076
rect 1200 4036 1212 4076
rect 1228 4036 1240 4076
rect 1256 4036 1268 4076
rect 1379 4036 1391 4076
rect 1409 4036 1421 4076
rect 1511 4056 1523 4076
rect 1531 4056 1543 4076
rect 1611 4056 1623 4076
rect 1631 4056 1643 4076
rect 1651 4056 1663 4076
rect 1731 4056 1743 4076
rect 1751 4056 1763 4076
rect 1818 4016 1830 4076
rect 1854 4018 1866 4076
rect 1971 4036 1983 4076
rect 1991 4036 2003 4076
rect 2011 4048 2023 4076
rect 2031 4036 2043 4076
rect 2154 4018 2166 4076
rect 2190 4016 2202 4076
rect 2258 4016 2270 4076
rect 2294 4018 2306 4076
rect 2411 4036 2423 4076
rect 2431 4036 2443 4076
rect 2451 4048 2463 4076
rect 2471 4036 2483 4076
rect 2559 4036 2571 4076
rect 2589 4036 2601 4076
rect 2659 4036 2671 4076
rect 2689 4036 2701 4076
rect 2778 4016 2790 4076
rect 2814 4018 2826 4076
rect 2918 4016 2930 4076
rect 2954 4018 2966 4076
rect 3071 4056 3083 4076
rect 3091 4056 3103 4076
rect 3194 4018 3206 4076
rect 3230 4016 3242 4076
rect 3311 4056 3323 4076
rect 3331 4056 3343 4076
rect 3411 4036 3423 4076
rect 3431 4036 3443 4076
rect 3451 4048 3463 4076
rect 3471 4036 3483 4076
rect 3539 4036 3551 4076
rect 3569 4036 3581 4076
rect 3671 4036 3683 4076
rect 3691 4056 3703 4076
rect 3711 4056 3723 4076
rect 3731 4056 3743 4076
rect 3819 4036 3831 4076
rect 3849 4036 3861 4076
rect 3951 4036 3963 4076
rect 3971 4036 3983 4076
rect 3991 4048 4003 4076
rect 4011 4036 4023 4076
rect 4098 4056 4110 4076
rect 4120 4036 4132 4076
rect 4148 4036 4160 4076
rect 4219 4036 4231 4076
rect 4249 4036 4261 4076
rect 4337 4036 4349 4076
rect 4357 4048 4369 4076
rect 4377 4036 4389 4076
rect 4397 4036 4409 4076
rect 4477 4036 4489 4076
rect 4497 4048 4509 4076
rect 4517 4036 4529 4076
rect 4537 4036 4549 4076
rect 4617 4056 4629 4076
rect 4637 4056 4649 4076
rect 4657 4056 4669 4076
rect 4677 4036 4689 4076
rect 4779 4036 4791 4076
rect 4809 4036 4821 4076
rect 4878 4016 4890 4076
rect 4914 4018 4926 4076
rect 5017 4056 5029 4076
rect 5037 4056 5049 4076
rect 5131 4056 5143 4076
rect 5151 4056 5163 4076
rect 5177 4036 5189 4076
rect 5199 4056 5211 4076
rect 5229 4056 5241 4076
rect 5257 4056 5269 4076
rect 5283 4056 5295 4076
rect 5305 4056 5317 4076
rect 5335 4056 5347 4076
rect 5367 4056 5379 4076
rect 5387 4036 5399 4076
rect 5417 4036 5429 4076
rect 5439 4056 5451 4076
rect 5469 4056 5481 4076
rect 5497 4056 5509 4076
rect 5523 4056 5535 4076
rect 5545 4056 5557 4076
rect 5575 4056 5587 4076
rect 5607 4056 5619 4076
rect 5627 4036 5639 4076
rect 5697 4036 5709 4076
rect 5717 4048 5729 4076
rect 5737 4036 5749 4076
rect 5757 4036 5769 4076
rect 79 3624 91 3664
rect 109 3624 121 3664
rect 214 3624 226 3682
rect 250 3624 262 3684
rect 391 3624 403 3644
rect 411 3624 423 3644
rect 431 3624 443 3644
rect 451 3624 465 3644
rect 551 3624 563 3664
rect 571 3624 583 3664
rect 591 3624 603 3652
rect 611 3624 623 3664
rect 699 3624 711 3664
rect 729 3624 741 3664
rect 797 3624 809 3664
rect 817 3624 829 3652
rect 837 3624 849 3664
rect 857 3624 869 3664
rect 992 3624 1004 3664
rect 1020 3624 1032 3664
rect 1048 3624 1060 3664
rect 1119 3624 1131 3664
rect 1149 3624 1161 3664
rect 1238 3624 1250 3684
rect 1274 3624 1286 3682
rect 1380 3624 1392 3664
rect 1408 3624 1420 3664
rect 1430 3624 1442 3644
rect 1517 3624 1529 3664
rect 1537 3624 1549 3652
rect 1557 3624 1569 3664
rect 1577 3624 1589 3664
rect 1657 3624 1669 3644
rect 1677 3624 1689 3644
rect 1779 3624 1791 3664
rect 1809 3624 1821 3664
rect 1879 3624 1891 3664
rect 1909 3624 1921 3664
rect 1997 3624 2009 3644
rect 2017 3624 2029 3644
rect 2037 3624 2049 3644
rect 2057 3624 2069 3664
rect 2139 3624 2151 3664
rect 2169 3624 2181 3664
rect 2258 3624 2270 3684
rect 2294 3624 2306 3682
rect 2411 3624 2423 3664
rect 2431 3624 2443 3664
rect 2451 3624 2463 3652
rect 2471 3624 2483 3664
rect 2539 3624 2551 3664
rect 2569 3624 2581 3664
rect 2657 3624 2669 3664
rect 2677 3624 2689 3652
rect 2697 3624 2709 3664
rect 2717 3624 2729 3664
rect 2811 3624 2823 3644
rect 2831 3624 2843 3644
rect 2911 3624 2923 3664
rect 2931 3624 2943 3664
rect 2951 3624 2963 3652
rect 2971 3624 2983 3664
rect 3039 3624 3051 3664
rect 3069 3624 3081 3664
rect 3199 3624 3211 3664
rect 3229 3624 3241 3664
rect 3311 3624 3323 3644
rect 3331 3624 3343 3644
rect 3398 3624 3410 3684
rect 3434 3624 3446 3682
rect 3537 3624 3549 3644
rect 3557 3624 3569 3644
rect 3651 3624 3663 3644
rect 3671 3624 3683 3644
rect 3691 3624 3703 3644
rect 3779 3624 3791 3664
rect 3809 3624 3821 3664
rect 3897 3624 3909 3644
rect 3917 3624 3929 3644
rect 4011 3624 4023 3644
rect 4031 3624 4043 3644
rect 4057 3624 4069 3664
rect 4079 3624 4091 3644
rect 4109 3624 4121 3644
rect 4137 3624 4149 3644
rect 4163 3624 4175 3644
rect 4185 3624 4197 3644
rect 4215 3624 4227 3644
rect 4247 3624 4259 3644
rect 4267 3624 4279 3664
rect 4351 3624 4363 3664
rect 4371 3636 4383 3664
rect 4391 3624 4403 3664
rect 4411 3624 4423 3654
rect 4431 3624 4443 3664
rect 4499 3624 4511 3664
rect 4529 3624 4541 3664
rect 4617 3624 4629 3644
rect 4637 3624 4649 3644
rect 4657 3624 4669 3644
rect 4737 3624 4749 3664
rect 4757 3624 4769 3652
rect 4777 3624 4789 3664
rect 4797 3624 4809 3664
rect 4877 3624 4889 3664
rect 4897 3624 4909 3664
rect 5019 3624 5031 3664
rect 5049 3624 5061 3664
rect 5117 3624 5129 3644
rect 5137 3624 5149 3644
rect 5231 3624 5243 3664
rect 5251 3624 5263 3664
rect 5271 3624 5283 3664
rect 5291 3624 5303 3664
rect 5311 3624 5323 3664
rect 5331 3624 5343 3664
rect 5351 3624 5363 3664
rect 5371 3624 5383 3664
rect 5391 3624 5403 3664
rect 5417 3624 5429 3664
rect 5439 3624 5451 3644
rect 5469 3624 5481 3644
rect 5497 3624 5509 3644
rect 5523 3624 5535 3644
rect 5545 3624 5557 3644
rect 5575 3624 5587 3644
rect 5607 3624 5619 3644
rect 5627 3624 5639 3664
rect 5719 3624 5731 3664
rect 5749 3624 5761 3664
rect 71 3556 83 3596
rect 91 3556 103 3596
rect 111 3568 123 3596
rect 131 3556 143 3596
rect 200 3556 212 3596
rect 228 3556 240 3596
rect 250 3576 262 3596
rect 337 3576 349 3596
rect 357 3576 369 3596
rect 437 3556 449 3596
rect 457 3568 469 3596
rect 477 3556 489 3596
rect 497 3556 509 3596
rect 578 3536 590 3596
rect 614 3538 626 3596
rect 759 3556 771 3596
rect 789 3556 801 3596
rect 879 3556 891 3596
rect 909 3556 921 3596
rect 977 3556 989 3596
rect 997 3568 1009 3596
rect 1017 3556 1029 3596
rect 1037 3556 1049 3596
rect 1154 3538 1166 3596
rect 1190 3536 1202 3596
rect 1259 3556 1271 3596
rect 1289 3556 1301 3596
rect 1414 3538 1426 3596
rect 1450 3536 1462 3596
rect 1517 3556 1529 3596
rect 1537 3568 1549 3596
rect 1557 3556 1569 3596
rect 1577 3556 1589 3596
rect 1678 3576 1690 3596
rect 1700 3556 1712 3596
rect 1728 3556 1740 3596
rect 1834 3538 1846 3596
rect 1870 3536 1882 3596
rect 1940 3556 1952 3596
rect 1968 3556 1980 3596
rect 1990 3576 2002 3596
rect 2091 3556 2103 3596
rect 2111 3556 2123 3596
rect 2131 3568 2143 3596
rect 2151 3556 2163 3596
rect 2237 3556 2249 3596
rect 2257 3568 2269 3596
rect 2277 3556 2289 3596
rect 2297 3556 2309 3596
rect 2398 3576 2410 3596
rect 2420 3556 2432 3596
rect 2448 3556 2460 3596
rect 2541 3556 2553 3596
rect 2561 3556 2573 3596
rect 2591 3556 2603 3596
rect 2659 3556 2671 3596
rect 2689 3556 2701 3596
rect 2791 3556 2803 3596
rect 2811 3556 2823 3596
rect 2831 3568 2843 3596
rect 2851 3556 2863 3596
rect 2949 3556 2961 3596
rect 2969 3556 2981 3596
rect 2991 3576 3003 3596
rect 3079 3556 3091 3596
rect 3109 3556 3121 3596
rect 3178 3536 3190 3596
rect 3214 3538 3226 3596
rect 3354 3538 3366 3596
rect 3390 3536 3402 3596
rect 3471 3556 3483 3596
rect 3491 3556 3503 3596
rect 3511 3568 3523 3596
rect 3531 3556 3543 3596
rect 3611 3556 3623 3596
rect 3631 3556 3643 3596
rect 3651 3568 3663 3596
rect 3671 3556 3683 3596
rect 3761 3556 3773 3596
rect 3781 3556 3793 3596
rect 3811 3556 3823 3596
rect 3877 3576 3889 3596
rect 3897 3576 3909 3596
rect 3917 3576 3929 3596
rect 4031 3556 4043 3596
rect 4051 3556 4063 3596
rect 4071 3568 4083 3596
rect 4091 3556 4103 3596
rect 4157 3576 4169 3596
rect 4177 3576 4189 3596
rect 4257 3556 4269 3596
rect 4277 3568 4289 3596
rect 4297 3556 4309 3596
rect 4317 3556 4329 3596
rect 4419 3556 4431 3596
rect 4449 3556 4461 3596
rect 4519 3556 4531 3596
rect 4549 3556 4561 3596
rect 4597 3556 4609 3596
rect 4619 3576 4631 3596
rect 4649 3576 4661 3596
rect 4677 3576 4689 3596
rect 4703 3576 4715 3596
rect 4725 3576 4737 3596
rect 4755 3576 4767 3596
rect 4787 3576 4799 3596
rect 4807 3556 4819 3596
rect 4899 3556 4911 3596
rect 4929 3556 4941 3596
rect 5011 3556 5023 3596
rect 5031 3556 5043 3596
rect 5051 3568 5063 3596
rect 5071 3556 5083 3596
rect 5159 3556 5171 3596
rect 5189 3556 5201 3596
rect 5241 3556 5253 3596
rect 5261 3576 5273 3596
rect 5293 3576 5305 3596
rect 5323 3576 5335 3596
rect 5345 3576 5357 3596
rect 5371 3576 5383 3596
rect 5399 3576 5411 3596
rect 5429 3576 5441 3596
rect 5451 3556 5463 3596
rect 5539 3556 5551 3596
rect 5569 3556 5581 3596
rect 5637 3556 5649 3596
rect 5657 3568 5669 3596
rect 5677 3556 5689 3596
rect 5697 3556 5709 3596
rect 71 3144 83 3164
rect 91 3144 103 3164
rect 171 3144 183 3184
rect 191 3144 203 3184
rect 211 3144 223 3172
rect 231 3144 243 3184
rect 311 3144 323 3164
rect 331 3144 343 3164
rect 399 3144 411 3184
rect 429 3144 441 3184
rect 520 3144 532 3184
rect 548 3144 560 3184
rect 570 3144 582 3164
rect 657 3144 669 3184
rect 687 3144 699 3184
rect 707 3144 719 3184
rect 839 3144 851 3184
rect 869 3144 881 3184
rect 974 3144 986 3202
rect 1010 3144 1022 3204
rect 1114 3144 1126 3202
rect 1150 3144 1162 3204
rect 1220 3144 1232 3184
rect 1248 3144 1260 3184
rect 1270 3144 1282 3164
rect 1371 3144 1383 3164
rect 1391 3144 1403 3164
rect 1494 3144 1506 3202
rect 1530 3144 1542 3204
rect 1634 3144 1646 3202
rect 1670 3144 1682 3204
rect 1758 3144 1770 3164
rect 1780 3144 1792 3184
rect 1808 3144 1820 3184
rect 1919 3144 1931 3184
rect 1949 3144 1961 3184
rect 2038 3144 2050 3164
rect 2060 3144 2072 3184
rect 2088 3144 2100 3184
rect 2159 3144 2171 3184
rect 2189 3144 2201 3184
rect 2301 3144 2313 3184
rect 2321 3144 2333 3184
rect 2351 3144 2363 3184
rect 2419 3144 2431 3184
rect 2449 3144 2461 3184
rect 2551 3144 2563 3184
rect 2571 3144 2583 3184
rect 2591 3144 2603 3172
rect 2611 3144 2623 3184
rect 2698 3144 2710 3164
rect 2720 3144 2732 3184
rect 2748 3144 2760 3184
rect 2818 3144 2830 3204
rect 2854 3144 2866 3202
rect 2958 3144 2970 3204
rect 2994 3144 3006 3202
rect 3119 3144 3131 3184
rect 3149 3144 3161 3184
rect 3259 3144 3271 3184
rect 3289 3144 3301 3184
rect 3357 3144 3369 3164
rect 3377 3144 3389 3164
rect 3494 3144 3506 3202
rect 3530 3144 3542 3204
rect 3600 3144 3612 3184
rect 3628 3144 3640 3184
rect 3650 3144 3662 3164
rect 3751 3144 3763 3184
rect 3771 3144 3783 3184
rect 3791 3144 3803 3172
rect 3811 3144 3823 3184
rect 3877 3144 3889 3164
rect 3897 3144 3909 3164
rect 3937 3144 3949 3184
rect 3959 3144 3971 3164
rect 3989 3144 4001 3164
rect 4017 3144 4029 3164
rect 4043 3144 4055 3164
rect 4065 3144 4077 3164
rect 4095 3144 4107 3164
rect 4127 3144 4139 3164
rect 4147 3144 4159 3184
rect 4217 3144 4229 3184
rect 4237 3144 4249 3172
rect 4257 3144 4269 3184
rect 4277 3144 4289 3184
rect 4357 3144 4369 3184
rect 4377 3144 4389 3172
rect 4397 3144 4409 3184
rect 4417 3144 4429 3184
rect 4457 3144 4469 3184
rect 4479 3144 4491 3164
rect 4509 3144 4521 3164
rect 4537 3144 4549 3164
rect 4563 3144 4575 3164
rect 4585 3144 4597 3164
rect 4615 3144 4627 3164
rect 4647 3144 4659 3164
rect 4667 3144 4679 3184
rect 4737 3144 4749 3184
rect 4757 3144 4769 3172
rect 4777 3144 4789 3184
rect 4797 3144 4809 3184
rect 4899 3144 4911 3184
rect 4929 3144 4941 3184
rect 5011 3144 5023 3184
rect 5031 3144 5043 3184
rect 5051 3144 5063 3172
rect 5071 3144 5083 3184
rect 5151 3144 5163 3164
rect 5171 3144 5183 3164
rect 5259 3144 5271 3184
rect 5289 3144 5301 3184
rect 5357 3144 5369 3164
rect 5377 3144 5389 3164
rect 5477 3144 5489 3184
rect 5497 3144 5509 3172
rect 5517 3144 5529 3184
rect 5537 3144 5549 3184
rect 5659 3144 5671 3184
rect 5689 3144 5701 3184
rect 101 3076 113 3116
rect 121 3076 133 3116
rect 151 3076 163 3116
rect 238 3056 250 3116
rect 274 3058 286 3116
rect 379 3076 391 3116
rect 409 3076 421 3116
rect 511 3076 523 3116
rect 531 3076 543 3116
rect 551 3088 563 3116
rect 571 3076 583 3116
rect 637 3076 649 3116
rect 657 3088 669 3116
rect 677 3076 689 3116
rect 697 3076 709 3116
rect 777 3076 789 3116
rect 797 3088 809 3116
rect 817 3076 829 3116
rect 837 3076 849 3116
rect 917 3076 929 3116
rect 937 3088 949 3116
rect 957 3076 969 3116
rect 977 3076 989 3116
rect 1079 3076 1091 3116
rect 1109 3076 1121 3116
rect 1211 3096 1223 3116
rect 1231 3096 1243 3116
rect 1251 3096 1263 3116
rect 1317 3076 1329 3116
rect 1337 3088 1349 3116
rect 1357 3076 1369 3116
rect 1377 3076 1389 3116
rect 1494 3058 1506 3116
rect 1530 3056 1542 3116
rect 1638 3096 1650 3116
rect 1660 3076 1672 3116
rect 1688 3076 1700 3116
rect 1771 3076 1783 3116
rect 1791 3076 1803 3116
rect 1811 3088 1823 3116
rect 1831 3076 1843 3116
rect 1897 3076 1909 3116
rect 1917 3088 1929 3116
rect 1937 3076 1949 3116
rect 1957 3076 1969 3116
rect 2071 3076 2083 3116
rect 2091 3076 2103 3116
rect 2111 3088 2123 3116
rect 2131 3076 2143 3116
rect 2211 3076 2223 3116
rect 2231 3076 2243 3116
rect 2251 3088 2263 3116
rect 2271 3076 2283 3116
rect 2378 3096 2390 3116
rect 2400 3076 2412 3116
rect 2428 3076 2440 3116
rect 2518 3096 2530 3116
rect 2540 3076 2552 3116
rect 2568 3076 2580 3116
rect 2672 3076 2684 3116
rect 2700 3076 2712 3116
rect 2728 3076 2740 3116
rect 2811 3076 2823 3116
rect 2831 3096 2843 3116
rect 2851 3096 2863 3116
rect 2871 3096 2883 3116
rect 2937 3096 2949 3116
rect 2957 3096 2969 3116
rect 2977 3096 2989 3116
rect 3079 3076 3091 3116
rect 3109 3076 3121 3116
rect 3221 3076 3233 3116
rect 3241 3076 3253 3116
rect 3271 3076 3283 3116
rect 3337 3096 3349 3116
rect 3357 3096 3369 3116
rect 3377 3096 3389 3116
rect 3397 3076 3409 3116
rect 3491 3076 3503 3116
rect 3511 3076 3523 3116
rect 3531 3088 3543 3116
rect 3551 3076 3563 3116
rect 3631 3076 3643 3116
rect 3651 3076 3663 3116
rect 3671 3088 3683 3116
rect 3691 3076 3703 3116
rect 3771 3076 3783 3116
rect 3791 3096 3803 3116
rect 3811 3096 3823 3116
rect 3831 3096 3843 3116
rect 3941 3076 3953 3116
rect 3961 3076 3973 3116
rect 3991 3076 4003 3116
rect 4057 3096 4069 3116
rect 4077 3096 4089 3116
rect 4097 3096 4109 3116
rect 4178 3056 4190 3116
rect 4214 3058 4226 3116
rect 4281 3076 4293 3116
rect 4301 3096 4313 3116
rect 4333 3096 4345 3116
rect 4363 3096 4375 3116
rect 4385 3096 4397 3116
rect 4411 3096 4423 3116
rect 4439 3096 4451 3116
rect 4469 3096 4481 3116
rect 4491 3076 4503 3116
rect 4577 3076 4589 3116
rect 4597 3088 4609 3116
rect 4617 3076 4629 3116
rect 4637 3076 4649 3116
rect 4717 3076 4729 3116
rect 4737 3088 4749 3116
rect 4757 3076 4769 3116
rect 4777 3076 4789 3116
rect 4879 3076 4891 3116
rect 4909 3076 4921 3116
rect 4979 3076 4991 3116
rect 5009 3076 5021 3116
rect 5061 3076 5073 3116
rect 5081 3096 5093 3116
rect 5113 3096 5125 3116
rect 5143 3096 5155 3116
rect 5165 3096 5177 3116
rect 5191 3096 5203 3116
rect 5219 3096 5231 3116
rect 5249 3096 5261 3116
rect 5271 3076 5283 3116
rect 5351 3076 5363 3116
rect 5371 3076 5383 3116
rect 5391 3076 5403 3116
rect 5411 3076 5423 3116
rect 5431 3076 5443 3116
rect 5451 3076 5463 3116
rect 5471 3076 5483 3116
rect 5491 3076 5503 3116
rect 5511 3076 5523 3116
rect 5537 3076 5549 3116
rect 5559 3096 5571 3116
rect 5589 3096 5601 3116
rect 5617 3096 5629 3116
rect 5643 3096 5655 3116
rect 5665 3096 5677 3116
rect 5695 3096 5707 3116
rect 5727 3096 5739 3116
rect 5747 3076 5759 3116
rect 79 2664 91 2704
rect 109 2664 121 2704
rect 177 2664 189 2704
rect 197 2664 209 2692
rect 217 2664 229 2704
rect 237 2664 249 2704
rect 331 2664 343 2684
rect 351 2664 363 2684
rect 420 2664 432 2704
rect 448 2664 460 2704
rect 470 2664 482 2684
rect 579 2664 591 2704
rect 609 2664 621 2704
rect 677 2664 689 2704
rect 707 2664 719 2704
rect 727 2664 739 2704
rect 819 2664 831 2704
rect 849 2664 861 2704
rect 940 2664 952 2704
rect 968 2664 980 2704
rect 990 2664 1002 2684
rect 1079 2664 1091 2704
rect 1109 2664 1121 2704
rect 1231 2664 1243 2704
rect 1251 2664 1263 2704
rect 1271 2664 1283 2692
rect 1291 2664 1303 2704
rect 1357 2664 1369 2704
rect 1377 2664 1389 2692
rect 1397 2664 1409 2704
rect 1417 2664 1429 2704
rect 1511 2664 1523 2704
rect 1531 2664 1543 2684
rect 1551 2664 1563 2684
rect 1571 2664 1583 2684
rect 1637 2664 1649 2684
rect 1657 2664 1669 2684
rect 1677 2664 1689 2684
rect 1781 2664 1793 2704
rect 1801 2664 1813 2704
rect 1831 2664 1843 2704
rect 1939 2664 1951 2704
rect 1969 2664 1981 2704
rect 2037 2664 2049 2704
rect 2057 2664 2069 2692
rect 2077 2664 2089 2704
rect 2097 2664 2109 2704
rect 2201 2664 2213 2704
rect 2221 2664 2233 2704
rect 2251 2664 2263 2704
rect 2339 2664 2351 2704
rect 2369 2664 2381 2704
rect 2457 2664 2469 2684
rect 2477 2664 2489 2684
rect 2497 2664 2509 2684
rect 2614 2664 2626 2722
rect 2650 2664 2662 2724
rect 2741 2664 2753 2704
rect 2761 2664 2773 2704
rect 2791 2664 2803 2704
rect 2877 2664 2889 2704
rect 2897 2664 2909 2692
rect 2917 2664 2929 2704
rect 2937 2664 2949 2704
rect 3054 2664 3066 2722
rect 3090 2664 3102 2724
rect 3159 2664 3171 2704
rect 3189 2664 3201 2704
rect 3291 2664 3303 2704
rect 3311 2664 3323 2704
rect 3331 2664 3343 2692
rect 3351 2664 3363 2704
rect 3441 2664 3453 2704
rect 3461 2664 3473 2704
rect 3491 2664 3503 2704
rect 3557 2664 3569 2684
rect 3577 2664 3589 2684
rect 3597 2664 3609 2684
rect 3678 2664 3690 2724
rect 3714 2664 3726 2722
rect 3819 2664 3831 2704
rect 3849 2664 3861 2704
rect 3951 2664 3963 2704
rect 3971 2664 3983 2704
rect 4051 2664 4063 2704
rect 4071 2664 4083 2704
rect 4091 2664 4103 2692
rect 4111 2664 4123 2704
rect 4179 2664 4191 2704
rect 4209 2664 4221 2704
rect 4297 2664 4309 2704
rect 4317 2664 4329 2704
rect 4397 2664 4409 2684
rect 4417 2664 4429 2684
rect 4457 2664 4469 2704
rect 4479 2664 4491 2684
rect 4509 2664 4521 2684
rect 4537 2664 4549 2684
rect 4563 2664 4575 2684
rect 4585 2664 4597 2684
rect 4615 2664 4627 2684
rect 4647 2664 4659 2684
rect 4667 2664 4679 2704
rect 4701 2664 4713 2704
rect 4721 2664 4733 2684
rect 4753 2664 4765 2684
rect 4783 2664 4795 2684
rect 4805 2664 4817 2684
rect 4831 2664 4843 2684
rect 4859 2664 4871 2684
rect 4889 2664 4901 2684
rect 4911 2664 4923 2704
rect 4997 2664 5009 2704
rect 5017 2664 5029 2692
rect 5037 2664 5049 2704
rect 5057 2664 5069 2704
rect 5139 2664 5151 2704
rect 5169 2664 5181 2704
rect 5257 2664 5269 2704
rect 5277 2664 5289 2704
rect 5297 2664 5309 2704
rect 5337 2664 5349 2704
rect 5359 2664 5371 2684
rect 5389 2664 5401 2684
rect 5417 2664 5429 2684
rect 5443 2664 5455 2684
rect 5465 2664 5477 2684
rect 5495 2664 5507 2684
rect 5527 2664 5539 2684
rect 5547 2664 5559 2704
rect 5617 2664 5629 2704
rect 5637 2664 5649 2692
rect 5657 2664 5669 2704
rect 5677 2664 5689 2704
rect 71 2616 83 2636
rect 91 2616 103 2636
rect 157 2616 169 2636
rect 177 2616 189 2636
rect 278 2616 290 2636
rect 300 2596 312 2636
rect 328 2596 340 2636
rect 398 2576 410 2636
rect 434 2578 446 2636
rect 537 2616 549 2636
rect 557 2616 569 2636
rect 637 2616 649 2636
rect 657 2616 669 2636
rect 677 2616 689 2636
rect 757 2596 769 2636
rect 777 2608 789 2636
rect 797 2596 809 2636
rect 817 2596 829 2636
rect 920 2596 932 2636
rect 948 2596 960 2636
rect 970 2616 982 2636
rect 1071 2596 1083 2636
rect 1091 2596 1103 2636
rect 1111 2608 1123 2636
rect 1131 2596 1143 2636
rect 1219 2596 1231 2636
rect 1249 2596 1261 2636
rect 1317 2596 1329 2636
rect 1347 2596 1359 2636
rect 1367 2596 1379 2636
rect 1494 2578 1506 2636
rect 1530 2576 1542 2636
rect 1597 2616 1609 2636
rect 1617 2616 1629 2636
rect 1697 2596 1709 2636
rect 1717 2608 1729 2636
rect 1737 2596 1749 2636
rect 1757 2596 1769 2636
rect 1851 2596 1863 2636
rect 1871 2596 1883 2636
rect 1891 2608 1903 2636
rect 1911 2596 1923 2636
rect 1977 2596 1989 2636
rect 1997 2608 2009 2636
rect 2017 2596 2029 2636
rect 2037 2596 2049 2636
rect 2154 2578 2166 2636
rect 2190 2576 2202 2636
rect 2278 2616 2290 2636
rect 2300 2596 2312 2636
rect 2328 2596 2340 2636
rect 2399 2596 2411 2636
rect 2429 2596 2441 2636
rect 2551 2596 2563 2636
rect 2571 2596 2583 2636
rect 2591 2608 2603 2636
rect 2611 2596 2623 2636
rect 2677 2596 2689 2636
rect 2697 2608 2709 2636
rect 2717 2596 2729 2636
rect 2737 2596 2749 2636
rect 2838 2616 2850 2636
rect 2860 2596 2872 2636
rect 2888 2596 2900 2636
rect 2971 2616 2983 2636
rect 2991 2616 3003 2636
rect 3057 2596 3069 2636
rect 3077 2608 3089 2636
rect 3097 2596 3109 2636
rect 3117 2596 3129 2636
rect 3219 2596 3231 2636
rect 3249 2596 3261 2636
rect 3374 2578 3386 2636
rect 3410 2576 3422 2636
rect 3477 2596 3489 2636
rect 3507 2596 3519 2636
rect 3527 2596 3539 2636
rect 3619 2596 3631 2636
rect 3649 2596 3661 2636
rect 3740 2596 3752 2636
rect 3768 2596 3780 2636
rect 3796 2596 3808 2636
rect 3897 2616 3909 2636
rect 3917 2616 3929 2636
rect 3937 2616 3949 2636
rect 3985 2616 3997 2636
rect 4005 2616 4017 2636
rect 4031 2596 4043 2636
rect 4067 2596 4079 2636
rect 4104 2596 4116 2636
rect 4135 2616 4147 2636
rect 4155 2616 4167 2636
rect 4175 2616 4187 2636
rect 4200 2616 4212 2636
rect 4220 2616 4232 2636
rect 4240 2616 4252 2636
rect 4270 2616 4282 2636
rect 4290 2616 4302 2636
rect 4310 2616 4322 2636
rect 4330 2616 4342 2636
rect 4358 2596 4370 2636
rect 4394 2596 4406 2636
rect 4430 2596 4442 2636
rect 4458 2596 4470 2636
rect 4494 2596 4506 2636
rect 4530 2596 4542 2636
rect 4558 2616 4570 2636
rect 4578 2616 4590 2636
rect 4598 2616 4610 2636
rect 4618 2616 4630 2636
rect 4648 2616 4660 2636
rect 4668 2616 4680 2636
rect 4688 2616 4700 2636
rect 4713 2616 4725 2636
rect 4733 2616 4745 2636
rect 4753 2616 4765 2636
rect 4784 2596 4796 2636
rect 4821 2596 4833 2636
rect 4857 2596 4869 2636
rect 4883 2616 4895 2636
rect 4903 2616 4915 2636
rect 4941 2596 4953 2636
rect 4961 2616 4973 2636
rect 4993 2616 5005 2636
rect 5023 2616 5035 2636
rect 5045 2616 5057 2636
rect 5071 2616 5083 2636
rect 5099 2616 5111 2636
rect 5129 2616 5141 2636
rect 5151 2596 5163 2636
rect 5231 2596 5243 2636
rect 5251 2596 5263 2636
rect 5271 2596 5283 2636
rect 5291 2596 5303 2636
rect 5311 2596 5323 2636
rect 5331 2596 5343 2636
rect 5351 2596 5363 2636
rect 5371 2596 5383 2636
rect 5391 2596 5403 2636
rect 5477 2596 5489 2636
rect 5497 2596 5509 2636
rect 5517 2596 5529 2636
rect 5537 2596 5549 2636
rect 5557 2596 5569 2636
rect 5577 2596 5589 2636
rect 5597 2596 5609 2636
rect 5617 2596 5629 2636
rect 5637 2596 5649 2636
rect 5717 2596 5729 2636
rect 5737 2596 5749 2636
rect 69 2184 81 2224
rect 89 2184 101 2224
rect 111 2184 123 2204
rect 214 2184 226 2242
rect 250 2184 262 2244
rect 319 2184 331 2224
rect 349 2184 361 2224
rect 437 2184 449 2224
rect 457 2184 469 2212
rect 477 2184 489 2224
rect 497 2184 509 2224
rect 591 2184 603 2224
rect 611 2184 623 2224
rect 631 2184 643 2212
rect 651 2184 663 2224
rect 774 2184 786 2242
rect 810 2184 822 2244
rect 899 2184 911 2224
rect 929 2184 941 2224
rect 1011 2184 1023 2224
rect 1031 2184 1043 2204
rect 1051 2184 1063 2204
rect 1071 2184 1083 2204
rect 1137 2184 1149 2224
rect 1157 2184 1169 2224
rect 1274 2184 1286 2242
rect 1310 2184 1322 2244
rect 1398 2184 1410 2204
rect 1420 2184 1432 2224
rect 1448 2184 1460 2224
rect 1551 2184 1563 2224
rect 1571 2184 1583 2224
rect 1591 2184 1603 2212
rect 1611 2184 1623 2224
rect 1698 2184 1710 2204
rect 1720 2184 1732 2224
rect 1748 2184 1760 2224
rect 1854 2184 1866 2242
rect 1890 2184 1902 2244
rect 1994 2184 2006 2242
rect 2030 2184 2042 2244
rect 2065 2184 2077 2204
rect 2085 2184 2097 2204
rect 2111 2184 2123 2224
rect 2147 2184 2159 2224
rect 2184 2184 2196 2224
rect 2215 2184 2227 2204
rect 2235 2184 2247 2204
rect 2255 2184 2267 2204
rect 2280 2184 2292 2204
rect 2300 2184 2312 2204
rect 2320 2184 2332 2204
rect 2350 2184 2362 2204
rect 2370 2184 2382 2204
rect 2390 2184 2402 2204
rect 2410 2184 2422 2204
rect 2438 2184 2450 2224
rect 2474 2184 2486 2224
rect 2510 2184 2522 2224
rect 2589 2184 2601 2224
rect 2609 2184 2621 2224
rect 2631 2184 2643 2204
rect 2717 2184 2729 2224
rect 2737 2184 2749 2212
rect 2757 2184 2769 2224
rect 2777 2184 2789 2224
rect 2857 2184 2869 2224
rect 2877 2184 2889 2212
rect 2897 2184 2909 2224
rect 2917 2184 2929 2224
rect 3019 2184 3031 2224
rect 3049 2184 3061 2224
rect 3139 2184 3151 2224
rect 3169 2184 3181 2224
rect 3278 2184 3290 2204
rect 3300 2184 3312 2224
rect 3328 2184 3340 2224
rect 3397 2184 3409 2204
rect 3417 2184 3429 2204
rect 3437 2184 3449 2204
rect 3537 2184 3549 2224
rect 3557 2184 3569 2212
rect 3577 2184 3589 2224
rect 3597 2184 3609 2224
rect 3679 2184 3691 2224
rect 3709 2184 3721 2224
rect 3797 2184 3809 2204
rect 3819 2184 3831 2224
rect 3839 2184 3851 2224
rect 3885 2184 3897 2204
rect 3905 2184 3917 2204
rect 3931 2184 3943 2224
rect 3967 2184 3979 2224
rect 4004 2184 4016 2224
rect 4035 2184 4047 2204
rect 4055 2184 4067 2204
rect 4075 2184 4087 2204
rect 4100 2184 4112 2204
rect 4120 2184 4132 2204
rect 4140 2184 4152 2204
rect 4170 2184 4182 2204
rect 4190 2184 4202 2204
rect 4210 2184 4222 2204
rect 4230 2184 4242 2204
rect 4258 2184 4270 2224
rect 4294 2184 4306 2224
rect 4330 2184 4342 2224
rect 4397 2184 4409 2224
rect 4427 2184 4439 2224
rect 4447 2184 4459 2224
rect 4540 2184 4552 2224
rect 4568 2184 4580 2224
rect 4596 2184 4608 2224
rect 4699 2184 4711 2224
rect 4729 2184 4741 2224
rect 4829 2184 4841 2224
rect 4849 2184 4861 2224
rect 4871 2184 4883 2204
rect 4937 2184 4949 2204
rect 4957 2184 4969 2204
rect 5040 2184 5052 2224
rect 5068 2184 5080 2224
rect 5096 2184 5108 2224
rect 5199 2184 5211 2224
rect 5229 2184 5241 2224
rect 5317 2184 5329 2224
rect 5337 2184 5349 2224
rect 5419 2184 5431 2224
rect 5449 2184 5461 2224
rect 5537 2184 5549 2204
rect 5557 2184 5569 2204
rect 5637 2192 5649 2212
rect 5657 2192 5669 2212
rect 5687 2192 5699 2224
rect 5717 2192 5729 2232
rect 89 2116 101 2156
rect 109 2116 121 2156
rect 131 2136 143 2156
rect 254 2098 266 2156
rect 290 2096 302 2156
rect 360 2116 372 2156
rect 388 2116 400 2156
rect 410 2136 422 2156
rect 511 2136 523 2156
rect 531 2136 543 2156
rect 611 2116 623 2156
rect 631 2116 643 2156
rect 651 2128 663 2156
rect 671 2116 683 2156
rect 758 2136 770 2156
rect 780 2116 792 2156
rect 808 2116 820 2156
rect 878 2096 890 2156
rect 914 2098 926 2156
rect 1074 2098 1086 2156
rect 1110 2096 1122 2156
rect 1191 2116 1203 2156
rect 1211 2116 1223 2156
rect 1231 2128 1243 2156
rect 1251 2116 1263 2156
rect 1331 2116 1343 2156
rect 1351 2116 1363 2156
rect 1371 2128 1383 2156
rect 1391 2116 1403 2156
rect 1478 2136 1490 2156
rect 1500 2116 1512 2156
rect 1528 2116 1540 2156
rect 1634 2098 1646 2156
rect 1670 2096 1682 2156
rect 1737 2116 1749 2156
rect 1757 2128 1769 2156
rect 1777 2116 1789 2156
rect 1797 2116 1809 2156
rect 1880 2116 1892 2156
rect 1908 2116 1920 2156
rect 1930 2136 1942 2156
rect 2091 2136 2103 2156
rect 2111 2136 2123 2156
rect 2131 2136 2143 2156
rect 2151 2136 2165 2156
rect 2274 2098 2286 2156
rect 2310 2096 2322 2156
rect 2345 2136 2357 2156
rect 2365 2136 2377 2156
rect 2391 2116 2403 2156
rect 2427 2116 2439 2156
rect 2464 2116 2476 2156
rect 2495 2136 2507 2156
rect 2515 2136 2527 2156
rect 2535 2136 2547 2156
rect 2560 2136 2572 2156
rect 2580 2136 2592 2156
rect 2600 2136 2612 2156
rect 2630 2136 2642 2156
rect 2650 2136 2662 2156
rect 2670 2136 2682 2156
rect 2690 2136 2702 2156
rect 2718 2116 2730 2156
rect 2754 2116 2766 2156
rect 2790 2116 2802 2156
rect 2857 2116 2869 2156
rect 2877 2128 2889 2156
rect 2897 2116 2909 2156
rect 2917 2116 2929 2156
rect 3019 2116 3031 2156
rect 3049 2116 3061 2156
rect 3119 2116 3131 2156
rect 3149 2116 3161 2156
rect 3257 2136 3269 2156
rect 3277 2136 3289 2156
rect 3297 2136 3309 2156
rect 3401 2116 3413 2156
rect 3421 2116 3433 2156
rect 3451 2116 3463 2156
rect 3520 2116 3532 2156
rect 3548 2116 3560 2156
rect 3570 2136 3582 2156
rect 3691 2116 3703 2156
rect 3711 2116 3723 2156
rect 3798 2096 3810 2156
rect 3834 2098 3846 2156
rect 3957 2116 3969 2156
rect 3977 2116 3989 2156
rect 4101 2116 4113 2156
rect 4121 2116 4133 2156
rect 4151 2116 4163 2156
rect 4239 2116 4251 2156
rect 4269 2116 4281 2156
rect 4351 2116 4363 2156
rect 4371 2116 4383 2156
rect 4391 2128 4403 2156
rect 4411 2116 4423 2156
rect 4477 2116 4489 2156
rect 4497 2128 4509 2156
rect 4517 2116 4529 2156
rect 4537 2116 4549 2156
rect 4619 2116 4631 2156
rect 4649 2116 4661 2156
rect 4739 2116 4751 2156
rect 4769 2116 4781 2156
rect 4891 2116 4903 2156
rect 4911 2116 4923 2156
rect 4931 2128 4943 2156
rect 4951 2116 4963 2156
rect 5031 2116 5043 2156
rect 5051 2116 5063 2156
rect 5071 2128 5083 2156
rect 5091 2116 5103 2156
rect 5157 2136 5169 2156
rect 5177 2136 5189 2156
rect 5257 2136 5269 2156
rect 5277 2136 5289 2156
rect 5297 2136 5309 2156
rect 5379 2116 5391 2156
rect 5409 2116 5421 2156
rect 5497 2136 5509 2156
rect 5517 2136 5529 2156
rect 5611 2136 5623 2156
rect 5631 2136 5643 2156
rect 5697 2116 5709 2156
rect 5717 2128 5729 2156
rect 5737 2116 5749 2156
rect 5757 2116 5769 2156
rect 94 1704 106 1762
rect 130 1704 142 1764
rect 200 1704 212 1744
rect 228 1704 240 1744
rect 250 1704 262 1724
rect 351 1704 363 1744
rect 371 1704 383 1744
rect 391 1704 403 1732
rect 411 1704 423 1744
rect 514 1704 526 1762
rect 550 1704 562 1764
rect 651 1704 663 1724
rect 671 1704 683 1724
rect 691 1704 703 1724
rect 760 1704 772 1744
rect 788 1704 800 1744
rect 810 1704 822 1724
rect 931 1704 943 1724
rect 951 1704 963 1724
rect 1051 1704 1063 1744
rect 1071 1704 1083 1744
rect 1091 1704 1103 1732
rect 1111 1704 1123 1744
rect 1191 1704 1203 1744
rect 1211 1704 1223 1744
rect 1231 1704 1243 1732
rect 1251 1704 1263 1744
rect 1331 1704 1343 1724
rect 1351 1704 1363 1724
rect 1431 1704 1443 1744
rect 1451 1704 1463 1744
rect 1471 1704 1483 1732
rect 1491 1704 1503 1744
rect 1557 1704 1569 1744
rect 1577 1704 1589 1732
rect 1597 1704 1609 1744
rect 1617 1704 1629 1744
rect 1711 1704 1723 1744
rect 1731 1704 1743 1744
rect 1751 1704 1763 1732
rect 1771 1704 1783 1744
rect 1859 1704 1871 1744
rect 1889 1704 1901 1744
rect 1979 1704 1991 1744
rect 2009 1704 2021 1744
rect 2111 1704 2123 1744
rect 2131 1704 2143 1744
rect 2151 1704 2163 1744
rect 2185 1704 2197 1724
rect 2205 1704 2217 1724
rect 2231 1704 2243 1744
rect 2267 1704 2279 1744
rect 2304 1704 2316 1744
rect 2335 1704 2347 1724
rect 2355 1704 2367 1724
rect 2375 1704 2387 1724
rect 2400 1704 2412 1724
rect 2420 1704 2432 1724
rect 2440 1704 2452 1724
rect 2470 1704 2482 1724
rect 2490 1704 2502 1724
rect 2510 1704 2522 1724
rect 2530 1704 2542 1724
rect 2558 1704 2570 1744
rect 2594 1704 2606 1744
rect 2630 1704 2642 1744
rect 2699 1704 2711 1744
rect 2729 1704 2741 1744
rect 2854 1704 2866 1762
rect 2890 1704 2902 1764
rect 2971 1704 2983 1744
rect 2991 1704 3003 1744
rect 3011 1704 3023 1732
rect 3031 1704 3043 1744
rect 3097 1704 3109 1724
rect 3117 1704 3129 1724
rect 3137 1704 3149 1724
rect 3217 1712 3229 1732
rect 3237 1712 3249 1732
rect 3267 1712 3279 1744
rect 3297 1712 3309 1752
rect 3391 1704 3403 1724
rect 3411 1704 3423 1724
rect 3477 1704 3489 1744
rect 3497 1704 3509 1734
rect 3517 1704 3529 1744
rect 3537 1716 3549 1744
rect 3557 1704 3569 1744
rect 3651 1704 3663 1744
rect 3671 1704 3683 1744
rect 3691 1704 3703 1732
rect 3711 1704 3723 1744
rect 3811 1704 3823 1744
rect 3831 1704 3843 1744
rect 3851 1704 3863 1732
rect 3871 1704 3883 1744
rect 3937 1704 3949 1744
rect 3957 1704 3969 1732
rect 3977 1704 3989 1744
rect 3997 1704 4009 1744
rect 4099 1704 4111 1744
rect 4129 1704 4141 1744
rect 4232 1704 4244 1744
rect 4260 1704 4272 1744
rect 4288 1704 4300 1744
rect 4379 1704 4391 1744
rect 4409 1704 4421 1744
rect 4477 1704 4489 1744
rect 4497 1704 4509 1732
rect 4517 1704 4529 1744
rect 4537 1704 4549 1744
rect 4641 1704 4653 1744
rect 4661 1704 4673 1744
rect 4691 1704 4703 1744
rect 4771 1704 4783 1724
rect 4791 1704 4803 1724
rect 4811 1704 4823 1724
rect 4899 1704 4911 1744
rect 4929 1704 4941 1744
rect 5032 1704 5044 1744
rect 5060 1704 5072 1744
rect 5088 1704 5100 1744
rect 5171 1704 5183 1724
rect 5191 1704 5203 1724
rect 5271 1704 5283 1724
rect 5291 1704 5303 1724
rect 5311 1704 5323 1724
rect 5377 1704 5389 1744
rect 5397 1704 5409 1732
rect 5417 1704 5429 1744
rect 5437 1704 5449 1744
rect 5531 1704 5543 1744
rect 5551 1704 5563 1744
rect 5571 1704 5583 1732
rect 5591 1704 5603 1744
rect 5657 1704 5669 1744
rect 5677 1704 5689 1744
rect 5697 1704 5709 1744
rect 78 1616 90 1676
rect 114 1618 126 1676
rect 254 1618 266 1676
rect 290 1616 302 1676
rect 360 1636 372 1676
rect 388 1636 400 1676
rect 410 1656 422 1676
rect 518 1656 530 1676
rect 540 1636 552 1676
rect 568 1636 580 1676
rect 639 1636 651 1676
rect 669 1636 681 1676
rect 757 1656 769 1676
rect 777 1656 789 1676
rect 871 1636 883 1676
rect 891 1636 903 1676
rect 911 1648 923 1676
rect 931 1636 943 1676
rect 1034 1618 1046 1676
rect 1070 1616 1082 1676
rect 1159 1636 1171 1676
rect 1189 1636 1201 1676
rect 1277 1656 1289 1676
rect 1297 1656 1309 1676
rect 1317 1656 1329 1676
rect 1409 1636 1421 1676
rect 1429 1636 1441 1676
rect 1451 1656 1463 1676
rect 1551 1656 1563 1676
rect 1571 1656 1583 1676
rect 1640 1636 1652 1676
rect 1668 1636 1680 1676
rect 1696 1636 1708 1676
rect 1765 1656 1777 1676
rect 1785 1656 1797 1676
rect 1811 1636 1823 1676
rect 1847 1636 1859 1676
rect 1884 1636 1896 1676
rect 1915 1656 1927 1676
rect 1935 1656 1947 1676
rect 1955 1656 1967 1676
rect 1980 1656 1992 1676
rect 2000 1656 2012 1676
rect 2020 1656 2032 1676
rect 2050 1656 2062 1676
rect 2070 1656 2082 1676
rect 2090 1656 2102 1676
rect 2110 1656 2122 1676
rect 2138 1636 2150 1676
rect 2174 1636 2186 1676
rect 2210 1636 2222 1676
rect 2297 1636 2309 1676
rect 2317 1648 2329 1676
rect 2337 1636 2349 1676
rect 2357 1636 2369 1676
rect 2439 1636 2451 1676
rect 2469 1636 2481 1676
rect 2571 1636 2583 1676
rect 2591 1636 2603 1676
rect 2611 1648 2623 1676
rect 2631 1636 2643 1676
rect 2719 1636 2731 1676
rect 2749 1636 2761 1676
rect 2831 1636 2843 1676
rect 2851 1636 2863 1676
rect 2871 1648 2883 1676
rect 2891 1636 2903 1676
rect 2971 1636 2983 1676
rect 2991 1636 3003 1676
rect 3011 1648 3023 1676
rect 3031 1636 3043 1676
rect 3058 1636 3070 1676
rect 3094 1636 3106 1676
rect 3130 1636 3142 1676
rect 3158 1656 3170 1676
rect 3178 1656 3190 1676
rect 3198 1656 3210 1676
rect 3218 1656 3230 1676
rect 3248 1656 3260 1676
rect 3268 1656 3280 1676
rect 3288 1656 3300 1676
rect 3313 1656 3325 1676
rect 3333 1656 3345 1676
rect 3353 1656 3365 1676
rect 3384 1636 3396 1676
rect 3421 1636 3433 1676
rect 3457 1636 3469 1676
rect 3483 1656 3495 1676
rect 3503 1656 3515 1676
rect 3598 1656 3610 1676
rect 3620 1636 3632 1676
rect 3648 1636 3660 1676
rect 3717 1636 3729 1676
rect 3737 1648 3749 1676
rect 3757 1636 3769 1676
rect 3777 1636 3789 1676
rect 3869 1636 3881 1676
rect 3889 1636 3901 1676
rect 3911 1656 3923 1676
rect 4001 1636 4013 1676
rect 4021 1636 4033 1676
rect 4051 1636 4063 1676
rect 4119 1636 4131 1676
rect 4149 1636 4161 1676
rect 4272 1636 4284 1676
rect 4300 1636 4312 1676
rect 4328 1636 4340 1676
rect 4432 1636 4444 1676
rect 4460 1636 4472 1676
rect 4488 1636 4500 1676
rect 4580 1636 4592 1676
rect 4608 1636 4620 1676
rect 4636 1636 4648 1676
rect 4739 1636 4751 1676
rect 4769 1636 4781 1676
rect 4857 1636 4869 1676
rect 4877 1648 4889 1676
rect 4897 1636 4909 1676
rect 4917 1636 4929 1676
rect 5021 1636 5033 1676
rect 5041 1636 5053 1676
rect 5071 1636 5083 1676
rect 5158 1616 5170 1676
rect 5194 1618 5206 1676
rect 5300 1636 5312 1676
rect 5328 1636 5340 1676
rect 5356 1636 5368 1676
rect 5459 1636 5471 1676
rect 5489 1636 5501 1676
rect 5578 1616 5590 1676
rect 5614 1618 5626 1676
rect 5751 1636 5763 1676
rect 5771 1636 5783 1676
rect 94 1224 106 1282
rect 130 1224 142 1284
rect 200 1224 212 1264
rect 228 1224 240 1264
rect 250 1224 262 1244
rect 374 1224 386 1282
rect 410 1224 422 1284
rect 491 1224 503 1264
rect 511 1224 523 1264
rect 531 1224 543 1252
rect 551 1224 563 1264
rect 631 1224 643 1264
rect 651 1224 663 1264
rect 671 1224 683 1252
rect 691 1224 703 1264
rect 801 1224 813 1264
rect 821 1224 833 1264
rect 851 1224 863 1264
rect 919 1224 931 1264
rect 949 1224 961 1264
rect 1051 1224 1063 1244
rect 1071 1224 1083 1244
rect 1138 1224 1150 1284
rect 1174 1224 1186 1282
rect 1279 1224 1291 1264
rect 1309 1224 1321 1264
rect 1419 1224 1431 1264
rect 1449 1224 1461 1264
rect 1539 1224 1551 1264
rect 1569 1224 1581 1264
rect 1694 1224 1706 1282
rect 1730 1224 1742 1284
rect 1799 1224 1811 1264
rect 1829 1224 1841 1264
rect 1954 1224 1966 1282
rect 1990 1224 2002 1284
rect 2071 1224 2083 1244
rect 2091 1224 2103 1244
rect 2214 1224 2226 1282
rect 2250 1224 2262 1284
rect 2354 1224 2366 1282
rect 2390 1224 2402 1284
rect 2457 1224 2469 1244
rect 2477 1224 2489 1244
rect 2591 1224 2603 1264
rect 2611 1224 2623 1264
rect 2631 1224 2643 1252
rect 2651 1224 2663 1264
rect 2720 1224 2732 1264
rect 2748 1224 2760 1264
rect 2770 1224 2782 1244
rect 2871 1224 2883 1264
rect 2891 1224 2903 1264
rect 2911 1224 2923 1252
rect 2931 1224 2943 1264
rect 3011 1224 3023 1264
rect 3031 1224 3043 1264
rect 3051 1224 3063 1252
rect 3071 1224 3083 1264
rect 3151 1224 3163 1264
rect 3171 1224 3183 1264
rect 3191 1224 3203 1252
rect 3211 1224 3223 1264
rect 3291 1224 3303 1244
rect 3311 1224 3323 1244
rect 3377 1224 3389 1244
rect 3397 1224 3409 1244
rect 3489 1224 3501 1264
rect 3509 1224 3521 1264
rect 3531 1224 3543 1244
rect 3638 1224 3650 1244
rect 3660 1224 3672 1264
rect 3688 1224 3700 1264
rect 3757 1224 3769 1264
rect 3777 1224 3789 1252
rect 3797 1224 3809 1264
rect 3817 1224 3829 1264
rect 3911 1224 3923 1244
rect 3931 1224 3943 1244
rect 4011 1224 4023 1264
rect 4031 1224 4043 1264
rect 4051 1224 4063 1252
rect 4071 1224 4083 1264
rect 4151 1224 4163 1264
rect 4171 1224 4183 1264
rect 4191 1224 4203 1252
rect 4211 1224 4223 1264
rect 4298 1224 4310 1244
rect 4320 1224 4332 1264
rect 4348 1224 4360 1264
rect 4431 1224 4443 1264
rect 4451 1224 4463 1264
rect 4471 1224 4483 1252
rect 4491 1224 4503 1264
rect 4577 1224 4589 1264
rect 4597 1224 4609 1252
rect 4617 1224 4629 1264
rect 4637 1224 4649 1264
rect 4719 1224 4731 1264
rect 4749 1224 4761 1264
rect 4837 1224 4849 1264
rect 4857 1224 4869 1252
rect 4877 1224 4889 1264
rect 4897 1224 4909 1264
rect 4977 1224 4989 1244
rect 4997 1224 5009 1244
rect 5017 1224 5029 1244
rect 5099 1224 5111 1264
rect 5129 1224 5141 1264
rect 5239 1224 5251 1264
rect 5269 1224 5281 1264
rect 5351 1224 5363 1264
rect 5371 1224 5383 1264
rect 5391 1224 5403 1252
rect 5411 1224 5423 1264
rect 5477 1224 5489 1264
rect 5497 1224 5509 1252
rect 5517 1224 5529 1264
rect 5537 1224 5549 1264
rect 5637 1224 5649 1264
rect 5657 1224 5669 1252
rect 5677 1224 5689 1264
rect 5697 1224 5709 1264
rect 71 1176 83 1196
rect 91 1176 103 1196
rect 160 1156 172 1196
rect 188 1156 200 1196
rect 210 1176 222 1196
rect 297 1156 309 1196
rect 317 1168 329 1196
rect 337 1156 349 1196
rect 357 1156 369 1196
rect 437 1156 449 1196
rect 457 1168 469 1196
rect 477 1156 489 1196
rect 497 1156 509 1196
rect 614 1138 626 1196
rect 650 1136 662 1196
rect 717 1156 729 1196
rect 737 1168 749 1196
rect 757 1156 769 1196
rect 777 1156 789 1196
rect 880 1156 892 1196
rect 908 1156 920 1196
rect 930 1176 942 1196
rect 1031 1156 1043 1196
rect 1051 1156 1063 1196
rect 1071 1168 1083 1196
rect 1091 1156 1103 1196
rect 1171 1176 1183 1196
rect 1191 1176 1203 1196
rect 1260 1156 1272 1196
rect 1288 1156 1300 1196
rect 1310 1176 1322 1196
rect 1411 1176 1423 1196
rect 1431 1176 1443 1196
rect 1511 1176 1523 1196
rect 1531 1176 1543 1196
rect 1551 1176 1563 1196
rect 1637 1176 1649 1196
rect 1657 1176 1669 1196
rect 1774 1138 1786 1196
rect 1810 1136 1822 1196
rect 1899 1156 1911 1196
rect 1929 1156 1941 1196
rect 2011 1156 2023 1196
rect 2031 1156 2043 1196
rect 2051 1168 2063 1196
rect 2071 1156 2083 1196
rect 2174 1138 2186 1196
rect 2210 1136 2222 1196
rect 2314 1138 2326 1196
rect 2350 1136 2362 1196
rect 2431 1156 2443 1196
rect 2451 1156 2463 1196
rect 2471 1168 2483 1196
rect 2491 1156 2503 1196
rect 2594 1138 2606 1196
rect 2630 1136 2642 1196
rect 2717 1176 2729 1196
rect 2737 1176 2749 1196
rect 2817 1176 2829 1196
rect 2837 1176 2849 1196
rect 2857 1176 2869 1196
rect 2937 1176 2949 1196
rect 2957 1176 2969 1196
rect 2977 1176 2989 1196
rect 3057 1156 3069 1196
rect 3087 1156 3099 1196
rect 3107 1156 3119 1196
rect 3211 1176 3223 1196
rect 3231 1176 3243 1196
rect 3251 1176 3263 1196
rect 3351 1176 3363 1196
rect 3371 1176 3383 1196
rect 3391 1176 3403 1196
rect 3471 1176 3483 1196
rect 3491 1176 3503 1196
rect 3571 1156 3583 1196
rect 3591 1156 3603 1196
rect 3611 1168 3623 1196
rect 3631 1156 3643 1196
rect 3711 1156 3723 1196
rect 3731 1156 3743 1196
rect 3751 1168 3763 1196
rect 3771 1156 3783 1196
rect 3839 1156 3851 1196
rect 3869 1156 3881 1196
rect 3959 1156 3971 1196
rect 3989 1156 4001 1196
rect 4077 1176 4089 1196
rect 4097 1176 4109 1196
rect 4117 1176 4129 1196
rect 4197 1176 4209 1196
rect 4217 1176 4229 1196
rect 4318 1176 4330 1196
rect 4340 1156 4352 1196
rect 4368 1156 4380 1196
rect 4471 1156 4483 1196
rect 4491 1156 4503 1196
rect 4511 1168 4523 1196
rect 4531 1156 4543 1196
rect 4618 1176 4630 1196
rect 4640 1156 4652 1196
rect 4668 1156 4680 1196
rect 4737 1156 4749 1196
rect 4757 1168 4769 1196
rect 4777 1156 4789 1196
rect 4797 1156 4809 1196
rect 4877 1176 4889 1196
rect 4899 1156 4911 1196
rect 4919 1156 4931 1196
rect 4997 1176 5009 1196
rect 5017 1176 5029 1196
rect 5097 1176 5109 1196
rect 5117 1176 5129 1196
rect 5219 1156 5231 1196
rect 5249 1156 5261 1196
rect 5351 1156 5363 1196
rect 5371 1156 5383 1196
rect 5391 1168 5403 1196
rect 5411 1156 5423 1196
rect 5477 1176 5489 1196
rect 5497 1176 5509 1196
rect 5517 1176 5529 1196
rect 5634 1138 5646 1196
rect 5670 1136 5682 1196
rect 5751 1176 5763 1196
rect 5771 1176 5783 1196
rect 94 744 106 802
rect 130 744 142 804
rect 200 744 212 784
rect 228 744 240 784
rect 250 744 262 764
rect 374 744 386 802
rect 410 744 422 804
rect 498 744 510 764
rect 520 744 532 784
rect 548 744 560 784
rect 654 744 666 802
rect 690 744 702 804
rect 760 744 772 784
rect 788 744 800 784
rect 810 744 822 764
rect 911 744 923 784
rect 931 744 943 784
rect 951 744 963 772
rect 971 744 983 784
rect 1074 744 1086 802
rect 1110 744 1122 804
rect 1177 744 1189 784
rect 1197 744 1209 772
rect 1217 744 1229 784
rect 1237 744 1249 784
rect 1354 744 1366 802
rect 1390 744 1402 804
rect 1457 744 1469 764
rect 1477 744 1489 764
rect 1559 744 1571 784
rect 1589 744 1601 784
rect 1734 744 1746 802
rect 1770 744 1782 804
rect 1874 744 1886 802
rect 1910 744 1922 804
rect 1978 744 1990 804
rect 2014 744 2026 802
rect 2117 744 2129 784
rect 2137 744 2149 772
rect 2157 744 2169 784
rect 2177 744 2189 784
rect 2257 744 2269 784
rect 2287 744 2299 784
rect 2307 744 2319 784
rect 2397 744 2409 764
rect 2417 744 2429 764
rect 2519 744 2531 784
rect 2549 744 2561 784
rect 2631 744 2643 784
rect 2651 744 2663 764
rect 2671 744 2683 764
rect 2691 744 2703 764
rect 2759 744 2771 784
rect 2789 744 2801 784
rect 2899 744 2911 784
rect 2929 744 2941 784
rect 3017 744 3029 764
rect 3037 744 3049 764
rect 3131 744 3143 764
rect 3151 744 3163 764
rect 3259 744 3271 784
rect 3289 744 3301 784
rect 3391 744 3403 764
rect 3411 744 3423 764
rect 3431 744 3443 764
rect 3511 744 3523 764
rect 3531 744 3543 764
rect 3551 744 3563 764
rect 3638 744 3650 764
rect 3660 744 3672 784
rect 3688 744 3700 784
rect 3771 744 3783 764
rect 3791 744 3803 764
rect 3871 744 3883 784
rect 3891 744 3903 784
rect 3911 744 3923 772
rect 3931 744 3943 784
rect 3999 744 4011 784
rect 4029 744 4041 784
rect 4131 744 4143 784
rect 4151 744 4163 784
rect 4171 744 4183 772
rect 4191 744 4203 784
rect 4271 744 4283 784
rect 4291 744 4303 784
rect 4311 744 4323 772
rect 4331 744 4343 784
rect 4417 744 4429 764
rect 4437 744 4449 764
rect 4531 744 4543 784
rect 4551 744 4563 784
rect 4571 744 4583 772
rect 4591 744 4603 784
rect 4660 744 4672 784
rect 4688 744 4700 784
rect 4710 744 4722 764
rect 4809 744 4821 784
rect 4829 744 4841 784
rect 4851 744 4863 764
rect 4931 744 4943 784
rect 4951 744 4963 784
rect 4971 744 4983 772
rect 4991 744 5003 784
rect 5060 744 5072 784
rect 5088 744 5100 784
rect 5110 744 5122 764
rect 5211 744 5223 784
rect 5231 744 5243 764
rect 5251 744 5263 764
rect 5271 744 5283 764
rect 5371 744 5383 764
rect 5391 744 5403 764
rect 5492 744 5504 784
rect 5520 744 5532 784
rect 5548 744 5560 784
rect 5637 744 5649 784
rect 5657 744 5669 772
rect 5677 744 5689 784
rect 5697 744 5709 784
rect 94 658 106 716
rect 130 656 142 716
rect 238 696 250 716
rect 260 676 272 716
rect 288 676 300 716
rect 394 658 406 716
rect 430 656 442 716
rect 511 676 523 716
rect 531 676 543 716
rect 551 688 563 716
rect 571 676 583 716
rect 640 676 652 716
rect 668 676 680 716
rect 690 696 702 716
rect 779 676 791 716
rect 809 676 821 716
rect 931 676 943 716
rect 951 676 963 716
rect 971 688 983 716
rect 991 676 1003 716
rect 1094 658 1106 716
rect 1130 656 1142 716
rect 1200 676 1212 716
rect 1228 676 1240 716
rect 1250 696 1262 716
rect 1358 696 1370 716
rect 1380 676 1392 716
rect 1408 676 1420 716
rect 1498 656 1510 716
rect 1534 658 1546 716
rect 1651 676 1663 716
rect 1671 676 1683 716
rect 1691 688 1703 716
rect 1711 676 1723 716
rect 1814 658 1826 716
rect 1850 656 1862 716
rect 1920 676 1932 716
rect 1948 676 1960 716
rect 1970 696 1982 716
rect 2071 696 2083 716
rect 2091 696 2103 716
rect 2111 696 2123 716
rect 2191 676 2203 716
rect 2211 696 2223 716
rect 2231 696 2243 716
rect 2251 696 2263 716
rect 2317 676 2329 716
rect 2347 676 2359 716
rect 2367 676 2379 716
rect 2459 676 2471 716
rect 2489 676 2501 716
rect 2599 676 2611 716
rect 2629 676 2641 716
rect 2711 696 2723 716
rect 2731 696 2743 716
rect 2751 696 2763 716
rect 2817 676 2829 716
rect 2837 688 2849 716
rect 2857 676 2869 716
rect 2877 676 2889 716
rect 2979 676 2991 716
rect 3009 676 3021 716
rect 3080 676 3092 716
rect 3108 676 3120 716
rect 3130 696 3142 716
rect 3254 658 3266 716
rect 3290 656 3302 716
rect 3359 676 3371 716
rect 3389 676 3401 716
rect 3491 676 3503 716
rect 3511 676 3523 716
rect 3531 688 3543 716
rect 3551 676 3563 716
rect 3619 676 3631 716
rect 3649 676 3661 716
rect 3751 676 3763 716
rect 3771 676 3783 716
rect 3791 688 3803 716
rect 3811 676 3823 716
rect 3877 676 3889 716
rect 3897 688 3909 716
rect 3917 676 3929 716
rect 3937 676 3949 716
rect 4020 676 4032 716
rect 4048 676 4060 716
rect 4070 696 4082 716
rect 4177 676 4189 716
rect 4197 688 4209 716
rect 4217 676 4229 716
rect 4237 676 4249 716
rect 4331 696 4343 716
rect 4351 696 4363 716
rect 4438 696 4450 716
rect 4460 676 4472 716
rect 4488 676 4500 716
rect 4571 676 4583 716
rect 4591 676 4603 716
rect 4611 688 4623 716
rect 4631 676 4643 716
rect 4711 676 4723 716
rect 4731 676 4743 716
rect 4751 688 4763 716
rect 4771 676 4783 716
rect 4857 676 4869 716
rect 4877 688 4889 716
rect 4897 676 4909 716
rect 4917 676 4929 716
rect 4997 696 5009 716
rect 5017 696 5029 716
rect 5117 696 5129 716
rect 5139 676 5151 716
rect 5159 676 5171 716
rect 5251 676 5263 716
rect 5271 676 5283 716
rect 5291 688 5303 716
rect 5311 676 5323 716
rect 5377 676 5389 716
rect 5397 688 5409 716
rect 5417 676 5429 716
rect 5437 676 5449 716
rect 5531 676 5543 716
rect 5551 676 5563 716
rect 5571 688 5583 716
rect 5591 676 5603 716
rect 5657 696 5669 716
rect 5677 696 5689 716
rect 5697 696 5709 716
rect 94 264 106 322
rect 130 264 142 324
rect 211 264 223 304
rect 231 264 243 304
rect 251 264 263 292
rect 271 264 283 304
rect 371 264 383 304
rect 391 264 403 304
rect 411 264 423 292
rect 431 264 443 304
rect 534 264 546 322
rect 570 264 582 324
rect 661 264 673 304
rect 681 264 693 304
rect 711 264 723 304
rect 814 264 826 322
rect 850 264 862 324
rect 938 264 950 284
rect 960 264 972 304
rect 988 264 1000 304
rect 1058 264 1070 324
rect 1094 264 1106 322
rect 1211 264 1223 304
rect 1231 264 1243 284
rect 1251 264 1263 284
rect 1271 264 1283 284
rect 1374 264 1386 322
rect 1410 264 1422 324
rect 1511 264 1523 284
rect 1531 264 1543 284
rect 1611 264 1623 304
rect 1631 264 1643 304
rect 1651 264 1663 292
rect 1671 264 1683 304
rect 1761 264 1773 304
rect 1781 264 1793 304
rect 1811 264 1823 304
rect 1877 264 1889 284
rect 1897 264 1909 284
rect 1917 264 1929 284
rect 2017 264 2029 284
rect 2037 264 2049 284
rect 2131 264 2143 304
rect 2151 264 2163 304
rect 2171 264 2183 292
rect 2191 264 2203 304
rect 2278 264 2290 284
rect 2300 264 2312 304
rect 2328 264 2340 304
rect 2411 264 2423 284
rect 2431 264 2443 284
rect 2534 264 2546 322
rect 2570 264 2582 324
rect 2637 264 2649 304
rect 2657 264 2669 292
rect 2677 264 2689 304
rect 2697 264 2709 304
rect 2791 264 2803 284
rect 2811 264 2823 284
rect 2891 264 2903 284
rect 2911 264 2923 284
rect 2931 264 2943 284
rect 2997 264 3009 284
rect 3017 264 3029 284
rect 3118 264 3130 284
rect 3140 264 3152 304
rect 3168 264 3180 304
rect 3260 264 3272 304
rect 3288 264 3300 304
rect 3310 264 3322 284
rect 3411 264 3423 284
rect 3431 264 3443 284
rect 3517 264 3529 304
rect 3537 264 3549 292
rect 3557 264 3569 304
rect 3577 264 3589 304
rect 3660 264 3672 304
rect 3688 264 3700 304
rect 3710 264 3722 284
rect 3834 264 3846 322
rect 3870 264 3882 324
rect 3939 264 3951 304
rect 3969 264 3981 304
rect 4114 264 4126 322
rect 4150 264 4162 324
rect 4231 264 4243 304
rect 4251 264 4263 304
rect 4271 264 4283 292
rect 4291 264 4303 304
rect 4371 264 4383 284
rect 4391 264 4403 284
rect 4479 264 4491 304
rect 4509 264 4521 304
rect 4591 264 4603 304
rect 4611 264 4623 304
rect 4631 264 4643 292
rect 4651 264 4663 304
rect 4731 264 4743 284
rect 4751 264 4763 284
rect 4831 264 4843 304
rect 4851 264 4863 304
rect 4871 264 4883 292
rect 4891 264 4903 304
rect 4957 272 4969 292
rect 4977 272 4989 292
rect 5007 272 5019 304
rect 5037 272 5049 312
rect 5131 264 5143 304
rect 5151 264 5163 304
rect 5171 264 5183 292
rect 5191 264 5203 304
rect 5277 264 5289 304
rect 5297 264 5309 292
rect 5317 264 5329 304
rect 5337 264 5349 304
rect 5458 264 5470 284
rect 5480 264 5492 304
rect 5508 264 5520 304
rect 5577 264 5589 304
rect 5597 264 5609 292
rect 5617 264 5629 304
rect 5637 264 5649 304
rect 5719 264 5731 304
rect 5749 264 5761 304
rect 94 178 106 236
rect 130 176 142 236
rect 200 196 212 236
rect 228 196 240 236
rect 250 216 262 236
rect 378 216 390 236
rect 400 196 412 236
rect 428 196 440 236
rect 511 196 523 236
rect 531 196 543 236
rect 551 208 563 236
rect 571 196 583 236
rect 637 196 649 236
rect 657 208 669 236
rect 677 196 689 236
rect 697 196 709 236
rect 814 178 826 236
rect 850 176 862 236
rect 917 216 929 236
rect 937 216 949 236
rect 1017 196 1029 236
rect 1037 208 1049 236
rect 1057 196 1069 236
rect 1077 196 1089 236
rect 1160 196 1172 236
rect 1188 196 1200 236
rect 1210 216 1222 236
rect 1297 216 1309 236
rect 1317 216 1329 236
rect 1337 216 1349 236
rect 1417 196 1429 236
rect 1447 196 1459 236
rect 1467 196 1479 236
rect 1571 216 1583 236
rect 1591 216 1603 236
rect 1671 196 1683 236
rect 1691 196 1703 236
rect 1711 208 1723 236
rect 1731 196 1743 236
rect 1819 196 1831 236
rect 1849 196 1861 236
rect 1918 176 1930 236
rect 1954 178 1966 236
rect 2114 178 2126 236
rect 2150 176 2162 236
rect 2217 216 2229 236
rect 2239 196 2251 236
rect 2259 196 2271 236
rect 2359 196 2371 236
rect 2389 196 2401 236
rect 2457 196 2469 236
rect 2487 196 2499 236
rect 2507 196 2519 236
rect 2618 216 2630 236
rect 2640 196 2652 236
rect 2668 196 2680 236
rect 2761 196 2773 236
rect 2781 196 2793 236
rect 2811 196 2823 236
rect 2899 196 2911 236
rect 2929 196 2941 236
rect 3039 196 3051 236
rect 3069 196 3081 236
rect 3174 178 3186 236
rect 3210 176 3222 236
rect 3291 216 3303 236
rect 3311 216 3323 236
rect 3377 196 3389 236
rect 3397 208 3409 236
rect 3417 196 3429 236
rect 3437 196 3449 236
rect 3531 216 3543 236
rect 3551 216 3563 236
rect 3639 196 3651 236
rect 3669 196 3681 236
rect 3749 196 3761 236
rect 3769 196 3781 236
rect 3791 216 3803 236
rect 3857 216 3869 236
rect 3879 196 3891 236
rect 3899 196 3911 236
rect 3999 196 4011 236
rect 4029 196 4041 236
rect 4117 196 4129 236
rect 4147 196 4159 236
rect 4167 196 4179 236
rect 4291 216 4303 236
rect 4311 216 4323 236
rect 4331 216 4343 236
rect 4399 196 4411 236
rect 4429 196 4441 236
rect 4554 178 4566 236
rect 4590 176 4602 236
rect 4691 196 4703 236
rect 4711 196 4723 236
rect 4731 208 4743 236
rect 4751 196 4763 236
rect 4819 196 4831 236
rect 4849 196 4861 236
rect 4951 196 4963 236
rect 4971 196 4983 236
rect 4991 208 5003 236
rect 5011 196 5023 236
rect 5077 216 5089 236
rect 5097 216 5109 236
rect 5117 216 5129 236
rect 5219 196 5231 236
rect 5249 196 5261 236
rect 5317 208 5329 228
rect 5337 208 5349 228
rect 5367 196 5379 228
rect 5397 188 5409 228
rect 5477 216 5489 236
rect 5497 216 5509 236
rect 5591 216 5603 236
rect 5611 216 5623 236
rect 5679 196 5691 236
rect 5709 196 5721 236
<< pdcontact >>
rect 76 5716 88 5756
rect 98 5676 110 5756
rect 126 5676 138 5756
rect 202 5676 214 5756
rect 230 5676 242 5756
rect 252 5716 264 5756
rect 371 5676 383 5756
rect 391 5676 403 5756
rect 411 5688 423 5756
rect 431 5684 443 5756
rect 497 5716 509 5756
rect 517 5716 529 5756
rect 537 5720 549 5756
rect 557 5716 569 5756
rect 656 5716 668 5756
rect 678 5676 690 5756
rect 706 5676 718 5756
rect 791 5716 803 5756
rect 811 5716 823 5756
rect 831 5716 843 5756
rect 911 5676 923 5756
rect 931 5676 943 5756
rect 951 5688 963 5756
rect 971 5684 983 5756
rect 1057 5676 1069 5756
rect 1085 5676 1097 5756
rect 1221 5677 1233 5756
rect 1241 5677 1253 5756
rect 1271 5676 1283 5756
rect 1347 5676 1359 5756
rect 1367 5676 1379 5756
rect 1391 5716 1403 5756
rect 1411 5716 1423 5756
rect 1491 5716 1503 5756
rect 1511 5720 1523 5756
rect 1531 5716 1543 5756
rect 1551 5716 1563 5756
rect 1651 5676 1663 5756
rect 1671 5676 1683 5756
rect 1691 5688 1703 5756
rect 1711 5684 1723 5756
rect 1791 5716 1803 5756
rect 1811 5720 1823 5756
rect 1831 5716 1843 5756
rect 1851 5716 1863 5756
rect 1917 5716 1929 5756
rect 1937 5716 1949 5756
rect 2036 5716 2048 5756
rect 2058 5676 2070 5756
rect 2086 5676 2098 5756
rect 2162 5676 2174 5756
rect 2190 5676 2202 5756
rect 2212 5716 2224 5756
rect 2297 5684 2309 5756
rect 2317 5688 2329 5756
rect 2337 5676 2349 5756
rect 2357 5676 2369 5756
rect 2451 5716 2463 5756
rect 2471 5716 2483 5756
rect 2491 5716 2503 5756
rect 2571 5716 2583 5756
rect 2591 5720 2603 5756
rect 2611 5716 2623 5756
rect 2631 5716 2643 5756
rect 2711 5716 2723 5756
rect 2731 5720 2743 5756
rect 2751 5716 2763 5756
rect 2771 5716 2783 5756
rect 2837 5716 2849 5756
rect 2857 5716 2869 5756
rect 2877 5716 2889 5756
rect 2971 5716 2983 5756
rect 2991 5716 3003 5756
rect 3076 5716 3088 5756
rect 3098 5676 3110 5756
rect 3126 5676 3138 5756
rect 3227 5676 3239 5756
rect 3247 5676 3259 5756
rect 3271 5716 3283 5756
rect 3291 5716 3303 5756
rect 3383 5676 3395 5756
rect 3411 5676 3423 5756
rect 3491 5716 3503 5756
rect 3511 5720 3523 5756
rect 3531 5716 3543 5756
rect 3551 5716 3563 5756
rect 3651 5716 3663 5756
rect 3671 5716 3683 5756
rect 3751 5716 3763 5756
rect 3771 5716 3783 5756
rect 3837 5716 3849 5756
rect 3857 5716 3869 5756
rect 3942 5676 3954 5756
rect 3970 5676 3982 5756
rect 3992 5716 4004 5756
rect 4077 5716 4089 5756
rect 4097 5716 4109 5756
rect 4137 5676 4149 5756
rect 4157 5736 4169 5756
rect 4187 5736 4199 5756
rect 4215 5716 4227 5756
rect 4241 5716 4253 5756
rect 4261 5716 4273 5756
rect 4293 5716 4305 5756
rect 4327 5716 4339 5756
rect 4347 5676 4359 5756
rect 4456 5716 4468 5756
rect 4478 5676 4490 5756
rect 4506 5676 4518 5756
rect 4591 5676 4603 5756
rect 4611 5676 4623 5756
rect 4631 5676 4643 5756
rect 4651 5676 4663 5756
rect 4671 5676 4683 5756
rect 4691 5676 4703 5756
rect 4711 5676 4723 5756
rect 4731 5676 4743 5756
rect 4751 5676 4763 5756
rect 4831 5716 4843 5756
rect 4851 5716 4863 5756
rect 4936 5716 4948 5756
rect 4958 5676 4970 5756
rect 4986 5676 4998 5756
rect 5071 5716 5083 5756
rect 5091 5716 5103 5756
rect 5111 5716 5123 5756
rect 5177 5716 5189 5756
rect 5197 5716 5209 5756
rect 5217 5716 5229 5756
rect 5302 5676 5314 5756
rect 5330 5676 5342 5756
rect 5352 5716 5364 5756
rect 5437 5716 5449 5756
rect 5457 5716 5469 5756
rect 5537 5716 5549 5756
rect 5557 5716 5569 5756
rect 5577 5716 5589 5756
rect 5657 5716 5669 5756
rect 5677 5716 5689 5756
rect 76 5304 88 5344
rect 98 5304 110 5384
rect 126 5304 138 5384
rect 231 5304 243 5344
rect 251 5304 263 5340
rect 271 5304 283 5344
rect 291 5304 303 5344
rect 371 5304 383 5344
rect 391 5304 403 5340
rect 411 5304 423 5344
rect 431 5304 443 5344
rect 511 5304 523 5344
rect 531 5304 543 5340
rect 551 5304 563 5344
rect 571 5304 583 5344
rect 657 5304 669 5344
rect 677 5304 689 5344
rect 697 5304 709 5340
rect 717 5304 729 5344
rect 802 5304 814 5384
rect 830 5304 842 5384
rect 852 5304 864 5344
rect 937 5304 949 5344
rect 957 5304 969 5344
rect 977 5304 989 5340
rect 997 5304 1009 5344
rect 1091 5304 1103 5384
rect 1111 5304 1123 5384
rect 1131 5304 1143 5372
rect 1151 5304 1163 5376
rect 1217 5304 1229 5344
rect 1237 5304 1249 5344
rect 1257 5304 1269 5340
rect 1277 5304 1289 5344
rect 1377 5304 1389 5384
rect 1405 5304 1417 5384
rect 1511 5304 1523 5344
rect 1531 5304 1543 5340
rect 1551 5304 1563 5344
rect 1571 5304 1583 5344
rect 1642 5304 1654 5384
rect 1670 5304 1682 5384
rect 1692 5304 1704 5344
rect 1791 5304 1803 5344
rect 1811 5304 1823 5340
rect 1831 5304 1843 5344
rect 1851 5304 1863 5344
rect 1931 5304 1943 5344
rect 1951 5304 1963 5340
rect 1971 5304 1983 5344
rect 1991 5304 2003 5344
rect 2057 5304 2069 5344
rect 2077 5304 2089 5344
rect 2097 5304 2109 5344
rect 2211 5304 2223 5344
rect 2231 5304 2243 5344
rect 2307 5304 2319 5384
rect 2327 5304 2339 5384
rect 2351 5304 2363 5344
rect 2371 5304 2383 5344
rect 2442 5304 2454 5384
rect 2470 5304 2482 5384
rect 2492 5304 2504 5344
rect 2611 5304 2623 5344
rect 2631 5304 2643 5340
rect 2651 5304 2663 5344
rect 2671 5304 2683 5344
rect 2751 5304 2763 5344
rect 2771 5304 2783 5340
rect 2791 5304 2803 5344
rect 2811 5304 2823 5344
rect 2882 5304 2894 5384
rect 2910 5304 2922 5384
rect 2932 5304 2944 5344
rect 3017 5304 3029 5344
rect 3037 5304 3049 5344
rect 3117 5304 3129 5344
rect 3137 5304 3149 5344
rect 3157 5304 3169 5344
rect 3257 5304 3269 5344
rect 3277 5304 3289 5344
rect 3297 5304 3309 5340
rect 3317 5304 3329 5344
rect 3397 5304 3409 5344
rect 3417 5304 3429 5344
rect 3437 5304 3449 5344
rect 3517 5304 3529 5384
rect 3547 5304 3559 5383
rect 3567 5304 3579 5383
rect 3671 5304 3683 5344
rect 3691 5304 3703 5340
rect 3711 5304 3723 5344
rect 3731 5304 3743 5344
rect 3811 5304 3823 5384
rect 3831 5304 3843 5384
rect 3851 5304 3863 5372
rect 3871 5304 3883 5376
rect 3937 5304 3949 5344
rect 3957 5304 3969 5344
rect 3977 5304 3989 5344
rect 4076 5304 4088 5344
rect 4098 5304 4110 5384
rect 4126 5304 4138 5384
rect 4211 5304 4223 5344
rect 4231 5304 4243 5344
rect 4251 5304 4263 5344
rect 4331 5304 4343 5344
rect 4351 5304 4363 5340
rect 4371 5304 4383 5344
rect 4391 5304 4403 5344
rect 4477 5304 4489 5376
rect 4497 5304 4509 5372
rect 4517 5304 4529 5384
rect 4537 5304 4549 5384
rect 4617 5304 4629 5344
rect 4637 5304 4649 5344
rect 4722 5304 4734 5384
rect 4750 5304 4762 5384
rect 4772 5304 4784 5344
rect 4817 5304 4829 5384
rect 4837 5304 4849 5324
rect 4867 5304 4879 5324
rect 4895 5304 4907 5344
rect 4921 5304 4933 5344
rect 4941 5304 4953 5344
rect 4973 5304 4985 5344
rect 5007 5304 5019 5344
rect 5027 5304 5039 5384
rect 5097 5304 5109 5344
rect 5117 5304 5129 5344
rect 5157 5304 5169 5384
rect 5177 5304 5189 5324
rect 5207 5304 5219 5324
rect 5235 5304 5247 5344
rect 5261 5304 5273 5344
rect 5281 5304 5293 5344
rect 5313 5304 5325 5344
rect 5347 5304 5359 5344
rect 5367 5304 5379 5384
rect 5442 5304 5454 5384
rect 5470 5304 5482 5384
rect 5492 5304 5504 5344
rect 5597 5304 5609 5344
rect 5617 5304 5629 5344
rect 5637 5304 5649 5344
rect 5717 5304 5729 5344
rect 5737 5304 5749 5344
rect 5757 5304 5769 5344
rect 71 5236 83 5276
rect 91 5240 103 5276
rect 111 5236 123 5276
rect 131 5236 143 5276
rect 197 5204 209 5276
rect 217 5208 229 5276
rect 237 5196 249 5276
rect 257 5196 269 5276
rect 337 5236 349 5276
rect 357 5236 369 5276
rect 451 5236 463 5276
rect 471 5240 483 5276
rect 491 5236 503 5276
rect 511 5236 523 5276
rect 577 5204 589 5276
rect 597 5208 609 5276
rect 617 5196 629 5276
rect 637 5196 649 5276
rect 731 5196 743 5276
rect 751 5196 763 5276
rect 771 5208 783 5276
rect 791 5204 803 5276
rect 857 5236 869 5276
rect 877 5236 889 5276
rect 897 5240 909 5276
rect 917 5236 929 5276
rect 1011 5236 1023 5276
rect 1031 5240 1043 5276
rect 1051 5236 1063 5276
rect 1071 5236 1083 5276
rect 1137 5236 1149 5276
rect 1157 5236 1169 5276
rect 1251 5236 1263 5276
rect 1271 5240 1283 5276
rect 1291 5236 1303 5276
rect 1311 5236 1323 5276
rect 1416 5236 1428 5276
rect 1438 5196 1450 5276
rect 1466 5196 1478 5276
rect 1551 5236 1563 5276
rect 1571 5236 1583 5276
rect 1656 5236 1668 5276
rect 1678 5196 1690 5276
rect 1706 5196 1718 5276
rect 1807 5208 1819 5268
rect 1827 5212 1839 5264
rect 1847 5208 1859 5268
rect 1871 5218 1883 5276
rect 1891 5216 1903 5264
rect 1911 5216 1923 5276
rect 1931 5216 1943 5276
rect 1951 5216 1963 5276
rect 2031 5196 2043 5276
rect 2051 5196 2063 5264
rect 2071 5198 2083 5276
rect 2091 5210 2103 5276
rect 2111 5198 2123 5276
rect 2177 5236 2189 5276
rect 2197 5236 2209 5276
rect 2217 5236 2229 5276
rect 2311 5236 2323 5276
rect 2331 5240 2343 5276
rect 2351 5236 2363 5276
rect 2371 5236 2383 5276
rect 2451 5196 2463 5276
rect 2471 5196 2483 5276
rect 2491 5208 2503 5276
rect 2511 5204 2523 5276
rect 2591 5236 2603 5276
rect 2611 5236 2623 5276
rect 2696 5236 2708 5276
rect 2718 5196 2730 5276
rect 2746 5196 2758 5276
rect 2856 5236 2868 5276
rect 2878 5196 2890 5276
rect 2906 5196 2918 5276
rect 2987 5196 2999 5276
rect 3007 5196 3019 5276
rect 3031 5236 3043 5276
rect 3051 5236 3063 5276
rect 3117 5196 3129 5276
rect 3145 5196 3157 5276
rect 3271 5236 3283 5276
rect 3291 5236 3303 5276
rect 3383 5196 3395 5276
rect 3411 5196 3423 5276
rect 3516 5236 3528 5276
rect 3538 5196 3550 5276
rect 3566 5196 3578 5276
rect 3637 5236 3649 5276
rect 3657 5236 3669 5276
rect 3677 5236 3689 5276
rect 3771 5236 3783 5276
rect 3791 5236 3803 5276
rect 3811 5236 3823 5276
rect 3911 5236 3923 5276
rect 3931 5236 3943 5276
rect 3951 5236 3963 5276
rect 4017 5236 4029 5276
rect 4037 5236 4049 5276
rect 4057 5240 4069 5276
rect 4077 5236 4089 5276
rect 4176 5236 4188 5276
rect 4198 5196 4210 5276
rect 4226 5196 4238 5276
rect 4322 5196 4334 5276
rect 4350 5196 4362 5276
rect 4372 5236 4384 5276
rect 4457 5236 4469 5276
rect 4477 5236 4489 5276
rect 4571 5236 4583 5276
rect 4591 5240 4603 5276
rect 4611 5236 4623 5276
rect 4631 5236 4643 5276
rect 4697 5204 4709 5276
rect 4717 5208 4729 5276
rect 4737 5196 4749 5276
rect 4757 5196 4769 5276
rect 4837 5196 4849 5276
rect 4865 5196 4877 5276
rect 4917 5196 4929 5276
rect 4937 5256 4949 5276
rect 4967 5256 4979 5276
rect 4995 5236 5007 5276
rect 5021 5236 5033 5276
rect 5041 5236 5053 5276
rect 5073 5236 5085 5276
rect 5107 5236 5119 5276
rect 5127 5196 5139 5276
rect 5202 5196 5214 5276
rect 5230 5196 5242 5276
rect 5252 5236 5264 5276
rect 5337 5236 5349 5276
rect 5357 5236 5369 5276
rect 5442 5196 5454 5276
rect 5470 5196 5482 5276
rect 5492 5236 5504 5276
rect 5591 5236 5603 5276
rect 5611 5236 5623 5276
rect 5631 5236 5643 5276
rect 5697 5236 5709 5276
rect 5717 5236 5729 5276
rect 5737 5236 5749 5276
rect 76 4824 88 4864
rect 98 4824 110 4904
rect 126 4824 138 4904
rect 211 4824 223 4864
rect 231 4824 243 4860
rect 251 4824 263 4864
rect 271 4824 283 4864
rect 337 4824 349 4864
rect 357 4824 369 4864
rect 377 4824 389 4860
rect 397 4824 409 4864
rect 482 4824 494 4904
rect 510 4824 522 4904
rect 532 4824 544 4864
rect 631 4824 643 4864
rect 651 4824 663 4864
rect 671 4824 683 4864
rect 756 4824 768 4864
rect 778 4824 790 4904
rect 806 4824 818 4904
rect 896 4824 908 4864
rect 918 4824 930 4904
rect 946 4824 958 4904
rect 1031 4824 1043 4904
rect 1051 4824 1063 4904
rect 1071 4824 1083 4892
rect 1091 4824 1103 4896
rect 1176 4824 1188 4864
rect 1198 4824 1210 4904
rect 1226 4824 1238 4904
rect 1311 4824 1323 4864
rect 1331 4824 1343 4864
rect 1411 4824 1423 4864
rect 1431 4824 1443 4864
rect 1451 4824 1463 4864
rect 1551 4824 1563 4864
rect 1571 4824 1583 4860
rect 1591 4824 1603 4864
rect 1611 4824 1623 4864
rect 1696 4824 1708 4864
rect 1718 4824 1730 4904
rect 1746 4824 1758 4904
rect 1817 4824 1829 4896
rect 1837 4824 1849 4892
rect 1857 4824 1869 4904
rect 1877 4824 1889 4904
rect 1957 4824 1969 4864
rect 1977 4824 1989 4864
rect 1997 4824 2009 4864
rect 2091 4824 2103 4904
rect 2111 4824 2123 4904
rect 2131 4824 2143 4892
rect 2151 4824 2163 4896
rect 2251 4824 2263 4864
rect 2271 4824 2283 4864
rect 2356 4824 2368 4864
rect 2378 4824 2390 4904
rect 2406 4824 2418 4904
rect 2491 4824 2503 4864
rect 2511 4824 2523 4860
rect 2531 4824 2543 4864
rect 2551 4824 2563 4864
rect 2631 4824 2643 4864
rect 2651 4824 2663 4864
rect 2751 4824 2763 4864
rect 2771 4824 2783 4864
rect 2791 4824 2803 4864
rect 2857 4824 2869 4864
rect 2877 4824 2889 4864
rect 2957 4824 2969 4864
rect 2977 4824 2989 4864
rect 2997 4824 3009 4860
rect 3017 4824 3029 4864
rect 3116 4824 3128 4864
rect 3138 4824 3150 4904
rect 3166 4824 3178 4904
rect 3256 4824 3268 4864
rect 3278 4824 3290 4904
rect 3306 4824 3318 4904
rect 3391 4824 3403 4904
rect 3411 4824 3423 4904
rect 3431 4824 3443 4892
rect 3451 4824 3463 4896
rect 3517 4824 3529 4904
rect 3547 4824 3559 4903
rect 3567 4824 3579 4903
rect 3683 4824 3695 4904
rect 3711 4824 3723 4904
rect 3791 4824 3803 4864
rect 3811 4824 3823 4860
rect 3831 4824 3843 4864
rect 3851 4824 3863 4864
rect 3931 4824 3943 4864
rect 3951 4824 3963 4864
rect 4017 4824 4029 4864
rect 4037 4824 4049 4864
rect 4057 4824 4069 4860
rect 4077 4824 4089 4864
rect 4157 4824 4169 4864
rect 4177 4824 4189 4864
rect 4197 4824 4209 4860
rect 4217 4824 4229 4864
rect 4307 4824 4319 4904
rect 4327 4824 4339 4904
rect 4351 4824 4363 4864
rect 4371 4824 4383 4864
rect 4457 4824 4469 4904
rect 4487 4824 4499 4903
rect 4507 4824 4519 4903
rect 4597 4824 4609 4904
rect 4625 4824 4637 4904
rect 4736 4824 4748 4864
rect 4758 4824 4770 4904
rect 4786 4824 4798 4904
rect 4817 4824 4829 4904
rect 4837 4824 4849 4844
rect 4867 4824 4879 4844
rect 4895 4824 4907 4864
rect 4921 4824 4933 4864
rect 4941 4824 4953 4864
rect 4973 4824 4985 4864
rect 5007 4824 5019 4864
rect 5027 4824 5039 4904
rect 5102 4824 5114 4904
rect 5130 4824 5142 4904
rect 5152 4824 5164 4864
rect 5197 4824 5209 4904
rect 5217 4824 5229 4844
rect 5247 4824 5259 4844
rect 5275 4824 5287 4864
rect 5301 4824 5313 4864
rect 5321 4824 5333 4864
rect 5353 4824 5365 4864
rect 5387 4824 5399 4864
rect 5407 4824 5419 4904
rect 5491 4824 5503 4864
rect 5511 4824 5523 4864
rect 5531 4824 5543 4864
rect 5597 4824 5609 4864
rect 5617 4824 5629 4864
rect 5637 4824 5649 4864
rect 5737 4824 5749 4864
rect 5757 4824 5769 4864
rect 5777 4824 5789 4864
rect 71 4716 83 4796
rect 91 4716 103 4796
rect 111 4728 123 4796
rect 131 4724 143 4796
rect 211 4756 223 4796
rect 231 4760 243 4796
rect 251 4756 263 4796
rect 271 4756 283 4796
rect 337 4724 349 4796
rect 357 4728 369 4796
rect 377 4716 389 4796
rect 397 4716 409 4796
rect 477 4756 489 4796
rect 497 4756 509 4796
rect 517 4756 529 4796
rect 611 4756 623 4796
rect 631 4760 643 4796
rect 651 4756 663 4796
rect 671 4756 683 4796
rect 771 4756 783 4796
rect 791 4760 803 4796
rect 811 4756 823 4796
rect 831 4756 843 4796
rect 897 4756 909 4796
rect 917 4756 929 4796
rect 997 4756 1009 4796
rect 1017 4756 1029 4796
rect 1111 4756 1123 4796
rect 1131 4756 1143 4796
rect 1216 4756 1228 4796
rect 1238 4716 1250 4796
rect 1266 4716 1278 4796
rect 1342 4716 1354 4796
rect 1370 4716 1382 4796
rect 1392 4756 1404 4796
rect 1477 4756 1489 4796
rect 1497 4756 1509 4796
rect 1577 4756 1589 4796
rect 1597 4756 1609 4796
rect 1617 4760 1629 4796
rect 1637 4756 1649 4796
rect 1736 4756 1748 4796
rect 1758 4716 1770 4796
rect 1786 4716 1798 4796
rect 1871 4756 1883 4796
rect 1891 4756 1903 4796
rect 1911 4756 1923 4796
rect 1982 4716 1994 4796
rect 2010 4716 2022 4796
rect 2032 4756 2044 4796
rect 2131 4756 2143 4796
rect 2151 4760 2163 4796
rect 2171 4756 2183 4796
rect 2191 4756 2203 4796
rect 2269 4716 2281 4796
rect 2289 4716 2301 4796
rect 2311 4756 2323 4796
rect 2377 4756 2389 4796
rect 2397 4756 2409 4796
rect 2417 4756 2429 4796
rect 2497 4756 2509 4796
rect 2517 4756 2529 4796
rect 2537 4756 2549 4796
rect 2629 4716 2641 4796
rect 2649 4716 2661 4796
rect 2671 4756 2683 4796
rect 2737 4756 2749 4796
rect 2757 4756 2769 4796
rect 2777 4760 2789 4796
rect 2797 4756 2809 4796
rect 2903 4716 2915 4796
rect 2931 4716 2943 4796
rect 3017 4716 3029 4796
rect 3047 4716 3069 4796
rect 3087 4716 3099 4796
rect 3191 4756 3203 4796
rect 3211 4756 3223 4796
rect 3231 4756 3243 4796
rect 3311 4756 3323 4796
rect 3331 4760 3343 4796
rect 3351 4756 3363 4796
rect 3371 4756 3383 4796
rect 3451 4716 3463 4796
rect 3471 4716 3483 4796
rect 3491 4728 3503 4796
rect 3511 4724 3523 4796
rect 3591 4756 3603 4796
rect 3611 4760 3623 4796
rect 3631 4756 3643 4796
rect 3651 4756 3663 4796
rect 3731 4716 3743 4796
rect 3751 4716 3763 4796
rect 3771 4728 3783 4796
rect 3791 4724 3803 4796
rect 3857 4756 3869 4796
rect 3877 4756 3889 4796
rect 3897 4760 3909 4796
rect 3917 4756 3929 4796
rect 3997 4756 4009 4796
rect 4017 4756 4029 4796
rect 4037 4760 4049 4796
rect 4057 4756 4069 4796
rect 4137 4756 4149 4796
rect 4157 4756 4169 4796
rect 4247 4716 4259 4796
rect 4267 4716 4279 4796
rect 4291 4756 4303 4796
rect 4311 4756 4323 4796
rect 4411 4756 4423 4796
rect 4431 4760 4443 4796
rect 4451 4756 4463 4796
rect 4471 4756 4483 4796
rect 4537 4756 4549 4796
rect 4557 4756 4569 4796
rect 4577 4760 4589 4796
rect 4597 4756 4609 4796
rect 4677 4756 4689 4796
rect 4697 4756 4709 4796
rect 4737 4716 4749 4796
rect 4757 4776 4769 4796
rect 4787 4776 4799 4796
rect 4815 4756 4827 4796
rect 4841 4756 4853 4796
rect 4861 4756 4873 4796
rect 4893 4756 4905 4796
rect 4927 4756 4939 4796
rect 4947 4716 4959 4796
rect 5022 4716 5034 4796
rect 5050 4716 5062 4796
rect 5072 4756 5084 4796
rect 5157 4756 5169 4796
rect 5177 4756 5189 4796
rect 5197 4756 5209 4796
rect 5277 4756 5289 4796
rect 5297 4756 5309 4796
rect 5317 4756 5329 4796
rect 5417 4756 5429 4796
rect 5437 4756 5449 4796
rect 5457 4756 5469 4796
rect 5537 4756 5549 4796
rect 5557 4756 5569 4796
rect 5577 4756 5589 4796
rect 5671 4756 5683 4796
rect 5691 4760 5703 4796
rect 5711 4756 5723 4796
rect 5731 4756 5743 4796
rect 76 4344 88 4384
rect 98 4344 110 4424
rect 126 4344 138 4424
rect 211 4344 223 4384
rect 231 4344 243 4380
rect 251 4344 263 4384
rect 271 4344 283 4384
rect 337 4344 349 4416
rect 357 4344 369 4412
rect 377 4344 389 4424
rect 397 4344 409 4424
rect 516 4344 528 4384
rect 538 4344 550 4424
rect 566 4344 578 4424
rect 656 4344 668 4384
rect 678 4344 690 4424
rect 706 4344 718 4424
rect 777 4344 789 4384
rect 797 4344 809 4384
rect 877 4344 889 4416
rect 897 4344 909 4412
rect 917 4344 929 4424
rect 937 4344 949 4424
rect 1031 4344 1043 4384
rect 1051 4344 1063 4384
rect 1131 4344 1143 4384
rect 1151 4344 1163 4380
rect 1171 4344 1183 4384
rect 1191 4344 1203 4384
rect 1271 4344 1283 4424
rect 1291 4344 1303 4424
rect 1311 4344 1323 4412
rect 1331 4344 1343 4416
rect 1411 4344 1423 4384
rect 1431 4344 1443 4384
rect 1502 4344 1514 4424
rect 1530 4344 1542 4424
rect 1552 4344 1564 4384
rect 1651 4344 1663 4384
rect 1671 4344 1683 4384
rect 1691 4344 1703 4384
rect 1771 4344 1783 4384
rect 1791 4344 1803 4380
rect 1811 4344 1823 4384
rect 1831 4344 1843 4384
rect 1923 4344 1935 4424
rect 1951 4344 1963 4424
rect 2031 4344 2043 4384
rect 2051 4344 2063 4380
rect 2071 4344 2083 4384
rect 2091 4344 2103 4384
rect 2191 4344 2203 4384
rect 2211 4344 2223 4380
rect 2231 4344 2243 4384
rect 2251 4344 2263 4384
rect 2331 4344 2343 4384
rect 2351 4344 2363 4384
rect 2371 4344 2383 4384
rect 2451 4344 2463 4384
rect 2471 4344 2483 4380
rect 2491 4344 2503 4384
rect 2511 4344 2523 4384
rect 2577 4344 2589 4384
rect 2597 4344 2609 4384
rect 2617 4344 2629 4380
rect 2637 4344 2649 4384
rect 2731 4344 2743 4384
rect 2751 4344 2763 4384
rect 2843 4344 2855 4424
rect 2871 4344 2883 4424
rect 2951 4344 2963 4384
rect 2971 4344 2983 4380
rect 2991 4344 3003 4384
rect 3011 4344 3023 4384
rect 3091 4344 3103 4384
rect 3111 4344 3123 4380
rect 3131 4344 3143 4384
rect 3151 4344 3163 4384
rect 3217 4344 3229 4384
rect 3237 4344 3249 4384
rect 3322 4344 3334 4424
rect 3350 4344 3362 4424
rect 3372 4344 3384 4384
rect 3467 4344 3479 4424
rect 3487 4344 3499 4424
rect 3511 4344 3523 4384
rect 3531 4344 3543 4384
rect 3617 4344 3629 4384
rect 3637 4344 3649 4384
rect 3657 4344 3669 4384
rect 3761 4344 3773 4423
rect 3781 4344 3793 4423
rect 3811 4344 3823 4424
rect 3877 4344 3889 4384
rect 3897 4344 3909 4384
rect 3917 4344 3929 4384
rect 4009 4344 4021 4424
rect 4029 4344 4041 4424
rect 4051 4344 4063 4384
rect 4117 4344 4129 4384
rect 4137 4344 4149 4384
rect 4161 4344 4173 4424
rect 4181 4344 4193 4424
rect 4271 4344 4283 4384
rect 4291 4344 4303 4384
rect 4311 4344 4323 4384
rect 4396 4344 4408 4384
rect 4418 4344 4430 4424
rect 4446 4344 4458 4424
rect 4517 4344 4529 4384
rect 4537 4344 4549 4384
rect 4557 4344 4569 4384
rect 4651 4344 4663 4384
rect 4671 4344 4683 4384
rect 4691 4344 4703 4384
rect 4757 4344 4769 4384
rect 4777 4344 4789 4384
rect 4857 4344 4869 4384
rect 4877 4344 4889 4384
rect 4897 4344 4909 4384
rect 4982 4344 4994 4424
rect 5010 4344 5022 4424
rect 5032 4344 5044 4384
rect 5077 4344 5089 4424
rect 5097 4344 5109 4364
rect 5127 4344 5139 4364
rect 5155 4344 5167 4384
rect 5181 4344 5193 4384
rect 5201 4344 5213 4384
rect 5233 4344 5245 4384
rect 5267 4344 5279 4384
rect 5287 4344 5299 4424
rect 5362 4344 5374 4424
rect 5390 4344 5402 4424
rect 5412 4344 5424 4384
rect 5497 4344 5509 4424
rect 5527 4344 5539 4423
rect 5547 4344 5559 4423
rect 5656 4344 5668 4384
rect 5678 4344 5690 4424
rect 5706 4344 5718 4424
rect 96 4276 108 4316
rect 118 4236 130 4316
rect 146 4236 158 4316
rect 236 4276 248 4316
rect 258 4236 270 4316
rect 286 4236 298 4316
rect 391 4276 403 4316
rect 411 4280 423 4316
rect 431 4276 443 4316
rect 451 4276 463 4316
rect 531 4276 543 4316
rect 551 4280 563 4316
rect 571 4276 583 4316
rect 591 4276 603 4316
rect 681 4237 693 4316
rect 701 4237 713 4316
rect 731 4236 743 4316
rect 816 4276 828 4316
rect 838 4236 850 4316
rect 866 4236 878 4316
rect 937 4276 949 4316
rect 957 4276 969 4316
rect 1051 4236 1063 4316
rect 1071 4236 1083 4316
rect 1091 4248 1103 4316
rect 1111 4244 1123 4316
rect 1211 4276 1223 4316
rect 1231 4280 1243 4316
rect 1251 4276 1263 4316
rect 1271 4276 1283 4316
rect 1351 4276 1363 4316
rect 1371 4276 1383 4316
rect 1391 4276 1403 4316
rect 1471 4276 1483 4316
rect 1491 4276 1503 4316
rect 1511 4276 1523 4316
rect 1603 4236 1615 4316
rect 1631 4236 1643 4316
rect 1711 4276 1723 4316
rect 1731 4280 1743 4316
rect 1751 4276 1763 4316
rect 1771 4276 1783 4316
rect 1851 4276 1863 4316
rect 1871 4280 1883 4316
rect 1891 4276 1903 4316
rect 1911 4276 1923 4316
rect 1977 4276 1989 4316
rect 1997 4276 2009 4316
rect 2017 4280 2029 4316
rect 2037 4276 2049 4316
rect 2117 4276 2129 4316
rect 2137 4276 2149 4316
rect 2157 4280 2169 4316
rect 2177 4276 2189 4316
rect 2283 4236 2295 4316
rect 2311 4236 2323 4316
rect 2416 4276 2428 4316
rect 2438 4236 2450 4316
rect 2466 4236 2478 4316
rect 2571 4276 2583 4316
rect 2591 4280 2603 4316
rect 2611 4276 2623 4316
rect 2631 4276 2643 4316
rect 2697 4276 2709 4316
rect 2717 4276 2729 4316
rect 2817 4276 2829 4316
rect 2837 4276 2849 4316
rect 2857 4280 2869 4316
rect 2877 4276 2889 4316
rect 2957 4276 2969 4316
rect 2977 4276 2989 4316
rect 2997 4276 3009 4316
rect 3077 4244 3089 4316
rect 3097 4248 3109 4316
rect 3117 4236 3129 4316
rect 3137 4236 3149 4316
rect 3217 4244 3229 4316
rect 3237 4248 3249 4316
rect 3257 4236 3269 4316
rect 3277 4236 3289 4316
rect 3362 4236 3374 4316
rect 3390 4236 3402 4316
rect 3412 4276 3424 4316
rect 3517 4276 3529 4316
rect 3537 4276 3549 4316
rect 3617 4276 3629 4316
rect 3637 4276 3649 4316
rect 3657 4280 3669 4316
rect 3677 4276 3689 4316
rect 3757 4276 3769 4316
rect 3777 4276 3789 4316
rect 3797 4280 3809 4316
rect 3817 4276 3829 4316
rect 3911 4276 3923 4316
rect 3931 4276 3943 4316
rect 3951 4276 3963 4316
rect 4051 4276 4063 4316
rect 4071 4276 4083 4316
rect 4091 4276 4103 4316
rect 4171 4276 4183 4316
rect 4191 4276 4203 4316
rect 4211 4276 4223 4316
rect 4296 4276 4308 4316
rect 4318 4236 4330 4316
rect 4346 4236 4358 4316
rect 4417 4236 4429 4316
rect 4447 4237 4459 4316
rect 4467 4237 4479 4316
rect 4576 4276 4588 4316
rect 4598 4236 4610 4316
rect 4626 4236 4638 4316
rect 4722 4236 4734 4316
rect 4750 4236 4762 4316
rect 4772 4276 4784 4316
rect 4857 4236 4869 4316
rect 4885 4236 4897 4316
rect 4977 4276 4989 4316
rect 4997 4276 5009 4316
rect 5097 4244 5109 4316
rect 5117 4248 5129 4316
rect 5137 4236 5149 4316
rect 5157 4236 5169 4316
rect 5242 4236 5254 4316
rect 5270 4236 5282 4316
rect 5292 4276 5304 4316
rect 5377 4276 5389 4316
rect 5397 4276 5409 4316
rect 5482 4236 5494 4316
rect 5510 4236 5522 4316
rect 5532 4276 5544 4316
rect 5581 4236 5593 4316
rect 5601 4276 5613 4316
rect 5635 4276 5647 4316
rect 5667 4276 5679 4316
rect 5687 4276 5699 4316
rect 5713 4276 5725 4316
rect 5741 4296 5753 4316
rect 5771 4296 5783 4316
rect 5791 4236 5803 4316
rect 71 3864 83 3904
rect 91 3864 103 3904
rect 182 3864 194 3944
rect 210 3864 222 3944
rect 232 3864 244 3904
rect 331 3864 343 3904
rect 351 3864 363 3904
rect 437 3864 449 3936
rect 457 3864 469 3932
rect 477 3864 489 3944
rect 497 3864 509 3944
rect 603 3864 615 3944
rect 631 3864 643 3944
rect 731 3864 743 3904
rect 751 3864 763 3904
rect 822 3864 834 3944
rect 850 3864 862 3944
rect 872 3864 884 3904
rect 957 3864 969 3904
rect 977 3864 989 3904
rect 1057 3864 1069 3904
rect 1077 3864 1089 3904
rect 1097 3864 1109 3900
rect 1117 3864 1129 3904
rect 1197 3864 1209 3942
rect 1217 3864 1229 3930
rect 1237 3864 1249 3942
rect 1257 3876 1269 3944
rect 1277 3864 1289 3944
rect 1377 3864 1389 3904
rect 1397 3864 1409 3904
rect 1417 3864 1429 3904
rect 1511 3864 1523 3904
rect 1531 3864 1543 3904
rect 1623 3864 1635 3944
rect 1651 3864 1663 3944
rect 1731 3864 1743 3904
rect 1751 3864 1763 3904
rect 1817 3864 1829 3904
rect 1837 3864 1849 3904
rect 1857 3864 1869 3900
rect 1877 3864 1889 3904
rect 1976 3864 1988 3904
rect 1998 3864 2010 3944
rect 2026 3864 2038 3944
rect 2131 3864 2143 3904
rect 2151 3864 2163 3900
rect 2171 3864 2183 3904
rect 2191 3864 2203 3904
rect 2257 3864 2269 3904
rect 2277 3864 2289 3904
rect 2297 3864 2309 3900
rect 2317 3864 2329 3904
rect 2416 3864 2428 3904
rect 2438 3864 2450 3944
rect 2466 3864 2478 3944
rect 2551 3864 2563 3904
rect 2571 3864 2583 3904
rect 2591 3864 2603 3904
rect 2657 3864 2669 3904
rect 2677 3864 2689 3904
rect 2697 3864 2709 3904
rect 2777 3864 2789 3904
rect 2797 3864 2809 3904
rect 2817 3864 2829 3900
rect 2837 3864 2849 3904
rect 2917 3864 2929 3904
rect 2937 3864 2949 3904
rect 2957 3864 2969 3900
rect 2977 3864 2989 3904
rect 3071 3864 3083 3904
rect 3091 3864 3103 3904
rect 3171 3864 3183 3904
rect 3191 3864 3203 3900
rect 3211 3864 3223 3904
rect 3231 3864 3243 3904
rect 3311 3864 3323 3904
rect 3331 3864 3343 3904
rect 3416 3864 3428 3904
rect 3438 3864 3450 3944
rect 3466 3864 3478 3944
rect 3537 3864 3549 3904
rect 3557 3864 3569 3904
rect 3577 3864 3589 3904
rect 3681 3864 3693 3943
rect 3701 3864 3713 3943
rect 3731 3864 3743 3944
rect 3817 3864 3829 3904
rect 3837 3864 3849 3904
rect 3857 3864 3869 3904
rect 3956 3864 3968 3904
rect 3978 3864 3990 3944
rect 4006 3864 4018 3944
rect 4091 3864 4103 3944
rect 4111 3864 4123 3944
rect 4131 3864 4143 3932
rect 4151 3864 4163 3936
rect 4217 3864 4229 3904
rect 4237 3864 4249 3904
rect 4257 3864 4269 3904
rect 4342 3864 4354 3944
rect 4370 3864 4382 3944
rect 4392 3864 4404 3904
rect 4482 3864 4494 3944
rect 4510 3864 4522 3944
rect 4532 3864 4544 3904
rect 4617 3864 4629 3944
rect 4647 3864 4659 3943
rect 4667 3864 4679 3943
rect 4771 3864 4783 3904
rect 4791 3864 4803 3904
rect 4811 3864 4823 3904
rect 4877 3864 4889 3904
rect 4897 3864 4909 3904
rect 4917 3864 4929 3900
rect 4937 3864 4949 3904
rect 5017 3864 5029 3904
rect 5037 3864 5049 3904
rect 5131 3864 5143 3904
rect 5151 3864 5163 3904
rect 5177 3864 5189 3944
rect 5197 3864 5209 3884
rect 5227 3864 5239 3884
rect 5255 3864 5267 3904
rect 5281 3864 5293 3904
rect 5301 3864 5313 3904
rect 5333 3864 5345 3904
rect 5367 3864 5379 3904
rect 5387 3864 5399 3944
rect 5417 3864 5429 3944
rect 5437 3864 5449 3884
rect 5467 3864 5479 3884
rect 5495 3864 5507 3904
rect 5521 3864 5533 3904
rect 5541 3864 5553 3904
rect 5573 3864 5585 3904
rect 5607 3864 5619 3904
rect 5627 3864 5639 3944
rect 5702 3864 5714 3944
rect 5730 3864 5742 3944
rect 5752 3864 5764 3904
rect 71 3796 83 3836
rect 91 3796 103 3836
rect 111 3796 123 3836
rect 191 3796 203 3836
rect 211 3800 223 3836
rect 231 3796 243 3836
rect 251 3796 263 3836
rect 327 3768 339 3828
rect 347 3772 359 3824
rect 367 3768 379 3828
rect 391 3778 403 3836
rect 411 3776 423 3824
rect 431 3776 443 3836
rect 451 3776 463 3836
rect 471 3776 483 3836
rect 556 3796 568 3836
rect 578 3756 590 3836
rect 606 3756 618 3836
rect 691 3796 703 3836
rect 711 3796 723 3836
rect 731 3796 743 3836
rect 802 3756 814 3836
rect 830 3756 842 3836
rect 852 3796 864 3836
rect 971 3756 983 3836
rect 991 3756 1003 3824
rect 1011 3758 1023 3836
rect 1031 3770 1043 3836
rect 1051 3758 1063 3836
rect 1117 3796 1129 3836
rect 1137 3796 1149 3836
rect 1157 3796 1169 3836
rect 1237 3796 1249 3836
rect 1257 3796 1269 3836
rect 1277 3800 1289 3836
rect 1297 3796 1309 3836
rect 1377 3764 1389 3836
rect 1397 3768 1409 3836
rect 1417 3756 1429 3836
rect 1437 3756 1449 3836
rect 1522 3756 1534 3836
rect 1550 3756 1562 3836
rect 1572 3796 1584 3836
rect 1657 3796 1669 3836
rect 1677 3796 1689 3836
rect 1771 3796 1783 3836
rect 1791 3796 1803 3836
rect 1811 3796 1823 3836
rect 1877 3796 1889 3836
rect 1897 3796 1909 3836
rect 1917 3796 1929 3836
rect 1997 3756 2009 3836
rect 2027 3757 2039 3836
rect 2047 3757 2059 3836
rect 2137 3796 2149 3836
rect 2157 3796 2169 3836
rect 2177 3796 2189 3836
rect 2257 3796 2269 3836
rect 2277 3796 2289 3836
rect 2297 3800 2309 3836
rect 2317 3796 2329 3836
rect 2416 3796 2428 3836
rect 2438 3756 2450 3836
rect 2466 3756 2478 3836
rect 2537 3796 2549 3836
rect 2557 3796 2569 3836
rect 2577 3796 2589 3836
rect 2662 3756 2674 3836
rect 2690 3756 2702 3836
rect 2712 3796 2724 3836
rect 2811 3796 2823 3836
rect 2831 3796 2843 3836
rect 2916 3796 2928 3836
rect 2938 3756 2950 3836
rect 2966 3756 2978 3836
rect 3037 3796 3049 3836
rect 3057 3796 3069 3836
rect 3077 3796 3089 3836
rect 3191 3796 3203 3836
rect 3211 3796 3223 3836
rect 3231 3796 3243 3836
rect 3311 3796 3323 3836
rect 3331 3796 3343 3836
rect 3397 3796 3409 3836
rect 3417 3796 3429 3836
rect 3437 3800 3449 3836
rect 3457 3796 3469 3836
rect 3537 3796 3549 3836
rect 3557 3796 3569 3836
rect 3663 3756 3675 3836
rect 3691 3756 3703 3836
rect 3777 3796 3789 3836
rect 3797 3796 3809 3836
rect 3817 3796 3829 3836
rect 3897 3796 3909 3836
rect 3917 3796 3929 3836
rect 4011 3796 4023 3836
rect 4031 3796 4043 3836
rect 4057 3756 4069 3836
rect 4077 3816 4089 3836
rect 4107 3816 4119 3836
rect 4135 3796 4147 3836
rect 4161 3796 4173 3836
rect 4181 3796 4193 3836
rect 4213 3796 4225 3836
rect 4247 3796 4259 3836
rect 4267 3756 4279 3836
rect 4361 3756 4373 3836
rect 4391 3756 4413 3836
rect 4431 3756 4443 3836
rect 4497 3796 4509 3836
rect 4517 3796 4529 3836
rect 4537 3796 4549 3836
rect 4617 3756 4629 3836
rect 4645 3756 4657 3836
rect 4742 3756 4754 3836
rect 4770 3756 4782 3836
rect 4792 3796 4804 3836
rect 4877 3756 4889 3836
rect 4897 3756 4909 3836
rect 5011 3796 5023 3836
rect 5031 3796 5043 3836
rect 5051 3796 5063 3836
rect 5117 3796 5129 3836
rect 5137 3796 5149 3836
rect 5231 3756 5243 3836
rect 5251 3756 5263 3836
rect 5271 3756 5283 3836
rect 5291 3756 5303 3836
rect 5311 3756 5323 3836
rect 5331 3756 5343 3836
rect 5351 3756 5363 3836
rect 5371 3756 5383 3836
rect 5391 3756 5403 3836
rect 5417 3756 5429 3836
rect 5437 3816 5449 3836
rect 5467 3816 5479 3836
rect 5495 3796 5507 3836
rect 5521 3796 5533 3836
rect 5541 3796 5553 3836
rect 5573 3796 5585 3836
rect 5607 3796 5619 3836
rect 5627 3756 5639 3836
rect 5711 3796 5723 3836
rect 5731 3796 5743 3836
rect 5751 3796 5763 3836
rect 76 3384 88 3424
rect 98 3384 110 3464
rect 126 3384 138 3464
rect 197 3384 209 3456
rect 217 3384 229 3452
rect 237 3384 249 3464
rect 257 3384 269 3464
rect 337 3384 349 3424
rect 357 3384 369 3424
rect 442 3384 454 3464
rect 470 3384 482 3464
rect 492 3384 504 3424
rect 577 3384 589 3424
rect 597 3384 609 3424
rect 617 3384 629 3420
rect 637 3384 649 3424
rect 751 3384 763 3424
rect 771 3384 783 3424
rect 791 3384 803 3424
rect 871 3384 883 3424
rect 891 3384 903 3424
rect 911 3384 923 3424
rect 982 3384 994 3464
rect 1010 3384 1022 3464
rect 1032 3384 1044 3424
rect 1131 3384 1143 3424
rect 1151 3384 1163 3420
rect 1171 3384 1183 3424
rect 1191 3384 1203 3424
rect 1257 3384 1269 3424
rect 1277 3384 1289 3424
rect 1297 3384 1309 3424
rect 1391 3384 1403 3424
rect 1411 3384 1423 3420
rect 1431 3384 1443 3424
rect 1451 3384 1463 3424
rect 1522 3384 1534 3464
rect 1550 3384 1562 3464
rect 1572 3384 1584 3424
rect 1671 3384 1683 3464
rect 1691 3384 1703 3464
rect 1711 3384 1723 3452
rect 1731 3384 1743 3456
rect 1811 3384 1823 3424
rect 1831 3384 1843 3420
rect 1851 3384 1863 3424
rect 1871 3384 1883 3424
rect 1937 3384 1949 3456
rect 1957 3384 1969 3452
rect 1977 3384 1989 3464
rect 1997 3384 2009 3464
rect 2096 3384 2108 3424
rect 2118 3384 2130 3464
rect 2146 3384 2158 3464
rect 2242 3384 2254 3464
rect 2270 3384 2282 3464
rect 2292 3384 2304 3424
rect 2391 3384 2403 3464
rect 2411 3384 2423 3464
rect 2431 3384 2443 3452
rect 2451 3384 2463 3456
rect 2527 3384 2539 3464
rect 2547 3384 2559 3464
rect 2571 3384 2583 3424
rect 2591 3384 2603 3424
rect 2657 3384 2669 3424
rect 2677 3384 2689 3424
rect 2697 3384 2709 3424
rect 2796 3384 2808 3424
rect 2818 3384 2830 3464
rect 2846 3384 2858 3464
rect 2949 3384 2961 3464
rect 2969 3384 2981 3464
rect 2991 3384 3003 3424
rect 3071 3384 3083 3424
rect 3091 3384 3103 3424
rect 3111 3384 3123 3424
rect 3177 3384 3189 3424
rect 3197 3384 3209 3424
rect 3217 3384 3229 3420
rect 3237 3384 3249 3424
rect 3331 3384 3343 3424
rect 3351 3384 3363 3420
rect 3371 3384 3383 3424
rect 3391 3384 3403 3424
rect 3476 3384 3488 3424
rect 3498 3384 3510 3464
rect 3526 3384 3538 3464
rect 3616 3384 3628 3424
rect 3638 3384 3650 3464
rect 3666 3384 3678 3464
rect 3747 3384 3759 3464
rect 3767 3384 3779 3464
rect 3791 3384 3803 3424
rect 3811 3384 3823 3424
rect 3877 3384 3889 3464
rect 3905 3384 3917 3464
rect 4036 3384 4048 3424
rect 4058 3384 4070 3464
rect 4086 3384 4098 3464
rect 4157 3384 4169 3424
rect 4177 3384 4189 3424
rect 4262 3384 4274 3464
rect 4290 3384 4302 3464
rect 4312 3384 4324 3424
rect 4411 3384 4423 3424
rect 4431 3384 4443 3424
rect 4451 3384 4463 3424
rect 4517 3384 4529 3424
rect 4537 3384 4549 3424
rect 4557 3384 4569 3424
rect 4597 3384 4609 3464
rect 4617 3384 4629 3404
rect 4647 3384 4659 3404
rect 4675 3384 4687 3424
rect 4701 3384 4713 3424
rect 4721 3384 4733 3424
rect 4753 3384 4765 3424
rect 4787 3384 4799 3424
rect 4807 3384 4819 3464
rect 4891 3384 4903 3424
rect 4911 3384 4923 3424
rect 4931 3384 4943 3424
rect 5016 3384 5028 3424
rect 5038 3384 5050 3464
rect 5066 3384 5078 3464
rect 5157 3384 5169 3424
rect 5177 3384 5189 3424
rect 5197 3384 5209 3424
rect 5241 3384 5253 3464
rect 5261 3384 5273 3424
rect 5295 3384 5307 3424
rect 5327 3384 5339 3424
rect 5347 3384 5359 3424
rect 5373 3384 5385 3424
rect 5401 3384 5413 3404
rect 5431 3384 5443 3404
rect 5451 3384 5463 3464
rect 5531 3384 5543 3424
rect 5551 3384 5563 3424
rect 5571 3384 5583 3424
rect 5642 3384 5654 3464
rect 5670 3384 5682 3464
rect 5692 3384 5704 3424
rect 71 3316 83 3356
rect 91 3316 103 3356
rect 176 3316 188 3356
rect 198 3276 210 3356
rect 226 3276 238 3356
rect 311 3316 323 3356
rect 331 3316 343 3356
rect 397 3316 409 3356
rect 417 3316 429 3356
rect 437 3316 449 3356
rect 517 3284 529 3356
rect 537 3288 549 3356
rect 557 3276 569 3356
rect 577 3276 589 3356
rect 657 3316 669 3356
rect 677 3316 689 3356
rect 701 3276 713 3356
rect 721 3276 733 3356
rect 831 3316 843 3356
rect 851 3316 863 3356
rect 871 3316 883 3356
rect 951 3316 963 3356
rect 971 3320 983 3356
rect 991 3316 1003 3356
rect 1011 3316 1023 3356
rect 1091 3316 1103 3356
rect 1111 3320 1123 3356
rect 1131 3316 1143 3356
rect 1151 3316 1163 3356
rect 1217 3284 1229 3356
rect 1237 3288 1249 3356
rect 1257 3276 1269 3356
rect 1277 3276 1289 3356
rect 1371 3316 1383 3356
rect 1391 3316 1403 3356
rect 1471 3316 1483 3356
rect 1491 3320 1503 3356
rect 1511 3316 1523 3356
rect 1531 3316 1543 3356
rect 1611 3316 1623 3356
rect 1631 3320 1643 3356
rect 1651 3316 1663 3356
rect 1671 3316 1683 3356
rect 1751 3276 1763 3356
rect 1771 3276 1783 3356
rect 1791 3288 1803 3356
rect 1811 3284 1823 3356
rect 1911 3316 1923 3356
rect 1931 3316 1943 3356
rect 1951 3316 1963 3356
rect 2031 3276 2043 3356
rect 2051 3276 2063 3356
rect 2071 3288 2083 3356
rect 2091 3284 2103 3356
rect 2157 3316 2169 3356
rect 2177 3316 2189 3356
rect 2197 3316 2209 3356
rect 2287 3276 2299 3356
rect 2307 3276 2319 3356
rect 2331 3316 2343 3356
rect 2351 3316 2363 3356
rect 2417 3316 2429 3356
rect 2437 3316 2449 3356
rect 2457 3316 2469 3356
rect 2556 3316 2568 3356
rect 2578 3276 2590 3356
rect 2606 3276 2618 3356
rect 2691 3276 2703 3356
rect 2711 3276 2723 3356
rect 2731 3288 2743 3356
rect 2751 3284 2763 3356
rect 2817 3316 2829 3356
rect 2837 3316 2849 3356
rect 2857 3320 2869 3356
rect 2877 3316 2889 3356
rect 2957 3316 2969 3356
rect 2977 3316 2989 3356
rect 2997 3320 3009 3356
rect 3017 3316 3029 3356
rect 3111 3316 3123 3356
rect 3131 3316 3143 3356
rect 3151 3316 3163 3356
rect 3251 3316 3263 3356
rect 3271 3316 3283 3356
rect 3291 3316 3303 3356
rect 3357 3316 3369 3356
rect 3377 3316 3389 3356
rect 3471 3316 3483 3356
rect 3491 3320 3503 3356
rect 3511 3316 3523 3356
rect 3531 3316 3543 3356
rect 3597 3284 3609 3356
rect 3617 3288 3629 3356
rect 3637 3276 3649 3356
rect 3657 3276 3669 3356
rect 3756 3316 3768 3356
rect 3778 3276 3790 3356
rect 3806 3276 3818 3356
rect 3877 3316 3889 3356
rect 3897 3316 3909 3356
rect 3937 3276 3949 3356
rect 3957 3336 3969 3356
rect 3987 3336 3999 3356
rect 4015 3316 4027 3356
rect 4041 3316 4053 3356
rect 4061 3316 4073 3356
rect 4093 3316 4105 3356
rect 4127 3316 4139 3356
rect 4147 3276 4159 3356
rect 4222 3276 4234 3356
rect 4250 3276 4262 3356
rect 4272 3316 4284 3356
rect 4362 3276 4374 3356
rect 4390 3276 4402 3356
rect 4412 3316 4424 3356
rect 4457 3276 4469 3356
rect 4477 3336 4489 3356
rect 4507 3336 4519 3356
rect 4535 3316 4547 3356
rect 4561 3316 4573 3356
rect 4581 3316 4593 3356
rect 4613 3316 4625 3356
rect 4647 3316 4659 3356
rect 4667 3276 4679 3356
rect 4742 3276 4754 3356
rect 4770 3276 4782 3356
rect 4792 3316 4804 3356
rect 4891 3316 4903 3356
rect 4911 3316 4923 3356
rect 4931 3316 4943 3356
rect 5016 3316 5028 3356
rect 5038 3276 5050 3356
rect 5066 3276 5078 3356
rect 5151 3316 5163 3356
rect 5171 3316 5183 3356
rect 5251 3316 5263 3356
rect 5271 3316 5283 3356
rect 5291 3316 5303 3356
rect 5357 3316 5369 3356
rect 5377 3316 5389 3356
rect 5482 3276 5494 3356
rect 5510 3276 5522 3356
rect 5532 3316 5544 3356
rect 5651 3316 5663 3356
rect 5671 3316 5683 3356
rect 5691 3316 5703 3356
rect 87 2904 99 2984
rect 107 2904 119 2984
rect 131 2904 143 2944
rect 151 2904 163 2944
rect 237 2904 249 2944
rect 257 2904 269 2944
rect 277 2904 289 2940
rect 297 2904 309 2944
rect 377 2904 389 2944
rect 397 2904 409 2944
rect 417 2904 429 2944
rect 516 2904 528 2944
rect 538 2904 550 2984
rect 566 2904 578 2984
rect 642 2904 654 2984
rect 670 2904 682 2984
rect 692 2904 704 2944
rect 782 2904 794 2984
rect 810 2904 822 2984
rect 832 2904 844 2944
rect 922 2904 934 2984
rect 950 2904 962 2984
rect 972 2904 984 2944
rect 1071 2904 1083 2944
rect 1091 2904 1103 2944
rect 1111 2904 1123 2944
rect 1223 2904 1235 2984
rect 1251 2904 1263 2984
rect 1322 2904 1334 2984
rect 1350 2904 1362 2984
rect 1372 2904 1384 2944
rect 1471 2904 1483 2944
rect 1491 2904 1503 2940
rect 1511 2904 1523 2944
rect 1531 2904 1543 2944
rect 1631 2904 1643 2984
rect 1651 2904 1663 2984
rect 1671 2904 1683 2972
rect 1691 2904 1703 2976
rect 1776 2904 1788 2944
rect 1798 2904 1810 2984
rect 1826 2904 1838 2984
rect 1902 2904 1914 2984
rect 1930 2904 1942 2984
rect 1952 2904 1964 2944
rect 2076 2904 2088 2944
rect 2098 2904 2110 2984
rect 2126 2904 2138 2984
rect 2216 2904 2228 2944
rect 2238 2904 2250 2984
rect 2266 2904 2278 2984
rect 2371 2904 2383 2984
rect 2391 2904 2403 2984
rect 2411 2904 2423 2972
rect 2431 2904 2443 2976
rect 2511 2904 2523 2984
rect 2531 2904 2543 2984
rect 2551 2904 2563 2972
rect 2571 2904 2583 2976
rect 2651 2904 2663 2984
rect 2671 2916 2683 2984
rect 2691 2904 2703 2982
rect 2711 2904 2723 2970
rect 2731 2904 2743 2982
rect 2821 2904 2833 2983
rect 2841 2904 2853 2983
rect 2871 2904 2883 2984
rect 2937 2904 2949 2984
rect 2965 2904 2977 2984
rect 3077 2904 3089 2944
rect 3097 2904 3109 2944
rect 3117 2904 3129 2944
rect 3207 2904 3219 2984
rect 3227 2904 3239 2984
rect 3251 2904 3263 2944
rect 3271 2904 3283 2944
rect 3337 2904 3349 2984
rect 3367 2904 3379 2983
rect 3387 2904 3399 2983
rect 3496 2904 3508 2944
rect 3518 2904 3530 2984
rect 3546 2904 3558 2984
rect 3636 2904 3648 2944
rect 3658 2904 3670 2984
rect 3686 2904 3698 2984
rect 3781 2904 3793 2983
rect 3801 2904 3813 2983
rect 3831 2904 3843 2984
rect 3927 2904 3939 2984
rect 3947 2904 3959 2984
rect 3971 2904 3983 2944
rect 3991 2904 4003 2944
rect 4057 2904 4069 2984
rect 4085 2904 4097 2984
rect 4177 2904 4189 2944
rect 4197 2904 4209 2944
rect 4217 2904 4229 2940
rect 4237 2904 4249 2944
rect 4281 2904 4293 2984
rect 4301 2904 4313 2944
rect 4335 2904 4347 2944
rect 4367 2904 4379 2944
rect 4387 2904 4399 2944
rect 4413 2904 4425 2944
rect 4441 2904 4453 2924
rect 4471 2904 4483 2924
rect 4491 2904 4503 2984
rect 4582 2904 4594 2984
rect 4610 2904 4622 2984
rect 4632 2904 4644 2944
rect 4722 2904 4734 2984
rect 4750 2904 4762 2984
rect 4772 2904 4784 2944
rect 4871 2904 4883 2944
rect 4891 2904 4903 2944
rect 4911 2904 4923 2944
rect 4977 2904 4989 2944
rect 4997 2904 5009 2944
rect 5017 2904 5029 2944
rect 5061 2904 5073 2984
rect 5081 2904 5093 2944
rect 5115 2904 5127 2944
rect 5147 2904 5159 2944
rect 5167 2904 5179 2944
rect 5193 2904 5205 2944
rect 5221 2904 5233 2924
rect 5251 2904 5263 2924
rect 5271 2904 5283 2984
rect 5351 2904 5363 2984
rect 5371 2904 5383 2984
rect 5391 2904 5403 2984
rect 5411 2904 5423 2984
rect 5431 2904 5443 2984
rect 5451 2904 5463 2984
rect 5471 2904 5483 2984
rect 5491 2904 5503 2984
rect 5511 2904 5523 2984
rect 5537 2904 5549 2984
rect 5557 2904 5569 2924
rect 5587 2904 5599 2924
rect 5615 2904 5627 2944
rect 5641 2904 5653 2944
rect 5661 2904 5673 2944
rect 5693 2904 5705 2944
rect 5727 2904 5739 2944
rect 5747 2904 5759 2984
rect 71 2836 83 2876
rect 91 2836 103 2876
rect 111 2836 123 2876
rect 182 2796 194 2876
rect 210 2796 222 2876
rect 232 2836 244 2876
rect 331 2836 343 2876
rect 351 2836 363 2876
rect 417 2804 429 2876
rect 437 2808 449 2876
rect 457 2796 469 2876
rect 477 2796 489 2876
rect 571 2836 583 2876
rect 591 2836 603 2876
rect 611 2836 623 2876
rect 677 2836 689 2876
rect 697 2836 709 2876
rect 721 2796 733 2876
rect 741 2796 753 2876
rect 817 2836 829 2876
rect 837 2836 849 2876
rect 857 2836 869 2876
rect 937 2804 949 2876
rect 957 2808 969 2876
rect 977 2796 989 2876
rect 997 2796 1009 2876
rect 1077 2836 1089 2876
rect 1097 2836 1109 2876
rect 1117 2836 1129 2876
rect 1236 2836 1248 2876
rect 1258 2796 1270 2876
rect 1286 2796 1298 2876
rect 1362 2796 1374 2876
rect 1390 2796 1402 2876
rect 1412 2836 1424 2876
rect 1521 2797 1533 2876
rect 1541 2797 1553 2876
rect 1571 2796 1583 2876
rect 1637 2796 1649 2876
rect 1665 2796 1677 2876
rect 1767 2796 1779 2876
rect 1787 2796 1799 2876
rect 1811 2836 1823 2876
rect 1831 2836 1843 2876
rect 1931 2836 1943 2876
rect 1951 2836 1963 2876
rect 1971 2836 1983 2876
rect 2042 2796 2054 2876
rect 2070 2796 2082 2876
rect 2092 2836 2104 2876
rect 2187 2796 2199 2876
rect 2207 2796 2219 2876
rect 2231 2836 2243 2876
rect 2251 2836 2263 2876
rect 2331 2836 2343 2876
rect 2351 2836 2363 2876
rect 2371 2836 2383 2876
rect 2457 2796 2469 2876
rect 2485 2796 2497 2876
rect 2591 2836 2603 2876
rect 2611 2840 2623 2876
rect 2631 2836 2643 2876
rect 2651 2836 2663 2876
rect 2727 2796 2739 2876
rect 2747 2796 2759 2876
rect 2771 2836 2783 2876
rect 2791 2836 2803 2876
rect 2882 2796 2894 2876
rect 2910 2796 2922 2876
rect 2932 2836 2944 2876
rect 3031 2836 3043 2876
rect 3051 2840 3063 2876
rect 3071 2836 3083 2876
rect 3091 2836 3103 2876
rect 3157 2836 3169 2876
rect 3177 2836 3189 2876
rect 3197 2836 3209 2876
rect 3296 2836 3308 2876
rect 3318 2796 3330 2876
rect 3346 2796 3358 2876
rect 3427 2796 3439 2876
rect 3447 2796 3459 2876
rect 3471 2836 3483 2876
rect 3491 2836 3503 2876
rect 3557 2796 3569 2876
rect 3585 2796 3597 2876
rect 3677 2836 3689 2876
rect 3697 2836 3709 2876
rect 3717 2840 3729 2876
rect 3737 2836 3749 2876
rect 3817 2836 3829 2876
rect 3837 2836 3849 2876
rect 3857 2836 3869 2876
rect 3951 2796 3963 2876
rect 3971 2796 3983 2876
rect 4056 2836 4068 2876
rect 4078 2796 4090 2876
rect 4106 2796 4118 2876
rect 4177 2836 4189 2876
rect 4197 2836 4209 2876
rect 4217 2836 4229 2876
rect 4297 2796 4309 2876
rect 4317 2796 4329 2876
rect 4397 2836 4409 2876
rect 4417 2836 4429 2876
rect 4457 2796 4469 2876
rect 4477 2856 4489 2876
rect 4507 2856 4519 2876
rect 4535 2836 4547 2876
rect 4561 2836 4573 2876
rect 4581 2836 4593 2876
rect 4613 2836 4625 2876
rect 4647 2836 4659 2876
rect 4667 2796 4679 2876
rect 4701 2796 4713 2876
rect 4721 2836 4733 2876
rect 4755 2836 4767 2876
rect 4787 2836 4799 2876
rect 4807 2836 4819 2876
rect 4833 2836 4845 2876
rect 4861 2856 4873 2876
rect 4891 2856 4903 2876
rect 4911 2796 4923 2876
rect 5002 2796 5014 2876
rect 5030 2796 5042 2876
rect 5052 2836 5064 2876
rect 5137 2836 5149 2876
rect 5157 2836 5169 2876
rect 5177 2836 5189 2876
rect 5257 2796 5269 2874
rect 5277 2796 5289 2876
rect 5297 2796 5309 2876
rect 5337 2796 5349 2876
rect 5357 2856 5369 2876
rect 5387 2856 5399 2876
rect 5415 2836 5427 2876
rect 5441 2836 5453 2876
rect 5461 2836 5473 2876
rect 5493 2836 5505 2876
rect 5527 2836 5539 2876
rect 5547 2796 5559 2876
rect 5622 2796 5634 2876
rect 5650 2796 5662 2876
rect 5672 2836 5684 2876
rect 71 2424 83 2464
rect 91 2424 103 2464
rect 157 2424 169 2464
rect 177 2424 189 2464
rect 271 2424 283 2504
rect 291 2424 303 2504
rect 311 2424 323 2492
rect 331 2424 343 2496
rect 397 2424 409 2464
rect 417 2424 429 2464
rect 437 2424 449 2460
rect 457 2424 469 2464
rect 537 2424 549 2464
rect 557 2424 569 2464
rect 637 2424 649 2504
rect 665 2424 677 2504
rect 762 2424 774 2504
rect 790 2424 802 2504
rect 812 2424 824 2464
rect 917 2424 929 2496
rect 937 2424 949 2492
rect 957 2424 969 2504
rect 977 2424 989 2504
rect 1076 2424 1088 2464
rect 1098 2424 1110 2504
rect 1126 2424 1138 2504
rect 1211 2424 1223 2464
rect 1231 2424 1243 2464
rect 1251 2424 1263 2464
rect 1317 2424 1329 2464
rect 1337 2424 1349 2464
rect 1361 2424 1373 2504
rect 1381 2424 1393 2504
rect 1471 2424 1483 2464
rect 1491 2424 1503 2460
rect 1511 2424 1523 2464
rect 1531 2424 1543 2464
rect 1597 2424 1609 2464
rect 1617 2424 1629 2464
rect 1702 2424 1714 2504
rect 1730 2424 1742 2504
rect 1752 2424 1764 2464
rect 1856 2424 1868 2464
rect 1878 2424 1890 2504
rect 1906 2424 1918 2504
rect 1982 2424 1994 2504
rect 2010 2424 2022 2504
rect 2032 2424 2044 2464
rect 2131 2424 2143 2464
rect 2151 2424 2163 2460
rect 2171 2424 2183 2464
rect 2191 2424 2203 2464
rect 2271 2424 2283 2504
rect 2291 2424 2303 2504
rect 2311 2424 2323 2492
rect 2331 2424 2343 2496
rect 2397 2424 2409 2464
rect 2417 2424 2429 2464
rect 2437 2424 2449 2464
rect 2556 2424 2568 2464
rect 2578 2424 2590 2504
rect 2606 2424 2618 2504
rect 2682 2424 2694 2504
rect 2710 2424 2722 2504
rect 2732 2424 2744 2464
rect 2831 2424 2843 2504
rect 2851 2424 2863 2504
rect 2871 2424 2883 2492
rect 2891 2424 2903 2496
rect 2971 2424 2983 2464
rect 2991 2424 3003 2464
rect 3062 2424 3074 2504
rect 3090 2424 3102 2504
rect 3112 2424 3124 2464
rect 3217 2424 3229 2464
rect 3237 2424 3249 2464
rect 3257 2424 3269 2464
rect 3351 2424 3363 2464
rect 3371 2424 3383 2460
rect 3391 2424 3403 2464
rect 3411 2424 3423 2464
rect 3477 2424 3489 2464
rect 3497 2424 3509 2464
rect 3521 2424 3533 2504
rect 3541 2424 3553 2504
rect 3617 2424 3629 2464
rect 3637 2424 3649 2464
rect 3657 2424 3669 2464
rect 3737 2424 3749 2502
rect 3757 2424 3769 2490
rect 3777 2424 3789 2502
rect 3797 2436 3809 2504
rect 3817 2424 3829 2504
rect 3897 2424 3909 2504
rect 3925 2424 3937 2504
rect 3985 2424 3997 2464
rect 4005 2424 4017 2464
rect 4030 2424 4042 2464
rect 4050 2424 4062 2464
rect 4070 2424 4082 2464
rect 4090 2424 4102 2464
rect 4110 2424 4122 2464
rect 4135 2424 4147 2444
rect 4155 2424 4167 2444
rect 4175 2424 4187 2444
rect 4200 2424 4212 2464
rect 4220 2424 4232 2464
rect 4240 2424 4252 2464
rect 4265 2424 4277 2464
rect 4285 2424 4297 2444
rect 4305 2424 4317 2444
rect 4325 2424 4337 2444
rect 4350 2424 4362 2447
rect 4370 2424 4382 2464
rect 4390 2424 4402 2464
rect 4410 2424 4422 2464
rect 4430 2424 4442 2464
rect 4458 2424 4470 2464
rect 4478 2424 4490 2464
rect 4498 2424 4510 2464
rect 4518 2424 4530 2464
rect 4538 2424 4550 2447
rect 4563 2424 4575 2444
rect 4583 2424 4595 2444
rect 4603 2424 4615 2444
rect 4623 2424 4635 2464
rect 4648 2424 4660 2464
rect 4668 2424 4680 2464
rect 4688 2424 4700 2464
rect 4713 2424 4725 2444
rect 4733 2424 4745 2444
rect 4753 2424 4765 2444
rect 4778 2424 4790 2464
rect 4798 2424 4810 2464
rect 4818 2424 4830 2464
rect 4838 2424 4850 2464
rect 4858 2424 4870 2464
rect 4883 2424 4895 2464
rect 4903 2424 4915 2464
rect 4941 2424 4953 2504
rect 4961 2424 4973 2464
rect 4995 2424 5007 2464
rect 5027 2424 5039 2464
rect 5047 2424 5059 2464
rect 5073 2424 5085 2464
rect 5101 2424 5113 2444
rect 5131 2424 5143 2444
rect 5151 2424 5163 2504
rect 5231 2424 5243 2504
rect 5251 2424 5263 2504
rect 5271 2424 5283 2504
rect 5291 2424 5303 2504
rect 5311 2424 5323 2504
rect 5331 2424 5343 2504
rect 5351 2424 5363 2504
rect 5371 2424 5383 2504
rect 5391 2424 5403 2504
rect 5477 2424 5489 2504
rect 5497 2424 5509 2504
rect 5517 2424 5529 2504
rect 5537 2424 5549 2504
rect 5557 2424 5569 2504
rect 5577 2424 5589 2504
rect 5597 2424 5609 2504
rect 5617 2424 5629 2504
rect 5637 2424 5649 2504
rect 5717 2424 5729 2504
rect 5737 2424 5749 2504
rect 69 2316 81 2396
rect 89 2316 101 2396
rect 111 2356 123 2396
rect 191 2356 203 2396
rect 211 2360 223 2396
rect 231 2356 243 2396
rect 251 2356 263 2396
rect 317 2356 329 2396
rect 337 2356 349 2396
rect 357 2356 369 2396
rect 442 2316 454 2396
rect 470 2316 482 2396
rect 492 2356 504 2396
rect 596 2356 608 2396
rect 618 2316 630 2396
rect 646 2316 658 2396
rect 751 2356 763 2396
rect 771 2360 783 2396
rect 791 2356 803 2396
rect 811 2356 823 2396
rect 891 2356 903 2396
rect 911 2356 923 2396
rect 931 2356 943 2396
rect 1021 2317 1033 2396
rect 1041 2317 1053 2396
rect 1071 2316 1083 2396
rect 1137 2316 1149 2396
rect 1157 2316 1169 2396
rect 1251 2356 1263 2396
rect 1271 2360 1283 2396
rect 1291 2356 1303 2396
rect 1311 2356 1323 2396
rect 1391 2316 1403 2396
rect 1411 2316 1423 2396
rect 1431 2328 1443 2396
rect 1451 2324 1463 2396
rect 1556 2356 1568 2396
rect 1578 2316 1590 2396
rect 1606 2316 1618 2396
rect 1691 2316 1703 2396
rect 1711 2316 1723 2396
rect 1731 2328 1743 2396
rect 1751 2324 1763 2396
rect 1831 2356 1843 2396
rect 1851 2360 1863 2396
rect 1871 2356 1883 2396
rect 1891 2356 1903 2396
rect 1971 2356 1983 2396
rect 1991 2360 2003 2396
rect 2011 2356 2023 2396
rect 2031 2356 2043 2396
rect 2065 2356 2077 2396
rect 2085 2356 2097 2396
rect 2110 2356 2122 2396
rect 2130 2356 2142 2396
rect 2150 2356 2162 2396
rect 2170 2356 2182 2396
rect 2190 2356 2202 2396
rect 2215 2376 2227 2396
rect 2235 2376 2247 2396
rect 2255 2376 2267 2396
rect 2280 2356 2292 2396
rect 2300 2356 2312 2396
rect 2320 2356 2332 2396
rect 2345 2356 2357 2396
rect 2365 2376 2377 2396
rect 2385 2376 2397 2396
rect 2405 2376 2417 2396
rect 2430 2373 2442 2396
rect 2450 2356 2462 2396
rect 2470 2356 2482 2396
rect 2490 2356 2502 2396
rect 2510 2356 2522 2396
rect 2589 2316 2601 2396
rect 2609 2316 2621 2396
rect 2631 2356 2643 2396
rect 2722 2316 2734 2396
rect 2750 2316 2762 2396
rect 2772 2356 2784 2396
rect 2862 2316 2874 2396
rect 2890 2316 2902 2396
rect 2912 2356 2924 2396
rect 3011 2356 3023 2396
rect 3031 2356 3043 2396
rect 3051 2356 3063 2396
rect 3137 2356 3149 2396
rect 3157 2356 3169 2396
rect 3177 2356 3189 2396
rect 3271 2316 3283 2396
rect 3291 2316 3303 2396
rect 3311 2328 3323 2396
rect 3331 2324 3343 2396
rect 3397 2316 3409 2396
rect 3425 2316 3437 2396
rect 3542 2316 3554 2396
rect 3570 2316 3582 2396
rect 3592 2356 3604 2396
rect 3677 2356 3689 2396
rect 3697 2356 3709 2396
rect 3717 2356 3729 2396
rect 3797 2356 3809 2396
rect 3819 2316 3831 2396
rect 3839 2316 3851 2396
rect 3885 2356 3897 2396
rect 3905 2356 3917 2396
rect 3930 2356 3942 2396
rect 3950 2356 3962 2396
rect 3970 2356 3982 2396
rect 3990 2356 4002 2396
rect 4010 2356 4022 2396
rect 4035 2376 4047 2396
rect 4055 2376 4067 2396
rect 4075 2376 4087 2396
rect 4100 2356 4112 2396
rect 4120 2356 4132 2396
rect 4140 2356 4152 2396
rect 4165 2356 4177 2396
rect 4185 2376 4197 2396
rect 4205 2376 4217 2396
rect 4225 2376 4237 2396
rect 4250 2373 4262 2396
rect 4270 2356 4282 2396
rect 4290 2356 4302 2396
rect 4310 2356 4322 2396
rect 4330 2356 4342 2396
rect 4397 2356 4409 2396
rect 4417 2356 4429 2396
rect 4441 2316 4453 2396
rect 4461 2316 4473 2396
rect 4537 2318 4549 2396
rect 4557 2330 4569 2396
rect 4577 2318 4589 2396
rect 4597 2316 4609 2384
rect 4617 2316 4629 2396
rect 4697 2356 4709 2396
rect 4717 2356 4729 2396
rect 4737 2356 4749 2396
rect 4829 2316 4841 2396
rect 4849 2316 4861 2396
rect 4871 2356 4883 2396
rect 4937 2356 4949 2396
rect 4957 2356 4969 2396
rect 5037 2318 5049 2396
rect 5057 2330 5069 2396
rect 5077 2318 5089 2396
rect 5097 2316 5109 2384
rect 5117 2316 5129 2396
rect 5197 2356 5209 2396
rect 5217 2356 5229 2396
rect 5237 2356 5249 2396
rect 5317 2316 5329 2396
rect 5337 2316 5349 2396
rect 5417 2356 5429 2396
rect 5437 2356 5449 2396
rect 5457 2356 5469 2396
rect 5537 2356 5549 2396
rect 5557 2356 5569 2396
rect 5637 2348 5649 2388
rect 5657 2348 5669 2388
rect 5687 2324 5699 2388
rect 5717 2316 5729 2396
rect 89 1944 101 2024
rect 109 1944 121 2024
rect 131 1944 143 1984
rect 231 1944 243 1984
rect 251 1944 263 1980
rect 271 1944 283 1984
rect 291 1944 303 1984
rect 357 1944 369 2016
rect 377 1944 389 2012
rect 397 1944 409 2024
rect 417 1944 429 2024
rect 511 1944 523 1984
rect 531 1944 543 1984
rect 616 1944 628 1984
rect 638 1944 650 2024
rect 666 1944 678 2024
rect 751 1944 763 2024
rect 771 1944 783 2024
rect 791 1944 803 2012
rect 811 1944 823 2016
rect 877 1944 889 1984
rect 897 1944 909 1984
rect 917 1944 929 1980
rect 937 1944 949 1984
rect 1051 1944 1063 1984
rect 1071 1944 1083 1980
rect 1091 1944 1103 1984
rect 1111 1944 1123 1984
rect 1196 1944 1208 1984
rect 1218 1944 1230 2024
rect 1246 1944 1258 2024
rect 1336 1944 1348 1984
rect 1358 1944 1370 2024
rect 1386 1944 1398 2024
rect 1471 1944 1483 2024
rect 1491 1944 1503 2024
rect 1511 1944 1523 2012
rect 1531 1944 1543 2016
rect 1611 1944 1623 1984
rect 1631 1944 1643 1980
rect 1651 1944 1663 1984
rect 1671 1944 1683 1984
rect 1742 1944 1754 2024
rect 1770 1944 1782 2024
rect 1792 1944 1804 1984
rect 1877 1944 1889 2016
rect 1897 1944 1909 2012
rect 1917 1944 1929 2024
rect 1937 1944 1949 2024
rect 2027 1952 2039 2012
rect 2047 1956 2059 2008
rect 2067 1952 2079 2012
rect 2091 1944 2103 2002
rect 2111 1956 2123 2004
rect 2131 1944 2143 2004
rect 2151 1944 2163 2004
rect 2171 1944 2183 2004
rect 2251 1944 2263 1984
rect 2271 1944 2283 1980
rect 2291 1944 2303 1984
rect 2311 1944 2323 1984
rect 2345 1944 2357 1984
rect 2365 1944 2377 1984
rect 2390 1944 2402 1984
rect 2410 1944 2422 1984
rect 2430 1944 2442 1984
rect 2450 1944 2462 1984
rect 2470 1944 2482 1984
rect 2495 1944 2507 1964
rect 2515 1944 2527 1964
rect 2535 1944 2547 1964
rect 2560 1944 2572 1984
rect 2580 1944 2592 1984
rect 2600 1944 2612 1984
rect 2625 1944 2637 1984
rect 2645 1944 2657 1964
rect 2665 1944 2677 1964
rect 2685 1944 2697 1964
rect 2710 1944 2722 1967
rect 2730 1944 2742 1984
rect 2750 1944 2762 1984
rect 2770 1944 2782 1984
rect 2790 1944 2802 1984
rect 2862 1944 2874 2024
rect 2890 1944 2902 2024
rect 2912 1944 2924 1984
rect 3011 1944 3023 1984
rect 3031 1944 3043 1984
rect 3051 1944 3063 1984
rect 3117 1944 3129 1984
rect 3137 1944 3149 1984
rect 3157 1944 3169 1984
rect 3257 1944 3269 2024
rect 3285 1944 3297 2024
rect 3387 1944 3399 2024
rect 3407 1944 3419 2024
rect 3431 1944 3443 1984
rect 3451 1944 3463 1984
rect 3517 1944 3529 2016
rect 3537 1944 3549 2012
rect 3557 1944 3569 2024
rect 3577 1944 3589 2024
rect 3691 1944 3703 2024
rect 3711 1944 3723 2024
rect 3797 1944 3809 1984
rect 3817 1944 3829 1984
rect 3837 1944 3849 1980
rect 3857 1944 3869 1984
rect 3957 1944 3969 2024
rect 3977 1944 3989 2024
rect 4087 1944 4099 2024
rect 4107 1944 4119 2024
rect 4131 1944 4143 1984
rect 4151 1944 4163 1984
rect 4231 1944 4243 1984
rect 4251 1944 4263 1984
rect 4271 1944 4283 1984
rect 4356 1944 4368 1984
rect 4378 1944 4390 2024
rect 4406 1944 4418 2024
rect 4482 1944 4494 2024
rect 4510 1944 4522 2024
rect 4532 1944 4544 1984
rect 4617 1944 4629 1984
rect 4637 1944 4649 1984
rect 4657 1944 4669 1984
rect 4737 1944 4749 1984
rect 4757 1944 4769 1984
rect 4777 1944 4789 1984
rect 4896 1944 4908 1984
rect 4918 1944 4930 2024
rect 4946 1944 4958 2024
rect 5036 1944 5048 1984
rect 5058 1944 5070 2024
rect 5086 1944 5098 2024
rect 5157 1944 5169 1984
rect 5177 1944 5189 1984
rect 5257 1944 5269 2024
rect 5285 1944 5297 2024
rect 5377 1944 5389 1984
rect 5397 1944 5409 1984
rect 5417 1944 5429 1984
rect 5497 1944 5509 1984
rect 5517 1944 5529 1984
rect 5611 1944 5623 1984
rect 5631 1944 5643 1984
rect 5702 1944 5714 2024
rect 5730 1944 5742 2024
rect 5752 1944 5764 1984
rect 71 1876 83 1916
rect 91 1880 103 1916
rect 111 1876 123 1916
rect 131 1876 143 1916
rect 197 1844 209 1916
rect 217 1848 229 1916
rect 237 1836 249 1916
rect 257 1836 269 1916
rect 356 1876 368 1916
rect 378 1836 390 1916
rect 406 1836 418 1916
rect 491 1876 503 1916
rect 511 1880 523 1916
rect 531 1876 543 1916
rect 551 1876 563 1916
rect 663 1836 675 1916
rect 691 1836 703 1916
rect 757 1844 769 1916
rect 777 1848 789 1916
rect 797 1836 809 1916
rect 817 1836 829 1916
rect 931 1876 943 1916
rect 951 1876 963 1916
rect 1056 1876 1068 1916
rect 1078 1836 1090 1916
rect 1106 1836 1118 1916
rect 1196 1876 1208 1916
rect 1218 1836 1230 1916
rect 1246 1836 1258 1916
rect 1331 1876 1343 1916
rect 1351 1876 1363 1916
rect 1436 1876 1448 1916
rect 1458 1836 1470 1916
rect 1486 1836 1498 1916
rect 1562 1836 1574 1916
rect 1590 1836 1602 1916
rect 1612 1876 1624 1916
rect 1716 1876 1728 1916
rect 1738 1836 1750 1916
rect 1766 1836 1778 1916
rect 1851 1876 1863 1916
rect 1871 1876 1883 1916
rect 1891 1876 1903 1916
rect 1971 1876 1983 1916
rect 1991 1876 2003 1916
rect 2011 1876 2023 1916
rect 2111 1836 2123 1916
rect 2131 1836 2143 1916
rect 2151 1836 2163 1914
rect 2185 1876 2197 1916
rect 2205 1876 2217 1916
rect 2230 1876 2242 1916
rect 2250 1876 2262 1916
rect 2270 1876 2282 1916
rect 2290 1876 2302 1916
rect 2310 1876 2322 1916
rect 2335 1896 2347 1916
rect 2355 1896 2367 1916
rect 2375 1896 2387 1916
rect 2400 1876 2412 1916
rect 2420 1876 2432 1916
rect 2440 1876 2452 1916
rect 2465 1876 2477 1916
rect 2485 1896 2497 1916
rect 2505 1896 2517 1916
rect 2525 1896 2537 1916
rect 2550 1893 2562 1916
rect 2570 1876 2582 1916
rect 2590 1876 2602 1916
rect 2610 1876 2622 1916
rect 2630 1876 2642 1916
rect 2697 1876 2709 1916
rect 2717 1876 2729 1916
rect 2737 1876 2749 1916
rect 2831 1876 2843 1916
rect 2851 1880 2863 1916
rect 2871 1876 2883 1916
rect 2891 1876 2903 1916
rect 2976 1876 2988 1916
rect 2998 1836 3010 1916
rect 3026 1836 3038 1916
rect 3097 1836 3109 1916
rect 3125 1836 3137 1916
rect 3217 1868 3229 1908
rect 3237 1868 3249 1908
rect 3267 1844 3279 1908
rect 3297 1836 3309 1916
rect 3391 1876 3403 1916
rect 3411 1876 3423 1916
rect 3477 1836 3489 1916
rect 3507 1836 3529 1916
rect 3547 1836 3559 1916
rect 3656 1876 3668 1916
rect 3678 1836 3690 1916
rect 3706 1836 3718 1916
rect 3816 1876 3828 1916
rect 3838 1836 3850 1916
rect 3866 1836 3878 1916
rect 3942 1836 3954 1916
rect 3970 1836 3982 1916
rect 3992 1876 4004 1916
rect 4091 1876 4103 1916
rect 4111 1876 4123 1916
rect 4131 1876 4143 1916
rect 4211 1836 4223 1916
rect 4231 1836 4243 1904
rect 4251 1838 4263 1916
rect 4271 1850 4283 1916
rect 4291 1838 4303 1916
rect 4371 1876 4383 1916
rect 4391 1876 4403 1916
rect 4411 1876 4423 1916
rect 4482 1836 4494 1916
rect 4510 1836 4522 1916
rect 4532 1876 4544 1916
rect 4627 1836 4639 1916
rect 4647 1836 4659 1916
rect 4671 1876 4683 1916
rect 4691 1876 4703 1916
rect 4783 1836 4795 1916
rect 4811 1836 4823 1916
rect 4891 1876 4903 1916
rect 4911 1876 4923 1916
rect 4931 1876 4943 1916
rect 5011 1836 5023 1916
rect 5031 1836 5043 1904
rect 5051 1838 5063 1916
rect 5071 1850 5083 1916
rect 5091 1838 5103 1916
rect 5171 1876 5183 1916
rect 5191 1876 5203 1916
rect 5283 1836 5295 1916
rect 5311 1836 5323 1916
rect 5382 1836 5394 1916
rect 5410 1836 5422 1916
rect 5432 1876 5444 1916
rect 5536 1876 5548 1916
rect 5558 1836 5570 1916
rect 5586 1836 5598 1916
rect 5657 1836 5669 1914
rect 5677 1836 5689 1916
rect 5697 1836 5709 1916
rect 77 1464 89 1504
rect 97 1464 109 1504
rect 117 1464 129 1500
rect 137 1464 149 1504
rect 231 1464 243 1504
rect 251 1464 263 1500
rect 271 1464 283 1504
rect 291 1464 303 1504
rect 357 1464 369 1536
rect 377 1464 389 1532
rect 397 1464 409 1544
rect 417 1464 429 1544
rect 511 1464 523 1544
rect 531 1464 543 1544
rect 551 1464 563 1532
rect 571 1464 583 1536
rect 637 1464 649 1504
rect 657 1464 669 1504
rect 677 1464 689 1504
rect 757 1464 769 1504
rect 777 1464 789 1504
rect 876 1464 888 1504
rect 898 1464 910 1544
rect 926 1464 938 1544
rect 1011 1464 1023 1504
rect 1031 1464 1043 1500
rect 1051 1464 1063 1504
rect 1071 1464 1083 1504
rect 1151 1464 1163 1504
rect 1171 1464 1183 1504
rect 1191 1464 1203 1504
rect 1277 1464 1289 1544
rect 1305 1464 1317 1544
rect 1409 1464 1421 1544
rect 1429 1464 1441 1544
rect 1451 1464 1463 1504
rect 1551 1464 1563 1504
rect 1571 1464 1583 1504
rect 1637 1464 1649 1542
rect 1657 1464 1669 1530
rect 1677 1464 1689 1542
rect 1697 1476 1709 1544
rect 1717 1464 1729 1544
rect 1765 1464 1777 1504
rect 1785 1464 1797 1504
rect 1810 1464 1822 1504
rect 1830 1464 1842 1504
rect 1850 1464 1862 1504
rect 1870 1464 1882 1504
rect 1890 1464 1902 1504
rect 1915 1464 1927 1484
rect 1935 1464 1947 1484
rect 1955 1464 1967 1484
rect 1980 1464 1992 1504
rect 2000 1464 2012 1504
rect 2020 1464 2032 1504
rect 2045 1464 2057 1504
rect 2065 1464 2077 1484
rect 2085 1464 2097 1484
rect 2105 1464 2117 1484
rect 2130 1464 2142 1487
rect 2150 1464 2162 1504
rect 2170 1464 2182 1504
rect 2190 1464 2202 1504
rect 2210 1464 2222 1504
rect 2302 1464 2314 1544
rect 2330 1464 2342 1544
rect 2352 1464 2364 1504
rect 2437 1464 2449 1504
rect 2457 1464 2469 1504
rect 2477 1464 2489 1504
rect 2576 1464 2588 1504
rect 2598 1464 2610 1544
rect 2626 1464 2638 1544
rect 2711 1464 2723 1504
rect 2731 1464 2743 1504
rect 2751 1464 2763 1504
rect 2836 1464 2848 1504
rect 2858 1464 2870 1544
rect 2886 1464 2898 1544
rect 2976 1464 2988 1504
rect 2998 1464 3010 1544
rect 3026 1464 3038 1544
rect 3058 1464 3070 1504
rect 3078 1464 3090 1504
rect 3098 1464 3110 1504
rect 3118 1464 3130 1504
rect 3138 1464 3150 1487
rect 3163 1464 3175 1484
rect 3183 1464 3195 1484
rect 3203 1464 3215 1484
rect 3223 1464 3235 1504
rect 3248 1464 3260 1504
rect 3268 1464 3280 1504
rect 3288 1464 3300 1504
rect 3313 1464 3325 1484
rect 3333 1464 3345 1484
rect 3353 1464 3365 1484
rect 3378 1464 3390 1504
rect 3398 1464 3410 1504
rect 3418 1464 3430 1504
rect 3438 1464 3450 1504
rect 3458 1464 3470 1504
rect 3483 1464 3495 1504
rect 3503 1464 3515 1504
rect 3591 1464 3603 1544
rect 3611 1464 3623 1544
rect 3631 1464 3643 1532
rect 3651 1464 3663 1536
rect 3722 1464 3734 1544
rect 3750 1464 3762 1544
rect 3772 1464 3784 1504
rect 3869 1464 3881 1544
rect 3889 1464 3901 1544
rect 3911 1464 3923 1504
rect 3987 1464 3999 1544
rect 4007 1464 4019 1544
rect 4031 1464 4043 1504
rect 4051 1464 4063 1504
rect 4117 1464 4129 1504
rect 4137 1464 4149 1504
rect 4157 1464 4169 1504
rect 4251 1464 4263 1544
rect 4271 1476 4283 1544
rect 4291 1464 4303 1542
rect 4311 1464 4323 1530
rect 4331 1464 4343 1542
rect 4411 1464 4423 1544
rect 4431 1476 4443 1544
rect 4451 1464 4463 1542
rect 4471 1464 4483 1530
rect 4491 1464 4503 1542
rect 4577 1464 4589 1542
rect 4597 1464 4609 1530
rect 4617 1464 4629 1542
rect 4637 1476 4649 1544
rect 4657 1464 4669 1544
rect 4737 1464 4749 1504
rect 4757 1464 4769 1504
rect 4777 1464 4789 1504
rect 4862 1464 4874 1544
rect 4890 1464 4902 1544
rect 4912 1464 4924 1504
rect 5007 1464 5019 1544
rect 5027 1464 5039 1544
rect 5051 1464 5063 1504
rect 5071 1464 5083 1504
rect 5157 1464 5169 1504
rect 5177 1464 5189 1504
rect 5197 1464 5209 1500
rect 5217 1464 5229 1504
rect 5297 1464 5309 1542
rect 5317 1464 5329 1530
rect 5337 1464 5349 1542
rect 5357 1476 5369 1544
rect 5377 1464 5389 1544
rect 5457 1464 5469 1504
rect 5477 1464 5489 1504
rect 5497 1464 5509 1504
rect 5577 1464 5589 1504
rect 5597 1464 5609 1504
rect 5617 1464 5629 1500
rect 5637 1464 5649 1504
rect 5751 1464 5763 1544
rect 5771 1464 5783 1544
rect 71 1396 83 1436
rect 91 1400 103 1436
rect 111 1396 123 1436
rect 131 1396 143 1436
rect 197 1364 209 1436
rect 217 1368 229 1436
rect 237 1356 249 1436
rect 257 1356 269 1436
rect 351 1396 363 1436
rect 371 1400 383 1436
rect 391 1396 403 1436
rect 411 1396 423 1436
rect 496 1396 508 1436
rect 518 1356 530 1436
rect 546 1356 558 1436
rect 636 1396 648 1436
rect 658 1356 670 1436
rect 686 1356 698 1436
rect 787 1356 799 1436
rect 807 1356 819 1436
rect 831 1396 843 1436
rect 851 1396 863 1436
rect 917 1396 929 1436
rect 937 1396 949 1436
rect 957 1396 969 1436
rect 1051 1396 1063 1436
rect 1071 1396 1083 1436
rect 1137 1396 1149 1436
rect 1157 1396 1169 1436
rect 1177 1400 1189 1436
rect 1197 1396 1209 1436
rect 1277 1396 1289 1436
rect 1297 1396 1309 1436
rect 1317 1396 1329 1436
rect 1411 1396 1423 1436
rect 1431 1396 1443 1436
rect 1451 1396 1463 1436
rect 1531 1396 1543 1436
rect 1551 1396 1563 1436
rect 1571 1396 1583 1436
rect 1671 1396 1683 1436
rect 1691 1400 1703 1436
rect 1711 1396 1723 1436
rect 1731 1396 1743 1436
rect 1797 1396 1809 1436
rect 1817 1396 1829 1436
rect 1837 1396 1849 1436
rect 1931 1396 1943 1436
rect 1951 1400 1963 1436
rect 1971 1396 1983 1436
rect 1991 1396 2003 1436
rect 2071 1396 2083 1436
rect 2091 1396 2103 1436
rect 2191 1396 2203 1436
rect 2211 1400 2223 1436
rect 2231 1396 2243 1436
rect 2251 1396 2263 1436
rect 2331 1396 2343 1436
rect 2351 1400 2363 1436
rect 2371 1396 2383 1436
rect 2391 1396 2403 1436
rect 2457 1396 2469 1436
rect 2477 1396 2489 1436
rect 2596 1396 2608 1436
rect 2618 1356 2630 1436
rect 2646 1356 2658 1436
rect 2717 1364 2729 1436
rect 2737 1368 2749 1436
rect 2757 1356 2769 1436
rect 2777 1356 2789 1436
rect 2876 1396 2888 1436
rect 2898 1356 2910 1436
rect 2926 1356 2938 1436
rect 3016 1396 3028 1436
rect 3038 1356 3050 1436
rect 3066 1356 3078 1436
rect 3156 1396 3168 1436
rect 3178 1356 3190 1436
rect 3206 1356 3218 1436
rect 3291 1396 3303 1436
rect 3311 1396 3323 1436
rect 3377 1396 3389 1436
rect 3397 1396 3409 1436
rect 3489 1356 3501 1436
rect 3509 1356 3521 1436
rect 3531 1396 3543 1436
rect 3631 1356 3643 1436
rect 3651 1356 3663 1436
rect 3671 1368 3683 1436
rect 3691 1364 3703 1436
rect 3762 1356 3774 1436
rect 3790 1356 3802 1436
rect 3812 1396 3824 1436
rect 3911 1396 3923 1436
rect 3931 1396 3943 1436
rect 4016 1396 4028 1436
rect 4038 1356 4050 1436
rect 4066 1356 4078 1436
rect 4156 1396 4168 1436
rect 4178 1356 4190 1436
rect 4206 1356 4218 1436
rect 4291 1356 4303 1436
rect 4311 1356 4323 1436
rect 4331 1368 4343 1436
rect 4351 1364 4363 1436
rect 4436 1396 4448 1436
rect 4458 1356 4470 1436
rect 4486 1356 4498 1436
rect 4582 1356 4594 1436
rect 4610 1356 4622 1436
rect 4632 1396 4644 1436
rect 4717 1396 4729 1436
rect 4737 1396 4749 1436
rect 4757 1396 4769 1436
rect 4842 1356 4854 1436
rect 4870 1356 4882 1436
rect 4892 1396 4904 1436
rect 4977 1356 4989 1436
rect 5005 1356 5017 1436
rect 5097 1396 5109 1436
rect 5117 1396 5129 1436
rect 5137 1396 5149 1436
rect 5231 1396 5243 1436
rect 5251 1396 5263 1436
rect 5271 1396 5283 1436
rect 5356 1396 5368 1436
rect 5378 1356 5390 1436
rect 5406 1356 5418 1436
rect 5482 1356 5494 1436
rect 5510 1356 5522 1436
rect 5532 1396 5544 1436
rect 5642 1356 5654 1436
rect 5670 1356 5682 1436
rect 5692 1396 5704 1436
rect 71 984 83 1024
rect 91 984 103 1024
rect 157 984 169 1056
rect 177 984 189 1052
rect 197 984 209 1064
rect 217 984 229 1064
rect 302 984 314 1064
rect 330 984 342 1064
rect 352 984 364 1024
rect 442 984 454 1064
rect 470 984 482 1064
rect 492 984 504 1024
rect 591 984 603 1024
rect 611 984 623 1020
rect 631 984 643 1024
rect 651 984 663 1024
rect 722 984 734 1064
rect 750 984 762 1064
rect 772 984 784 1024
rect 877 984 889 1056
rect 897 984 909 1052
rect 917 984 929 1064
rect 937 984 949 1064
rect 1036 984 1048 1024
rect 1058 984 1070 1064
rect 1086 984 1098 1064
rect 1171 984 1183 1024
rect 1191 984 1203 1024
rect 1257 984 1269 1056
rect 1277 984 1289 1052
rect 1297 984 1309 1064
rect 1317 984 1329 1064
rect 1411 984 1423 1024
rect 1431 984 1443 1024
rect 1523 984 1535 1064
rect 1551 984 1563 1064
rect 1637 984 1649 1024
rect 1657 984 1669 1024
rect 1751 984 1763 1024
rect 1771 984 1783 1020
rect 1791 984 1803 1024
rect 1811 984 1823 1024
rect 1891 984 1903 1024
rect 1911 984 1923 1024
rect 1931 984 1943 1024
rect 2016 984 2028 1024
rect 2038 984 2050 1064
rect 2066 984 2078 1064
rect 2151 984 2163 1024
rect 2171 984 2183 1020
rect 2191 984 2203 1024
rect 2211 984 2223 1024
rect 2291 984 2303 1024
rect 2311 984 2323 1020
rect 2331 984 2343 1024
rect 2351 984 2363 1024
rect 2436 984 2448 1024
rect 2458 984 2470 1064
rect 2486 984 2498 1064
rect 2571 984 2583 1024
rect 2591 984 2603 1020
rect 2611 984 2623 1024
rect 2631 984 2643 1024
rect 2717 984 2729 1024
rect 2737 984 2749 1024
rect 2817 984 2829 1064
rect 2845 984 2857 1064
rect 2937 984 2949 1064
rect 2965 984 2977 1064
rect 3057 984 3069 1024
rect 3077 984 3089 1024
rect 3101 984 3113 1064
rect 3121 984 3133 1064
rect 3223 984 3235 1064
rect 3251 984 3263 1064
rect 3363 984 3375 1064
rect 3391 984 3403 1064
rect 3471 984 3483 1024
rect 3491 984 3503 1024
rect 3576 984 3588 1024
rect 3598 984 3610 1064
rect 3626 984 3638 1064
rect 3716 984 3728 1024
rect 3738 984 3750 1064
rect 3766 984 3778 1064
rect 3837 984 3849 1024
rect 3857 984 3869 1024
rect 3877 984 3889 1024
rect 3957 984 3969 1024
rect 3977 984 3989 1024
rect 3997 984 4009 1024
rect 4077 984 4089 1064
rect 4105 984 4117 1064
rect 4197 984 4209 1024
rect 4217 984 4229 1024
rect 4311 984 4323 1064
rect 4331 984 4343 1064
rect 4351 984 4363 1052
rect 4371 984 4383 1056
rect 4476 984 4488 1024
rect 4498 984 4510 1064
rect 4526 984 4538 1064
rect 4611 984 4623 1064
rect 4631 984 4643 1064
rect 4651 984 4663 1052
rect 4671 984 4683 1056
rect 4742 984 4754 1064
rect 4770 984 4782 1064
rect 4792 984 4804 1024
rect 4877 984 4889 1024
rect 4899 984 4911 1064
rect 4919 984 4931 1064
rect 4997 984 5009 1024
rect 5017 984 5029 1024
rect 5097 984 5109 1024
rect 5117 984 5129 1024
rect 5211 984 5223 1024
rect 5231 984 5243 1024
rect 5251 984 5263 1024
rect 5356 984 5368 1024
rect 5378 984 5390 1064
rect 5406 984 5418 1064
rect 5477 984 5489 1064
rect 5505 984 5517 1064
rect 5611 984 5623 1024
rect 5631 984 5643 1020
rect 5651 984 5663 1024
rect 5671 984 5683 1024
rect 5751 984 5763 1024
rect 5771 984 5783 1024
rect 71 916 83 956
rect 91 920 103 956
rect 111 916 123 956
rect 131 916 143 956
rect 197 884 209 956
rect 217 888 229 956
rect 237 876 249 956
rect 257 876 269 956
rect 351 916 363 956
rect 371 920 383 956
rect 391 916 403 956
rect 411 916 423 956
rect 491 876 503 956
rect 511 876 523 956
rect 531 888 543 956
rect 551 884 563 956
rect 631 916 643 956
rect 651 920 663 956
rect 671 916 683 956
rect 691 916 703 956
rect 757 884 769 956
rect 777 888 789 956
rect 797 876 809 956
rect 817 876 829 956
rect 916 916 928 956
rect 938 876 950 956
rect 966 876 978 956
rect 1051 916 1063 956
rect 1071 920 1083 956
rect 1091 916 1103 956
rect 1111 916 1123 956
rect 1182 876 1194 956
rect 1210 876 1222 956
rect 1232 916 1244 956
rect 1331 916 1343 956
rect 1351 920 1363 956
rect 1371 916 1383 956
rect 1391 916 1403 956
rect 1457 916 1469 956
rect 1477 916 1489 956
rect 1557 916 1569 956
rect 1577 916 1589 956
rect 1597 916 1609 956
rect 1711 916 1723 956
rect 1731 920 1743 956
rect 1751 916 1763 956
rect 1771 916 1783 956
rect 1851 916 1863 956
rect 1871 920 1883 956
rect 1891 916 1903 956
rect 1911 916 1923 956
rect 1977 916 1989 956
rect 1997 916 2009 956
rect 2017 920 2029 956
rect 2037 916 2049 956
rect 2122 876 2134 956
rect 2150 876 2162 956
rect 2172 916 2184 956
rect 2257 916 2269 956
rect 2277 916 2289 956
rect 2301 876 2313 956
rect 2321 876 2333 956
rect 2397 916 2409 956
rect 2417 916 2429 956
rect 2511 916 2523 956
rect 2531 916 2543 956
rect 2551 916 2563 956
rect 2641 877 2653 956
rect 2661 877 2673 956
rect 2691 876 2703 956
rect 2757 916 2769 956
rect 2777 916 2789 956
rect 2797 916 2809 956
rect 2891 916 2903 956
rect 2911 916 2923 956
rect 2931 916 2943 956
rect 3017 916 3029 956
rect 3037 916 3049 956
rect 3131 916 3143 956
rect 3151 916 3163 956
rect 3251 916 3263 956
rect 3271 916 3283 956
rect 3291 916 3303 956
rect 3403 876 3415 956
rect 3431 876 3443 956
rect 3523 876 3535 956
rect 3551 876 3563 956
rect 3631 876 3643 956
rect 3651 876 3663 956
rect 3671 888 3683 956
rect 3691 884 3703 956
rect 3771 916 3783 956
rect 3791 916 3803 956
rect 3876 916 3888 956
rect 3898 876 3910 956
rect 3926 876 3938 956
rect 3997 916 4009 956
rect 4017 916 4029 956
rect 4037 916 4049 956
rect 4136 916 4148 956
rect 4158 876 4170 956
rect 4186 876 4198 956
rect 4276 916 4288 956
rect 4298 876 4310 956
rect 4326 876 4338 956
rect 4417 916 4429 956
rect 4437 916 4449 956
rect 4536 916 4548 956
rect 4558 876 4570 956
rect 4586 876 4598 956
rect 4657 884 4669 956
rect 4677 888 4689 956
rect 4697 876 4709 956
rect 4717 876 4729 956
rect 4809 876 4821 956
rect 4829 876 4841 956
rect 4851 916 4863 956
rect 4936 916 4948 956
rect 4958 876 4970 956
rect 4986 876 4998 956
rect 5057 884 5069 956
rect 5077 888 5089 956
rect 5097 876 5109 956
rect 5117 876 5129 956
rect 5221 877 5233 956
rect 5241 877 5253 956
rect 5271 876 5283 956
rect 5371 916 5383 956
rect 5391 916 5403 956
rect 5471 876 5483 956
rect 5491 876 5503 944
rect 5511 878 5523 956
rect 5531 890 5543 956
rect 5551 878 5563 956
rect 5642 876 5654 956
rect 5670 876 5682 956
rect 5692 916 5704 956
rect 71 504 83 544
rect 91 504 103 540
rect 111 504 123 544
rect 131 504 143 544
rect 231 504 243 584
rect 251 504 263 584
rect 271 504 283 572
rect 291 504 303 576
rect 371 504 383 544
rect 391 504 403 540
rect 411 504 423 544
rect 431 504 443 544
rect 516 504 528 544
rect 538 504 550 584
rect 566 504 578 584
rect 637 504 649 576
rect 657 504 669 572
rect 677 504 689 584
rect 697 504 709 584
rect 777 504 789 544
rect 797 504 809 544
rect 817 504 829 544
rect 936 504 948 544
rect 958 504 970 584
rect 986 504 998 584
rect 1071 504 1083 544
rect 1091 504 1103 540
rect 1111 504 1123 544
rect 1131 504 1143 544
rect 1197 504 1209 576
rect 1217 504 1229 572
rect 1237 504 1249 584
rect 1257 504 1269 584
rect 1351 504 1363 584
rect 1371 504 1383 584
rect 1391 504 1403 572
rect 1411 504 1423 576
rect 1497 504 1509 544
rect 1517 504 1529 544
rect 1537 504 1549 540
rect 1557 504 1569 544
rect 1656 504 1668 544
rect 1678 504 1690 584
rect 1706 504 1718 584
rect 1791 504 1803 544
rect 1811 504 1823 540
rect 1831 504 1843 544
rect 1851 504 1863 544
rect 1917 504 1929 576
rect 1937 504 1949 572
rect 1957 504 1969 584
rect 1977 504 1989 584
rect 2083 504 2095 584
rect 2111 504 2123 584
rect 2201 504 2213 583
rect 2221 504 2233 583
rect 2251 504 2263 584
rect 2317 504 2329 544
rect 2337 504 2349 544
rect 2361 504 2373 584
rect 2381 504 2393 584
rect 2457 504 2469 544
rect 2477 504 2489 544
rect 2497 504 2509 544
rect 2591 504 2603 544
rect 2611 504 2623 544
rect 2631 504 2643 544
rect 2723 504 2735 584
rect 2751 504 2763 584
rect 2822 504 2834 584
rect 2850 504 2862 584
rect 2872 504 2884 544
rect 2971 504 2983 544
rect 2991 504 3003 544
rect 3011 504 3023 544
rect 3077 504 3089 576
rect 3097 504 3109 572
rect 3117 504 3129 584
rect 3137 504 3149 584
rect 3231 504 3243 544
rect 3251 504 3263 540
rect 3271 504 3283 544
rect 3291 504 3303 544
rect 3357 504 3369 544
rect 3377 504 3389 544
rect 3397 504 3409 544
rect 3496 504 3508 544
rect 3518 504 3530 584
rect 3546 504 3558 584
rect 3617 504 3629 544
rect 3637 504 3649 544
rect 3657 504 3669 544
rect 3756 504 3768 544
rect 3778 504 3790 584
rect 3806 504 3818 584
rect 3882 504 3894 584
rect 3910 504 3922 584
rect 3932 504 3944 544
rect 4017 504 4029 576
rect 4037 504 4049 572
rect 4057 504 4069 584
rect 4077 504 4089 584
rect 4182 504 4194 584
rect 4210 504 4222 584
rect 4232 504 4244 544
rect 4331 504 4343 544
rect 4351 504 4363 544
rect 4431 504 4443 584
rect 4451 504 4463 584
rect 4471 504 4483 572
rect 4491 504 4503 576
rect 4576 504 4588 544
rect 4598 504 4610 584
rect 4626 504 4638 584
rect 4716 504 4728 544
rect 4738 504 4750 584
rect 4766 504 4778 584
rect 4862 504 4874 584
rect 4890 504 4902 584
rect 4912 504 4924 544
rect 4997 504 5009 544
rect 5017 504 5029 544
rect 5117 504 5129 544
rect 5139 504 5151 584
rect 5159 504 5171 584
rect 5256 504 5268 544
rect 5278 504 5290 584
rect 5306 504 5318 584
rect 5382 504 5394 584
rect 5410 504 5422 584
rect 5432 504 5444 544
rect 5536 504 5548 544
rect 5558 504 5570 584
rect 5586 504 5598 584
rect 5657 504 5669 584
rect 5685 504 5697 584
rect 71 436 83 476
rect 91 440 103 476
rect 111 436 123 476
rect 131 436 143 476
rect 216 436 228 476
rect 238 396 250 476
rect 266 396 278 476
rect 376 436 388 476
rect 398 396 410 476
rect 426 396 438 476
rect 511 436 523 476
rect 531 440 543 476
rect 551 436 563 476
rect 571 436 583 476
rect 647 396 659 476
rect 667 396 679 476
rect 691 436 703 476
rect 711 436 723 476
rect 791 436 803 476
rect 811 440 823 476
rect 831 436 843 476
rect 851 436 863 476
rect 931 396 943 476
rect 951 396 963 476
rect 971 408 983 476
rect 991 404 1003 476
rect 1057 436 1069 476
rect 1077 436 1089 476
rect 1097 440 1109 476
rect 1117 436 1129 476
rect 1221 397 1233 476
rect 1241 397 1253 476
rect 1271 396 1283 476
rect 1351 436 1363 476
rect 1371 440 1383 476
rect 1391 436 1403 476
rect 1411 436 1423 476
rect 1511 436 1523 476
rect 1531 436 1543 476
rect 1616 436 1628 476
rect 1638 396 1650 476
rect 1666 396 1678 476
rect 1747 396 1759 476
rect 1767 396 1779 476
rect 1791 436 1803 476
rect 1811 436 1823 476
rect 1877 396 1889 476
rect 1905 396 1917 476
rect 2017 436 2029 476
rect 2037 436 2049 476
rect 2136 436 2148 476
rect 2158 396 2170 476
rect 2186 396 2198 476
rect 2271 396 2283 476
rect 2291 396 2303 476
rect 2311 408 2323 476
rect 2331 404 2343 476
rect 2411 436 2423 476
rect 2431 436 2443 476
rect 2511 436 2523 476
rect 2531 440 2543 476
rect 2551 436 2563 476
rect 2571 436 2583 476
rect 2642 396 2654 476
rect 2670 396 2682 476
rect 2692 436 2704 476
rect 2791 436 2803 476
rect 2811 436 2823 476
rect 2903 396 2915 476
rect 2931 396 2943 476
rect 2997 436 3009 476
rect 3017 436 3029 476
rect 3111 396 3123 476
rect 3131 396 3143 476
rect 3151 408 3163 476
rect 3171 404 3183 476
rect 3257 404 3269 476
rect 3277 408 3289 476
rect 3297 396 3309 476
rect 3317 396 3329 476
rect 3411 436 3423 476
rect 3431 436 3443 476
rect 3522 396 3534 476
rect 3550 396 3562 476
rect 3572 436 3584 476
rect 3657 404 3669 476
rect 3677 408 3689 476
rect 3697 396 3709 476
rect 3717 396 3729 476
rect 3811 436 3823 476
rect 3831 440 3843 476
rect 3851 436 3863 476
rect 3871 436 3883 476
rect 3937 436 3949 476
rect 3957 436 3969 476
rect 3977 436 3989 476
rect 4091 436 4103 476
rect 4111 440 4123 476
rect 4131 436 4143 476
rect 4151 436 4163 476
rect 4236 436 4248 476
rect 4258 396 4270 476
rect 4286 396 4298 476
rect 4371 436 4383 476
rect 4391 436 4403 476
rect 4471 436 4483 476
rect 4491 436 4503 476
rect 4511 436 4523 476
rect 4596 436 4608 476
rect 4618 396 4630 476
rect 4646 396 4658 476
rect 4731 436 4743 476
rect 4751 436 4763 476
rect 4836 436 4848 476
rect 4858 396 4870 476
rect 4886 396 4898 476
rect 4957 428 4969 468
rect 4977 428 4989 468
rect 5007 404 5019 468
rect 5037 396 5049 476
rect 5136 436 5148 476
rect 5158 396 5170 476
rect 5186 396 5198 476
rect 5282 396 5294 476
rect 5310 396 5322 476
rect 5332 436 5344 476
rect 5451 396 5463 476
rect 5471 396 5483 476
rect 5491 408 5503 476
rect 5511 404 5523 476
rect 5582 396 5594 476
rect 5610 396 5622 476
rect 5632 436 5644 476
rect 5717 436 5729 476
rect 5737 436 5749 476
rect 5757 436 5769 476
rect 71 24 83 64
rect 91 24 103 60
rect 111 24 123 64
rect 131 24 143 64
rect 197 24 209 96
rect 217 24 229 92
rect 237 24 249 104
rect 257 24 269 104
rect 371 24 383 104
rect 391 24 403 104
rect 411 24 423 92
rect 431 24 443 96
rect 516 24 528 64
rect 538 24 550 104
rect 566 24 578 104
rect 642 24 654 104
rect 670 24 682 104
rect 692 24 704 64
rect 791 24 803 64
rect 811 24 823 60
rect 831 24 843 64
rect 851 24 863 64
rect 917 24 929 64
rect 937 24 949 64
rect 1022 24 1034 104
rect 1050 24 1062 104
rect 1072 24 1084 64
rect 1157 24 1169 96
rect 1177 24 1189 92
rect 1197 24 1209 104
rect 1217 24 1229 104
rect 1297 24 1309 104
rect 1325 24 1337 104
rect 1417 24 1429 64
rect 1437 24 1449 64
rect 1461 24 1473 104
rect 1481 24 1493 104
rect 1571 24 1583 64
rect 1591 24 1603 64
rect 1676 24 1688 64
rect 1698 24 1710 104
rect 1726 24 1738 104
rect 1811 24 1823 64
rect 1831 24 1843 64
rect 1851 24 1863 64
rect 1917 24 1929 64
rect 1937 24 1949 64
rect 1957 24 1969 60
rect 1977 24 1989 64
rect 2091 24 2103 64
rect 2111 24 2123 60
rect 2131 24 2143 64
rect 2151 24 2163 64
rect 2217 24 2229 64
rect 2239 24 2251 104
rect 2259 24 2271 104
rect 2351 24 2363 64
rect 2371 24 2383 64
rect 2391 24 2403 64
rect 2457 24 2469 64
rect 2477 24 2489 64
rect 2501 24 2513 104
rect 2521 24 2533 104
rect 2611 24 2623 104
rect 2631 24 2643 104
rect 2651 24 2663 92
rect 2671 24 2683 96
rect 2747 24 2759 104
rect 2767 24 2779 104
rect 2791 24 2803 64
rect 2811 24 2823 64
rect 2897 24 2909 64
rect 2917 24 2929 64
rect 2937 24 2949 64
rect 3031 24 3043 64
rect 3051 24 3063 64
rect 3071 24 3083 64
rect 3151 24 3163 64
rect 3171 24 3183 60
rect 3191 24 3203 64
rect 3211 24 3223 64
rect 3291 24 3303 64
rect 3311 24 3323 64
rect 3382 24 3394 104
rect 3410 24 3422 104
rect 3432 24 3444 64
rect 3531 24 3543 64
rect 3551 24 3563 64
rect 3631 24 3643 64
rect 3651 24 3663 64
rect 3671 24 3683 64
rect 3749 24 3761 104
rect 3769 24 3781 104
rect 3791 24 3803 64
rect 3857 24 3869 64
rect 3879 24 3891 104
rect 3899 24 3911 104
rect 3991 24 4003 64
rect 4011 24 4023 64
rect 4031 24 4043 64
rect 4117 24 4129 64
rect 4137 24 4149 64
rect 4161 24 4173 104
rect 4181 24 4193 104
rect 4303 24 4315 104
rect 4331 24 4343 104
rect 4397 24 4409 64
rect 4417 24 4429 64
rect 4437 24 4449 64
rect 4531 24 4543 64
rect 4551 24 4563 60
rect 4571 24 4583 64
rect 4591 24 4603 64
rect 4696 24 4708 64
rect 4718 24 4730 104
rect 4746 24 4758 104
rect 4817 24 4829 64
rect 4837 24 4849 64
rect 4857 24 4869 64
rect 4956 24 4968 64
rect 4978 24 4990 104
rect 5006 24 5018 104
rect 5077 24 5089 104
rect 5105 24 5117 104
rect 5211 24 5223 64
rect 5231 24 5243 64
rect 5251 24 5263 64
rect 5317 32 5329 72
rect 5337 32 5349 72
rect 5367 32 5379 96
rect 5397 24 5409 104
rect 5477 24 5489 64
rect 5497 24 5509 64
rect 5591 24 5603 64
rect 5611 24 5623 64
rect 5677 24 5689 64
rect 5697 24 5709 64
rect 5717 24 5729 64
<< psubstratepcontact >>
rect 4 5524 5816 5536
rect 4 5044 5816 5056
rect 4 4564 5816 4576
rect 4 4084 5816 4096
rect 4 3604 5816 3616
rect 4 3124 5816 3136
rect 4 2644 5816 2656
rect 4 2164 5816 2176
rect 4 1684 5816 1696
rect 4 1204 5816 1216
rect 4 724 5816 736
rect 4 244 5816 256
<< nsubstratencontact >>
rect 4 5764 5816 5776
rect 4 5284 5816 5296
rect 4 4804 5816 4816
rect 4 4324 5816 4336
rect 4 3844 5816 3856
rect 4 3364 5816 3376
rect 4 2884 5816 2896
rect 4 2404 5816 2416
rect 4 1924 5816 1936
rect 4 1444 5816 1456
rect 4 964 5816 976
rect 4 484 5816 496
rect 4 4 5816 16
<< polysilicon >>
rect 90 5756 94 5760
rect 112 5756 116 5760
rect 120 5756 124 5760
rect 216 5756 220 5760
rect 224 5756 228 5760
rect 246 5756 250 5760
rect 385 5756 389 5760
rect 405 5756 409 5760
rect 425 5756 429 5760
rect 511 5756 515 5760
rect 531 5756 535 5760
rect 551 5756 555 5760
rect 670 5756 674 5760
rect 692 5756 696 5760
rect 700 5756 704 5760
rect 805 5756 809 5760
rect 825 5756 829 5760
rect 925 5756 929 5760
rect 945 5756 949 5760
rect 965 5756 969 5760
rect 1071 5756 1075 5760
rect 1079 5756 1083 5760
rect 1235 5756 1239 5760
rect 1255 5756 1259 5760
rect 1265 5756 1269 5760
rect 1361 5756 1365 5760
rect 1383 5756 1387 5760
rect 1405 5756 1409 5760
rect 1505 5756 1509 5760
rect 1525 5756 1529 5760
rect 1545 5756 1549 5760
rect 1665 5756 1669 5760
rect 1685 5756 1689 5760
rect 1705 5756 1709 5760
rect 1805 5756 1809 5760
rect 1825 5756 1829 5760
rect 1845 5756 1849 5760
rect 1931 5756 1935 5760
rect 2050 5756 2054 5760
rect 2072 5756 2076 5760
rect 2080 5756 2084 5760
rect 2176 5756 2180 5760
rect 2184 5756 2188 5760
rect 2206 5756 2210 5760
rect 2311 5756 2315 5760
rect 2331 5756 2335 5760
rect 2351 5756 2355 5760
rect 2465 5756 2469 5760
rect 2485 5756 2489 5760
rect 2585 5756 2589 5760
rect 2605 5756 2609 5760
rect 2625 5756 2629 5760
rect 2725 5756 2729 5760
rect 2745 5756 2749 5760
rect 2765 5756 2769 5760
rect 2851 5756 2855 5760
rect 2871 5756 2875 5760
rect 2985 5756 2989 5760
rect 3090 5756 3094 5760
rect 3112 5756 3116 5760
rect 3120 5756 3124 5760
rect 3241 5756 3245 5760
rect 3263 5756 3267 5760
rect 3285 5756 3289 5760
rect 3397 5756 3401 5760
rect 3405 5756 3409 5760
rect 3505 5756 3509 5760
rect 3525 5756 3529 5760
rect 3545 5756 3549 5760
rect 3665 5756 3669 5760
rect 3765 5756 3769 5760
rect 3851 5756 3855 5760
rect 3956 5756 3960 5760
rect 3964 5756 3968 5760
rect 3986 5756 3990 5760
rect 4091 5756 4095 5760
rect 4151 5756 4155 5760
rect 4173 5756 4177 5760
rect 4181 5756 4185 5760
rect 4201 5756 4205 5760
rect 4209 5756 4213 5760
rect 4255 5756 4259 5760
rect 4275 5756 4279 5760
rect 4287 5756 4291 5760
rect 4307 5756 4311 5760
rect 4321 5756 4325 5760
rect 4341 5756 4345 5760
rect 4470 5756 4474 5760
rect 4492 5756 4496 5760
rect 4500 5756 4504 5760
rect 4605 5756 4609 5760
rect 4625 5756 4629 5760
rect 4645 5756 4649 5760
rect 4665 5756 4669 5760
rect 4685 5756 4689 5760
rect 4705 5756 4709 5760
rect 4725 5756 4729 5760
rect 4745 5756 4749 5760
rect 4845 5756 4849 5760
rect 4950 5756 4954 5760
rect 4972 5756 4976 5760
rect 4980 5756 4984 5760
rect 5085 5756 5089 5760
rect 5105 5756 5109 5760
rect 5191 5756 5195 5760
rect 5211 5756 5215 5760
rect 5316 5756 5320 5760
rect 5324 5756 5328 5760
rect 5346 5756 5350 5760
rect 5451 5756 5455 5760
rect 5551 5756 5555 5760
rect 5571 5756 5575 5760
rect 5671 5756 5675 5760
rect 90 5673 94 5716
rect 87 5661 94 5673
rect 85 5584 89 5661
rect 112 5619 116 5676
rect 120 5672 124 5676
rect 216 5672 220 5676
rect 120 5664 138 5672
rect 134 5653 138 5664
rect 202 5664 220 5672
rect 202 5653 206 5664
rect 105 5607 114 5619
rect 105 5584 109 5607
rect 134 5596 138 5641
rect 125 5589 138 5596
rect 202 5596 206 5641
rect 224 5619 228 5676
rect 246 5673 250 5716
rect 511 5708 515 5716
rect 500 5704 515 5708
rect 531 5704 535 5716
rect 246 5661 253 5673
rect 226 5607 235 5619
rect 202 5589 215 5596
rect 125 5584 129 5589
rect 211 5584 215 5589
rect 231 5584 235 5607
rect 251 5584 255 5661
rect 385 5619 389 5676
rect 405 5662 409 5676
rect 425 5662 429 5676
rect 500 5673 506 5704
rect 520 5700 535 5704
rect 520 5693 526 5700
rect 405 5656 420 5662
rect 425 5656 441 5662
rect 506 5661 516 5673
rect 414 5633 420 5656
rect 385 5607 394 5619
rect 392 5564 396 5607
rect 414 5584 418 5621
rect 434 5619 441 5656
rect 434 5594 441 5607
rect 512 5604 516 5661
rect 520 5604 524 5681
rect 551 5673 555 5716
rect 670 5673 674 5716
rect 528 5661 535 5673
rect 547 5661 555 5673
rect 667 5661 674 5673
rect 528 5604 532 5661
rect 422 5588 441 5594
rect 422 5584 426 5588
rect 665 5584 669 5661
rect 692 5619 696 5676
rect 700 5672 704 5676
rect 700 5664 718 5672
rect 714 5653 718 5664
rect 685 5607 694 5619
rect 685 5584 689 5607
rect 714 5596 718 5641
rect 805 5639 809 5716
rect 806 5627 809 5639
rect 803 5611 809 5627
rect 825 5639 829 5716
rect 825 5627 834 5639
rect 825 5611 831 5627
rect 803 5604 817 5611
rect 705 5589 718 5596
rect 705 5584 709 5589
rect 813 5584 817 5604
rect 823 5604 831 5611
rect 925 5619 929 5676
rect 945 5662 949 5676
rect 965 5662 969 5676
rect 945 5656 960 5662
rect 965 5656 981 5662
rect 954 5633 960 5656
rect 925 5607 934 5619
rect 823 5584 827 5604
rect 932 5564 936 5607
rect 954 5584 958 5621
rect 974 5619 981 5656
rect 1071 5653 1075 5676
rect 1066 5641 1075 5653
rect 1079 5653 1083 5676
rect 1235 5671 1239 5676
rect 1255 5653 1259 5676
rect 1265 5672 1269 5676
rect 1265 5667 1278 5672
rect 1079 5641 1094 5653
rect 974 5594 981 5607
rect 962 5588 981 5594
rect 962 5584 966 5588
rect 1071 5564 1075 5641
rect 1091 5564 1095 5641
rect 1225 5592 1235 5604
rect 1225 5584 1229 5592
rect 1255 5577 1259 5641
rect 1245 5571 1259 5577
rect 1274 5633 1278 5667
rect 1274 5576 1278 5621
rect 1361 5602 1365 5676
rect 1383 5639 1387 5716
rect 1405 5653 1409 5716
rect 1505 5673 1509 5716
rect 1525 5704 1529 5716
rect 1545 5708 1549 5716
rect 1545 5704 1560 5708
rect 1525 5700 1540 5704
rect 1534 5693 1540 5700
rect 1505 5661 1513 5673
rect 1525 5661 1532 5673
rect 1405 5641 1414 5653
rect 1386 5627 1399 5639
rect 1361 5590 1373 5602
rect 1375 5584 1379 5590
rect 1395 5584 1399 5627
rect 1405 5584 1409 5641
rect 1528 5604 1532 5661
rect 1536 5604 1540 5681
rect 1554 5673 1560 5704
rect 1544 5661 1554 5673
rect 1544 5604 1548 5661
rect 1665 5619 1669 5676
rect 1685 5662 1689 5676
rect 1705 5662 1709 5676
rect 1805 5673 1809 5716
rect 1825 5704 1829 5716
rect 1845 5708 1849 5716
rect 1845 5704 1860 5708
rect 1825 5700 1840 5704
rect 1834 5693 1840 5700
rect 1685 5656 1700 5662
rect 1705 5656 1721 5662
rect 1805 5661 1813 5673
rect 1825 5661 1832 5673
rect 1694 5633 1700 5656
rect 1665 5607 1674 5619
rect 1265 5571 1278 5576
rect 1245 5564 1249 5571
rect 1265 5564 1269 5571
rect 1672 5564 1676 5607
rect 1694 5584 1698 5621
rect 1714 5619 1721 5656
rect 1714 5594 1721 5607
rect 1828 5604 1832 5661
rect 1836 5604 1840 5681
rect 1854 5673 1860 5704
rect 1844 5661 1854 5673
rect 1844 5604 1848 5661
rect 1931 5633 1935 5716
rect 2050 5673 2054 5716
rect 2047 5661 2054 5673
rect 1926 5621 1935 5633
rect 1702 5588 1721 5594
rect 1702 5584 1706 5588
rect 1931 5564 1935 5621
rect 2045 5584 2049 5661
rect 2072 5619 2076 5676
rect 2080 5672 2084 5676
rect 2176 5672 2180 5676
rect 2080 5664 2098 5672
rect 2094 5653 2098 5664
rect 2162 5664 2180 5672
rect 2162 5653 2166 5664
rect 2065 5607 2074 5619
rect 2065 5584 2069 5607
rect 2094 5596 2098 5641
rect 2085 5589 2098 5596
rect 2162 5596 2166 5641
rect 2184 5619 2188 5676
rect 2206 5673 2210 5716
rect 2206 5661 2213 5673
rect 2311 5662 2315 5676
rect 2331 5662 2335 5676
rect 2186 5607 2195 5619
rect 2162 5589 2175 5596
rect 2085 5584 2089 5589
rect 2171 5584 2175 5589
rect 2191 5584 2195 5607
rect 2211 5584 2215 5661
rect 2299 5656 2315 5662
rect 2320 5656 2335 5662
rect 2299 5619 2306 5656
rect 2320 5633 2326 5656
rect 2299 5594 2306 5607
rect 2299 5588 2318 5594
rect 2314 5584 2318 5588
rect 2322 5584 2326 5621
rect 2351 5619 2355 5676
rect 2465 5639 2469 5716
rect 2466 5627 2469 5639
rect 2346 5607 2355 5619
rect 2463 5611 2469 5627
rect 2485 5639 2489 5716
rect 2585 5673 2589 5716
rect 2605 5704 2609 5716
rect 2625 5708 2629 5716
rect 2625 5704 2640 5708
rect 2605 5700 2620 5704
rect 2614 5693 2620 5700
rect 2585 5661 2593 5673
rect 2605 5661 2612 5673
rect 2485 5627 2494 5639
rect 2485 5611 2491 5627
rect 2344 5564 2348 5607
rect 2463 5604 2477 5611
rect 2473 5584 2477 5604
rect 2483 5604 2491 5611
rect 2608 5604 2612 5661
rect 2616 5604 2620 5681
rect 2634 5673 2640 5704
rect 2725 5673 2729 5716
rect 2745 5704 2749 5716
rect 2765 5708 2769 5716
rect 2765 5704 2780 5708
rect 2745 5700 2760 5704
rect 2754 5693 2760 5700
rect 2624 5661 2634 5673
rect 2725 5661 2733 5673
rect 2745 5661 2752 5673
rect 2624 5604 2628 5661
rect 2748 5604 2752 5661
rect 2756 5604 2760 5681
rect 2774 5673 2780 5704
rect 2764 5661 2774 5673
rect 2764 5604 2768 5661
rect 2851 5639 2855 5716
rect 2846 5627 2855 5639
rect 2849 5611 2855 5627
rect 2871 5639 2875 5716
rect 2871 5627 2874 5639
rect 2985 5633 2989 5716
rect 3090 5673 3094 5716
rect 3087 5661 3094 5673
rect 2871 5611 2877 5627
rect 2849 5604 2857 5611
rect 2483 5584 2487 5604
rect 2853 5584 2857 5604
rect 2863 5604 2877 5611
rect 2985 5621 2994 5633
rect 2863 5584 2867 5604
rect 2985 5564 2989 5621
rect 3085 5584 3089 5661
rect 3112 5619 3116 5676
rect 3120 5672 3124 5676
rect 3120 5664 3138 5672
rect 3134 5653 3138 5664
rect 3105 5607 3114 5619
rect 3105 5584 3109 5607
rect 3134 5596 3138 5641
rect 3125 5589 3138 5596
rect 3241 5602 3245 5676
rect 3263 5639 3267 5716
rect 3285 5653 3289 5716
rect 3397 5653 3401 5676
rect 3285 5641 3294 5653
rect 3386 5641 3401 5653
rect 3405 5653 3409 5676
rect 3505 5673 3509 5716
rect 3525 5704 3529 5716
rect 3545 5708 3549 5716
rect 3545 5704 3560 5708
rect 3525 5700 3540 5704
rect 3534 5693 3540 5700
rect 3505 5661 3513 5673
rect 3525 5661 3532 5673
rect 3405 5641 3414 5653
rect 3266 5627 3279 5639
rect 3241 5590 3253 5602
rect 3125 5584 3129 5589
rect 3255 5584 3259 5590
rect 3275 5584 3279 5627
rect 3285 5584 3289 5641
rect 3385 5564 3389 5641
rect 3405 5564 3409 5641
rect 3528 5604 3532 5661
rect 3536 5604 3540 5681
rect 3554 5673 3560 5704
rect 3544 5661 3554 5673
rect 3544 5604 3548 5661
rect 3665 5633 3669 5716
rect 3765 5633 3769 5716
rect 3851 5633 3855 5716
rect 3956 5672 3960 5676
rect 3942 5664 3960 5672
rect 3942 5653 3946 5664
rect 3665 5621 3674 5633
rect 3765 5621 3774 5633
rect 3846 5621 3855 5633
rect 3665 5564 3669 5621
rect 3765 5564 3769 5621
rect 3851 5564 3855 5621
rect 3942 5596 3946 5641
rect 3964 5619 3968 5676
rect 3986 5673 3990 5716
rect 3986 5661 3993 5673
rect 3966 5607 3975 5619
rect 3942 5589 3955 5596
rect 3951 5584 3955 5589
rect 3971 5584 3975 5607
rect 3991 5584 3995 5661
rect 4091 5633 4095 5716
rect 4173 5713 4177 5736
rect 4169 5706 4177 5713
rect 4169 5677 4173 5706
rect 4181 5696 4185 5736
rect 4201 5684 4205 5716
rect 4209 5712 4213 5716
rect 4209 5710 4245 5712
rect 4209 5708 4233 5710
rect 4086 5621 4095 5633
rect 4091 5564 4095 5621
rect 4151 5664 4155 5676
rect 4169 5671 4177 5677
rect 4151 5652 4153 5664
rect 4151 5584 4155 5652
rect 4173 5625 4177 5671
rect 4173 5564 4177 5613
rect 4201 5589 4207 5684
rect 4183 5585 4207 5589
rect 4183 5564 4187 5585
rect 4203 5580 4221 5581
rect 4203 5576 4233 5580
rect 4203 5564 4207 5576
rect 4241 5572 4245 5698
rect 4255 5690 4259 5716
rect 4275 5710 4279 5716
rect 4211 5568 4245 5572
rect 4211 5564 4215 5568
rect 4257 5564 4261 5678
rect 4273 5588 4277 5698
rect 4287 5676 4291 5716
rect 4282 5664 4285 5676
rect 4282 5600 4286 5664
rect 4307 5657 4311 5716
rect 4302 5649 4311 5657
rect 4302 5620 4306 5649
rect 4321 5634 4325 5716
rect 4341 5633 4345 5676
rect 4470 5673 4474 5716
rect 4467 5661 4474 5673
rect 4282 5596 4315 5600
rect 4281 5576 4283 5588
rect 4279 5564 4283 5576
rect 4289 5576 4291 5588
rect 4289 5564 4293 5576
rect 4311 5564 4315 5596
rect 4321 5564 4325 5622
rect 4341 5584 4345 5621
rect 4465 5584 4469 5661
rect 4492 5619 4496 5676
rect 4500 5672 4504 5676
rect 4500 5664 4518 5672
rect 4514 5653 4518 5664
rect 4485 5607 4494 5619
rect 4485 5584 4489 5607
rect 4514 5596 4518 5641
rect 4505 5589 4518 5596
rect 4605 5616 4609 5676
rect 4625 5616 4629 5676
rect 4645 5616 4649 5676
rect 4665 5616 4669 5676
rect 4685 5616 4689 5676
rect 4705 5616 4709 5676
rect 4725 5619 4729 5676
rect 4745 5619 4749 5676
rect 4605 5604 4618 5616
rect 4645 5604 4658 5616
rect 4685 5604 4698 5616
rect 4725 5607 4734 5619
rect 4746 5607 4749 5619
rect 4505 5584 4509 5589
rect 4605 5584 4609 5604
rect 4625 5584 4629 5604
rect 4645 5584 4649 5604
rect 4665 5584 4669 5604
rect 4685 5584 4689 5604
rect 4705 5584 4709 5604
rect 4725 5584 4729 5607
rect 4745 5584 4749 5607
rect 4845 5633 4849 5716
rect 4950 5673 4954 5716
rect 4947 5661 4954 5673
rect 4845 5621 4854 5633
rect 4845 5564 4849 5621
rect 4945 5584 4949 5661
rect 4972 5619 4976 5676
rect 4980 5672 4984 5676
rect 4980 5664 4998 5672
rect 4994 5653 4998 5664
rect 4965 5607 4974 5619
rect 4965 5584 4969 5607
rect 4994 5596 4998 5641
rect 5085 5639 5089 5716
rect 5086 5627 5089 5639
rect 5083 5611 5089 5627
rect 5105 5639 5109 5716
rect 5191 5639 5195 5716
rect 5105 5627 5114 5639
rect 5186 5627 5195 5639
rect 5105 5611 5111 5627
rect 5083 5604 5097 5611
rect 4985 5589 4998 5596
rect 4985 5584 4989 5589
rect 5093 5584 5097 5604
rect 5103 5604 5111 5611
rect 5189 5611 5195 5627
rect 5211 5639 5215 5716
rect 5316 5672 5320 5676
rect 5302 5664 5320 5672
rect 5302 5653 5306 5664
rect 5211 5627 5214 5639
rect 5211 5611 5217 5627
rect 5189 5604 5197 5611
rect 5103 5584 5107 5604
rect 5193 5584 5197 5604
rect 5203 5604 5217 5611
rect 5203 5584 5207 5604
rect 5302 5596 5306 5641
rect 5324 5619 5328 5676
rect 5346 5673 5350 5716
rect 5346 5661 5353 5673
rect 5326 5607 5335 5619
rect 5302 5589 5315 5596
rect 5311 5584 5315 5589
rect 5331 5584 5335 5607
rect 5351 5584 5355 5661
rect 5451 5633 5455 5716
rect 5551 5639 5555 5716
rect 5446 5621 5455 5633
rect 5546 5627 5555 5639
rect 5451 5564 5455 5621
rect 5549 5611 5555 5627
rect 5571 5639 5575 5716
rect 5571 5627 5574 5639
rect 5671 5633 5675 5716
rect 5571 5611 5577 5627
rect 5666 5621 5675 5633
rect 5549 5604 5557 5611
rect 5553 5584 5557 5604
rect 5563 5604 5577 5611
rect 5563 5584 5567 5604
rect 5671 5564 5675 5621
rect 85 5540 89 5544
rect 105 5540 109 5544
rect 125 5540 129 5544
rect 211 5540 215 5544
rect 231 5540 235 5544
rect 251 5540 255 5544
rect 392 5540 396 5544
rect 414 5540 418 5544
rect 422 5540 426 5544
rect 512 5540 516 5544
rect 520 5540 524 5544
rect 528 5540 532 5544
rect 665 5540 669 5544
rect 685 5540 689 5544
rect 705 5540 709 5544
rect 813 5540 817 5544
rect 823 5540 827 5544
rect 932 5540 936 5544
rect 954 5540 958 5544
rect 962 5540 966 5544
rect 1071 5540 1075 5544
rect 1091 5540 1095 5544
rect 1225 5540 1229 5544
rect 1245 5540 1249 5544
rect 1265 5540 1269 5544
rect 1375 5540 1379 5544
rect 1395 5540 1399 5544
rect 1405 5540 1409 5544
rect 1528 5540 1532 5544
rect 1536 5540 1540 5544
rect 1544 5540 1548 5544
rect 1672 5540 1676 5544
rect 1694 5540 1698 5544
rect 1702 5540 1706 5544
rect 1828 5540 1832 5544
rect 1836 5540 1840 5544
rect 1844 5540 1848 5544
rect 1931 5540 1935 5544
rect 2045 5540 2049 5544
rect 2065 5540 2069 5544
rect 2085 5540 2089 5544
rect 2171 5540 2175 5544
rect 2191 5540 2195 5544
rect 2211 5540 2215 5544
rect 2314 5540 2318 5544
rect 2322 5540 2326 5544
rect 2344 5540 2348 5544
rect 2473 5540 2477 5544
rect 2483 5540 2487 5544
rect 2608 5540 2612 5544
rect 2616 5540 2620 5544
rect 2624 5540 2628 5544
rect 2748 5540 2752 5544
rect 2756 5540 2760 5544
rect 2764 5540 2768 5544
rect 2853 5540 2857 5544
rect 2863 5540 2867 5544
rect 2985 5540 2989 5544
rect 3085 5540 3089 5544
rect 3105 5540 3109 5544
rect 3125 5540 3129 5544
rect 3255 5540 3259 5544
rect 3275 5540 3279 5544
rect 3285 5540 3289 5544
rect 3385 5540 3389 5544
rect 3405 5540 3409 5544
rect 3528 5540 3532 5544
rect 3536 5540 3540 5544
rect 3544 5540 3548 5544
rect 3665 5540 3669 5544
rect 3765 5540 3769 5544
rect 3851 5540 3855 5544
rect 3951 5540 3955 5544
rect 3971 5540 3975 5544
rect 3991 5540 3995 5544
rect 4091 5540 4095 5544
rect 4151 5540 4155 5544
rect 4173 5540 4177 5544
rect 4183 5540 4187 5544
rect 4203 5540 4207 5544
rect 4211 5540 4215 5544
rect 4257 5540 4261 5544
rect 4279 5540 4283 5544
rect 4289 5540 4293 5544
rect 4311 5540 4315 5544
rect 4321 5540 4325 5544
rect 4341 5540 4345 5544
rect 4465 5540 4469 5544
rect 4485 5540 4489 5544
rect 4505 5540 4509 5544
rect 4605 5540 4609 5544
rect 4625 5540 4629 5544
rect 4645 5540 4649 5544
rect 4665 5540 4669 5544
rect 4685 5540 4689 5544
rect 4705 5540 4709 5544
rect 4725 5540 4729 5544
rect 4745 5540 4749 5544
rect 4845 5540 4849 5544
rect 4945 5540 4949 5544
rect 4965 5540 4969 5544
rect 4985 5540 4989 5544
rect 5093 5540 5097 5544
rect 5103 5540 5107 5544
rect 5193 5540 5197 5544
rect 5203 5540 5207 5544
rect 5311 5540 5315 5544
rect 5331 5540 5335 5544
rect 5351 5540 5355 5544
rect 5451 5540 5455 5544
rect 5553 5540 5557 5544
rect 5563 5540 5567 5544
rect 5671 5540 5675 5544
rect 85 5516 89 5520
rect 105 5516 109 5520
rect 125 5516 129 5520
rect 268 5516 272 5520
rect 276 5516 280 5520
rect 284 5516 288 5520
rect 408 5516 412 5520
rect 416 5516 420 5520
rect 424 5516 428 5520
rect 548 5516 552 5520
rect 556 5516 560 5520
rect 564 5516 568 5520
rect 672 5516 676 5520
rect 680 5516 684 5520
rect 688 5516 692 5520
rect 811 5516 815 5520
rect 831 5516 835 5520
rect 851 5516 855 5520
rect 952 5516 956 5520
rect 960 5516 964 5520
rect 968 5516 972 5520
rect 1112 5516 1116 5520
rect 1134 5516 1138 5520
rect 1142 5516 1146 5520
rect 1232 5516 1236 5520
rect 1240 5516 1244 5520
rect 1248 5516 1252 5520
rect 1391 5516 1395 5520
rect 1411 5516 1415 5520
rect 1548 5516 1552 5520
rect 1556 5516 1560 5520
rect 1564 5516 1568 5520
rect 1651 5516 1655 5520
rect 1671 5516 1675 5520
rect 1691 5516 1695 5520
rect 1828 5516 1832 5520
rect 1836 5516 1840 5520
rect 1844 5516 1848 5520
rect 1968 5516 1972 5520
rect 1976 5516 1980 5520
rect 1984 5516 1988 5520
rect 2073 5516 2077 5520
rect 2083 5516 2087 5520
rect 2225 5516 2229 5520
rect 2335 5516 2339 5520
rect 2355 5516 2359 5520
rect 2365 5516 2369 5520
rect 2451 5516 2455 5520
rect 2471 5516 2475 5520
rect 2491 5516 2495 5520
rect 2648 5516 2652 5520
rect 2656 5516 2660 5520
rect 2664 5516 2668 5520
rect 2788 5516 2792 5520
rect 2796 5516 2800 5520
rect 2804 5516 2808 5520
rect 2891 5516 2895 5520
rect 2911 5516 2915 5520
rect 2931 5516 2935 5520
rect 3031 5516 3035 5520
rect 3133 5516 3137 5520
rect 3143 5516 3147 5520
rect 3272 5516 3276 5520
rect 3280 5516 3284 5520
rect 3288 5516 3292 5520
rect 3413 5516 3417 5520
rect 3423 5516 3427 5520
rect 3531 5516 3535 5520
rect 3551 5516 3555 5520
rect 3571 5516 3575 5520
rect 3708 5516 3712 5520
rect 3716 5516 3720 5520
rect 3724 5516 3728 5520
rect 3832 5516 3836 5520
rect 3854 5516 3858 5520
rect 3862 5516 3866 5520
rect 3953 5516 3957 5520
rect 3963 5516 3967 5520
rect 4085 5516 4089 5520
rect 4105 5516 4109 5520
rect 4125 5516 4129 5520
rect 4233 5516 4237 5520
rect 4243 5516 4247 5520
rect 4368 5516 4372 5520
rect 4376 5516 4380 5520
rect 4384 5516 4388 5520
rect 4494 5516 4498 5520
rect 4502 5516 4506 5520
rect 4524 5516 4528 5520
rect 4631 5516 4635 5520
rect 4731 5516 4735 5520
rect 4751 5516 4755 5520
rect 4771 5516 4775 5520
rect 4831 5516 4835 5520
rect 4853 5516 4857 5520
rect 4863 5516 4867 5520
rect 4883 5516 4887 5520
rect 4891 5516 4895 5520
rect 4937 5516 4941 5520
rect 4959 5516 4963 5520
rect 4969 5516 4973 5520
rect 4991 5516 4995 5520
rect 5001 5516 5005 5520
rect 5021 5516 5025 5520
rect 5111 5516 5115 5520
rect 5171 5516 5175 5520
rect 5193 5516 5197 5520
rect 5203 5516 5207 5520
rect 5223 5516 5227 5520
rect 5231 5516 5235 5520
rect 5277 5516 5281 5520
rect 5299 5516 5303 5520
rect 5309 5516 5313 5520
rect 5331 5516 5335 5520
rect 5341 5516 5345 5520
rect 5361 5516 5365 5520
rect 5451 5516 5455 5520
rect 5471 5516 5475 5520
rect 5491 5516 5495 5520
rect 5613 5516 5617 5520
rect 5623 5516 5627 5520
rect 5733 5516 5737 5520
rect 5743 5516 5747 5520
rect 85 5399 89 5476
rect 105 5453 109 5476
rect 125 5471 129 5476
rect 125 5464 138 5471
rect 105 5441 114 5453
rect 87 5387 94 5399
rect 90 5344 94 5387
rect 112 5384 116 5441
rect 134 5419 138 5464
rect 811 5471 815 5476
rect 802 5464 815 5471
rect 134 5396 138 5407
rect 268 5399 272 5456
rect 120 5388 138 5396
rect 120 5384 124 5388
rect 245 5387 253 5399
rect 265 5387 272 5399
rect 245 5344 249 5387
rect 276 5379 280 5456
rect 284 5399 288 5456
rect 408 5399 412 5456
rect 284 5387 294 5399
rect 385 5387 393 5399
rect 405 5387 412 5399
rect 274 5360 280 5367
rect 265 5356 280 5360
rect 294 5356 300 5387
rect 265 5344 269 5356
rect 285 5352 300 5356
rect 285 5344 289 5352
rect 385 5344 389 5387
rect 416 5379 420 5456
rect 424 5399 428 5456
rect 548 5399 552 5456
rect 424 5387 434 5399
rect 525 5387 533 5399
rect 545 5387 552 5399
rect 414 5360 420 5367
rect 405 5356 420 5360
rect 434 5356 440 5387
rect 405 5344 409 5356
rect 425 5352 440 5356
rect 425 5344 429 5352
rect 525 5344 529 5387
rect 556 5379 560 5456
rect 564 5399 568 5456
rect 672 5399 676 5456
rect 564 5387 574 5399
rect 666 5387 676 5399
rect 554 5360 560 5367
rect 545 5356 560 5360
rect 574 5356 580 5387
rect 545 5344 549 5356
rect 565 5352 580 5356
rect 660 5356 666 5387
rect 680 5379 684 5456
rect 688 5399 692 5456
rect 802 5419 806 5464
rect 831 5453 835 5476
rect 826 5441 835 5453
rect 688 5387 695 5399
rect 707 5387 715 5399
rect 802 5396 806 5407
rect 802 5388 820 5396
rect 680 5360 686 5367
rect 680 5356 695 5360
rect 660 5352 675 5356
rect 565 5344 569 5352
rect 671 5344 675 5352
rect 691 5344 695 5356
rect 711 5344 715 5387
rect 816 5384 820 5388
rect 824 5384 828 5441
rect 851 5399 855 5476
rect 952 5399 956 5456
rect 846 5387 853 5399
rect 946 5387 956 5399
rect 846 5344 850 5387
rect 940 5356 946 5387
rect 960 5379 964 5456
rect 968 5399 972 5456
rect 1112 5453 1116 5496
rect 1105 5441 1114 5453
rect 968 5387 975 5399
rect 987 5387 995 5399
rect 960 5360 966 5367
rect 960 5356 975 5360
rect 940 5352 955 5356
rect 951 5344 955 5352
rect 971 5344 975 5356
rect 991 5344 995 5387
rect 1105 5384 1109 5441
rect 1134 5439 1138 5476
rect 1142 5472 1146 5476
rect 1142 5466 1161 5472
rect 1154 5453 1161 5466
rect 1134 5404 1140 5427
rect 1154 5404 1161 5441
rect 1125 5398 1140 5404
rect 1145 5398 1161 5404
rect 1232 5399 1236 5456
rect 1125 5384 1129 5398
rect 1145 5384 1149 5398
rect 1226 5387 1236 5399
rect 1220 5356 1226 5387
rect 1240 5379 1244 5456
rect 1248 5399 1252 5456
rect 1391 5419 1395 5496
rect 1411 5419 1415 5496
rect 1651 5471 1655 5476
rect 1642 5464 1655 5471
rect 1386 5407 1395 5419
rect 1248 5387 1255 5399
rect 1267 5387 1275 5399
rect 1240 5360 1246 5367
rect 1240 5356 1255 5360
rect 1220 5352 1235 5356
rect 1231 5344 1235 5352
rect 1251 5344 1255 5356
rect 1271 5344 1275 5387
rect 1391 5384 1395 5407
rect 1399 5407 1414 5419
rect 1399 5384 1403 5407
rect 1548 5399 1552 5456
rect 1525 5387 1533 5399
rect 1545 5387 1552 5399
rect 1525 5344 1529 5387
rect 1556 5379 1560 5456
rect 1564 5399 1568 5456
rect 1642 5419 1646 5464
rect 1671 5453 1675 5476
rect 1666 5441 1675 5453
rect 1564 5387 1574 5399
rect 1642 5396 1646 5407
rect 1642 5388 1660 5396
rect 1554 5360 1560 5367
rect 1545 5356 1560 5360
rect 1574 5356 1580 5387
rect 1656 5384 1660 5388
rect 1664 5384 1668 5441
rect 1691 5399 1695 5476
rect 2073 5456 2077 5476
rect 1828 5399 1832 5456
rect 1686 5387 1693 5399
rect 1805 5387 1813 5399
rect 1825 5387 1832 5399
rect 1545 5344 1549 5356
rect 1565 5352 1580 5356
rect 1565 5344 1569 5352
rect 1686 5344 1690 5387
rect 1805 5344 1809 5387
rect 1836 5379 1840 5456
rect 1844 5399 1848 5456
rect 1968 5399 1972 5456
rect 1844 5387 1854 5399
rect 1945 5387 1953 5399
rect 1965 5387 1972 5399
rect 1834 5360 1840 5367
rect 1825 5356 1840 5360
rect 1854 5356 1860 5387
rect 1825 5344 1829 5356
rect 1845 5352 1860 5356
rect 1845 5344 1849 5352
rect 1945 5344 1949 5387
rect 1976 5379 1980 5456
rect 1984 5399 1988 5456
rect 2069 5449 2077 5456
rect 2083 5456 2087 5476
rect 2083 5449 2097 5456
rect 2069 5433 2075 5449
rect 2066 5421 2075 5433
rect 1984 5387 1994 5399
rect 1974 5360 1980 5367
rect 1965 5356 1980 5360
rect 1994 5356 2000 5387
rect 1965 5344 1969 5356
rect 1985 5352 2000 5356
rect 1985 5344 1989 5352
rect 2071 5344 2075 5421
rect 2091 5433 2097 5449
rect 2225 5439 2229 5496
rect 2335 5470 2339 5476
rect 2321 5458 2333 5470
rect 2091 5421 2094 5433
rect 2225 5427 2234 5439
rect 2091 5344 2095 5421
rect 2225 5344 2229 5427
rect 2321 5384 2325 5458
rect 2355 5433 2359 5476
rect 2346 5421 2359 5433
rect 2343 5344 2347 5421
rect 2365 5419 2369 5476
rect 2451 5471 2455 5476
rect 2442 5464 2455 5471
rect 2442 5419 2446 5464
rect 2471 5453 2475 5476
rect 2466 5441 2475 5453
rect 2365 5407 2374 5419
rect 2365 5344 2369 5407
rect 2442 5396 2446 5407
rect 2442 5388 2460 5396
rect 2456 5384 2460 5388
rect 2464 5384 2468 5441
rect 2491 5399 2495 5476
rect 2891 5471 2895 5476
rect 2882 5464 2895 5471
rect 2648 5399 2652 5456
rect 2486 5387 2493 5399
rect 2625 5387 2633 5399
rect 2645 5387 2652 5399
rect 2486 5344 2490 5387
rect 2625 5344 2629 5387
rect 2656 5379 2660 5456
rect 2664 5399 2668 5456
rect 2788 5399 2792 5456
rect 2664 5387 2674 5399
rect 2765 5387 2773 5399
rect 2785 5387 2792 5399
rect 2654 5360 2660 5367
rect 2645 5356 2660 5360
rect 2674 5356 2680 5387
rect 2645 5344 2649 5356
rect 2665 5352 2680 5356
rect 2665 5344 2669 5352
rect 2765 5344 2769 5387
rect 2796 5379 2800 5456
rect 2804 5399 2808 5456
rect 2882 5419 2886 5464
rect 2911 5453 2915 5476
rect 2906 5441 2915 5453
rect 2804 5387 2814 5399
rect 2882 5396 2886 5407
rect 2882 5388 2900 5396
rect 2794 5360 2800 5367
rect 2785 5356 2800 5360
rect 2814 5356 2820 5387
rect 2896 5384 2900 5388
rect 2904 5384 2908 5441
rect 2931 5399 2935 5476
rect 3031 5439 3035 5496
rect 3133 5456 3137 5476
rect 3026 5427 3035 5439
rect 3129 5449 3137 5456
rect 3143 5456 3147 5476
rect 3531 5489 3535 5496
rect 3551 5489 3555 5496
rect 3522 5484 3535 5489
rect 3413 5456 3417 5476
rect 3143 5449 3157 5456
rect 3129 5433 3135 5449
rect 2926 5387 2933 5399
rect 2785 5344 2789 5356
rect 2805 5352 2820 5356
rect 2805 5344 2809 5352
rect 2926 5344 2930 5387
rect 3031 5344 3035 5427
rect 3126 5421 3135 5433
rect 3131 5344 3135 5421
rect 3151 5433 3157 5449
rect 3151 5421 3154 5433
rect 3151 5344 3155 5421
rect 3272 5399 3276 5456
rect 3266 5387 3276 5399
rect 3260 5356 3266 5387
rect 3280 5379 3284 5456
rect 3288 5399 3292 5456
rect 3409 5449 3417 5456
rect 3423 5456 3427 5476
rect 3423 5449 3437 5456
rect 3409 5433 3415 5449
rect 3406 5421 3415 5433
rect 3288 5387 3295 5399
rect 3307 5387 3315 5399
rect 3280 5360 3286 5367
rect 3280 5356 3295 5360
rect 3260 5352 3275 5356
rect 3271 5344 3275 5352
rect 3291 5344 3295 5356
rect 3311 5344 3315 5387
rect 3411 5344 3415 5421
rect 3431 5433 3437 5449
rect 3522 5439 3526 5484
rect 3431 5421 3434 5433
rect 3431 5344 3435 5421
rect 3522 5393 3526 5427
rect 3541 5483 3555 5489
rect 3541 5419 3545 5483
rect 3571 5468 3575 5476
rect 3565 5456 3575 5468
rect 3522 5388 3535 5393
rect 3531 5384 3535 5388
rect 3541 5384 3545 5407
rect 3708 5399 3712 5456
rect 3561 5384 3565 5389
rect 3685 5387 3693 5399
rect 3705 5387 3712 5399
rect 3685 5344 3689 5387
rect 3716 5379 3720 5456
rect 3724 5399 3728 5456
rect 3832 5453 3836 5496
rect 3825 5441 3834 5453
rect 3724 5387 3734 5399
rect 3714 5360 3720 5367
rect 3705 5356 3720 5360
rect 3734 5356 3740 5387
rect 3825 5384 3829 5441
rect 3854 5439 3858 5476
rect 3862 5472 3866 5476
rect 3862 5466 3881 5472
rect 3874 5453 3881 5466
rect 3953 5456 3957 5476
rect 3949 5449 3957 5456
rect 3963 5456 3967 5476
rect 3963 5449 3977 5456
rect 3854 5404 3860 5427
rect 3874 5404 3881 5441
rect 3949 5433 3955 5449
rect 3946 5421 3955 5433
rect 3845 5398 3860 5404
rect 3865 5398 3881 5404
rect 3845 5384 3849 5398
rect 3865 5384 3869 5398
rect 3705 5344 3709 5356
rect 3725 5352 3740 5356
rect 3725 5344 3729 5352
rect 3951 5344 3955 5421
rect 3971 5433 3977 5449
rect 3971 5421 3974 5433
rect 3971 5344 3975 5421
rect 4085 5399 4089 5476
rect 4105 5453 4109 5476
rect 4125 5471 4129 5476
rect 4125 5464 4138 5471
rect 4105 5441 4114 5453
rect 4087 5387 4094 5399
rect 4090 5344 4094 5387
rect 4112 5384 4116 5441
rect 4134 5419 4138 5464
rect 4233 5456 4237 5476
rect 4223 5449 4237 5456
rect 4243 5456 4247 5476
rect 4494 5472 4498 5476
rect 4479 5466 4498 5472
rect 4243 5449 4251 5456
rect 4223 5433 4229 5449
rect 4226 5421 4229 5433
rect 4134 5396 4138 5407
rect 4120 5388 4138 5396
rect 4120 5384 4124 5388
rect 4225 5344 4229 5421
rect 4245 5433 4251 5449
rect 4245 5421 4254 5433
rect 4245 5344 4249 5421
rect 4368 5399 4372 5456
rect 4345 5387 4353 5399
rect 4365 5387 4372 5399
rect 4345 5344 4349 5387
rect 4376 5379 4380 5456
rect 4384 5399 4388 5456
rect 4479 5453 4486 5466
rect 4479 5404 4486 5441
rect 4502 5439 4506 5476
rect 4524 5453 4528 5496
rect 4526 5441 4535 5453
rect 4500 5404 4506 5427
rect 4384 5387 4394 5399
rect 4479 5398 4495 5404
rect 4500 5398 4515 5404
rect 4374 5360 4380 5367
rect 4365 5356 4380 5360
rect 4394 5356 4400 5387
rect 4491 5384 4495 5398
rect 4511 5384 4515 5398
rect 4531 5384 4535 5441
rect 4631 5439 4635 5496
rect 4731 5471 4735 5476
rect 4626 5427 4635 5439
rect 4365 5344 4369 5356
rect 4385 5352 4400 5356
rect 4385 5344 4389 5352
rect 4631 5344 4635 5427
rect 4722 5464 4735 5471
rect 4722 5419 4726 5464
rect 4751 5453 4755 5476
rect 4746 5441 4755 5453
rect 4722 5396 4726 5407
rect 4722 5388 4740 5396
rect 4736 5384 4740 5388
rect 4744 5384 4748 5441
rect 4771 5399 4775 5476
rect 4831 5408 4835 5476
rect 4853 5447 4857 5496
rect 4863 5475 4867 5496
rect 4883 5484 4887 5496
rect 4891 5492 4895 5496
rect 4891 5488 4925 5492
rect 4883 5480 4913 5484
rect 4883 5479 4901 5480
rect 4863 5471 4887 5475
rect 4766 5387 4773 5399
rect 4831 5396 4833 5408
rect 4766 5344 4770 5387
rect 4831 5384 4835 5396
rect 4853 5389 4857 5435
rect 4849 5383 4857 5389
rect 4849 5354 4853 5383
rect 4881 5376 4887 5471
rect 4849 5347 4857 5354
rect 4853 5324 4857 5347
rect 4861 5324 4865 5364
rect 4881 5344 4885 5376
rect 4921 5362 4925 5488
rect 4937 5382 4941 5496
rect 4959 5484 4963 5496
rect 4961 5472 4963 5484
rect 4969 5484 4973 5496
rect 4969 5472 4971 5484
rect 4889 5350 4913 5352
rect 4889 5348 4925 5350
rect 4889 5344 4893 5348
rect 4935 5344 4939 5370
rect 4953 5362 4957 5472
rect 4991 5464 4995 5496
rect 4962 5460 4995 5464
rect 4962 5396 4966 5460
rect 4982 5411 4986 5440
rect 5001 5438 5005 5496
rect 5021 5439 5025 5476
rect 5111 5439 5115 5496
rect 5106 5427 5115 5439
rect 4982 5403 4991 5411
rect 4962 5384 4965 5396
rect 4955 5344 4959 5350
rect 4967 5344 4971 5384
rect 4987 5344 4991 5403
rect 5001 5344 5005 5426
rect 5021 5384 5025 5427
rect 5111 5344 5115 5427
rect 5171 5408 5175 5476
rect 5193 5447 5197 5496
rect 5203 5475 5207 5496
rect 5223 5484 5227 5496
rect 5231 5492 5235 5496
rect 5231 5488 5265 5492
rect 5223 5480 5253 5484
rect 5223 5479 5241 5480
rect 5203 5471 5227 5475
rect 5171 5396 5173 5408
rect 5171 5384 5175 5396
rect 5193 5389 5197 5435
rect 5189 5383 5197 5389
rect 5189 5354 5193 5383
rect 5221 5376 5227 5471
rect 5189 5347 5197 5354
rect 5193 5324 5197 5347
rect 5201 5324 5205 5364
rect 5221 5344 5225 5376
rect 5261 5362 5265 5488
rect 5277 5382 5281 5496
rect 5299 5484 5303 5496
rect 5301 5472 5303 5484
rect 5309 5484 5313 5496
rect 5309 5472 5311 5484
rect 5229 5350 5253 5352
rect 5229 5348 5265 5350
rect 5229 5344 5233 5348
rect 5275 5344 5279 5370
rect 5293 5362 5297 5472
rect 5331 5464 5335 5496
rect 5302 5460 5335 5464
rect 5302 5396 5306 5460
rect 5322 5411 5326 5440
rect 5341 5438 5345 5496
rect 5361 5439 5365 5476
rect 5451 5471 5455 5476
rect 5442 5464 5455 5471
rect 5322 5403 5331 5411
rect 5302 5384 5305 5396
rect 5295 5344 5299 5350
rect 5307 5344 5311 5384
rect 5327 5344 5331 5403
rect 5341 5344 5345 5426
rect 5361 5384 5365 5427
rect 5442 5419 5446 5464
rect 5471 5453 5475 5476
rect 5466 5441 5475 5453
rect 5442 5396 5446 5407
rect 5442 5388 5460 5396
rect 5456 5384 5460 5388
rect 5464 5384 5468 5441
rect 5491 5399 5495 5476
rect 5613 5456 5617 5476
rect 5609 5449 5617 5456
rect 5623 5456 5627 5476
rect 5733 5456 5737 5476
rect 5623 5449 5637 5456
rect 5609 5433 5615 5449
rect 5606 5421 5615 5433
rect 5486 5387 5493 5399
rect 5486 5344 5490 5387
rect 5611 5344 5615 5421
rect 5631 5433 5637 5449
rect 5729 5449 5737 5456
rect 5743 5456 5747 5476
rect 5743 5449 5757 5456
rect 5729 5433 5735 5449
rect 5631 5421 5634 5433
rect 5726 5421 5735 5433
rect 5631 5344 5635 5421
rect 5731 5344 5735 5421
rect 5751 5433 5757 5449
rect 5751 5421 5754 5433
rect 5751 5344 5755 5421
rect 90 5300 94 5304
rect 112 5300 116 5304
rect 120 5300 124 5304
rect 245 5300 249 5304
rect 265 5300 269 5304
rect 285 5300 289 5304
rect 385 5300 389 5304
rect 405 5300 409 5304
rect 425 5300 429 5304
rect 525 5300 529 5304
rect 545 5300 549 5304
rect 565 5300 569 5304
rect 671 5300 675 5304
rect 691 5300 695 5304
rect 711 5300 715 5304
rect 816 5300 820 5304
rect 824 5300 828 5304
rect 846 5300 850 5304
rect 951 5300 955 5304
rect 971 5300 975 5304
rect 991 5300 995 5304
rect 1105 5300 1109 5304
rect 1125 5300 1129 5304
rect 1145 5300 1149 5304
rect 1231 5300 1235 5304
rect 1251 5300 1255 5304
rect 1271 5300 1275 5304
rect 1391 5300 1395 5304
rect 1399 5300 1403 5304
rect 1525 5300 1529 5304
rect 1545 5300 1549 5304
rect 1565 5300 1569 5304
rect 1656 5300 1660 5304
rect 1664 5300 1668 5304
rect 1686 5300 1690 5304
rect 1805 5300 1809 5304
rect 1825 5300 1829 5304
rect 1845 5300 1849 5304
rect 1945 5300 1949 5304
rect 1965 5300 1969 5304
rect 1985 5300 1989 5304
rect 2071 5300 2075 5304
rect 2091 5300 2095 5304
rect 2225 5300 2229 5304
rect 2321 5300 2325 5304
rect 2343 5300 2347 5304
rect 2365 5300 2369 5304
rect 2456 5300 2460 5304
rect 2464 5300 2468 5304
rect 2486 5300 2490 5304
rect 2625 5300 2629 5304
rect 2645 5300 2649 5304
rect 2665 5300 2669 5304
rect 2765 5300 2769 5304
rect 2785 5300 2789 5304
rect 2805 5300 2809 5304
rect 2896 5300 2900 5304
rect 2904 5300 2908 5304
rect 2926 5300 2930 5304
rect 3031 5300 3035 5304
rect 3131 5300 3135 5304
rect 3151 5300 3155 5304
rect 3271 5300 3275 5304
rect 3291 5300 3295 5304
rect 3311 5300 3315 5304
rect 3411 5300 3415 5304
rect 3431 5300 3435 5304
rect 3531 5300 3535 5304
rect 3541 5300 3545 5304
rect 3561 5300 3565 5304
rect 3685 5300 3689 5304
rect 3705 5300 3709 5304
rect 3725 5300 3729 5304
rect 3825 5300 3829 5304
rect 3845 5300 3849 5304
rect 3865 5300 3869 5304
rect 3951 5300 3955 5304
rect 3971 5300 3975 5304
rect 4090 5300 4094 5304
rect 4112 5300 4116 5304
rect 4120 5300 4124 5304
rect 4225 5300 4229 5304
rect 4245 5300 4249 5304
rect 4345 5300 4349 5304
rect 4365 5300 4369 5304
rect 4385 5300 4389 5304
rect 4491 5300 4495 5304
rect 4511 5300 4515 5304
rect 4531 5300 4535 5304
rect 4631 5300 4635 5304
rect 4736 5300 4740 5304
rect 4744 5300 4748 5304
rect 4766 5300 4770 5304
rect 4831 5300 4835 5304
rect 4853 5300 4857 5304
rect 4861 5300 4865 5304
rect 4881 5300 4885 5304
rect 4889 5300 4893 5304
rect 4935 5300 4939 5304
rect 4955 5300 4959 5304
rect 4967 5300 4971 5304
rect 4987 5300 4991 5304
rect 5001 5300 5005 5304
rect 5021 5300 5025 5304
rect 5111 5300 5115 5304
rect 5171 5300 5175 5304
rect 5193 5300 5197 5304
rect 5201 5300 5205 5304
rect 5221 5300 5225 5304
rect 5229 5300 5233 5304
rect 5275 5300 5279 5304
rect 5295 5300 5299 5304
rect 5307 5300 5311 5304
rect 5327 5300 5331 5304
rect 5341 5300 5345 5304
rect 5361 5300 5365 5304
rect 5456 5300 5460 5304
rect 5464 5300 5468 5304
rect 5486 5300 5490 5304
rect 5611 5300 5615 5304
rect 5631 5300 5635 5304
rect 5731 5300 5735 5304
rect 5751 5300 5755 5304
rect 85 5276 89 5280
rect 105 5276 109 5280
rect 125 5276 129 5280
rect 211 5276 215 5280
rect 231 5276 235 5280
rect 251 5276 255 5280
rect 351 5276 355 5280
rect 465 5276 469 5280
rect 485 5276 489 5280
rect 505 5276 509 5280
rect 591 5276 595 5280
rect 611 5276 615 5280
rect 631 5276 635 5280
rect 745 5276 749 5280
rect 765 5276 769 5280
rect 785 5276 789 5280
rect 871 5276 875 5280
rect 891 5276 895 5280
rect 911 5276 915 5280
rect 1025 5276 1029 5280
rect 1045 5276 1049 5280
rect 1065 5276 1069 5280
rect 1151 5276 1155 5280
rect 1265 5276 1269 5280
rect 1285 5276 1289 5280
rect 1305 5276 1309 5280
rect 1430 5276 1434 5280
rect 1452 5276 1456 5280
rect 1460 5276 1464 5280
rect 1565 5276 1569 5280
rect 1670 5276 1674 5280
rect 1692 5276 1696 5280
rect 1700 5276 1704 5280
rect 1885 5276 1889 5280
rect 1905 5276 1909 5280
rect 1925 5276 1929 5280
rect 1945 5276 1949 5280
rect 2045 5276 2049 5280
rect 2065 5276 2069 5280
rect 2085 5276 2089 5280
rect 2105 5276 2109 5280
rect 2191 5276 2195 5280
rect 2211 5276 2215 5280
rect 2325 5276 2329 5280
rect 2345 5276 2349 5280
rect 2365 5276 2369 5280
rect 2465 5276 2469 5280
rect 2485 5276 2489 5280
rect 2505 5276 2509 5280
rect 2605 5276 2609 5280
rect 2710 5276 2714 5280
rect 2732 5276 2736 5280
rect 2740 5276 2744 5280
rect 2870 5276 2874 5280
rect 2892 5276 2896 5280
rect 2900 5276 2904 5280
rect 3001 5276 3005 5280
rect 3023 5276 3027 5280
rect 3045 5276 3049 5280
rect 3131 5276 3135 5280
rect 3139 5276 3143 5280
rect 3285 5276 3289 5280
rect 3397 5276 3401 5280
rect 3405 5276 3409 5280
rect 3530 5276 3534 5280
rect 3552 5276 3556 5280
rect 3560 5276 3564 5280
rect 3651 5276 3655 5280
rect 3671 5276 3675 5280
rect 3785 5276 3789 5280
rect 3805 5276 3809 5280
rect 3925 5276 3929 5280
rect 3945 5276 3949 5280
rect 4031 5276 4035 5280
rect 4051 5276 4055 5280
rect 4071 5276 4075 5280
rect 4190 5276 4194 5280
rect 4212 5276 4216 5280
rect 4220 5276 4224 5280
rect 4336 5276 4340 5280
rect 4344 5276 4348 5280
rect 4366 5276 4370 5280
rect 4471 5276 4475 5280
rect 4585 5276 4589 5280
rect 4605 5276 4609 5280
rect 4625 5276 4629 5280
rect 4711 5276 4715 5280
rect 4731 5276 4735 5280
rect 4751 5276 4755 5280
rect 4851 5276 4855 5280
rect 4859 5276 4863 5280
rect 4931 5276 4935 5280
rect 4953 5276 4957 5280
rect 4961 5276 4965 5280
rect 4981 5276 4985 5280
rect 4989 5276 4993 5280
rect 5035 5276 5039 5280
rect 5055 5276 5059 5280
rect 5067 5276 5071 5280
rect 5087 5276 5091 5280
rect 5101 5276 5105 5280
rect 5121 5276 5125 5280
rect 5216 5276 5220 5280
rect 5224 5276 5228 5280
rect 5246 5276 5250 5280
rect 5351 5276 5355 5280
rect 5456 5276 5460 5280
rect 5464 5276 5468 5280
rect 5486 5276 5490 5280
rect 5605 5276 5609 5280
rect 5625 5276 5629 5280
rect 5711 5276 5715 5280
rect 5731 5276 5735 5280
rect 85 5193 89 5236
rect 105 5224 109 5236
rect 125 5228 129 5236
rect 125 5224 140 5228
rect 105 5220 120 5224
rect 114 5213 120 5220
rect 85 5181 93 5193
rect 105 5181 112 5193
rect 108 5124 112 5181
rect 116 5124 120 5201
rect 134 5193 140 5224
rect 124 5181 134 5193
rect 211 5182 215 5196
rect 231 5182 235 5196
rect 124 5124 128 5181
rect 199 5176 215 5182
rect 220 5176 235 5182
rect 199 5139 206 5176
rect 220 5153 226 5176
rect 199 5114 206 5127
rect 199 5108 218 5114
rect 214 5104 218 5108
rect 222 5104 226 5141
rect 251 5139 255 5196
rect 351 5153 355 5236
rect 465 5193 469 5236
rect 485 5224 489 5236
rect 505 5228 509 5236
rect 505 5224 520 5228
rect 485 5220 500 5224
rect 494 5213 500 5220
rect 465 5181 473 5193
rect 485 5181 492 5193
rect 346 5141 355 5153
rect 246 5127 255 5139
rect 244 5084 248 5127
rect 351 5084 355 5141
rect 488 5124 492 5181
rect 496 5124 500 5201
rect 514 5193 520 5224
rect 871 5228 875 5236
rect 860 5224 875 5228
rect 891 5224 895 5236
rect 504 5181 514 5193
rect 591 5182 595 5196
rect 611 5182 615 5196
rect 504 5124 508 5181
rect 579 5176 595 5182
rect 600 5176 615 5182
rect 579 5139 586 5176
rect 600 5153 606 5176
rect 579 5114 586 5127
rect 579 5108 598 5114
rect 594 5104 598 5108
rect 602 5104 606 5141
rect 631 5139 635 5196
rect 626 5127 635 5139
rect 745 5139 749 5196
rect 765 5182 769 5196
rect 785 5182 789 5196
rect 860 5193 866 5224
rect 880 5220 895 5224
rect 880 5213 886 5220
rect 765 5176 780 5182
rect 785 5176 801 5182
rect 866 5181 876 5193
rect 774 5153 780 5176
rect 745 5127 754 5139
rect 624 5084 628 5127
rect 752 5084 756 5127
rect 774 5104 778 5141
rect 794 5139 801 5176
rect 794 5114 801 5127
rect 872 5124 876 5181
rect 880 5124 884 5201
rect 911 5193 915 5236
rect 888 5181 895 5193
rect 907 5181 915 5193
rect 1025 5193 1029 5236
rect 1045 5224 1049 5236
rect 1065 5228 1069 5236
rect 1065 5224 1080 5228
rect 1045 5220 1060 5224
rect 1054 5213 1060 5220
rect 1025 5181 1033 5193
rect 1045 5181 1052 5193
rect 888 5124 892 5181
rect 1048 5124 1052 5181
rect 1056 5124 1060 5201
rect 1074 5193 1080 5224
rect 1064 5181 1074 5193
rect 1064 5124 1068 5181
rect 1151 5153 1155 5236
rect 1265 5193 1269 5236
rect 1285 5224 1289 5236
rect 1305 5228 1309 5236
rect 1305 5224 1320 5228
rect 1285 5220 1300 5224
rect 1294 5213 1300 5220
rect 1265 5181 1273 5193
rect 1285 5181 1292 5193
rect 1146 5141 1155 5153
rect 782 5108 801 5114
rect 782 5104 786 5108
rect 1151 5084 1155 5141
rect 1288 5124 1292 5181
rect 1296 5124 1300 5201
rect 1314 5193 1320 5224
rect 1430 5193 1434 5236
rect 1304 5181 1314 5193
rect 1427 5181 1434 5193
rect 1304 5124 1308 5181
rect 1425 5104 1429 5181
rect 1452 5139 1456 5196
rect 1460 5192 1464 5196
rect 1460 5184 1478 5192
rect 1474 5173 1478 5184
rect 1445 5127 1454 5139
rect 1445 5104 1449 5127
rect 1474 5116 1478 5161
rect 1465 5109 1478 5116
rect 1565 5153 1569 5236
rect 1670 5193 1674 5236
rect 1821 5268 1825 5272
rect 1841 5268 1845 5272
rect 1885 5212 1889 5216
rect 1905 5212 1909 5216
rect 1885 5208 1909 5212
rect 1821 5200 1825 5208
rect 1841 5200 1845 5208
rect 1821 5196 1871 5200
rect 1667 5181 1674 5193
rect 1565 5141 1574 5153
rect 1465 5104 1469 5109
rect 1565 5084 1569 5141
rect 1665 5104 1669 5181
rect 1692 5139 1696 5196
rect 1700 5192 1704 5196
rect 1700 5184 1718 5192
rect 1714 5173 1718 5184
rect 1865 5173 1871 5196
rect 1865 5161 1874 5173
rect 1685 5127 1694 5139
rect 1685 5104 1689 5127
rect 1714 5116 1718 5161
rect 1705 5109 1718 5116
rect 1705 5104 1709 5109
rect 1865 5106 1871 5161
rect 1905 5139 1909 5208
rect 1906 5127 1909 5139
rect 1865 5100 1889 5106
rect 1885 5084 1889 5100
rect 1905 5084 1909 5127
rect 1925 5212 1929 5216
rect 1945 5212 1949 5216
rect 1925 5208 1949 5212
rect 1925 5173 1929 5208
rect 2045 5173 2049 5196
rect 1925 5161 1934 5173
rect 2046 5161 2049 5173
rect 1925 5084 1929 5161
rect 2040 5113 2046 5161
rect 2065 5139 2069 5196
rect 2085 5174 2089 5196
rect 2105 5174 2109 5196
rect 2085 5168 2098 5174
rect 2105 5173 2125 5174
rect 2105 5168 2113 5173
rect 2094 5139 2098 5168
rect 2067 5127 2069 5139
rect 2065 5125 2069 5127
rect 2065 5118 2078 5125
rect 2040 5109 2070 5113
rect 2066 5104 2070 5109
rect 2074 5104 2078 5118
rect 2094 5104 2098 5127
rect 2113 5119 2119 5161
rect 2191 5159 2195 5236
rect 2186 5147 2195 5159
rect 2189 5131 2195 5147
rect 2211 5159 2215 5236
rect 2325 5193 2329 5236
rect 2345 5224 2349 5236
rect 2365 5228 2369 5236
rect 2365 5224 2380 5228
rect 2345 5220 2360 5224
rect 2354 5213 2360 5220
rect 2325 5181 2333 5193
rect 2345 5181 2352 5193
rect 2211 5147 2214 5159
rect 2211 5131 2217 5147
rect 2189 5124 2197 5131
rect 2102 5112 2119 5119
rect 2102 5104 2106 5112
rect 2193 5104 2197 5124
rect 2203 5124 2217 5131
rect 2348 5124 2352 5181
rect 2356 5124 2360 5201
rect 2374 5193 2380 5224
rect 2364 5181 2374 5193
rect 2364 5124 2368 5181
rect 2465 5139 2469 5196
rect 2485 5182 2489 5196
rect 2505 5182 2509 5196
rect 2485 5176 2500 5182
rect 2505 5176 2521 5182
rect 2494 5153 2500 5176
rect 2465 5127 2474 5139
rect 2203 5104 2207 5124
rect 2472 5084 2476 5127
rect 2494 5104 2498 5141
rect 2514 5139 2521 5176
rect 2605 5153 2609 5236
rect 2710 5193 2714 5236
rect 2707 5181 2714 5193
rect 2605 5141 2614 5153
rect 2514 5114 2521 5127
rect 2502 5108 2521 5114
rect 2502 5104 2506 5108
rect 2605 5084 2609 5141
rect 2705 5104 2709 5181
rect 2732 5139 2736 5196
rect 2740 5192 2744 5196
rect 2870 5193 2874 5236
rect 2740 5184 2758 5192
rect 2754 5173 2758 5184
rect 2867 5181 2874 5193
rect 2725 5127 2734 5139
rect 2725 5104 2729 5127
rect 2754 5116 2758 5161
rect 2745 5109 2758 5116
rect 2745 5104 2749 5109
rect 2865 5104 2869 5181
rect 2892 5139 2896 5196
rect 2900 5192 2904 5196
rect 2900 5184 2918 5192
rect 2914 5173 2918 5184
rect 2885 5127 2894 5139
rect 2885 5104 2889 5127
rect 2914 5116 2918 5161
rect 2905 5109 2918 5116
rect 3001 5122 3005 5196
rect 3023 5159 3027 5236
rect 3045 5173 3049 5236
rect 3131 5173 3135 5196
rect 3045 5161 3054 5173
rect 3126 5161 3135 5173
rect 3139 5173 3143 5196
rect 3139 5161 3154 5173
rect 3026 5147 3039 5159
rect 3001 5110 3013 5122
rect 2905 5104 2909 5109
rect 3015 5104 3019 5110
rect 3035 5104 3039 5147
rect 3045 5104 3049 5161
rect 3131 5084 3135 5161
rect 3151 5084 3155 5161
rect 3285 5153 3289 5236
rect 3397 5173 3401 5196
rect 3386 5161 3401 5173
rect 3405 5173 3409 5196
rect 3530 5193 3534 5236
rect 3527 5181 3534 5193
rect 3405 5161 3414 5173
rect 3285 5141 3294 5153
rect 3285 5084 3289 5141
rect 3385 5084 3389 5161
rect 3405 5084 3409 5161
rect 3525 5104 3529 5181
rect 3552 5139 3556 5196
rect 3560 5192 3564 5196
rect 3560 5184 3578 5192
rect 3574 5173 3578 5184
rect 3545 5127 3554 5139
rect 3545 5104 3549 5127
rect 3574 5116 3578 5161
rect 3651 5159 3655 5236
rect 3646 5147 3655 5159
rect 3649 5131 3655 5147
rect 3671 5159 3675 5236
rect 3785 5159 3789 5236
rect 3671 5147 3674 5159
rect 3786 5147 3789 5159
rect 3671 5131 3677 5147
rect 3649 5124 3657 5131
rect 3565 5109 3578 5116
rect 3565 5104 3569 5109
rect 3653 5104 3657 5124
rect 3663 5124 3677 5131
rect 3783 5131 3789 5147
rect 3805 5159 3809 5236
rect 3925 5159 3929 5236
rect 3805 5147 3814 5159
rect 3926 5147 3929 5159
rect 3805 5131 3811 5147
rect 3783 5124 3797 5131
rect 3663 5104 3667 5124
rect 3793 5104 3797 5124
rect 3803 5124 3811 5131
rect 3923 5131 3929 5147
rect 3945 5159 3949 5236
rect 4031 5228 4035 5236
rect 4020 5224 4035 5228
rect 4051 5224 4055 5236
rect 4020 5193 4026 5224
rect 4040 5220 4055 5224
rect 4040 5213 4046 5220
rect 4026 5181 4036 5193
rect 3945 5147 3954 5159
rect 3945 5131 3951 5147
rect 3923 5124 3937 5131
rect 3803 5104 3807 5124
rect 3933 5104 3937 5124
rect 3943 5124 3951 5131
rect 4032 5124 4036 5181
rect 4040 5124 4044 5201
rect 4071 5193 4075 5236
rect 4190 5193 4194 5236
rect 4048 5181 4055 5193
rect 4067 5181 4075 5193
rect 4187 5181 4194 5193
rect 4048 5124 4052 5181
rect 3943 5104 3947 5124
rect 4185 5104 4189 5181
rect 4212 5139 4216 5196
rect 4220 5192 4224 5196
rect 4336 5192 4340 5196
rect 4220 5184 4238 5192
rect 4234 5173 4238 5184
rect 4322 5184 4340 5192
rect 4322 5173 4326 5184
rect 4205 5127 4214 5139
rect 4205 5104 4209 5127
rect 4234 5116 4238 5161
rect 4225 5109 4238 5116
rect 4322 5116 4326 5161
rect 4344 5139 4348 5196
rect 4366 5193 4370 5236
rect 4366 5181 4373 5193
rect 4346 5127 4355 5139
rect 4322 5109 4335 5116
rect 4225 5104 4229 5109
rect 4331 5104 4335 5109
rect 4351 5104 4355 5127
rect 4371 5104 4375 5181
rect 4471 5153 4475 5236
rect 4585 5193 4589 5236
rect 4605 5224 4609 5236
rect 4625 5228 4629 5236
rect 4625 5224 4640 5228
rect 4605 5220 4620 5224
rect 4614 5213 4620 5220
rect 4585 5181 4593 5193
rect 4605 5181 4612 5193
rect 4466 5141 4475 5153
rect 4471 5084 4475 5141
rect 4608 5124 4612 5181
rect 4616 5124 4620 5201
rect 4634 5193 4640 5224
rect 4953 5233 4957 5256
rect 4949 5226 4957 5233
rect 4949 5197 4953 5226
rect 4961 5216 4965 5256
rect 4981 5204 4985 5236
rect 4989 5232 4993 5236
rect 4989 5230 5025 5232
rect 4989 5228 5013 5230
rect 4624 5181 4634 5193
rect 4711 5182 4715 5196
rect 4731 5182 4735 5196
rect 4624 5124 4628 5181
rect 4699 5176 4715 5182
rect 4720 5176 4735 5182
rect 4699 5139 4706 5176
rect 4720 5153 4726 5176
rect 4699 5114 4706 5127
rect 4699 5108 4718 5114
rect 4714 5104 4718 5108
rect 4722 5104 4726 5141
rect 4751 5139 4755 5196
rect 4851 5173 4855 5196
rect 4846 5161 4855 5173
rect 4859 5173 4863 5196
rect 4931 5184 4935 5196
rect 4949 5191 4957 5197
rect 4859 5161 4874 5173
rect 4931 5172 4933 5184
rect 4746 5127 4755 5139
rect 4744 5084 4748 5127
rect 4851 5084 4855 5161
rect 4871 5084 4875 5161
rect 4931 5104 4935 5172
rect 4953 5145 4957 5191
rect 4953 5084 4957 5133
rect 4981 5109 4987 5204
rect 4963 5105 4987 5109
rect 4963 5084 4967 5105
rect 4983 5100 5001 5101
rect 4983 5096 5013 5100
rect 4983 5084 4987 5096
rect 5021 5092 5025 5218
rect 5035 5210 5039 5236
rect 5055 5230 5059 5236
rect 4991 5088 5025 5092
rect 4991 5084 4995 5088
rect 5037 5084 5041 5198
rect 5053 5108 5057 5218
rect 5067 5196 5071 5236
rect 5062 5184 5065 5196
rect 5062 5120 5066 5184
rect 5087 5177 5091 5236
rect 5082 5169 5091 5177
rect 5082 5140 5086 5169
rect 5101 5154 5105 5236
rect 5121 5153 5125 5196
rect 5216 5192 5220 5196
rect 5202 5184 5220 5192
rect 5202 5173 5206 5184
rect 5062 5116 5095 5120
rect 5061 5096 5063 5108
rect 5059 5084 5063 5096
rect 5069 5096 5071 5108
rect 5069 5084 5073 5096
rect 5091 5084 5095 5116
rect 5101 5084 5105 5142
rect 5121 5104 5125 5141
rect 5202 5116 5206 5161
rect 5224 5139 5228 5196
rect 5246 5193 5250 5236
rect 5246 5181 5253 5193
rect 5226 5127 5235 5139
rect 5202 5109 5215 5116
rect 5211 5104 5215 5109
rect 5231 5104 5235 5127
rect 5251 5104 5255 5181
rect 5351 5153 5355 5236
rect 5456 5192 5460 5196
rect 5442 5184 5460 5192
rect 5442 5173 5446 5184
rect 5346 5141 5355 5153
rect 5351 5084 5355 5141
rect 5442 5116 5446 5161
rect 5464 5139 5468 5196
rect 5486 5193 5490 5236
rect 5486 5181 5493 5193
rect 5466 5127 5475 5139
rect 5442 5109 5455 5116
rect 5451 5104 5455 5109
rect 5471 5104 5475 5127
rect 5491 5104 5495 5181
rect 5605 5159 5609 5236
rect 5606 5147 5609 5159
rect 5603 5131 5609 5147
rect 5625 5159 5629 5236
rect 5711 5159 5715 5236
rect 5625 5147 5634 5159
rect 5706 5147 5715 5159
rect 5625 5131 5631 5147
rect 5603 5124 5617 5131
rect 5613 5104 5617 5124
rect 5623 5124 5631 5131
rect 5709 5131 5715 5147
rect 5731 5159 5735 5236
rect 5731 5147 5734 5159
rect 5731 5131 5737 5147
rect 5709 5124 5717 5131
rect 5623 5104 5627 5124
rect 5713 5104 5717 5124
rect 5723 5124 5737 5131
rect 5723 5104 5727 5124
rect 108 5060 112 5064
rect 116 5060 120 5064
rect 124 5060 128 5064
rect 214 5060 218 5064
rect 222 5060 226 5064
rect 244 5060 248 5064
rect 351 5060 355 5064
rect 488 5060 492 5064
rect 496 5060 500 5064
rect 504 5060 508 5064
rect 594 5060 598 5064
rect 602 5060 606 5064
rect 624 5060 628 5064
rect 752 5060 756 5064
rect 774 5060 778 5064
rect 782 5060 786 5064
rect 872 5060 876 5064
rect 880 5060 884 5064
rect 888 5060 892 5064
rect 1048 5060 1052 5064
rect 1056 5060 1060 5064
rect 1064 5060 1068 5064
rect 1151 5060 1155 5064
rect 1288 5060 1292 5064
rect 1296 5060 1300 5064
rect 1304 5060 1308 5064
rect 1425 5060 1429 5064
rect 1445 5060 1449 5064
rect 1465 5060 1469 5064
rect 1565 5060 1569 5064
rect 1665 5060 1669 5064
rect 1685 5060 1689 5064
rect 1705 5060 1709 5064
rect 1885 5060 1889 5064
rect 1905 5060 1909 5064
rect 1925 5060 1929 5064
rect 2066 5060 2070 5064
rect 2074 5060 2078 5064
rect 2094 5060 2098 5064
rect 2102 5060 2106 5064
rect 2193 5060 2197 5064
rect 2203 5060 2207 5064
rect 2348 5060 2352 5064
rect 2356 5060 2360 5064
rect 2364 5060 2368 5064
rect 2472 5060 2476 5064
rect 2494 5060 2498 5064
rect 2502 5060 2506 5064
rect 2605 5060 2609 5064
rect 2705 5060 2709 5064
rect 2725 5060 2729 5064
rect 2745 5060 2749 5064
rect 2865 5060 2869 5064
rect 2885 5060 2889 5064
rect 2905 5060 2909 5064
rect 3015 5060 3019 5064
rect 3035 5060 3039 5064
rect 3045 5060 3049 5064
rect 3131 5060 3135 5064
rect 3151 5060 3155 5064
rect 3285 5060 3289 5064
rect 3385 5060 3389 5064
rect 3405 5060 3409 5064
rect 3525 5060 3529 5064
rect 3545 5060 3549 5064
rect 3565 5060 3569 5064
rect 3653 5060 3657 5064
rect 3663 5060 3667 5064
rect 3793 5060 3797 5064
rect 3803 5060 3807 5064
rect 3933 5060 3937 5064
rect 3943 5060 3947 5064
rect 4032 5060 4036 5064
rect 4040 5060 4044 5064
rect 4048 5060 4052 5064
rect 4185 5060 4189 5064
rect 4205 5060 4209 5064
rect 4225 5060 4229 5064
rect 4331 5060 4335 5064
rect 4351 5060 4355 5064
rect 4371 5060 4375 5064
rect 4471 5060 4475 5064
rect 4608 5060 4612 5064
rect 4616 5060 4620 5064
rect 4624 5060 4628 5064
rect 4714 5060 4718 5064
rect 4722 5060 4726 5064
rect 4744 5060 4748 5064
rect 4851 5060 4855 5064
rect 4871 5060 4875 5064
rect 4931 5060 4935 5064
rect 4953 5060 4957 5064
rect 4963 5060 4967 5064
rect 4983 5060 4987 5064
rect 4991 5060 4995 5064
rect 5037 5060 5041 5064
rect 5059 5060 5063 5064
rect 5069 5060 5073 5064
rect 5091 5060 5095 5064
rect 5101 5060 5105 5064
rect 5121 5060 5125 5064
rect 5211 5060 5215 5064
rect 5231 5060 5235 5064
rect 5251 5060 5255 5064
rect 5351 5060 5355 5064
rect 5451 5060 5455 5064
rect 5471 5060 5475 5064
rect 5491 5060 5495 5064
rect 5613 5060 5617 5064
rect 5623 5060 5627 5064
rect 5713 5060 5717 5064
rect 5723 5060 5727 5064
rect 85 5036 89 5040
rect 105 5036 109 5040
rect 125 5036 129 5040
rect 248 5036 252 5040
rect 256 5036 260 5040
rect 264 5036 268 5040
rect 352 5036 356 5040
rect 360 5036 364 5040
rect 368 5036 372 5040
rect 491 5036 495 5040
rect 511 5036 515 5040
rect 531 5036 535 5040
rect 653 5036 657 5040
rect 663 5036 667 5040
rect 765 5036 769 5040
rect 785 5036 789 5040
rect 805 5036 809 5040
rect 905 5036 909 5040
rect 925 5036 929 5040
rect 945 5036 949 5040
rect 1052 5036 1056 5040
rect 1074 5036 1078 5040
rect 1082 5036 1086 5040
rect 1185 5036 1189 5040
rect 1205 5036 1209 5040
rect 1225 5036 1229 5040
rect 1325 5036 1329 5040
rect 1433 5036 1437 5040
rect 1443 5036 1447 5040
rect 1588 5036 1592 5040
rect 1596 5036 1600 5040
rect 1604 5036 1608 5040
rect 1705 5036 1709 5040
rect 1725 5036 1729 5040
rect 1745 5036 1749 5040
rect 1834 5036 1838 5040
rect 1842 5036 1846 5040
rect 1864 5036 1868 5040
rect 1973 5036 1977 5040
rect 1983 5036 1987 5040
rect 2112 5036 2116 5040
rect 2134 5036 2138 5040
rect 2142 5036 2146 5040
rect 2265 5036 2269 5040
rect 2365 5036 2369 5040
rect 2385 5036 2389 5040
rect 2405 5036 2409 5040
rect 2528 5036 2532 5040
rect 2536 5036 2540 5040
rect 2544 5036 2548 5040
rect 2645 5036 2649 5040
rect 2773 5036 2777 5040
rect 2783 5036 2787 5040
rect 2871 5036 2875 5040
rect 2972 5036 2976 5040
rect 2980 5036 2984 5040
rect 2988 5036 2992 5040
rect 3125 5036 3129 5040
rect 3145 5036 3149 5040
rect 3165 5036 3169 5040
rect 3265 5036 3269 5040
rect 3285 5036 3289 5040
rect 3305 5036 3309 5040
rect 3412 5036 3416 5040
rect 3434 5036 3438 5040
rect 3442 5036 3446 5040
rect 3531 5036 3535 5040
rect 3551 5036 3555 5040
rect 3571 5036 3575 5040
rect 3685 5036 3689 5040
rect 3705 5036 3709 5040
rect 3828 5036 3832 5040
rect 3836 5036 3840 5040
rect 3844 5036 3848 5040
rect 3945 5036 3949 5040
rect 4032 5036 4036 5040
rect 4040 5036 4044 5040
rect 4048 5036 4052 5040
rect 4172 5036 4176 5040
rect 4180 5036 4184 5040
rect 4188 5036 4192 5040
rect 4335 5036 4339 5040
rect 4355 5036 4359 5040
rect 4365 5036 4369 5040
rect 4471 5036 4475 5040
rect 4491 5036 4495 5040
rect 4511 5036 4515 5040
rect 4611 5036 4615 5040
rect 4631 5036 4635 5040
rect 4745 5036 4749 5040
rect 4765 5036 4769 5040
rect 4785 5036 4789 5040
rect 4831 5036 4835 5040
rect 4853 5036 4857 5040
rect 4863 5036 4867 5040
rect 4883 5036 4887 5040
rect 4891 5036 4895 5040
rect 4937 5036 4941 5040
rect 4959 5036 4963 5040
rect 4969 5036 4973 5040
rect 4991 5036 4995 5040
rect 5001 5036 5005 5040
rect 5021 5036 5025 5040
rect 5111 5036 5115 5040
rect 5131 5036 5135 5040
rect 5151 5036 5155 5040
rect 5211 5036 5215 5040
rect 5233 5036 5237 5040
rect 5243 5036 5247 5040
rect 5263 5036 5267 5040
rect 5271 5036 5275 5040
rect 5317 5036 5321 5040
rect 5339 5036 5343 5040
rect 5349 5036 5353 5040
rect 5371 5036 5375 5040
rect 5381 5036 5385 5040
rect 5401 5036 5405 5040
rect 5513 5036 5517 5040
rect 5523 5036 5527 5040
rect 5613 5036 5617 5040
rect 5623 5036 5627 5040
rect 5753 5036 5757 5040
rect 5763 5036 5767 5040
rect 85 4919 89 4996
rect 105 4973 109 4996
rect 125 4991 129 4996
rect 125 4984 138 4991
rect 105 4961 114 4973
rect 87 4907 94 4919
rect 90 4864 94 4907
rect 112 4904 116 4961
rect 134 4939 138 4984
rect 491 4991 495 4996
rect 482 4984 495 4991
rect 134 4916 138 4927
rect 248 4919 252 4976
rect 120 4908 138 4916
rect 120 4904 124 4908
rect 225 4907 233 4919
rect 245 4907 252 4919
rect 225 4864 229 4907
rect 256 4899 260 4976
rect 264 4919 268 4976
rect 352 4919 356 4976
rect 264 4907 274 4919
rect 346 4907 356 4919
rect 254 4880 260 4887
rect 245 4876 260 4880
rect 274 4876 280 4907
rect 245 4864 249 4876
rect 265 4872 280 4876
rect 340 4876 346 4907
rect 360 4899 364 4976
rect 368 4919 372 4976
rect 482 4939 486 4984
rect 511 4973 515 4996
rect 506 4961 515 4973
rect 368 4907 375 4919
rect 387 4907 395 4919
rect 482 4916 486 4927
rect 482 4908 500 4916
rect 360 4880 366 4887
rect 360 4876 375 4880
rect 340 4872 355 4876
rect 265 4864 269 4872
rect 351 4864 355 4872
rect 371 4864 375 4876
rect 391 4864 395 4907
rect 496 4904 500 4908
rect 504 4904 508 4961
rect 531 4919 535 4996
rect 653 4976 657 4996
rect 643 4969 657 4976
rect 663 4976 667 4996
rect 663 4969 671 4976
rect 643 4953 649 4969
rect 646 4941 649 4953
rect 526 4907 533 4919
rect 526 4864 530 4907
rect 645 4864 649 4941
rect 665 4953 671 4969
rect 665 4941 674 4953
rect 665 4864 669 4941
rect 765 4919 769 4996
rect 785 4973 789 4996
rect 805 4991 809 4996
rect 805 4984 818 4991
rect 785 4961 794 4973
rect 767 4907 774 4919
rect 770 4864 774 4907
rect 792 4904 796 4961
rect 814 4939 818 4984
rect 814 4916 818 4927
rect 905 4919 909 4996
rect 925 4973 929 4996
rect 945 4991 949 4996
rect 945 4984 958 4991
rect 925 4961 934 4973
rect 800 4908 818 4916
rect 800 4904 804 4908
rect 907 4907 914 4919
rect 910 4864 914 4907
rect 932 4904 936 4961
rect 954 4939 958 4984
rect 1052 4973 1056 5016
rect 1045 4961 1054 4973
rect 954 4916 958 4927
rect 940 4908 958 4916
rect 940 4904 944 4908
rect 1045 4904 1049 4961
rect 1074 4959 1078 4996
rect 1082 4992 1086 4996
rect 1082 4986 1101 4992
rect 1094 4973 1101 4986
rect 1074 4924 1080 4947
rect 1094 4924 1101 4961
rect 1065 4918 1080 4924
rect 1085 4918 1101 4924
rect 1185 4919 1189 4996
rect 1205 4973 1209 4996
rect 1225 4991 1229 4996
rect 1225 4984 1238 4991
rect 1205 4961 1214 4973
rect 1065 4904 1069 4918
rect 1085 4904 1089 4918
rect 1187 4907 1194 4919
rect 1190 4864 1194 4907
rect 1212 4904 1216 4961
rect 1234 4939 1238 4984
rect 1325 4959 1329 5016
rect 1433 4976 1437 4996
rect 1423 4969 1437 4976
rect 1443 4976 1447 4996
rect 1443 4969 1451 4976
rect 1325 4947 1334 4959
rect 1423 4953 1429 4969
rect 1234 4916 1238 4927
rect 1220 4908 1238 4916
rect 1220 4904 1224 4908
rect 1325 4864 1329 4947
rect 1426 4941 1429 4953
rect 1425 4864 1429 4941
rect 1445 4953 1451 4969
rect 1445 4941 1454 4953
rect 1445 4864 1449 4941
rect 1588 4919 1592 4976
rect 1565 4907 1573 4919
rect 1585 4907 1592 4919
rect 1565 4864 1569 4907
rect 1596 4899 1600 4976
rect 1604 4919 1608 4976
rect 1705 4919 1709 4996
rect 1725 4973 1729 4996
rect 1745 4991 1749 4996
rect 1834 4992 1838 4996
rect 1745 4984 1758 4991
rect 1725 4961 1734 4973
rect 1604 4907 1614 4919
rect 1707 4907 1714 4919
rect 1594 4880 1600 4887
rect 1585 4876 1600 4880
rect 1614 4876 1620 4907
rect 1585 4864 1589 4876
rect 1605 4872 1620 4876
rect 1605 4864 1609 4872
rect 1710 4864 1714 4907
rect 1732 4904 1736 4961
rect 1754 4939 1758 4984
rect 1819 4986 1838 4992
rect 1819 4973 1826 4986
rect 1754 4916 1758 4927
rect 1819 4924 1826 4961
rect 1842 4959 1846 4996
rect 1864 4973 1868 5016
rect 1973 4976 1977 4996
rect 1866 4961 1875 4973
rect 1840 4924 1846 4947
rect 1819 4918 1835 4924
rect 1840 4918 1855 4924
rect 1740 4908 1758 4916
rect 1740 4904 1744 4908
rect 1831 4904 1835 4918
rect 1851 4904 1855 4918
rect 1871 4904 1875 4961
rect 1969 4969 1977 4976
rect 1983 4976 1987 4996
rect 1983 4969 1997 4976
rect 2112 4973 2116 5016
rect 1969 4953 1975 4969
rect 1966 4941 1975 4953
rect 1971 4864 1975 4941
rect 1991 4953 1997 4969
rect 2105 4961 2114 4973
rect 1991 4941 1994 4953
rect 1991 4864 1995 4941
rect 2105 4904 2109 4961
rect 2134 4959 2138 4996
rect 2142 4992 2146 4996
rect 2142 4986 2161 4992
rect 2154 4973 2161 4986
rect 2134 4924 2140 4947
rect 2154 4924 2161 4961
rect 2125 4918 2140 4924
rect 2145 4918 2161 4924
rect 2265 4959 2269 5016
rect 2265 4947 2274 4959
rect 2125 4904 2129 4918
rect 2145 4904 2149 4918
rect 2265 4864 2269 4947
rect 2365 4919 2369 4996
rect 2385 4973 2389 4996
rect 2405 4991 2409 4996
rect 2405 4984 2418 4991
rect 2385 4961 2394 4973
rect 2367 4907 2374 4919
rect 2370 4864 2374 4907
rect 2392 4904 2396 4961
rect 2414 4939 2418 4984
rect 2414 4916 2418 4927
rect 2528 4919 2532 4976
rect 2400 4908 2418 4916
rect 2400 4904 2404 4908
rect 2505 4907 2513 4919
rect 2525 4907 2532 4919
rect 2505 4864 2509 4907
rect 2536 4899 2540 4976
rect 2544 4919 2548 4976
rect 2645 4959 2649 5016
rect 2773 4976 2777 4996
rect 2763 4969 2777 4976
rect 2783 4976 2787 4996
rect 2783 4969 2791 4976
rect 2645 4947 2654 4959
rect 2763 4953 2769 4969
rect 2544 4907 2554 4919
rect 2534 4880 2540 4887
rect 2525 4876 2540 4880
rect 2554 4876 2560 4907
rect 2525 4864 2529 4876
rect 2545 4872 2560 4876
rect 2545 4864 2549 4872
rect 2645 4864 2649 4947
rect 2766 4941 2769 4953
rect 2765 4864 2769 4941
rect 2785 4953 2791 4969
rect 2871 4959 2875 5016
rect 2785 4941 2794 4953
rect 2866 4947 2875 4959
rect 2785 4864 2789 4941
rect 2871 4864 2875 4947
rect 2972 4919 2976 4976
rect 2966 4907 2976 4919
rect 2960 4876 2966 4907
rect 2980 4899 2984 4976
rect 2988 4919 2992 4976
rect 3125 4919 3129 4996
rect 3145 4973 3149 4996
rect 3165 4991 3169 4996
rect 3165 4984 3178 4991
rect 3145 4961 3154 4973
rect 2988 4907 2995 4919
rect 3007 4907 3015 4919
rect 3127 4907 3134 4919
rect 2980 4880 2986 4887
rect 2980 4876 2995 4880
rect 2960 4872 2975 4876
rect 2971 4864 2975 4872
rect 2991 4864 2995 4876
rect 3011 4864 3015 4907
rect 3130 4864 3134 4907
rect 3152 4904 3156 4961
rect 3174 4939 3178 4984
rect 3174 4916 3178 4927
rect 3265 4919 3269 4996
rect 3285 4973 3289 4996
rect 3305 4991 3309 4996
rect 3305 4984 3318 4991
rect 3285 4961 3294 4973
rect 3160 4908 3178 4916
rect 3160 4904 3164 4908
rect 3267 4907 3274 4919
rect 3270 4864 3274 4907
rect 3292 4904 3296 4961
rect 3314 4939 3318 4984
rect 3412 4973 3416 5016
rect 3531 5009 3535 5016
rect 3551 5009 3555 5016
rect 3522 5004 3535 5009
rect 3405 4961 3414 4973
rect 3314 4916 3318 4927
rect 3300 4908 3318 4916
rect 3300 4904 3304 4908
rect 3405 4904 3409 4961
rect 3434 4959 3438 4996
rect 3442 4992 3446 4996
rect 3442 4986 3461 4992
rect 3454 4973 3461 4986
rect 3434 4924 3440 4947
rect 3454 4924 3461 4961
rect 3522 4959 3526 5004
rect 3425 4918 3440 4924
rect 3445 4918 3461 4924
rect 3425 4904 3429 4918
rect 3445 4904 3449 4918
rect 3522 4913 3526 4947
rect 3541 5003 3555 5009
rect 3541 4939 3545 5003
rect 3571 4988 3575 4996
rect 3565 4976 3575 4988
rect 3685 4939 3689 5016
rect 3705 4939 3709 5016
rect 3686 4927 3701 4939
rect 3522 4908 3535 4913
rect 3531 4904 3535 4908
rect 3541 4904 3545 4927
rect 3561 4904 3565 4909
rect 3697 4904 3701 4927
rect 3705 4927 3714 4939
rect 3705 4904 3709 4927
rect 3828 4919 3832 4976
rect 3805 4907 3813 4919
rect 3825 4907 3832 4919
rect 3805 4864 3809 4907
rect 3836 4899 3840 4976
rect 3844 4919 3848 4976
rect 3945 4959 3949 5016
rect 4471 5009 4475 5016
rect 4491 5009 4495 5016
rect 4462 5004 4475 5009
rect 4335 4990 4339 4996
rect 4321 4978 4333 4990
rect 3945 4947 3954 4959
rect 3844 4907 3854 4919
rect 3834 4880 3840 4887
rect 3825 4876 3840 4880
rect 3854 4876 3860 4907
rect 3825 4864 3829 4876
rect 3845 4872 3860 4876
rect 3845 4864 3849 4872
rect 3945 4864 3949 4947
rect 4032 4919 4036 4976
rect 4026 4907 4036 4919
rect 4020 4876 4026 4907
rect 4040 4899 4044 4976
rect 4048 4919 4052 4976
rect 4172 4919 4176 4976
rect 4048 4907 4055 4919
rect 4067 4907 4075 4919
rect 4166 4907 4176 4919
rect 4040 4880 4046 4887
rect 4040 4876 4055 4880
rect 4020 4872 4035 4876
rect 4031 4864 4035 4872
rect 4051 4864 4055 4876
rect 4071 4864 4075 4907
rect 4160 4876 4166 4907
rect 4180 4899 4184 4976
rect 4188 4919 4192 4976
rect 4188 4907 4195 4919
rect 4207 4907 4215 4919
rect 4180 4880 4186 4887
rect 4180 4876 4195 4880
rect 4160 4872 4175 4876
rect 4171 4864 4175 4872
rect 4191 4864 4195 4876
rect 4211 4864 4215 4907
rect 4321 4904 4325 4978
rect 4355 4953 4359 4996
rect 4346 4941 4359 4953
rect 4343 4864 4347 4941
rect 4365 4939 4369 4996
rect 4462 4959 4466 5004
rect 4365 4927 4374 4939
rect 4365 4864 4369 4927
rect 4462 4913 4466 4947
rect 4481 5003 4495 5009
rect 4481 4939 4485 5003
rect 4511 4988 4515 4996
rect 4505 4976 4515 4988
rect 4611 4939 4615 5016
rect 4631 4939 4635 5016
rect 4606 4927 4615 4939
rect 4462 4908 4475 4913
rect 4471 4904 4475 4908
rect 4481 4904 4485 4927
rect 4501 4904 4505 4909
rect 4611 4904 4615 4927
rect 4619 4927 4634 4939
rect 4619 4904 4623 4927
rect 4745 4919 4749 4996
rect 4765 4973 4769 4996
rect 4785 4991 4789 4996
rect 4785 4984 4798 4991
rect 4765 4961 4774 4973
rect 4747 4907 4754 4919
rect 4750 4864 4754 4907
rect 4772 4904 4776 4961
rect 4794 4939 4798 4984
rect 4831 4928 4835 4996
rect 4853 4967 4857 5016
rect 4863 4995 4867 5016
rect 4883 5004 4887 5016
rect 4891 5012 4895 5016
rect 4891 5008 4925 5012
rect 4883 5000 4913 5004
rect 4883 4999 4901 5000
rect 4863 4991 4887 4995
rect 4794 4916 4798 4927
rect 4780 4908 4798 4916
rect 4831 4916 4833 4928
rect 4780 4904 4784 4908
rect 4831 4904 4835 4916
rect 4853 4909 4857 4955
rect 4849 4903 4857 4909
rect 4849 4874 4853 4903
rect 4881 4896 4887 4991
rect 4849 4867 4857 4874
rect 4853 4844 4857 4867
rect 4861 4844 4865 4884
rect 4881 4864 4885 4896
rect 4921 4882 4925 5008
rect 4937 4902 4941 5016
rect 4959 5004 4963 5016
rect 4961 4992 4963 5004
rect 4969 5004 4973 5016
rect 4969 4992 4971 5004
rect 4889 4870 4913 4872
rect 4889 4868 4925 4870
rect 4889 4864 4893 4868
rect 4935 4864 4939 4890
rect 4953 4882 4957 4992
rect 4991 4984 4995 5016
rect 4962 4980 4995 4984
rect 4962 4916 4966 4980
rect 4982 4931 4986 4960
rect 5001 4958 5005 5016
rect 5021 4959 5025 4996
rect 5111 4991 5115 4996
rect 5102 4984 5115 4991
rect 4982 4923 4991 4931
rect 4962 4904 4965 4916
rect 4955 4864 4959 4870
rect 4967 4864 4971 4904
rect 4987 4864 4991 4923
rect 5001 4864 5005 4946
rect 5021 4904 5025 4947
rect 5102 4939 5106 4984
rect 5131 4973 5135 4996
rect 5126 4961 5135 4973
rect 5102 4916 5106 4927
rect 5102 4908 5120 4916
rect 5116 4904 5120 4908
rect 5124 4904 5128 4961
rect 5151 4919 5155 4996
rect 5211 4928 5215 4996
rect 5233 4967 5237 5016
rect 5243 4995 5247 5016
rect 5263 5004 5267 5016
rect 5271 5012 5275 5016
rect 5271 5008 5305 5012
rect 5263 5000 5293 5004
rect 5263 4999 5281 5000
rect 5243 4991 5267 4995
rect 5146 4907 5153 4919
rect 5211 4916 5213 4928
rect 5146 4864 5150 4907
rect 5211 4904 5215 4916
rect 5233 4909 5237 4955
rect 5229 4903 5237 4909
rect 5229 4874 5233 4903
rect 5261 4896 5267 4991
rect 5229 4867 5237 4874
rect 5233 4844 5237 4867
rect 5241 4844 5245 4884
rect 5261 4864 5265 4896
rect 5301 4882 5305 5008
rect 5317 4902 5321 5016
rect 5339 5004 5343 5016
rect 5341 4992 5343 5004
rect 5349 5004 5353 5016
rect 5349 4992 5351 5004
rect 5269 4870 5293 4872
rect 5269 4868 5305 4870
rect 5269 4864 5273 4868
rect 5315 4864 5319 4890
rect 5333 4882 5337 4992
rect 5371 4984 5375 5016
rect 5342 4980 5375 4984
rect 5342 4916 5346 4980
rect 5362 4931 5366 4960
rect 5381 4958 5385 5016
rect 5401 4959 5405 4996
rect 5513 4976 5517 4996
rect 5503 4969 5517 4976
rect 5523 4976 5527 4996
rect 5613 4976 5617 4996
rect 5523 4969 5531 4976
rect 5503 4953 5509 4969
rect 5362 4923 5371 4931
rect 5342 4904 5345 4916
rect 5335 4864 5339 4870
rect 5347 4864 5351 4904
rect 5367 4864 5371 4923
rect 5381 4864 5385 4946
rect 5401 4904 5405 4947
rect 5506 4941 5509 4953
rect 5505 4864 5509 4941
rect 5525 4953 5531 4969
rect 5609 4969 5617 4976
rect 5623 4976 5627 4996
rect 5753 4976 5757 4996
rect 5623 4969 5637 4976
rect 5609 4953 5615 4969
rect 5525 4941 5534 4953
rect 5606 4941 5615 4953
rect 5525 4864 5529 4941
rect 5611 4864 5615 4941
rect 5631 4953 5637 4969
rect 5749 4969 5757 4976
rect 5763 4976 5767 4996
rect 5763 4969 5777 4976
rect 5749 4953 5755 4969
rect 5631 4941 5634 4953
rect 5746 4941 5755 4953
rect 5631 4864 5635 4941
rect 5751 4864 5755 4941
rect 5771 4953 5777 4969
rect 5771 4941 5774 4953
rect 5771 4864 5775 4941
rect 90 4820 94 4824
rect 112 4820 116 4824
rect 120 4820 124 4824
rect 225 4820 229 4824
rect 245 4820 249 4824
rect 265 4820 269 4824
rect 351 4820 355 4824
rect 371 4820 375 4824
rect 391 4820 395 4824
rect 496 4820 500 4824
rect 504 4820 508 4824
rect 526 4820 530 4824
rect 645 4820 649 4824
rect 665 4820 669 4824
rect 770 4820 774 4824
rect 792 4820 796 4824
rect 800 4820 804 4824
rect 910 4820 914 4824
rect 932 4820 936 4824
rect 940 4820 944 4824
rect 1045 4820 1049 4824
rect 1065 4820 1069 4824
rect 1085 4820 1089 4824
rect 1190 4820 1194 4824
rect 1212 4820 1216 4824
rect 1220 4820 1224 4824
rect 1325 4820 1329 4824
rect 1425 4820 1429 4824
rect 1445 4820 1449 4824
rect 1565 4820 1569 4824
rect 1585 4820 1589 4824
rect 1605 4820 1609 4824
rect 1710 4820 1714 4824
rect 1732 4820 1736 4824
rect 1740 4820 1744 4824
rect 1831 4820 1835 4824
rect 1851 4820 1855 4824
rect 1871 4820 1875 4824
rect 1971 4820 1975 4824
rect 1991 4820 1995 4824
rect 2105 4820 2109 4824
rect 2125 4820 2129 4824
rect 2145 4820 2149 4824
rect 2265 4820 2269 4824
rect 2370 4820 2374 4824
rect 2392 4820 2396 4824
rect 2400 4820 2404 4824
rect 2505 4820 2509 4824
rect 2525 4820 2529 4824
rect 2545 4820 2549 4824
rect 2645 4820 2649 4824
rect 2765 4820 2769 4824
rect 2785 4820 2789 4824
rect 2871 4820 2875 4824
rect 2971 4820 2975 4824
rect 2991 4820 2995 4824
rect 3011 4820 3015 4824
rect 3130 4820 3134 4824
rect 3152 4820 3156 4824
rect 3160 4820 3164 4824
rect 3270 4820 3274 4824
rect 3292 4820 3296 4824
rect 3300 4820 3304 4824
rect 3405 4820 3409 4824
rect 3425 4820 3429 4824
rect 3445 4820 3449 4824
rect 3531 4820 3535 4824
rect 3541 4820 3545 4824
rect 3561 4820 3565 4824
rect 3697 4820 3701 4824
rect 3705 4820 3709 4824
rect 3805 4820 3809 4824
rect 3825 4820 3829 4824
rect 3845 4820 3849 4824
rect 3945 4820 3949 4824
rect 4031 4820 4035 4824
rect 4051 4820 4055 4824
rect 4071 4820 4075 4824
rect 4171 4820 4175 4824
rect 4191 4820 4195 4824
rect 4211 4820 4215 4824
rect 4321 4820 4325 4824
rect 4343 4820 4347 4824
rect 4365 4820 4369 4824
rect 4471 4820 4475 4824
rect 4481 4820 4485 4824
rect 4501 4820 4505 4824
rect 4611 4820 4615 4824
rect 4619 4820 4623 4824
rect 4750 4820 4754 4824
rect 4772 4820 4776 4824
rect 4780 4820 4784 4824
rect 4831 4820 4835 4824
rect 4853 4820 4857 4824
rect 4861 4820 4865 4824
rect 4881 4820 4885 4824
rect 4889 4820 4893 4824
rect 4935 4820 4939 4824
rect 4955 4820 4959 4824
rect 4967 4820 4971 4824
rect 4987 4820 4991 4824
rect 5001 4820 5005 4824
rect 5021 4820 5025 4824
rect 5116 4820 5120 4824
rect 5124 4820 5128 4824
rect 5146 4820 5150 4824
rect 5211 4820 5215 4824
rect 5233 4820 5237 4824
rect 5241 4820 5245 4824
rect 5261 4820 5265 4824
rect 5269 4820 5273 4824
rect 5315 4820 5319 4824
rect 5335 4820 5339 4824
rect 5347 4820 5351 4824
rect 5367 4820 5371 4824
rect 5381 4820 5385 4824
rect 5401 4820 5405 4824
rect 5505 4820 5509 4824
rect 5525 4820 5529 4824
rect 5611 4820 5615 4824
rect 5631 4820 5635 4824
rect 5751 4820 5755 4824
rect 5771 4820 5775 4824
rect 85 4796 89 4800
rect 105 4796 109 4800
rect 125 4796 129 4800
rect 225 4796 229 4800
rect 245 4796 249 4800
rect 265 4796 269 4800
rect 351 4796 355 4800
rect 371 4796 375 4800
rect 391 4796 395 4800
rect 491 4796 495 4800
rect 511 4796 515 4800
rect 625 4796 629 4800
rect 645 4796 649 4800
rect 665 4796 669 4800
rect 785 4796 789 4800
rect 805 4796 809 4800
rect 825 4796 829 4800
rect 911 4796 915 4800
rect 1011 4796 1015 4800
rect 1125 4796 1129 4800
rect 1230 4796 1234 4800
rect 1252 4796 1256 4800
rect 1260 4796 1264 4800
rect 1356 4796 1360 4800
rect 1364 4796 1368 4800
rect 1386 4796 1390 4800
rect 1491 4796 1495 4800
rect 1591 4796 1595 4800
rect 1611 4796 1615 4800
rect 1631 4796 1635 4800
rect 1750 4796 1754 4800
rect 1772 4796 1776 4800
rect 1780 4796 1784 4800
rect 1885 4796 1889 4800
rect 1905 4796 1909 4800
rect 1996 4796 2000 4800
rect 2004 4796 2008 4800
rect 2026 4796 2030 4800
rect 2145 4796 2149 4800
rect 2165 4796 2169 4800
rect 2185 4796 2189 4800
rect 2283 4796 2287 4800
rect 2305 4796 2309 4800
rect 2391 4796 2395 4800
rect 2411 4796 2415 4800
rect 2511 4796 2515 4800
rect 2531 4796 2535 4800
rect 2643 4796 2647 4800
rect 2665 4796 2669 4800
rect 2751 4796 2755 4800
rect 2771 4796 2775 4800
rect 2791 4796 2795 4800
rect 2917 4796 2921 4800
rect 2925 4796 2929 4800
rect 3031 4796 3035 4800
rect 3041 4796 3045 4800
rect 3071 4796 3075 4800
rect 3081 4796 3085 4800
rect 3205 4796 3209 4800
rect 3225 4796 3229 4800
rect 3325 4796 3329 4800
rect 3345 4796 3349 4800
rect 3365 4796 3369 4800
rect 3465 4796 3469 4800
rect 3485 4796 3489 4800
rect 3505 4796 3509 4800
rect 3605 4796 3609 4800
rect 3625 4796 3629 4800
rect 3645 4796 3649 4800
rect 3745 4796 3749 4800
rect 3765 4796 3769 4800
rect 3785 4796 3789 4800
rect 3871 4796 3875 4800
rect 3891 4796 3895 4800
rect 3911 4796 3915 4800
rect 4011 4796 4015 4800
rect 4031 4796 4035 4800
rect 4051 4796 4055 4800
rect 4151 4796 4155 4800
rect 4261 4796 4265 4800
rect 4283 4796 4287 4800
rect 4305 4796 4309 4800
rect 4425 4796 4429 4800
rect 4445 4796 4449 4800
rect 4465 4796 4469 4800
rect 4551 4796 4555 4800
rect 4571 4796 4575 4800
rect 4591 4796 4595 4800
rect 4691 4796 4695 4800
rect 4751 4796 4755 4800
rect 4773 4796 4777 4800
rect 4781 4796 4785 4800
rect 4801 4796 4805 4800
rect 4809 4796 4813 4800
rect 4855 4796 4859 4800
rect 4875 4796 4879 4800
rect 4887 4796 4891 4800
rect 4907 4796 4911 4800
rect 4921 4796 4925 4800
rect 4941 4796 4945 4800
rect 5036 4796 5040 4800
rect 5044 4796 5048 4800
rect 5066 4796 5070 4800
rect 5171 4796 5175 4800
rect 5191 4796 5195 4800
rect 5291 4796 5295 4800
rect 5311 4796 5315 4800
rect 5431 4796 5435 4800
rect 5451 4796 5455 4800
rect 5551 4796 5555 4800
rect 5571 4796 5575 4800
rect 5685 4796 5689 4800
rect 5705 4796 5709 4800
rect 5725 4796 5729 4800
rect 85 4659 89 4716
rect 105 4702 109 4716
rect 125 4702 129 4716
rect 225 4713 229 4756
rect 245 4744 249 4756
rect 265 4748 269 4756
rect 265 4744 280 4748
rect 245 4740 260 4744
rect 254 4733 260 4740
rect 105 4696 120 4702
rect 125 4696 141 4702
rect 225 4701 233 4713
rect 245 4701 252 4713
rect 114 4673 120 4696
rect 85 4647 94 4659
rect 92 4604 96 4647
rect 114 4624 118 4661
rect 134 4659 141 4696
rect 134 4634 141 4647
rect 248 4644 252 4701
rect 256 4644 260 4721
rect 274 4713 280 4744
rect 264 4701 274 4713
rect 351 4702 355 4716
rect 371 4702 375 4716
rect 264 4644 268 4701
rect 339 4696 355 4702
rect 360 4696 375 4702
rect 339 4659 346 4696
rect 360 4673 366 4696
rect 122 4628 141 4634
rect 122 4624 126 4628
rect 339 4634 346 4647
rect 339 4628 358 4634
rect 354 4624 358 4628
rect 362 4624 366 4661
rect 391 4659 395 4716
rect 491 4679 495 4756
rect 486 4667 495 4679
rect 386 4647 395 4659
rect 489 4651 495 4667
rect 511 4679 515 4756
rect 625 4713 629 4756
rect 645 4744 649 4756
rect 665 4748 669 4756
rect 665 4744 680 4748
rect 645 4740 660 4744
rect 654 4733 660 4740
rect 625 4701 633 4713
rect 645 4701 652 4713
rect 511 4667 514 4679
rect 511 4651 517 4667
rect 384 4604 388 4647
rect 489 4644 497 4651
rect 493 4624 497 4644
rect 503 4644 517 4651
rect 648 4644 652 4701
rect 656 4644 660 4721
rect 674 4713 680 4744
rect 785 4713 789 4756
rect 805 4744 809 4756
rect 825 4748 829 4756
rect 825 4744 840 4748
rect 805 4740 820 4744
rect 814 4733 820 4740
rect 664 4701 674 4713
rect 785 4701 793 4713
rect 805 4701 812 4713
rect 664 4644 668 4701
rect 808 4644 812 4701
rect 816 4644 820 4721
rect 834 4713 840 4744
rect 824 4701 834 4713
rect 824 4644 828 4701
rect 911 4673 915 4756
rect 1011 4673 1015 4756
rect 906 4661 915 4673
rect 1006 4661 1015 4673
rect 503 4624 507 4644
rect 911 4604 915 4661
rect 1011 4604 1015 4661
rect 1125 4673 1129 4756
rect 1230 4713 1234 4756
rect 1227 4701 1234 4713
rect 1125 4661 1134 4673
rect 1125 4604 1129 4661
rect 1225 4624 1229 4701
rect 1252 4659 1256 4716
rect 1260 4712 1264 4716
rect 1356 4712 1360 4716
rect 1260 4704 1278 4712
rect 1274 4693 1278 4704
rect 1342 4704 1360 4712
rect 1342 4693 1346 4704
rect 1245 4647 1254 4659
rect 1245 4624 1249 4647
rect 1274 4636 1278 4681
rect 1265 4629 1278 4636
rect 1342 4636 1346 4681
rect 1364 4659 1368 4716
rect 1386 4713 1390 4756
rect 1386 4701 1393 4713
rect 1366 4647 1375 4659
rect 1342 4629 1355 4636
rect 1265 4624 1269 4629
rect 1351 4624 1355 4629
rect 1371 4624 1375 4647
rect 1391 4624 1395 4701
rect 1491 4673 1495 4756
rect 1591 4748 1595 4756
rect 1580 4744 1595 4748
rect 1611 4744 1615 4756
rect 1580 4713 1586 4744
rect 1600 4740 1615 4744
rect 1600 4733 1606 4740
rect 1586 4701 1596 4713
rect 1486 4661 1495 4673
rect 1491 4604 1495 4661
rect 1592 4644 1596 4701
rect 1600 4644 1604 4721
rect 1631 4713 1635 4756
rect 1750 4713 1754 4756
rect 1608 4701 1615 4713
rect 1627 4701 1635 4713
rect 1747 4701 1754 4713
rect 1608 4644 1612 4701
rect 1745 4624 1749 4701
rect 1772 4659 1776 4716
rect 1780 4712 1784 4716
rect 1780 4704 1798 4712
rect 1794 4693 1798 4704
rect 1765 4647 1774 4659
rect 1765 4624 1769 4647
rect 1794 4636 1798 4681
rect 1885 4679 1889 4756
rect 1886 4667 1889 4679
rect 1883 4651 1889 4667
rect 1905 4679 1909 4756
rect 1996 4712 2000 4716
rect 1982 4704 2000 4712
rect 1982 4693 1986 4704
rect 1905 4667 1914 4679
rect 1905 4651 1911 4667
rect 1883 4644 1897 4651
rect 1785 4629 1798 4636
rect 1785 4624 1789 4629
rect 1893 4624 1897 4644
rect 1903 4644 1911 4651
rect 1903 4624 1907 4644
rect 1982 4636 1986 4681
rect 2004 4659 2008 4716
rect 2026 4713 2030 4756
rect 2145 4713 2149 4756
rect 2165 4744 2169 4756
rect 2185 4748 2189 4756
rect 2185 4744 2200 4748
rect 2165 4740 2180 4744
rect 2174 4733 2180 4740
rect 2026 4701 2033 4713
rect 2145 4701 2153 4713
rect 2165 4701 2172 4713
rect 2006 4647 2015 4659
rect 1982 4629 1995 4636
rect 1991 4624 1995 4629
rect 2011 4624 2015 4647
rect 2031 4624 2035 4701
rect 2168 4644 2172 4701
rect 2176 4644 2180 4721
rect 2194 4713 2200 4744
rect 2184 4701 2194 4713
rect 2283 4710 2287 4716
rect 2184 4644 2188 4701
rect 2283 4698 2285 4710
rect 2305 4693 2309 4756
rect 2305 4681 2314 4693
rect 2283 4630 2285 4642
rect 2283 4624 2287 4630
rect 2305 4604 2309 4681
rect 2391 4679 2395 4756
rect 2386 4667 2395 4679
rect 2389 4651 2395 4667
rect 2411 4679 2415 4756
rect 2511 4679 2515 4756
rect 2411 4667 2414 4679
rect 2506 4667 2515 4679
rect 2411 4651 2417 4667
rect 2389 4644 2397 4651
rect 2393 4624 2397 4644
rect 2403 4644 2417 4651
rect 2509 4651 2515 4667
rect 2531 4679 2535 4756
rect 2643 4710 2647 4716
rect 2643 4698 2645 4710
rect 2665 4693 2669 4756
rect 2751 4748 2755 4756
rect 2740 4744 2755 4748
rect 2771 4744 2775 4756
rect 2740 4713 2746 4744
rect 2760 4740 2775 4744
rect 2760 4733 2766 4740
rect 2746 4701 2756 4713
rect 2665 4681 2674 4693
rect 2531 4667 2534 4679
rect 2531 4651 2537 4667
rect 2509 4644 2517 4651
rect 2403 4624 2407 4644
rect 2513 4624 2517 4644
rect 2523 4644 2537 4651
rect 2523 4624 2527 4644
rect 2643 4630 2645 4642
rect 2643 4624 2647 4630
rect 2665 4604 2669 4681
rect 2752 4644 2756 4701
rect 2760 4644 2764 4721
rect 2791 4713 2795 4756
rect 2768 4701 2775 4713
rect 2787 4701 2795 4713
rect 2768 4644 2772 4701
rect 2917 4693 2921 4716
rect 2906 4681 2921 4693
rect 2925 4693 2929 4716
rect 3031 4712 3035 4716
rect 3021 4708 3035 4712
rect 3041 4712 3045 4716
rect 3041 4708 3055 4712
rect 3021 4693 3026 4708
rect 2925 4681 2934 4693
rect 2905 4604 2909 4681
rect 2925 4604 2929 4681
rect 3020 4635 3026 4681
rect 3049 4659 3055 4708
rect 3071 4659 3075 4716
rect 3081 4712 3085 4716
rect 3081 4708 3095 4712
rect 3091 4693 3095 4708
rect 3091 4681 3093 4693
rect 3046 4647 3055 4659
rect 3020 4631 3035 4635
rect 3031 4624 3035 4631
rect 3051 4624 3055 4647
rect 3071 4624 3075 4647
rect 3091 4624 3095 4681
rect 3205 4679 3209 4756
rect 3206 4667 3209 4679
rect 3203 4651 3209 4667
rect 3225 4679 3229 4756
rect 3325 4713 3329 4756
rect 3345 4744 3349 4756
rect 3365 4748 3369 4756
rect 3365 4744 3380 4748
rect 3345 4740 3360 4744
rect 3354 4733 3360 4740
rect 3325 4701 3333 4713
rect 3345 4701 3352 4713
rect 3225 4667 3234 4679
rect 3225 4651 3231 4667
rect 3203 4644 3217 4651
rect 3213 4624 3217 4644
rect 3223 4644 3231 4651
rect 3348 4644 3352 4701
rect 3356 4644 3360 4721
rect 3374 4713 3380 4744
rect 3364 4701 3374 4713
rect 3364 4644 3368 4701
rect 3465 4659 3469 4716
rect 3485 4702 3489 4716
rect 3505 4702 3509 4716
rect 3605 4713 3609 4756
rect 3625 4744 3629 4756
rect 3645 4748 3649 4756
rect 3645 4744 3660 4748
rect 3625 4740 3640 4744
rect 3634 4733 3640 4740
rect 3485 4696 3500 4702
rect 3505 4696 3521 4702
rect 3605 4701 3613 4713
rect 3625 4701 3632 4713
rect 3494 4673 3500 4696
rect 3465 4647 3474 4659
rect 3223 4624 3227 4644
rect 3472 4604 3476 4647
rect 3494 4624 3498 4661
rect 3514 4659 3521 4696
rect 3514 4634 3521 4647
rect 3628 4644 3632 4701
rect 3636 4644 3640 4721
rect 3654 4713 3660 4744
rect 3871 4748 3875 4756
rect 3860 4744 3875 4748
rect 3891 4744 3895 4756
rect 3644 4701 3654 4713
rect 3644 4644 3648 4701
rect 3745 4659 3749 4716
rect 3765 4702 3769 4716
rect 3785 4702 3789 4716
rect 3860 4713 3866 4744
rect 3880 4740 3895 4744
rect 3880 4733 3886 4740
rect 3765 4696 3780 4702
rect 3785 4696 3801 4702
rect 3866 4701 3876 4713
rect 3774 4673 3780 4696
rect 3745 4647 3754 4659
rect 3502 4628 3521 4634
rect 3502 4624 3506 4628
rect 3752 4604 3756 4647
rect 3774 4624 3778 4661
rect 3794 4659 3801 4696
rect 3794 4634 3801 4647
rect 3872 4644 3876 4701
rect 3880 4644 3884 4721
rect 3911 4713 3915 4756
rect 4011 4748 4015 4756
rect 4000 4744 4015 4748
rect 4031 4744 4035 4756
rect 4000 4713 4006 4744
rect 4020 4740 4035 4744
rect 4020 4733 4026 4740
rect 3888 4701 3895 4713
rect 3907 4701 3915 4713
rect 4006 4701 4016 4713
rect 3888 4644 3892 4701
rect 4012 4644 4016 4701
rect 4020 4644 4024 4721
rect 4051 4713 4055 4756
rect 4028 4701 4035 4713
rect 4047 4701 4055 4713
rect 4028 4644 4032 4701
rect 4151 4673 4155 4756
rect 4146 4661 4155 4673
rect 3782 4628 3801 4634
rect 3782 4624 3786 4628
rect 4151 4604 4155 4661
rect 4261 4642 4265 4716
rect 4283 4679 4287 4756
rect 4305 4693 4309 4756
rect 4425 4713 4429 4756
rect 4445 4744 4449 4756
rect 4465 4748 4469 4756
rect 4551 4748 4555 4756
rect 4465 4744 4480 4748
rect 4445 4740 4460 4744
rect 4454 4733 4460 4740
rect 4425 4701 4433 4713
rect 4445 4701 4452 4713
rect 4305 4681 4314 4693
rect 4286 4667 4299 4679
rect 4261 4630 4273 4642
rect 4275 4624 4279 4630
rect 4295 4624 4299 4667
rect 4305 4624 4309 4681
rect 4448 4644 4452 4701
rect 4456 4644 4460 4721
rect 4474 4713 4480 4744
rect 4540 4744 4555 4748
rect 4571 4744 4575 4756
rect 4540 4713 4546 4744
rect 4560 4740 4575 4744
rect 4560 4733 4566 4740
rect 4464 4701 4474 4713
rect 4546 4701 4556 4713
rect 4464 4644 4468 4701
rect 4552 4644 4556 4701
rect 4560 4644 4564 4721
rect 4591 4713 4595 4756
rect 4568 4701 4575 4713
rect 4587 4701 4595 4713
rect 4568 4644 4572 4701
rect 4691 4673 4695 4756
rect 4773 4753 4777 4776
rect 4769 4746 4777 4753
rect 4769 4717 4773 4746
rect 4781 4736 4785 4776
rect 4801 4724 4805 4756
rect 4809 4752 4813 4756
rect 4809 4750 4845 4752
rect 4809 4748 4833 4750
rect 4686 4661 4695 4673
rect 4691 4604 4695 4661
rect 4751 4704 4755 4716
rect 4769 4711 4777 4717
rect 4751 4692 4753 4704
rect 4751 4624 4755 4692
rect 4773 4665 4777 4711
rect 4773 4604 4777 4653
rect 4801 4629 4807 4724
rect 4783 4625 4807 4629
rect 4783 4604 4787 4625
rect 4803 4620 4821 4621
rect 4803 4616 4833 4620
rect 4803 4604 4807 4616
rect 4841 4612 4845 4738
rect 4855 4730 4859 4756
rect 4875 4750 4879 4756
rect 4811 4608 4845 4612
rect 4811 4604 4815 4608
rect 4857 4604 4861 4718
rect 4873 4628 4877 4738
rect 4887 4716 4891 4756
rect 4882 4704 4885 4716
rect 4882 4640 4886 4704
rect 4907 4697 4911 4756
rect 4902 4689 4911 4697
rect 4902 4660 4906 4689
rect 4921 4674 4925 4756
rect 4941 4673 4945 4716
rect 5036 4712 5040 4716
rect 5022 4704 5040 4712
rect 5022 4693 5026 4704
rect 4882 4636 4915 4640
rect 4881 4616 4883 4628
rect 4879 4604 4883 4616
rect 4889 4616 4891 4628
rect 4889 4604 4893 4616
rect 4911 4604 4915 4636
rect 4921 4604 4925 4662
rect 4941 4624 4945 4661
rect 5022 4636 5026 4681
rect 5044 4659 5048 4716
rect 5066 4713 5070 4756
rect 5066 4701 5073 4713
rect 5046 4647 5055 4659
rect 5022 4629 5035 4636
rect 5031 4624 5035 4629
rect 5051 4624 5055 4647
rect 5071 4624 5075 4701
rect 5171 4679 5175 4756
rect 5166 4667 5175 4679
rect 5169 4651 5175 4667
rect 5191 4679 5195 4756
rect 5291 4679 5295 4756
rect 5191 4667 5194 4679
rect 5286 4667 5295 4679
rect 5191 4651 5197 4667
rect 5169 4644 5177 4651
rect 5173 4624 5177 4644
rect 5183 4644 5197 4651
rect 5289 4651 5295 4667
rect 5311 4679 5315 4756
rect 5431 4679 5435 4756
rect 5311 4667 5314 4679
rect 5426 4667 5435 4679
rect 5311 4651 5317 4667
rect 5289 4644 5297 4651
rect 5183 4624 5187 4644
rect 5293 4624 5297 4644
rect 5303 4644 5317 4651
rect 5429 4651 5435 4667
rect 5451 4679 5455 4756
rect 5551 4679 5555 4756
rect 5451 4667 5454 4679
rect 5546 4667 5555 4679
rect 5451 4651 5457 4667
rect 5429 4644 5437 4651
rect 5303 4624 5307 4644
rect 5433 4624 5437 4644
rect 5443 4644 5457 4651
rect 5549 4651 5555 4667
rect 5571 4679 5575 4756
rect 5685 4713 5689 4756
rect 5705 4744 5709 4756
rect 5725 4748 5729 4756
rect 5725 4744 5740 4748
rect 5705 4740 5720 4744
rect 5714 4733 5720 4740
rect 5685 4701 5693 4713
rect 5705 4701 5712 4713
rect 5571 4667 5574 4679
rect 5571 4651 5577 4667
rect 5549 4644 5557 4651
rect 5443 4624 5447 4644
rect 5553 4624 5557 4644
rect 5563 4644 5577 4651
rect 5708 4644 5712 4701
rect 5716 4644 5720 4721
rect 5734 4713 5740 4744
rect 5724 4701 5734 4713
rect 5724 4644 5728 4701
rect 5563 4624 5567 4644
rect 92 4580 96 4584
rect 114 4580 118 4584
rect 122 4580 126 4584
rect 248 4580 252 4584
rect 256 4580 260 4584
rect 264 4580 268 4584
rect 354 4580 358 4584
rect 362 4580 366 4584
rect 384 4580 388 4584
rect 493 4580 497 4584
rect 503 4580 507 4584
rect 648 4580 652 4584
rect 656 4580 660 4584
rect 664 4580 668 4584
rect 808 4580 812 4584
rect 816 4580 820 4584
rect 824 4580 828 4584
rect 911 4580 915 4584
rect 1011 4580 1015 4584
rect 1125 4580 1129 4584
rect 1225 4580 1229 4584
rect 1245 4580 1249 4584
rect 1265 4580 1269 4584
rect 1351 4580 1355 4584
rect 1371 4580 1375 4584
rect 1391 4580 1395 4584
rect 1491 4580 1495 4584
rect 1592 4580 1596 4584
rect 1600 4580 1604 4584
rect 1608 4580 1612 4584
rect 1745 4580 1749 4584
rect 1765 4580 1769 4584
rect 1785 4580 1789 4584
rect 1893 4580 1897 4584
rect 1903 4580 1907 4584
rect 1991 4580 1995 4584
rect 2011 4580 2015 4584
rect 2031 4580 2035 4584
rect 2168 4580 2172 4584
rect 2176 4580 2180 4584
rect 2184 4580 2188 4584
rect 2283 4580 2287 4584
rect 2305 4580 2309 4584
rect 2393 4580 2397 4584
rect 2403 4580 2407 4584
rect 2513 4580 2517 4584
rect 2523 4580 2527 4584
rect 2643 4580 2647 4584
rect 2665 4580 2669 4584
rect 2752 4580 2756 4584
rect 2760 4580 2764 4584
rect 2768 4580 2772 4584
rect 2905 4580 2909 4584
rect 2925 4580 2929 4584
rect 3031 4580 3035 4584
rect 3051 4580 3055 4584
rect 3071 4580 3075 4584
rect 3091 4580 3095 4584
rect 3213 4580 3217 4584
rect 3223 4580 3227 4584
rect 3348 4580 3352 4584
rect 3356 4580 3360 4584
rect 3364 4580 3368 4584
rect 3472 4580 3476 4584
rect 3494 4580 3498 4584
rect 3502 4580 3506 4584
rect 3628 4580 3632 4584
rect 3636 4580 3640 4584
rect 3644 4580 3648 4584
rect 3752 4580 3756 4584
rect 3774 4580 3778 4584
rect 3782 4580 3786 4584
rect 3872 4580 3876 4584
rect 3880 4580 3884 4584
rect 3888 4580 3892 4584
rect 4012 4580 4016 4584
rect 4020 4580 4024 4584
rect 4028 4580 4032 4584
rect 4151 4580 4155 4584
rect 4275 4580 4279 4584
rect 4295 4580 4299 4584
rect 4305 4580 4309 4584
rect 4448 4580 4452 4584
rect 4456 4580 4460 4584
rect 4464 4580 4468 4584
rect 4552 4580 4556 4584
rect 4560 4580 4564 4584
rect 4568 4580 4572 4584
rect 4691 4580 4695 4584
rect 4751 4580 4755 4584
rect 4773 4580 4777 4584
rect 4783 4580 4787 4584
rect 4803 4580 4807 4584
rect 4811 4580 4815 4584
rect 4857 4580 4861 4584
rect 4879 4580 4883 4584
rect 4889 4580 4893 4584
rect 4911 4580 4915 4584
rect 4921 4580 4925 4584
rect 4941 4580 4945 4584
rect 5031 4580 5035 4584
rect 5051 4580 5055 4584
rect 5071 4580 5075 4584
rect 5173 4580 5177 4584
rect 5183 4580 5187 4584
rect 5293 4580 5297 4584
rect 5303 4580 5307 4584
rect 5433 4580 5437 4584
rect 5443 4580 5447 4584
rect 5553 4580 5557 4584
rect 5563 4580 5567 4584
rect 5708 4580 5712 4584
rect 5716 4580 5720 4584
rect 5724 4580 5728 4584
rect 85 4556 89 4560
rect 105 4556 109 4560
rect 125 4556 129 4560
rect 248 4556 252 4560
rect 256 4556 260 4560
rect 264 4556 268 4560
rect 354 4556 358 4560
rect 362 4556 366 4560
rect 384 4556 388 4560
rect 525 4556 529 4560
rect 545 4556 549 4560
rect 565 4556 569 4560
rect 665 4556 669 4560
rect 685 4556 689 4560
rect 705 4556 709 4560
rect 791 4556 795 4560
rect 894 4556 898 4560
rect 902 4556 906 4560
rect 924 4556 928 4560
rect 1045 4556 1049 4560
rect 1168 4556 1172 4560
rect 1176 4556 1180 4560
rect 1184 4556 1188 4560
rect 1292 4556 1296 4560
rect 1314 4556 1318 4560
rect 1322 4556 1326 4560
rect 1425 4556 1429 4560
rect 1511 4556 1515 4560
rect 1531 4556 1535 4560
rect 1551 4556 1555 4560
rect 1673 4556 1677 4560
rect 1683 4556 1687 4560
rect 1808 4556 1812 4560
rect 1816 4556 1820 4560
rect 1824 4556 1828 4560
rect 1925 4556 1929 4560
rect 1945 4556 1949 4560
rect 2068 4556 2072 4560
rect 2076 4556 2080 4560
rect 2084 4556 2088 4560
rect 2228 4556 2232 4560
rect 2236 4556 2240 4560
rect 2244 4556 2248 4560
rect 2353 4556 2357 4560
rect 2363 4556 2367 4560
rect 2488 4556 2492 4560
rect 2496 4556 2500 4560
rect 2504 4556 2508 4560
rect 2592 4556 2596 4560
rect 2600 4556 2604 4560
rect 2608 4556 2612 4560
rect 2745 4556 2749 4560
rect 2845 4556 2849 4560
rect 2865 4556 2869 4560
rect 2988 4556 2992 4560
rect 2996 4556 3000 4560
rect 3004 4556 3008 4560
rect 3128 4556 3132 4560
rect 3136 4556 3140 4560
rect 3144 4556 3148 4560
rect 3231 4556 3235 4560
rect 3331 4556 3335 4560
rect 3351 4556 3355 4560
rect 3371 4556 3375 4560
rect 3495 4556 3499 4560
rect 3515 4556 3519 4560
rect 3525 4556 3529 4560
rect 3633 4556 3637 4560
rect 3643 4556 3647 4560
rect 3765 4556 3769 4560
rect 3785 4556 3789 4560
rect 3805 4556 3809 4560
rect 3893 4556 3897 4560
rect 3903 4556 3907 4560
rect 4023 4556 4027 4560
rect 4045 4556 4049 4560
rect 4131 4556 4135 4560
rect 4141 4556 4145 4560
rect 4161 4556 4165 4560
rect 4293 4556 4297 4560
rect 4303 4556 4307 4560
rect 4405 4556 4409 4560
rect 4425 4556 4429 4560
rect 4445 4556 4449 4560
rect 4533 4556 4537 4560
rect 4543 4556 4547 4560
rect 4673 4556 4677 4560
rect 4683 4556 4687 4560
rect 4771 4556 4775 4560
rect 4873 4556 4877 4560
rect 4883 4556 4887 4560
rect 4991 4556 4995 4560
rect 5011 4556 5015 4560
rect 5031 4556 5035 4560
rect 5091 4556 5095 4560
rect 5113 4556 5117 4560
rect 5123 4556 5127 4560
rect 5143 4556 5147 4560
rect 5151 4556 5155 4560
rect 5197 4556 5201 4560
rect 5219 4556 5223 4560
rect 5229 4556 5233 4560
rect 5251 4556 5255 4560
rect 5261 4556 5265 4560
rect 5281 4556 5285 4560
rect 5371 4556 5375 4560
rect 5391 4556 5395 4560
rect 5411 4556 5415 4560
rect 5511 4556 5515 4560
rect 5531 4556 5535 4560
rect 5551 4556 5555 4560
rect 5665 4556 5669 4560
rect 5685 4556 5689 4560
rect 5705 4556 5709 4560
rect 85 4439 89 4516
rect 105 4493 109 4516
rect 125 4511 129 4516
rect 125 4504 138 4511
rect 105 4481 114 4493
rect 87 4427 94 4439
rect 90 4384 94 4427
rect 112 4424 116 4481
rect 134 4459 138 4504
rect 354 4512 358 4516
rect 339 4506 358 4512
rect 134 4436 138 4447
rect 248 4439 252 4496
rect 120 4428 138 4436
rect 120 4424 124 4428
rect 225 4427 233 4439
rect 245 4427 252 4439
rect 225 4384 229 4427
rect 256 4419 260 4496
rect 264 4439 268 4496
rect 339 4493 346 4506
rect 339 4444 346 4481
rect 362 4479 366 4516
rect 384 4493 388 4536
rect 386 4481 395 4493
rect 360 4444 366 4467
rect 264 4427 274 4439
rect 339 4438 355 4444
rect 360 4438 375 4444
rect 254 4400 260 4407
rect 245 4396 260 4400
rect 274 4396 280 4427
rect 351 4424 355 4438
rect 371 4424 375 4438
rect 391 4424 395 4481
rect 525 4439 529 4516
rect 545 4493 549 4516
rect 565 4511 569 4516
rect 565 4504 578 4511
rect 545 4481 554 4493
rect 527 4427 534 4439
rect 245 4384 249 4396
rect 265 4392 280 4396
rect 265 4384 269 4392
rect 530 4384 534 4427
rect 552 4424 556 4481
rect 574 4459 578 4504
rect 574 4436 578 4447
rect 665 4439 669 4516
rect 685 4493 689 4516
rect 705 4511 709 4516
rect 705 4504 718 4511
rect 685 4481 694 4493
rect 560 4428 578 4436
rect 560 4424 564 4428
rect 667 4427 674 4439
rect 670 4384 674 4427
rect 692 4424 696 4481
rect 714 4459 718 4504
rect 791 4479 795 4536
rect 894 4512 898 4516
rect 879 4506 898 4512
rect 879 4493 886 4506
rect 786 4467 795 4479
rect 714 4436 718 4447
rect 700 4428 718 4436
rect 700 4424 704 4428
rect 791 4384 795 4467
rect 879 4444 886 4481
rect 902 4479 906 4516
rect 924 4493 928 4536
rect 926 4481 935 4493
rect 900 4444 906 4467
rect 879 4438 895 4444
rect 900 4438 915 4444
rect 891 4424 895 4438
rect 911 4424 915 4438
rect 931 4424 935 4481
rect 1045 4479 1049 4536
rect 1045 4467 1054 4479
rect 1045 4384 1049 4467
rect 1168 4439 1172 4496
rect 1145 4427 1153 4439
rect 1165 4427 1172 4439
rect 1145 4384 1149 4427
rect 1176 4419 1180 4496
rect 1184 4439 1188 4496
rect 1292 4493 1296 4536
rect 1285 4481 1294 4493
rect 1184 4427 1194 4439
rect 1174 4400 1180 4407
rect 1165 4396 1180 4400
rect 1194 4396 1200 4427
rect 1285 4424 1289 4481
rect 1314 4479 1318 4516
rect 1322 4512 1326 4516
rect 1322 4506 1341 4512
rect 1334 4493 1341 4506
rect 1314 4444 1320 4467
rect 1334 4444 1341 4481
rect 1305 4438 1320 4444
rect 1325 4438 1341 4444
rect 1425 4479 1429 4536
rect 1511 4511 1515 4516
rect 1502 4504 1515 4511
rect 1425 4467 1434 4479
rect 1305 4424 1309 4438
rect 1325 4424 1329 4438
rect 1165 4384 1169 4396
rect 1185 4392 1200 4396
rect 1185 4384 1189 4392
rect 1425 4384 1429 4467
rect 1502 4459 1506 4504
rect 1531 4493 1535 4516
rect 1526 4481 1535 4493
rect 1502 4436 1506 4447
rect 1502 4428 1520 4436
rect 1516 4424 1520 4428
rect 1524 4424 1528 4481
rect 1551 4439 1555 4516
rect 1673 4496 1677 4516
rect 1663 4489 1677 4496
rect 1683 4496 1687 4516
rect 1683 4489 1691 4496
rect 1663 4473 1669 4489
rect 1666 4461 1669 4473
rect 1546 4427 1553 4439
rect 1546 4384 1550 4427
rect 1665 4384 1669 4461
rect 1685 4473 1691 4489
rect 1685 4461 1694 4473
rect 1685 4384 1689 4461
rect 1808 4439 1812 4496
rect 1785 4427 1793 4439
rect 1805 4427 1812 4439
rect 1785 4384 1789 4427
rect 1816 4419 1820 4496
rect 1824 4439 1828 4496
rect 1925 4459 1929 4536
rect 1945 4459 1949 4536
rect 2353 4496 2357 4516
rect 1926 4447 1941 4459
rect 1824 4427 1834 4439
rect 1814 4400 1820 4407
rect 1805 4396 1820 4400
rect 1834 4396 1840 4427
rect 1937 4424 1941 4447
rect 1945 4447 1954 4459
rect 1945 4424 1949 4447
rect 2068 4439 2072 4496
rect 2045 4427 2053 4439
rect 2065 4427 2072 4439
rect 1805 4384 1809 4396
rect 1825 4392 1840 4396
rect 1825 4384 1829 4392
rect 2045 4384 2049 4427
rect 2076 4419 2080 4496
rect 2084 4439 2088 4496
rect 2228 4439 2232 4496
rect 2084 4427 2094 4439
rect 2205 4427 2213 4439
rect 2225 4427 2232 4439
rect 2074 4400 2080 4407
rect 2065 4396 2080 4400
rect 2094 4396 2100 4427
rect 2065 4384 2069 4396
rect 2085 4392 2100 4396
rect 2085 4384 2089 4392
rect 2205 4384 2209 4427
rect 2236 4419 2240 4496
rect 2244 4439 2248 4496
rect 2343 4489 2357 4496
rect 2363 4496 2367 4516
rect 2363 4489 2371 4496
rect 2343 4473 2349 4489
rect 2346 4461 2349 4473
rect 2244 4427 2254 4439
rect 2234 4400 2240 4407
rect 2225 4396 2240 4400
rect 2254 4396 2260 4427
rect 2225 4384 2229 4396
rect 2245 4392 2260 4396
rect 2245 4384 2249 4392
rect 2345 4384 2349 4461
rect 2365 4473 2371 4489
rect 2365 4461 2374 4473
rect 2365 4384 2369 4461
rect 2488 4439 2492 4496
rect 2465 4427 2473 4439
rect 2485 4427 2492 4439
rect 2465 4384 2469 4427
rect 2496 4419 2500 4496
rect 2504 4439 2508 4496
rect 2592 4439 2596 4496
rect 2504 4427 2514 4439
rect 2586 4427 2596 4439
rect 2494 4400 2500 4407
rect 2485 4396 2500 4400
rect 2514 4396 2520 4427
rect 2485 4384 2489 4396
rect 2505 4392 2520 4396
rect 2580 4396 2586 4427
rect 2600 4419 2604 4496
rect 2608 4439 2612 4496
rect 2745 4479 2749 4536
rect 2745 4467 2754 4479
rect 2608 4427 2615 4439
rect 2627 4427 2635 4439
rect 2600 4400 2606 4407
rect 2600 4396 2615 4400
rect 2580 4392 2595 4396
rect 2505 4384 2509 4392
rect 2591 4384 2595 4392
rect 2611 4384 2615 4396
rect 2631 4384 2635 4427
rect 2745 4384 2749 4467
rect 2845 4459 2849 4536
rect 2865 4459 2869 4536
rect 2846 4447 2861 4459
rect 2857 4424 2861 4447
rect 2865 4447 2874 4459
rect 2865 4424 2869 4447
rect 2988 4439 2992 4496
rect 2965 4427 2973 4439
rect 2985 4427 2992 4439
rect 2965 4384 2969 4427
rect 2996 4419 3000 4496
rect 3004 4439 3008 4496
rect 3128 4439 3132 4496
rect 3004 4427 3014 4439
rect 3105 4427 3113 4439
rect 3125 4427 3132 4439
rect 2994 4400 3000 4407
rect 2985 4396 3000 4400
rect 3014 4396 3020 4427
rect 2985 4384 2989 4396
rect 3005 4392 3020 4396
rect 3005 4384 3009 4392
rect 3105 4384 3109 4427
rect 3136 4419 3140 4496
rect 3144 4439 3148 4496
rect 3231 4479 3235 4536
rect 3785 4529 3789 4536
rect 3805 4529 3809 4536
rect 3785 4523 3799 4529
rect 3805 4524 3818 4529
rect 3331 4511 3335 4516
rect 3226 4467 3235 4479
rect 3144 4427 3154 4439
rect 3134 4400 3140 4407
rect 3125 4396 3140 4400
rect 3154 4396 3160 4427
rect 3125 4384 3129 4396
rect 3145 4392 3160 4396
rect 3145 4384 3149 4392
rect 3231 4384 3235 4467
rect 3322 4504 3335 4511
rect 3322 4459 3326 4504
rect 3351 4493 3355 4516
rect 3346 4481 3355 4493
rect 3322 4436 3326 4447
rect 3322 4428 3340 4436
rect 3336 4424 3340 4428
rect 3344 4424 3348 4481
rect 3371 4439 3375 4516
rect 3495 4510 3499 4516
rect 3481 4498 3493 4510
rect 3366 4427 3373 4439
rect 3366 4384 3370 4427
rect 3481 4424 3485 4498
rect 3515 4473 3519 4516
rect 3506 4461 3519 4473
rect 3503 4384 3507 4461
rect 3525 4459 3529 4516
rect 3633 4496 3637 4516
rect 3629 4489 3637 4496
rect 3643 4496 3647 4516
rect 3765 4508 3769 4516
rect 3765 4496 3775 4508
rect 3643 4489 3657 4496
rect 3629 4473 3635 4489
rect 3626 4461 3635 4473
rect 3525 4447 3534 4459
rect 3525 4384 3529 4447
rect 3631 4384 3635 4461
rect 3651 4473 3657 4489
rect 3651 4461 3654 4473
rect 3651 4384 3655 4461
rect 3795 4459 3799 4523
rect 3814 4479 3818 4524
rect 3893 4496 3897 4516
rect 3889 4489 3897 4496
rect 3903 4496 3907 4516
rect 4023 4510 4027 4516
rect 4023 4498 4025 4510
rect 3903 4489 3917 4496
rect 3889 4473 3895 4489
rect 3775 4424 3779 4429
rect 3795 4424 3799 4447
rect 3814 4433 3818 4467
rect 3886 4461 3895 4473
rect 3805 4428 3818 4433
rect 3805 4424 3809 4428
rect 3891 4384 3895 4461
rect 3911 4473 3917 4489
rect 3911 4461 3914 4473
rect 3911 4384 3915 4461
rect 4045 4459 4049 4536
rect 4131 4459 4135 4516
rect 4141 4473 4145 4516
rect 4161 4510 4165 4516
rect 4167 4498 4179 4510
rect 4141 4461 4154 4473
rect 4045 4447 4054 4459
rect 4126 4447 4135 4459
rect 4023 4430 4025 4442
rect 4023 4424 4027 4430
rect 4045 4384 4049 4447
rect 4131 4384 4135 4447
rect 4153 4384 4157 4461
rect 4175 4424 4179 4498
rect 4293 4496 4297 4516
rect 4283 4489 4297 4496
rect 4303 4496 4307 4516
rect 4303 4489 4311 4496
rect 4283 4473 4289 4489
rect 4286 4461 4289 4473
rect 4285 4384 4289 4461
rect 4305 4473 4311 4489
rect 4305 4461 4314 4473
rect 4305 4384 4309 4461
rect 4405 4439 4409 4516
rect 4425 4493 4429 4516
rect 4445 4511 4449 4516
rect 4445 4504 4458 4511
rect 4425 4481 4434 4493
rect 4407 4427 4414 4439
rect 4410 4384 4414 4427
rect 4432 4424 4436 4481
rect 4454 4459 4458 4504
rect 4533 4496 4537 4516
rect 4529 4489 4537 4496
rect 4543 4496 4547 4516
rect 4673 4496 4677 4516
rect 4543 4489 4557 4496
rect 4529 4473 4535 4489
rect 4526 4461 4535 4473
rect 4454 4436 4458 4447
rect 4440 4428 4458 4436
rect 4440 4424 4444 4428
rect 4531 4384 4535 4461
rect 4551 4473 4557 4489
rect 4663 4489 4677 4496
rect 4683 4496 4687 4516
rect 4683 4489 4691 4496
rect 4663 4473 4669 4489
rect 4551 4461 4554 4473
rect 4666 4461 4669 4473
rect 4551 4384 4555 4461
rect 4665 4384 4669 4461
rect 4685 4473 4691 4489
rect 4771 4479 4775 4536
rect 4873 4496 4877 4516
rect 4685 4461 4694 4473
rect 4766 4467 4775 4479
rect 4869 4489 4877 4496
rect 4883 4496 4887 4516
rect 4991 4511 4995 4516
rect 4982 4504 4995 4511
rect 4883 4489 4897 4496
rect 4869 4473 4875 4489
rect 4685 4384 4689 4461
rect 4771 4384 4775 4467
rect 4866 4461 4875 4473
rect 4871 4384 4875 4461
rect 4891 4473 4897 4489
rect 4891 4461 4894 4473
rect 4891 4384 4895 4461
rect 4982 4459 4986 4504
rect 5011 4493 5015 4516
rect 5006 4481 5015 4493
rect 4982 4436 4986 4447
rect 4982 4428 5000 4436
rect 4996 4424 5000 4428
rect 5004 4424 5008 4481
rect 5031 4439 5035 4516
rect 5091 4448 5095 4516
rect 5113 4487 5117 4536
rect 5123 4515 5127 4536
rect 5143 4524 5147 4536
rect 5151 4532 5155 4536
rect 5151 4528 5185 4532
rect 5143 4520 5173 4524
rect 5143 4519 5161 4520
rect 5123 4511 5147 4515
rect 5026 4427 5033 4439
rect 5091 4436 5093 4448
rect 5026 4384 5030 4427
rect 5091 4424 5095 4436
rect 5113 4429 5117 4475
rect 5109 4423 5117 4429
rect 5109 4394 5113 4423
rect 5141 4416 5147 4511
rect 5109 4387 5117 4394
rect 5113 4364 5117 4387
rect 5121 4364 5125 4404
rect 5141 4384 5145 4416
rect 5181 4402 5185 4528
rect 5197 4422 5201 4536
rect 5219 4524 5223 4536
rect 5221 4512 5223 4524
rect 5229 4524 5233 4536
rect 5229 4512 5231 4524
rect 5149 4390 5173 4392
rect 5149 4388 5185 4390
rect 5149 4384 5153 4388
rect 5195 4384 5199 4410
rect 5213 4402 5217 4512
rect 5251 4504 5255 4536
rect 5222 4500 5255 4504
rect 5222 4436 5226 4500
rect 5242 4451 5246 4480
rect 5261 4478 5265 4536
rect 5511 4529 5515 4536
rect 5531 4529 5535 4536
rect 5502 4524 5515 4529
rect 5281 4479 5285 4516
rect 5371 4511 5375 4516
rect 5362 4504 5375 4511
rect 5242 4443 5251 4451
rect 5222 4424 5225 4436
rect 5215 4384 5219 4390
rect 5227 4384 5231 4424
rect 5247 4384 5251 4443
rect 5261 4384 5265 4466
rect 5281 4424 5285 4467
rect 5362 4459 5366 4504
rect 5391 4493 5395 4516
rect 5386 4481 5395 4493
rect 5362 4436 5366 4447
rect 5362 4428 5380 4436
rect 5376 4424 5380 4428
rect 5384 4424 5388 4481
rect 5411 4439 5415 4516
rect 5502 4479 5506 4524
rect 5406 4427 5413 4439
rect 5502 4433 5506 4467
rect 5521 4523 5535 4529
rect 5521 4459 5525 4523
rect 5551 4508 5555 4516
rect 5545 4496 5555 4508
rect 5502 4428 5515 4433
rect 5406 4384 5410 4427
rect 5511 4424 5515 4428
rect 5521 4424 5525 4447
rect 5665 4439 5669 4516
rect 5685 4493 5689 4516
rect 5705 4511 5709 4516
rect 5705 4504 5718 4511
rect 5685 4481 5694 4493
rect 5541 4424 5545 4429
rect 5667 4427 5674 4439
rect 5670 4384 5674 4427
rect 5692 4424 5696 4481
rect 5714 4459 5718 4504
rect 5714 4436 5718 4447
rect 5700 4428 5718 4436
rect 5700 4424 5704 4428
rect 90 4340 94 4344
rect 112 4340 116 4344
rect 120 4340 124 4344
rect 225 4340 229 4344
rect 245 4340 249 4344
rect 265 4340 269 4344
rect 351 4340 355 4344
rect 371 4340 375 4344
rect 391 4340 395 4344
rect 530 4340 534 4344
rect 552 4340 556 4344
rect 560 4340 564 4344
rect 670 4340 674 4344
rect 692 4340 696 4344
rect 700 4340 704 4344
rect 791 4340 795 4344
rect 891 4340 895 4344
rect 911 4340 915 4344
rect 931 4340 935 4344
rect 1045 4340 1049 4344
rect 1145 4340 1149 4344
rect 1165 4340 1169 4344
rect 1185 4340 1189 4344
rect 1285 4340 1289 4344
rect 1305 4340 1309 4344
rect 1325 4340 1329 4344
rect 1425 4340 1429 4344
rect 1516 4340 1520 4344
rect 1524 4340 1528 4344
rect 1546 4340 1550 4344
rect 1665 4340 1669 4344
rect 1685 4340 1689 4344
rect 1785 4340 1789 4344
rect 1805 4340 1809 4344
rect 1825 4340 1829 4344
rect 1937 4340 1941 4344
rect 1945 4340 1949 4344
rect 2045 4340 2049 4344
rect 2065 4340 2069 4344
rect 2085 4340 2089 4344
rect 2205 4340 2209 4344
rect 2225 4340 2229 4344
rect 2245 4340 2249 4344
rect 2345 4340 2349 4344
rect 2365 4340 2369 4344
rect 2465 4340 2469 4344
rect 2485 4340 2489 4344
rect 2505 4340 2509 4344
rect 2591 4340 2595 4344
rect 2611 4340 2615 4344
rect 2631 4340 2635 4344
rect 2745 4340 2749 4344
rect 2857 4340 2861 4344
rect 2865 4340 2869 4344
rect 2965 4340 2969 4344
rect 2985 4340 2989 4344
rect 3005 4340 3009 4344
rect 3105 4340 3109 4344
rect 3125 4340 3129 4344
rect 3145 4340 3149 4344
rect 3231 4340 3235 4344
rect 3336 4340 3340 4344
rect 3344 4340 3348 4344
rect 3366 4340 3370 4344
rect 3481 4340 3485 4344
rect 3503 4340 3507 4344
rect 3525 4340 3529 4344
rect 3631 4340 3635 4344
rect 3651 4340 3655 4344
rect 3775 4340 3779 4344
rect 3795 4340 3799 4344
rect 3805 4340 3809 4344
rect 3891 4340 3895 4344
rect 3911 4340 3915 4344
rect 4023 4340 4027 4344
rect 4045 4340 4049 4344
rect 4131 4340 4135 4344
rect 4153 4340 4157 4344
rect 4175 4340 4179 4344
rect 4285 4340 4289 4344
rect 4305 4340 4309 4344
rect 4410 4340 4414 4344
rect 4432 4340 4436 4344
rect 4440 4340 4444 4344
rect 4531 4340 4535 4344
rect 4551 4340 4555 4344
rect 4665 4340 4669 4344
rect 4685 4340 4689 4344
rect 4771 4340 4775 4344
rect 4871 4340 4875 4344
rect 4891 4340 4895 4344
rect 4996 4340 5000 4344
rect 5004 4340 5008 4344
rect 5026 4340 5030 4344
rect 5091 4340 5095 4344
rect 5113 4340 5117 4344
rect 5121 4340 5125 4344
rect 5141 4340 5145 4344
rect 5149 4340 5153 4344
rect 5195 4340 5199 4344
rect 5215 4340 5219 4344
rect 5227 4340 5231 4344
rect 5247 4340 5251 4344
rect 5261 4340 5265 4344
rect 5281 4340 5285 4344
rect 5376 4340 5380 4344
rect 5384 4340 5388 4344
rect 5406 4340 5410 4344
rect 5511 4340 5515 4344
rect 5521 4340 5525 4344
rect 5541 4340 5545 4344
rect 5670 4340 5674 4344
rect 5692 4340 5696 4344
rect 5700 4340 5704 4344
rect 110 4316 114 4320
rect 132 4316 136 4320
rect 140 4316 144 4320
rect 250 4316 254 4320
rect 272 4316 276 4320
rect 280 4316 284 4320
rect 405 4316 409 4320
rect 425 4316 429 4320
rect 445 4316 449 4320
rect 545 4316 549 4320
rect 565 4316 569 4320
rect 585 4316 589 4320
rect 695 4316 699 4320
rect 715 4316 719 4320
rect 725 4316 729 4320
rect 830 4316 834 4320
rect 852 4316 856 4320
rect 860 4316 864 4320
rect 951 4316 955 4320
rect 1065 4316 1069 4320
rect 1085 4316 1089 4320
rect 1105 4316 1109 4320
rect 1225 4316 1229 4320
rect 1245 4316 1249 4320
rect 1265 4316 1269 4320
rect 1365 4316 1369 4320
rect 1385 4316 1389 4320
rect 1485 4316 1489 4320
rect 1505 4316 1509 4320
rect 1617 4316 1621 4320
rect 1625 4316 1629 4320
rect 1725 4316 1729 4320
rect 1745 4316 1749 4320
rect 1765 4316 1769 4320
rect 1865 4316 1869 4320
rect 1885 4316 1889 4320
rect 1905 4316 1909 4320
rect 1991 4316 1995 4320
rect 2011 4316 2015 4320
rect 2031 4316 2035 4320
rect 2131 4316 2135 4320
rect 2151 4316 2155 4320
rect 2171 4316 2175 4320
rect 2297 4316 2301 4320
rect 2305 4316 2309 4320
rect 2430 4316 2434 4320
rect 2452 4316 2456 4320
rect 2460 4316 2464 4320
rect 2585 4316 2589 4320
rect 2605 4316 2609 4320
rect 2625 4316 2629 4320
rect 2711 4316 2715 4320
rect 2831 4316 2835 4320
rect 2851 4316 2855 4320
rect 2871 4316 2875 4320
rect 2971 4316 2975 4320
rect 2991 4316 2995 4320
rect 3091 4316 3095 4320
rect 3111 4316 3115 4320
rect 3131 4316 3135 4320
rect 3231 4316 3235 4320
rect 3251 4316 3255 4320
rect 3271 4316 3275 4320
rect 3376 4316 3380 4320
rect 3384 4316 3388 4320
rect 3406 4316 3410 4320
rect 3531 4316 3535 4320
rect 3631 4316 3635 4320
rect 3651 4316 3655 4320
rect 3671 4316 3675 4320
rect 3771 4316 3775 4320
rect 3791 4316 3795 4320
rect 3811 4316 3815 4320
rect 3925 4316 3929 4320
rect 3945 4316 3949 4320
rect 4065 4316 4069 4320
rect 4085 4316 4089 4320
rect 4185 4316 4189 4320
rect 4205 4316 4209 4320
rect 4310 4316 4314 4320
rect 4332 4316 4336 4320
rect 4340 4316 4344 4320
rect 4431 4316 4435 4320
rect 4441 4316 4445 4320
rect 4461 4316 4465 4320
rect 4590 4316 4594 4320
rect 4612 4316 4616 4320
rect 4620 4316 4624 4320
rect 4736 4316 4740 4320
rect 4744 4316 4748 4320
rect 4766 4316 4770 4320
rect 4871 4316 4875 4320
rect 4879 4316 4883 4320
rect 4991 4316 4995 4320
rect 5111 4316 5115 4320
rect 5131 4316 5135 4320
rect 5151 4316 5155 4320
rect 5256 4316 5260 4320
rect 5264 4316 5268 4320
rect 5286 4316 5290 4320
rect 5391 4316 5395 4320
rect 5496 4316 5500 4320
rect 5504 4316 5508 4320
rect 5526 4316 5530 4320
rect 5595 4316 5599 4320
rect 5615 4316 5619 4320
rect 5629 4316 5633 4320
rect 5649 4316 5653 4320
rect 5661 4316 5665 4320
rect 5681 4316 5685 4320
rect 5727 4316 5731 4320
rect 5735 4316 5739 4320
rect 5755 4316 5759 4320
rect 5763 4316 5767 4320
rect 5785 4316 5789 4320
rect 110 4233 114 4276
rect 107 4221 114 4233
rect 105 4144 109 4221
rect 132 4179 136 4236
rect 140 4232 144 4236
rect 250 4233 254 4276
rect 140 4224 158 4232
rect 154 4213 158 4224
rect 247 4221 254 4233
rect 125 4167 134 4179
rect 125 4144 129 4167
rect 154 4156 158 4201
rect 145 4149 158 4156
rect 145 4144 149 4149
rect 245 4144 249 4221
rect 272 4179 276 4236
rect 280 4232 284 4236
rect 405 4233 409 4276
rect 425 4264 429 4276
rect 445 4268 449 4276
rect 445 4264 460 4268
rect 425 4260 440 4264
rect 434 4253 440 4260
rect 280 4224 298 4232
rect 294 4213 298 4224
rect 405 4221 413 4233
rect 425 4221 432 4233
rect 265 4167 274 4179
rect 265 4144 269 4167
rect 294 4156 298 4201
rect 428 4164 432 4221
rect 436 4164 440 4241
rect 454 4233 460 4264
rect 545 4233 549 4276
rect 565 4264 569 4276
rect 585 4268 589 4276
rect 585 4264 600 4268
rect 565 4260 580 4264
rect 574 4253 580 4260
rect 444 4221 454 4233
rect 545 4221 553 4233
rect 565 4221 572 4233
rect 444 4164 448 4221
rect 568 4164 572 4221
rect 576 4164 580 4241
rect 594 4233 600 4264
rect 584 4221 594 4233
rect 695 4231 699 4236
rect 584 4164 588 4221
rect 715 4213 719 4236
rect 725 4232 729 4236
rect 830 4233 834 4276
rect 725 4227 738 4232
rect 285 4149 298 4156
rect 285 4144 289 4149
rect 685 4152 695 4164
rect 685 4144 689 4152
rect 715 4137 719 4201
rect 705 4131 719 4137
rect 734 4193 738 4227
rect 827 4221 834 4233
rect 734 4136 738 4181
rect 825 4144 829 4221
rect 852 4179 856 4236
rect 860 4232 864 4236
rect 860 4224 878 4232
rect 874 4213 878 4224
rect 845 4167 854 4179
rect 845 4144 849 4167
rect 874 4156 878 4201
rect 951 4193 955 4276
rect 946 4181 955 4193
rect 865 4149 878 4156
rect 865 4144 869 4149
rect 725 4131 738 4136
rect 705 4124 709 4131
rect 725 4124 729 4131
rect 951 4124 955 4181
rect 1065 4179 1069 4236
rect 1085 4222 1089 4236
rect 1105 4222 1109 4236
rect 1225 4233 1229 4276
rect 1245 4264 1249 4276
rect 1265 4268 1269 4276
rect 1265 4264 1280 4268
rect 1245 4260 1260 4264
rect 1254 4253 1260 4260
rect 1085 4216 1100 4222
rect 1105 4216 1121 4222
rect 1225 4221 1233 4233
rect 1245 4221 1252 4233
rect 1094 4193 1100 4216
rect 1065 4167 1074 4179
rect 1072 4124 1076 4167
rect 1094 4144 1098 4181
rect 1114 4179 1121 4216
rect 1114 4154 1121 4167
rect 1248 4164 1252 4221
rect 1256 4164 1260 4241
rect 1274 4233 1280 4264
rect 1264 4221 1274 4233
rect 1264 4164 1268 4221
rect 1365 4199 1369 4276
rect 1366 4187 1369 4199
rect 1363 4171 1369 4187
rect 1385 4199 1389 4276
rect 1485 4199 1489 4276
rect 1385 4187 1394 4199
rect 1486 4187 1489 4199
rect 1385 4171 1391 4187
rect 1363 4164 1377 4171
rect 1102 4148 1121 4154
rect 1102 4144 1106 4148
rect 1373 4144 1377 4164
rect 1383 4164 1391 4171
rect 1483 4171 1489 4187
rect 1505 4199 1509 4276
rect 1617 4213 1621 4236
rect 1606 4201 1621 4213
rect 1625 4213 1629 4236
rect 1725 4233 1729 4276
rect 1745 4264 1749 4276
rect 1765 4268 1769 4276
rect 1765 4264 1780 4268
rect 1745 4260 1760 4264
rect 1754 4253 1760 4260
rect 1725 4221 1733 4233
rect 1745 4221 1752 4233
rect 1625 4201 1634 4213
rect 1505 4187 1514 4199
rect 1505 4171 1511 4187
rect 1483 4164 1497 4171
rect 1383 4144 1387 4164
rect 1493 4144 1497 4164
rect 1503 4164 1511 4171
rect 1503 4144 1507 4164
rect 1605 4124 1609 4201
rect 1625 4124 1629 4201
rect 1748 4164 1752 4221
rect 1756 4164 1760 4241
rect 1774 4233 1780 4264
rect 1865 4233 1869 4276
rect 1885 4264 1889 4276
rect 1905 4268 1909 4276
rect 1991 4268 1995 4276
rect 1905 4264 1920 4268
rect 1885 4260 1900 4264
rect 1894 4253 1900 4260
rect 1764 4221 1774 4233
rect 1865 4221 1873 4233
rect 1885 4221 1892 4233
rect 1764 4164 1768 4221
rect 1888 4164 1892 4221
rect 1896 4164 1900 4241
rect 1914 4233 1920 4264
rect 1980 4264 1995 4268
rect 2011 4264 2015 4276
rect 1980 4233 1986 4264
rect 2000 4260 2015 4264
rect 2000 4253 2006 4260
rect 1904 4221 1914 4233
rect 1986 4221 1996 4233
rect 1904 4164 1908 4221
rect 1992 4164 1996 4221
rect 2000 4164 2004 4241
rect 2031 4233 2035 4276
rect 2131 4268 2135 4276
rect 2120 4264 2135 4268
rect 2151 4264 2155 4276
rect 2120 4233 2126 4264
rect 2140 4260 2155 4264
rect 2140 4253 2146 4260
rect 2008 4221 2015 4233
rect 2027 4221 2035 4233
rect 2126 4221 2136 4233
rect 2008 4164 2012 4221
rect 2132 4164 2136 4221
rect 2140 4164 2144 4241
rect 2171 4233 2175 4276
rect 2148 4221 2155 4233
rect 2167 4221 2175 4233
rect 2148 4164 2152 4221
rect 2297 4213 2301 4236
rect 2286 4201 2301 4213
rect 2305 4213 2309 4236
rect 2430 4233 2434 4276
rect 2427 4221 2434 4233
rect 2305 4201 2314 4213
rect 2285 4124 2289 4201
rect 2305 4124 2309 4201
rect 2425 4144 2429 4221
rect 2452 4179 2456 4236
rect 2460 4232 2464 4236
rect 2585 4233 2589 4276
rect 2605 4264 2609 4276
rect 2625 4268 2629 4276
rect 2625 4264 2640 4268
rect 2605 4260 2620 4264
rect 2614 4253 2620 4260
rect 2460 4224 2478 4232
rect 2474 4213 2478 4224
rect 2585 4221 2593 4233
rect 2605 4221 2612 4233
rect 2445 4167 2454 4179
rect 2445 4144 2449 4167
rect 2474 4156 2478 4201
rect 2608 4164 2612 4221
rect 2616 4164 2620 4241
rect 2634 4233 2640 4264
rect 2624 4221 2634 4233
rect 2624 4164 2628 4221
rect 2711 4193 2715 4276
rect 2831 4268 2835 4276
rect 2820 4264 2835 4268
rect 2851 4264 2855 4276
rect 2820 4233 2826 4264
rect 2840 4260 2855 4264
rect 2840 4253 2846 4260
rect 2826 4221 2836 4233
rect 2706 4181 2715 4193
rect 2465 4149 2478 4156
rect 2465 4144 2469 4149
rect 2711 4124 2715 4181
rect 2832 4164 2836 4221
rect 2840 4164 2844 4241
rect 2871 4233 2875 4276
rect 2848 4221 2855 4233
rect 2867 4221 2875 4233
rect 2848 4164 2852 4221
rect 2971 4199 2975 4276
rect 2966 4187 2975 4199
rect 2969 4171 2975 4187
rect 2991 4199 2995 4276
rect 3091 4222 3095 4236
rect 3111 4222 3115 4236
rect 3079 4216 3095 4222
rect 3100 4216 3115 4222
rect 2991 4187 2994 4199
rect 2991 4171 2997 4187
rect 3079 4179 3086 4216
rect 3100 4193 3106 4216
rect 2969 4164 2977 4171
rect 2973 4144 2977 4164
rect 2983 4164 2997 4171
rect 2983 4144 2987 4164
rect 3079 4154 3086 4167
rect 3079 4148 3098 4154
rect 3094 4144 3098 4148
rect 3102 4144 3106 4181
rect 3131 4179 3135 4236
rect 3231 4222 3235 4236
rect 3251 4222 3255 4236
rect 3219 4216 3235 4222
rect 3240 4216 3255 4222
rect 3219 4179 3226 4216
rect 3240 4193 3246 4216
rect 3126 4167 3135 4179
rect 3124 4124 3128 4167
rect 3219 4154 3226 4167
rect 3219 4148 3238 4154
rect 3234 4144 3238 4148
rect 3242 4144 3246 4181
rect 3271 4179 3275 4236
rect 3376 4232 3380 4236
rect 3362 4224 3380 4232
rect 3362 4213 3366 4224
rect 3266 4167 3275 4179
rect 3264 4124 3268 4167
rect 3362 4156 3366 4201
rect 3384 4179 3388 4236
rect 3406 4233 3410 4276
rect 3406 4221 3413 4233
rect 3386 4167 3395 4179
rect 3362 4149 3375 4156
rect 3371 4144 3375 4149
rect 3391 4144 3395 4167
rect 3411 4144 3415 4221
rect 3531 4193 3535 4276
rect 3631 4268 3635 4276
rect 3620 4264 3635 4268
rect 3651 4264 3655 4276
rect 3620 4233 3626 4264
rect 3640 4260 3655 4264
rect 3640 4253 3646 4260
rect 3626 4221 3636 4233
rect 3526 4181 3535 4193
rect 3531 4124 3535 4181
rect 3632 4164 3636 4221
rect 3640 4164 3644 4241
rect 3671 4233 3675 4276
rect 3771 4268 3775 4276
rect 3760 4264 3775 4268
rect 3791 4264 3795 4276
rect 3760 4233 3766 4264
rect 3780 4260 3795 4264
rect 3780 4253 3786 4260
rect 3648 4221 3655 4233
rect 3667 4221 3675 4233
rect 3766 4221 3776 4233
rect 3648 4164 3652 4221
rect 3772 4164 3776 4221
rect 3780 4164 3784 4241
rect 3811 4233 3815 4276
rect 3788 4221 3795 4233
rect 3807 4221 3815 4233
rect 3788 4164 3792 4221
rect 3925 4199 3929 4276
rect 3926 4187 3929 4199
rect 3923 4171 3929 4187
rect 3945 4199 3949 4276
rect 4065 4199 4069 4276
rect 3945 4187 3954 4199
rect 4066 4187 4069 4199
rect 3945 4171 3951 4187
rect 3923 4164 3937 4171
rect 3933 4144 3937 4164
rect 3943 4164 3951 4171
rect 4063 4171 4069 4187
rect 4085 4199 4089 4276
rect 4185 4199 4189 4276
rect 4085 4187 4094 4199
rect 4186 4187 4189 4199
rect 4085 4171 4091 4187
rect 4063 4164 4077 4171
rect 3943 4144 3947 4164
rect 4073 4144 4077 4164
rect 4083 4164 4091 4171
rect 4183 4171 4189 4187
rect 4205 4199 4209 4276
rect 4310 4233 4314 4276
rect 4307 4221 4314 4233
rect 4205 4187 4214 4199
rect 4205 4171 4211 4187
rect 4183 4164 4197 4171
rect 4083 4144 4087 4164
rect 4193 4144 4197 4164
rect 4203 4164 4211 4171
rect 4203 4144 4207 4164
rect 4305 4144 4309 4221
rect 4332 4179 4336 4236
rect 4340 4232 4344 4236
rect 4431 4232 4435 4236
rect 4340 4224 4358 4232
rect 4354 4213 4358 4224
rect 4422 4227 4435 4232
rect 4325 4167 4334 4179
rect 4325 4144 4329 4167
rect 4354 4156 4358 4201
rect 4422 4193 4426 4227
rect 4441 4213 4445 4236
rect 4461 4231 4465 4236
rect 4590 4233 4594 4276
rect 4587 4221 4594 4233
rect 4345 4149 4358 4156
rect 4345 4144 4349 4149
rect 4422 4136 4426 4181
rect 4441 4137 4445 4201
rect 4465 4152 4475 4164
rect 4471 4144 4475 4152
rect 4585 4144 4589 4221
rect 4612 4179 4616 4236
rect 4620 4232 4624 4236
rect 4736 4232 4740 4236
rect 4620 4224 4638 4232
rect 4634 4213 4638 4224
rect 4722 4224 4740 4232
rect 4722 4213 4726 4224
rect 4605 4167 4614 4179
rect 4605 4144 4609 4167
rect 4634 4156 4638 4201
rect 4625 4149 4638 4156
rect 4722 4156 4726 4201
rect 4744 4179 4748 4236
rect 4766 4233 4770 4276
rect 4766 4221 4773 4233
rect 4746 4167 4755 4179
rect 4722 4149 4735 4156
rect 4625 4144 4629 4149
rect 4731 4144 4735 4149
rect 4751 4144 4755 4167
rect 4771 4144 4775 4221
rect 4871 4213 4875 4236
rect 4866 4201 4875 4213
rect 4879 4213 4883 4236
rect 4879 4201 4894 4213
rect 4422 4131 4435 4136
rect 4441 4131 4455 4137
rect 4431 4124 4435 4131
rect 4451 4124 4455 4131
rect 4871 4124 4875 4201
rect 4891 4124 4895 4201
rect 4991 4193 4995 4276
rect 5111 4222 5115 4236
rect 5131 4222 5135 4236
rect 4986 4181 4995 4193
rect 4991 4124 4995 4181
rect 5099 4216 5115 4222
rect 5120 4216 5135 4222
rect 5099 4179 5106 4216
rect 5120 4193 5126 4216
rect 5099 4154 5106 4167
rect 5099 4148 5118 4154
rect 5114 4144 5118 4148
rect 5122 4144 5126 4181
rect 5151 4179 5155 4236
rect 5256 4232 5260 4236
rect 5242 4224 5260 4232
rect 5242 4213 5246 4224
rect 5146 4167 5155 4179
rect 5144 4124 5148 4167
rect 5242 4156 5246 4201
rect 5264 4179 5268 4236
rect 5286 4233 5290 4276
rect 5286 4221 5293 4233
rect 5266 4167 5275 4179
rect 5242 4149 5255 4156
rect 5251 4144 5255 4149
rect 5271 4144 5275 4167
rect 5291 4144 5295 4221
rect 5391 4193 5395 4276
rect 5496 4232 5500 4236
rect 5482 4224 5500 4232
rect 5482 4213 5486 4224
rect 5386 4181 5395 4193
rect 5391 4124 5395 4181
rect 5482 4156 5486 4201
rect 5504 4179 5508 4236
rect 5526 4233 5530 4276
rect 5526 4221 5533 4233
rect 5506 4167 5515 4179
rect 5482 4149 5495 4156
rect 5491 4144 5495 4149
rect 5511 4144 5515 4167
rect 5531 4144 5535 4221
rect 5595 4193 5599 4236
rect 5615 4194 5619 4276
rect 5629 4217 5633 4276
rect 5649 4236 5653 4276
rect 5661 4270 5665 4276
rect 5655 4224 5658 4236
rect 5629 4209 5638 4217
rect 5595 4144 5599 4181
rect 5615 4124 5619 4182
rect 5634 4180 5638 4209
rect 5654 4160 5658 4224
rect 5625 4156 5658 4160
rect 5625 4124 5629 4156
rect 5663 4148 5667 4258
rect 5681 4250 5685 4276
rect 5727 4272 5731 4276
rect 5695 4270 5731 4272
rect 5707 4268 5731 4270
rect 5649 4136 5651 4148
rect 5647 4124 5651 4136
rect 5657 4136 5659 4148
rect 5657 4124 5661 4136
rect 5679 4124 5683 4238
rect 5695 4132 5699 4258
rect 5735 4244 5739 4276
rect 5755 4256 5759 4296
rect 5763 4273 5767 4296
rect 5763 4266 5771 4273
rect 5733 4149 5739 4244
rect 5767 4237 5771 4266
rect 5763 4231 5771 4237
rect 5763 4185 5767 4231
rect 5785 4224 5789 4236
rect 5787 4212 5789 4224
rect 5733 4145 5757 4149
rect 5719 4140 5737 4141
rect 5707 4136 5737 4140
rect 5695 4128 5729 4132
rect 5725 4124 5729 4128
rect 5733 4124 5737 4136
rect 5753 4124 5757 4145
rect 5763 4124 5767 4173
rect 5785 4144 5789 4212
rect 105 4100 109 4104
rect 125 4100 129 4104
rect 145 4100 149 4104
rect 245 4100 249 4104
rect 265 4100 269 4104
rect 285 4100 289 4104
rect 428 4100 432 4104
rect 436 4100 440 4104
rect 444 4100 448 4104
rect 568 4100 572 4104
rect 576 4100 580 4104
rect 584 4100 588 4104
rect 685 4100 689 4104
rect 705 4100 709 4104
rect 725 4100 729 4104
rect 825 4100 829 4104
rect 845 4100 849 4104
rect 865 4100 869 4104
rect 951 4100 955 4104
rect 1072 4100 1076 4104
rect 1094 4100 1098 4104
rect 1102 4100 1106 4104
rect 1248 4100 1252 4104
rect 1256 4100 1260 4104
rect 1264 4100 1268 4104
rect 1373 4100 1377 4104
rect 1383 4100 1387 4104
rect 1493 4100 1497 4104
rect 1503 4100 1507 4104
rect 1605 4100 1609 4104
rect 1625 4100 1629 4104
rect 1748 4100 1752 4104
rect 1756 4100 1760 4104
rect 1764 4100 1768 4104
rect 1888 4100 1892 4104
rect 1896 4100 1900 4104
rect 1904 4100 1908 4104
rect 1992 4100 1996 4104
rect 2000 4100 2004 4104
rect 2008 4100 2012 4104
rect 2132 4100 2136 4104
rect 2140 4100 2144 4104
rect 2148 4100 2152 4104
rect 2285 4100 2289 4104
rect 2305 4100 2309 4104
rect 2425 4100 2429 4104
rect 2445 4100 2449 4104
rect 2465 4100 2469 4104
rect 2608 4100 2612 4104
rect 2616 4100 2620 4104
rect 2624 4100 2628 4104
rect 2711 4100 2715 4104
rect 2832 4100 2836 4104
rect 2840 4100 2844 4104
rect 2848 4100 2852 4104
rect 2973 4100 2977 4104
rect 2983 4100 2987 4104
rect 3094 4100 3098 4104
rect 3102 4100 3106 4104
rect 3124 4100 3128 4104
rect 3234 4100 3238 4104
rect 3242 4100 3246 4104
rect 3264 4100 3268 4104
rect 3371 4100 3375 4104
rect 3391 4100 3395 4104
rect 3411 4100 3415 4104
rect 3531 4100 3535 4104
rect 3632 4100 3636 4104
rect 3640 4100 3644 4104
rect 3648 4100 3652 4104
rect 3772 4100 3776 4104
rect 3780 4100 3784 4104
rect 3788 4100 3792 4104
rect 3933 4100 3937 4104
rect 3943 4100 3947 4104
rect 4073 4100 4077 4104
rect 4083 4100 4087 4104
rect 4193 4100 4197 4104
rect 4203 4100 4207 4104
rect 4305 4100 4309 4104
rect 4325 4100 4329 4104
rect 4345 4100 4349 4104
rect 4431 4100 4435 4104
rect 4451 4100 4455 4104
rect 4471 4100 4475 4104
rect 4585 4100 4589 4104
rect 4605 4100 4609 4104
rect 4625 4100 4629 4104
rect 4731 4100 4735 4104
rect 4751 4100 4755 4104
rect 4771 4100 4775 4104
rect 4871 4100 4875 4104
rect 4891 4100 4895 4104
rect 4991 4100 4995 4104
rect 5114 4100 5118 4104
rect 5122 4100 5126 4104
rect 5144 4100 5148 4104
rect 5251 4100 5255 4104
rect 5271 4100 5275 4104
rect 5291 4100 5295 4104
rect 5391 4100 5395 4104
rect 5491 4100 5495 4104
rect 5511 4100 5515 4104
rect 5531 4100 5535 4104
rect 5595 4100 5599 4104
rect 5615 4100 5619 4104
rect 5625 4100 5629 4104
rect 5647 4100 5651 4104
rect 5657 4100 5661 4104
rect 5679 4100 5683 4104
rect 5725 4100 5729 4104
rect 5733 4100 5737 4104
rect 5753 4100 5757 4104
rect 5763 4100 5767 4104
rect 5785 4100 5789 4104
rect 85 4076 89 4080
rect 191 4076 195 4080
rect 211 4076 215 4080
rect 231 4076 235 4080
rect 345 4076 349 4080
rect 454 4076 458 4080
rect 462 4076 466 4080
rect 484 4076 488 4080
rect 605 4076 609 4080
rect 625 4076 629 4080
rect 745 4076 749 4080
rect 831 4076 835 4080
rect 851 4076 855 4080
rect 871 4076 875 4080
rect 971 4076 975 4080
rect 1072 4076 1076 4080
rect 1080 4076 1084 4080
rect 1088 4076 1092 4080
rect 1214 4076 1218 4080
rect 1222 4076 1226 4080
rect 1242 4076 1246 4080
rect 1250 4076 1254 4080
rect 1393 4076 1397 4080
rect 1403 4076 1407 4080
rect 1525 4076 1529 4080
rect 1625 4076 1629 4080
rect 1645 4076 1649 4080
rect 1745 4076 1749 4080
rect 1832 4076 1836 4080
rect 1840 4076 1844 4080
rect 1848 4076 1852 4080
rect 1985 4076 1989 4080
rect 2005 4076 2009 4080
rect 2025 4076 2029 4080
rect 2168 4076 2172 4080
rect 2176 4076 2180 4080
rect 2184 4076 2188 4080
rect 2272 4076 2276 4080
rect 2280 4076 2284 4080
rect 2288 4076 2292 4080
rect 2425 4076 2429 4080
rect 2445 4076 2449 4080
rect 2465 4076 2469 4080
rect 2573 4076 2577 4080
rect 2583 4076 2587 4080
rect 2673 4076 2677 4080
rect 2683 4076 2687 4080
rect 2792 4076 2796 4080
rect 2800 4076 2804 4080
rect 2808 4076 2812 4080
rect 2932 4076 2936 4080
rect 2940 4076 2944 4080
rect 2948 4076 2952 4080
rect 3085 4076 3089 4080
rect 3208 4076 3212 4080
rect 3216 4076 3220 4080
rect 3224 4076 3228 4080
rect 3325 4076 3329 4080
rect 3425 4076 3429 4080
rect 3445 4076 3449 4080
rect 3465 4076 3469 4080
rect 3553 4076 3557 4080
rect 3563 4076 3567 4080
rect 3685 4076 3689 4080
rect 3705 4076 3709 4080
rect 3725 4076 3729 4080
rect 3833 4076 3837 4080
rect 3843 4076 3847 4080
rect 3965 4076 3969 4080
rect 3985 4076 3989 4080
rect 4005 4076 4009 4080
rect 4112 4076 4116 4080
rect 4134 4076 4138 4080
rect 4142 4076 4146 4080
rect 4233 4076 4237 4080
rect 4243 4076 4247 4080
rect 4351 4076 4355 4080
rect 4371 4076 4375 4080
rect 4391 4076 4395 4080
rect 4491 4076 4495 4080
rect 4511 4076 4515 4080
rect 4531 4076 4535 4080
rect 4631 4076 4635 4080
rect 4651 4076 4655 4080
rect 4671 4076 4675 4080
rect 4793 4076 4797 4080
rect 4803 4076 4807 4080
rect 4892 4076 4896 4080
rect 4900 4076 4904 4080
rect 4908 4076 4912 4080
rect 5031 4076 5035 4080
rect 5145 4076 5149 4080
rect 5191 4076 5195 4080
rect 5213 4076 5217 4080
rect 5223 4076 5227 4080
rect 5243 4076 5247 4080
rect 5251 4076 5255 4080
rect 5297 4076 5301 4080
rect 5319 4076 5323 4080
rect 5329 4076 5333 4080
rect 5351 4076 5355 4080
rect 5361 4076 5365 4080
rect 5381 4076 5385 4080
rect 5431 4076 5435 4080
rect 5453 4076 5457 4080
rect 5463 4076 5467 4080
rect 5483 4076 5487 4080
rect 5491 4076 5495 4080
rect 5537 4076 5541 4080
rect 5559 4076 5563 4080
rect 5569 4076 5573 4080
rect 5591 4076 5595 4080
rect 5601 4076 5605 4080
rect 5621 4076 5625 4080
rect 5711 4076 5715 4080
rect 5731 4076 5735 4080
rect 5751 4076 5755 4080
rect 85 3999 89 4056
rect 191 4031 195 4036
rect 182 4024 195 4031
rect 85 3987 94 3999
rect 85 3904 89 3987
rect 182 3979 186 4024
rect 211 4013 215 4036
rect 206 4001 215 4013
rect 182 3956 186 3967
rect 182 3948 200 3956
rect 196 3944 200 3948
rect 204 3944 208 4001
rect 231 3959 235 4036
rect 345 3999 349 4056
rect 454 4032 458 4036
rect 439 4026 458 4032
rect 439 4013 446 4026
rect 345 3987 354 3999
rect 226 3947 233 3959
rect 226 3904 230 3947
rect 345 3904 349 3987
rect 439 3964 446 4001
rect 462 3999 466 4036
rect 484 4013 488 4056
rect 486 4001 495 4013
rect 460 3964 466 3987
rect 439 3958 455 3964
rect 460 3958 475 3964
rect 451 3944 455 3958
rect 471 3944 475 3958
rect 491 3944 495 4001
rect 605 3979 609 4056
rect 625 3979 629 4056
rect 745 3999 749 4056
rect 831 4031 835 4036
rect 822 4024 835 4031
rect 745 3987 754 3999
rect 606 3967 621 3979
rect 617 3944 621 3967
rect 625 3967 634 3979
rect 625 3944 629 3967
rect 745 3904 749 3987
rect 822 3979 826 4024
rect 851 4013 855 4036
rect 846 4001 855 4013
rect 822 3956 826 3967
rect 822 3948 840 3956
rect 836 3944 840 3948
rect 844 3944 848 4001
rect 871 3959 875 4036
rect 971 3999 975 4056
rect 1214 4028 1218 4036
rect 1201 4021 1218 4028
rect 966 3987 975 3999
rect 866 3947 873 3959
rect 866 3904 870 3947
rect 971 3904 975 3987
rect 1072 3959 1076 4016
rect 1066 3947 1076 3959
rect 1060 3916 1066 3947
rect 1080 3939 1084 4016
rect 1088 3959 1092 4016
rect 1201 3979 1207 4021
rect 1222 4013 1226 4036
rect 1242 4022 1246 4036
rect 1250 4031 1254 4036
rect 1250 4027 1280 4031
rect 1242 4015 1255 4022
rect 1251 4013 1255 4015
rect 1251 4001 1253 4013
rect 1222 3972 1226 4001
rect 1207 3967 1215 3972
rect 1195 3966 1215 3967
rect 1222 3966 1235 3972
rect 1088 3947 1095 3959
rect 1107 3947 1115 3959
rect 1080 3920 1086 3927
rect 1080 3916 1095 3920
rect 1060 3912 1075 3916
rect 1071 3904 1075 3912
rect 1091 3904 1095 3916
rect 1111 3904 1115 3947
rect 1211 3944 1215 3966
rect 1231 3944 1235 3966
rect 1251 3944 1255 4001
rect 1274 3979 1280 4027
rect 1393 4016 1397 4036
rect 1389 4009 1397 4016
rect 1403 4016 1407 4036
rect 1403 4009 1417 4016
rect 1389 3993 1395 4009
rect 1386 3981 1395 3993
rect 1271 3967 1274 3979
rect 1271 3944 1275 3967
rect 1391 3904 1395 3981
rect 1411 3993 1417 4009
rect 1525 3999 1529 4056
rect 1411 3981 1414 3993
rect 1525 3987 1534 3999
rect 1411 3904 1415 3981
rect 1525 3904 1529 3987
rect 1625 3979 1629 4056
rect 1645 3979 1649 4056
rect 1745 3999 1749 4056
rect 1745 3987 1754 3999
rect 1626 3967 1641 3979
rect 1637 3944 1641 3967
rect 1645 3967 1654 3979
rect 1645 3944 1649 3967
rect 1745 3904 1749 3987
rect 1832 3959 1836 4016
rect 1826 3947 1836 3959
rect 1820 3916 1826 3947
rect 1840 3939 1844 4016
rect 1848 3959 1852 4016
rect 1985 3959 1989 4036
rect 2005 4013 2009 4036
rect 2025 4031 2029 4036
rect 2025 4024 2038 4031
rect 2005 4001 2014 4013
rect 1848 3947 1855 3959
rect 1867 3947 1875 3959
rect 1987 3947 1994 3959
rect 1840 3920 1846 3927
rect 1840 3916 1855 3920
rect 1820 3912 1835 3916
rect 1831 3904 1835 3912
rect 1851 3904 1855 3916
rect 1871 3904 1875 3947
rect 1990 3904 1994 3947
rect 2012 3944 2016 4001
rect 2034 3979 2038 4024
rect 2034 3956 2038 3967
rect 2168 3959 2172 4016
rect 2020 3948 2038 3956
rect 2020 3944 2024 3948
rect 2145 3947 2153 3959
rect 2165 3947 2172 3959
rect 2145 3904 2149 3947
rect 2176 3939 2180 4016
rect 2184 3959 2188 4016
rect 2272 3959 2276 4016
rect 2184 3947 2194 3959
rect 2266 3947 2276 3959
rect 2174 3920 2180 3927
rect 2165 3916 2180 3920
rect 2194 3916 2200 3947
rect 2165 3904 2169 3916
rect 2185 3912 2200 3916
rect 2260 3916 2266 3947
rect 2280 3939 2284 4016
rect 2288 3959 2292 4016
rect 2425 3959 2429 4036
rect 2445 4013 2449 4036
rect 2465 4031 2469 4036
rect 2465 4024 2478 4031
rect 2445 4001 2454 4013
rect 2288 3947 2295 3959
rect 2307 3947 2315 3959
rect 2427 3947 2434 3959
rect 2280 3920 2286 3927
rect 2280 3916 2295 3920
rect 2260 3912 2275 3916
rect 2185 3904 2189 3912
rect 2271 3904 2275 3912
rect 2291 3904 2295 3916
rect 2311 3904 2315 3947
rect 2430 3904 2434 3947
rect 2452 3944 2456 4001
rect 2474 3979 2478 4024
rect 2573 4016 2577 4036
rect 2563 4009 2577 4016
rect 2583 4016 2587 4036
rect 2673 4016 2677 4036
rect 2583 4009 2591 4016
rect 2563 3993 2569 4009
rect 2566 3981 2569 3993
rect 2474 3956 2478 3967
rect 2460 3948 2478 3956
rect 2460 3944 2464 3948
rect 2565 3904 2569 3981
rect 2585 3993 2591 4009
rect 2669 4009 2677 4016
rect 2683 4016 2687 4036
rect 2683 4009 2697 4016
rect 2669 3993 2675 4009
rect 2585 3981 2594 3993
rect 2666 3981 2675 3993
rect 2585 3904 2589 3981
rect 2671 3904 2675 3981
rect 2691 3993 2697 4009
rect 2691 3981 2694 3993
rect 2691 3904 2695 3981
rect 2792 3959 2796 4016
rect 2786 3947 2796 3959
rect 2780 3916 2786 3947
rect 2800 3939 2804 4016
rect 2808 3959 2812 4016
rect 2932 3959 2936 4016
rect 2808 3947 2815 3959
rect 2827 3947 2835 3959
rect 2926 3947 2936 3959
rect 2800 3920 2806 3927
rect 2800 3916 2815 3920
rect 2780 3912 2795 3916
rect 2791 3904 2795 3912
rect 2811 3904 2815 3916
rect 2831 3904 2835 3947
rect 2920 3916 2926 3947
rect 2940 3939 2944 4016
rect 2948 3959 2952 4016
rect 3085 3999 3089 4056
rect 3085 3987 3094 3999
rect 2948 3947 2955 3959
rect 2967 3947 2975 3959
rect 2940 3920 2946 3927
rect 2940 3916 2955 3920
rect 2920 3912 2935 3916
rect 2931 3904 2935 3912
rect 2951 3904 2955 3916
rect 2971 3904 2975 3947
rect 3085 3904 3089 3987
rect 3208 3959 3212 4016
rect 3185 3947 3193 3959
rect 3205 3947 3212 3959
rect 3185 3904 3189 3947
rect 3216 3939 3220 4016
rect 3224 3959 3228 4016
rect 3325 3999 3329 4056
rect 3705 4049 3709 4056
rect 3725 4049 3729 4056
rect 3705 4043 3719 4049
rect 3725 4044 3738 4049
rect 3325 3987 3334 3999
rect 3224 3947 3234 3959
rect 3214 3920 3220 3927
rect 3205 3916 3220 3920
rect 3234 3916 3240 3947
rect 3205 3904 3209 3916
rect 3225 3912 3240 3916
rect 3225 3904 3229 3912
rect 3325 3904 3329 3987
rect 3425 3959 3429 4036
rect 3445 4013 3449 4036
rect 3465 4031 3469 4036
rect 3465 4024 3478 4031
rect 3445 4001 3454 4013
rect 3427 3947 3434 3959
rect 3430 3904 3434 3947
rect 3452 3944 3456 4001
rect 3474 3979 3478 4024
rect 3553 4016 3557 4036
rect 3549 4009 3557 4016
rect 3563 4016 3567 4036
rect 3685 4028 3689 4036
rect 3685 4016 3695 4028
rect 3563 4009 3577 4016
rect 3549 3993 3555 4009
rect 3546 3981 3555 3993
rect 3474 3956 3478 3967
rect 3460 3948 3478 3956
rect 3460 3944 3464 3948
rect 3551 3904 3555 3981
rect 3571 3993 3577 4009
rect 3571 3981 3574 3993
rect 3571 3904 3575 3981
rect 3715 3979 3719 4043
rect 3734 3999 3738 4044
rect 3833 4016 3837 4036
rect 3829 4009 3837 4016
rect 3843 4016 3847 4036
rect 3843 4009 3857 4016
rect 3829 3993 3835 4009
rect 3695 3944 3699 3949
rect 3715 3944 3719 3967
rect 3734 3953 3738 3987
rect 3826 3981 3835 3993
rect 3725 3948 3738 3953
rect 3725 3944 3729 3948
rect 3831 3904 3835 3981
rect 3851 3993 3857 4009
rect 3851 3981 3854 3993
rect 3851 3904 3855 3981
rect 3965 3959 3969 4036
rect 3985 4013 3989 4036
rect 4005 4031 4009 4036
rect 4005 4024 4018 4031
rect 3985 4001 3994 4013
rect 3967 3947 3974 3959
rect 3970 3904 3974 3947
rect 3992 3944 3996 4001
rect 4014 3979 4018 4024
rect 4112 4013 4116 4056
rect 4631 4049 4635 4056
rect 4651 4049 4655 4056
rect 4622 4044 4635 4049
rect 4105 4001 4114 4013
rect 4014 3956 4018 3967
rect 4000 3948 4018 3956
rect 4000 3944 4004 3948
rect 4105 3944 4109 4001
rect 4134 3999 4138 4036
rect 4142 4032 4146 4036
rect 4142 4026 4161 4032
rect 4154 4013 4161 4026
rect 4233 4016 4237 4036
rect 4229 4009 4237 4016
rect 4243 4016 4247 4036
rect 4351 4031 4355 4036
rect 4342 4024 4355 4031
rect 4243 4009 4257 4016
rect 4134 3964 4140 3987
rect 4154 3964 4161 4001
rect 4229 3993 4235 4009
rect 4226 3981 4235 3993
rect 4125 3958 4140 3964
rect 4145 3958 4161 3964
rect 4125 3944 4129 3958
rect 4145 3944 4149 3958
rect 4231 3904 4235 3981
rect 4251 3993 4257 4009
rect 4251 3981 4254 3993
rect 4251 3904 4255 3981
rect 4342 3979 4346 4024
rect 4371 4013 4375 4036
rect 4366 4001 4375 4013
rect 4342 3956 4346 3967
rect 4342 3948 4360 3956
rect 4356 3944 4360 3948
rect 4364 3944 4368 4001
rect 4391 3959 4395 4036
rect 4491 4031 4495 4036
rect 4482 4024 4495 4031
rect 4482 3979 4486 4024
rect 4511 4013 4515 4036
rect 4506 4001 4515 4013
rect 4386 3947 4393 3959
rect 4482 3956 4486 3967
rect 4482 3948 4500 3956
rect 4386 3904 4390 3947
rect 4496 3944 4500 3948
rect 4504 3944 4508 4001
rect 4531 3959 4535 4036
rect 4622 3999 4626 4044
rect 4526 3947 4533 3959
rect 4622 3953 4626 3987
rect 4641 4043 4655 4049
rect 4641 3979 4645 4043
rect 4671 4028 4675 4036
rect 4665 4016 4675 4028
rect 4793 4016 4797 4036
rect 4783 4009 4797 4016
rect 4803 4016 4807 4036
rect 4803 4009 4811 4016
rect 4783 3993 4789 4009
rect 4786 3981 4789 3993
rect 4622 3948 4635 3953
rect 4526 3904 4530 3947
rect 4631 3944 4635 3948
rect 4641 3944 4645 3967
rect 4661 3944 4665 3949
rect 4785 3904 4789 3981
rect 4805 3993 4811 4009
rect 4805 3981 4814 3993
rect 4805 3904 4809 3981
rect 4892 3959 4896 4016
rect 4886 3947 4896 3959
rect 4880 3916 4886 3947
rect 4900 3939 4904 4016
rect 4908 3959 4912 4016
rect 5031 3999 5035 4056
rect 5026 3987 5035 3999
rect 4908 3947 4915 3959
rect 4927 3947 4935 3959
rect 4900 3920 4906 3927
rect 4900 3916 4915 3920
rect 4880 3912 4895 3916
rect 4891 3904 4895 3912
rect 4911 3904 4915 3916
rect 4931 3904 4935 3947
rect 5031 3904 5035 3987
rect 5145 3999 5149 4056
rect 5145 3987 5154 3999
rect 5145 3904 5149 3987
rect 5191 3968 5195 4036
rect 5213 4007 5217 4056
rect 5223 4035 5227 4056
rect 5243 4044 5247 4056
rect 5251 4052 5255 4056
rect 5251 4048 5285 4052
rect 5243 4040 5273 4044
rect 5243 4039 5261 4040
rect 5223 4031 5247 4035
rect 5191 3956 5193 3968
rect 5191 3944 5195 3956
rect 5213 3949 5217 3995
rect 5209 3943 5217 3949
rect 5209 3914 5213 3943
rect 5241 3936 5247 4031
rect 5209 3907 5217 3914
rect 5213 3884 5217 3907
rect 5221 3884 5225 3924
rect 5241 3904 5245 3936
rect 5281 3922 5285 4048
rect 5297 3942 5301 4056
rect 5319 4044 5323 4056
rect 5321 4032 5323 4044
rect 5329 4044 5333 4056
rect 5329 4032 5331 4044
rect 5249 3910 5273 3912
rect 5249 3908 5285 3910
rect 5249 3904 5253 3908
rect 5295 3904 5299 3930
rect 5313 3922 5317 4032
rect 5351 4024 5355 4056
rect 5322 4020 5355 4024
rect 5322 3956 5326 4020
rect 5342 3971 5346 4000
rect 5361 3998 5365 4056
rect 5381 3999 5385 4036
rect 5342 3963 5351 3971
rect 5322 3944 5325 3956
rect 5315 3904 5319 3910
rect 5327 3904 5331 3944
rect 5347 3904 5351 3963
rect 5361 3904 5365 3986
rect 5381 3944 5385 3987
rect 5431 3968 5435 4036
rect 5453 4007 5457 4056
rect 5463 4035 5467 4056
rect 5483 4044 5487 4056
rect 5491 4052 5495 4056
rect 5491 4048 5525 4052
rect 5483 4040 5513 4044
rect 5483 4039 5501 4040
rect 5463 4031 5487 4035
rect 5431 3956 5433 3968
rect 5431 3944 5435 3956
rect 5453 3949 5457 3995
rect 5449 3943 5457 3949
rect 5449 3914 5453 3943
rect 5481 3936 5487 4031
rect 5449 3907 5457 3914
rect 5453 3884 5457 3907
rect 5461 3884 5465 3924
rect 5481 3904 5485 3936
rect 5521 3922 5525 4048
rect 5537 3942 5541 4056
rect 5559 4044 5563 4056
rect 5561 4032 5563 4044
rect 5569 4044 5573 4056
rect 5569 4032 5571 4044
rect 5489 3910 5513 3912
rect 5489 3908 5525 3910
rect 5489 3904 5493 3908
rect 5535 3904 5539 3930
rect 5553 3922 5557 4032
rect 5591 4024 5595 4056
rect 5562 4020 5595 4024
rect 5562 3956 5566 4020
rect 5582 3971 5586 4000
rect 5601 3998 5605 4056
rect 5621 3999 5625 4036
rect 5711 4031 5715 4036
rect 5702 4024 5715 4031
rect 5582 3963 5591 3971
rect 5562 3944 5565 3956
rect 5555 3904 5559 3910
rect 5567 3904 5571 3944
rect 5587 3904 5591 3963
rect 5601 3904 5605 3986
rect 5621 3944 5625 3987
rect 5702 3979 5706 4024
rect 5731 4013 5735 4036
rect 5726 4001 5735 4013
rect 5702 3956 5706 3967
rect 5702 3948 5720 3956
rect 5716 3944 5720 3948
rect 5724 3944 5728 4001
rect 5751 3959 5755 4036
rect 5746 3947 5753 3959
rect 5746 3904 5750 3947
rect 85 3860 89 3864
rect 196 3860 200 3864
rect 204 3860 208 3864
rect 226 3860 230 3864
rect 345 3860 349 3864
rect 451 3860 455 3864
rect 471 3860 475 3864
rect 491 3860 495 3864
rect 617 3860 621 3864
rect 625 3860 629 3864
rect 745 3860 749 3864
rect 836 3860 840 3864
rect 844 3860 848 3864
rect 866 3860 870 3864
rect 971 3860 975 3864
rect 1071 3860 1075 3864
rect 1091 3860 1095 3864
rect 1111 3860 1115 3864
rect 1211 3860 1215 3864
rect 1231 3860 1235 3864
rect 1251 3860 1255 3864
rect 1271 3860 1275 3864
rect 1391 3860 1395 3864
rect 1411 3860 1415 3864
rect 1525 3860 1529 3864
rect 1637 3860 1641 3864
rect 1645 3860 1649 3864
rect 1745 3860 1749 3864
rect 1831 3860 1835 3864
rect 1851 3860 1855 3864
rect 1871 3860 1875 3864
rect 1990 3860 1994 3864
rect 2012 3860 2016 3864
rect 2020 3860 2024 3864
rect 2145 3860 2149 3864
rect 2165 3860 2169 3864
rect 2185 3860 2189 3864
rect 2271 3860 2275 3864
rect 2291 3860 2295 3864
rect 2311 3860 2315 3864
rect 2430 3860 2434 3864
rect 2452 3860 2456 3864
rect 2460 3860 2464 3864
rect 2565 3860 2569 3864
rect 2585 3860 2589 3864
rect 2671 3860 2675 3864
rect 2691 3860 2695 3864
rect 2791 3860 2795 3864
rect 2811 3860 2815 3864
rect 2831 3860 2835 3864
rect 2931 3860 2935 3864
rect 2951 3860 2955 3864
rect 2971 3860 2975 3864
rect 3085 3860 3089 3864
rect 3185 3860 3189 3864
rect 3205 3860 3209 3864
rect 3225 3860 3229 3864
rect 3325 3860 3329 3864
rect 3430 3860 3434 3864
rect 3452 3860 3456 3864
rect 3460 3860 3464 3864
rect 3551 3860 3555 3864
rect 3571 3860 3575 3864
rect 3695 3860 3699 3864
rect 3715 3860 3719 3864
rect 3725 3860 3729 3864
rect 3831 3860 3835 3864
rect 3851 3860 3855 3864
rect 3970 3860 3974 3864
rect 3992 3860 3996 3864
rect 4000 3860 4004 3864
rect 4105 3860 4109 3864
rect 4125 3860 4129 3864
rect 4145 3860 4149 3864
rect 4231 3860 4235 3864
rect 4251 3860 4255 3864
rect 4356 3860 4360 3864
rect 4364 3860 4368 3864
rect 4386 3860 4390 3864
rect 4496 3860 4500 3864
rect 4504 3860 4508 3864
rect 4526 3860 4530 3864
rect 4631 3860 4635 3864
rect 4641 3860 4645 3864
rect 4661 3860 4665 3864
rect 4785 3860 4789 3864
rect 4805 3860 4809 3864
rect 4891 3860 4895 3864
rect 4911 3860 4915 3864
rect 4931 3860 4935 3864
rect 5031 3860 5035 3864
rect 5145 3860 5149 3864
rect 5191 3860 5195 3864
rect 5213 3860 5217 3864
rect 5221 3860 5225 3864
rect 5241 3860 5245 3864
rect 5249 3860 5253 3864
rect 5295 3860 5299 3864
rect 5315 3860 5319 3864
rect 5327 3860 5331 3864
rect 5347 3860 5351 3864
rect 5361 3860 5365 3864
rect 5381 3860 5385 3864
rect 5431 3860 5435 3864
rect 5453 3860 5457 3864
rect 5461 3860 5465 3864
rect 5481 3860 5485 3864
rect 5489 3860 5493 3864
rect 5535 3860 5539 3864
rect 5555 3860 5559 3864
rect 5567 3860 5571 3864
rect 5587 3860 5591 3864
rect 5601 3860 5605 3864
rect 5621 3860 5625 3864
rect 5716 3860 5720 3864
rect 5724 3860 5728 3864
rect 5746 3860 5750 3864
rect 85 3836 89 3840
rect 105 3836 109 3840
rect 205 3836 209 3840
rect 225 3836 229 3840
rect 245 3836 249 3840
rect 405 3836 409 3840
rect 425 3836 429 3840
rect 445 3836 449 3840
rect 465 3836 469 3840
rect 570 3836 574 3840
rect 592 3836 596 3840
rect 600 3836 604 3840
rect 705 3836 709 3840
rect 725 3836 729 3840
rect 816 3836 820 3840
rect 824 3836 828 3840
rect 846 3836 850 3840
rect 985 3836 989 3840
rect 1005 3836 1009 3840
rect 1025 3836 1029 3840
rect 1045 3836 1049 3840
rect 1131 3836 1135 3840
rect 1151 3836 1155 3840
rect 1251 3836 1255 3840
rect 1271 3836 1275 3840
rect 1291 3836 1295 3840
rect 1391 3836 1395 3840
rect 1411 3836 1415 3840
rect 1431 3836 1435 3840
rect 1536 3836 1540 3840
rect 1544 3836 1548 3840
rect 1566 3836 1570 3840
rect 1671 3836 1675 3840
rect 1785 3836 1789 3840
rect 1805 3836 1809 3840
rect 1891 3836 1895 3840
rect 1911 3836 1915 3840
rect 2011 3836 2015 3840
rect 2021 3836 2025 3840
rect 2041 3836 2045 3840
rect 2151 3836 2155 3840
rect 2171 3836 2175 3840
rect 2271 3836 2275 3840
rect 2291 3836 2295 3840
rect 2311 3836 2315 3840
rect 2430 3836 2434 3840
rect 2452 3836 2456 3840
rect 2460 3836 2464 3840
rect 2551 3836 2555 3840
rect 2571 3836 2575 3840
rect 2676 3836 2680 3840
rect 2684 3836 2688 3840
rect 2706 3836 2710 3840
rect 2825 3836 2829 3840
rect 2930 3836 2934 3840
rect 2952 3836 2956 3840
rect 2960 3836 2964 3840
rect 3051 3836 3055 3840
rect 3071 3836 3075 3840
rect 3205 3836 3209 3840
rect 3225 3836 3229 3840
rect 3325 3836 3329 3840
rect 3411 3836 3415 3840
rect 3431 3836 3435 3840
rect 3451 3836 3455 3840
rect 3551 3836 3555 3840
rect 3677 3836 3681 3840
rect 3685 3836 3689 3840
rect 3791 3836 3795 3840
rect 3811 3836 3815 3840
rect 3911 3836 3915 3840
rect 4025 3836 4029 3840
rect 4071 3836 4075 3840
rect 4093 3836 4097 3840
rect 4101 3836 4105 3840
rect 4121 3836 4125 3840
rect 4129 3836 4133 3840
rect 4175 3836 4179 3840
rect 4195 3836 4199 3840
rect 4207 3836 4211 3840
rect 4227 3836 4231 3840
rect 4241 3836 4245 3840
rect 4261 3836 4265 3840
rect 4375 3836 4379 3840
rect 4385 3836 4389 3840
rect 4415 3836 4419 3840
rect 4425 3836 4429 3840
rect 4511 3836 4515 3840
rect 4531 3836 4535 3840
rect 4631 3836 4635 3840
rect 4639 3836 4643 3840
rect 4756 3836 4760 3840
rect 4764 3836 4768 3840
rect 4786 3836 4790 3840
rect 4891 3836 4895 3840
rect 5025 3836 5029 3840
rect 5045 3836 5049 3840
rect 5131 3836 5135 3840
rect 5245 3836 5249 3840
rect 5265 3836 5269 3840
rect 5285 3836 5289 3840
rect 5305 3836 5309 3840
rect 5325 3836 5329 3840
rect 5345 3836 5349 3840
rect 5365 3836 5369 3840
rect 5385 3836 5389 3840
rect 5431 3836 5435 3840
rect 5453 3836 5457 3840
rect 5461 3836 5465 3840
rect 5481 3836 5485 3840
rect 5489 3836 5493 3840
rect 5535 3836 5539 3840
rect 5555 3836 5559 3840
rect 5567 3836 5571 3840
rect 5587 3836 5591 3840
rect 5601 3836 5605 3840
rect 5621 3836 5625 3840
rect 5725 3836 5729 3840
rect 5745 3836 5749 3840
rect 341 3828 345 3832
rect 361 3828 365 3832
rect 85 3719 89 3796
rect 86 3707 89 3719
rect 83 3691 89 3707
rect 105 3719 109 3796
rect 205 3753 209 3796
rect 225 3784 229 3796
rect 245 3788 249 3796
rect 245 3784 260 3788
rect 225 3780 240 3784
rect 234 3773 240 3780
rect 205 3741 213 3753
rect 225 3741 232 3753
rect 105 3707 114 3719
rect 105 3691 111 3707
rect 83 3684 97 3691
rect 93 3664 97 3684
rect 103 3684 111 3691
rect 228 3684 232 3741
rect 236 3684 240 3761
rect 254 3753 260 3784
rect 405 3772 409 3776
rect 425 3772 429 3776
rect 405 3768 429 3772
rect 341 3760 345 3768
rect 361 3760 365 3768
rect 341 3756 391 3760
rect 244 3741 254 3753
rect 244 3684 248 3741
rect 385 3733 391 3756
rect 385 3721 394 3733
rect 103 3664 107 3684
rect 385 3666 391 3721
rect 425 3699 429 3768
rect 426 3687 429 3699
rect 385 3660 409 3666
rect 405 3644 409 3660
rect 425 3644 429 3687
rect 445 3772 449 3776
rect 465 3772 469 3776
rect 445 3768 469 3772
rect 445 3733 449 3768
rect 570 3753 574 3796
rect 567 3741 574 3753
rect 445 3721 454 3733
rect 445 3644 449 3721
rect 565 3664 569 3741
rect 592 3699 596 3756
rect 600 3752 604 3756
rect 600 3744 618 3752
rect 614 3733 618 3744
rect 585 3687 594 3699
rect 585 3664 589 3687
rect 614 3676 618 3721
rect 705 3719 709 3796
rect 706 3707 709 3719
rect 703 3691 709 3707
rect 725 3719 729 3796
rect 816 3752 820 3756
rect 802 3744 820 3752
rect 802 3733 806 3744
rect 725 3707 734 3719
rect 725 3691 731 3707
rect 703 3684 717 3691
rect 605 3669 618 3676
rect 605 3664 609 3669
rect 713 3664 717 3684
rect 723 3684 731 3691
rect 723 3664 727 3684
rect 802 3676 806 3721
rect 824 3699 828 3756
rect 846 3753 850 3796
rect 846 3741 853 3753
rect 826 3687 835 3699
rect 802 3669 815 3676
rect 811 3664 815 3669
rect 831 3664 835 3687
rect 851 3664 855 3741
rect 985 3733 989 3756
rect 986 3721 989 3733
rect 980 3673 986 3721
rect 1005 3699 1009 3756
rect 1025 3734 1029 3756
rect 1045 3734 1049 3756
rect 1025 3728 1038 3734
rect 1045 3733 1065 3734
rect 1045 3728 1053 3733
rect 1034 3699 1038 3728
rect 1007 3687 1009 3699
rect 1005 3685 1009 3687
rect 1005 3678 1018 3685
rect 980 3669 1010 3673
rect 1006 3664 1010 3669
rect 1014 3664 1018 3678
rect 1034 3664 1038 3687
rect 1053 3679 1059 3721
rect 1131 3719 1135 3796
rect 1126 3707 1135 3719
rect 1129 3691 1135 3707
rect 1151 3719 1155 3796
rect 1251 3788 1255 3796
rect 1240 3784 1255 3788
rect 1271 3784 1275 3796
rect 1240 3753 1246 3784
rect 1260 3780 1275 3784
rect 1260 3773 1266 3780
rect 1246 3741 1256 3753
rect 1151 3707 1154 3719
rect 1151 3691 1157 3707
rect 1129 3684 1137 3691
rect 1042 3672 1059 3679
rect 1042 3664 1046 3672
rect 1133 3664 1137 3684
rect 1143 3684 1157 3691
rect 1252 3684 1256 3741
rect 1260 3684 1264 3761
rect 1291 3753 1295 3796
rect 1268 3741 1275 3753
rect 1287 3741 1295 3753
rect 1391 3742 1395 3756
rect 1411 3742 1415 3756
rect 1268 3684 1272 3741
rect 1379 3736 1395 3742
rect 1400 3736 1415 3742
rect 1379 3699 1386 3736
rect 1400 3713 1406 3736
rect 1143 3664 1147 3684
rect 1379 3674 1386 3687
rect 1379 3668 1398 3674
rect 1394 3664 1398 3668
rect 1402 3664 1406 3701
rect 1431 3699 1435 3756
rect 1536 3752 1540 3756
rect 1522 3744 1540 3752
rect 1522 3733 1526 3744
rect 1426 3687 1435 3699
rect 1424 3644 1428 3687
rect 1522 3676 1526 3721
rect 1544 3699 1548 3756
rect 1566 3753 1570 3796
rect 1566 3741 1573 3753
rect 1546 3687 1555 3699
rect 1522 3669 1535 3676
rect 1531 3664 1535 3669
rect 1551 3664 1555 3687
rect 1571 3664 1575 3741
rect 1671 3713 1675 3796
rect 1785 3719 1789 3796
rect 1666 3701 1675 3713
rect 1786 3707 1789 3719
rect 1671 3644 1675 3701
rect 1783 3691 1789 3707
rect 1805 3719 1809 3796
rect 1891 3719 1895 3796
rect 1805 3707 1814 3719
rect 1886 3707 1895 3719
rect 1805 3691 1811 3707
rect 1783 3684 1797 3691
rect 1793 3664 1797 3684
rect 1803 3684 1811 3691
rect 1889 3691 1895 3707
rect 1911 3719 1915 3796
rect 2011 3752 2015 3756
rect 2002 3747 2015 3752
rect 1911 3707 1914 3719
rect 2002 3713 2006 3747
rect 2021 3733 2025 3756
rect 2041 3751 2045 3756
rect 1911 3691 1917 3707
rect 1889 3684 1897 3691
rect 1803 3664 1807 3684
rect 1893 3664 1897 3684
rect 1903 3684 1917 3691
rect 1903 3664 1907 3684
rect 2002 3656 2006 3701
rect 2021 3657 2025 3721
rect 2151 3719 2155 3796
rect 2146 3707 2155 3719
rect 2149 3691 2155 3707
rect 2171 3719 2175 3796
rect 2271 3788 2275 3796
rect 2260 3784 2275 3788
rect 2291 3784 2295 3796
rect 2260 3753 2266 3784
rect 2280 3780 2295 3784
rect 2280 3773 2286 3780
rect 2266 3741 2276 3753
rect 2171 3707 2174 3719
rect 2171 3691 2177 3707
rect 2149 3684 2157 3691
rect 2045 3672 2055 3684
rect 2051 3664 2055 3672
rect 2153 3664 2157 3684
rect 2163 3684 2177 3691
rect 2272 3684 2276 3741
rect 2280 3684 2284 3761
rect 2311 3753 2315 3796
rect 2430 3753 2434 3796
rect 2288 3741 2295 3753
rect 2307 3741 2315 3753
rect 2427 3741 2434 3753
rect 2288 3684 2292 3741
rect 2163 3664 2167 3684
rect 2002 3651 2015 3656
rect 2021 3651 2035 3657
rect 2011 3644 2015 3651
rect 2031 3644 2035 3651
rect 2425 3664 2429 3741
rect 2452 3699 2456 3756
rect 2460 3752 2464 3756
rect 2460 3744 2478 3752
rect 2474 3733 2478 3744
rect 2445 3687 2454 3699
rect 2445 3664 2449 3687
rect 2474 3676 2478 3721
rect 2551 3719 2555 3796
rect 2546 3707 2555 3719
rect 2549 3691 2555 3707
rect 2571 3719 2575 3796
rect 2676 3752 2680 3756
rect 2662 3744 2680 3752
rect 2662 3733 2666 3744
rect 2571 3707 2574 3719
rect 2571 3691 2577 3707
rect 2549 3684 2557 3691
rect 2465 3669 2478 3676
rect 2465 3664 2469 3669
rect 2553 3664 2557 3684
rect 2563 3684 2577 3691
rect 2563 3664 2567 3684
rect 2662 3676 2666 3721
rect 2684 3699 2688 3756
rect 2706 3753 2710 3796
rect 2706 3741 2713 3753
rect 2686 3687 2695 3699
rect 2662 3669 2675 3676
rect 2671 3664 2675 3669
rect 2691 3664 2695 3687
rect 2711 3664 2715 3741
rect 2825 3713 2829 3796
rect 2930 3753 2934 3796
rect 2927 3741 2934 3753
rect 2825 3701 2834 3713
rect 2825 3644 2829 3701
rect 2925 3664 2929 3741
rect 2952 3699 2956 3756
rect 2960 3752 2964 3756
rect 2960 3744 2978 3752
rect 2974 3733 2978 3744
rect 2945 3687 2954 3699
rect 2945 3664 2949 3687
rect 2974 3676 2978 3721
rect 3051 3719 3055 3796
rect 3046 3707 3055 3719
rect 3049 3691 3055 3707
rect 3071 3719 3075 3796
rect 3205 3719 3209 3796
rect 3071 3707 3074 3719
rect 3206 3707 3209 3719
rect 3071 3691 3077 3707
rect 3049 3684 3057 3691
rect 2965 3669 2978 3676
rect 2965 3664 2969 3669
rect 3053 3664 3057 3684
rect 3063 3684 3077 3691
rect 3203 3691 3209 3707
rect 3225 3719 3229 3796
rect 3225 3707 3234 3719
rect 3325 3713 3329 3796
rect 3411 3788 3415 3796
rect 3400 3784 3415 3788
rect 3431 3784 3435 3796
rect 3400 3753 3406 3784
rect 3420 3780 3435 3784
rect 3420 3773 3426 3780
rect 3406 3741 3416 3753
rect 3225 3691 3231 3707
rect 3203 3684 3217 3691
rect 3063 3664 3067 3684
rect 3213 3664 3217 3684
rect 3223 3684 3231 3691
rect 3325 3701 3334 3713
rect 3223 3664 3227 3684
rect 3325 3644 3329 3701
rect 3412 3684 3416 3741
rect 3420 3684 3424 3761
rect 3451 3753 3455 3796
rect 3428 3741 3435 3753
rect 3447 3741 3455 3753
rect 3428 3684 3432 3741
rect 3551 3713 3555 3796
rect 3677 3733 3681 3756
rect 3666 3721 3681 3733
rect 3685 3733 3689 3756
rect 3685 3721 3694 3733
rect 3546 3701 3555 3713
rect 3551 3644 3555 3701
rect 3665 3644 3669 3721
rect 3685 3644 3689 3721
rect 3791 3719 3795 3796
rect 3786 3707 3795 3719
rect 3789 3691 3795 3707
rect 3811 3719 3815 3796
rect 3811 3707 3814 3719
rect 3911 3713 3915 3796
rect 3811 3691 3817 3707
rect 3906 3701 3915 3713
rect 3789 3684 3797 3691
rect 3793 3664 3797 3684
rect 3803 3684 3817 3691
rect 3803 3664 3807 3684
rect 3911 3644 3915 3701
rect 4025 3713 4029 3796
rect 4093 3793 4097 3816
rect 4089 3786 4097 3793
rect 4089 3757 4093 3786
rect 4101 3776 4105 3816
rect 4121 3764 4125 3796
rect 4129 3792 4133 3796
rect 4129 3790 4165 3792
rect 4129 3788 4153 3790
rect 4071 3744 4075 3756
rect 4089 3751 4097 3757
rect 4071 3732 4073 3744
rect 4025 3701 4034 3713
rect 4025 3644 4029 3701
rect 4071 3664 4075 3732
rect 4093 3705 4097 3751
rect 4093 3644 4097 3693
rect 4121 3669 4127 3764
rect 4103 3665 4127 3669
rect 4103 3644 4107 3665
rect 4123 3660 4141 3661
rect 4123 3656 4153 3660
rect 4123 3644 4127 3656
rect 4161 3652 4165 3778
rect 4175 3770 4179 3796
rect 4195 3790 4199 3796
rect 4131 3648 4165 3652
rect 4131 3644 4135 3648
rect 4177 3644 4181 3758
rect 4193 3668 4197 3778
rect 4207 3756 4211 3796
rect 4202 3744 4205 3756
rect 4202 3680 4206 3744
rect 4227 3737 4231 3796
rect 4222 3729 4231 3737
rect 4222 3700 4226 3729
rect 4241 3714 4245 3796
rect 4261 3713 4265 3756
rect 4375 3752 4379 3756
rect 4365 3748 4379 3752
rect 4365 3733 4369 3748
rect 4367 3721 4369 3733
rect 4202 3676 4235 3680
rect 4201 3656 4203 3668
rect 4199 3644 4203 3656
rect 4209 3656 4211 3668
rect 4209 3644 4213 3656
rect 4231 3644 4235 3676
rect 4241 3644 4245 3702
rect 4261 3664 4265 3701
rect 4365 3664 4369 3721
rect 4385 3699 4389 3756
rect 4415 3752 4419 3756
rect 4405 3748 4419 3752
rect 4425 3752 4429 3756
rect 4425 3748 4439 3752
rect 4405 3699 4411 3748
rect 4434 3733 4439 3748
rect 4405 3687 4414 3699
rect 4385 3664 4389 3687
rect 4405 3664 4409 3687
rect 4434 3675 4440 3721
rect 4511 3719 4515 3796
rect 4506 3707 4515 3719
rect 4509 3691 4515 3707
rect 4531 3719 4535 3796
rect 4631 3733 4635 3756
rect 4626 3721 4635 3733
rect 4639 3733 4643 3756
rect 4756 3752 4760 3756
rect 4742 3744 4760 3752
rect 4742 3733 4746 3744
rect 4639 3721 4654 3733
rect 4531 3707 4534 3719
rect 4531 3691 4537 3707
rect 4509 3684 4517 3691
rect 4425 3671 4440 3675
rect 4425 3664 4429 3671
rect 4513 3664 4517 3684
rect 4523 3684 4537 3691
rect 4523 3664 4527 3684
rect 4631 3644 4635 3721
rect 4651 3644 4655 3721
rect 4742 3676 4746 3721
rect 4764 3699 4768 3756
rect 4786 3753 4790 3796
rect 4786 3741 4793 3753
rect 4766 3687 4775 3699
rect 4742 3669 4755 3676
rect 4751 3664 4755 3669
rect 4771 3664 4775 3687
rect 4791 3664 4795 3741
rect 4891 3699 4895 3756
rect 5025 3719 5029 3796
rect 5026 3707 5029 3719
rect 4886 3687 4895 3699
rect 4891 3664 4895 3687
rect 5023 3691 5029 3707
rect 5045 3719 5049 3796
rect 5045 3707 5054 3719
rect 5131 3713 5135 3796
rect 5453 3793 5457 3816
rect 5449 3786 5457 3793
rect 5449 3757 5453 3786
rect 5461 3776 5465 3816
rect 5481 3764 5485 3796
rect 5489 3792 5493 3796
rect 5489 3790 5525 3792
rect 5489 3788 5513 3790
rect 5045 3691 5051 3707
rect 5126 3701 5135 3713
rect 5023 3684 5037 3691
rect 5033 3664 5037 3684
rect 5043 3684 5051 3691
rect 5043 3664 5047 3684
rect 5131 3644 5135 3701
rect 5245 3696 5249 3756
rect 5265 3696 5269 3756
rect 5285 3696 5289 3756
rect 5305 3696 5309 3756
rect 5325 3696 5329 3756
rect 5345 3696 5349 3756
rect 5365 3699 5369 3756
rect 5385 3699 5389 3756
rect 5245 3684 5258 3696
rect 5285 3684 5298 3696
rect 5325 3684 5338 3696
rect 5365 3687 5374 3699
rect 5386 3687 5389 3699
rect 5245 3664 5249 3684
rect 5265 3664 5269 3684
rect 5285 3664 5289 3684
rect 5305 3664 5309 3684
rect 5325 3664 5329 3684
rect 5345 3664 5349 3684
rect 5365 3664 5369 3687
rect 5385 3664 5389 3687
rect 5431 3744 5435 3756
rect 5449 3751 5457 3757
rect 5431 3732 5433 3744
rect 5431 3664 5435 3732
rect 5453 3705 5457 3751
rect 5453 3644 5457 3693
rect 5481 3669 5487 3764
rect 5463 3665 5487 3669
rect 5463 3644 5467 3665
rect 5483 3660 5501 3661
rect 5483 3656 5513 3660
rect 5483 3644 5487 3656
rect 5521 3652 5525 3778
rect 5535 3770 5539 3796
rect 5555 3790 5559 3796
rect 5491 3648 5525 3652
rect 5491 3644 5495 3648
rect 5537 3644 5541 3758
rect 5553 3668 5557 3778
rect 5567 3756 5571 3796
rect 5562 3744 5565 3756
rect 5562 3680 5566 3744
rect 5587 3737 5591 3796
rect 5582 3729 5591 3737
rect 5582 3700 5586 3729
rect 5601 3714 5605 3796
rect 5621 3713 5625 3756
rect 5725 3719 5729 3796
rect 5562 3676 5595 3680
rect 5561 3656 5563 3668
rect 5559 3644 5563 3656
rect 5569 3656 5571 3668
rect 5569 3644 5573 3656
rect 5591 3644 5595 3676
rect 5601 3644 5605 3702
rect 5726 3707 5729 3719
rect 5621 3664 5625 3701
rect 5723 3691 5729 3707
rect 5745 3719 5749 3796
rect 5745 3707 5754 3719
rect 5745 3691 5751 3707
rect 5723 3684 5737 3691
rect 5733 3664 5737 3684
rect 5743 3684 5751 3691
rect 5743 3664 5747 3684
rect 93 3620 97 3624
rect 103 3620 107 3624
rect 228 3620 232 3624
rect 236 3620 240 3624
rect 244 3620 248 3624
rect 405 3620 409 3624
rect 425 3620 429 3624
rect 445 3620 449 3624
rect 565 3620 569 3624
rect 585 3620 589 3624
rect 605 3620 609 3624
rect 713 3620 717 3624
rect 723 3620 727 3624
rect 811 3620 815 3624
rect 831 3620 835 3624
rect 851 3620 855 3624
rect 1006 3620 1010 3624
rect 1014 3620 1018 3624
rect 1034 3620 1038 3624
rect 1042 3620 1046 3624
rect 1133 3620 1137 3624
rect 1143 3620 1147 3624
rect 1252 3620 1256 3624
rect 1260 3620 1264 3624
rect 1268 3620 1272 3624
rect 1394 3620 1398 3624
rect 1402 3620 1406 3624
rect 1424 3620 1428 3624
rect 1531 3620 1535 3624
rect 1551 3620 1555 3624
rect 1571 3620 1575 3624
rect 1671 3620 1675 3624
rect 1793 3620 1797 3624
rect 1803 3620 1807 3624
rect 1893 3620 1897 3624
rect 1903 3620 1907 3624
rect 2011 3620 2015 3624
rect 2031 3620 2035 3624
rect 2051 3620 2055 3624
rect 2153 3620 2157 3624
rect 2163 3620 2167 3624
rect 2272 3620 2276 3624
rect 2280 3620 2284 3624
rect 2288 3620 2292 3624
rect 2425 3620 2429 3624
rect 2445 3620 2449 3624
rect 2465 3620 2469 3624
rect 2553 3620 2557 3624
rect 2563 3620 2567 3624
rect 2671 3620 2675 3624
rect 2691 3620 2695 3624
rect 2711 3620 2715 3624
rect 2825 3620 2829 3624
rect 2925 3620 2929 3624
rect 2945 3620 2949 3624
rect 2965 3620 2969 3624
rect 3053 3620 3057 3624
rect 3063 3620 3067 3624
rect 3213 3620 3217 3624
rect 3223 3620 3227 3624
rect 3325 3620 3329 3624
rect 3412 3620 3416 3624
rect 3420 3620 3424 3624
rect 3428 3620 3432 3624
rect 3551 3620 3555 3624
rect 3665 3620 3669 3624
rect 3685 3620 3689 3624
rect 3793 3620 3797 3624
rect 3803 3620 3807 3624
rect 3911 3620 3915 3624
rect 4025 3620 4029 3624
rect 4071 3620 4075 3624
rect 4093 3620 4097 3624
rect 4103 3620 4107 3624
rect 4123 3620 4127 3624
rect 4131 3620 4135 3624
rect 4177 3620 4181 3624
rect 4199 3620 4203 3624
rect 4209 3620 4213 3624
rect 4231 3620 4235 3624
rect 4241 3620 4245 3624
rect 4261 3620 4265 3624
rect 4365 3620 4369 3624
rect 4385 3620 4389 3624
rect 4405 3620 4409 3624
rect 4425 3620 4429 3624
rect 4513 3620 4517 3624
rect 4523 3620 4527 3624
rect 4631 3620 4635 3624
rect 4651 3620 4655 3624
rect 4751 3620 4755 3624
rect 4771 3620 4775 3624
rect 4791 3620 4795 3624
rect 4891 3620 4895 3624
rect 5033 3620 5037 3624
rect 5043 3620 5047 3624
rect 5131 3620 5135 3624
rect 5245 3620 5249 3624
rect 5265 3620 5269 3624
rect 5285 3620 5289 3624
rect 5305 3620 5309 3624
rect 5325 3620 5329 3624
rect 5345 3620 5349 3624
rect 5365 3620 5369 3624
rect 5385 3620 5389 3624
rect 5431 3620 5435 3624
rect 5453 3620 5457 3624
rect 5463 3620 5467 3624
rect 5483 3620 5487 3624
rect 5491 3620 5495 3624
rect 5537 3620 5541 3624
rect 5559 3620 5563 3624
rect 5569 3620 5573 3624
rect 5591 3620 5595 3624
rect 5601 3620 5605 3624
rect 5621 3620 5625 3624
rect 5733 3620 5737 3624
rect 5743 3620 5747 3624
rect 85 3596 89 3600
rect 105 3596 109 3600
rect 125 3596 129 3600
rect 214 3596 218 3600
rect 222 3596 226 3600
rect 244 3596 248 3600
rect 351 3596 355 3600
rect 451 3596 455 3600
rect 471 3596 475 3600
rect 491 3596 495 3600
rect 592 3596 596 3600
rect 600 3596 604 3600
rect 608 3596 612 3600
rect 773 3596 777 3600
rect 783 3596 787 3600
rect 893 3596 897 3600
rect 903 3596 907 3600
rect 991 3596 995 3600
rect 1011 3596 1015 3600
rect 1031 3596 1035 3600
rect 1168 3596 1172 3600
rect 1176 3596 1180 3600
rect 1184 3596 1188 3600
rect 1273 3596 1277 3600
rect 1283 3596 1287 3600
rect 1428 3596 1432 3600
rect 1436 3596 1440 3600
rect 1444 3596 1448 3600
rect 1531 3596 1535 3600
rect 1551 3596 1555 3600
rect 1571 3596 1575 3600
rect 1692 3596 1696 3600
rect 1714 3596 1718 3600
rect 1722 3596 1726 3600
rect 1848 3596 1852 3600
rect 1856 3596 1860 3600
rect 1864 3596 1868 3600
rect 1954 3596 1958 3600
rect 1962 3596 1966 3600
rect 1984 3596 1988 3600
rect 2105 3596 2109 3600
rect 2125 3596 2129 3600
rect 2145 3596 2149 3600
rect 2251 3596 2255 3600
rect 2271 3596 2275 3600
rect 2291 3596 2295 3600
rect 2412 3596 2416 3600
rect 2434 3596 2438 3600
rect 2442 3596 2446 3600
rect 2555 3596 2559 3600
rect 2575 3596 2579 3600
rect 2585 3596 2589 3600
rect 2673 3596 2677 3600
rect 2683 3596 2687 3600
rect 2805 3596 2809 3600
rect 2825 3596 2829 3600
rect 2845 3596 2849 3600
rect 2963 3596 2967 3600
rect 2985 3596 2989 3600
rect 3093 3596 3097 3600
rect 3103 3596 3107 3600
rect 3192 3596 3196 3600
rect 3200 3596 3204 3600
rect 3208 3596 3212 3600
rect 3368 3596 3372 3600
rect 3376 3596 3380 3600
rect 3384 3596 3388 3600
rect 3485 3596 3489 3600
rect 3505 3596 3509 3600
rect 3525 3596 3529 3600
rect 3625 3596 3629 3600
rect 3645 3596 3649 3600
rect 3665 3596 3669 3600
rect 3775 3596 3779 3600
rect 3795 3596 3799 3600
rect 3805 3596 3809 3600
rect 3891 3596 3895 3600
rect 3911 3596 3915 3600
rect 4045 3596 4049 3600
rect 4065 3596 4069 3600
rect 4085 3596 4089 3600
rect 4171 3596 4175 3600
rect 4271 3596 4275 3600
rect 4291 3596 4295 3600
rect 4311 3596 4315 3600
rect 4433 3596 4437 3600
rect 4443 3596 4447 3600
rect 4533 3596 4537 3600
rect 4543 3596 4547 3600
rect 4611 3596 4615 3600
rect 4633 3596 4637 3600
rect 4643 3596 4647 3600
rect 4663 3596 4667 3600
rect 4671 3596 4675 3600
rect 4717 3596 4721 3600
rect 4739 3596 4743 3600
rect 4749 3596 4753 3600
rect 4771 3596 4775 3600
rect 4781 3596 4785 3600
rect 4801 3596 4805 3600
rect 4913 3596 4917 3600
rect 4923 3596 4927 3600
rect 5025 3596 5029 3600
rect 5045 3596 5049 3600
rect 5065 3596 5069 3600
rect 5173 3596 5177 3600
rect 5183 3596 5187 3600
rect 5255 3596 5259 3600
rect 5275 3596 5279 3600
rect 5285 3596 5289 3600
rect 5307 3596 5311 3600
rect 5317 3596 5321 3600
rect 5339 3596 5343 3600
rect 5385 3596 5389 3600
rect 5393 3596 5397 3600
rect 5413 3596 5417 3600
rect 5423 3596 5427 3600
rect 5445 3596 5449 3600
rect 5553 3596 5557 3600
rect 5563 3596 5567 3600
rect 5651 3596 5655 3600
rect 5671 3596 5675 3600
rect 5691 3596 5695 3600
rect 85 3479 89 3556
rect 105 3533 109 3556
rect 125 3551 129 3556
rect 214 3552 218 3556
rect 125 3544 138 3551
rect 105 3521 114 3533
rect 87 3467 94 3479
rect 90 3424 94 3467
rect 112 3464 116 3521
rect 134 3499 138 3544
rect 199 3546 218 3552
rect 199 3533 206 3546
rect 134 3476 138 3487
rect 199 3484 206 3521
rect 222 3519 226 3556
rect 244 3533 248 3576
rect 246 3521 255 3533
rect 220 3484 226 3507
rect 199 3478 215 3484
rect 220 3478 235 3484
rect 120 3468 138 3476
rect 120 3464 124 3468
rect 211 3464 215 3478
rect 231 3464 235 3478
rect 251 3464 255 3521
rect 351 3519 355 3576
rect 451 3551 455 3556
rect 346 3507 355 3519
rect 351 3424 355 3507
rect 442 3544 455 3551
rect 442 3499 446 3544
rect 471 3533 475 3556
rect 466 3521 475 3533
rect 442 3476 446 3487
rect 442 3468 460 3476
rect 456 3464 460 3468
rect 464 3464 468 3521
rect 491 3479 495 3556
rect 773 3536 777 3556
rect 592 3479 596 3536
rect 486 3467 493 3479
rect 586 3467 596 3479
rect 486 3424 490 3467
rect 580 3436 586 3467
rect 600 3459 604 3536
rect 608 3479 612 3536
rect 763 3529 777 3536
rect 783 3536 787 3556
rect 893 3536 897 3556
rect 783 3529 791 3536
rect 763 3513 769 3529
rect 766 3501 769 3513
rect 608 3467 615 3479
rect 627 3467 635 3479
rect 600 3440 606 3447
rect 600 3436 615 3440
rect 580 3432 595 3436
rect 591 3424 595 3432
rect 611 3424 615 3436
rect 631 3424 635 3467
rect 765 3424 769 3501
rect 785 3513 791 3529
rect 883 3529 897 3536
rect 903 3536 907 3556
rect 991 3551 995 3556
rect 982 3544 995 3551
rect 903 3529 911 3536
rect 883 3513 889 3529
rect 785 3501 794 3513
rect 886 3501 889 3513
rect 785 3424 789 3501
rect 885 3424 889 3501
rect 905 3513 911 3529
rect 905 3501 914 3513
rect 905 3424 909 3501
rect 982 3499 986 3544
rect 1011 3533 1015 3556
rect 1006 3521 1015 3533
rect 982 3476 986 3487
rect 982 3468 1000 3476
rect 996 3464 1000 3468
rect 1004 3464 1008 3521
rect 1031 3479 1035 3556
rect 1273 3536 1277 3556
rect 1168 3479 1172 3536
rect 1026 3467 1033 3479
rect 1145 3467 1153 3479
rect 1165 3467 1172 3479
rect 1026 3424 1030 3467
rect 1145 3424 1149 3467
rect 1176 3459 1180 3536
rect 1184 3479 1188 3536
rect 1269 3529 1277 3536
rect 1283 3536 1287 3556
rect 1531 3551 1535 3556
rect 1522 3544 1535 3551
rect 1283 3529 1297 3536
rect 1269 3513 1275 3529
rect 1266 3501 1275 3513
rect 1184 3467 1194 3479
rect 1174 3440 1180 3447
rect 1165 3436 1180 3440
rect 1194 3436 1200 3467
rect 1165 3424 1169 3436
rect 1185 3432 1200 3436
rect 1185 3424 1189 3432
rect 1271 3424 1275 3501
rect 1291 3513 1297 3529
rect 1291 3501 1294 3513
rect 1291 3424 1295 3501
rect 1428 3479 1432 3536
rect 1405 3467 1413 3479
rect 1425 3467 1432 3479
rect 1405 3424 1409 3467
rect 1436 3459 1440 3536
rect 1444 3479 1448 3536
rect 1522 3499 1526 3544
rect 1551 3533 1555 3556
rect 1546 3521 1555 3533
rect 1444 3467 1454 3479
rect 1522 3476 1526 3487
rect 1522 3468 1540 3476
rect 1434 3440 1440 3447
rect 1425 3436 1440 3440
rect 1454 3436 1460 3467
rect 1536 3464 1540 3468
rect 1544 3464 1548 3521
rect 1571 3479 1575 3556
rect 1692 3533 1696 3576
rect 1685 3521 1694 3533
rect 1566 3467 1573 3479
rect 1425 3424 1429 3436
rect 1445 3432 1460 3436
rect 1445 3424 1449 3432
rect 1566 3424 1570 3467
rect 1685 3464 1689 3521
rect 1714 3519 1718 3556
rect 1722 3552 1726 3556
rect 1722 3546 1741 3552
rect 1734 3533 1741 3546
rect 1954 3552 1958 3556
rect 1939 3546 1958 3552
rect 1714 3484 1720 3507
rect 1734 3484 1741 3521
rect 1705 3478 1720 3484
rect 1725 3478 1741 3484
rect 1848 3479 1852 3536
rect 1705 3464 1709 3478
rect 1725 3464 1729 3478
rect 1825 3467 1833 3479
rect 1845 3467 1852 3479
rect 1825 3424 1829 3467
rect 1856 3459 1860 3536
rect 1864 3479 1868 3536
rect 1939 3533 1946 3546
rect 1939 3484 1946 3521
rect 1962 3519 1966 3556
rect 1984 3533 1988 3576
rect 1986 3521 1995 3533
rect 1960 3484 1966 3507
rect 1864 3467 1874 3479
rect 1939 3478 1955 3484
rect 1960 3478 1975 3484
rect 1854 3440 1860 3447
rect 1845 3436 1860 3440
rect 1874 3436 1880 3467
rect 1951 3464 1955 3478
rect 1971 3464 1975 3478
rect 1991 3464 1995 3521
rect 2105 3479 2109 3556
rect 2125 3533 2129 3556
rect 2145 3551 2149 3556
rect 2251 3551 2255 3556
rect 2145 3544 2158 3551
rect 2125 3521 2134 3533
rect 2107 3467 2114 3479
rect 1845 3424 1849 3436
rect 1865 3432 1880 3436
rect 1865 3424 1869 3432
rect 2110 3424 2114 3467
rect 2132 3464 2136 3521
rect 2154 3499 2158 3544
rect 2242 3544 2255 3551
rect 2242 3499 2246 3544
rect 2271 3533 2275 3556
rect 2266 3521 2275 3533
rect 2154 3476 2158 3487
rect 2140 3468 2158 3476
rect 2242 3476 2246 3487
rect 2242 3468 2260 3476
rect 2140 3464 2144 3468
rect 2256 3464 2260 3468
rect 2264 3464 2268 3521
rect 2291 3479 2295 3556
rect 2412 3533 2416 3576
rect 2405 3521 2414 3533
rect 2286 3467 2293 3479
rect 2286 3424 2290 3467
rect 2405 3464 2409 3521
rect 2434 3519 2438 3556
rect 2442 3552 2446 3556
rect 2442 3546 2461 3552
rect 2555 3550 2559 3556
rect 2454 3533 2461 3546
rect 2541 3538 2553 3550
rect 2434 3484 2440 3507
rect 2454 3484 2461 3521
rect 2425 3478 2440 3484
rect 2445 3478 2461 3484
rect 2425 3464 2429 3478
rect 2445 3464 2449 3478
rect 2541 3464 2545 3538
rect 2575 3513 2579 3556
rect 2566 3501 2579 3513
rect 2563 3424 2567 3501
rect 2585 3499 2589 3556
rect 2673 3536 2677 3556
rect 2669 3529 2677 3536
rect 2683 3536 2687 3556
rect 2683 3529 2697 3536
rect 2669 3513 2675 3529
rect 2666 3501 2675 3513
rect 2585 3487 2594 3499
rect 2585 3424 2589 3487
rect 2671 3424 2675 3501
rect 2691 3513 2697 3529
rect 2691 3501 2694 3513
rect 2691 3424 2695 3501
rect 2805 3479 2809 3556
rect 2825 3533 2829 3556
rect 2845 3551 2849 3556
rect 2845 3544 2858 3551
rect 2825 3521 2834 3533
rect 2807 3467 2814 3479
rect 2810 3424 2814 3467
rect 2832 3464 2836 3521
rect 2854 3499 2858 3544
rect 2963 3550 2967 3556
rect 2963 3538 2965 3550
rect 2985 3499 2989 3576
rect 3093 3536 3097 3556
rect 3083 3529 3097 3536
rect 3103 3536 3107 3556
rect 3103 3529 3111 3536
rect 3083 3513 3089 3529
rect 3086 3501 3089 3513
rect 2985 3487 2994 3499
rect 2854 3476 2858 3487
rect 2840 3468 2858 3476
rect 2963 3470 2965 3482
rect 2840 3464 2844 3468
rect 2963 3464 2967 3470
rect 2985 3424 2989 3487
rect 3085 3424 3089 3501
rect 3105 3513 3111 3529
rect 3105 3501 3114 3513
rect 3105 3424 3109 3501
rect 3192 3479 3196 3536
rect 3186 3467 3196 3479
rect 3180 3436 3186 3467
rect 3200 3459 3204 3536
rect 3208 3479 3212 3536
rect 3368 3479 3372 3536
rect 3208 3467 3215 3479
rect 3227 3467 3235 3479
rect 3200 3440 3206 3447
rect 3200 3436 3215 3440
rect 3180 3432 3195 3436
rect 3191 3424 3195 3432
rect 3211 3424 3215 3436
rect 3231 3424 3235 3467
rect 3345 3467 3353 3479
rect 3365 3467 3372 3479
rect 3345 3424 3349 3467
rect 3376 3459 3380 3536
rect 3384 3479 3388 3536
rect 3485 3479 3489 3556
rect 3505 3533 3509 3556
rect 3525 3551 3529 3556
rect 3525 3544 3538 3551
rect 3505 3521 3514 3533
rect 3384 3467 3394 3479
rect 3487 3467 3494 3479
rect 3374 3440 3380 3447
rect 3365 3436 3380 3440
rect 3394 3436 3400 3467
rect 3365 3424 3369 3436
rect 3385 3432 3400 3436
rect 3385 3424 3389 3432
rect 3490 3424 3494 3467
rect 3512 3464 3516 3521
rect 3534 3499 3538 3544
rect 3534 3476 3538 3487
rect 3625 3479 3629 3556
rect 3645 3533 3649 3556
rect 3665 3551 3669 3556
rect 3665 3544 3678 3551
rect 3775 3550 3779 3556
rect 3645 3521 3654 3533
rect 3520 3468 3538 3476
rect 3520 3464 3524 3468
rect 3627 3467 3634 3479
rect 3630 3424 3634 3467
rect 3652 3464 3656 3521
rect 3674 3499 3678 3544
rect 3761 3538 3773 3550
rect 3674 3476 3678 3487
rect 3660 3468 3678 3476
rect 3660 3464 3664 3468
rect 3761 3464 3765 3538
rect 3795 3513 3799 3556
rect 3786 3501 3799 3513
rect 3783 3424 3787 3501
rect 3805 3499 3809 3556
rect 3891 3499 3895 3576
rect 3911 3499 3915 3576
rect 3805 3487 3814 3499
rect 3886 3487 3895 3499
rect 3805 3424 3809 3487
rect 3891 3464 3895 3487
rect 3899 3487 3914 3499
rect 3899 3464 3903 3487
rect 4045 3479 4049 3556
rect 4065 3533 4069 3556
rect 4085 3551 4089 3556
rect 4085 3544 4098 3551
rect 4065 3521 4074 3533
rect 4047 3467 4054 3479
rect 4050 3424 4054 3467
rect 4072 3464 4076 3521
rect 4094 3499 4098 3544
rect 4171 3519 4175 3576
rect 4271 3551 4275 3556
rect 4166 3507 4175 3519
rect 4094 3476 4098 3487
rect 4080 3468 4098 3476
rect 4080 3464 4084 3468
rect 4171 3424 4175 3507
rect 4262 3544 4275 3551
rect 4262 3499 4266 3544
rect 4291 3533 4295 3556
rect 4286 3521 4295 3533
rect 4262 3476 4266 3487
rect 4262 3468 4280 3476
rect 4276 3464 4280 3468
rect 4284 3464 4288 3521
rect 4311 3479 4315 3556
rect 4433 3536 4437 3556
rect 4423 3529 4437 3536
rect 4443 3536 4447 3556
rect 4533 3536 4537 3556
rect 4443 3529 4451 3536
rect 4423 3513 4429 3529
rect 4426 3501 4429 3513
rect 4306 3467 4313 3479
rect 4306 3424 4310 3467
rect 4425 3424 4429 3501
rect 4445 3513 4451 3529
rect 4529 3529 4537 3536
rect 4543 3536 4547 3556
rect 4543 3529 4557 3536
rect 4529 3513 4535 3529
rect 4445 3501 4454 3513
rect 4526 3501 4535 3513
rect 4445 3424 4449 3501
rect 4531 3424 4535 3501
rect 4551 3513 4557 3529
rect 4551 3501 4554 3513
rect 4551 3424 4555 3501
rect 4611 3488 4615 3556
rect 4633 3527 4637 3576
rect 4643 3555 4647 3576
rect 4663 3564 4667 3576
rect 4671 3572 4675 3576
rect 4671 3568 4705 3572
rect 4663 3560 4693 3564
rect 4663 3559 4681 3560
rect 4643 3551 4667 3555
rect 4611 3476 4613 3488
rect 4611 3464 4615 3476
rect 4633 3469 4637 3515
rect 4629 3463 4637 3469
rect 4629 3434 4633 3463
rect 4661 3456 4667 3551
rect 4629 3427 4637 3434
rect 4633 3404 4637 3427
rect 4641 3404 4645 3444
rect 4661 3424 4665 3456
rect 4701 3442 4705 3568
rect 4717 3462 4721 3576
rect 4739 3564 4743 3576
rect 4741 3552 4743 3564
rect 4749 3564 4753 3576
rect 4749 3552 4751 3564
rect 4669 3430 4693 3432
rect 4669 3428 4705 3430
rect 4669 3424 4673 3428
rect 4715 3424 4719 3450
rect 4733 3442 4737 3552
rect 4771 3544 4775 3576
rect 4742 3540 4775 3544
rect 4742 3476 4746 3540
rect 4762 3491 4766 3520
rect 4781 3518 4785 3576
rect 4801 3519 4805 3556
rect 4913 3536 4917 3556
rect 4903 3529 4917 3536
rect 4923 3536 4927 3556
rect 4923 3529 4931 3536
rect 4903 3513 4909 3529
rect 4762 3483 4771 3491
rect 4742 3464 4745 3476
rect 4735 3424 4739 3430
rect 4747 3424 4751 3464
rect 4767 3424 4771 3483
rect 4781 3424 4785 3506
rect 4801 3464 4805 3507
rect 4906 3501 4909 3513
rect 4905 3424 4909 3501
rect 4925 3513 4931 3529
rect 4925 3501 4934 3513
rect 4925 3424 4929 3501
rect 5025 3479 5029 3556
rect 5045 3533 5049 3556
rect 5065 3551 5069 3556
rect 5065 3544 5078 3551
rect 5045 3521 5054 3533
rect 5027 3467 5034 3479
rect 5030 3424 5034 3467
rect 5052 3464 5056 3521
rect 5074 3499 5078 3544
rect 5173 3536 5177 3556
rect 5169 3529 5177 3536
rect 5183 3536 5187 3556
rect 5183 3529 5197 3536
rect 5169 3513 5175 3529
rect 5166 3501 5175 3513
rect 5074 3476 5078 3487
rect 5060 3468 5078 3476
rect 5060 3464 5064 3468
rect 5171 3424 5175 3501
rect 5191 3513 5197 3529
rect 5255 3519 5259 3556
rect 5191 3501 5194 3513
rect 5275 3518 5279 3576
rect 5285 3544 5289 3576
rect 5307 3564 5311 3576
rect 5309 3552 5311 3564
rect 5317 3564 5321 3576
rect 5317 3552 5319 3564
rect 5285 3540 5318 3544
rect 5191 3424 5195 3501
rect 5255 3464 5259 3507
rect 5275 3424 5279 3506
rect 5294 3491 5298 3520
rect 5289 3483 5298 3491
rect 5289 3424 5293 3483
rect 5314 3476 5318 3540
rect 5315 3464 5318 3476
rect 5309 3424 5313 3464
rect 5323 3442 5327 3552
rect 5339 3462 5343 3576
rect 5385 3572 5389 3576
rect 5355 3568 5389 3572
rect 5321 3424 5325 3430
rect 5341 3424 5345 3450
rect 5355 3442 5359 3568
rect 5393 3564 5397 3576
rect 5367 3560 5397 3564
rect 5379 3559 5397 3560
rect 5413 3555 5417 3576
rect 5393 3551 5417 3555
rect 5393 3456 5399 3551
rect 5423 3527 5427 3576
rect 5423 3469 5427 3515
rect 5445 3488 5449 3556
rect 5553 3536 5557 3556
rect 5543 3529 5557 3536
rect 5563 3536 5567 3556
rect 5651 3551 5655 3556
rect 5642 3544 5655 3551
rect 5563 3529 5571 3536
rect 5543 3513 5549 3529
rect 5546 3501 5549 3513
rect 5447 3476 5449 3488
rect 5423 3463 5431 3469
rect 5445 3464 5449 3476
rect 5367 3430 5391 3432
rect 5355 3428 5391 3430
rect 5387 3424 5391 3428
rect 5395 3424 5399 3456
rect 5415 3404 5419 3444
rect 5427 3434 5431 3463
rect 5423 3427 5431 3434
rect 5423 3404 5427 3427
rect 5545 3424 5549 3501
rect 5565 3513 5571 3529
rect 5565 3501 5574 3513
rect 5565 3424 5569 3501
rect 5642 3499 5646 3544
rect 5671 3533 5675 3556
rect 5666 3521 5675 3533
rect 5642 3476 5646 3487
rect 5642 3468 5660 3476
rect 5656 3464 5660 3468
rect 5664 3464 5668 3521
rect 5691 3479 5695 3556
rect 5686 3467 5693 3479
rect 5686 3424 5690 3467
rect 90 3380 94 3384
rect 112 3380 116 3384
rect 120 3380 124 3384
rect 211 3380 215 3384
rect 231 3380 235 3384
rect 251 3380 255 3384
rect 351 3380 355 3384
rect 456 3380 460 3384
rect 464 3380 468 3384
rect 486 3380 490 3384
rect 591 3380 595 3384
rect 611 3380 615 3384
rect 631 3380 635 3384
rect 765 3380 769 3384
rect 785 3380 789 3384
rect 885 3380 889 3384
rect 905 3380 909 3384
rect 996 3380 1000 3384
rect 1004 3380 1008 3384
rect 1026 3380 1030 3384
rect 1145 3380 1149 3384
rect 1165 3380 1169 3384
rect 1185 3380 1189 3384
rect 1271 3380 1275 3384
rect 1291 3380 1295 3384
rect 1405 3380 1409 3384
rect 1425 3380 1429 3384
rect 1445 3380 1449 3384
rect 1536 3380 1540 3384
rect 1544 3380 1548 3384
rect 1566 3380 1570 3384
rect 1685 3380 1689 3384
rect 1705 3380 1709 3384
rect 1725 3380 1729 3384
rect 1825 3380 1829 3384
rect 1845 3380 1849 3384
rect 1865 3380 1869 3384
rect 1951 3380 1955 3384
rect 1971 3380 1975 3384
rect 1991 3380 1995 3384
rect 2110 3380 2114 3384
rect 2132 3380 2136 3384
rect 2140 3380 2144 3384
rect 2256 3380 2260 3384
rect 2264 3380 2268 3384
rect 2286 3380 2290 3384
rect 2405 3380 2409 3384
rect 2425 3380 2429 3384
rect 2445 3380 2449 3384
rect 2541 3380 2545 3384
rect 2563 3380 2567 3384
rect 2585 3380 2589 3384
rect 2671 3380 2675 3384
rect 2691 3380 2695 3384
rect 2810 3380 2814 3384
rect 2832 3380 2836 3384
rect 2840 3380 2844 3384
rect 2963 3380 2967 3384
rect 2985 3380 2989 3384
rect 3085 3380 3089 3384
rect 3105 3380 3109 3384
rect 3191 3380 3195 3384
rect 3211 3380 3215 3384
rect 3231 3380 3235 3384
rect 3345 3380 3349 3384
rect 3365 3380 3369 3384
rect 3385 3380 3389 3384
rect 3490 3380 3494 3384
rect 3512 3380 3516 3384
rect 3520 3380 3524 3384
rect 3630 3380 3634 3384
rect 3652 3380 3656 3384
rect 3660 3380 3664 3384
rect 3761 3380 3765 3384
rect 3783 3380 3787 3384
rect 3805 3380 3809 3384
rect 3891 3380 3895 3384
rect 3899 3380 3903 3384
rect 4050 3380 4054 3384
rect 4072 3380 4076 3384
rect 4080 3380 4084 3384
rect 4171 3380 4175 3384
rect 4276 3380 4280 3384
rect 4284 3380 4288 3384
rect 4306 3380 4310 3384
rect 4425 3380 4429 3384
rect 4445 3380 4449 3384
rect 4531 3380 4535 3384
rect 4551 3380 4555 3384
rect 4611 3380 4615 3384
rect 4633 3380 4637 3384
rect 4641 3380 4645 3384
rect 4661 3380 4665 3384
rect 4669 3380 4673 3384
rect 4715 3380 4719 3384
rect 4735 3380 4739 3384
rect 4747 3380 4751 3384
rect 4767 3380 4771 3384
rect 4781 3380 4785 3384
rect 4801 3380 4805 3384
rect 4905 3380 4909 3384
rect 4925 3380 4929 3384
rect 5030 3380 5034 3384
rect 5052 3380 5056 3384
rect 5060 3380 5064 3384
rect 5171 3380 5175 3384
rect 5191 3380 5195 3384
rect 5255 3380 5259 3384
rect 5275 3380 5279 3384
rect 5289 3380 5293 3384
rect 5309 3380 5313 3384
rect 5321 3380 5325 3384
rect 5341 3380 5345 3384
rect 5387 3380 5391 3384
rect 5395 3380 5399 3384
rect 5415 3380 5419 3384
rect 5423 3380 5427 3384
rect 5445 3380 5449 3384
rect 5545 3380 5549 3384
rect 5565 3380 5569 3384
rect 5656 3380 5660 3384
rect 5664 3380 5668 3384
rect 5686 3380 5690 3384
rect 85 3356 89 3360
rect 190 3356 194 3360
rect 212 3356 216 3360
rect 220 3356 224 3360
rect 325 3356 329 3360
rect 411 3356 415 3360
rect 431 3356 435 3360
rect 531 3356 535 3360
rect 551 3356 555 3360
rect 571 3356 575 3360
rect 671 3356 675 3360
rect 693 3356 697 3360
rect 715 3356 719 3360
rect 845 3356 849 3360
rect 865 3356 869 3360
rect 965 3356 969 3360
rect 985 3356 989 3360
rect 1005 3356 1009 3360
rect 1105 3356 1109 3360
rect 1125 3356 1129 3360
rect 1145 3356 1149 3360
rect 1231 3356 1235 3360
rect 1251 3356 1255 3360
rect 1271 3356 1275 3360
rect 1385 3356 1389 3360
rect 1485 3356 1489 3360
rect 1505 3356 1509 3360
rect 1525 3356 1529 3360
rect 1625 3356 1629 3360
rect 1645 3356 1649 3360
rect 1665 3356 1669 3360
rect 1765 3356 1769 3360
rect 1785 3356 1789 3360
rect 1805 3356 1809 3360
rect 1925 3356 1929 3360
rect 1945 3356 1949 3360
rect 2045 3356 2049 3360
rect 2065 3356 2069 3360
rect 2085 3356 2089 3360
rect 2171 3356 2175 3360
rect 2191 3356 2195 3360
rect 2301 3356 2305 3360
rect 2323 3356 2327 3360
rect 2345 3356 2349 3360
rect 2431 3356 2435 3360
rect 2451 3356 2455 3360
rect 2570 3356 2574 3360
rect 2592 3356 2596 3360
rect 2600 3356 2604 3360
rect 2705 3356 2709 3360
rect 2725 3356 2729 3360
rect 2745 3356 2749 3360
rect 2831 3356 2835 3360
rect 2851 3356 2855 3360
rect 2871 3356 2875 3360
rect 2971 3356 2975 3360
rect 2991 3356 2995 3360
rect 3011 3356 3015 3360
rect 3125 3356 3129 3360
rect 3145 3356 3149 3360
rect 3265 3356 3269 3360
rect 3285 3356 3289 3360
rect 3371 3356 3375 3360
rect 3485 3356 3489 3360
rect 3505 3356 3509 3360
rect 3525 3356 3529 3360
rect 3611 3356 3615 3360
rect 3631 3356 3635 3360
rect 3651 3356 3655 3360
rect 3770 3356 3774 3360
rect 3792 3356 3796 3360
rect 3800 3356 3804 3360
rect 3891 3356 3895 3360
rect 3951 3356 3955 3360
rect 3973 3356 3977 3360
rect 3981 3356 3985 3360
rect 4001 3356 4005 3360
rect 4009 3356 4013 3360
rect 4055 3356 4059 3360
rect 4075 3356 4079 3360
rect 4087 3356 4091 3360
rect 4107 3356 4111 3360
rect 4121 3356 4125 3360
rect 4141 3356 4145 3360
rect 4236 3356 4240 3360
rect 4244 3356 4248 3360
rect 4266 3356 4270 3360
rect 4376 3356 4380 3360
rect 4384 3356 4388 3360
rect 4406 3356 4410 3360
rect 4471 3356 4475 3360
rect 4493 3356 4497 3360
rect 4501 3356 4505 3360
rect 4521 3356 4525 3360
rect 4529 3356 4533 3360
rect 4575 3356 4579 3360
rect 4595 3356 4599 3360
rect 4607 3356 4611 3360
rect 4627 3356 4631 3360
rect 4641 3356 4645 3360
rect 4661 3356 4665 3360
rect 4756 3356 4760 3360
rect 4764 3356 4768 3360
rect 4786 3356 4790 3360
rect 4905 3356 4909 3360
rect 4925 3356 4929 3360
rect 5030 3356 5034 3360
rect 5052 3356 5056 3360
rect 5060 3356 5064 3360
rect 5165 3356 5169 3360
rect 5265 3356 5269 3360
rect 5285 3356 5289 3360
rect 5371 3356 5375 3360
rect 5496 3356 5500 3360
rect 5504 3356 5508 3360
rect 5526 3356 5530 3360
rect 5665 3356 5669 3360
rect 5685 3356 5689 3360
rect 85 3233 89 3316
rect 190 3273 194 3316
rect 187 3261 194 3273
rect 85 3221 94 3233
rect 85 3164 89 3221
rect 185 3184 189 3261
rect 212 3219 216 3276
rect 220 3272 224 3276
rect 220 3264 238 3272
rect 234 3253 238 3264
rect 205 3207 214 3219
rect 205 3184 209 3207
rect 234 3196 238 3241
rect 225 3189 238 3196
rect 325 3233 329 3316
rect 411 3239 415 3316
rect 325 3221 334 3233
rect 406 3227 415 3239
rect 225 3184 229 3189
rect 325 3164 329 3221
rect 409 3211 415 3227
rect 431 3239 435 3316
rect 531 3262 535 3276
rect 551 3262 555 3276
rect 519 3256 535 3262
rect 540 3256 555 3262
rect 431 3227 434 3239
rect 431 3211 437 3227
rect 519 3219 526 3256
rect 540 3233 546 3256
rect 409 3204 417 3211
rect 413 3184 417 3204
rect 423 3204 437 3211
rect 423 3184 427 3204
rect 519 3194 526 3207
rect 519 3188 538 3194
rect 534 3184 538 3188
rect 542 3184 546 3221
rect 571 3219 575 3276
rect 671 3253 675 3316
rect 666 3241 675 3253
rect 566 3207 575 3219
rect 564 3164 568 3207
rect 671 3184 675 3241
rect 693 3239 697 3316
rect 681 3227 694 3239
rect 681 3184 685 3227
rect 715 3202 719 3276
rect 845 3239 849 3316
rect 846 3227 849 3239
rect 843 3211 849 3227
rect 865 3239 869 3316
rect 965 3273 969 3316
rect 985 3304 989 3316
rect 1005 3308 1009 3316
rect 1005 3304 1020 3308
rect 985 3300 1000 3304
rect 994 3293 1000 3300
rect 965 3261 973 3273
rect 985 3261 992 3273
rect 865 3227 874 3239
rect 865 3211 871 3227
rect 843 3204 857 3211
rect 707 3190 719 3202
rect 701 3184 705 3190
rect 853 3184 857 3204
rect 863 3204 871 3211
rect 988 3204 992 3261
rect 996 3204 1000 3281
rect 1014 3273 1020 3304
rect 1105 3273 1109 3316
rect 1125 3304 1129 3316
rect 1145 3308 1149 3316
rect 1145 3304 1160 3308
rect 1125 3300 1140 3304
rect 1134 3293 1140 3300
rect 1004 3261 1014 3273
rect 1105 3261 1113 3273
rect 1125 3261 1132 3273
rect 1004 3204 1008 3261
rect 1128 3204 1132 3261
rect 1136 3204 1140 3281
rect 1154 3273 1160 3304
rect 1144 3261 1154 3273
rect 1231 3262 1235 3276
rect 1251 3262 1255 3276
rect 1144 3204 1148 3261
rect 1219 3256 1235 3262
rect 1240 3256 1255 3262
rect 1219 3219 1226 3256
rect 1240 3233 1246 3256
rect 863 3184 867 3204
rect 1219 3194 1226 3207
rect 1219 3188 1238 3194
rect 1234 3184 1238 3188
rect 1242 3184 1246 3221
rect 1271 3219 1275 3276
rect 1266 3207 1275 3219
rect 1385 3233 1389 3316
rect 1485 3273 1489 3316
rect 1505 3304 1509 3316
rect 1525 3308 1529 3316
rect 1525 3304 1540 3308
rect 1505 3300 1520 3304
rect 1514 3293 1520 3300
rect 1485 3261 1493 3273
rect 1505 3261 1512 3273
rect 1385 3221 1394 3233
rect 1264 3164 1268 3207
rect 1385 3164 1389 3221
rect 1508 3204 1512 3261
rect 1516 3204 1520 3281
rect 1534 3273 1540 3304
rect 1625 3273 1629 3316
rect 1645 3304 1649 3316
rect 1665 3308 1669 3316
rect 1665 3304 1680 3308
rect 1645 3300 1660 3304
rect 1654 3293 1660 3300
rect 1524 3261 1534 3273
rect 1625 3261 1633 3273
rect 1645 3261 1652 3273
rect 1524 3204 1528 3261
rect 1648 3204 1652 3261
rect 1656 3204 1660 3281
rect 1674 3273 1680 3304
rect 1664 3261 1674 3273
rect 1664 3204 1668 3261
rect 1765 3219 1769 3276
rect 1785 3262 1789 3276
rect 1805 3262 1809 3276
rect 1785 3256 1800 3262
rect 1805 3256 1821 3262
rect 1794 3233 1800 3256
rect 1765 3207 1774 3219
rect 1772 3164 1776 3207
rect 1794 3184 1798 3221
rect 1814 3219 1821 3256
rect 1925 3239 1929 3316
rect 1926 3227 1929 3239
rect 1923 3211 1929 3227
rect 1945 3239 1949 3316
rect 1945 3227 1954 3239
rect 1945 3211 1951 3227
rect 1814 3194 1821 3207
rect 1923 3204 1937 3211
rect 1802 3188 1821 3194
rect 1802 3184 1806 3188
rect 1933 3184 1937 3204
rect 1943 3204 1951 3211
rect 2045 3219 2049 3276
rect 2065 3262 2069 3276
rect 2085 3262 2089 3276
rect 2065 3256 2080 3262
rect 2085 3256 2101 3262
rect 2074 3233 2080 3256
rect 2045 3207 2054 3219
rect 1943 3184 1947 3204
rect 2052 3164 2056 3207
rect 2074 3184 2078 3221
rect 2094 3219 2101 3256
rect 2171 3239 2175 3316
rect 2166 3227 2175 3239
rect 2169 3211 2175 3227
rect 2191 3239 2195 3316
rect 2191 3227 2194 3239
rect 2191 3211 2197 3227
rect 2094 3194 2101 3207
rect 2169 3204 2177 3211
rect 2082 3188 2101 3194
rect 2082 3184 2086 3188
rect 2173 3184 2177 3204
rect 2183 3204 2197 3211
rect 2183 3184 2187 3204
rect 2301 3202 2305 3276
rect 2323 3239 2327 3316
rect 2345 3253 2349 3316
rect 2345 3241 2354 3253
rect 2326 3227 2339 3239
rect 2301 3190 2313 3202
rect 2315 3184 2319 3190
rect 2335 3184 2339 3227
rect 2345 3184 2349 3241
rect 2431 3239 2435 3316
rect 2426 3227 2435 3239
rect 2429 3211 2435 3227
rect 2451 3239 2455 3316
rect 2570 3273 2574 3316
rect 2831 3308 2835 3316
rect 2820 3304 2835 3308
rect 2851 3304 2855 3316
rect 2567 3261 2574 3273
rect 2451 3227 2454 3239
rect 2451 3211 2457 3227
rect 2429 3204 2437 3211
rect 2433 3184 2437 3204
rect 2443 3204 2457 3211
rect 2443 3184 2447 3204
rect 2565 3184 2569 3261
rect 2592 3219 2596 3276
rect 2600 3272 2604 3276
rect 2600 3264 2618 3272
rect 2614 3253 2618 3264
rect 2585 3207 2594 3219
rect 2585 3184 2589 3207
rect 2614 3196 2618 3241
rect 2705 3219 2709 3276
rect 2725 3262 2729 3276
rect 2745 3262 2749 3276
rect 2820 3273 2826 3304
rect 2840 3300 2855 3304
rect 2840 3293 2846 3300
rect 2725 3256 2740 3262
rect 2745 3256 2761 3262
rect 2826 3261 2836 3273
rect 2734 3233 2740 3256
rect 2705 3207 2714 3219
rect 2605 3189 2618 3196
rect 2605 3184 2609 3189
rect 2712 3164 2716 3207
rect 2734 3184 2738 3221
rect 2754 3219 2761 3256
rect 2754 3194 2761 3207
rect 2832 3204 2836 3261
rect 2840 3204 2844 3281
rect 2871 3273 2875 3316
rect 2971 3308 2975 3316
rect 2960 3304 2975 3308
rect 2991 3304 2995 3316
rect 2960 3273 2966 3304
rect 2980 3300 2995 3304
rect 2980 3293 2986 3300
rect 2848 3261 2855 3273
rect 2867 3261 2875 3273
rect 2966 3261 2976 3273
rect 2848 3204 2852 3261
rect 2972 3204 2976 3261
rect 2980 3204 2984 3281
rect 3011 3273 3015 3316
rect 2988 3261 2995 3273
rect 3007 3261 3015 3273
rect 2988 3204 2992 3261
rect 3125 3239 3129 3316
rect 3126 3227 3129 3239
rect 3123 3211 3129 3227
rect 3145 3239 3149 3316
rect 3265 3239 3269 3316
rect 3145 3227 3154 3239
rect 3266 3227 3269 3239
rect 3145 3211 3151 3227
rect 3123 3204 3137 3211
rect 2742 3188 2761 3194
rect 2742 3184 2746 3188
rect 3133 3184 3137 3204
rect 3143 3204 3151 3211
rect 3263 3211 3269 3227
rect 3285 3239 3289 3316
rect 3285 3227 3294 3239
rect 3371 3233 3375 3316
rect 3485 3273 3489 3316
rect 3505 3304 3509 3316
rect 3525 3308 3529 3316
rect 3525 3304 3540 3308
rect 3505 3300 3520 3304
rect 3514 3293 3520 3300
rect 3485 3261 3493 3273
rect 3505 3261 3512 3273
rect 3285 3211 3291 3227
rect 3366 3221 3375 3233
rect 3263 3204 3277 3211
rect 3143 3184 3147 3204
rect 3273 3184 3277 3204
rect 3283 3204 3291 3211
rect 3283 3184 3287 3204
rect 3371 3164 3375 3221
rect 3508 3204 3512 3261
rect 3516 3204 3520 3281
rect 3534 3273 3540 3304
rect 3524 3261 3534 3273
rect 3611 3262 3615 3276
rect 3631 3262 3635 3276
rect 3524 3204 3528 3261
rect 3599 3256 3615 3262
rect 3620 3256 3635 3262
rect 3599 3219 3606 3256
rect 3620 3233 3626 3256
rect 3599 3194 3606 3207
rect 3599 3188 3618 3194
rect 3614 3184 3618 3188
rect 3622 3184 3626 3221
rect 3651 3219 3655 3276
rect 3770 3273 3774 3316
rect 3767 3261 3774 3273
rect 3646 3207 3655 3219
rect 3644 3164 3648 3207
rect 3765 3184 3769 3261
rect 3792 3219 3796 3276
rect 3800 3272 3804 3276
rect 3800 3264 3818 3272
rect 3814 3253 3818 3264
rect 3785 3207 3794 3219
rect 3785 3184 3789 3207
rect 3814 3196 3818 3241
rect 3891 3233 3895 3316
rect 3973 3313 3977 3336
rect 3969 3306 3977 3313
rect 3969 3277 3973 3306
rect 3981 3296 3985 3336
rect 4001 3284 4005 3316
rect 4009 3312 4013 3316
rect 4009 3310 4045 3312
rect 4009 3308 4033 3310
rect 3886 3221 3895 3233
rect 3805 3189 3818 3196
rect 3805 3184 3809 3189
rect 3891 3164 3895 3221
rect 3951 3264 3955 3276
rect 3969 3271 3977 3277
rect 3951 3252 3953 3264
rect 3951 3184 3955 3252
rect 3973 3225 3977 3271
rect 3973 3164 3977 3213
rect 4001 3189 4007 3284
rect 3983 3185 4007 3189
rect 3983 3164 3987 3185
rect 4003 3180 4021 3181
rect 4003 3176 4033 3180
rect 4003 3164 4007 3176
rect 4041 3172 4045 3298
rect 4055 3290 4059 3316
rect 4075 3310 4079 3316
rect 4011 3168 4045 3172
rect 4011 3164 4015 3168
rect 4057 3164 4061 3278
rect 4073 3188 4077 3298
rect 4087 3276 4091 3316
rect 4082 3264 4085 3276
rect 4082 3200 4086 3264
rect 4107 3257 4111 3316
rect 4102 3249 4111 3257
rect 4102 3220 4106 3249
rect 4121 3234 4125 3316
rect 4141 3233 4145 3276
rect 4236 3272 4240 3276
rect 4222 3264 4240 3272
rect 4222 3253 4226 3264
rect 4082 3196 4115 3200
rect 4081 3176 4083 3188
rect 4079 3164 4083 3176
rect 4089 3176 4091 3188
rect 4089 3164 4093 3176
rect 4111 3164 4115 3196
rect 4121 3164 4125 3222
rect 4141 3184 4145 3221
rect 4222 3196 4226 3241
rect 4244 3219 4248 3276
rect 4266 3273 4270 3316
rect 4266 3261 4273 3273
rect 4376 3272 4380 3276
rect 4362 3264 4380 3272
rect 4246 3207 4255 3219
rect 4222 3189 4235 3196
rect 4231 3184 4235 3189
rect 4251 3184 4255 3207
rect 4271 3184 4275 3261
rect 4362 3253 4366 3264
rect 4362 3196 4366 3241
rect 4384 3219 4388 3276
rect 4406 3273 4410 3316
rect 4493 3313 4497 3336
rect 4489 3306 4497 3313
rect 4489 3277 4493 3306
rect 4501 3296 4505 3336
rect 4521 3284 4525 3316
rect 4529 3312 4533 3316
rect 4529 3310 4565 3312
rect 4529 3308 4553 3310
rect 4406 3261 4413 3273
rect 4471 3264 4475 3276
rect 4489 3271 4497 3277
rect 4386 3207 4395 3219
rect 4362 3189 4375 3196
rect 4371 3184 4375 3189
rect 4391 3184 4395 3207
rect 4411 3184 4415 3261
rect 4471 3252 4473 3264
rect 4471 3184 4475 3252
rect 4493 3225 4497 3271
rect 4493 3164 4497 3213
rect 4521 3189 4527 3284
rect 4503 3185 4527 3189
rect 4503 3164 4507 3185
rect 4523 3180 4541 3181
rect 4523 3176 4553 3180
rect 4523 3164 4527 3176
rect 4561 3172 4565 3298
rect 4575 3290 4579 3316
rect 4595 3310 4599 3316
rect 4531 3168 4565 3172
rect 4531 3164 4535 3168
rect 4577 3164 4581 3278
rect 4593 3188 4597 3298
rect 4607 3276 4611 3316
rect 4602 3264 4605 3276
rect 4602 3200 4606 3264
rect 4627 3257 4631 3316
rect 4622 3249 4631 3257
rect 4622 3220 4626 3249
rect 4641 3234 4645 3316
rect 4661 3233 4665 3276
rect 4756 3272 4760 3276
rect 4742 3264 4760 3272
rect 4742 3253 4746 3264
rect 4602 3196 4635 3200
rect 4601 3176 4603 3188
rect 4599 3164 4603 3176
rect 4609 3176 4611 3188
rect 4609 3164 4613 3176
rect 4631 3164 4635 3196
rect 4641 3164 4645 3222
rect 4661 3184 4665 3221
rect 4742 3196 4746 3241
rect 4764 3219 4768 3276
rect 4786 3273 4790 3316
rect 4786 3261 4793 3273
rect 4766 3207 4775 3219
rect 4742 3189 4755 3196
rect 4751 3184 4755 3189
rect 4771 3184 4775 3207
rect 4791 3184 4795 3261
rect 4905 3239 4909 3316
rect 4906 3227 4909 3239
rect 4903 3211 4909 3227
rect 4925 3239 4929 3316
rect 5030 3273 5034 3316
rect 5027 3261 5034 3273
rect 4925 3227 4934 3239
rect 4925 3211 4931 3227
rect 4903 3204 4917 3211
rect 4913 3184 4917 3204
rect 4923 3204 4931 3211
rect 4923 3184 4927 3204
rect 5025 3184 5029 3261
rect 5052 3219 5056 3276
rect 5060 3272 5064 3276
rect 5060 3264 5078 3272
rect 5074 3253 5078 3264
rect 5045 3207 5054 3219
rect 5045 3184 5049 3207
rect 5074 3196 5078 3241
rect 5065 3189 5078 3196
rect 5165 3233 5169 3316
rect 5265 3239 5269 3316
rect 5165 3221 5174 3233
rect 5266 3227 5269 3239
rect 5065 3184 5069 3189
rect 5165 3164 5169 3221
rect 5263 3211 5269 3227
rect 5285 3239 5289 3316
rect 5285 3227 5294 3239
rect 5371 3233 5375 3316
rect 5496 3272 5500 3276
rect 5482 3264 5500 3272
rect 5482 3253 5486 3264
rect 5285 3211 5291 3227
rect 5366 3221 5375 3233
rect 5263 3204 5277 3211
rect 5273 3184 5277 3204
rect 5283 3204 5291 3211
rect 5283 3184 5287 3204
rect 5371 3164 5375 3221
rect 5482 3196 5486 3241
rect 5504 3219 5508 3276
rect 5526 3273 5530 3316
rect 5526 3261 5533 3273
rect 5506 3207 5515 3219
rect 5482 3189 5495 3196
rect 5491 3184 5495 3189
rect 5511 3184 5515 3207
rect 5531 3184 5535 3261
rect 5665 3239 5669 3316
rect 5666 3227 5669 3239
rect 5663 3211 5669 3227
rect 5685 3239 5689 3316
rect 5685 3227 5694 3239
rect 5685 3211 5691 3227
rect 5663 3204 5677 3211
rect 5673 3184 5677 3204
rect 5683 3204 5691 3211
rect 5683 3184 5687 3204
rect 85 3140 89 3144
rect 185 3140 189 3144
rect 205 3140 209 3144
rect 225 3140 229 3144
rect 325 3140 329 3144
rect 413 3140 417 3144
rect 423 3140 427 3144
rect 534 3140 538 3144
rect 542 3140 546 3144
rect 564 3140 568 3144
rect 671 3140 675 3144
rect 681 3140 685 3144
rect 701 3140 705 3144
rect 853 3140 857 3144
rect 863 3140 867 3144
rect 988 3140 992 3144
rect 996 3140 1000 3144
rect 1004 3140 1008 3144
rect 1128 3140 1132 3144
rect 1136 3140 1140 3144
rect 1144 3140 1148 3144
rect 1234 3140 1238 3144
rect 1242 3140 1246 3144
rect 1264 3140 1268 3144
rect 1385 3140 1389 3144
rect 1508 3140 1512 3144
rect 1516 3140 1520 3144
rect 1524 3140 1528 3144
rect 1648 3140 1652 3144
rect 1656 3140 1660 3144
rect 1664 3140 1668 3144
rect 1772 3140 1776 3144
rect 1794 3140 1798 3144
rect 1802 3140 1806 3144
rect 1933 3140 1937 3144
rect 1943 3140 1947 3144
rect 2052 3140 2056 3144
rect 2074 3140 2078 3144
rect 2082 3140 2086 3144
rect 2173 3140 2177 3144
rect 2183 3140 2187 3144
rect 2315 3140 2319 3144
rect 2335 3140 2339 3144
rect 2345 3140 2349 3144
rect 2433 3140 2437 3144
rect 2443 3140 2447 3144
rect 2565 3140 2569 3144
rect 2585 3140 2589 3144
rect 2605 3140 2609 3144
rect 2712 3140 2716 3144
rect 2734 3140 2738 3144
rect 2742 3140 2746 3144
rect 2832 3140 2836 3144
rect 2840 3140 2844 3144
rect 2848 3140 2852 3144
rect 2972 3140 2976 3144
rect 2980 3140 2984 3144
rect 2988 3140 2992 3144
rect 3133 3140 3137 3144
rect 3143 3140 3147 3144
rect 3273 3140 3277 3144
rect 3283 3140 3287 3144
rect 3371 3140 3375 3144
rect 3508 3140 3512 3144
rect 3516 3140 3520 3144
rect 3524 3140 3528 3144
rect 3614 3140 3618 3144
rect 3622 3140 3626 3144
rect 3644 3140 3648 3144
rect 3765 3140 3769 3144
rect 3785 3140 3789 3144
rect 3805 3140 3809 3144
rect 3891 3140 3895 3144
rect 3951 3140 3955 3144
rect 3973 3140 3977 3144
rect 3983 3140 3987 3144
rect 4003 3140 4007 3144
rect 4011 3140 4015 3144
rect 4057 3140 4061 3144
rect 4079 3140 4083 3144
rect 4089 3140 4093 3144
rect 4111 3140 4115 3144
rect 4121 3140 4125 3144
rect 4141 3140 4145 3144
rect 4231 3140 4235 3144
rect 4251 3140 4255 3144
rect 4271 3140 4275 3144
rect 4371 3140 4375 3144
rect 4391 3140 4395 3144
rect 4411 3140 4415 3144
rect 4471 3140 4475 3144
rect 4493 3140 4497 3144
rect 4503 3140 4507 3144
rect 4523 3140 4527 3144
rect 4531 3140 4535 3144
rect 4577 3140 4581 3144
rect 4599 3140 4603 3144
rect 4609 3140 4613 3144
rect 4631 3140 4635 3144
rect 4641 3140 4645 3144
rect 4661 3140 4665 3144
rect 4751 3140 4755 3144
rect 4771 3140 4775 3144
rect 4791 3140 4795 3144
rect 4913 3140 4917 3144
rect 4923 3140 4927 3144
rect 5025 3140 5029 3144
rect 5045 3140 5049 3144
rect 5065 3140 5069 3144
rect 5165 3140 5169 3144
rect 5273 3140 5277 3144
rect 5283 3140 5287 3144
rect 5371 3140 5375 3144
rect 5491 3140 5495 3144
rect 5511 3140 5515 3144
rect 5531 3140 5535 3144
rect 5673 3140 5677 3144
rect 5683 3140 5687 3144
rect 115 3116 119 3120
rect 135 3116 139 3120
rect 145 3116 149 3120
rect 252 3116 256 3120
rect 260 3116 264 3120
rect 268 3116 272 3120
rect 393 3116 397 3120
rect 403 3116 407 3120
rect 525 3116 529 3120
rect 545 3116 549 3120
rect 565 3116 569 3120
rect 651 3116 655 3120
rect 671 3116 675 3120
rect 691 3116 695 3120
rect 791 3116 795 3120
rect 811 3116 815 3120
rect 831 3116 835 3120
rect 931 3116 935 3120
rect 951 3116 955 3120
rect 971 3116 975 3120
rect 1093 3116 1097 3120
rect 1103 3116 1107 3120
rect 1225 3116 1229 3120
rect 1245 3116 1249 3120
rect 1331 3116 1335 3120
rect 1351 3116 1355 3120
rect 1371 3116 1375 3120
rect 1508 3116 1512 3120
rect 1516 3116 1520 3120
rect 1524 3116 1528 3120
rect 1652 3116 1656 3120
rect 1674 3116 1678 3120
rect 1682 3116 1686 3120
rect 1785 3116 1789 3120
rect 1805 3116 1809 3120
rect 1825 3116 1829 3120
rect 1911 3116 1915 3120
rect 1931 3116 1935 3120
rect 1951 3116 1955 3120
rect 2085 3116 2089 3120
rect 2105 3116 2109 3120
rect 2125 3116 2129 3120
rect 2225 3116 2229 3120
rect 2245 3116 2249 3120
rect 2265 3116 2269 3120
rect 2392 3116 2396 3120
rect 2414 3116 2418 3120
rect 2422 3116 2426 3120
rect 2532 3116 2536 3120
rect 2554 3116 2558 3120
rect 2562 3116 2566 3120
rect 2686 3116 2690 3120
rect 2694 3116 2698 3120
rect 2714 3116 2718 3120
rect 2722 3116 2726 3120
rect 2825 3116 2829 3120
rect 2845 3116 2849 3120
rect 2865 3116 2869 3120
rect 2951 3116 2955 3120
rect 2971 3116 2975 3120
rect 3093 3116 3097 3120
rect 3103 3116 3107 3120
rect 3235 3116 3239 3120
rect 3255 3116 3259 3120
rect 3265 3116 3269 3120
rect 3351 3116 3355 3120
rect 3371 3116 3375 3120
rect 3391 3116 3395 3120
rect 3505 3116 3509 3120
rect 3525 3116 3529 3120
rect 3545 3116 3549 3120
rect 3645 3116 3649 3120
rect 3665 3116 3669 3120
rect 3685 3116 3689 3120
rect 3785 3116 3789 3120
rect 3805 3116 3809 3120
rect 3825 3116 3829 3120
rect 3955 3116 3959 3120
rect 3975 3116 3979 3120
rect 3985 3116 3989 3120
rect 4071 3116 4075 3120
rect 4091 3116 4095 3120
rect 4192 3116 4196 3120
rect 4200 3116 4204 3120
rect 4208 3116 4212 3120
rect 4295 3116 4299 3120
rect 4315 3116 4319 3120
rect 4325 3116 4329 3120
rect 4347 3116 4351 3120
rect 4357 3116 4361 3120
rect 4379 3116 4383 3120
rect 4425 3116 4429 3120
rect 4433 3116 4437 3120
rect 4453 3116 4457 3120
rect 4463 3116 4467 3120
rect 4485 3116 4489 3120
rect 4591 3116 4595 3120
rect 4611 3116 4615 3120
rect 4631 3116 4635 3120
rect 4731 3116 4735 3120
rect 4751 3116 4755 3120
rect 4771 3116 4775 3120
rect 4893 3116 4897 3120
rect 4903 3116 4907 3120
rect 4993 3116 4997 3120
rect 5003 3116 5007 3120
rect 5075 3116 5079 3120
rect 5095 3116 5099 3120
rect 5105 3116 5109 3120
rect 5127 3116 5131 3120
rect 5137 3116 5141 3120
rect 5159 3116 5163 3120
rect 5205 3116 5209 3120
rect 5213 3116 5217 3120
rect 5233 3116 5237 3120
rect 5243 3116 5247 3120
rect 5265 3116 5269 3120
rect 5365 3116 5369 3120
rect 5385 3116 5389 3120
rect 5405 3116 5409 3120
rect 5425 3116 5429 3120
rect 5445 3116 5449 3120
rect 5465 3116 5469 3120
rect 5485 3116 5489 3120
rect 5505 3116 5509 3120
rect 5551 3116 5555 3120
rect 5573 3116 5577 3120
rect 5583 3116 5587 3120
rect 5603 3116 5607 3120
rect 5611 3116 5615 3120
rect 5657 3116 5661 3120
rect 5679 3116 5683 3120
rect 5689 3116 5693 3120
rect 5711 3116 5715 3120
rect 5721 3116 5725 3120
rect 5741 3116 5745 3120
rect 115 3070 119 3076
rect 101 3058 113 3070
rect 101 2984 105 3058
rect 135 3033 139 3076
rect 126 3021 139 3033
rect 123 2944 127 3021
rect 145 3019 149 3076
rect 393 3056 397 3076
rect 145 3007 154 3019
rect 145 2944 149 3007
rect 252 2999 256 3056
rect 246 2987 256 2999
rect 240 2956 246 2987
rect 260 2979 264 3056
rect 268 2999 272 3056
rect 389 3049 397 3056
rect 403 3056 407 3076
rect 403 3049 417 3056
rect 389 3033 395 3049
rect 386 3021 395 3033
rect 268 2987 275 2999
rect 287 2987 295 2999
rect 260 2960 266 2967
rect 260 2956 275 2960
rect 240 2952 255 2956
rect 251 2944 255 2952
rect 271 2944 275 2956
rect 291 2944 295 2987
rect 391 2944 395 3021
rect 411 3033 417 3049
rect 411 3021 414 3033
rect 411 2944 415 3021
rect 525 2999 529 3076
rect 545 3053 549 3076
rect 565 3071 569 3076
rect 651 3071 655 3076
rect 565 3064 578 3071
rect 545 3041 554 3053
rect 527 2987 534 2999
rect 530 2944 534 2987
rect 552 2984 556 3041
rect 574 3019 578 3064
rect 642 3064 655 3071
rect 642 3019 646 3064
rect 671 3053 675 3076
rect 666 3041 675 3053
rect 574 2996 578 3007
rect 560 2988 578 2996
rect 642 2996 646 3007
rect 642 2988 660 2996
rect 560 2984 564 2988
rect 656 2984 660 2988
rect 664 2984 668 3041
rect 691 2999 695 3076
rect 791 3071 795 3076
rect 782 3064 795 3071
rect 782 3019 786 3064
rect 811 3053 815 3076
rect 806 3041 815 3053
rect 686 2987 693 2999
rect 782 2996 786 3007
rect 782 2988 800 2996
rect 686 2944 690 2987
rect 796 2984 800 2988
rect 804 2984 808 3041
rect 831 2999 835 3076
rect 931 3071 935 3076
rect 922 3064 935 3071
rect 922 3019 926 3064
rect 951 3053 955 3076
rect 946 3041 955 3053
rect 826 2987 833 2999
rect 922 2996 926 3007
rect 922 2988 940 2996
rect 826 2944 830 2987
rect 936 2984 940 2988
rect 944 2984 948 3041
rect 971 2999 975 3076
rect 1093 3056 1097 3076
rect 1083 3049 1097 3056
rect 1103 3056 1107 3076
rect 1103 3049 1111 3056
rect 1083 3033 1089 3049
rect 1086 3021 1089 3033
rect 966 2987 973 2999
rect 966 2944 970 2987
rect 1085 2944 1089 3021
rect 1105 3033 1111 3049
rect 1105 3021 1114 3033
rect 1105 2944 1109 3021
rect 1225 3019 1229 3096
rect 1245 3019 1249 3096
rect 1331 3071 1335 3076
rect 1322 3064 1335 3071
rect 1322 3019 1326 3064
rect 1351 3053 1355 3076
rect 1346 3041 1355 3053
rect 1226 3007 1241 3019
rect 1237 2984 1241 3007
rect 1245 3007 1254 3019
rect 1245 2984 1249 3007
rect 1322 2996 1326 3007
rect 1322 2988 1340 2996
rect 1336 2984 1340 2988
rect 1344 2984 1348 3041
rect 1371 2999 1375 3076
rect 1508 2999 1512 3056
rect 1366 2987 1373 2999
rect 1485 2987 1493 2999
rect 1505 2987 1512 2999
rect 1366 2944 1370 2987
rect 1485 2944 1489 2987
rect 1516 2979 1520 3056
rect 1524 2999 1528 3056
rect 1652 3053 1656 3096
rect 1645 3041 1654 3053
rect 1524 2987 1534 2999
rect 1514 2960 1520 2967
rect 1505 2956 1520 2960
rect 1534 2956 1540 2987
rect 1645 2984 1649 3041
rect 1674 3039 1678 3076
rect 1682 3072 1686 3076
rect 1682 3066 1701 3072
rect 1694 3053 1701 3066
rect 1674 3004 1680 3027
rect 1694 3004 1701 3041
rect 1665 2998 1680 3004
rect 1685 2998 1701 3004
rect 1785 2999 1789 3076
rect 1805 3053 1809 3076
rect 1825 3071 1829 3076
rect 1911 3071 1915 3076
rect 1825 3064 1838 3071
rect 1805 3041 1814 3053
rect 1665 2984 1669 2998
rect 1685 2984 1689 2998
rect 1787 2987 1794 2999
rect 1505 2944 1509 2956
rect 1525 2952 1540 2956
rect 1525 2944 1529 2952
rect 1790 2944 1794 2987
rect 1812 2984 1816 3041
rect 1834 3019 1838 3064
rect 1902 3064 1915 3071
rect 1902 3019 1906 3064
rect 1931 3053 1935 3076
rect 1926 3041 1935 3053
rect 1834 2996 1838 3007
rect 1820 2988 1838 2996
rect 1902 2996 1906 3007
rect 1902 2988 1920 2996
rect 1820 2984 1824 2988
rect 1916 2984 1920 2988
rect 1924 2984 1928 3041
rect 1951 2999 1955 3076
rect 2085 2999 2089 3076
rect 2105 3053 2109 3076
rect 2125 3071 2129 3076
rect 2125 3064 2138 3071
rect 2105 3041 2114 3053
rect 1946 2987 1953 2999
rect 2087 2987 2094 2999
rect 1946 2944 1950 2987
rect 2090 2944 2094 2987
rect 2112 2984 2116 3041
rect 2134 3019 2138 3064
rect 2134 2996 2138 3007
rect 2225 2999 2229 3076
rect 2245 3053 2249 3076
rect 2265 3071 2269 3076
rect 2265 3064 2278 3071
rect 2245 3041 2254 3053
rect 2120 2988 2138 2996
rect 2120 2984 2124 2988
rect 2227 2987 2234 2999
rect 2230 2944 2234 2987
rect 2252 2984 2256 3041
rect 2274 3019 2278 3064
rect 2392 3053 2396 3096
rect 2385 3041 2394 3053
rect 2274 2996 2278 3007
rect 2260 2988 2278 2996
rect 2260 2984 2264 2988
rect 2385 2984 2389 3041
rect 2414 3039 2418 3076
rect 2422 3072 2426 3076
rect 2422 3066 2441 3072
rect 2434 3053 2441 3066
rect 2532 3053 2536 3096
rect 2845 3089 2849 3096
rect 2865 3089 2869 3096
rect 2845 3083 2859 3089
rect 2865 3084 2878 3089
rect 2525 3041 2534 3053
rect 2414 3004 2420 3027
rect 2434 3004 2441 3041
rect 2405 2998 2420 3004
rect 2425 2998 2441 3004
rect 2405 2984 2409 2998
rect 2425 2984 2429 2998
rect 2525 2984 2529 3041
rect 2554 3039 2558 3076
rect 2562 3072 2566 3076
rect 2562 3066 2581 3072
rect 2686 3071 2690 3076
rect 2574 3053 2581 3066
rect 2660 3067 2690 3071
rect 2554 3004 2560 3027
rect 2574 3004 2581 3041
rect 2660 3019 2666 3067
rect 2694 3062 2698 3076
rect 2685 3055 2698 3062
rect 2685 3053 2689 3055
rect 2714 3053 2718 3076
rect 2722 3068 2726 3076
rect 2825 3068 2829 3076
rect 2722 3061 2739 3068
rect 2687 3041 2689 3053
rect 2666 3007 2669 3019
rect 2545 2998 2560 3004
rect 2565 2998 2581 3004
rect 2545 2984 2549 2998
rect 2565 2984 2569 2998
rect 2665 2984 2669 3007
rect 2685 2984 2689 3041
rect 2714 3012 2718 3041
rect 2733 3019 2739 3061
rect 2825 3056 2835 3068
rect 2855 3019 2859 3083
rect 2874 3039 2878 3084
rect 2705 3006 2718 3012
rect 2725 3007 2733 3012
rect 2725 3006 2745 3007
rect 2705 2984 2709 3006
rect 2725 2984 2729 3006
rect 2835 2984 2839 2989
rect 2855 2984 2859 3007
rect 2874 2993 2878 3027
rect 2951 3019 2955 3096
rect 2971 3019 2975 3096
rect 3351 3089 3355 3096
rect 3371 3089 3375 3096
rect 3342 3084 3355 3089
rect 3093 3056 3097 3076
rect 3089 3049 3097 3056
rect 3103 3056 3107 3076
rect 3235 3070 3239 3076
rect 3221 3058 3233 3070
rect 3103 3049 3117 3056
rect 3089 3033 3095 3049
rect 3086 3021 3095 3033
rect 2946 3007 2955 3019
rect 2865 2988 2878 2993
rect 2865 2984 2869 2988
rect 2951 2984 2955 3007
rect 2959 3007 2974 3019
rect 2959 2984 2963 3007
rect 3091 2944 3095 3021
rect 3111 3033 3117 3049
rect 3111 3021 3114 3033
rect 3111 2944 3115 3021
rect 3221 2984 3225 3058
rect 3255 3033 3259 3076
rect 3246 3021 3259 3033
rect 3243 2944 3247 3021
rect 3265 3019 3269 3076
rect 3342 3039 3346 3084
rect 3265 3007 3274 3019
rect 3265 2944 3269 3007
rect 3342 2993 3346 3027
rect 3361 3083 3375 3089
rect 3361 3019 3365 3083
rect 3805 3089 3809 3096
rect 3825 3089 3829 3096
rect 3805 3083 3819 3089
rect 3825 3084 3838 3089
rect 3391 3068 3395 3076
rect 3385 3056 3395 3068
rect 3342 2988 3355 2993
rect 3351 2984 3355 2988
rect 3361 2984 3365 3007
rect 3505 2999 3509 3076
rect 3525 3053 3529 3076
rect 3545 3071 3549 3076
rect 3545 3064 3558 3071
rect 3525 3041 3534 3053
rect 3381 2984 3385 2989
rect 3507 2987 3514 2999
rect 3510 2944 3514 2987
rect 3532 2984 3536 3041
rect 3554 3019 3558 3064
rect 3554 2996 3558 3007
rect 3645 2999 3649 3076
rect 3665 3053 3669 3076
rect 3685 3071 3689 3076
rect 3685 3064 3698 3071
rect 3665 3041 3674 3053
rect 3540 2988 3558 2996
rect 3540 2984 3544 2988
rect 3647 2987 3654 2999
rect 3650 2944 3654 2987
rect 3672 2984 3676 3041
rect 3694 3019 3698 3064
rect 3785 3068 3789 3076
rect 3785 3056 3795 3068
rect 3815 3019 3819 3083
rect 3834 3039 3838 3084
rect 3955 3070 3959 3076
rect 3941 3058 3953 3070
rect 3694 2996 3698 3007
rect 3680 2988 3698 2996
rect 3680 2984 3684 2988
rect 3795 2984 3799 2989
rect 3815 2984 3819 3007
rect 3834 2993 3838 3027
rect 3825 2988 3838 2993
rect 3825 2984 3829 2988
rect 3941 2984 3945 3058
rect 3975 3033 3979 3076
rect 3966 3021 3979 3033
rect 3963 2944 3967 3021
rect 3985 3019 3989 3076
rect 4071 3019 4075 3096
rect 4091 3019 4095 3096
rect 3985 3007 3994 3019
rect 4066 3007 4075 3019
rect 3985 2944 3989 3007
rect 4071 2984 4075 3007
rect 4079 3007 4094 3019
rect 4079 2984 4083 3007
rect 4192 2999 4196 3056
rect 4186 2987 4196 2999
rect 4180 2956 4186 2987
rect 4200 2979 4204 3056
rect 4208 2999 4212 3056
rect 4295 3039 4299 3076
rect 4315 3038 4319 3096
rect 4325 3064 4329 3096
rect 4347 3084 4351 3096
rect 4349 3072 4351 3084
rect 4357 3084 4361 3096
rect 4357 3072 4359 3084
rect 4325 3060 4358 3064
rect 4208 2987 4215 2999
rect 4227 2987 4235 2999
rect 4200 2960 4206 2967
rect 4200 2956 4215 2960
rect 4180 2952 4195 2956
rect 4191 2944 4195 2952
rect 4211 2944 4215 2956
rect 4231 2944 4235 2987
rect 4295 2984 4299 3027
rect 4315 2944 4319 3026
rect 4334 3011 4338 3040
rect 4329 3003 4338 3011
rect 4329 2944 4333 3003
rect 4354 2996 4358 3060
rect 4355 2984 4358 2996
rect 4349 2944 4353 2984
rect 4363 2962 4367 3072
rect 4379 2982 4383 3096
rect 4425 3092 4429 3096
rect 4395 3088 4429 3092
rect 4361 2944 4365 2950
rect 4381 2944 4385 2970
rect 4395 2962 4399 3088
rect 4433 3084 4437 3096
rect 4407 3080 4437 3084
rect 4419 3079 4437 3080
rect 4453 3075 4457 3096
rect 4433 3071 4457 3075
rect 4433 2976 4439 3071
rect 4463 3047 4467 3096
rect 4463 2989 4467 3035
rect 4485 3008 4489 3076
rect 4591 3071 4595 3076
rect 4582 3064 4595 3071
rect 4582 3019 4586 3064
rect 4611 3053 4615 3076
rect 4606 3041 4615 3053
rect 4487 2996 4489 3008
rect 4463 2983 4471 2989
rect 4485 2984 4489 2996
rect 4582 2996 4586 3007
rect 4582 2988 4600 2996
rect 4596 2984 4600 2988
rect 4604 2984 4608 3041
rect 4631 2999 4635 3076
rect 4731 3071 4735 3076
rect 4722 3064 4735 3071
rect 4722 3019 4726 3064
rect 4751 3053 4755 3076
rect 4746 3041 4755 3053
rect 4626 2987 4633 2999
rect 4722 2996 4726 3007
rect 4722 2988 4740 2996
rect 4407 2950 4431 2952
rect 4395 2948 4431 2950
rect 4427 2944 4431 2948
rect 4435 2944 4439 2976
rect 4455 2924 4459 2964
rect 4467 2954 4471 2983
rect 4463 2947 4471 2954
rect 4463 2924 4467 2947
rect 4626 2944 4630 2987
rect 4736 2984 4740 2988
rect 4744 2984 4748 3041
rect 4771 2999 4775 3076
rect 4893 3056 4897 3076
rect 4883 3049 4897 3056
rect 4903 3056 4907 3076
rect 4993 3056 4997 3076
rect 4903 3049 4911 3056
rect 4883 3033 4889 3049
rect 4886 3021 4889 3033
rect 4766 2987 4773 2999
rect 4766 2944 4770 2987
rect 4885 2944 4889 3021
rect 4905 3033 4911 3049
rect 4989 3049 4997 3056
rect 5003 3056 5007 3076
rect 5003 3049 5017 3056
rect 4989 3033 4995 3049
rect 4905 3021 4914 3033
rect 4986 3021 4995 3033
rect 4905 2944 4909 3021
rect 4991 2944 4995 3021
rect 5011 3033 5017 3049
rect 5075 3039 5079 3076
rect 5011 3021 5014 3033
rect 5095 3038 5099 3096
rect 5105 3064 5109 3096
rect 5127 3084 5131 3096
rect 5129 3072 5131 3084
rect 5137 3084 5141 3096
rect 5137 3072 5139 3084
rect 5105 3060 5138 3064
rect 5011 2944 5015 3021
rect 5075 2984 5079 3027
rect 5095 2944 5099 3026
rect 5114 3011 5118 3040
rect 5109 3003 5118 3011
rect 5109 2944 5113 3003
rect 5134 2996 5138 3060
rect 5135 2984 5138 2996
rect 5129 2944 5133 2984
rect 5143 2962 5147 3072
rect 5159 2982 5163 3096
rect 5205 3092 5209 3096
rect 5175 3088 5209 3092
rect 5141 2944 5145 2950
rect 5161 2944 5165 2970
rect 5175 2962 5179 3088
rect 5213 3084 5217 3096
rect 5187 3080 5217 3084
rect 5199 3079 5217 3080
rect 5233 3075 5237 3096
rect 5213 3071 5237 3075
rect 5213 2976 5219 3071
rect 5243 3047 5247 3096
rect 5243 2989 5247 3035
rect 5265 3008 5269 3076
rect 5267 2996 5269 3008
rect 5243 2983 5251 2989
rect 5265 2984 5269 2996
rect 5365 3056 5369 3076
rect 5385 3056 5389 3076
rect 5405 3056 5409 3076
rect 5425 3056 5429 3076
rect 5445 3056 5449 3076
rect 5465 3056 5469 3076
rect 5365 3044 5378 3056
rect 5405 3044 5418 3056
rect 5445 3044 5458 3056
rect 5485 3053 5489 3076
rect 5505 3053 5509 3076
rect 5365 2984 5369 3044
rect 5385 2984 5389 3044
rect 5405 2984 5409 3044
rect 5425 2984 5429 3044
rect 5445 2984 5449 3044
rect 5465 2984 5469 3044
rect 5485 3041 5494 3053
rect 5506 3041 5509 3053
rect 5485 2984 5489 3041
rect 5505 2984 5509 3041
rect 5551 3008 5555 3076
rect 5573 3047 5577 3096
rect 5583 3075 5587 3096
rect 5603 3084 5607 3096
rect 5611 3092 5615 3096
rect 5611 3088 5645 3092
rect 5603 3080 5633 3084
rect 5603 3079 5621 3080
rect 5583 3071 5607 3075
rect 5551 2996 5553 3008
rect 5551 2984 5555 2996
rect 5573 2989 5577 3035
rect 5187 2950 5211 2952
rect 5175 2948 5211 2950
rect 5207 2944 5211 2948
rect 5215 2944 5219 2976
rect 5235 2924 5239 2964
rect 5247 2954 5251 2983
rect 5243 2947 5251 2954
rect 5243 2924 5247 2947
rect 5569 2983 5577 2989
rect 5569 2954 5573 2983
rect 5601 2976 5607 3071
rect 5569 2947 5577 2954
rect 5573 2924 5577 2947
rect 5581 2924 5585 2964
rect 5601 2944 5605 2976
rect 5641 2962 5645 3088
rect 5657 2982 5661 3096
rect 5679 3084 5683 3096
rect 5681 3072 5683 3084
rect 5689 3084 5693 3096
rect 5689 3072 5691 3084
rect 5609 2950 5633 2952
rect 5609 2948 5645 2950
rect 5609 2944 5613 2948
rect 5655 2944 5659 2970
rect 5673 2962 5677 3072
rect 5711 3064 5715 3096
rect 5682 3060 5715 3064
rect 5682 2996 5686 3060
rect 5702 3011 5706 3040
rect 5721 3038 5725 3096
rect 5741 3039 5745 3076
rect 5702 3003 5711 3011
rect 5682 2984 5685 2996
rect 5675 2944 5679 2950
rect 5687 2944 5691 2984
rect 5707 2944 5711 3003
rect 5721 2944 5725 3026
rect 5741 2984 5745 3027
rect 101 2900 105 2904
rect 123 2900 127 2904
rect 145 2900 149 2904
rect 251 2900 255 2904
rect 271 2900 275 2904
rect 291 2900 295 2904
rect 391 2900 395 2904
rect 411 2900 415 2904
rect 530 2900 534 2904
rect 552 2900 556 2904
rect 560 2900 564 2904
rect 656 2900 660 2904
rect 664 2900 668 2904
rect 686 2900 690 2904
rect 796 2900 800 2904
rect 804 2900 808 2904
rect 826 2900 830 2904
rect 936 2900 940 2904
rect 944 2900 948 2904
rect 966 2900 970 2904
rect 1085 2900 1089 2904
rect 1105 2900 1109 2904
rect 1237 2900 1241 2904
rect 1245 2900 1249 2904
rect 1336 2900 1340 2904
rect 1344 2900 1348 2904
rect 1366 2900 1370 2904
rect 1485 2900 1489 2904
rect 1505 2900 1509 2904
rect 1525 2900 1529 2904
rect 1645 2900 1649 2904
rect 1665 2900 1669 2904
rect 1685 2900 1689 2904
rect 1790 2900 1794 2904
rect 1812 2900 1816 2904
rect 1820 2900 1824 2904
rect 1916 2900 1920 2904
rect 1924 2900 1928 2904
rect 1946 2900 1950 2904
rect 2090 2900 2094 2904
rect 2112 2900 2116 2904
rect 2120 2900 2124 2904
rect 2230 2900 2234 2904
rect 2252 2900 2256 2904
rect 2260 2900 2264 2904
rect 2385 2900 2389 2904
rect 2405 2900 2409 2904
rect 2425 2900 2429 2904
rect 2525 2900 2529 2904
rect 2545 2900 2549 2904
rect 2565 2900 2569 2904
rect 2665 2900 2669 2904
rect 2685 2900 2689 2904
rect 2705 2900 2709 2904
rect 2725 2900 2729 2904
rect 2835 2900 2839 2904
rect 2855 2900 2859 2904
rect 2865 2900 2869 2904
rect 2951 2900 2955 2904
rect 2959 2900 2963 2904
rect 3091 2900 3095 2904
rect 3111 2900 3115 2904
rect 3221 2900 3225 2904
rect 3243 2900 3247 2904
rect 3265 2900 3269 2904
rect 3351 2900 3355 2904
rect 3361 2900 3365 2904
rect 3381 2900 3385 2904
rect 3510 2900 3514 2904
rect 3532 2900 3536 2904
rect 3540 2900 3544 2904
rect 3650 2900 3654 2904
rect 3672 2900 3676 2904
rect 3680 2900 3684 2904
rect 3795 2900 3799 2904
rect 3815 2900 3819 2904
rect 3825 2900 3829 2904
rect 3941 2900 3945 2904
rect 3963 2900 3967 2904
rect 3985 2900 3989 2904
rect 4071 2900 4075 2904
rect 4079 2900 4083 2904
rect 4191 2900 4195 2904
rect 4211 2900 4215 2904
rect 4231 2900 4235 2904
rect 4295 2900 4299 2904
rect 4315 2900 4319 2904
rect 4329 2900 4333 2904
rect 4349 2900 4353 2904
rect 4361 2900 4365 2904
rect 4381 2900 4385 2904
rect 4427 2900 4431 2904
rect 4435 2900 4439 2904
rect 4455 2900 4459 2904
rect 4463 2900 4467 2904
rect 4485 2900 4489 2904
rect 4596 2900 4600 2904
rect 4604 2900 4608 2904
rect 4626 2900 4630 2904
rect 4736 2900 4740 2904
rect 4744 2900 4748 2904
rect 4766 2900 4770 2904
rect 4885 2900 4889 2904
rect 4905 2900 4909 2904
rect 4991 2900 4995 2904
rect 5011 2900 5015 2904
rect 5075 2900 5079 2904
rect 5095 2900 5099 2904
rect 5109 2900 5113 2904
rect 5129 2900 5133 2904
rect 5141 2900 5145 2904
rect 5161 2900 5165 2904
rect 5207 2900 5211 2904
rect 5215 2900 5219 2904
rect 5235 2900 5239 2904
rect 5243 2900 5247 2904
rect 5265 2900 5269 2904
rect 5365 2900 5369 2904
rect 5385 2900 5389 2904
rect 5405 2900 5409 2904
rect 5425 2900 5429 2904
rect 5445 2900 5449 2904
rect 5465 2900 5469 2904
rect 5485 2900 5489 2904
rect 5505 2900 5509 2904
rect 5551 2900 5555 2904
rect 5573 2900 5577 2904
rect 5581 2900 5585 2904
rect 5601 2900 5605 2904
rect 5609 2900 5613 2904
rect 5655 2900 5659 2904
rect 5675 2900 5679 2904
rect 5687 2900 5691 2904
rect 5707 2900 5711 2904
rect 5721 2900 5725 2904
rect 5741 2900 5745 2904
rect 85 2876 89 2880
rect 105 2876 109 2880
rect 196 2876 200 2880
rect 204 2876 208 2880
rect 226 2876 230 2880
rect 345 2876 349 2880
rect 431 2876 435 2880
rect 451 2876 455 2880
rect 471 2876 475 2880
rect 585 2876 589 2880
rect 605 2876 609 2880
rect 691 2876 695 2880
rect 713 2876 717 2880
rect 735 2876 739 2880
rect 831 2876 835 2880
rect 851 2876 855 2880
rect 951 2876 955 2880
rect 971 2876 975 2880
rect 991 2876 995 2880
rect 1091 2876 1095 2880
rect 1111 2876 1115 2880
rect 1250 2876 1254 2880
rect 1272 2876 1276 2880
rect 1280 2876 1284 2880
rect 1376 2876 1380 2880
rect 1384 2876 1388 2880
rect 1406 2876 1410 2880
rect 1535 2876 1539 2880
rect 1555 2876 1559 2880
rect 1565 2876 1569 2880
rect 1651 2876 1655 2880
rect 1659 2876 1663 2880
rect 1781 2876 1785 2880
rect 1803 2876 1807 2880
rect 1825 2876 1829 2880
rect 1945 2876 1949 2880
rect 1965 2876 1969 2880
rect 2056 2876 2060 2880
rect 2064 2876 2068 2880
rect 2086 2876 2090 2880
rect 2201 2876 2205 2880
rect 2223 2876 2227 2880
rect 2245 2876 2249 2880
rect 2345 2876 2349 2880
rect 2365 2876 2369 2880
rect 2471 2876 2475 2880
rect 2479 2876 2483 2880
rect 2605 2876 2609 2880
rect 2625 2876 2629 2880
rect 2645 2876 2649 2880
rect 2741 2876 2745 2880
rect 2763 2876 2767 2880
rect 2785 2876 2789 2880
rect 2896 2876 2900 2880
rect 2904 2876 2908 2880
rect 2926 2876 2930 2880
rect 3045 2876 3049 2880
rect 3065 2876 3069 2880
rect 3085 2876 3089 2880
rect 3171 2876 3175 2880
rect 3191 2876 3195 2880
rect 3310 2876 3314 2880
rect 3332 2876 3336 2880
rect 3340 2876 3344 2880
rect 3441 2876 3445 2880
rect 3463 2876 3467 2880
rect 3485 2876 3489 2880
rect 3571 2876 3575 2880
rect 3579 2876 3583 2880
rect 3691 2876 3695 2880
rect 3711 2876 3715 2880
rect 3731 2876 3735 2880
rect 3831 2876 3835 2880
rect 3851 2876 3855 2880
rect 3965 2876 3969 2880
rect 4070 2876 4074 2880
rect 4092 2876 4096 2880
rect 4100 2876 4104 2880
rect 4191 2876 4195 2880
rect 4211 2876 4215 2880
rect 4311 2876 4315 2880
rect 4411 2876 4415 2880
rect 4471 2876 4475 2880
rect 4493 2876 4497 2880
rect 4501 2876 4505 2880
rect 4521 2876 4525 2880
rect 4529 2876 4533 2880
rect 4575 2876 4579 2880
rect 4595 2876 4599 2880
rect 4607 2876 4611 2880
rect 4627 2876 4631 2880
rect 4641 2876 4645 2880
rect 4661 2876 4665 2880
rect 4715 2876 4719 2880
rect 4735 2876 4739 2880
rect 4749 2876 4753 2880
rect 4769 2876 4773 2880
rect 4781 2876 4785 2880
rect 4801 2876 4805 2880
rect 4847 2876 4851 2880
rect 4855 2876 4859 2880
rect 4875 2876 4879 2880
rect 4883 2876 4887 2880
rect 4905 2876 4909 2880
rect 5016 2876 5020 2880
rect 5024 2876 5028 2880
rect 5046 2876 5050 2880
rect 5151 2876 5155 2880
rect 5171 2876 5175 2880
rect 5271 2876 5275 2880
rect 5291 2876 5295 2880
rect 5351 2876 5355 2880
rect 5373 2876 5377 2880
rect 5381 2876 5385 2880
rect 5401 2876 5405 2880
rect 5409 2876 5413 2880
rect 5455 2876 5459 2880
rect 5475 2876 5479 2880
rect 5487 2876 5491 2880
rect 5507 2876 5511 2880
rect 5521 2876 5525 2880
rect 5541 2876 5545 2880
rect 5636 2876 5640 2880
rect 5644 2876 5648 2880
rect 5666 2876 5670 2880
rect 85 2759 89 2836
rect 86 2747 89 2759
rect 83 2731 89 2747
rect 105 2759 109 2836
rect 196 2792 200 2796
rect 182 2784 200 2792
rect 182 2773 186 2784
rect 105 2747 114 2759
rect 105 2731 111 2747
rect 83 2724 97 2731
rect 93 2704 97 2724
rect 103 2724 111 2731
rect 103 2704 107 2724
rect 182 2716 186 2761
rect 204 2739 208 2796
rect 226 2793 230 2836
rect 226 2781 233 2793
rect 206 2727 215 2739
rect 182 2709 195 2716
rect 191 2704 195 2709
rect 211 2704 215 2727
rect 231 2704 235 2781
rect 345 2753 349 2836
rect 431 2782 435 2796
rect 451 2782 455 2796
rect 419 2776 435 2782
rect 440 2776 455 2782
rect 345 2741 354 2753
rect 345 2684 349 2741
rect 419 2739 426 2776
rect 440 2753 446 2776
rect 419 2714 426 2727
rect 419 2708 438 2714
rect 434 2704 438 2708
rect 442 2704 446 2741
rect 471 2739 475 2796
rect 585 2759 589 2836
rect 586 2747 589 2759
rect 466 2727 475 2739
rect 583 2731 589 2747
rect 605 2759 609 2836
rect 691 2773 695 2836
rect 686 2761 695 2773
rect 605 2747 614 2759
rect 605 2731 611 2747
rect 464 2684 468 2727
rect 583 2724 597 2731
rect 593 2704 597 2724
rect 603 2724 611 2731
rect 603 2704 607 2724
rect 691 2704 695 2761
rect 713 2759 717 2836
rect 701 2747 714 2759
rect 701 2704 705 2747
rect 735 2722 739 2796
rect 831 2759 835 2836
rect 826 2747 835 2759
rect 829 2731 835 2747
rect 851 2759 855 2836
rect 951 2782 955 2796
rect 971 2782 975 2796
rect 939 2776 955 2782
rect 960 2776 975 2782
rect 851 2747 854 2759
rect 851 2731 857 2747
rect 939 2739 946 2776
rect 960 2753 966 2776
rect 829 2724 837 2731
rect 727 2710 739 2722
rect 721 2704 725 2710
rect 833 2704 837 2724
rect 843 2724 857 2731
rect 843 2704 847 2724
rect 939 2714 946 2727
rect 939 2708 958 2714
rect 954 2704 958 2708
rect 962 2704 966 2741
rect 991 2739 995 2796
rect 1091 2759 1095 2836
rect 1086 2747 1095 2759
rect 986 2727 995 2739
rect 1089 2731 1095 2747
rect 1111 2759 1115 2836
rect 1250 2793 1254 2836
rect 1247 2781 1254 2793
rect 1111 2747 1114 2759
rect 1111 2731 1117 2747
rect 984 2684 988 2727
rect 1089 2724 1097 2731
rect 1093 2704 1097 2724
rect 1103 2724 1117 2731
rect 1103 2704 1107 2724
rect 1245 2704 1249 2781
rect 1272 2739 1276 2796
rect 1280 2792 1284 2796
rect 1376 2792 1380 2796
rect 1280 2784 1298 2792
rect 1294 2773 1298 2784
rect 1362 2784 1380 2792
rect 1362 2773 1366 2784
rect 1265 2727 1274 2739
rect 1265 2704 1269 2727
rect 1294 2716 1298 2761
rect 1285 2709 1298 2716
rect 1362 2716 1366 2761
rect 1384 2739 1388 2796
rect 1406 2793 1410 2836
rect 1406 2781 1413 2793
rect 1535 2791 1539 2796
rect 1386 2727 1395 2739
rect 1362 2709 1375 2716
rect 1285 2704 1289 2709
rect 1371 2704 1375 2709
rect 1391 2704 1395 2727
rect 1411 2704 1415 2781
rect 1555 2773 1559 2796
rect 1565 2792 1569 2796
rect 1565 2787 1578 2792
rect 1525 2712 1535 2724
rect 1525 2704 1529 2712
rect 1555 2697 1559 2761
rect 1545 2691 1559 2697
rect 1574 2753 1578 2787
rect 1651 2773 1655 2796
rect 1646 2761 1655 2773
rect 1659 2773 1663 2796
rect 1659 2761 1674 2773
rect 1574 2696 1578 2741
rect 1565 2691 1578 2696
rect 1545 2684 1549 2691
rect 1565 2684 1569 2691
rect 1651 2684 1655 2761
rect 1671 2684 1675 2761
rect 1781 2722 1785 2796
rect 1803 2759 1807 2836
rect 1825 2773 1829 2836
rect 1825 2761 1834 2773
rect 1806 2747 1819 2759
rect 1781 2710 1793 2722
rect 1795 2704 1799 2710
rect 1815 2704 1819 2747
rect 1825 2704 1829 2761
rect 1945 2759 1949 2836
rect 1946 2747 1949 2759
rect 1943 2731 1949 2747
rect 1965 2759 1969 2836
rect 2056 2792 2060 2796
rect 2042 2784 2060 2792
rect 2042 2773 2046 2784
rect 1965 2747 1974 2759
rect 1965 2731 1971 2747
rect 1943 2724 1957 2731
rect 1953 2704 1957 2724
rect 1963 2724 1971 2731
rect 1963 2704 1967 2724
rect 2042 2716 2046 2761
rect 2064 2739 2068 2796
rect 2086 2793 2090 2836
rect 2086 2781 2093 2793
rect 2066 2727 2075 2739
rect 2042 2709 2055 2716
rect 2051 2704 2055 2709
rect 2071 2704 2075 2727
rect 2091 2704 2095 2781
rect 2201 2722 2205 2796
rect 2223 2759 2227 2836
rect 2245 2773 2249 2836
rect 2245 2761 2254 2773
rect 2226 2747 2239 2759
rect 2201 2710 2213 2722
rect 2215 2704 2219 2710
rect 2235 2704 2239 2747
rect 2245 2704 2249 2761
rect 2345 2759 2349 2836
rect 2346 2747 2349 2759
rect 2343 2731 2349 2747
rect 2365 2759 2369 2836
rect 2471 2773 2475 2796
rect 2466 2761 2475 2773
rect 2479 2773 2483 2796
rect 2605 2793 2609 2836
rect 2625 2824 2629 2836
rect 2645 2828 2649 2836
rect 2645 2824 2660 2828
rect 2625 2820 2640 2824
rect 2634 2813 2640 2820
rect 2605 2781 2613 2793
rect 2625 2781 2632 2793
rect 2479 2761 2494 2773
rect 2365 2747 2374 2759
rect 2365 2731 2371 2747
rect 2343 2724 2357 2731
rect 2353 2704 2357 2724
rect 2363 2724 2371 2731
rect 2363 2704 2367 2724
rect 2471 2684 2475 2761
rect 2491 2684 2495 2761
rect 2628 2724 2632 2781
rect 2636 2724 2640 2801
rect 2654 2793 2660 2824
rect 2644 2781 2654 2793
rect 2644 2724 2648 2781
rect 2741 2722 2745 2796
rect 2763 2759 2767 2836
rect 2785 2773 2789 2836
rect 2896 2792 2900 2796
rect 2882 2784 2900 2792
rect 2882 2773 2886 2784
rect 2785 2761 2794 2773
rect 2766 2747 2779 2759
rect 2741 2710 2753 2722
rect 2755 2704 2759 2710
rect 2775 2704 2779 2747
rect 2785 2704 2789 2761
rect 2882 2716 2886 2761
rect 2904 2739 2908 2796
rect 2926 2793 2930 2836
rect 3045 2793 3049 2836
rect 3065 2824 3069 2836
rect 3085 2828 3089 2836
rect 3085 2824 3100 2828
rect 3065 2820 3080 2824
rect 3074 2813 3080 2820
rect 2926 2781 2933 2793
rect 3045 2781 3053 2793
rect 3065 2781 3072 2793
rect 2906 2727 2915 2739
rect 2882 2709 2895 2716
rect 2891 2704 2895 2709
rect 2911 2704 2915 2727
rect 2931 2704 2935 2781
rect 3068 2724 3072 2781
rect 3076 2724 3080 2801
rect 3094 2793 3100 2824
rect 3084 2781 3094 2793
rect 3084 2724 3088 2781
rect 3171 2759 3175 2836
rect 3166 2747 3175 2759
rect 3169 2731 3175 2747
rect 3191 2759 3195 2836
rect 3310 2793 3314 2836
rect 3307 2781 3314 2793
rect 3191 2747 3194 2759
rect 3191 2731 3197 2747
rect 3169 2724 3177 2731
rect 3173 2704 3177 2724
rect 3183 2724 3197 2731
rect 3183 2704 3187 2724
rect 3305 2704 3309 2781
rect 3332 2739 3336 2796
rect 3340 2792 3344 2796
rect 3340 2784 3358 2792
rect 3354 2773 3358 2784
rect 3325 2727 3334 2739
rect 3325 2704 3329 2727
rect 3354 2716 3358 2761
rect 3345 2709 3358 2716
rect 3441 2722 3445 2796
rect 3463 2759 3467 2836
rect 3485 2773 3489 2836
rect 3691 2828 3695 2836
rect 3680 2824 3695 2828
rect 3711 2824 3715 2836
rect 3571 2773 3575 2796
rect 3485 2761 3494 2773
rect 3566 2761 3575 2773
rect 3579 2773 3583 2796
rect 3680 2793 3686 2824
rect 3700 2820 3715 2824
rect 3700 2813 3706 2820
rect 3686 2781 3696 2793
rect 3579 2761 3594 2773
rect 3466 2747 3479 2759
rect 3441 2710 3453 2722
rect 3345 2704 3349 2709
rect 3455 2704 3459 2710
rect 3475 2704 3479 2747
rect 3485 2704 3489 2761
rect 3571 2684 3575 2761
rect 3591 2684 3595 2761
rect 3692 2724 3696 2781
rect 3700 2724 3704 2801
rect 3731 2793 3735 2836
rect 3708 2781 3715 2793
rect 3727 2781 3735 2793
rect 3708 2724 3712 2781
rect 3831 2759 3835 2836
rect 3826 2747 3835 2759
rect 3829 2731 3835 2747
rect 3851 2759 3855 2836
rect 3851 2747 3854 2759
rect 3851 2731 3857 2747
rect 3829 2724 3837 2731
rect 3833 2704 3837 2724
rect 3843 2724 3857 2731
rect 3965 2739 3969 2796
rect 4070 2793 4074 2836
rect 4067 2781 4074 2793
rect 3965 2727 3974 2739
rect 3843 2704 3847 2724
rect 3965 2704 3969 2727
rect 4065 2704 4069 2781
rect 4092 2739 4096 2796
rect 4100 2792 4104 2796
rect 4100 2784 4118 2792
rect 4114 2773 4118 2784
rect 4085 2727 4094 2739
rect 4085 2704 4089 2727
rect 4114 2716 4118 2761
rect 4191 2759 4195 2836
rect 4186 2747 4195 2759
rect 4189 2731 4195 2747
rect 4211 2759 4215 2836
rect 4211 2747 4214 2759
rect 4211 2731 4217 2747
rect 4311 2739 4315 2796
rect 4411 2753 4415 2836
rect 4493 2833 4497 2856
rect 4489 2826 4497 2833
rect 4489 2797 4493 2826
rect 4501 2816 4505 2856
rect 4521 2804 4525 2836
rect 4529 2832 4533 2836
rect 4529 2830 4565 2832
rect 4529 2828 4553 2830
rect 4406 2741 4415 2753
rect 4189 2724 4197 2731
rect 4105 2709 4118 2716
rect 4105 2704 4109 2709
rect 4193 2704 4197 2724
rect 4203 2724 4217 2731
rect 4306 2727 4315 2739
rect 4203 2704 4207 2724
rect 4311 2704 4315 2727
rect 4411 2684 4415 2741
rect 4471 2784 4475 2796
rect 4489 2791 4497 2797
rect 4471 2772 4473 2784
rect 4471 2704 4475 2772
rect 4493 2745 4497 2791
rect 4493 2684 4497 2733
rect 4521 2709 4527 2804
rect 4503 2705 4527 2709
rect 4503 2684 4507 2705
rect 4523 2700 4541 2701
rect 4523 2696 4553 2700
rect 4523 2684 4527 2696
rect 4561 2692 4565 2818
rect 4575 2810 4579 2836
rect 4595 2830 4599 2836
rect 4531 2688 4565 2692
rect 4531 2684 4535 2688
rect 4577 2684 4581 2798
rect 4593 2708 4597 2818
rect 4607 2796 4611 2836
rect 4602 2784 4605 2796
rect 4602 2720 4606 2784
rect 4627 2777 4631 2836
rect 4622 2769 4631 2777
rect 4622 2740 4626 2769
rect 4641 2754 4645 2836
rect 4661 2753 4665 2796
rect 4715 2753 4719 2796
rect 4735 2754 4739 2836
rect 4749 2777 4753 2836
rect 4769 2796 4773 2836
rect 4781 2830 4785 2836
rect 4775 2784 4778 2796
rect 4749 2769 4758 2777
rect 4602 2716 4635 2720
rect 4601 2696 4603 2708
rect 4599 2684 4603 2696
rect 4609 2696 4611 2708
rect 4609 2684 4613 2696
rect 4631 2684 4635 2716
rect 4641 2684 4645 2742
rect 4661 2704 4665 2741
rect 4715 2704 4719 2741
rect 4735 2684 4739 2742
rect 4754 2740 4758 2769
rect 4774 2720 4778 2784
rect 4745 2716 4778 2720
rect 4745 2684 4749 2716
rect 4783 2708 4787 2818
rect 4801 2810 4805 2836
rect 4847 2832 4851 2836
rect 4815 2830 4851 2832
rect 4827 2828 4851 2830
rect 4769 2696 4771 2708
rect 4767 2684 4771 2696
rect 4777 2696 4779 2708
rect 4777 2684 4781 2696
rect 4799 2684 4803 2798
rect 4815 2692 4819 2818
rect 4855 2804 4859 2836
rect 4875 2816 4879 2856
rect 4883 2833 4887 2856
rect 4883 2826 4891 2833
rect 4853 2709 4859 2804
rect 4887 2797 4891 2826
rect 4883 2791 4891 2797
rect 4883 2745 4887 2791
rect 4905 2784 4909 2796
rect 5016 2792 5020 2796
rect 4907 2772 4909 2784
rect 5002 2784 5020 2792
rect 5002 2773 5006 2784
rect 4853 2705 4877 2709
rect 4839 2700 4857 2701
rect 4827 2696 4857 2700
rect 4815 2688 4849 2692
rect 4845 2684 4849 2688
rect 4853 2684 4857 2696
rect 4873 2684 4877 2705
rect 4883 2684 4887 2733
rect 4905 2704 4909 2772
rect 5002 2716 5006 2761
rect 5024 2739 5028 2796
rect 5046 2793 5050 2836
rect 5046 2781 5053 2793
rect 5026 2727 5035 2739
rect 5002 2709 5015 2716
rect 5011 2704 5015 2709
rect 5031 2704 5035 2727
rect 5051 2704 5055 2781
rect 5151 2759 5155 2836
rect 5146 2747 5155 2759
rect 5149 2731 5155 2747
rect 5171 2759 5175 2836
rect 5373 2833 5377 2856
rect 5369 2826 5377 2833
rect 5369 2797 5373 2826
rect 5381 2816 5385 2856
rect 5401 2804 5405 2836
rect 5409 2832 5413 2836
rect 5409 2830 5445 2832
rect 5409 2828 5433 2830
rect 5271 2792 5275 2796
rect 5291 2792 5295 2796
rect 5271 2788 5295 2792
rect 5171 2747 5174 2759
rect 5171 2731 5177 2747
rect 5271 2739 5275 2788
rect 5149 2724 5157 2731
rect 5153 2704 5157 2724
rect 5163 2724 5177 2731
rect 5266 2727 5275 2739
rect 5163 2704 5167 2724
rect 5271 2712 5275 2727
rect 5351 2784 5355 2796
rect 5369 2791 5377 2797
rect 5351 2772 5353 2784
rect 5271 2708 5295 2712
rect 5271 2704 5275 2708
rect 5291 2704 5295 2708
rect 5351 2704 5355 2772
rect 5373 2745 5377 2791
rect 5373 2684 5377 2733
rect 5401 2709 5407 2804
rect 5383 2705 5407 2709
rect 5383 2684 5387 2705
rect 5403 2700 5421 2701
rect 5403 2696 5433 2700
rect 5403 2684 5407 2696
rect 5441 2692 5445 2818
rect 5455 2810 5459 2836
rect 5475 2830 5479 2836
rect 5411 2688 5445 2692
rect 5411 2684 5415 2688
rect 5457 2684 5461 2798
rect 5473 2708 5477 2818
rect 5487 2796 5491 2836
rect 5482 2784 5485 2796
rect 5482 2720 5486 2784
rect 5507 2777 5511 2836
rect 5502 2769 5511 2777
rect 5502 2740 5506 2769
rect 5521 2754 5525 2836
rect 5541 2753 5545 2796
rect 5636 2792 5640 2796
rect 5622 2784 5640 2792
rect 5622 2773 5626 2784
rect 5482 2716 5515 2720
rect 5481 2696 5483 2708
rect 5479 2684 5483 2696
rect 5489 2696 5491 2708
rect 5489 2684 5493 2696
rect 5511 2684 5515 2716
rect 5521 2684 5525 2742
rect 5541 2704 5545 2741
rect 5622 2716 5626 2761
rect 5644 2739 5648 2796
rect 5666 2793 5670 2836
rect 5666 2781 5673 2793
rect 5646 2727 5655 2739
rect 5622 2709 5635 2716
rect 5631 2704 5635 2709
rect 5651 2704 5655 2727
rect 5671 2704 5675 2781
rect 93 2660 97 2664
rect 103 2660 107 2664
rect 191 2660 195 2664
rect 211 2660 215 2664
rect 231 2660 235 2664
rect 345 2660 349 2664
rect 434 2660 438 2664
rect 442 2660 446 2664
rect 464 2660 468 2664
rect 593 2660 597 2664
rect 603 2660 607 2664
rect 691 2660 695 2664
rect 701 2660 705 2664
rect 721 2660 725 2664
rect 833 2660 837 2664
rect 843 2660 847 2664
rect 954 2660 958 2664
rect 962 2660 966 2664
rect 984 2660 988 2664
rect 1093 2660 1097 2664
rect 1103 2660 1107 2664
rect 1245 2660 1249 2664
rect 1265 2660 1269 2664
rect 1285 2660 1289 2664
rect 1371 2660 1375 2664
rect 1391 2660 1395 2664
rect 1411 2660 1415 2664
rect 1525 2660 1529 2664
rect 1545 2660 1549 2664
rect 1565 2660 1569 2664
rect 1651 2660 1655 2664
rect 1671 2660 1675 2664
rect 1795 2660 1799 2664
rect 1815 2660 1819 2664
rect 1825 2660 1829 2664
rect 1953 2660 1957 2664
rect 1963 2660 1967 2664
rect 2051 2660 2055 2664
rect 2071 2660 2075 2664
rect 2091 2660 2095 2664
rect 2215 2660 2219 2664
rect 2235 2660 2239 2664
rect 2245 2660 2249 2664
rect 2353 2660 2357 2664
rect 2363 2660 2367 2664
rect 2471 2660 2475 2664
rect 2491 2660 2495 2664
rect 2628 2660 2632 2664
rect 2636 2660 2640 2664
rect 2644 2660 2648 2664
rect 2755 2660 2759 2664
rect 2775 2660 2779 2664
rect 2785 2660 2789 2664
rect 2891 2660 2895 2664
rect 2911 2660 2915 2664
rect 2931 2660 2935 2664
rect 3068 2660 3072 2664
rect 3076 2660 3080 2664
rect 3084 2660 3088 2664
rect 3173 2660 3177 2664
rect 3183 2660 3187 2664
rect 3305 2660 3309 2664
rect 3325 2660 3329 2664
rect 3345 2660 3349 2664
rect 3455 2660 3459 2664
rect 3475 2660 3479 2664
rect 3485 2660 3489 2664
rect 3571 2660 3575 2664
rect 3591 2660 3595 2664
rect 3692 2660 3696 2664
rect 3700 2660 3704 2664
rect 3708 2660 3712 2664
rect 3833 2660 3837 2664
rect 3843 2660 3847 2664
rect 3965 2660 3969 2664
rect 4065 2660 4069 2664
rect 4085 2660 4089 2664
rect 4105 2660 4109 2664
rect 4193 2660 4197 2664
rect 4203 2660 4207 2664
rect 4311 2660 4315 2664
rect 4411 2660 4415 2664
rect 4471 2660 4475 2664
rect 4493 2660 4497 2664
rect 4503 2660 4507 2664
rect 4523 2660 4527 2664
rect 4531 2660 4535 2664
rect 4577 2660 4581 2664
rect 4599 2660 4603 2664
rect 4609 2660 4613 2664
rect 4631 2660 4635 2664
rect 4641 2660 4645 2664
rect 4661 2660 4665 2664
rect 4715 2660 4719 2664
rect 4735 2660 4739 2664
rect 4745 2660 4749 2664
rect 4767 2660 4771 2664
rect 4777 2660 4781 2664
rect 4799 2660 4803 2664
rect 4845 2660 4849 2664
rect 4853 2660 4857 2664
rect 4873 2660 4877 2664
rect 4883 2660 4887 2664
rect 4905 2660 4909 2664
rect 5011 2660 5015 2664
rect 5031 2660 5035 2664
rect 5051 2660 5055 2664
rect 5153 2660 5157 2664
rect 5163 2660 5167 2664
rect 5271 2660 5275 2664
rect 5291 2660 5295 2664
rect 5351 2660 5355 2664
rect 5373 2660 5377 2664
rect 5383 2660 5387 2664
rect 5403 2660 5407 2664
rect 5411 2660 5415 2664
rect 5457 2660 5461 2664
rect 5479 2660 5483 2664
rect 5489 2660 5493 2664
rect 5511 2660 5515 2664
rect 5521 2660 5525 2664
rect 5541 2660 5545 2664
rect 5631 2660 5635 2664
rect 5651 2660 5655 2664
rect 5671 2660 5675 2664
rect 85 2636 89 2640
rect 171 2636 175 2640
rect 292 2636 296 2640
rect 314 2636 318 2640
rect 322 2636 326 2640
rect 412 2636 416 2640
rect 420 2636 424 2640
rect 428 2636 432 2640
rect 551 2636 555 2640
rect 651 2636 655 2640
rect 671 2636 675 2640
rect 771 2636 775 2640
rect 791 2636 795 2640
rect 811 2636 815 2640
rect 934 2636 938 2640
rect 942 2636 946 2640
rect 964 2636 968 2640
rect 1085 2636 1089 2640
rect 1105 2636 1109 2640
rect 1125 2636 1129 2640
rect 1233 2636 1237 2640
rect 1243 2636 1247 2640
rect 1331 2636 1335 2640
rect 1341 2636 1345 2640
rect 1361 2636 1365 2640
rect 1508 2636 1512 2640
rect 1516 2636 1520 2640
rect 1524 2636 1528 2640
rect 1611 2636 1615 2640
rect 1711 2636 1715 2640
rect 1731 2636 1735 2640
rect 1751 2636 1755 2640
rect 1865 2636 1869 2640
rect 1885 2636 1889 2640
rect 1905 2636 1909 2640
rect 1991 2636 1995 2640
rect 2011 2636 2015 2640
rect 2031 2636 2035 2640
rect 2168 2636 2172 2640
rect 2176 2636 2180 2640
rect 2184 2636 2188 2640
rect 2292 2636 2296 2640
rect 2314 2636 2318 2640
rect 2322 2636 2326 2640
rect 2413 2636 2417 2640
rect 2423 2636 2427 2640
rect 2565 2636 2569 2640
rect 2585 2636 2589 2640
rect 2605 2636 2609 2640
rect 2691 2636 2695 2640
rect 2711 2636 2715 2640
rect 2731 2636 2735 2640
rect 2852 2636 2856 2640
rect 2874 2636 2878 2640
rect 2882 2636 2886 2640
rect 2985 2636 2989 2640
rect 3071 2636 3075 2640
rect 3091 2636 3095 2640
rect 3111 2636 3115 2640
rect 3233 2636 3237 2640
rect 3243 2636 3247 2640
rect 3388 2636 3392 2640
rect 3396 2636 3400 2640
rect 3404 2636 3408 2640
rect 3491 2636 3495 2640
rect 3501 2636 3505 2640
rect 3521 2636 3525 2640
rect 3633 2636 3637 2640
rect 3643 2636 3647 2640
rect 3754 2636 3758 2640
rect 3762 2636 3766 2640
rect 3782 2636 3786 2640
rect 3790 2636 3794 2640
rect 3911 2636 3915 2640
rect 3931 2636 3935 2640
rect 3999 2636 4003 2640
rect 4047 2636 4051 2640
rect 4059 2636 4063 2640
rect 4084 2636 4088 2640
rect 4096 2636 4100 2640
rect 4149 2636 4153 2640
rect 4169 2636 4173 2640
rect 4214 2636 4218 2640
rect 4234 2636 4238 2640
rect 4284 2636 4288 2640
rect 4304 2636 4308 2640
rect 4324 2636 4328 2640
rect 4374 2636 4378 2640
rect 4386 2636 4390 2640
rect 4410 2636 4414 2640
rect 4422 2636 4426 2640
rect 4474 2636 4478 2640
rect 4486 2636 4490 2640
rect 4510 2636 4514 2640
rect 4522 2636 4526 2640
rect 4572 2636 4576 2640
rect 4592 2636 4596 2640
rect 4612 2636 4616 2640
rect 4662 2636 4666 2640
rect 4682 2636 4686 2640
rect 4727 2636 4731 2640
rect 4747 2636 4751 2640
rect 4800 2636 4804 2640
rect 4812 2636 4816 2640
rect 4837 2636 4841 2640
rect 4849 2636 4853 2640
rect 4897 2636 4901 2640
rect 4955 2636 4959 2640
rect 4975 2636 4979 2640
rect 4985 2636 4989 2640
rect 5007 2636 5011 2640
rect 5017 2636 5021 2640
rect 5039 2636 5043 2640
rect 5085 2636 5089 2640
rect 5093 2636 5097 2640
rect 5113 2636 5117 2640
rect 5123 2636 5127 2640
rect 5145 2636 5149 2640
rect 5245 2636 5249 2640
rect 5265 2636 5269 2640
rect 5285 2636 5289 2640
rect 5305 2636 5309 2640
rect 5325 2636 5329 2640
rect 5345 2636 5349 2640
rect 5365 2636 5369 2640
rect 5385 2636 5389 2640
rect 5491 2636 5495 2640
rect 5511 2636 5515 2640
rect 5531 2636 5535 2640
rect 5551 2636 5555 2640
rect 5571 2636 5575 2640
rect 5591 2636 5595 2640
rect 5611 2636 5615 2640
rect 5631 2636 5635 2640
rect 5731 2636 5735 2640
rect 85 2559 89 2616
rect 171 2559 175 2616
rect 292 2573 296 2616
rect 85 2547 94 2559
rect 166 2547 175 2559
rect 85 2464 89 2547
rect 171 2464 175 2547
rect 285 2561 294 2573
rect 285 2504 289 2561
rect 314 2559 318 2596
rect 322 2592 326 2596
rect 322 2586 341 2592
rect 334 2573 341 2586
rect 314 2524 320 2547
rect 334 2524 341 2561
rect 305 2518 320 2524
rect 325 2518 341 2524
rect 412 2519 416 2576
rect 305 2504 309 2518
rect 325 2504 329 2518
rect 406 2507 416 2519
rect 400 2476 406 2507
rect 420 2499 424 2576
rect 428 2519 432 2576
rect 551 2559 555 2616
rect 546 2547 555 2559
rect 428 2507 435 2519
rect 447 2507 455 2519
rect 420 2480 426 2487
rect 420 2476 435 2480
rect 400 2472 415 2476
rect 411 2464 415 2472
rect 431 2464 435 2476
rect 451 2464 455 2507
rect 551 2464 555 2547
rect 651 2539 655 2616
rect 671 2539 675 2616
rect 771 2591 775 2596
rect 762 2584 775 2591
rect 762 2539 766 2584
rect 791 2573 795 2596
rect 786 2561 795 2573
rect 646 2527 655 2539
rect 651 2504 655 2527
rect 659 2527 674 2539
rect 659 2504 663 2527
rect 762 2516 766 2527
rect 762 2508 780 2516
rect 776 2504 780 2508
rect 784 2504 788 2561
rect 811 2519 815 2596
rect 934 2592 938 2596
rect 919 2586 938 2592
rect 919 2573 926 2586
rect 919 2524 926 2561
rect 942 2559 946 2596
rect 964 2573 968 2616
rect 966 2561 975 2573
rect 940 2524 946 2547
rect 806 2507 813 2519
rect 919 2518 935 2524
rect 940 2518 955 2524
rect 806 2464 810 2507
rect 931 2504 935 2518
rect 951 2504 955 2518
rect 971 2504 975 2561
rect 1085 2519 1089 2596
rect 1105 2573 1109 2596
rect 1125 2591 1129 2596
rect 1125 2584 1138 2591
rect 1105 2561 1114 2573
rect 1087 2507 1094 2519
rect 1090 2464 1094 2507
rect 1112 2504 1116 2561
rect 1134 2539 1138 2584
rect 1233 2576 1237 2596
rect 1223 2569 1237 2576
rect 1243 2576 1247 2596
rect 1243 2569 1251 2576
rect 1223 2553 1229 2569
rect 1226 2541 1229 2553
rect 1134 2516 1138 2527
rect 1120 2508 1138 2516
rect 1120 2504 1124 2508
rect 1225 2464 1229 2541
rect 1245 2553 1251 2569
rect 1245 2541 1254 2553
rect 1245 2464 1249 2541
rect 1331 2539 1335 2596
rect 1341 2553 1345 2596
rect 1361 2590 1365 2596
rect 1367 2578 1379 2590
rect 1341 2541 1354 2553
rect 1326 2527 1335 2539
rect 1331 2464 1335 2527
rect 1353 2464 1357 2541
rect 1375 2504 1379 2578
rect 1508 2519 1512 2576
rect 1485 2507 1493 2519
rect 1505 2507 1512 2519
rect 1485 2464 1489 2507
rect 1516 2499 1520 2576
rect 1524 2519 1528 2576
rect 1611 2559 1615 2616
rect 1711 2591 1715 2596
rect 1606 2547 1615 2559
rect 1524 2507 1534 2519
rect 1514 2480 1520 2487
rect 1505 2476 1520 2480
rect 1534 2476 1540 2507
rect 1505 2464 1509 2476
rect 1525 2472 1540 2476
rect 1525 2464 1529 2472
rect 1611 2464 1615 2547
rect 1702 2584 1715 2591
rect 1702 2539 1706 2584
rect 1731 2573 1735 2596
rect 1726 2561 1735 2573
rect 1702 2516 1706 2527
rect 1702 2508 1720 2516
rect 1716 2504 1720 2508
rect 1724 2504 1728 2561
rect 1751 2519 1755 2596
rect 1865 2519 1869 2596
rect 1885 2573 1889 2596
rect 1905 2591 1909 2596
rect 1991 2591 1995 2596
rect 1905 2584 1918 2591
rect 1885 2561 1894 2573
rect 1746 2507 1753 2519
rect 1867 2507 1874 2519
rect 1746 2464 1750 2507
rect 1870 2464 1874 2507
rect 1892 2504 1896 2561
rect 1914 2539 1918 2584
rect 1982 2584 1995 2591
rect 1982 2539 1986 2584
rect 2011 2573 2015 2596
rect 2006 2561 2015 2573
rect 1914 2516 1918 2527
rect 1900 2508 1918 2516
rect 1982 2516 1986 2527
rect 1982 2508 2000 2516
rect 1900 2504 1904 2508
rect 1996 2504 2000 2508
rect 2004 2504 2008 2561
rect 2031 2519 2035 2596
rect 2168 2519 2172 2576
rect 2026 2507 2033 2519
rect 2145 2507 2153 2519
rect 2165 2507 2172 2519
rect 2026 2464 2030 2507
rect 2145 2464 2149 2507
rect 2176 2499 2180 2576
rect 2184 2519 2188 2576
rect 2292 2573 2296 2616
rect 2285 2561 2294 2573
rect 2184 2507 2194 2519
rect 2174 2480 2180 2487
rect 2165 2476 2180 2480
rect 2194 2476 2200 2507
rect 2285 2504 2289 2561
rect 2314 2559 2318 2596
rect 2322 2592 2326 2596
rect 2322 2586 2341 2592
rect 2334 2573 2341 2586
rect 2413 2576 2417 2596
rect 2409 2569 2417 2576
rect 2423 2576 2427 2596
rect 2423 2569 2437 2576
rect 2314 2524 2320 2547
rect 2334 2524 2341 2561
rect 2409 2553 2415 2569
rect 2406 2541 2415 2553
rect 2305 2518 2320 2524
rect 2325 2518 2341 2524
rect 2305 2504 2309 2518
rect 2325 2504 2329 2518
rect 2165 2464 2169 2476
rect 2185 2472 2200 2476
rect 2185 2464 2189 2472
rect 2411 2464 2415 2541
rect 2431 2553 2437 2569
rect 2431 2541 2434 2553
rect 2431 2464 2435 2541
rect 2565 2519 2569 2596
rect 2585 2573 2589 2596
rect 2605 2591 2609 2596
rect 2691 2591 2695 2596
rect 2605 2584 2618 2591
rect 2585 2561 2594 2573
rect 2567 2507 2574 2519
rect 2570 2464 2574 2507
rect 2592 2504 2596 2561
rect 2614 2539 2618 2584
rect 2682 2584 2695 2591
rect 2682 2539 2686 2584
rect 2711 2573 2715 2596
rect 2706 2561 2715 2573
rect 2614 2516 2618 2527
rect 2600 2508 2618 2516
rect 2682 2516 2686 2527
rect 2682 2508 2700 2516
rect 2600 2504 2604 2508
rect 2696 2504 2700 2508
rect 2704 2504 2708 2561
rect 2731 2519 2735 2596
rect 2852 2573 2856 2616
rect 2845 2561 2854 2573
rect 2726 2507 2733 2519
rect 2726 2464 2730 2507
rect 2845 2504 2849 2561
rect 2874 2559 2878 2596
rect 2882 2592 2886 2596
rect 2882 2586 2901 2592
rect 2894 2573 2901 2586
rect 2874 2524 2880 2547
rect 2894 2524 2901 2561
rect 2865 2518 2880 2524
rect 2885 2518 2901 2524
rect 2985 2559 2989 2616
rect 3071 2591 3075 2596
rect 3062 2584 3075 2591
rect 2985 2547 2994 2559
rect 2865 2504 2869 2518
rect 2885 2504 2889 2518
rect 2985 2464 2989 2547
rect 3062 2539 3066 2584
rect 3091 2573 3095 2596
rect 3086 2561 3095 2573
rect 3062 2516 3066 2527
rect 3062 2508 3080 2516
rect 3076 2504 3080 2508
rect 3084 2504 3088 2561
rect 3111 2519 3115 2596
rect 3233 2576 3237 2596
rect 3229 2569 3237 2576
rect 3243 2576 3247 2596
rect 3243 2569 3257 2576
rect 3229 2553 3235 2569
rect 3226 2541 3235 2553
rect 3106 2507 3113 2519
rect 3106 2464 3110 2507
rect 3231 2464 3235 2541
rect 3251 2553 3257 2569
rect 3251 2541 3254 2553
rect 3251 2464 3255 2541
rect 3388 2519 3392 2576
rect 3365 2507 3373 2519
rect 3385 2507 3392 2519
rect 3365 2464 3369 2507
rect 3396 2499 3400 2576
rect 3404 2519 3408 2576
rect 3491 2539 3495 2596
rect 3501 2553 3505 2596
rect 3521 2590 3525 2596
rect 3527 2578 3539 2590
rect 3501 2541 3514 2553
rect 3486 2527 3495 2539
rect 3404 2507 3414 2519
rect 3394 2480 3400 2487
rect 3385 2476 3400 2480
rect 3414 2476 3420 2507
rect 3385 2464 3389 2476
rect 3405 2472 3420 2476
rect 3405 2464 3409 2472
rect 3491 2464 3495 2527
rect 3513 2464 3517 2541
rect 3535 2504 3539 2578
rect 3633 2576 3637 2596
rect 3629 2569 3637 2576
rect 3643 2576 3647 2596
rect 3754 2588 3758 2596
rect 3741 2581 3758 2588
rect 3643 2569 3657 2576
rect 3629 2553 3635 2569
rect 3626 2541 3635 2553
rect 3631 2464 3635 2541
rect 3651 2553 3657 2569
rect 3651 2541 3654 2553
rect 3651 2464 3655 2541
rect 3741 2539 3747 2581
rect 3762 2573 3766 2596
rect 3782 2582 3786 2596
rect 3790 2591 3794 2596
rect 3790 2587 3820 2591
rect 3782 2575 3795 2582
rect 3791 2573 3795 2575
rect 3791 2561 3793 2573
rect 3762 2532 3766 2561
rect 3747 2527 3755 2532
rect 3735 2526 3755 2527
rect 3762 2526 3775 2532
rect 3751 2504 3755 2526
rect 3771 2504 3775 2526
rect 3791 2504 3795 2561
rect 3814 2539 3820 2587
rect 3911 2539 3915 2616
rect 3931 2539 3935 2616
rect 3999 2572 4003 2616
rect 4047 2584 4051 2596
rect 4059 2592 4063 2596
rect 4059 2588 4080 2592
rect 4047 2580 4070 2584
rect 3999 2560 4046 2572
rect 3811 2527 3814 2539
rect 3906 2527 3915 2539
rect 3811 2504 3815 2527
rect 3911 2504 3915 2527
rect 3919 2527 3934 2539
rect 3919 2504 3923 2527
rect 3999 2464 4003 2560
rect 4066 2552 4070 2580
rect 4044 2546 4070 2552
rect 4076 2572 4080 2588
rect 4084 2584 4088 2596
rect 4096 2592 4100 2596
rect 4096 2588 4120 2592
rect 4084 2580 4106 2584
rect 4076 2560 4078 2572
rect 4044 2515 4048 2546
rect 4044 2503 4045 2515
rect 4076 2506 4080 2560
rect 4100 2540 4106 2580
rect 4044 2464 4048 2503
rect 4065 2500 4080 2506
rect 4065 2482 4069 2500
rect 4094 2490 4100 2528
rect 4084 2484 4100 2490
rect 4064 2464 4068 2470
rect 4084 2464 4088 2484
rect 4115 2482 4120 2588
rect 4136 2545 4141 2578
rect 4149 2568 4153 2616
rect 4169 2590 4173 2616
rect 4214 2590 4218 2616
rect 4234 2608 4238 2616
rect 4234 2596 4258 2608
rect 4206 2578 4214 2584
rect 4149 2562 4175 2568
rect 4136 2533 4150 2545
rect 4104 2470 4109 2482
rect 4104 2464 4108 2470
rect 4149 2444 4153 2533
rect 4170 2484 4175 2562
rect 4206 2528 4210 2578
rect 4234 2557 4238 2596
rect 4284 2571 4288 2616
rect 4304 2587 4308 2616
rect 4279 2559 4288 2571
rect 4324 2567 4328 2616
rect 4374 2570 4378 2596
rect 4300 2563 4328 2567
rect 4364 2566 4378 2570
rect 4231 2545 4238 2557
rect 4206 2522 4218 2528
rect 4169 2472 4194 2484
rect 4169 2444 4173 2472
rect 4214 2464 4218 2522
rect 4234 2464 4238 2545
rect 4279 2464 4283 2559
rect 4300 2541 4304 2563
rect 4299 2444 4303 2529
rect 4319 2444 4323 2555
rect 4364 2531 4368 2566
rect 4364 2464 4368 2519
rect 4386 2511 4390 2596
rect 4410 2590 4414 2596
rect 4384 2464 4388 2499
rect 4402 2494 4406 2578
rect 4422 2553 4426 2596
rect 4474 2553 4478 2596
rect 4486 2590 4490 2596
rect 4426 2541 4428 2553
rect 4404 2464 4408 2482
rect 4424 2464 4428 2541
rect 4472 2541 4474 2553
rect 4472 2464 4476 2541
rect 4494 2494 4498 2578
rect 4510 2511 4514 2596
rect 4522 2570 4526 2596
rect 4522 2566 4536 2570
rect 4532 2531 4536 2566
rect 4572 2567 4576 2616
rect 4592 2587 4596 2616
rect 4612 2571 4616 2616
rect 4662 2608 4666 2616
rect 4642 2596 4666 2608
rect 4572 2563 4600 2567
rect 4492 2464 4496 2482
rect 4512 2464 4516 2499
rect 4532 2464 4536 2519
rect 4577 2444 4581 2555
rect 4596 2541 4600 2563
rect 4612 2559 4621 2571
rect 4597 2444 4601 2529
rect 4617 2464 4621 2559
rect 4662 2557 4666 2596
rect 4682 2590 4686 2616
rect 4727 2590 4731 2616
rect 4686 2578 4694 2584
rect 4662 2545 4669 2557
rect 4662 2464 4666 2545
rect 4690 2528 4694 2578
rect 4747 2568 4751 2616
rect 4800 2592 4804 2596
rect 4682 2522 4694 2528
rect 4725 2562 4751 2568
rect 4780 2588 4804 2592
rect 4682 2464 4686 2522
rect 4725 2484 4730 2562
rect 4759 2545 4764 2578
rect 4750 2533 4764 2545
rect 4706 2472 4731 2484
rect 4727 2444 4731 2472
rect 4747 2444 4751 2533
rect 4780 2482 4785 2588
rect 4812 2584 4816 2596
rect 4837 2592 4841 2596
rect 4794 2580 4816 2584
rect 4820 2588 4841 2592
rect 4794 2540 4800 2580
rect 4820 2572 4824 2588
rect 4849 2584 4853 2596
rect 4822 2560 4824 2572
rect 4800 2490 4806 2528
rect 4820 2506 4824 2560
rect 4830 2580 4853 2584
rect 4830 2552 4834 2580
rect 4897 2572 4901 2616
rect 4854 2560 4901 2572
rect 4830 2546 4856 2552
rect 4852 2515 4856 2546
rect 4820 2500 4835 2506
rect 4855 2503 4856 2515
rect 4800 2484 4816 2490
rect 4791 2470 4796 2482
rect 4792 2464 4796 2470
rect 4812 2464 4816 2484
rect 4831 2482 4835 2500
rect 4832 2464 4836 2470
rect 4852 2464 4856 2503
rect 4897 2464 4901 2560
rect 4955 2559 4959 2596
rect 4975 2558 4979 2616
rect 4985 2584 4989 2616
rect 5007 2604 5011 2616
rect 5009 2592 5011 2604
rect 5017 2604 5021 2616
rect 5017 2592 5019 2604
rect 4985 2580 5018 2584
rect 4955 2504 4959 2547
rect 4975 2464 4979 2546
rect 4994 2531 4998 2560
rect 4989 2523 4998 2531
rect 4989 2464 4993 2523
rect 5014 2516 5018 2580
rect 5015 2504 5018 2516
rect 5009 2464 5013 2504
rect 5023 2482 5027 2592
rect 5039 2502 5043 2616
rect 5085 2612 5089 2616
rect 5055 2608 5089 2612
rect 5021 2464 5025 2470
rect 5041 2464 5045 2490
rect 5055 2482 5059 2608
rect 5093 2604 5097 2616
rect 5067 2600 5097 2604
rect 5079 2599 5097 2600
rect 5113 2595 5117 2616
rect 5093 2591 5117 2595
rect 5093 2496 5099 2591
rect 5123 2567 5127 2616
rect 5123 2509 5127 2555
rect 5145 2528 5149 2596
rect 5147 2516 5149 2528
rect 5123 2503 5131 2509
rect 5145 2504 5149 2516
rect 5245 2576 5249 2596
rect 5265 2576 5269 2596
rect 5285 2576 5289 2596
rect 5305 2576 5309 2596
rect 5325 2576 5329 2596
rect 5345 2576 5349 2596
rect 5245 2564 5258 2576
rect 5285 2564 5298 2576
rect 5325 2564 5338 2576
rect 5365 2573 5369 2596
rect 5385 2573 5389 2596
rect 5245 2504 5249 2564
rect 5265 2504 5269 2564
rect 5285 2504 5289 2564
rect 5305 2504 5309 2564
rect 5325 2504 5329 2564
rect 5345 2504 5349 2564
rect 5365 2561 5374 2573
rect 5386 2561 5389 2573
rect 5365 2504 5369 2561
rect 5385 2504 5389 2561
rect 5491 2573 5495 2596
rect 5511 2573 5515 2596
rect 5531 2576 5535 2596
rect 5551 2576 5555 2596
rect 5571 2576 5575 2596
rect 5591 2576 5595 2596
rect 5611 2576 5615 2596
rect 5631 2576 5635 2596
rect 5491 2561 5494 2573
rect 5506 2561 5515 2573
rect 5542 2564 5555 2576
rect 5582 2564 5595 2576
rect 5622 2564 5635 2576
rect 5731 2573 5735 2596
rect 5491 2504 5495 2561
rect 5511 2504 5515 2561
rect 5531 2504 5535 2564
rect 5551 2504 5555 2564
rect 5571 2504 5575 2564
rect 5591 2504 5595 2564
rect 5611 2504 5615 2564
rect 5631 2504 5635 2564
rect 5726 2561 5735 2573
rect 5731 2504 5735 2561
rect 5067 2470 5091 2472
rect 5055 2468 5091 2470
rect 5087 2464 5091 2468
rect 5095 2464 5099 2496
rect 5115 2444 5119 2484
rect 5127 2474 5131 2503
rect 5123 2467 5131 2474
rect 5123 2444 5127 2467
rect 85 2420 89 2424
rect 171 2420 175 2424
rect 285 2420 289 2424
rect 305 2420 309 2424
rect 325 2420 329 2424
rect 411 2420 415 2424
rect 431 2420 435 2424
rect 451 2420 455 2424
rect 551 2420 555 2424
rect 651 2420 655 2424
rect 659 2420 663 2424
rect 776 2420 780 2424
rect 784 2420 788 2424
rect 806 2420 810 2424
rect 931 2420 935 2424
rect 951 2420 955 2424
rect 971 2420 975 2424
rect 1090 2420 1094 2424
rect 1112 2420 1116 2424
rect 1120 2420 1124 2424
rect 1225 2420 1229 2424
rect 1245 2420 1249 2424
rect 1331 2420 1335 2424
rect 1353 2420 1357 2424
rect 1375 2420 1379 2424
rect 1485 2420 1489 2424
rect 1505 2420 1509 2424
rect 1525 2420 1529 2424
rect 1611 2420 1615 2424
rect 1716 2420 1720 2424
rect 1724 2420 1728 2424
rect 1746 2420 1750 2424
rect 1870 2420 1874 2424
rect 1892 2420 1896 2424
rect 1900 2420 1904 2424
rect 1996 2420 2000 2424
rect 2004 2420 2008 2424
rect 2026 2420 2030 2424
rect 2145 2420 2149 2424
rect 2165 2420 2169 2424
rect 2185 2420 2189 2424
rect 2285 2420 2289 2424
rect 2305 2420 2309 2424
rect 2325 2420 2329 2424
rect 2411 2420 2415 2424
rect 2431 2420 2435 2424
rect 2570 2420 2574 2424
rect 2592 2420 2596 2424
rect 2600 2420 2604 2424
rect 2696 2420 2700 2424
rect 2704 2420 2708 2424
rect 2726 2420 2730 2424
rect 2845 2420 2849 2424
rect 2865 2420 2869 2424
rect 2885 2420 2889 2424
rect 2985 2420 2989 2424
rect 3076 2420 3080 2424
rect 3084 2420 3088 2424
rect 3106 2420 3110 2424
rect 3231 2420 3235 2424
rect 3251 2420 3255 2424
rect 3365 2420 3369 2424
rect 3385 2420 3389 2424
rect 3405 2420 3409 2424
rect 3491 2420 3495 2424
rect 3513 2420 3517 2424
rect 3535 2420 3539 2424
rect 3631 2420 3635 2424
rect 3651 2420 3655 2424
rect 3751 2420 3755 2424
rect 3771 2420 3775 2424
rect 3791 2420 3795 2424
rect 3811 2420 3815 2424
rect 3911 2420 3915 2424
rect 3919 2420 3923 2424
rect 3999 2420 4003 2424
rect 4044 2420 4048 2424
rect 4064 2420 4068 2424
rect 4084 2420 4088 2424
rect 4104 2420 4108 2424
rect 4149 2420 4153 2424
rect 4169 2420 4173 2424
rect 4214 2420 4218 2424
rect 4234 2420 4238 2424
rect 4279 2420 4283 2424
rect 4299 2420 4303 2424
rect 4319 2420 4323 2424
rect 4364 2420 4368 2424
rect 4384 2420 4388 2424
rect 4404 2420 4408 2424
rect 4424 2420 4428 2424
rect 4472 2420 4476 2424
rect 4492 2420 4496 2424
rect 4512 2420 4516 2424
rect 4532 2420 4536 2424
rect 4577 2420 4581 2424
rect 4597 2420 4601 2424
rect 4617 2420 4621 2424
rect 4662 2420 4666 2424
rect 4682 2420 4686 2424
rect 4727 2420 4731 2424
rect 4747 2420 4751 2424
rect 4792 2420 4796 2424
rect 4812 2420 4816 2424
rect 4832 2420 4836 2424
rect 4852 2420 4856 2424
rect 4897 2420 4901 2424
rect 4955 2420 4959 2424
rect 4975 2420 4979 2424
rect 4989 2420 4993 2424
rect 5009 2420 5013 2424
rect 5021 2420 5025 2424
rect 5041 2420 5045 2424
rect 5087 2420 5091 2424
rect 5095 2420 5099 2424
rect 5115 2420 5119 2424
rect 5123 2420 5127 2424
rect 5145 2420 5149 2424
rect 5245 2420 5249 2424
rect 5265 2420 5269 2424
rect 5285 2420 5289 2424
rect 5305 2420 5309 2424
rect 5325 2420 5329 2424
rect 5345 2420 5349 2424
rect 5365 2420 5369 2424
rect 5385 2420 5389 2424
rect 5491 2420 5495 2424
rect 5511 2420 5515 2424
rect 5531 2420 5535 2424
rect 5551 2420 5555 2424
rect 5571 2420 5575 2424
rect 5591 2420 5595 2424
rect 5611 2420 5615 2424
rect 5631 2420 5635 2424
rect 5731 2420 5735 2424
rect 83 2396 87 2400
rect 105 2396 109 2400
rect 205 2396 209 2400
rect 225 2396 229 2400
rect 245 2396 249 2400
rect 331 2396 335 2400
rect 351 2396 355 2400
rect 456 2396 460 2400
rect 464 2396 468 2400
rect 486 2396 490 2400
rect 610 2396 614 2400
rect 632 2396 636 2400
rect 640 2396 644 2400
rect 765 2396 769 2400
rect 785 2396 789 2400
rect 805 2396 809 2400
rect 905 2396 909 2400
rect 925 2396 929 2400
rect 1035 2396 1039 2400
rect 1055 2396 1059 2400
rect 1065 2396 1069 2400
rect 1151 2396 1155 2400
rect 1265 2396 1269 2400
rect 1285 2396 1289 2400
rect 1305 2396 1309 2400
rect 1405 2396 1409 2400
rect 1425 2396 1429 2400
rect 1445 2396 1449 2400
rect 1570 2396 1574 2400
rect 1592 2396 1596 2400
rect 1600 2396 1604 2400
rect 1705 2396 1709 2400
rect 1725 2396 1729 2400
rect 1745 2396 1749 2400
rect 1845 2396 1849 2400
rect 1865 2396 1869 2400
rect 1885 2396 1889 2400
rect 1985 2396 1989 2400
rect 2005 2396 2009 2400
rect 2025 2396 2029 2400
rect 2079 2396 2083 2400
rect 2124 2396 2128 2400
rect 2144 2396 2148 2400
rect 2164 2396 2168 2400
rect 2184 2396 2188 2400
rect 2229 2396 2233 2400
rect 2249 2396 2253 2400
rect 2294 2396 2298 2400
rect 2314 2396 2318 2400
rect 2359 2396 2363 2400
rect 2379 2396 2383 2400
rect 2399 2396 2403 2400
rect 2444 2396 2448 2400
rect 2464 2396 2468 2400
rect 2484 2396 2488 2400
rect 2504 2396 2508 2400
rect 2603 2396 2607 2400
rect 2625 2396 2629 2400
rect 2736 2396 2740 2400
rect 2744 2396 2748 2400
rect 2766 2396 2770 2400
rect 2876 2396 2880 2400
rect 2884 2396 2888 2400
rect 2906 2396 2910 2400
rect 3025 2396 3029 2400
rect 3045 2396 3049 2400
rect 3151 2396 3155 2400
rect 3171 2396 3175 2400
rect 3285 2396 3289 2400
rect 3305 2396 3309 2400
rect 3325 2396 3329 2400
rect 3411 2396 3415 2400
rect 3419 2396 3423 2400
rect 3556 2396 3560 2400
rect 3564 2396 3568 2400
rect 3586 2396 3590 2400
rect 3691 2396 3695 2400
rect 3711 2396 3715 2400
rect 3811 2396 3815 2400
rect 3833 2396 3837 2400
rect 3899 2396 3903 2400
rect 3944 2396 3948 2400
rect 3964 2396 3968 2400
rect 3984 2396 3988 2400
rect 4004 2396 4008 2400
rect 4049 2396 4053 2400
rect 4069 2396 4073 2400
rect 4114 2396 4118 2400
rect 4134 2396 4138 2400
rect 4179 2396 4183 2400
rect 4199 2396 4203 2400
rect 4219 2396 4223 2400
rect 4264 2396 4268 2400
rect 4284 2396 4288 2400
rect 4304 2396 4308 2400
rect 4324 2396 4328 2400
rect 4411 2396 4415 2400
rect 4433 2396 4437 2400
rect 4455 2396 4459 2400
rect 4551 2396 4555 2400
rect 4571 2396 4575 2400
rect 4591 2396 4595 2400
rect 4611 2396 4615 2400
rect 4711 2396 4715 2400
rect 4731 2396 4735 2400
rect 4843 2396 4847 2400
rect 4865 2396 4869 2400
rect 4951 2396 4955 2400
rect 5051 2396 5055 2400
rect 5071 2396 5075 2400
rect 5091 2396 5095 2400
rect 5111 2396 5115 2400
rect 5211 2396 5215 2400
rect 5231 2396 5235 2400
rect 5331 2396 5335 2400
rect 5431 2396 5435 2400
rect 5451 2396 5455 2400
rect 5551 2396 5555 2400
rect 5651 2396 5685 2400
rect 5701 2396 5705 2400
rect 5711 2396 5715 2400
rect 83 2310 87 2316
rect 83 2298 85 2310
rect 105 2293 109 2356
rect 205 2313 209 2356
rect 225 2344 229 2356
rect 245 2348 249 2356
rect 245 2344 260 2348
rect 225 2340 240 2344
rect 234 2333 240 2340
rect 205 2301 213 2313
rect 225 2301 232 2313
rect 105 2281 114 2293
rect 83 2230 85 2242
rect 83 2224 87 2230
rect 105 2204 109 2281
rect 228 2244 232 2301
rect 236 2244 240 2321
rect 254 2313 260 2344
rect 244 2301 254 2313
rect 244 2244 248 2301
rect 331 2279 335 2356
rect 326 2267 335 2279
rect 329 2251 335 2267
rect 351 2279 355 2356
rect 456 2312 460 2316
rect 442 2304 460 2312
rect 442 2293 446 2304
rect 351 2267 354 2279
rect 351 2251 357 2267
rect 329 2244 337 2251
rect 333 2224 337 2244
rect 343 2244 357 2251
rect 343 2224 347 2244
rect 442 2236 446 2281
rect 464 2259 468 2316
rect 486 2313 490 2356
rect 610 2313 614 2356
rect 486 2301 493 2313
rect 607 2301 614 2313
rect 466 2247 475 2259
rect 442 2229 455 2236
rect 451 2224 455 2229
rect 471 2224 475 2247
rect 491 2224 495 2301
rect 605 2224 609 2301
rect 632 2259 636 2316
rect 640 2312 644 2316
rect 765 2313 769 2356
rect 785 2344 789 2356
rect 805 2348 809 2356
rect 805 2344 820 2348
rect 785 2340 800 2344
rect 794 2333 800 2340
rect 640 2304 658 2312
rect 654 2293 658 2304
rect 765 2301 773 2313
rect 785 2301 792 2313
rect 625 2247 634 2259
rect 625 2224 629 2247
rect 654 2236 658 2281
rect 788 2244 792 2301
rect 796 2244 800 2321
rect 814 2313 820 2344
rect 804 2301 814 2313
rect 804 2244 808 2301
rect 905 2279 909 2356
rect 906 2267 909 2279
rect 903 2251 909 2267
rect 925 2279 929 2356
rect 1035 2311 1039 2316
rect 1055 2293 1059 2316
rect 1065 2312 1069 2316
rect 1065 2307 1078 2312
rect 925 2267 934 2279
rect 925 2251 931 2267
rect 903 2244 917 2251
rect 645 2229 658 2236
rect 645 2224 649 2229
rect 913 2224 917 2244
rect 923 2244 931 2251
rect 923 2224 927 2244
rect 1025 2232 1035 2244
rect 1025 2224 1029 2232
rect 1055 2217 1059 2281
rect 1045 2211 1059 2217
rect 1074 2273 1078 2307
rect 1074 2216 1078 2261
rect 1151 2259 1155 2316
rect 1265 2313 1269 2356
rect 1285 2344 1289 2356
rect 1305 2348 1309 2356
rect 1305 2344 1320 2348
rect 1285 2340 1300 2344
rect 1294 2333 1300 2340
rect 1265 2301 1273 2313
rect 1285 2301 1292 2313
rect 1146 2247 1155 2259
rect 1151 2224 1155 2247
rect 1288 2244 1292 2301
rect 1296 2244 1300 2321
rect 1314 2313 1320 2344
rect 1304 2301 1314 2313
rect 1304 2244 1308 2301
rect 1405 2259 1409 2316
rect 1425 2302 1429 2316
rect 1445 2302 1449 2316
rect 1570 2313 1574 2356
rect 1425 2296 1440 2302
rect 1445 2296 1461 2302
rect 1567 2301 1574 2313
rect 1434 2273 1440 2296
rect 1405 2247 1414 2259
rect 1065 2211 1078 2216
rect 1045 2204 1049 2211
rect 1065 2204 1069 2211
rect 1412 2204 1416 2247
rect 1434 2224 1438 2261
rect 1454 2259 1461 2296
rect 1454 2234 1461 2247
rect 1442 2228 1461 2234
rect 1442 2224 1446 2228
rect 1565 2224 1569 2301
rect 1592 2259 1596 2316
rect 1600 2312 1604 2316
rect 1600 2304 1618 2312
rect 1614 2293 1618 2304
rect 1585 2247 1594 2259
rect 1585 2224 1589 2247
rect 1614 2236 1618 2281
rect 1705 2259 1709 2316
rect 1725 2302 1729 2316
rect 1745 2302 1749 2316
rect 1845 2313 1849 2356
rect 1865 2344 1869 2356
rect 1885 2348 1889 2356
rect 1885 2344 1900 2348
rect 1865 2340 1880 2344
rect 1874 2333 1880 2340
rect 1725 2296 1740 2302
rect 1745 2296 1761 2302
rect 1845 2301 1853 2313
rect 1865 2301 1872 2313
rect 1734 2273 1740 2296
rect 1705 2247 1714 2259
rect 1605 2229 1618 2236
rect 1605 2224 1609 2229
rect 1712 2204 1716 2247
rect 1734 2224 1738 2261
rect 1754 2259 1761 2296
rect 1754 2234 1761 2247
rect 1868 2244 1872 2301
rect 1876 2244 1880 2321
rect 1894 2313 1900 2344
rect 1985 2313 1989 2356
rect 2005 2344 2009 2356
rect 2025 2348 2029 2356
rect 2025 2344 2040 2348
rect 2005 2340 2020 2344
rect 2014 2333 2020 2340
rect 1884 2301 1894 2313
rect 1985 2301 1993 2313
rect 2005 2301 2012 2313
rect 1884 2244 1888 2301
rect 2008 2244 2012 2301
rect 2016 2244 2020 2321
rect 2034 2313 2040 2344
rect 2024 2301 2034 2313
rect 2024 2244 2028 2301
rect 2079 2260 2083 2356
rect 2124 2317 2128 2356
rect 2144 2350 2148 2356
rect 2145 2320 2149 2338
rect 2164 2336 2168 2356
rect 2184 2350 2188 2356
rect 2184 2338 2189 2350
rect 2164 2330 2180 2336
rect 2124 2305 2125 2317
rect 2145 2314 2160 2320
rect 2124 2274 2128 2305
rect 2124 2268 2150 2274
rect 2079 2248 2126 2260
rect 1742 2228 1761 2234
rect 1742 2224 1746 2228
rect 2079 2204 2083 2248
rect 2146 2240 2150 2268
rect 2127 2236 2150 2240
rect 2156 2260 2160 2314
rect 2174 2292 2180 2330
rect 2156 2248 2158 2260
rect 2127 2224 2131 2236
rect 2156 2232 2160 2248
rect 2180 2240 2186 2280
rect 2139 2228 2160 2232
rect 2164 2236 2186 2240
rect 2139 2224 2143 2228
rect 2164 2224 2168 2236
rect 2195 2232 2200 2338
rect 2229 2287 2233 2376
rect 2249 2348 2253 2376
rect 2249 2336 2274 2348
rect 2216 2275 2230 2287
rect 2216 2242 2221 2275
rect 2250 2258 2255 2336
rect 2294 2298 2298 2356
rect 2176 2228 2200 2232
rect 2229 2252 2255 2258
rect 2286 2292 2298 2298
rect 2176 2224 2180 2228
rect 2229 2204 2233 2252
rect 2286 2242 2290 2292
rect 2314 2275 2318 2356
rect 2311 2263 2318 2275
rect 2286 2236 2294 2242
rect 2249 2204 2253 2230
rect 2294 2204 2298 2230
rect 2314 2224 2318 2263
rect 2359 2261 2363 2356
rect 2379 2291 2383 2376
rect 2359 2249 2368 2261
rect 2380 2257 2384 2279
rect 2399 2265 2403 2376
rect 2444 2301 2448 2356
rect 2464 2321 2468 2356
rect 2484 2338 2488 2356
rect 2380 2253 2408 2257
rect 2314 2212 2338 2224
rect 2314 2204 2318 2212
rect 2364 2204 2368 2249
rect 2384 2204 2388 2233
rect 2404 2204 2408 2253
rect 2444 2254 2448 2289
rect 2444 2250 2458 2254
rect 2454 2224 2458 2250
rect 2466 2224 2470 2309
rect 2482 2242 2486 2326
rect 2504 2279 2508 2356
rect 2603 2310 2607 2316
rect 2603 2298 2605 2310
rect 2506 2267 2508 2279
rect 2625 2293 2629 2356
rect 2736 2312 2740 2316
rect 2722 2304 2740 2312
rect 2722 2293 2726 2304
rect 2625 2281 2634 2293
rect 2490 2224 2494 2230
rect 2502 2224 2506 2267
rect 2603 2230 2605 2242
rect 2603 2224 2607 2230
rect 2625 2204 2629 2281
rect 2722 2236 2726 2281
rect 2744 2259 2748 2316
rect 2766 2313 2770 2356
rect 2766 2301 2773 2313
rect 2876 2312 2880 2316
rect 2862 2304 2880 2312
rect 2746 2247 2755 2259
rect 2722 2229 2735 2236
rect 2731 2224 2735 2229
rect 2751 2224 2755 2247
rect 2771 2224 2775 2301
rect 2862 2293 2866 2304
rect 2862 2236 2866 2281
rect 2884 2259 2888 2316
rect 2906 2313 2910 2356
rect 2906 2301 2913 2313
rect 2886 2247 2895 2259
rect 2862 2229 2875 2236
rect 2871 2224 2875 2229
rect 2891 2224 2895 2247
rect 2911 2224 2915 2301
rect 3025 2279 3029 2356
rect 3026 2267 3029 2279
rect 3023 2251 3029 2267
rect 3045 2279 3049 2356
rect 3151 2279 3155 2356
rect 3045 2267 3054 2279
rect 3146 2267 3155 2279
rect 3045 2251 3051 2267
rect 3023 2244 3037 2251
rect 3033 2224 3037 2244
rect 3043 2244 3051 2251
rect 3149 2251 3155 2267
rect 3171 2279 3175 2356
rect 3171 2267 3174 2279
rect 3171 2251 3177 2267
rect 3149 2244 3157 2251
rect 3043 2224 3047 2244
rect 3153 2224 3157 2244
rect 3163 2244 3177 2251
rect 3285 2259 3289 2316
rect 3305 2302 3309 2316
rect 3325 2302 3329 2316
rect 3305 2296 3320 2302
rect 3325 2296 3341 2302
rect 3314 2273 3320 2296
rect 3285 2247 3294 2259
rect 3163 2224 3167 2244
rect 3292 2204 3296 2247
rect 3314 2224 3318 2261
rect 3334 2259 3341 2296
rect 3411 2293 3415 2316
rect 3406 2281 3415 2293
rect 3419 2293 3423 2316
rect 3556 2312 3560 2316
rect 3542 2304 3560 2312
rect 3542 2293 3546 2304
rect 3419 2281 3434 2293
rect 3334 2234 3341 2247
rect 3322 2228 3341 2234
rect 3322 2224 3326 2228
rect 3411 2204 3415 2281
rect 3431 2204 3435 2281
rect 3542 2236 3546 2281
rect 3564 2259 3568 2316
rect 3586 2313 3590 2356
rect 3586 2301 3593 2313
rect 3566 2247 3575 2259
rect 3542 2229 3555 2236
rect 3551 2224 3555 2229
rect 3571 2224 3575 2247
rect 3591 2224 3595 2301
rect 3691 2279 3695 2356
rect 3686 2267 3695 2279
rect 3689 2251 3695 2267
rect 3711 2279 3715 2356
rect 3811 2293 3815 2356
rect 3833 2310 3837 2316
rect 3835 2298 3837 2310
rect 3806 2281 3815 2293
rect 3711 2267 3714 2279
rect 3711 2251 3717 2267
rect 3689 2244 3697 2251
rect 3693 2224 3697 2244
rect 3703 2244 3717 2251
rect 3703 2224 3707 2244
rect 3811 2204 3815 2281
rect 3899 2260 3903 2356
rect 3944 2317 3948 2356
rect 3964 2350 3968 2356
rect 3965 2320 3969 2338
rect 3984 2336 3988 2356
rect 4004 2350 4008 2356
rect 4004 2338 4009 2350
rect 3984 2330 4000 2336
rect 3944 2305 3945 2317
rect 3965 2314 3980 2320
rect 3944 2274 3948 2305
rect 3944 2268 3970 2274
rect 3899 2248 3946 2260
rect 3835 2230 3837 2242
rect 3833 2224 3837 2230
rect 3899 2204 3903 2248
rect 3966 2240 3970 2268
rect 3947 2236 3970 2240
rect 3976 2260 3980 2314
rect 3994 2292 4000 2330
rect 3976 2248 3978 2260
rect 3947 2224 3951 2236
rect 3976 2232 3980 2248
rect 4000 2240 4006 2280
rect 3959 2228 3980 2232
rect 3984 2236 4006 2240
rect 3959 2224 3963 2228
rect 3984 2224 3988 2236
rect 4015 2232 4020 2338
rect 4049 2287 4053 2376
rect 4069 2348 4073 2376
rect 4069 2336 4094 2348
rect 4036 2275 4050 2287
rect 4036 2242 4041 2275
rect 4070 2258 4075 2336
rect 4114 2298 4118 2356
rect 3996 2228 4020 2232
rect 4049 2252 4075 2258
rect 4106 2292 4118 2298
rect 3996 2224 4000 2228
rect 4049 2204 4053 2252
rect 4106 2242 4110 2292
rect 4134 2275 4138 2356
rect 4131 2263 4138 2275
rect 4106 2236 4114 2242
rect 4069 2204 4073 2230
rect 4114 2204 4118 2230
rect 4134 2224 4138 2263
rect 4179 2261 4183 2356
rect 4199 2291 4203 2376
rect 4179 2249 4188 2261
rect 4200 2257 4204 2279
rect 4219 2265 4223 2376
rect 4264 2301 4268 2356
rect 4284 2321 4288 2356
rect 4304 2338 4308 2356
rect 4200 2253 4228 2257
rect 4134 2212 4158 2224
rect 4134 2204 4138 2212
rect 4184 2204 4188 2249
rect 4204 2204 4208 2233
rect 4224 2204 4228 2253
rect 4264 2254 4268 2289
rect 4264 2250 4278 2254
rect 4274 2224 4278 2250
rect 4286 2224 4290 2309
rect 4302 2242 4306 2326
rect 4324 2279 4328 2356
rect 4411 2293 4415 2356
rect 4406 2281 4415 2293
rect 4326 2267 4328 2279
rect 4310 2224 4314 2230
rect 4322 2224 4326 2267
rect 4411 2224 4415 2281
rect 4433 2279 4437 2356
rect 4421 2267 4434 2279
rect 4421 2224 4425 2267
rect 4455 2242 4459 2316
rect 4551 2294 4555 2316
rect 4571 2294 4575 2316
rect 4535 2293 4555 2294
rect 4547 2288 4555 2293
rect 4562 2288 4575 2294
rect 4447 2230 4459 2242
rect 4541 2239 4547 2281
rect 4562 2259 4566 2288
rect 4591 2259 4595 2316
rect 4611 2293 4615 2316
rect 4611 2281 4614 2293
rect 4591 2247 4593 2259
rect 4541 2232 4558 2239
rect 4441 2224 4445 2230
rect 4554 2224 4558 2232
rect 4562 2224 4566 2247
rect 4591 2245 4595 2247
rect 4582 2238 4595 2245
rect 4582 2224 4586 2238
rect 4614 2233 4620 2281
rect 4711 2279 4715 2356
rect 4706 2267 4715 2279
rect 4709 2251 4715 2267
rect 4731 2279 4735 2356
rect 4843 2310 4847 2316
rect 4843 2298 4845 2310
rect 4865 2293 4869 2356
rect 4865 2281 4874 2293
rect 4731 2267 4734 2279
rect 4731 2251 4737 2267
rect 4709 2244 4717 2251
rect 4590 2229 4620 2233
rect 4590 2224 4594 2229
rect 4713 2224 4717 2244
rect 4723 2244 4737 2251
rect 4723 2224 4727 2244
rect 4843 2230 4845 2242
rect 4843 2224 4847 2230
rect 4865 2204 4869 2281
rect 4951 2273 4955 2356
rect 5051 2294 5055 2316
rect 5071 2294 5075 2316
rect 5035 2293 5055 2294
rect 5047 2288 5055 2293
rect 5062 2288 5075 2294
rect 4946 2261 4955 2273
rect 4951 2204 4955 2261
rect 5041 2239 5047 2281
rect 5062 2259 5066 2288
rect 5091 2259 5095 2316
rect 5111 2293 5115 2316
rect 5111 2281 5114 2293
rect 5091 2247 5093 2259
rect 5041 2232 5058 2239
rect 5054 2224 5058 2232
rect 5062 2224 5066 2247
rect 5091 2245 5095 2247
rect 5082 2238 5095 2245
rect 5082 2224 5086 2238
rect 5114 2233 5120 2281
rect 5211 2279 5215 2356
rect 5206 2267 5215 2279
rect 5209 2251 5215 2267
rect 5231 2279 5235 2356
rect 5651 2388 5655 2396
rect 5671 2388 5675 2392
rect 5681 2388 5685 2396
rect 5231 2267 5234 2279
rect 5231 2251 5237 2267
rect 5331 2259 5335 2316
rect 5431 2279 5435 2356
rect 5426 2267 5435 2279
rect 5209 2244 5217 2251
rect 5090 2229 5120 2233
rect 5090 2224 5094 2229
rect 5213 2224 5217 2244
rect 5223 2244 5237 2251
rect 5326 2247 5335 2259
rect 5223 2224 5227 2244
rect 5331 2224 5335 2247
rect 5429 2251 5435 2267
rect 5451 2279 5455 2356
rect 5451 2267 5454 2279
rect 5551 2273 5555 2356
rect 5651 2344 5655 2348
rect 5451 2251 5457 2267
rect 5546 2261 5555 2273
rect 5429 2244 5437 2251
rect 5433 2224 5437 2244
rect 5443 2244 5457 2251
rect 5443 2224 5447 2244
rect 5551 2204 5555 2261
rect 5643 2340 5655 2344
rect 5643 2259 5647 2340
rect 5671 2303 5675 2308
rect 5681 2304 5685 2308
rect 5662 2299 5675 2303
rect 5662 2293 5667 2299
rect 5701 2294 5705 2316
rect 5675 2290 5705 2294
rect 5711 2293 5715 2316
rect 5643 2221 5647 2247
rect 5661 2250 5666 2281
rect 5711 2281 5714 2293
rect 5661 2244 5675 2250
rect 5671 2232 5675 2244
rect 5681 2232 5685 2278
rect 5701 2232 5705 2236
rect 5711 2232 5715 2281
rect 5643 2216 5655 2221
rect 5651 2212 5655 2216
rect 5651 2184 5655 2192
rect 5671 2188 5675 2192
rect 5681 2188 5685 2192
rect 5701 2184 5705 2192
rect 5711 2188 5715 2192
rect 83 2180 87 2184
rect 105 2180 109 2184
rect 228 2180 232 2184
rect 236 2180 240 2184
rect 244 2180 248 2184
rect 333 2180 337 2184
rect 343 2180 347 2184
rect 451 2180 455 2184
rect 471 2180 475 2184
rect 491 2180 495 2184
rect 605 2180 609 2184
rect 625 2180 629 2184
rect 645 2180 649 2184
rect 788 2180 792 2184
rect 796 2180 800 2184
rect 804 2180 808 2184
rect 913 2180 917 2184
rect 923 2180 927 2184
rect 1025 2180 1029 2184
rect 1045 2180 1049 2184
rect 1065 2180 1069 2184
rect 1151 2180 1155 2184
rect 1288 2180 1292 2184
rect 1296 2180 1300 2184
rect 1304 2180 1308 2184
rect 1412 2180 1416 2184
rect 1434 2180 1438 2184
rect 1442 2180 1446 2184
rect 1565 2180 1569 2184
rect 1585 2180 1589 2184
rect 1605 2180 1609 2184
rect 1712 2180 1716 2184
rect 1734 2180 1738 2184
rect 1742 2180 1746 2184
rect 1868 2180 1872 2184
rect 1876 2180 1880 2184
rect 1884 2180 1888 2184
rect 2008 2180 2012 2184
rect 2016 2180 2020 2184
rect 2024 2180 2028 2184
rect 2079 2180 2083 2184
rect 2127 2180 2131 2184
rect 2139 2180 2143 2184
rect 2164 2180 2168 2184
rect 2176 2180 2180 2184
rect 2229 2180 2233 2184
rect 2249 2180 2253 2184
rect 2294 2180 2298 2184
rect 2314 2180 2318 2184
rect 2364 2180 2368 2184
rect 2384 2180 2388 2184
rect 2404 2180 2408 2184
rect 2454 2180 2458 2184
rect 2466 2180 2470 2184
rect 2490 2180 2494 2184
rect 2502 2180 2506 2184
rect 2603 2180 2607 2184
rect 2625 2180 2629 2184
rect 2731 2180 2735 2184
rect 2751 2180 2755 2184
rect 2771 2180 2775 2184
rect 2871 2180 2875 2184
rect 2891 2180 2895 2184
rect 2911 2180 2915 2184
rect 3033 2180 3037 2184
rect 3043 2180 3047 2184
rect 3153 2180 3157 2184
rect 3163 2180 3167 2184
rect 3292 2180 3296 2184
rect 3314 2180 3318 2184
rect 3322 2180 3326 2184
rect 3411 2180 3415 2184
rect 3431 2180 3435 2184
rect 3551 2180 3555 2184
rect 3571 2180 3575 2184
rect 3591 2180 3595 2184
rect 3693 2180 3697 2184
rect 3703 2180 3707 2184
rect 3811 2180 3815 2184
rect 3833 2180 3837 2184
rect 3899 2180 3903 2184
rect 3947 2180 3951 2184
rect 3959 2180 3963 2184
rect 3984 2180 3988 2184
rect 3996 2180 4000 2184
rect 4049 2180 4053 2184
rect 4069 2180 4073 2184
rect 4114 2180 4118 2184
rect 4134 2180 4138 2184
rect 4184 2180 4188 2184
rect 4204 2180 4208 2184
rect 4224 2180 4228 2184
rect 4274 2180 4278 2184
rect 4286 2180 4290 2184
rect 4310 2180 4314 2184
rect 4322 2180 4326 2184
rect 4411 2180 4415 2184
rect 4421 2180 4425 2184
rect 4441 2180 4445 2184
rect 4554 2180 4558 2184
rect 4562 2180 4566 2184
rect 4582 2180 4586 2184
rect 4590 2180 4594 2184
rect 4713 2180 4717 2184
rect 4723 2180 4727 2184
rect 4843 2180 4847 2184
rect 4865 2180 4869 2184
rect 4951 2180 4955 2184
rect 5054 2180 5058 2184
rect 5062 2180 5066 2184
rect 5082 2180 5086 2184
rect 5090 2180 5094 2184
rect 5213 2180 5217 2184
rect 5223 2180 5227 2184
rect 5331 2180 5335 2184
rect 5433 2180 5437 2184
rect 5443 2180 5447 2184
rect 5551 2180 5555 2184
rect 5651 2180 5705 2184
rect 103 2156 107 2160
rect 125 2156 129 2160
rect 268 2156 272 2160
rect 276 2156 280 2160
rect 284 2156 288 2160
rect 374 2156 378 2160
rect 382 2156 386 2160
rect 404 2156 408 2160
rect 525 2156 529 2160
rect 625 2156 629 2160
rect 645 2156 649 2160
rect 665 2156 669 2160
rect 772 2156 776 2160
rect 794 2156 798 2160
rect 802 2156 806 2160
rect 892 2156 896 2160
rect 900 2156 904 2160
rect 908 2156 912 2160
rect 1088 2156 1092 2160
rect 1096 2156 1100 2160
rect 1104 2156 1108 2160
rect 1205 2156 1209 2160
rect 1225 2156 1229 2160
rect 1245 2156 1249 2160
rect 1345 2156 1349 2160
rect 1365 2156 1369 2160
rect 1385 2156 1389 2160
rect 1492 2156 1496 2160
rect 1514 2156 1518 2160
rect 1522 2156 1526 2160
rect 1648 2156 1652 2160
rect 1656 2156 1660 2160
rect 1664 2156 1668 2160
rect 1751 2156 1755 2160
rect 1771 2156 1775 2160
rect 1791 2156 1795 2160
rect 1894 2156 1898 2160
rect 1902 2156 1906 2160
rect 1924 2156 1928 2160
rect 2105 2156 2109 2160
rect 2125 2156 2129 2160
rect 2145 2156 2149 2160
rect 2288 2156 2292 2160
rect 2296 2156 2300 2160
rect 2304 2156 2308 2160
rect 2359 2156 2363 2160
rect 2407 2156 2411 2160
rect 2419 2156 2423 2160
rect 2444 2156 2448 2160
rect 2456 2156 2460 2160
rect 2509 2156 2513 2160
rect 2529 2156 2533 2160
rect 2574 2156 2578 2160
rect 2594 2156 2598 2160
rect 2644 2156 2648 2160
rect 2664 2156 2668 2160
rect 2684 2156 2688 2160
rect 2734 2156 2738 2160
rect 2746 2156 2750 2160
rect 2770 2156 2774 2160
rect 2782 2156 2786 2160
rect 2871 2156 2875 2160
rect 2891 2156 2895 2160
rect 2911 2156 2915 2160
rect 3033 2156 3037 2160
rect 3043 2156 3047 2160
rect 3133 2156 3137 2160
rect 3143 2156 3147 2160
rect 3271 2156 3275 2160
rect 3291 2156 3295 2160
rect 3415 2156 3419 2160
rect 3435 2156 3439 2160
rect 3445 2156 3449 2160
rect 3534 2156 3538 2160
rect 3542 2156 3546 2160
rect 3564 2156 3568 2160
rect 3705 2156 3709 2160
rect 3812 2156 3816 2160
rect 3820 2156 3824 2160
rect 3828 2156 3832 2160
rect 3971 2156 3975 2160
rect 4115 2156 4119 2160
rect 4135 2156 4139 2160
rect 4145 2156 4149 2160
rect 4253 2156 4257 2160
rect 4263 2156 4267 2160
rect 4365 2156 4369 2160
rect 4385 2156 4389 2160
rect 4405 2156 4409 2160
rect 4491 2156 4495 2160
rect 4511 2156 4515 2160
rect 4531 2156 4535 2160
rect 4633 2156 4637 2160
rect 4643 2156 4647 2160
rect 4753 2156 4757 2160
rect 4763 2156 4767 2160
rect 4905 2156 4909 2160
rect 4925 2156 4929 2160
rect 4945 2156 4949 2160
rect 5045 2156 5049 2160
rect 5065 2156 5069 2160
rect 5085 2156 5089 2160
rect 5171 2156 5175 2160
rect 5271 2156 5275 2160
rect 5291 2156 5295 2160
rect 5393 2156 5397 2160
rect 5403 2156 5407 2160
rect 5511 2156 5515 2160
rect 5625 2156 5629 2160
rect 5711 2156 5715 2160
rect 5731 2156 5735 2160
rect 5751 2156 5755 2160
rect 103 2110 107 2116
rect 103 2098 105 2110
rect 125 2059 129 2136
rect 374 2112 378 2116
rect 359 2106 378 2112
rect 125 2047 134 2059
rect 103 2030 105 2042
rect 103 2024 107 2030
rect 125 1984 129 2047
rect 268 2039 272 2096
rect 245 2027 253 2039
rect 265 2027 272 2039
rect 245 1984 249 2027
rect 276 2019 280 2096
rect 284 2039 288 2096
rect 359 2093 366 2106
rect 359 2044 366 2081
rect 382 2079 386 2116
rect 404 2093 408 2136
rect 406 2081 415 2093
rect 380 2044 386 2067
rect 284 2027 294 2039
rect 359 2038 375 2044
rect 380 2038 395 2044
rect 274 2000 280 2007
rect 265 1996 280 2000
rect 294 1996 300 2027
rect 371 2024 375 2038
rect 391 2024 395 2038
rect 411 2024 415 2081
rect 525 2079 529 2136
rect 525 2067 534 2079
rect 265 1984 269 1996
rect 285 1992 300 1996
rect 285 1984 289 1992
rect 525 1984 529 2067
rect 625 2039 629 2116
rect 645 2093 649 2116
rect 665 2111 669 2116
rect 665 2104 678 2111
rect 645 2081 654 2093
rect 627 2027 634 2039
rect 630 1984 634 2027
rect 652 2024 656 2081
rect 674 2059 678 2104
rect 772 2093 776 2136
rect 765 2081 774 2093
rect 674 2036 678 2047
rect 660 2028 678 2036
rect 660 2024 664 2028
rect 765 2024 769 2081
rect 794 2079 798 2116
rect 802 2112 806 2116
rect 802 2106 821 2112
rect 814 2093 821 2106
rect 794 2044 800 2067
rect 814 2044 821 2081
rect 785 2038 800 2044
rect 805 2038 821 2044
rect 892 2039 896 2096
rect 785 2024 789 2038
rect 805 2024 809 2038
rect 886 2027 896 2039
rect 880 1996 886 2027
rect 900 2019 904 2096
rect 908 2039 912 2096
rect 1088 2039 1092 2096
rect 908 2027 915 2039
rect 927 2027 935 2039
rect 900 2000 906 2007
rect 900 1996 915 2000
rect 880 1992 895 1996
rect 891 1984 895 1992
rect 911 1984 915 1996
rect 931 1984 935 2027
rect 1065 2027 1073 2039
rect 1085 2027 1092 2039
rect 1065 1984 1069 2027
rect 1096 2019 1100 2096
rect 1104 2039 1108 2096
rect 1205 2039 1209 2116
rect 1225 2093 1229 2116
rect 1245 2111 1249 2116
rect 1245 2104 1258 2111
rect 1225 2081 1234 2093
rect 1104 2027 1114 2039
rect 1207 2027 1214 2039
rect 1094 2000 1100 2007
rect 1085 1996 1100 2000
rect 1114 1996 1120 2027
rect 1085 1984 1089 1996
rect 1105 1992 1120 1996
rect 1105 1984 1109 1992
rect 1210 1984 1214 2027
rect 1232 2024 1236 2081
rect 1254 2059 1258 2104
rect 1254 2036 1258 2047
rect 1345 2039 1349 2116
rect 1365 2093 1369 2116
rect 1385 2111 1389 2116
rect 1385 2104 1398 2111
rect 1365 2081 1374 2093
rect 1240 2028 1258 2036
rect 1240 2024 1244 2028
rect 1347 2027 1354 2039
rect 1350 1984 1354 2027
rect 1372 2024 1376 2081
rect 1394 2059 1398 2104
rect 1492 2093 1496 2136
rect 1485 2081 1494 2093
rect 1394 2036 1398 2047
rect 1380 2028 1398 2036
rect 1380 2024 1384 2028
rect 1485 2024 1489 2081
rect 1514 2079 1518 2116
rect 1522 2112 1526 2116
rect 1522 2106 1541 2112
rect 1534 2093 1541 2106
rect 1751 2111 1755 2116
rect 1742 2104 1755 2111
rect 1514 2044 1520 2067
rect 1534 2044 1541 2081
rect 1505 2038 1520 2044
rect 1525 2038 1541 2044
rect 1648 2039 1652 2096
rect 1505 2024 1509 2038
rect 1525 2024 1529 2038
rect 1625 2027 1633 2039
rect 1645 2027 1652 2039
rect 1625 1984 1629 2027
rect 1656 2019 1660 2096
rect 1664 2039 1668 2096
rect 1742 2059 1746 2104
rect 1771 2093 1775 2116
rect 1766 2081 1775 2093
rect 1664 2027 1674 2039
rect 1742 2036 1746 2047
rect 1742 2028 1760 2036
rect 1654 2000 1660 2007
rect 1645 1996 1660 2000
rect 1674 1996 1680 2027
rect 1756 2024 1760 2028
rect 1764 2024 1768 2081
rect 1791 2039 1795 2116
rect 1894 2112 1898 2116
rect 1879 2106 1898 2112
rect 1879 2093 1886 2106
rect 1879 2044 1886 2081
rect 1902 2079 1906 2116
rect 1924 2093 1928 2136
rect 2105 2120 2109 2136
rect 2085 2114 2109 2120
rect 1926 2081 1935 2093
rect 1900 2044 1906 2067
rect 1786 2027 1793 2039
rect 1879 2038 1895 2044
rect 1900 2038 1915 2044
rect 1645 1984 1649 1996
rect 1665 1992 1680 1996
rect 1665 1984 1669 1992
rect 1786 1984 1790 2027
rect 1891 2024 1895 2038
rect 1911 2024 1915 2038
rect 1931 2024 1935 2081
rect 2085 2059 2091 2114
rect 2125 2093 2129 2136
rect 2126 2081 2129 2093
rect 2085 2047 2094 2059
rect 2085 2024 2091 2047
rect 2041 2020 2091 2024
rect 2041 2012 2045 2020
rect 2061 2012 2065 2020
rect 2125 2012 2129 2081
rect 2105 2008 2129 2012
rect 2105 2004 2109 2008
rect 2125 2004 2129 2008
rect 2145 2059 2149 2136
rect 2145 2047 2154 2059
rect 2145 2012 2149 2047
rect 2288 2039 2292 2096
rect 2265 2027 2273 2039
rect 2285 2027 2292 2039
rect 2145 2008 2169 2012
rect 2145 2004 2149 2008
rect 2165 2004 2169 2008
rect 2041 1948 2045 1952
rect 2061 1948 2065 1952
rect 2265 1984 2269 2027
rect 2296 2019 2300 2096
rect 2304 2039 2308 2096
rect 2359 2092 2363 2136
rect 2407 2104 2411 2116
rect 2419 2112 2423 2116
rect 2419 2108 2440 2112
rect 2407 2100 2430 2104
rect 2359 2080 2406 2092
rect 2304 2027 2314 2039
rect 2294 2000 2300 2007
rect 2285 1996 2300 2000
rect 2314 1996 2320 2027
rect 2285 1984 2289 1996
rect 2305 1992 2320 1996
rect 2305 1984 2309 1992
rect 2359 1984 2363 2080
rect 2426 2072 2430 2100
rect 2404 2066 2430 2072
rect 2436 2092 2440 2108
rect 2444 2104 2448 2116
rect 2456 2112 2460 2116
rect 2456 2108 2480 2112
rect 2444 2100 2466 2104
rect 2436 2080 2438 2092
rect 2404 2035 2408 2066
rect 2404 2023 2405 2035
rect 2436 2026 2440 2080
rect 2460 2060 2466 2100
rect 2404 1984 2408 2023
rect 2425 2020 2440 2026
rect 2425 2002 2429 2020
rect 2454 2010 2460 2048
rect 2444 2004 2460 2010
rect 2424 1984 2428 1990
rect 2444 1984 2448 2004
rect 2475 2002 2480 2108
rect 2496 2065 2501 2098
rect 2509 2088 2513 2136
rect 2529 2110 2533 2136
rect 2574 2110 2578 2136
rect 2594 2128 2598 2136
rect 2594 2116 2618 2128
rect 2566 2098 2574 2104
rect 2509 2082 2535 2088
rect 2496 2053 2510 2065
rect 2464 1990 2469 2002
rect 2464 1984 2468 1990
rect 2509 1964 2513 2053
rect 2530 2004 2535 2082
rect 2566 2048 2570 2098
rect 2594 2077 2598 2116
rect 2644 2091 2648 2136
rect 2664 2107 2668 2136
rect 2639 2079 2648 2091
rect 2684 2087 2688 2136
rect 2734 2090 2738 2116
rect 2660 2083 2688 2087
rect 2724 2086 2738 2090
rect 2591 2065 2598 2077
rect 2566 2042 2578 2048
rect 2529 1992 2554 2004
rect 2529 1964 2533 1992
rect 2574 1984 2578 2042
rect 2594 1984 2598 2065
rect 2639 1984 2643 2079
rect 2660 2061 2664 2083
rect 2659 1964 2663 2049
rect 2679 1964 2683 2075
rect 2724 2051 2728 2086
rect 2724 1984 2728 2039
rect 2746 2031 2750 2116
rect 2770 2110 2774 2116
rect 2744 1984 2748 2019
rect 2762 2014 2766 2098
rect 2782 2073 2786 2116
rect 2871 2111 2875 2116
rect 2862 2104 2875 2111
rect 2786 2061 2788 2073
rect 2764 1984 2768 2002
rect 2784 1984 2788 2061
rect 2862 2059 2866 2104
rect 2891 2093 2895 2116
rect 2886 2081 2895 2093
rect 2862 2036 2866 2047
rect 2862 2028 2880 2036
rect 2876 2024 2880 2028
rect 2884 2024 2888 2081
rect 2911 2039 2915 2116
rect 3033 2096 3037 2116
rect 3023 2089 3037 2096
rect 3043 2096 3047 2116
rect 3133 2096 3137 2116
rect 3043 2089 3051 2096
rect 3023 2073 3029 2089
rect 3026 2061 3029 2073
rect 2906 2027 2913 2039
rect 2906 1984 2910 2027
rect 3025 1984 3029 2061
rect 3045 2073 3051 2089
rect 3129 2089 3137 2096
rect 3143 2096 3147 2116
rect 3143 2089 3157 2096
rect 3129 2073 3135 2089
rect 3045 2061 3054 2073
rect 3126 2061 3135 2073
rect 3045 1984 3049 2061
rect 3131 1984 3135 2061
rect 3151 2073 3157 2089
rect 3151 2061 3154 2073
rect 3151 1984 3155 2061
rect 3271 2059 3275 2136
rect 3291 2059 3295 2136
rect 3415 2110 3419 2116
rect 3401 2098 3413 2110
rect 3266 2047 3275 2059
rect 3271 2024 3275 2047
rect 3279 2047 3294 2059
rect 3279 2024 3283 2047
rect 3401 2024 3405 2098
rect 3435 2073 3439 2116
rect 3426 2061 3439 2073
rect 3423 1984 3427 2061
rect 3445 2059 3449 2116
rect 3534 2112 3538 2116
rect 3519 2106 3538 2112
rect 3519 2093 3526 2106
rect 3445 2047 3454 2059
rect 3445 1984 3449 2047
rect 3519 2044 3526 2081
rect 3542 2079 3546 2116
rect 3564 2093 3568 2136
rect 3705 2093 3709 2116
rect 3566 2081 3575 2093
rect 3540 2044 3546 2067
rect 3519 2038 3535 2044
rect 3540 2038 3555 2044
rect 3531 2024 3535 2038
rect 3551 2024 3555 2038
rect 3571 2024 3575 2081
rect 3705 2081 3714 2093
rect 3705 2024 3709 2081
rect 3812 2039 3816 2096
rect 3806 2027 3816 2039
rect 3800 1996 3806 2027
rect 3820 2019 3824 2096
rect 3828 2039 3832 2096
rect 3971 2093 3975 2116
rect 4115 2110 4119 2116
rect 3966 2081 3975 2093
rect 3828 2027 3835 2039
rect 3847 2027 3855 2039
rect 3820 2000 3826 2007
rect 3820 1996 3835 2000
rect 3800 1992 3815 1996
rect 3811 1984 3815 1992
rect 3831 1984 3835 1996
rect 3851 1984 3855 2027
rect 3971 2024 3975 2081
rect 4101 2098 4113 2110
rect 4101 2024 4105 2098
rect 4135 2073 4139 2116
rect 4126 2061 4139 2073
rect 4123 1984 4127 2061
rect 4145 2059 4149 2116
rect 4253 2096 4257 2116
rect 4243 2089 4257 2096
rect 4263 2096 4267 2116
rect 4263 2089 4271 2096
rect 4243 2073 4249 2089
rect 4246 2061 4249 2073
rect 4145 2047 4154 2059
rect 4145 1984 4149 2047
rect 4245 1984 4249 2061
rect 4265 2073 4271 2089
rect 4265 2061 4274 2073
rect 4265 1984 4269 2061
rect 4365 2039 4369 2116
rect 4385 2093 4389 2116
rect 4405 2111 4409 2116
rect 4491 2111 4495 2116
rect 4405 2104 4418 2111
rect 4385 2081 4394 2093
rect 4367 2027 4374 2039
rect 4370 1984 4374 2027
rect 4392 2024 4396 2081
rect 4414 2059 4418 2104
rect 4482 2104 4495 2111
rect 4482 2059 4486 2104
rect 4511 2093 4515 2116
rect 4506 2081 4515 2093
rect 4414 2036 4418 2047
rect 4400 2028 4418 2036
rect 4482 2036 4486 2047
rect 4482 2028 4500 2036
rect 4400 2024 4404 2028
rect 4496 2024 4500 2028
rect 4504 2024 4508 2081
rect 4531 2039 4535 2116
rect 4633 2096 4637 2116
rect 4629 2089 4637 2096
rect 4643 2096 4647 2116
rect 4753 2096 4757 2116
rect 4643 2089 4657 2096
rect 4629 2073 4635 2089
rect 4626 2061 4635 2073
rect 4526 2027 4533 2039
rect 4526 1984 4530 2027
rect 4631 1984 4635 2061
rect 4651 2073 4657 2089
rect 4749 2089 4757 2096
rect 4763 2096 4767 2116
rect 4763 2089 4777 2096
rect 4749 2073 4755 2089
rect 4651 2061 4654 2073
rect 4746 2061 4755 2073
rect 4651 1984 4655 2061
rect 4751 1984 4755 2061
rect 4771 2073 4777 2089
rect 4771 2061 4774 2073
rect 4771 1984 4775 2061
rect 4905 2039 4909 2116
rect 4925 2093 4929 2116
rect 4945 2111 4949 2116
rect 4945 2104 4958 2111
rect 4925 2081 4934 2093
rect 4907 2027 4914 2039
rect 4910 1984 4914 2027
rect 4932 2024 4936 2081
rect 4954 2059 4958 2104
rect 4954 2036 4958 2047
rect 5045 2039 5049 2116
rect 5065 2093 5069 2116
rect 5085 2111 5089 2116
rect 5085 2104 5098 2111
rect 5065 2081 5074 2093
rect 4940 2028 4958 2036
rect 4940 2024 4944 2028
rect 5047 2027 5054 2039
rect 5050 1984 5054 2027
rect 5072 2024 5076 2081
rect 5094 2059 5098 2104
rect 5171 2079 5175 2136
rect 5166 2067 5175 2079
rect 5094 2036 5098 2047
rect 5080 2028 5098 2036
rect 5080 2024 5084 2028
rect 5171 1984 5175 2067
rect 5271 2059 5275 2136
rect 5291 2059 5295 2136
rect 5393 2096 5397 2116
rect 5389 2089 5397 2096
rect 5403 2096 5407 2116
rect 5403 2089 5417 2096
rect 5389 2073 5395 2089
rect 5386 2061 5395 2073
rect 5266 2047 5275 2059
rect 5271 2024 5275 2047
rect 5279 2047 5294 2059
rect 5279 2024 5283 2047
rect 5391 1984 5395 2061
rect 5411 2073 5417 2089
rect 5511 2079 5515 2136
rect 5411 2061 5414 2073
rect 5506 2067 5515 2079
rect 5411 1984 5415 2061
rect 5511 1984 5515 2067
rect 5625 2079 5629 2136
rect 5711 2111 5715 2116
rect 5702 2104 5715 2111
rect 5625 2067 5634 2079
rect 5625 1984 5629 2067
rect 5702 2059 5706 2104
rect 5731 2093 5735 2116
rect 5726 2081 5735 2093
rect 5702 2036 5706 2047
rect 5702 2028 5720 2036
rect 5716 2024 5720 2028
rect 5724 2024 5728 2081
rect 5751 2039 5755 2116
rect 5746 2027 5753 2039
rect 5746 1984 5750 2027
rect 103 1940 107 1944
rect 125 1940 129 1944
rect 245 1940 249 1944
rect 265 1940 269 1944
rect 285 1940 289 1944
rect 371 1940 375 1944
rect 391 1940 395 1944
rect 411 1940 415 1944
rect 525 1940 529 1944
rect 630 1940 634 1944
rect 652 1940 656 1944
rect 660 1940 664 1944
rect 765 1940 769 1944
rect 785 1940 789 1944
rect 805 1940 809 1944
rect 891 1940 895 1944
rect 911 1940 915 1944
rect 931 1940 935 1944
rect 1065 1940 1069 1944
rect 1085 1940 1089 1944
rect 1105 1940 1109 1944
rect 1210 1940 1214 1944
rect 1232 1940 1236 1944
rect 1240 1940 1244 1944
rect 1350 1940 1354 1944
rect 1372 1940 1376 1944
rect 1380 1940 1384 1944
rect 1485 1940 1489 1944
rect 1505 1940 1509 1944
rect 1525 1940 1529 1944
rect 1625 1940 1629 1944
rect 1645 1940 1649 1944
rect 1665 1940 1669 1944
rect 1756 1940 1760 1944
rect 1764 1940 1768 1944
rect 1786 1940 1790 1944
rect 1891 1940 1895 1944
rect 1911 1940 1915 1944
rect 1931 1940 1935 1944
rect 2105 1940 2109 1944
rect 2125 1940 2129 1944
rect 2145 1940 2149 1944
rect 2165 1940 2169 1944
rect 2265 1940 2269 1944
rect 2285 1940 2289 1944
rect 2305 1940 2309 1944
rect 2359 1940 2363 1944
rect 2404 1940 2408 1944
rect 2424 1940 2428 1944
rect 2444 1940 2448 1944
rect 2464 1940 2468 1944
rect 2509 1940 2513 1944
rect 2529 1940 2533 1944
rect 2574 1940 2578 1944
rect 2594 1940 2598 1944
rect 2639 1940 2643 1944
rect 2659 1940 2663 1944
rect 2679 1940 2683 1944
rect 2724 1940 2728 1944
rect 2744 1940 2748 1944
rect 2764 1940 2768 1944
rect 2784 1940 2788 1944
rect 2876 1940 2880 1944
rect 2884 1940 2888 1944
rect 2906 1940 2910 1944
rect 3025 1940 3029 1944
rect 3045 1940 3049 1944
rect 3131 1940 3135 1944
rect 3151 1940 3155 1944
rect 3271 1940 3275 1944
rect 3279 1940 3283 1944
rect 3401 1940 3405 1944
rect 3423 1940 3427 1944
rect 3445 1940 3449 1944
rect 3531 1940 3535 1944
rect 3551 1940 3555 1944
rect 3571 1940 3575 1944
rect 3705 1940 3709 1944
rect 3811 1940 3815 1944
rect 3831 1940 3835 1944
rect 3851 1940 3855 1944
rect 3971 1940 3975 1944
rect 4101 1940 4105 1944
rect 4123 1940 4127 1944
rect 4145 1940 4149 1944
rect 4245 1940 4249 1944
rect 4265 1940 4269 1944
rect 4370 1940 4374 1944
rect 4392 1940 4396 1944
rect 4400 1940 4404 1944
rect 4496 1940 4500 1944
rect 4504 1940 4508 1944
rect 4526 1940 4530 1944
rect 4631 1940 4635 1944
rect 4651 1940 4655 1944
rect 4751 1940 4755 1944
rect 4771 1940 4775 1944
rect 4910 1940 4914 1944
rect 4932 1940 4936 1944
rect 4940 1940 4944 1944
rect 5050 1940 5054 1944
rect 5072 1940 5076 1944
rect 5080 1940 5084 1944
rect 5171 1940 5175 1944
rect 5271 1940 5275 1944
rect 5279 1940 5283 1944
rect 5391 1940 5395 1944
rect 5411 1940 5415 1944
rect 5511 1940 5515 1944
rect 5625 1940 5629 1944
rect 5716 1940 5720 1944
rect 5724 1940 5728 1944
rect 5746 1940 5750 1944
rect 85 1916 89 1920
rect 105 1916 109 1920
rect 125 1916 129 1920
rect 211 1916 215 1920
rect 231 1916 235 1920
rect 251 1916 255 1920
rect 370 1916 374 1920
rect 392 1916 396 1920
rect 400 1916 404 1920
rect 505 1916 509 1920
rect 525 1916 529 1920
rect 545 1916 549 1920
rect 677 1916 681 1920
rect 685 1916 689 1920
rect 771 1916 775 1920
rect 791 1916 795 1920
rect 811 1916 815 1920
rect 945 1916 949 1920
rect 1070 1916 1074 1920
rect 1092 1916 1096 1920
rect 1100 1916 1104 1920
rect 1210 1916 1214 1920
rect 1232 1916 1236 1920
rect 1240 1916 1244 1920
rect 1345 1916 1349 1920
rect 1450 1916 1454 1920
rect 1472 1916 1476 1920
rect 1480 1916 1484 1920
rect 1576 1916 1580 1920
rect 1584 1916 1588 1920
rect 1606 1916 1610 1920
rect 1730 1916 1734 1920
rect 1752 1916 1756 1920
rect 1760 1916 1764 1920
rect 1865 1916 1869 1920
rect 1885 1916 1889 1920
rect 1985 1916 1989 1920
rect 2005 1916 2009 1920
rect 2125 1916 2129 1920
rect 2145 1916 2149 1920
rect 2199 1916 2203 1920
rect 2244 1916 2248 1920
rect 2264 1916 2268 1920
rect 2284 1916 2288 1920
rect 2304 1916 2308 1920
rect 2349 1916 2353 1920
rect 2369 1916 2373 1920
rect 2414 1916 2418 1920
rect 2434 1916 2438 1920
rect 2479 1916 2483 1920
rect 2499 1916 2503 1920
rect 2519 1916 2523 1920
rect 2564 1916 2568 1920
rect 2584 1916 2588 1920
rect 2604 1916 2608 1920
rect 2624 1916 2628 1920
rect 2711 1916 2715 1920
rect 2731 1916 2735 1920
rect 2845 1916 2849 1920
rect 2865 1916 2869 1920
rect 2885 1916 2889 1920
rect 2990 1916 2994 1920
rect 3012 1916 3016 1920
rect 3020 1916 3024 1920
rect 3111 1916 3115 1920
rect 3119 1916 3123 1920
rect 3231 1916 3265 1920
rect 3281 1916 3285 1920
rect 3291 1916 3295 1920
rect 3405 1916 3409 1920
rect 3491 1916 3495 1920
rect 3501 1916 3505 1920
rect 3531 1916 3535 1920
rect 3541 1916 3545 1920
rect 3670 1916 3674 1920
rect 3692 1916 3696 1920
rect 3700 1916 3704 1920
rect 3830 1916 3834 1920
rect 3852 1916 3856 1920
rect 3860 1916 3864 1920
rect 3956 1916 3960 1920
rect 3964 1916 3968 1920
rect 3986 1916 3990 1920
rect 4105 1916 4109 1920
rect 4125 1916 4129 1920
rect 4225 1916 4229 1920
rect 4245 1916 4249 1920
rect 4265 1916 4269 1920
rect 4285 1916 4289 1920
rect 4385 1916 4389 1920
rect 4405 1916 4409 1920
rect 4496 1916 4500 1920
rect 4504 1916 4508 1920
rect 4526 1916 4530 1920
rect 4641 1916 4645 1920
rect 4663 1916 4667 1920
rect 4685 1916 4689 1920
rect 4797 1916 4801 1920
rect 4805 1916 4809 1920
rect 4905 1916 4909 1920
rect 4925 1916 4929 1920
rect 5025 1916 5029 1920
rect 5045 1916 5049 1920
rect 5065 1916 5069 1920
rect 5085 1916 5089 1920
rect 5185 1916 5189 1920
rect 5297 1916 5301 1920
rect 5305 1916 5309 1920
rect 5396 1916 5400 1920
rect 5404 1916 5408 1920
rect 5426 1916 5430 1920
rect 5550 1916 5554 1920
rect 5572 1916 5576 1920
rect 5580 1916 5584 1920
rect 5671 1916 5675 1920
rect 5691 1916 5695 1920
rect 85 1833 89 1876
rect 105 1864 109 1876
rect 125 1868 129 1876
rect 125 1864 140 1868
rect 105 1860 120 1864
rect 114 1853 120 1860
rect 85 1821 93 1833
rect 105 1821 112 1833
rect 108 1764 112 1821
rect 116 1764 120 1841
rect 134 1833 140 1864
rect 124 1821 134 1833
rect 211 1822 215 1836
rect 231 1822 235 1836
rect 124 1764 128 1821
rect 199 1816 215 1822
rect 220 1816 235 1822
rect 199 1779 206 1816
rect 220 1793 226 1816
rect 199 1754 206 1767
rect 199 1748 218 1754
rect 214 1744 218 1748
rect 222 1744 226 1781
rect 251 1779 255 1836
rect 370 1833 374 1876
rect 367 1821 374 1833
rect 246 1767 255 1779
rect 244 1724 248 1767
rect 365 1744 369 1821
rect 392 1779 396 1836
rect 400 1832 404 1836
rect 505 1833 509 1876
rect 525 1864 529 1876
rect 545 1868 549 1876
rect 545 1864 560 1868
rect 525 1860 540 1864
rect 534 1853 540 1860
rect 400 1824 418 1832
rect 414 1813 418 1824
rect 505 1821 513 1833
rect 525 1821 532 1833
rect 385 1767 394 1779
rect 385 1744 389 1767
rect 414 1756 418 1801
rect 528 1764 532 1821
rect 536 1764 540 1841
rect 554 1833 560 1864
rect 544 1821 554 1833
rect 544 1764 548 1821
rect 677 1813 681 1836
rect 666 1801 681 1813
rect 685 1813 689 1836
rect 771 1822 775 1836
rect 791 1822 795 1836
rect 759 1816 775 1822
rect 780 1816 795 1822
rect 685 1801 694 1813
rect 405 1749 418 1756
rect 405 1744 409 1749
rect 665 1724 669 1801
rect 685 1724 689 1801
rect 759 1779 766 1816
rect 780 1793 786 1816
rect 759 1754 766 1767
rect 759 1748 778 1754
rect 774 1744 778 1748
rect 782 1744 786 1781
rect 811 1779 815 1836
rect 806 1767 815 1779
rect 945 1793 949 1876
rect 1070 1833 1074 1876
rect 1067 1821 1074 1833
rect 945 1781 954 1793
rect 804 1724 808 1767
rect 945 1724 949 1781
rect 1065 1744 1069 1821
rect 1092 1779 1096 1836
rect 1100 1832 1104 1836
rect 1210 1833 1214 1876
rect 1100 1824 1118 1832
rect 1114 1813 1118 1824
rect 1207 1821 1214 1833
rect 1085 1767 1094 1779
rect 1085 1744 1089 1767
rect 1114 1756 1118 1801
rect 1105 1749 1118 1756
rect 1105 1744 1109 1749
rect 1205 1744 1209 1821
rect 1232 1779 1236 1836
rect 1240 1832 1244 1836
rect 1240 1824 1258 1832
rect 1254 1813 1258 1824
rect 1225 1767 1234 1779
rect 1225 1744 1229 1767
rect 1254 1756 1258 1801
rect 1245 1749 1258 1756
rect 1345 1793 1349 1876
rect 1450 1833 1454 1876
rect 1447 1821 1454 1833
rect 1345 1781 1354 1793
rect 1245 1744 1249 1749
rect 1345 1724 1349 1781
rect 1445 1744 1449 1821
rect 1472 1779 1476 1836
rect 1480 1832 1484 1836
rect 1576 1832 1580 1836
rect 1480 1824 1498 1832
rect 1494 1813 1498 1824
rect 1562 1824 1580 1832
rect 1562 1813 1566 1824
rect 1465 1767 1474 1779
rect 1465 1744 1469 1767
rect 1494 1756 1498 1801
rect 1485 1749 1498 1756
rect 1562 1756 1566 1801
rect 1584 1779 1588 1836
rect 1606 1833 1610 1876
rect 1730 1833 1734 1876
rect 1606 1821 1613 1833
rect 1727 1821 1734 1833
rect 1586 1767 1595 1779
rect 1562 1749 1575 1756
rect 1485 1744 1489 1749
rect 1571 1744 1575 1749
rect 1591 1744 1595 1767
rect 1611 1744 1615 1821
rect 1725 1744 1729 1821
rect 1752 1779 1756 1836
rect 1760 1832 1764 1836
rect 1760 1824 1778 1832
rect 1774 1813 1778 1824
rect 1745 1767 1754 1779
rect 1745 1744 1749 1767
rect 1774 1756 1778 1801
rect 1865 1799 1869 1876
rect 1866 1787 1869 1799
rect 1863 1771 1869 1787
rect 1885 1799 1889 1876
rect 1985 1799 1989 1876
rect 1885 1787 1894 1799
rect 1986 1787 1989 1799
rect 1885 1771 1891 1787
rect 1863 1764 1877 1771
rect 1765 1749 1778 1756
rect 1765 1744 1769 1749
rect 1873 1744 1877 1764
rect 1883 1764 1891 1771
rect 1983 1771 1989 1787
rect 2005 1799 2009 1876
rect 2125 1832 2129 1836
rect 2145 1832 2149 1836
rect 2125 1828 2149 1832
rect 2005 1787 2014 1799
rect 2005 1771 2011 1787
rect 1983 1764 1997 1771
rect 1883 1744 1887 1764
rect 1993 1744 1997 1764
rect 2003 1764 2011 1771
rect 2145 1779 2149 1828
rect 2199 1780 2203 1876
rect 2244 1837 2248 1876
rect 2264 1870 2268 1876
rect 2265 1840 2269 1858
rect 2284 1856 2288 1876
rect 2304 1870 2308 1876
rect 2304 1858 2309 1870
rect 2284 1850 2300 1856
rect 2244 1825 2245 1837
rect 2265 1834 2280 1840
rect 2244 1794 2248 1825
rect 2244 1788 2270 1794
rect 2145 1767 2154 1779
rect 2199 1768 2246 1780
rect 2003 1744 2007 1764
rect 2145 1752 2149 1767
rect 2125 1748 2149 1752
rect 2125 1744 2129 1748
rect 2145 1744 2149 1748
rect 2199 1724 2203 1768
rect 2266 1760 2270 1788
rect 2247 1756 2270 1760
rect 2276 1780 2280 1834
rect 2294 1812 2300 1850
rect 2276 1768 2278 1780
rect 2247 1744 2251 1756
rect 2276 1752 2280 1768
rect 2300 1760 2306 1800
rect 2259 1748 2280 1752
rect 2284 1756 2306 1760
rect 2259 1744 2263 1748
rect 2284 1744 2288 1756
rect 2315 1752 2320 1858
rect 2349 1807 2353 1896
rect 2369 1868 2373 1896
rect 2369 1856 2394 1868
rect 2336 1795 2350 1807
rect 2336 1762 2341 1795
rect 2370 1778 2375 1856
rect 2414 1818 2418 1876
rect 2296 1748 2320 1752
rect 2349 1772 2375 1778
rect 2406 1812 2418 1818
rect 2296 1744 2300 1748
rect 2349 1724 2353 1772
rect 2406 1762 2410 1812
rect 2434 1795 2438 1876
rect 2431 1783 2438 1795
rect 2406 1756 2414 1762
rect 2369 1724 2373 1750
rect 2414 1724 2418 1750
rect 2434 1744 2438 1783
rect 2479 1781 2483 1876
rect 2499 1811 2503 1896
rect 2479 1769 2488 1781
rect 2500 1777 2504 1799
rect 2519 1785 2523 1896
rect 2564 1821 2568 1876
rect 2584 1841 2588 1876
rect 2604 1858 2608 1876
rect 2500 1773 2528 1777
rect 2434 1732 2458 1744
rect 2434 1724 2438 1732
rect 2484 1724 2488 1769
rect 2504 1724 2508 1753
rect 2524 1724 2528 1773
rect 2564 1774 2568 1809
rect 2564 1770 2578 1774
rect 2574 1744 2578 1770
rect 2586 1744 2590 1829
rect 2602 1762 2606 1846
rect 2624 1799 2628 1876
rect 2711 1799 2715 1876
rect 2626 1787 2628 1799
rect 2706 1787 2715 1799
rect 2610 1744 2614 1750
rect 2622 1744 2626 1787
rect 2709 1771 2715 1787
rect 2731 1799 2735 1876
rect 2845 1833 2849 1876
rect 2865 1864 2869 1876
rect 2885 1868 2889 1876
rect 2885 1864 2900 1868
rect 2865 1860 2880 1864
rect 2874 1853 2880 1860
rect 2845 1821 2853 1833
rect 2865 1821 2872 1833
rect 2731 1787 2734 1799
rect 2731 1771 2737 1787
rect 2709 1764 2717 1771
rect 2713 1744 2717 1764
rect 2723 1764 2737 1771
rect 2868 1764 2872 1821
rect 2876 1764 2880 1841
rect 2894 1833 2900 1864
rect 2990 1833 2994 1876
rect 3231 1908 3235 1916
rect 3251 1908 3255 1912
rect 3261 1908 3265 1916
rect 3231 1864 3235 1868
rect 3223 1860 3235 1864
rect 2884 1821 2894 1833
rect 2987 1821 2994 1833
rect 2884 1764 2888 1821
rect 2723 1744 2727 1764
rect 2985 1744 2989 1821
rect 3012 1779 3016 1836
rect 3020 1832 3024 1836
rect 3020 1824 3038 1832
rect 3034 1813 3038 1824
rect 3111 1813 3115 1836
rect 3106 1801 3115 1813
rect 3119 1813 3123 1836
rect 3119 1801 3134 1813
rect 3005 1767 3014 1779
rect 3005 1744 3009 1767
rect 3034 1756 3038 1801
rect 3025 1749 3038 1756
rect 3025 1744 3029 1749
rect 3111 1724 3115 1801
rect 3131 1724 3135 1801
rect 3223 1779 3227 1860
rect 3251 1823 3255 1828
rect 3261 1824 3265 1828
rect 3242 1819 3255 1823
rect 3242 1813 3247 1819
rect 3281 1814 3285 1836
rect 3255 1810 3285 1814
rect 3291 1813 3295 1836
rect 3223 1741 3227 1767
rect 3241 1770 3246 1801
rect 3291 1801 3294 1813
rect 3241 1764 3255 1770
rect 3251 1752 3255 1764
rect 3261 1752 3265 1798
rect 3281 1752 3285 1756
rect 3291 1752 3295 1801
rect 3405 1793 3409 1876
rect 3491 1832 3495 1836
rect 3481 1828 3495 1832
rect 3501 1832 3505 1836
rect 3501 1828 3515 1832
rect 3481 1813 3486 1828
rect 3405 1781 3414 1793
rect 3223 1736 3235 1741
rect 3231 1732 3235 1736
rect 3405 1724 3409 1781
rect 3480 1755 3486 1801
rect 3509 1779 3515 1828
rect 3531 1779 3535 1836
rect 3541 1832 3545 1836
rect 3670 1833 3674 1876
rect 3541 1828 3555 1832
rect 3551 1813 3555 1828
rect 3667 1821 3674 1833
rect 3551 1801 3553 1813
rect 3506 1767 3515 1779
rect 3480 1751 3495 1755
rect 3491 1744 3495 1751
rect 3511 1744 3515 1767
rect 3531 1744 3535 1767
rect 3551 1744 3555 1801
rect 3665 1744 3669 1821
rect 3692 1779 3696 1836
rect 3700 1832 3704 1836
rect 3830 1833 3834 1876
rect 3700 1824 3718 1832
rect 3714 1813 3718 1824
rect 3827 1821 3834 1833
rect 3685 1767 3694 1779
rect 3685 1744 3689 1767
rect 3714 1756 3718 1801
rect 3705 1749 3718 1756
rect 3705 1744 3709 1749
rect 3825 1744 3829 1821
rect 3852 1779 3856 1836
rect 3860 1832 3864 1836
rect 3956 1832 3960 1836
rect 3860 1824 3878 1832
rect 3874 1813 3878 1824
rect 3942 1824 3960 1832
rect 3942 1813 3946 1824
rect 3845 1767 3854 1779
rect 3845 1744 3849 1767
rect 3874 1756 3878 1801
rect 3865 1749 3878 1756
rect 3942 1756 3946 1801
rect 3964 1779 3968 1836
rect 3986 1833 3990 1876
rect 3986 1821 3993 1833
rect 3966 1767 3975 1779
rect 3942 1749 3955 1756
rect 3865 1744 3869 1749
rect 3951 1744 3955 1749
rect 3971 1744 3975 1767
rect 3991 1744 3995 1821
rect 4105 1799 4109 1876
rect 4106 1787 4109 1799
rect 4103 1771 4109 1787
rect 4125 1799 4129 1876
rect 4225 1813 4229 1836
rect 4226 1801 4229 1813
rect 4125 1787 4134 1799
rect 4125 1771 4131 1787
rect 4103 1764 4117 1771
rect 4113 1744 4117 1764
rect 4123 1764 4131 1771
rect 4123 1744 4127 1764
rect 4220 1753 4226 1801
rect 4245 1779 4249 1836
rect 4265 1814 4269 1836
rect 4285 1814 4289 1836
rect 4265 1808 4278 1814
rect 4285 1813 4305 1814
rect 4285 1808 4293 1813
rect 4274 1779 4278 1808
rect 4247 1767 4249 1779
rect 4245 1765 4249 1767
rect 4245 1758 4258 1765
rect 4220 1749 4250 1753
rect 4246 1744 4250 1749
rect 4254 1744 4258 1758
rect 4274 1744 4278 1767
rect 4293 1759 4299 1801
rect 4385 1799 4389 1876
rect 4386 1787 4389 1799
rect 4383 1771 4389 1787
rect 4405 1799 4409 1876
rect 4496 1832 4500 1836
rect 4482 1824 4500 1832
rect 4482 1813 4486 1824
rect 4405 1787 4414 1799
rect 4405 1771 4411 1787
rect 4383 1764 4397 1771
rect 4282 1752 4299 1759
rect 4282 1744 4286 1752
rect 4393 1744 4397 1764
rect 4403 1764 4411 1771
rect 4403 1744 4407 1764
rect 4482 1756 4486 1801
rect 4504 1779 4508 1836
rect 4526 1833 4530 1876
rect 4526 1821 4533 1833
rect 4506 1767 4515 1779
rect 4482 1749 4495 1756
rect 4491 1744 4495 1749
rect 4511 1744 4515 1767
rect 4531 1744 4535 1821
rect 4641 1762 4645 1836
rect 4663 1799 4667 1876
rect 4685 1813 4689 1876
rect 4797 1813 4801 1836
rect 4685 1801 4694 1813
rect 4786 1801 4801 1813
rect 4805 1813 4809 1836
rect 4805 1801 4814 1813
rect 4666 1787 4679 1799
rect 4641 1750 4653 1762
rect 4655 1744 4659 1750
rect 4675 1744 4679 1787
rect 4685 1744 4689 1801
rect 3231 1704 3235 1712
rect 3251 1708 3255 1712
rect 3261 1708 3265 1712
rect 3281 1704 3285 1712
rect 3291 1708 3295 1712
rect 4785 1724 4789 1801
rect 4805 1724 4809 1801
rect 4905 1799 4909 1876
rect 4906 1787 4909 1799
rect 4903 1771 4909 1787
rect 4925 1799 4929 1876
rect 5025 1813 5029 1836
rect 5026 1801 5029 1813
rect 4925 1787 4934 1799
rect 4925 1771 4931 1787
rect 4903 1764 4917 1771
rect 4913 1744 4917 1764
rect 4923 1764 4931 1771
rect 4923 1744 4927 1764
rect 5020 1753 5026 1801
rect 5045 1779 5049 1836
rect 5065 1814 5069 1836
rect 5085 1814 5089 1836
rect 5065 1808 5078 1814
rect 5085 1813 5105 1814
rect 5085 1808 5093 1813
rect 5074 1779 5078 1808
rect 5047 1767 5049 1779
rect 5045 1765 5049 1767
rect 5045 1758 5058 1765
rect 5020 1749 5050 1753
rect 5046 1744 5050 1749
rect 5054 1744 5058 1758
rect 5074 1744 5078 1767
rect 5093 1759 5099 1801
rect 5082 1752 5099 1759
rect 5185 1793 5189 1876
rect 5297 1813 5301 1836
rect 5286 1801 5301 1813
rect 5305 1813 5309 1836
rect 5396 1832 5400 1836
rect 5382 1824 5400 1832
rect 5382 1813 5386 1824
rect 5305 1801 5314 1813
rect 5185 1781 5194 1793
rect 5082 1744 5086 1752
rect 5185 1724 5189 1781
rect 5285 1724 5289 1801
rect 5305 1724 5309 1801
rect 5382 1756 5386 1801
rect 5404 1779 5408 1836
rect 5426 1833 5430 1876
rect 5550 1833 5554 1876
rect 5426 1821 5433 1833
rect 5547 1821 5554 1833
rect 5406 1767 5415 1779
rect 5382 1749 5395 1756
rect 5391 1744 5395 1749
rect 5411 1744 5415 1767
rect 5431 1744 5435 1821
rect 5545 1744 5549 1821
rect 5572 1779 5576 1836
rect 5580 1832 5584 1836
rect 5671 1832 5675 1836
rect 5691 1832 5695 1836
rect 5580 1824 5598 1832
rect 5594 1813 5598 1824
rect 5671 1828 5695 1832
rect 5565 1767 5574 1779
rect 5565 1744 5569 1767
rect 5594 1756 5598 1801
rect 5671 1779 5675 1828
rect 5666 1767 5675 1779
rect 5585 1749 5598 1756
rect 5671 1752 5675 1767
rect 5585 1744 5589 1749
rect 5671 1748 5695 1752
rect 5671 1744 5675 1748
rect 5691 1744 5695 1748
rect 108 1700 112 1704
rect 116 1700 120 1704
rect 124 1700 128 1704
rect 214 1700 218 1704
rect 222 1700 226 1704
rect 244 1700 248 1704
rect 365 1700 369 1704
rect 385 1700 389 1704
rect 405 1700 409 1704
rect 528 1700 532 1704
rect 536 1700 540 1704
rect 544 1700 548 1704
rect 665 1700 669 1704
rect 685 1700 689 1704
rect 774 1700 778 1704
rect 782 1700 786 1704
rect 804 1700 808 1704
rect 945 1700 949 1704
rect 1065 1700 1069 1704
rect 1085 1700 1089 1704
rect 1105 1700 1109 1704
rect 1205 1700 1209 1704
rect 1225 1700 1229 1704
rect 1245 1700 1249 1704
rect 1345 1700 1349 1704
rect 1445 1700 1449 1704
rect 1465 1700 1469 1704
rect 1485 1700 1489 1704
rect 1571 1700 1575 1704
rect 1591 1700 1595 1704
rect 1611 1700 1615 1704
rect 1725 1700 1729 1704
rect 1745 1700 1749 1704
rect 1765 1700 1769 1704
rect 1873 1700 1877 1704
rect 1883 1700 1887 1704
rect 1993 1700 1997 1704
rect 2003 1700 2007 1704
rect 2125 1700 2129 1704
rect 2145 1700 2149 1704
rect 2199 1700 2203 1704
rect 2247 1700 2251 1704
rect 2259 1700 2263 1704
rect 2284 1700 2288 1704
rect 2296 1700 2300 1704
rect 2349 1700 2353 1704
rect 2369 1700 2373 1704
rect 2414 1700 2418 1704
rect 2434 1700 2438 1704
rect 2484 1700 2488 1704
rect 2504 1700 2508 1704
rect 2524 1700 2528 1704
rect 2574 1700 2578 1704
rect 2586 1700 2590 1704
rect 2610 1700 2614 1704
rect 2622 1700 2626 1704
rect 2713 1700 2717 1704
rect 2723 1700 2727 1704
rect 2868 1700 2872 1704
rect 2876 1700 2880 1704
rect 2884 1700 2888 1704
rect 2985 1700 2989 1704
rect 3005 1700 3009 1704
rect 3025 1700 3029 1704
rect 3111 1700 3115 1704
rect 3131 1700 3135 1704
rect 3231 1700 3285 1704
rect 3405 1700 3409 1704
rect 3491 1700 3495 1704
rect 3511 1700 3515 1704
rect 3531 1700 3535 1704
rect 3551 1700 3555 1704
rect 3665 1700 3669 1704
rect 3685 1700 3689 1704
rect 3705 1700 3709 1704
rect 3825 1700 3829 1704
rect 3845 1700 3849 1704
rect 3865 1700 3869 1704
rect 3951 1700 3955 1704
rect 3971 1700 3975 1704
rect 3991 1700 3995 1704
rect 4113 1700 4117 1704
rect 4123 1700 4127 1704
rect 4246 1700 4250 1704
rect 4254 1700 4258 1704
rect 4274 1700 4278 1704
rect 4282 1700 4286 1704
rect 4393 1700 4397 1704
rect 4403 1700 4407 1704
rect 4491 1700 4495 1704
rect 4511 1700 4515 1704
rect 4531 1700 4535 1704
rect 4655 1700 4659 1704
rect 4675 1700 4679 1704
rect 4685 1700 4689 1704
rect 4785 1700 4789 1704
rect 4805 1700 4809 1704
rect 4913 1700 4917 1704
rect 4923 1700 4927 1704
rect 5046 1700 5050 1704
rect 5054 1700 5058 1704
rect 5074 1700 5078 1704
rect 5082 1700 5086 1704
rect 5185 1700 5189 1704
rect 5285 1700 5289 1704
rect 5305 1700 5309 1704
rect 5391 1700 5395 1704
rect 5411 1700 5415 1704
rect 5431 1700 5435 1704
rect 5545 1700 5549 1704
rect 5565 1700 5569 1704
rect 5585 1700 5589 1704
rect 5671 1700 5675 1704
rect 5691 1700 5695 1704
rect 92 1676 96 1680
rect 100 1676 104 1680
rect 108 1676 112 1680
rect 268 1676 272 1680
rect 276 1676 280 1680
rect 284 1676 288 1680
rect 374 1676 378 1680
rect 382 1676 386 1680
rect 404 1676 408 1680
rect 532 1676 536 1680
rect 554 1676 558 1680
rect 562 1676 566 1680
rect 653 1676 657 1680
rect 663 1676 667 1680
rect 771 1676 775 1680
rect 885 1676 889 1680
rect 905 1676 909 1680
rect 925 1676 929 1680
rect 1048 1676 1052 1680
rect 1056 1676 1060 1680
rect 1064 1676 1068 1680
rect 1173 1676 1177 1680
rect 1183 1676 1187 1680
rect 1291 1676 1295 1680
rect 1311 1676 1315 1680
rect 1423 1676 1427 1680
rect 1445 1676 1449 1680
rect 1565 1676 1569 1680
rect 1654 1676 1658 1680
rect 1662 1676 1666 1680
rect 1682 1676 1686 1680
rect 1690 1676 1694 1680
rect 1779 1676 1783 1680
rect 1827 1676 1831 1680
rect 1839 1676 1843 1680
rect 1864 1676 1868 1680
rect 1876 1676 1880 1680
rect 1929 1676 1933 1680
rect 1949 1676 1953 1680
rect 1994 1676 1998 1680
rect 2014 1676 2018 1680
rect 2064 1676 2068 1680
rect 2084 1676 2088 1680
rect 2104 1676 2108 1680
rect 2154 1676 2158 1680
rect 2166 1676 2170 1680
rect 2190 1676 2194 1680
rect 2202 1676 2206 1680
rect 2311 1676 2315 1680
rect 2331 1676 2335 1680
rect 2351 1676 2355 1680
rect 2453 1676 2457 1680
rect 2463 1676 2467 1680
rect 2585 1676 2589 1680
rect 2605 1676 2609 1680
rect 2625 1676 2629 1680
rect 2733 1676 2737 1680
rect 2743 1676 2747 1680
rect 2845 1676 2849 1680
rect 2865 1676 2869 1680
rect 2885 1676 2889 1680
rect 2985 1676 2989 1680
rect 3005 1676 3009 1680
rect 3025 1676 3029 1680
rect 3074 1676 3078 1680
rect 3086 1676 3090 1680
rect 3110 1676 3114 1680
rect 3122 1676 3126 1680
rect 3172 1676 3176 1680
rect 3192 1676 3196 1680
rect 3212 1676 3216 1680
rect 3262 1676 3266 1680
rect 3282 1676 3286 1680
rect 3327 1676 3331 1680
rect 3347 1676 3351 1680
rect 3400 1676 3404 1680
rect 3412 1676 3416 1680
rect 3437 1676 3441 1680
rect 3449 1676 3453 1680
rect 3497 1676 3501 1680
rect 3612 1676 3616 1680
rect 3634 1676 3638 1680
rect 3642 1676 3646 1680
rect 3731 1676 3735 1680
rect 3751 1676 3755 1680
rect 3771 1676 3775 1680
rect 3883 1676 3887 1680
rect 3905 1676 3909 1680
rect 4015 1676 4019 1680
rect 4035 1676 4039 1680
rect 4045 1676 4049 1680
rect 4133 1676 4137 1680
rect 4143 1676 4147 1680
rect 4286 1676 4290 1680
rect 4294 1676 4298 1680
rect 4314 1676 4318 1680
rect 4322 1676 4326 1680
rect 4446 1676 4450 1680
rect 4454 1676 4458 1680
rect 4474 1676 4478 1680
rect 4482 1676 4486 1680
rect 4594 1676 4598 1680
rect 4602 1676 4606 1680
rect 4622 1676 4626 1680
rect 4630 1676 4634 1680
rect 4753 1676 4757 1680
rect 4763 1676 4767 1680
rect 4871 1676 4875 1680
rect 4891 1676 4895 1680
rect 4911 1676 4915 1680
rect 5035 1676 5039 1680
rect 5055 1676 5059 1680
rect 5065 1676 5069 1680
rect 5172 1676 5176 1680
rect 5180 1676 5184 1680
rect 5188 1676 5192 1680
rect 5314 1676 5318 1680
rect 5322 1676 5326 1680
rect 5342 1676 5346 1680
rect 5350 1676 5354 1680
rect 5473 1676 5477 1680
rect 5483 1676 5487 1680
rect 5592 1676 5596 1680
rect 5600 1676 5604 1680
rect 5608 1676 5612 1680
rect 5765 1676 5769 1680
rect 374 1632 378 1636
rect 359 1626 378 1632
rect 92 1559 96 1616
rect 86 1547 96 1559
rect 80 1516 86 1547
rect 100 1539 104 1616
rect 108 1559 112 1616
rect 268 1559 272 1616
rect 108 1547 115 1559
rect 127 1547 135 1559
rect 100 1520 106 1527
rect 100 1516 115 1520
rect 80 1512 95 1516
rect 91 1504 95 1512
rect 111 1504 115 1516
rect 131 1504 135 1547
rect 245 1547 253 1559
rect 265 1547 272 1559
rect 245 1504 249 1547
rect 276 1539 280 1616
rect 284 1559 288 1616
rect 359 1613 366 1626
rect 359 1564 366 1601
rect 382 1599 386 1636
rect 404 1613 408 1656
rect 532 1613 536 1656
rect 406 1601 415 1613
rect 380 1564 386 1587
rect 284 1547 294 1559
rect 359 1558 375 1564
rect 380 1558 395 1564
rect 274 1520 280 1527
rect 265 1516 280 1520
rect 294 1516 300 1547
rect 371 1544 375 1558
rect 391 1544 395 1558
rect 411 1544 415 1601
rect 525 1601 534 1613
rect 525 1544 529 1601
rect 554 1599 558 1636
rect 562 1632 566 1636
rect 562 1626 581 1632
rect 574 1613 581 1626
rect 653 1616 657 1636
rect 649 1609 657 1616
rect 663 1616 667 1636
rect 663 1609 677 1616
rect 554 1564 560 1587
rect 574 1564 581 1601
rect 649 1593 655 1609
rect 646 1581 655 1593
rect 545 1558 560 1564
rect 565 1558 581 1564
rect 545 1544 549 1558
rect 565 1544 569 1558
rect 265 1504 269 1516
rect 285 1512 300 1516
rect 285 1504 289 1512
rect 651 1504 655 1581
rect 671 1593 677 1609
rect 771 1599 775 1656
rect 671 1581 674 1593
rect 766 1587 775 1599
rect 671 1504 675 1581
rect 771 1504 775 1587
rect 885 1559 889 1636
rect 905 1613 909 1636
rect 925 1631 929 1636
rect 925 1624 938 1631
rect 905 1601 914 1613
rect 887 1547 894 1559
rect 890 1504 894 1547
rect 912 1544 916 1601
rect 934 1579 938 1624
rect 1173 1616 1177 1636
rect 934 1556 938 1567
rect 1048 1559 1052 1616
rect 920 1548 938 1556
rect 920 1544 924 1548
rect 1025 1547 1033 1559
rect 1045 1547 1052 1559
rect 1025 1504 1029 1547
rect 1056 1539 1060 1616
rect 1064 1559 1068 1616
rect 1163 1609 1177 1616
rect 1183 1616 1187 1636
rect 1183 1609 1191 1616
rect 1163 1593 1169 1609
rect 1166 1581 1169 1593
rect 1064 1547 1074 1559
rect 1054 1520 1060 1527
rect 1045 1516 1060 1520
rect 1074 1516 1080 1547
rect 1045 1504 1049 1516
rect 1065 1512 1080 1516
rect 1065 1504 1069 1512
rect 1165 1504 1169 1581
rect 1185 1593 1191 1609
rect 1185 1581 1194 1593
rect 1185 1504 1189 1581
rect 1291 1579 1295 1656
rect 1311 1579 1315 1656
rect 1423 1630 1427 1636
rect 1423 1618 1425 1630
rect 1445 1579 1449 1656
rect 1565 1599 1569 1656
rect 1654 1628 1658 1636
rect 1641 1621 1658 1628
rect 1565 1587 1574 1599
rect 1286 1567 1295 1579
rect 1291 1544 1295 1567
rect 1299 1567 1314 1579
rect 1445 1567 1454 1579
rect 1299 1544 1303 1567
rect 1423 1550 1425 1562
rect 1423 1544 1427 1550
rect 1445 1504 1449 1567
rect 1565 1504 1569 1587
rect 1641 1579 1647 1621
rect 1662 1613 1666 1636
rect 1682 1622 1686 1636
rect 1690 1631 1694 1636
rect 1690 1627 1720 1631
rect 1682 1615 1695 1622
rect 1691 1613 1695 1615
rect 1691 1601 1693 1613
rect 1662 1572 1666 1601
rect 1647 1567 1655 1572
rect 1635 1566 1655 1567
rect 1662 1566 1675 1572
rect 1651 1544 1655 1566
rect 1671 1544 1675 1566
rect 1691 1544 1695 1601
rect 1714 1579 1720 1627
rect 1779 1612 1783 1656
rect 1827 1624 1831 1636
rect 1839 1632 1843 1636
rect 1839 1628 1860 1632
rect 1827 1620 1850 1624
rect 1779 1600 1826 1612
rect 1711 1567 1714 1579
rect 1711 1544 1715 1567
rect 1779 1504 1783 1600
rect 1846 1592 1850 1620
rect 1824 1586 1850 1592
rect 1856 1612 1860 1628
rect 1864 1624 1868 1636
rect 1876 1632 1880 1636
rect 1876 1628 1900 1632
rect 1864 1620 1886 1624
rect 1856 1600 1858 1612
rect 1824 1555 1828 1586
rect 1824 1543 1825 1555
rect 1856 1546 1860 1600
rect 1880 1580 1886 1620
rect 1824 1504 1828 1543
rect 1845 1540 1860 1546
rect 1845 1522 1849 1540
rect 1874 1530 1880 1568
rect 1864 1524 1880 1530
rect 1844 1504 1848 1510
rect 1864 1504 1868 1524
rect 1895 1522 1900 1628
rect 1916 1585 1921 1618
rect 1929 1608 1933 1656
rect 1949 1630 1953 1656
rect 1994 1630 1998 1656
rect 2014 1648 2018 1656
rect 2014 1636 2038 1648
rect 1986 1618 1994 1624
rect 1929 1602 1955 1608
rect 1916 1573 1930 1585
rect 1884 1510 1889 1522
rect 1884 1504 1888 1510
rect 1929 1484 1933 1573
rect 1950 1524 1955 1602
rect 1986 1568 1990 1618
rect 2014 1597 2018 1636
rect 2064 1611 2068 1656
rect 2084 1627 2088 1656
rect 2059 1599 2068 1611
rect 2104 1607 2108 1656
rect 2154 1610 2158 1636
rect 2080 1603 2108 1607
rect 2144 1606 2158 1610
rect 2011 1585 2018 1597
rect 1986 1562 1998 1568
rect 1949 1512 1974 1524
rect 1949 1484 1953 1512
rect 1994 1504 1998 1562
rect 2014 1504 2018 1585
rect 2059 1504 2063 1599
rect 2080 1581 2084 1603
rect 2079 1484 2083 1569
rect 2099 1484 2103 1595
rect 2144 1571 2148 1606
rect 2144 1504 2148 1559
rect 2166 1551 2170 1636
rect 2190 1630 2194 1636
rect 2164 1504 2168 1539
rect 2182 1534 2186 1618
rect 2202 1593 2206 1636
rect 2311 1631 2315 1636
rect 2302 1624 2315 1631
rect 2206 1581 2208 1593
rect 2184 1504 2188 1522
rect 2204 1504 2208 1581
rect 2302 1579 2306 1624
rect 2331 1613 2335 1636
rect 2326 1601 2335 1613
rect 2302 1556 2306 1567
rect 2302 1548 2320 1556
rect 2316 1544 2320 1548
rect 2324 1544 2328 1601
rect 2351 1559 2355 1636
rect 2453 1616 2457 1636
rect 2449 1609 2457 1616
rect 2463 1616 2467 1636
rect 2463 1609 2477 1616
rect 2449 1593 2455 1609
rect 2446 1581 2455 1593
rect 2346 1547 2353 1559
rect 2346 1504 2350 1547
rect 2451 1504 2455 1581
rect 2471 1593 2477 1609
rect 2471 1581 2474 1593
rect 2471 1504 2475 1581
rect 2585 1559 2589 1636
rect 2605 1613 2609 1636
rect 2625 1631 2629 1636
rect 2625 1624 2638 1631
rect 2605 1601 2614 1613
rect 2587 1547 2594 1559
rect 2590 1504 2594 1547
rect 2612 1544 2616 1601
rect 2634 1579 2638 1624
rect 2733 1616 2737 1636
rect 2723 1609 2737 1616
rect 2743 1616 2747 1636
rect 2743 1609 2751 1616
rect 2723 1593 2729 1609
rect 2726 1581 2729 1593
rect 2634 1556 2638 1567
rect 2620 1548 2638 1556
rect 2620 1544 2624 1548
rect 2725 1504 2729 1581
rect 2745 1593 2751 1609
rect 2745 1581 2754 1593
rect 2745 1504 2749 1581
rect 2845 1559 2849 1636
rect 2865 1613 2869 1636
rect 2885 1631 2889 1636
rect 2885 1624 2898 1631
rect 2865 1601 2874 1613
rect 2847 1547 2854 1559
rect 2850 1504 2854 1547
rect 2872 1544 2876 1601
rect 2894 1579 2898 1624
rect 2894 1556 2898 1567
rect 2985 1559 2989 1636
rect 3005 1613 3009 1636
rect 3025 1631 3029 1636
rect 3025 1624 3038 1631
rect 3005 1601 3014 1613
rect 2880 1548 2898 1556
rect 2880 1544 2884 1548
rect 2987 1547 2994 1559
rect 2990 1504 2994 1547
rect 3012 1544 3016 1601
rect 3034 1579 3038 1624
rect 3074 1593 3078 1636
rect 3086 1630 3090 1636
rect 3072 1581 3074 1593
rect 3034 1556 3038 1567
rect 3020 1548 3038 1556
rect 3020 1544 3024 1548
rect 3072 1504 3076 1581
rect 3094 1534 3098 1618
rect 3110 1551 3114 1636
rect 3122 1610 3126 1636
rect 3122 1606 3136 1610
rect 3132 1571 3136 1606
rect 3172 1607 3176 1656
rect 3192 1627 3196 1656
rect 3212 1611 3216 1656
rect 3262 1648 3266 1656
rect 3242 1636 3266 1648
rect 3172 1603 3200 1607
rect 3092 1504 3096 1522
rect 3112 1504 3116 1539
rect 3132 1504 3136 1559
rect 3177 1484 3181 1595
rect 3196 1581 3200 1603
rect 3212 1599 3221 1611
rect 3197 1484 3201 1569
rect 3217 1504 3221 1599
rect 3262 1597 3266 1636
rect 3282 1630 3286 1656
rect 3327 1630 3331 1656
rect 3286 1618 3294 1624
rect 3262 1585 3269 1597
rect 3262 1504 3266 1585
rect 3290 1568 3294 1618
rect 3347 1608 3351 1656
rect 3400 1632 3404 1636
rect 3282 1562 3294 1568
rect 3325 1602 3351 1608
rect 3380 1628 3404 1632
rect 3282 1504 3286 1562
rect 3325 1524 3330 1602
rect 3359 1585 3364 1618
rect 3350 1573 3364 1585
rect 3306 1512 3331 1524
rect 3327 1484 3331 1512
rect 3347 1484 3351 1573
rect 3380 1522 3385 1628
rect 3412 1624 3416 1636
rect 3437 1632 3441 1636
rect 3394 1620 3416 1624
rect 3420 1628 3441 1632
rect 3394 1580 3400 1620
rect 3420 1612 3424 1628
rect 3449 1624 3453 1636
rect 3422 1600 3424 1612
rect 3400 1530 3406 1568
rect 3420 1546 3424 1600
rect 3430 1620 3453 1624
rect 3430 1592 3434 1620
rect 3497 1612 3501 1656
rect 3612 1613 3616 1656
rect 3454 1600 3501 1612
rect 3430 1586 3456 1592
rect 3452 1555 3456 1586
rect 3420 1540 3435 1546
rect 3455 1543 3456 1555
rect 3400 1524 3416 1530
rect 3391 1510 3396 1522
rect 3392 1504 3396 1510
rect 3412 1504 3416 1524
rect 3431 1522 3435 1540
rect 3432 1504 3436 1510
rect 3452 1504 3456 1543
rect 3497 1504 3501 1600
rect 3605 1601 3614 1613
rect 3605 1544 3609 1601
rect 3634 1599 3638 1636
rect 3642 1632 3646 1636
rect 3642 1626 3661 1632
rect 3731 1631 3735 1636
rect 3654 1613 3661 1626
rect 3722 1624 3735 1631
rect 3634 1564 3640 1587
rect 3654 1564 3661 1601
rect 3722 1579 3726 1624
rect 3751 1613 3755 1636
rect 3746 1601 3755 1613
rect 3625 1558 3640 1564
rect 3645 1558 3661 1564
rect 3625 1544 3629 1558
rect 3645 1544 3649 1558
rect 3722 1556 3726 1567
rect 3722 1548 3740 1556
rect 3736 1544 3740 1548
rect 3744 1544 3748 1601
rect 3771 1559 3775 1636
rect 3883 1630 3887 1636
rect 3883 1618 3885 1630
rect 3905 1579 3909 1656
rect 4015 1630 4019 1636
rect 4001 1618 4013 1630
rect 3905 1567 3914 1579
rect 3766 1547 3773 1559
rect 3883 1550 3885 1562
rect 3766 1504 3770 1547
rect 3883 1544 3887 1550
rect 3905 1504 3909 1567
rect 4001 1544 4005 1618
rect 4035 1593 4039 1636
rect 4026 1581 4039 1593
rect 4023 1504 4027 1581
rect 4045 1579 4049 1636
rect 4133 1616 4137 1636
rect 4129 1609 4137 1616
rect 4143 1616 4147 1636
rect 4286 1631 4290 1636
rect 4260 1627 4290 1631
rect 4143 1609 4157 1616
rect 4129 1593 4135 1609
rect 4126 1581 4135 1593
rect 4045 1567 4054 1579
rect 4045 1504 4049 1567
rect 4131 1504 4135 1581
rect 4151 1593 4157 1609
rect 4151 1581 4154 1593
rect 4151 1504 4155 1581
rect 4260 1579 4266 1627
rect 4294 1622 4298 1636
rect 4285 1615 4298 1622
rect 4285 1613 4289 1615
rect 4314 1613 4318 1636
rect 4322 1628 4326 1636
rect 4446 1631 4450 1636
rect 4322 1621 4339 1628
rect 4287 1601 4289 1613
rect 4266 1567 4269 1579
rect 4265 1544 4269 1567
rect 4285 1544 4289 1601
rect 4314 1572 4318 1601
rect 4333 1579 4339 1621
rect 4420 1627 4450 1631
rect 4420 1579 4426 1627
rect 4454 1622 4458 1636
rect 4445 1615 4458 1622
rect 4445 1613 4449 1615
rect 4474 1613 4478 1636
rect 4482 1628 4486 1636
rect 4594 1628 4598 1636
rect 4482 1621 4499 1628
rect 4447 1601 4449 1613
rect 4305 1566 4318 1572
rect 4325 1567 4333 1572
rect 4426 1567 4429 1579
rect 4325 1566 4345 1567
rect 4305 1544 4309 1566
rect 4325 1544 4329 1566
rect 4425 1544 4429 1567
rect 4445 1544 4449 1601
rect 4474 1572 4478 1601
rect 4493 1579 4499 1621
rect 4581 1621 4598 1628
rect 4581 1579 4587 1621
rect 4602 1613 4606 1636
rect 4622 1622 4626 1636
rect 4630 1631 4634 1636
rect 4630 1627 4660 1631
rect 4622 1615 4635 1622
rect 4631 1613 4635 1615
rect 4631 1601 4633 1613
rect 4465 1566 4478 1572
rect 4485 1567 4493 1572
rect 4485 1566 4505 1567
rect 4602 1572 4606 1601
rect 4587 1567 4595 1572
rect 4575 1566 4595 1567
rect 4602 1566 4615 1572
rect 4465 1544 4469 1566
rect 4485 1544 4489 1566
rect 4591 1544 4595 1566
rect 4611 1544 4615 1566
rect 4631 1544 4635 1601
rect 4654 1579 4660 1627
rect 4753 1616 4757 1636
rect 4749 1609 4757 1616
rect 4763 1616 4767 1636
rect 4871 1631 4875 1636
rect 4862 1624 4875 1631
rect 4763 1609 4777 1616
rect 4749 1593 4755 1609
rect 4746 1581 4755 1593
rect 4651 1567 4654 1579
rect 4651 1544 4655 1567
rect 4751 1504 4755 1581
rect 4771 1593 4777 1609
rect 4771 1581 4774 1593
rect 4771 1504 4775 1581
rect 4862 1579 4866 1624
rect 4891 1613 4895 1636
rect 4886 1601 4895 1613
rect 4862 1556 4866 1567
rect 4862 1548 4880 1556
rect 4876 1544 4880 1548
rect 4884 1544 4888 1601
rect 4911 1559 4915 1636
rect 5035 1630 5039 1636
rect 5021 1618 5033 1630
rect 4906 1547 4913 1559
rect 4906 1504 4910 1547
rect 5021 1544 5025 1618
rect 5055 1593 5059 1636
rect 5046 1581 5059 1593
rect 5043 1504 5047 1581
rect 5065 1579 5069 1636
rect 5314 1628 5318 1636
rect 5301 1621 5318 1628
rect 5065 1567 5074 1579
rect 5065 1504 5069 1567
rect 5172 1559 5176 1616
rect 5166 1547 5176 1559
rect 5160 1516 5166 1547
rect 5180 1539 5184 1616
rect 5188 1559 5192 1616
rect 5301 1579 5307 1621
rect 5322 1613 5326 1636
rect 5342 1622 5346 1636
rect 5350 1631 5354 1636
rect 5350 1627 5380 1631
rect 5342 1615 5355 1622
rect 5351 1613 5355 1615
rect 5351 1601 5353 1613
rect 5322 1572 5326 1601
rect 5307 1567 5315 1572
rect 5295 1566 5315 1567
rect 5322 1566 5335 1572
rect 5188 1547 5195 1559
rect 5207 1547 5215 1559
rect 5180 1520 5186 1527
rect 5180 1516 5195 1520
rect 5160 1512 5175 1516
rect 5171 1504 5175 1512
rect 5191 1504 5195 1516
rect 5211 1504 5215 1547
rect 5311 1544 5315 1566
rect 5331 1544 5335 1566
rect 5351 1544 5355 1601
rect 5374 1579 5380 1627
rect 5473 1616 5477 1636
rect 5469 1609 5477 1616
rect 5483 1616 5487 1636
rect 5483 1609 5497 1616
rect 5469 1593 5475 1609
rect 5466 1581 5475 1593
rect 5371 1567 5374 1579
rect 5371 1544 5375 1567
rect 5471 1504 5475 1581
rect 5491 1593 5497 1609
rect 5491 1581 5494 1593
rect 5491 1504 5495 1581
rect 5592 1559 5596 1616
rect 5586 1547 5596 1559
rect 5580 1516 5586 1547
rect 5600 1539 5604 1616
rect 5608 1559 5612 1616
rect 5765 1613 5769 1636
rect 5765 1601 5774 1613
rect 5608 1547 5615 1559
rect 5627 1547 5635 1559
rect 5600 1520 5606 1527
rect 5600 1516 5615 1520
rect 5580 1512 5595 1516
rect 5591 1504 5595 1512
rect 5611 1504 5615 1516
rect 5631 1504 5635 1547
rect 5765 1544 5769 1601
rect 91 1460 95 1464
rect 111 1460 115 1464
rect 131 1460 135 1464
rect 245 1460 249 1464
rect 265 1460 269 1464
rect 285 1460 289 1464
rect 371 1460 375 1464
rect 391 1460 395 1464
rect 411 1460 415 1464
rect 525 1460 529 1464
rect 545 1460 549 1464
rect 565 1460 569 1464
rect 651 1460 655 1464
rect 671 1460 675 1464
rect 771 1460 775 1464
rect 890 1460 894 1464
rect 912 1460 916 1464
rect 920 1460 924 1464
rect 1025 1460 1029 1464
rect 1045 1460 1049 1464
rect 1065 1460 1069 1464
rect 1165 1460 1169 1464
rect 1185 1460 1189 1464
rect 1291 1460 1295 1464
rect 1299 1460 1303 1464
rect 1423 1460 1427 1464
rect 1445 1460 1449 1464
rect 1565 1460 1569 1464
rect 1651 1460 1655 1464
rect 1671 1460 1675 1464
rect 1691 1460 1695 1464
rect 1711 1460 1715 1464
rect 1779 1460 1783 1464
rect 1824 1460 1828 1464
rect 1844 1460 1848 1464
rect 1864 1460 1868 1464
rect 1884 1460 1888 1464
rect 1929 1460 1933 1464
rect 1949 1460 1953 1464
rect 1994 1460 1998 1464
rect 2014 1460 2018 1464
rect 2059 1460 2063 1464
rect 2079 1460 2083 1464
rect 2099 1460 2103 1464
rect 2144 1460 2148 1464
rect 2164 1460 2168 1464
rect 2184 1460 2188 1464
rect 2204 1460 2208 1464
rect 2316 1460 2320 1464
rect 2324 1460 2328 1464
rect 2346 1460 2350 1464
rect 2451 1460 2455 1464
rect 2471 1460 2475 1464
rect 2590 1460 2594 1464
rect 2612 1460 2616 1464
rect 2620 1460 2624 1464
rect 2725 1460 2729 1464
rect 2745 1460 2749 1464
rect 2850 1460 2854 1464
rect 2872 1460 2876 1464
rect 2880 1460 2884 1464
rect 2990 1460 2994 1464
rect 3012 1460 3016 1464
rect 3020 1460 3024 1464
rect 3072 1460 3076 1464
rect 3092 1460 3096 1464
rect 3112 1460 3116 1464
rect 3132 1460 3136 1464
rect 3177 1460 3181 1464
rect 3197 1460 3201 1464
rect 3217 1460 3221 1464
rect 3262 1460 3266 1464
rect 3282 1460 3286 1464
rect 3327 1460 3331 1464
rect 3347 1460 3351 1464
rect 3392 1460 3396 1464
rect 3412 1460 3416 1464
rect 3432 1460 3436 1464
rect 3452 1460 3456 1464
rect 3497 1460 3501 1464
rect 3605 1460 3609 1464
rect 3625 1460 3629 1464
rect 3645 1460 3649 1464
rect 3736 1460 3740 1464
rect 3744 1460 3748 1464
rect 3766 1460 3770 1464
rect 3883 1460 3887 1464
rect 3905 1460 3909 1464
rect 4001 1460 4005 1464
rect 4023 1460 4027 1464
rect 4045 1460 4049 1464
rect 4131 1460 4135 1464
rect 4151 1460 4155 1464
rect 4265 1460 4269 1464
rect 4285 1460 4289 1464
rect 4305 1460 4309 1464
rect 4325 1460 4329 1464
rect 4425 1460 4429 1464
rect 4445 1460 4449 1464
rect 4465 1460 4469 1464
rect 4485 1460 4489 1464
rect 4591 1460 4595 1464
rect 4611 1460 4615 1464
rect 4631 1460 4635 1464
rect 4651 1460 4655 1464
rect 4751 1460 4755 1464
rect 4771 1460 4775 1464
rect 4876 1460 4880 1464
rect 4884 1460 4888 1464
rect 4906 1460 4910 1464
rect 5021 1460 5025 1464
rect 5043 1460 5047 1464
rect 5065 1460 5069 1464
rect 5171 1460 5175 1464
rect 5191 1460 5195 1464
rect 5211 1460 5215 1464
rect 5311 1460 5315 1464
rect 5331 1460 5335 1464
rect 5351 1460 5355 1464
rect 5371 1460 5375 1464
rect 5471 1460 5475 1464
rect 5491 1460 5495 1464
rect 5591 1460 5595 1464
rect 5611 1460 5615 1464
rect 5631 1460 5635 1464
rect 5765 1460 5769 1464
rect 85 1436 89 1440
rect 105 1436 109 1440
rect 125 1436 129 1440
rect 211 1436 215 1440
rect 231 1436 235 1440
rect 251 1436 255 1440
rect 365 1436 369 1440
rect 385 1436 389 1440
rect 405 1436 409 1440
rect 510 1436 514 1440
rect 532 1436 536 1440
rect 540 1436 544 1440
rect 650 1436 654 1440
rect 672 1436 676 1440
rect 680 1436 684 1440
rect 801 1436 805 1440
rect 823 1436 827 1440
rect 845 1436 849 1440
rect 931 1436 935 1440
rect 951 1436 955 1440
rect 1065 1436 1069 1440
rect 1151 1436 1155 1440
rect 1171 1436 1175 1440
rect 1191 1436 1195 1440
rect 1291 1436 1295 1440
rect 1311 1436 1315 1440
rect 1425 1436 1429 1440
rect 1445 1436 1449 1440
rect 1545 1436 1549 1440
rect 1565 1436 1569 1440
rect 1685 1436 1689 1440
rect 1705 1436 1709 1440
rect 1725 1436 1729 1440
rect 1811 1436 1815 1440
rect 1831 1436 1835 1440
rect 1945 1436 1949 1440
rect 1965 1436 1969 1440
rect 1985 1436 1989 1440
rect 2085 1436 2089 1440
rect 2205 1436 2209 1440
rect 2225 1436 2229 1440
rect 2245 1436 2249 1440
rect 2345 1436 2349 1440
rect 2365 1436 2369 1440
rect 2385 1436 2389 1440
rect 2471 1436 2475 1440
rect 2610 1436 2614 1440
rect 2632 1436 2636 1440
rect 2640 1436 2644 1440
rect 2731 1436 2735 1440
rect 2751 1436 2755 1440
rect 2771 1436 2775 1440
rect 2890 1436 2894 1440
rect 2912 1436 2916 1440
rect 2920 1436 2924 1440
rect 3030 1436 3034 1440
rect 3052 1436 3056 1440
rect 3060 1436 3064 1440
rect 3170 1436 3174 1440
rect 3192 1436 3196 1440
rect 3200 1436 3204 1440
rect 3305 1436 3309 1440
rect 3391 1436 3395 1440
rect 3503 1436 3507 1440
rect 3525 1436 3529 1440
rect 3645 1436 3649 1440
rect 3665 1436 3669 1440
rect 3685 1436 3689 1440
rect 3776 1436 3780 1440
rect 3784 1436 3788 1440
rect 3806 1436 3810 1440
rect 3925 1436 3929 1440
rect 4030 1436 4034 1440
rect 4052 1436 4056 1440
rect 4060 1436 4064 1440
rect 4170 1436 4174 1440
rect 4192 1436 4196 1440
rect 4200 1436 4204 1440
rect 4305 1436 4309 1440
rect 4325 1436 4329 1440
rect 4345 1436 4349 1440
rect 4450 1436 4454 1440
rect 4472 1436 4476 1440
rect 4480 1436 4484 1440
rect 4596 1436 4600 1440
rect 4604 1436 4608 1440
rect 4626 1436 4630 1440
rect 4731 1436 4735 1440
rect 4751 1436 4755 1440
rect 4856 1436 4860 1440
rect 4864 1436 4868 1440
rect 4886 1436 4890 1440
rect 4991 1436 4995 1440
rect 4999 1436 5003 1440
rect 5111 1436 5115 1440
rect 5131 1436 5135 1440
rect 5245 1436 5249 1440
rect 5265 1436 5269 1440
rect 5370 1436 5374 1440
rect 5392 1436 5396 1440
rect 5400 1436 5404 1440
rect 5496 1436 5500 1440
rect 5504 1436 5508 1440
rect 5526 1436 5530 1440
rect 5656 1436 5660 1440
rect 5664 1436 5668 1440
rect 5686 1436 5690 1440
rect 85 1353 89 1396
rect 105 1384 109 1396
rect 125 1388 129 1396
rect 125 1384 140 1388
rect 105 1380 120 1384
rect 114 1373 120 1380
rect 85 1341 93 1353
rect 105 1341 112 1353
rect 108 1284 112 1341
rect 116 1284 120 1361
rect 134 1353 140 1384
rect 124 1341 134 1353
rect 211 1342 215 1356
rect 231 1342 235 1356
rect 124 1284 128 1341
rect 199 1336 215 1342
rect 220 1336 235 1342
rect 199 1299 206 1336
rect 220 1313 226 1336
rect 199 1274 206 1287
rect 199 1268 218 1274
rect 214 1264 218 1268
rect 222 1264 226 1301
rect 251 1299 255 1356
rect 365 1353 369 1396
rect 385 1384 389 1396
rect 405 1388 409 1396
rect 405 1384 420 1388
rect 385 1380 400 1384
rect 394 1373 400 1380
rect 365 1341 373 1353
rect 385 1341 392 1353
rect 246 1287 255 1299
rect 244 1244 248 1287
rect 388 1284 392 1341
rect 396 1284 400 1361
rect 414 1353 420 1384
rect 510 1353 514 1396
rect 404 1341 414 1353
rect 507 1341 514 1353
rect 404 1284 408 1341
rect 505 1264 509 1341
rect 532 1299 536 1356
rect 540 1352 544 1356
rect 650 1353 654 1396
rect 540 1344 558 1352
rect 554 1333 558 1344
rect 647 1341 654 1353
rect 525 1287 534 1299
rect 525 1264 529 1287
rect 554 1276 558 1321
rect 545 1269 558 1276
rect 545 1264 549 1269
rect 645 1264 649 1341
rect 672 1299 676 1356
rect 680 1352 684 1356
rect 680 1344 698 1352
rect 694 1333 698 1344
rect 665 1287 674 1299
rect 665 1264 669 1287
rect 694 1276 698 1321
rect 685 1269 698 1276
rect 801 1282 805 1356
rect 823 1319 827 1396
rect 845 1333 849 1396
rect 845 1321 854 1333
rect 826 1307 839 1319
rect 801 1270 813 1282
rect 685 1264 689 1269
rect 815 1264 819 1270
rect 835 1264 839 1307
rect 845 1264 849 1321
rect 931 1319 935 1396
rect 926 1307 935 1319
rect 929 1291 935 1307
rect 951 1319 955 1396
rect 951 1307 954 1319
rect 1065 1313 1069 1396
rect 1151 1388 1155 1396
rect 1140 1384 1155 1388
rect 1171 1384 1175 1396
rect 1140 1353 1146 1384
rect 1160 1380 1175 1384
rect 1160 1373 1166 1380
rect 1146 1341 1156 1353
rect 951 1291 957 1307
rect 929 1284 937 1291
rect 933 1264 937 1284
rect 943 1284 957 1291
rect 1065 1301 1074 1313
rect 943 1264 947 1284
rect 1065 1244 1069 1301
rect 1152 1284 1156 1341
rect 1160 1284 1164 1361
rect 1191 1353 1195 1396
rect 1168 1341 1175 1353
rect 1187 1341 1195 1353
rect 1168 1284 1172 1341
rect 1291 1319 1295 1396
rect 1286 1307 1295 1319
rect 1289 1291 1295 1307
rect 1311 1319 1315 1396
rect 1425 1319 1429 1396
rect 1311 1307 1314 1319
rect 1426 1307 1429 1319
rect 1311 1291 1317 1307
rect 1289 1284 1297 1291
rect 1293 1264 1297 1284
rect 1303 1284 1317 1291
rect 1423 1291 1429 1307
rect 1445 1319 1449 1396
rect 1545 1319 1549 1396
rect 1445 1307 1454 1319
rect 1546 1307 1549 1319
rect 1445 1291 1451 1307
rect 1423 1284 1437 1291
rect 1303 1264 1307 1284
rect 1433 1264 1437 1284
rect 1443 1284 1451 1291
rect 1543 1291 1549 1307
rect 1565 1319 1569 1396
rect 1685 1353 1689 1396
rect 1705 1384 1709 1396
rect 1725 1388 1729 1396
rect 1725 1384 1740 1388
rect 1705 1380 1720 1384
rect 1714 1373 1720 1380
rect 1685 1341 1693 1353
rect 1705 1341 1712 1353
rect 1565 1307 1574 1319
rect 1565 1291 1571 1307
rect 1543 1284 1557 1291
rect 1443 1264 1447 1284
rect 1553 1264 1557 1284
rect 1563 1284 1571 1291
rect 1708 1284 1712 1341
rect 1716 1284 1720 1361
rect 1734 1353 1740 1384
rect 1724 1341 1734 1353
rect 1724 1284 1728 1341
rect 1811 1319 1815 1396
rect 1806 1307 1815 1319
rect 1809 1291 1815 1307
rect 1831 1319 1835 1396
rect 1945 1353 1949 1396
rect 1965 1384 1969 1396
rect 1985 1388 1989 1396
rect 1985 1384 2000 1388
rect 1965 1380 1980 1384
rect 1974 1373 1980 1380
rect 1945 1341 1953 1353
rect 1965 1341 1972 1353
rect 1831 1307 1834 1319
rect 1831 1291 1837 1307
rect 1809 1284 1817 1291
rect 1563 1264 1567 1284
rect 1813 1264 1817 1284
rect 1823 1284 1837 1291
rect 1968 1284 1972 1341
rect 1976 1284 1980 1361
rect 1994 1353 2000 1384
rect 1984 1341 1994 1353
rect 1984 1284 1988 1341
rect 2085 1313 2089 1396
rect 2205 1353 2209 1396
rect 2225 1384 2229 1396
rect 2245 1388 2249 1396
rect 2245 1384 2260 1388
rect 2225 1380 2240 1384
rect 2234 1373 2240 1380
rect 2205 1341 2213 1353
rect 2225 1341 2232 1353
rect 2085 1301 2094 1313
rect 1823 1264 1827 1284
rect 2085 1244 2089 1301
rect 2228 1284 2232 1341
rect 2236 1284 2240 1361
rect 2254 1353 2260 1384
rect 2345 1353 2349 1396
rect 2365 1384 2369 1396
rect 2385 1388 2389 1396
rect 2385 1384 2400 1388
rect 2365 1380 2380 1384
rect 2374 1373 2380 1380
rect 2244 1341 2254 1353
rect 2345 1341 2353 1353
rect 2365 1341 2372 1353
rect 2244 1284 2248 1341
rect 2368 1284 2372 1341
rect 2376 1284 2380 1361
rect 2394 1353 2400 1384
rect 2384 1341 2394 1353
rect 2384 1284 2388 1341
rect 2471 1313 2475 1396
rect 2610 1353 2614 1396
rect 2607 1341 2614 1353
rect 2466 1301 2475 1313
rect 2471 1244 2475 1301
rect 2605 1264 2609 1341
rect 2632 1299 2636 1356
rect 2640 1352 2644 1356
rect 2640 1344 2658 1352
rect 2654 1333 2658 1344
rect 2731 1342 2735 1356
rect 2751 1342 2755 1356
rect 2719 1336 2735 1342
rect 2740 1336 2755 1342
rect 2625 1287 2634 1299
rect 2625 1264 2629 1287
rect 2654 1276 2658 1321
rect 2719 1299 2726 1336
rect 2740 1313 2746 1336
rect 2645 1269 2658 1276
rect 2719 1274 2726 1287
rect 2645 1264 2649 1269
rect 2719 1268 2738 1274
rect 2734 1264 2738 1268
rect 2742 1264 2746 1301
rect 2771 1299 2775 1356
rect 2890 1353 2894 1396
rect 2887 1341 2894 1353
rect 2766 1287 2775 1299
rect 2764 1244 2768 1287
rect 2885 1264 2889 1341
rect 2912 1299 2916 1356
rect 2920 1352 2924 1356
rect 3030 1353 3034 1396
rect 2920 1344 2938 1352
rect 2934 1333 2938 1344
rect 3027 1341 3034 1353
rect 2905 1287 2914 1299
rect 2905 1264 2909 1287
rect 2934 1276 2938 1321
rect 2925 1269 2938 1276
rect 2925 1264 2929 1269
rect 3025 1264 3029 1341
rect 3052 1299 3056 1356
rect 3060 1352 3064 1356
rect 3170 1353 3174 1396
rect 3060 1344 3078 1352
rect 3074 1333 3078 1344
rect 3167 1341 3174 1353
rect 3045 1287 3054 1299
rect 3045 1264 3049 1287
rect 3074 1276 3078 1321
rect 3065 1269 3078 1276
rect 3065 1264 3069 1269
rect 3165 1264 3169 1341
rect 3192 1299 3196 1356
rect 3200 1352 3204 1356
rect 3200 1344 3218 1352
rect 3214 1333 3218 1344
rect 3185 1287 3194 1299
rect 3185 1264 3189 1287
rect 3214 1276 3218 1321
rect 3205 1269 3218 1276
rect 3305 1313 3309 1396
rect 3391 1313 3395 1396
rect 3503 1350 3507 1356
rect 3503 1338 3505 1350
rect 3305 1301 3314 1313
rect 3386 1301 3395 1313
rect 3205 1264 3209 1269
rect 3305 1244 3309 1301
rect 3391 1244 3395 1301
rect 3525 1333 3529 1396
rect 3525 1321 3534 1333
rect 3503 1270 3505 1282
rect 3503 1264 3507 1270
rect 3525 1244 3529 1321
rect 3645 1299 3649 1356
rect 3665 1342 3669 1356
rect 3685 1342 3689 1356
rect 3776 1352 3780 1356
rect 3762 1344 3780 1352
rect 3665 1336 3680 1342
rect 3685 1336 3701 1342
rect 3674 1313 3680 1336
rect 3645 1287 3654 1299
rect 3652 1244 3656 1287
rect 3674 1264 3678 1301
rect 3694 1299 3701 1336
rect 3762 1333 3766 1344
rect 3694 1274 3701 1287
rect 3682 1268 3701 1274
rect 3762 1276 3766 1321
rect 3784 1299 3788 1356
rect 3806 1353 3810 1396
rect 3806 1341 3813 1353
rect 3786 1287 3795 1299
rect 3762 1269 3775 1276
rect 3682 1264 3686 1268
rect 3771 1264 3775 1269
rect 3791 1264 3795 1287
rect 3811 1264 3815 1341
rect 3925 1313 3929 1396
rect 4030 1353 4034 1396
rect 4027 1341 4034 1353
rect 3925 1301 3934 1313
rect 3925 1244 3929 1301
rect 4025 1264 4029 1341
rect 4052 1299 4056 1356
rect 4060 1352 4064 1356
rect 4170 1353 4174 1396
rect 4060 1344 4078 1352
rect 4074 1333 4078 1344
rect 4167 1341 4174 1353
rect 4045 1287 4054 1299
rect 4045 1264 4049 1287
rect 4074 1276 4078 1321
rect 4065 1269 4078 1276
rect 4065 1264 4069 1269
rect 4165 1264 4169 1341
rect 4192 1299 4196 1356
rect 4200 1352 4204 1356
rect 4200 1344 4218 1352
rect 4214 1333 4218 1344
rect 4185 1287 4194 1299
rect 4185 1264 4189 1287
rect 4214 1276 4218 1321
rect 4305 1299 4309 1356
rect 4325 1342 4329 1356
rect 4345 1342 4349 1356
rect 4450 1353 4454 1396
rect 4325 1336 4340 1342
rect 4345 1336 4361 1342
rect 4447 1341 4454 1353
rect 4334 1313 4340 1336
rect 4305 1287 4314 1299
rect 4205 1269 4218 1276
rect 4205 1264 4209 1269
rect 4312 1244 4316 1287
rect 4334 1264 4338 1301
rect 4354 1299 4361 1336
rect 4354 1274 4361 1287
rect 4342 1268 4361 1274
rect 4342 1264 4346 1268
rect 4445 1264 4449 1341
rect 4472 1299 4476 1356
rect 4480 1352 4484 1356
rect 4596 1352 4600 1356
rect 4480 1344 4498 1352
rect 4494 1333 4498 1344
rect 4582 1344 4600 1352
rect 4582 1333 4586 1344
rect 4465 1287 4474 1299
rect 4465 1264 4469 1287
rect 4494 1276 4498 1321
rect 4485 1269 4498 1276
rect 4582 1276 4586 1321
rect 4604 1299 4608 1356
rect 4626 1353 4630 1396
rect 4626 1341 4633 1353
rect 4606 1287 4615 1299
rect 4582 1269 4595 1276
rect 4485 1264 4489 1269
rect 4591 1264 4595 1269
rect 4611 1264 4615 1287
rect 4631 1264 4635 1341
rect 4731 1319 4735 1396
rect 4726 1307 4735 1319
rect 4729 1291 4735 1307
rect 4751 1319 4755 1396
rect 4856 1352 4860 1356
rect 4842 1344 4860 1352
rect 4842 1333 4846 1344
rect 4751 1307 4754 1319
rect 4751 1291 4757 1307
rect 4729 1284 4737 1291
rect 4733 1264 4737 1284
rect 4743 1284 4757 1291
rect 4743 1264 4747 1284
rect 4842 1276 4846 1321
rect 4864 1299 4868 1356
rect 4886 1353 4890 1396
rect 4886 1341 4893 1353
rect 4866 1287 4875 1299
rect 4842 1269 4855 1276
rect 4851 1264 4855 1269
rect 4871 1264 4875 1287
rect 4891 1264 4895 1341
rect 4991 1333 4995 1356
rect 4986 1321 4995 1333
rect 4999 1333 5003 1356
rect 4999 1321 5014 1333
rect 4991 1244 4995 1321
rect 5011 1244 5015 1321
rect 5111 1319 5115 1396
rect 5106 1307 5115 1319
rect 5109 1291 5115 1307
rect 5131 1319 5135 1396
rect 5245 1319 5249 1396
rect 5131 1307 5134 1319
rect 5246 1307 5249 1319
rect 5131 1291 5137 1307
rect 5109 1284 5117 1291
rect 5113 1264 5117 1284
rect 5123 1284 5137 1291
rect 5243 1291 5249 1307
rect 5265 1319 5269 1396
rect 5370 1353 5374 1396
rect 5367 1341 5374 1353
rect 5265 1307 5274 1319
rect 5265 1291 5271 1307
rect 5243 1284 5257 1291
rect 5123 1264 5127 1284
rect 5253 1264 5257 1284
rect 5263 1284 5271 1291
rect 5263 1264 5267 1284
rect 5365 1264 5369 1341
rect 5392 1299 5396 1356
rect 5400 1352 5404 1356
rect 5496 1352 5500 1356
rect 5400 1344 5418 1352
rect 5414 1333 5418 1344
rect 5482 1344 5500 1352
rect 5482 1333 5486 1344
rect 5385 1287 5394 1299
rect 5385 1264 5389 1287
rect 5414 1276 5418 1321
rect 5405 1269 5418 1276
rect 5482 1276 5486 1321
rect 5504 1299 5508 1356
rect 5526 1353 5530 1396
rect 5526 1341 5533 1353
rect 5656 1352 5660 1356
rect 5642 1344 5660 1352
rect 5506 1287 5515 1299
rect 5482 1269 5495 1276
rect 5405 1264 5409 1269
rect 5491 1264 5495 1269
rect 5511 1264 5515 1287
rect 5531 1264 5535 1341
rect 5642 1333 5646 1344
rect 5642 1276 5646 1321
rect 5664 1299 5668 1356
rect 5686 1353 5690 1396
rect 5686 1341 5693 1353
rect 5666 1287 5675 1299
rect 5642 1269 5655 1276
rect 5651 1264 5655 1269
rect 5671 1264 5675 1287
rect 5691 1264 5695 1341
rect 108 1220 112 1224
rect 116 1220 120 1224
rect 124 1220 128 1224
rect 214 1220 218 1224
rect 222 1220 226 1224
rect 244 1220 248 1224
rect 388 1220 392 1224
rect 396 1220 400 1224
rect 404 1220 408 1224
rect 505 1220 509 1224
rect 525 1220 529 1224
rect 545 1220 549 1224
rect 645 1220 649 1224
rect 665 1220 669 1224
rect 685 1220 689 1224
rect 815 1220 819 1224
rect 835 1220 839 1224
rect 845 1220 849 1224
rect 933 1220 937 1224
rect 943 1220 947 1224
rect 1065 1220 1069 1224
rect 1152 1220 1156 1224
rect 1160 1220 1164 1224
rect 1168 1220 1172 1224
rect 1293 1220 1297 1224
rect 1303 1220 1307 1224
rect 1433 1220 1437 1224
rect 1443 1220 1447 1224
rect 1553 1220 1557 1224
rect 1563 1220 1567 1224
rect 1708 1220 1712 1224
rect 1716 1220 1720 1224
rect 1724 1220 1728 1224
rect 1813 1220 1817 1224
rect 1823 1220 1827 1224
rect 1968 1220 1972 1224
rect 1976 1220 1980 1224
rect 1984 1220 1988 1224
rect 2085 1220 2089 1224
rect 2228 1220 2232 1224
rect 2236 1220 2240 1224
rect 2244 1220 2248 1224
rect 2368 1220 2372 1224
rect 2376 1220 2380 1224
rect 2384 1220 2388 1224
rect 2471 1220 2475 1224
rect 2605 1220 2609 1224
rect 2625 1220 2629 1224
rect 2645 1220 2649 1224
rect 2734 1220 2738 1224
rect 2742 1220 2746 1224
rect 2764 1220 2768 1224
rect 2885 1220 2889 1224
rect 2905 1220 2909 1224
rect 2925 1220 2929 1224
rect 3025 1220 3029 1224
rect 3045 1220 3049 1224
rect 3065 1220 3069 1224
rect 3165 1220 3169 1224
rect 3185 1220 3189 1224
rect 3205 1220 3209 1224
rect 3305 1220 3309 1224
rect 3391 1220 3395 1224
rect 3503 1220 3507 1224
rect 3525 1220 3529 1224
rect 3652 1220 3656 1224
rect 3674 1220 3678 1224
rect 3682 1220 3686 1224
rect 3771 1220 3775 1224
rect 3791 1220 3795 1224
rect 3811 1220 3815 1224
rect 3925 1220 3929 1224
rect 4025 1220 4029 1224
rect 4045 1220 4049 1224
rect 4065 1220 4069 1224
rect 4165 1220 4169 1224
rect 4185 1220 4189 1224
rect 4205 1220 4209 1224
rect 4312 1220 4316 1224
rect 4334 1220 4338 1224
rect 4342 1220 4346 1224
rect 4445 1220 4449 1224
rect 4465 1220 4469 1224
rect 4485 1220 4489 1224
rect 4591 1220 4595 1224
rect 4611 1220 4615 1224
rect 4631 1220 4635 1224
rect 4733 1220 4737 1224
rect 4743 1220 4747 1224
rect 4851 1220 4855 1224
rect 4871 1220 4875 1224
rect 4891 1220 4895 1224
rect 4991 1220 4995 1224
rect 5011 1220 5015 1224
rect 5113 1220 5117 1224
rect 5123 1220 5127 1224
rect 5253 1220 5257 1224
rect 5263 1220 5267 1224
rect 5365 1220 5369 1224
rect 5385 1220 5389 1224
rect 5405 1220 5409 1224
rect 5491 1220 5495 1224
rect 5511 1220 5515 1224
rect 5531 1220 5535 1224
rect 5651 1220 5655 1224
rect 5671 1220 5675 1224
rect 5691 1220 5695 1224
rect 85 1196 89 1200
rect 174 1196 178 1200
rect 182 1196 186 1200
rect 204 1196 208 1200
rect 311 1196 315 1200
rect 331 1196 335 1200
rect 351 1196 355 1200
rect 451 1196 455 1200
rect 471 1196 475 1200
rect 491 1196 495 1200
rect 628 1196 632 1200
rect 636 1196 640 1200
rect 644 1196 648 1200
rect 731 1196 735 1200
rect 751 1196 755 1200
rect 771 1196 775 1200
rect 894 1196 898 1200
rect 902 1196 906 1200
rect 924 1196 928 1200
rect 1045 1196 1049 1200
rect 1065 1196 1069 1200
rect 1085 1196 1089 1200
rect 1185 1196 1189 1200
rect 1274 1196 1278 1200
rect 1282 1196 1286 1200
rect 1304 1196 1308 1200
rect 1425 1196 1429 1200
rect 1525 1196 1529 1200
rect 1545 1196 1549 1200
rect 1651 1196 1655 1200
rect 1788 1196 1792 1200
rect 1796 1196 1800 1200
rect 1804 1196 1808 1200
rect 1913 1196 1917 1200
rect 1923 1196 1927 1200
rect 2025 1196 2029 1200
rect 2045 1196 2049 1200
rect 2065 1196 2069 1200
rect 2188 1196 2192 1200
rect 2196 1196 2200 1200
rect 2204 1196 2208 1200
rect 2328 1196 2332 1200
rect 2336 1196 2340 1200
rect 2344 1196 2348 1200
rect 2445 1196 2449 1200
rect 2465 1196 2469 1200
rect 2485 1196 2489 1200
rect 2608 1196 2612 1200
rect 2616 1196 2620 1200
rect 2624 1196 2628 1200
rect 2731 1196 2735 1200
rect 2831 1196 2835 1200
rect 2851 1196 2855 1200
rect 2951 1196 2955 1200
rect 2971 1196 2975 1200
rect 3071 1196 3075 1200
rect 3081 1196 3085 1200
rect 3101 1196 3105 1200
rect 3225 1196 3229 1200
rect 3245 1196 3249 1200
rect 3365 1196 3369 1200
rect 3385 1196 3389 1200
rect 3485 1196 3489 1200
rect 3585 1196 3589 1200
rect 3605 1196 3609 1200
rect 3625 1196 3629 1200
rect 3725 1196 3729 1200
rect 3745 1196 3749 1200
rect 3765 1196 3769 1200
rect 3853 1196 3857 1200
rect 3863 1196 3867 1200
rect 3973 1196 3977 1200
rect 3983 1196 3987 1200
rect 4091 1196 4095 1200
rect 4111 1196 4115 1200
rect 4211 1196 4215 1200
rect 4332 1196 4336 1200
rect 4354 1196 4358 1200
rect 4362 1196 4366 1200
rect 4485 1196 4489 1200
rect 4505 1196 4509 1200
rect 4525 1196 4529 1200
rect 4632 1196 4636 1200
rect 4654 1196 4658 1200
rect 4662 1196 4666 1200
rect 4751 1196 4755 1200
rect 4771 1196 4775 1200
rect 4791 1196 4795 1200
rect 4891 1196 4895 1200
rect 4913 1196 4917 1200
rect 5011 1196 5015 1200
rect 5111 1196 5115 1200
rect 5233 1196 5237 1200
rect 5243 1196 5247 1200
rect 5365 1196 5369 1200
rect 5385 1196 5389 1200
rect 5405 1196 5409 1200
rect 5491 1196 5495 1200
rect 5511 1196 5515 1200
rect 5648 1196 5652 1200
rect 5656 1196 5660 1200
rect 5664 1196 5668 1200
rect 5765 1196 5769 1200
rect 85 1119 89 1176
rect 174 1152 178 1156
rect 159 1146 178 1152
rect 159 1133 166 1146
rect 85 1107 94 1119
rect 85 1024 89 1107
rect 159 1084 166 1121
rect 182 1119 186 1156
rect 204 1133 208 1176
rect 311 1151 315 1156
rect 302 1144 315 1151
rect 206 1121 215 1133
rect 180 1084 186 1107
rect 159 1078 175 1084
rect 180 1078 195 1084
rect 171 1064 175 1078
rect 191 1064 195 1078
rect 211 1064 215 1121
rect 302 1099 306 1144
rect 331 1133 335 1156
rect 326 1121 335 1133
rect 302 1076 306 1087
rect 302 1068 320 1076
rect 316 1064 320 1068
rect 324 1064 328 1121
rect 351 1079 355 1156
rect 451 1151 455 1156
rect 442 1144 455 1151
rect 442 1099 446 1144
rect 471 1133 475 1156
rect 466 1121 475 1133
rect 346 1067 353 1079
rect 442 1076 446 1087
rect 442 1068 460 1076
rect 346 1024 350 1067
rect 456 1064 460 1068
rect 464 1064 468 1121
rect 491 1079 495 1156
rect 731 1151 735 1156
rect 722 1144 735 1151
rect 628 1079 632 1136
rect 486 1067 493 1079
rect 605 1067 613 1079
rect 625 1067 632 1079
rect 486 1024 490 1067
rect 605 1024 609 1067
rect 636 1059 640 1136
rect 644 1079 648 1136
rect 722 1099 726 1144
rect 751 1133 755 1156
rect 746 1121 755 1133
rect 644 1067 654 1079
rect 722 1076 726 1087
rect 722 1068 740 1076
rect 634 1040 640 1047
rect 625 1036 640 1040
rect 654 1036 660 1067
rect 736 1064 740 1068
rect 744 1064 748 1121
rect 771 1079 775 1156
rect 894 1152 898 1156
rect 879 1146 898 1152
rect 879 1133 886 1146
rect 879 1084 886 1121
rect 902 1119 906 1156
rect 924 1133 928 1176
rect 926 1121 935 1133
rect 900 1084 906 1107
rect 766 1067 773 1079
rect 879 1078 895 1084
rect 900 1078 915 1084
rect 625 1024 629 1036
rect 645 1032 660 1036
rect 645 1024 649 1032
rect 766 1024 770 1067
rect 891 1064 895 1078
rect 911 1064 915 1078
rect 931 1064 935 1121
rect 1045 1079 1049 1156
rect 1065 1133 1069 1156
rect 1085 1151 1089 1156
rect 1085 1144 1098 1151
rect 1065 1121 1074 1133
rect 1047 1067 1054 1079
rect 1050 1024 1054 1067
rect 1072 1064 1076 1121
rect 1094 1099 1098 1144
rect 1185 1119 1189 1176
rect 1274 1152 1278 1156
rect 1259 1146 1278 1152
rect 1259 1133 1266 1146
rect 1185 1107 1194 1119
rect 1094 1076 1098 1087
rect 1080 1068 1098 1076
rect 1080 1064 1084 1068
rect 1185 1024 1189 1107
rect 1259 1084 1266 1121
rect 1282 1119 1286 1156
rect 1304 1133 1308 1176
rect 1306 1121 1315 1133
rect 1280 1084 1286 1107
rect 1259 1078 1275 1084
rect 1280 1078 1295 1084
rect 1271 1064 1275 1078
rect 1291 1064 1295 1078
rect 1311 1064 1315 1121
rect 1425 1119 1429 1176
rect 1425 1107 1434 1119
rect 1425 1024 1429 1107
rect 1525 1099 1529 1176
rect 1545 1099 1549 1176
rect 1651 1119 1655 1176
rect 1913 1136 1917 1156
rect 1646 1107 1655 1119
rect 1526 1087 1541 1099
rect 1537 1064 1541 1087
rect 1545 1087 1554 1099
rect 1545 1064 1549 1087
rect 1651 1024 1655 1107
rect 1788 1079 1792 1136
rect 1765 1067 1773 1079
rect 1785 1067 1792 1079
rect 1765 1024 1769 1067
rect 1796 1059 1800 1136
rect 1804 1079 1808 1136
rect 1903 1129 1917 1136
rect 1923 1136 1927 1156
rect 1923 1129 1931 1136
rect 1903 1113 1909 1129
rect 1906 1101 1909 1113
rect 1804 1067 1814 1079
rect 1794 1040 1800 1047
rect 1785 1036 1800 1040
rect 1814 1036 1820 1067
rect 1785 1024 1789 1036
rect 1805 1032 1820 1036
rect 1805 1024 1809 1032
rect 1905 1024 1909 1101
rect 1925 1113 1931 1129
rect 1925 1101 1934 1113
rect 1925 1024 1929 1101
rect 2025 1079 2029 1156
rect 2045 1133 2049 1156
rect 2065 1151 2069 1156
rect 2065 1144 2078 1151
rect 2045 1121 2054 1133
rect 2027 1067 2034 1079
rect 2030 1024 2034 1067
rect 2052 1064 2056 1121
rect 2074 1099 2078 1144
rect 2074 1076 2078 1087
rect 2188 1079 2192 1136
rect 2060 1068 2078 1076
rect 2060 1064 2064 1068
rect 2165 1067 2173 1079
rect 2185 1067 2192 1079
rect 2165 1024 2169 1067
rect 2196 1059 2200 1136
rect 2204 1079 2208 1136
rect 2328 1079 2332 1136
rect 2204 1067 2214 1079
rect 2305 1067 2313 1079
rect 2325 1067 2332 1079
rect 2194 1040 2200 1047
rect 2185 1036 2200 1040
rect 2214 1036 2220 1067
rect 2185 1024 2189 1036
rect 2205 1032 2220 1036
rect 2205 1024 2209 1032
rect 2305 1024 2309 1067
rect 2336 1059 2340 1136
rect 2344 1079 2348 1136
rect 2445 1079 2449 1156
rect 2465 1133 2469 1156
rect 2485 1151 2489 1156
rect 2485 1144 2498 1151
rect 2465 1121 2474 1133
rect 2344 1067 2354 1079
rect 2447 1067 2454 1079
rect 2334 1040 2340 1047
rect 2325 1036 2340 1040
rect 2354 1036 2360 1067
rect 2325 1024 2329 1036
rect 2345 1032 2360 1036
rect 2345 1024 2349 1032
rect 2450 1024 2454 1067
rect 2472 1064 2476 1121
rect 2494 1099 2498 1144
rect 2494 1076 2498 1087
rect 2608 1079 2612 1136
rect 2480 1068 2498 1076
rect 2480 1064 2484 1068
rect 2585 1067 2593 1079
rect 2605 1067 2612 1079
rect 2585 1024 2589 1067
rect 2616 1059 2620 1136
rect 2624 1079 2628 1136
rect 2731 1119 2735 1176
rect 2726 1107 2735 1119
rect 2624 1067 2634 1079
rect 2614 1040 2620 1047
rect 2605 1036 2620 1040
rect 2634 1036 2640 1067
rect 2605 1024 2609 1036
rect 2625 1032 2640 1036
rect 2625 1024 2629 1032
rect 2731 1024 2735 1107
rect 2831 1099 2835 1176
rect 2851 1099 2855 1176
rect 2951 1099 2955 1176
rect 2971 1099 2975 1176
rect 3071 1099 3075 1156
rect 3081 1113 3085 1156
rect 3101 1150 3105 1156
rect 3107 1138 3119 1150
rect 3081 1101 3094 1113
rect 2826 1087 2835 1099
rect 2831 1064 2835 1087
rect 2839 1087 2854 1099
rect 2946 1087 2955 1099
rect 2839 1064 2843 1087
rect 2951 1064 2955 1087
rect 2959 1087 2974 1099
rect 3066 1087 3075 1099
rect 2959 1064 2963 1087
rect 3071 1024 3075 1087
rect 3093 1024 3097 1101
rect 3115 1064 3119 1138
rect 3225 1099 3229 1176
rect 3245 1099 3249 1176
rect 3365 1099 3369 1176
rect 3385 1099 3389 1176
rect 3485 1119 3489 1176
rect 3485 1107 3494 1119
rect 3226 1087 3241 1099
rect 3237 1064 3241 1087
rect 3245 1087 3254 1099
rect 3366 1087 3381 1099
rect 3245 1064 3249 1087
rect 3377 1064 3381 1087
rect 3385 1087 3394 1099
rect 3385 1064 3389 1087
rect 3485 1024 3489 1107
rect 3585 1079 3589 1156
rect 3605 1133 3609 1156
rect 3625 1151 3629 1156
rect 3625 1144 3638 1151
rect 3605 1121 3614 1133
rect 3587 1067 3594 1079
rect 3590 1024 3594 1067
rect 3612 1064 3616 1121
rect 3634 1099 3638 1144
rect 3634 1076 3638 1087
rect 3725 1079 3729 1156
rect 3745 1133 3749 1156
rect 3765 1151 3769 1156
rect 3765 1144 3778 1151
rect 3745 1121 3754 1133
rect 3620 1068 3638 1076
rect 3620 1064 3624 1068
rect 3727 1067 3734 1079
rect 3730 1024 3734 1067
rect 3752 1064 3756 1121
rect 3774 1099 3778 1144
rect 3853 1136 3857 1156
rect 3849 1129 3857 1136
rect 3863 1136 3867 1156
rect 3973 1136 3977 1156
rect 3863 1129 3877 1136
rect 3849 1113 3855 1129
rect 3846 1101 3855 1113
rect 3774 1076 3778 1087
rect 3760 1068 3778 1076
rect 3760 1064 3764 1068
rect 3851 1024 3855 1101
rect 3871 1113 3877 1129
rect 3969 1129 3977 1136
rect 3983 1136 3987 1156
rect 3983 1129 3997 1136
rect 3969 1113 3975 1129
rect 3871 1101 3874 1113
rect 3966 1101 3975 1113
rect 3871 1024 3875 1101
rect 3971 1024 3975 1101
rect 3991 1113 3997 1129
rect 3991 1101 3994 1113
rect 3991 1024 3995 1101
rect 4091 1099 4095 1176
rect 4111 1099 4115 1176
rect 4211 1119 4215 1176
rect 4332 1133 4336 1176
rect 4206 1107 4215 1119
rect 4086 1087 4095 1099
rect 4091 1064 4095 1087
rect 4099 1087 4114 1099
rect 4099 1064 4103 1087
rect 4211 1024 4215 1107
rect 4325 1121 4334 1133
rect 4325 1064 4329 1121
rect 4354 1119 4358 1156
rect 4362 1152 4366 1156
rect 4362 1146 4381 1152
rect 4374 1133 4381 1146
rect 4354 1084 4360 1107
rect 4374 1084 4381 1121
rect 4345 1078 4360 1084
rect 4365 1078 4381 1084
rect 4485 1079 4489 1156
rect 4505 1133 4509 1156
rect 4525 1151 4529 1156
rect 4525 1144 4538 1151
rect 4505 1121 4514 1133
rect 4345 1064 4349 1078
rect 4365 1064 4369 1078
rect 4487 1067 4494 1079
rect 4490 1024 4494 1067
rect 4512 1064 4516 1121
rect 4534 1099 4538 1144
rect 4632 1133 4636 1176
rect 4625 1121 4634 1133
rect 4534 1076 4538 1087
rect 4520 1068 4538 1076
rect 4520 1064 4524 1068
rect 4625 1064 4629 1121
rect 4654 1119 4658 1156
rect 4662 1152 4666 1156
rect 4662 1146 4681 1152
rect 4751 1151 4755 1156
rect 4674 1133 4681 1146
rect 4742 1144 4755 1151
rect 4654 1084 4660 1107
rect 4674 1084 4681 1121
rect 4742 1099 4746 1144
rect 4771 1133 4775 1156
rect 4766 1121 4775 1133
rect 4645 1078 4660 1084
rect 4665 1078 4681 1084
rect 4645 1064 4649 1078
rect 4665 1064 4669 1078
rect 4742 1076 4746 1087
rect 4742 1068 4760 1076
rect 4756 1064 4760 1068
rect 4764 1064 4768 1121
rect 4791 1079 4795 1156
rect 4891 1099 4895 1176
rect 4913 1150 4917 1156
rect 4915 1138 4917 1150
rect 5011 1119 5015 1176
rect 5111 1119 5115 1176
rect 5233 1136 5237 1156
rect 5006 1107 5015 1119
rect 5106 1107 5115 1119
rect 5223 1129 5237 1136
rect 5243 1136 5247 1156
rect 5243 1129 5251 1136
rect 5223 1113 5229 1129
rect 4886 1087 4895 1099
rect 4786 1067 4793 1079
rect 4786 1024 4790 1067
rect 4891 1024 4895 1087
rect 4915 1070 4917 1082
rect 4913 1064 4917 1070
rect 5011 1024 5015 1107
rect 5111 1024 5115 1107
rect 5226 1101 5229 1113
rect 5225 1024 5229 1101
rect 5245 1113 5251 1129
rect 5245 1101 5254 1113
rect 5245 1024 5249 1101
rect 5365 1079 5369 1156
rect 5385 1133 5389 1156
rect 5405 1151 5409 1156
rect 5405 1144 5418 1151
rect 5385 1121 5394 1133
rect 5367 1067 5374 1079
rect 5370 1024 5374 1067
rect 5392 1064 5396 1121
rect 5414 1099 5418 1144
rect 5491 1099 5495 1176
rect 5511 1099 5515 1176
rect 5486 1087 5495 1099
rect 5414 1076 5418 1087
rect 5400 1068 5418 1076
rect 5400 1064 5404 1068
rect 5491 1064 5495 1087
rect 5499 1087 5514 1099
rect 5499 1064 5503 1087
rect 5648 1079 5652 1136
rect 5625 1067 5633 1079
rect 5645 1067 5652 1079
rect 5625 1024 5629 1067
rect 5656 1059 5660 1136
rect 5664 1079 5668 1136
rect 5765 1119 5769 1176
rect 5765 1107 5774 1119
rect 5664 1067 5674 1079
rect 5654 1040 5660 1047
rect 5645 1036 5660 1040
rect 5674 1036 5680 1067
rect 5645 1024 5649 1036
rect 5665 1032 5680 1036
rect 5665 1024 5669 1032
rect 5765 1024 5769 1107
rect 85 980 89 984
rect 171 980 175 984
rect 191 980 195 984
rect 211 980 215 984
rect 316 980 320 984
rect 324 980 328 984
rect 346 980 350 984
rect 456 980 460 984
rect 464 980 468 984
rect 486 980 490 984
rect 605 980 609 984
rect 625 980 629 984
rect 645 980 649 984
rect 736 980 740 984
rect 744 980 748 984
rect 766 980 770 984
rect 891 980 895 984
rect 911 980 915 984
rect 931 980 935 984
rect 1050 980 1054 984
rect 1072 980 1076 984
rect 1080 980 1084 984
rect 1185 980 1189 984
rect 1271 980 1275 984
rect 1291 980 1295 984
rect 1311 980 1315 984
rect 1425 980 1429 984
rect 1537 980 1541 984
rect 1545 980 1549 984
rect 1651 980 1655 984
rect 1765 980 1769 984
rect 1785 980 1789 984
rect 1805 980 1809 984
rect 1905 980 1909 984
rect 1925 980 1929 984
rect 2030 980 2034 984
rect 2052 980 2056 984
rect 2060 980 2064 984
rect 2165 980 2169 984
rect 2185 980 2189 984
rect 2205 980 2209 984
rect 2305 980 2309 984
rect 2325 980 2329 984
rect 2345 980 2349 984
rect 2450 980 2454 984
rect 2472 980 2476 984
rect 2480 980 2484 984
rect 2585 980 2589 984
rect 2605 980 2609 984
rect 2625 980 2629 984
rect 2731 980 2735 984
rect 2831 980 2835 984
rect 2839 980 2843 984
rect 2951 980 2955 984
rect 2959 980 2963 984
rect 3071 980 3075 984
rect 3093 980 3097 984
rect 3115 980 3119 984
rect 3237 980 3241 984
rect 3245 980 3249 984
rect 3377 980 3381 984
rect 3385 980 3389 984
rect 3485 980 3489 984
rect 3590 980 3594 984
rect 3612 980 3616 984
rect 3620 980 3624 984
rect 3730 980 3734 984
rect 3752 980 3756 984
rect 3760 980 3764 984
rect 3851 980 3855 984
rect 3871 980 3875 984
rect 3971 980 3975 984
rect 3991 980 3995 984
rect 4091 980 4095 984
rect 4099 980 4103 984
rect 4211 980 4215 984
rect 4325 980 4329 984
rect 4345 980 4349 984
rect 4365 980 4369 984
rect 4490 980 4494 984
rect 4512 980 4516 984
rect 4520 980 4524 984
rect 4625 980 4629 984
rect 4645 980 4649 984
rect 4665 980 4669 984
rect 4756 980 4760 984
rect 4764 980 4768 984
rect 4786 980 4790 984
rect 4891 980 4895 984
rect 4913 980 4917 984
rect 5011 980 5015 984
rect 5111 980 5115 984
rect 5225 980 5229 984
rect 5245 980 5249 984
rect 5370 980 5374 984
rect 5392 980 5396 984
rect 5400 980 5404 984
rect 5491 980 5495 984
rect 5499 980 5503 984
rect 5625 980 5629 984
rect 5645 980 5649 984
rect 5665 980 5669 984
rect 5765 980 5769 984
rect 85 956 89 960
rect 105 956 109 960
rect 125 956 129 960
rect 211 956 215 960
rect 231 956 235 960
rect 251 956 255 960
rect 365 956 369 960
rect 385 956 389 960
rect 405 956 409 960
rect 505 956 509 960
rect 525 956 529 960
rect 545 956 549 960
rect 645 956 649 960
rect 665 956 669 960
rect 685 956 689 960
rect 771 956 775 960
rect 791 956 795 960
rect 811 956 815 960
rect 930 956 934 960
rect 952 956 956 960
rect 960 956 964 960
rect 1065 956 1069 960
rect 1085 956 1089 960
rect 1105 956 1109 960
rect 1196 956 1200 960
rect 1204 956 1208 960
rect 1226 956 1230 960
rect 1345 956 1349 960
rect 1365 956 1369 960
rect 1385 956 1389 960
rect 1471 956 1475 960
rect 1571 956 1575 960
rect 1591 956 1595 960
rect 1725 956 1729 960
rect 1745 956 1749 960
rect 1765 956 1769 960
rect 1865 956 1869 960
rect 1885 956 1889 960
rect 1905 956 1909 960
rect 1991 956 1995 960
rect 2011 956 2015 960
rect 2031 956 2035 960
rect 2136 956 2140 960
rect 2144 956 2148 960
rect 2166 956 2170 960
rect 2271 956 2275 960
rect 2293 956 2297 960
rect 2315 956 2319 960
rect 2411 956 2415 960
rect 2525 956 2529 960
rect 2545 956 2549 960
rect 2655 956 2659 960
rect 2675 956 2679 960
rect 2685 956 2689 960
rect 2771 956 2775 960
rect 2791 956 2795 960
rect 2905 956 2909 960
rect 2925 956 2929 960
rect 3031 956 3035 960
rect 3145 956 3149 960
rect 3265 956 3269 960
rect 3285 956 3289 960
rect 3417 956 3421 960
rect 3425 956 3429 960
rect 3537 956 3541 960
rect 3545 956 3549 960
rect 3645 956 3649 960
rect 3665 956 3669 960
rect 3685 956 3689 960
rect 3785 956 3789 960
rect 3890 956 3894 960
rect 3912 956 3916 960
rect 3920 956 3924 960
rect 4011 956 4015 960
rect 4031 956 4035 960
rect 4150 956 4154 960
rect 4172 956 4176 960
rect 4180 956 4184 960
rect 4290 956 4294 960
rect 4312 956 4316 960
rect 4320 956 4324 960
rect 4431 956 4435 960
rect 4550 956 4554 960
rect 4572 956 4576 960
rect 4580 956 4584 960
rect 4671 956 4675 960
rect 4691 956 4695 960
rect 4711 956 4715 960
rect 4823 956 4827 960
rect 4845 956 4849 960
rect 4950 956 4954 960
rect 4972 956 4976 960
rect 4980 956 4984 960
rect 5071 956 5075 960
rect 5091 956 5095 960
rect 5111 956 5115 960
rect 5235 956 5239 960
rect 5255 956 5259 960
rect 5265 956 5269 960
rect 5385 956 5389 960
rect 5485 956 5489 960
rect 5505 956 5509 960
rect 5525 956 5529 960
rect 5545 956 5549 960
rect 5656 956 5660 960
rect 5664 956 5668 960
rect 5686 956 5690 960
rect 85 873 89 916
rect 105 904 109 916
rect 125 908 129 916
rect 125 904 140 908
rect 105 900 120 904
rect 114 893 120 900
rect 85 861 93 873
rect 105 861 112 873
rect 108 804 112 861
rect 116 804 120 881
rect 134 873 140 904
rect 124 861 134 873
rect 211 862 215 876
rect 231 862 235 876
rect 124 804 128 861
rect 199 856 215 862
rect 220 856 235 862
rect 199 819 206 856
rect 220 833 226 856
rect 199 794 206 807
rect 199 788 218 794
rect 214 784 218 788
rect 222 784 226 821
rect 251 819 255 876
rect 365 873 369 916
rect 385 904 389 916
rect 405 908 409 916
rect 405 904 420 908
rect 385 900 400 904
rect 394 893 400 900
rect 365 861 373 873
rect 385 861 392 873
rect 246 807 255 819
rect 244 764 248 807
rect 388 804 392 861
rect 396 804 400 881
rect 414 873 420 904
rect 404 861 414 873
rect 404 804 408 861
rect 505 819 509 876
rect 525 862 529 876
rect 545 862 549 876
rect 645 873 649 916
rect 665 904 669 916
rect 685 908 689 916
rect 685 904 700 908
rect 665 900 680 904
rect 674 893 680 900
rect 525 856 540 862
rect 545 856 561 862
rect 645 861 653 873
rect 665 861 672 873
rect 534 833 540 856
rect 505 807 514 819
rect 512 764 516 807
rect 534 784 538 821
rect 554 819 561 856
rect 554 794 561 807
rect 668 804 672 861
rect 676 804 680 881
rect 694 873 700 904
rect 684 861 694 873
rect 771 862 775 876
rect 791 862 795 876
rect 684 804 688 861
rect 759 856 775 862
rect 780 856 795 862
rect 759 819 766 856
rect 780 833 786 856
rect 542 788 561 794
rect 542 784 546 788
rect 759 794 766 807
rect 759 788 778 794
rect 774 784 778 788
rect 782 784 786 821
rect 811 819 815 876
rect 930 873 934 916
rect 927 861 934 873
rect 806 807 815 819
rect 804 764 808 807
rect 925 784 929 861
rect 952 819 956 876
rect 960 872 964 876
rect 1065 873 1069 916
rect 1085 904 1089 916
rect 1105 908 1109 916
rect 1105 904 1120 908
rect 1085 900 1100 904
rect 1094 893 1100 900
rect 960 864 978 872
rect 974 853 978 864
rect 1065 861 1073 873
rect 1085 861 1092 873
rect 945 807 954 819
rect 945 784 949 807
rect 974 796 978 841
rect 1088 804 1092 861
rect 1096 804 1100 881
rect 1114 873 1120 904
rect 1104 861 1114 873
rect 1196 872 1200 876
rect 1182 864 1200 872
rect 1104 804 1108 861
rect 1182 853 1186 864
rect 965 789 978 796
rect 965 784 969 789
rect 1182 796 1186 841
rect 1204 819 1208 876
rect 1226 873 1230 916
rect 1345 873 1349 916
rect 1365 904 1369 916
rect 1385 908 1389 916
rect 1385 904 1400 908
rect 1365 900 1380 904
rect 1374 893 1380 900
rect 1226 861 1233 873
rect 1345 861 1353 873
rect 1365 861 1372 873
rect 1206 807 1215 819
rect 1182 789 1195 796
rect 1191 784 1195 789
rect 1211 784 1215 807
rect 1231 784 1235 861
rect 1368 804 1372 861
rect 1376 804 1380 881
rect 1394 873 1400 904
rect 1384 861 1394 873
rect 1384 804 1388 861
rect 1471 833 1475 916
rect 1571 839 1575 916
rect 1466 821 1475 833
rect 1566 827 1575 839
rect 1471 764 1475 821
rect 1569 811 1575 827
rect 1591 839 1595 916
rect 1725 873 1729 916
rect 1745 904 1749 916
rect 1765 908 1769 916
rect 1765 904 1780 908
rect 1745 900 1760 904
rect 1754 893 1760 900
rect 1725 861 1733 873
rect 1745 861 1752 873
rect 1591 827 1594 839
rect 1591 811 1597 827
rect 1569 804 1577 811
rect 1573 784 1577 804
rect 1583 804 1597 811
rect 1748 804 1752 861
rect 1756 804 1760 881
rect 1774 873 1780 904
rect 1865 873 1869 916
rect 1885 904 1889 916
rect 1905 908 1909 916
rect 1991 908 1995 916
rect 1905 904 1920 908
rect 1885 900 1900 904
rect 1894 893 1900 900
rect 1764 861 1774 873
rect 1865 861 1873 873
rect 1885 861 1892 873
rect 1764 804 1768 861
rect 1888 804 1892 861
rect 1896 804 1900 881
rect 1914 873 1920 904
rect 1980 904 1995 908
rect 2011 904 2015 916
rect 1980 873 1986 904
rect 2000 900 2015 904
rect 2000 893 2006 900
rect 1904 861 1914 873
rect 1986 861 1996 873
rect 1904 804 1908 861
rect 1992 804 1996 861
rect 2000 804 2004 881
rect 2031 873 2035 916
rect 2008 861 2015 873
rect 2027 861 2035 873
rect 2136 872 2140 876
rect 2122 864 2140 872
rect 2008 804 2012 861
rect 2122 853 2126 864
rect 1583 784 1587 804
rect 2122 796 2126 841
rect 2144 819 2148 876
rect 2166 873 2170 916
rect 2166 861 2173 873
rect 2146 807 2155 819
rect 2122 789 2135 796
rect 2131 784 2135 789
rect 2151 784 2155 807
rect 2171 784 2175 861
rect 2271 853 2275 916
rect 2266 841 2275 853
rect 2271 784 2275 841
rect 2293 839 2297 916
rect 2281 827 2294 839
rect 2281 784 2285 827
rect 2315 802 2319 876
rect 2411 833 2415 916
rect 2525 839 2529 916
rect 2406 821 2415 833
rect 2526 827 2529 839
rect 2307 790 2319 802
rect 2301 784 2305 790
rect 2411 764 2415 821
rect 2523 811 2529 827
rect 2545 839 2549 916
rect 2655 871 2659 876
rect 2675 853 2679 876
rect 2685 872 2689 876
rect 2685 867 2698 872
rect 2545 827 2554 839
rect 2545 811 2551 827
rect 2523 804 2537 811
rect 2533 784 2537 804
rect 2543 804 2551 811
rect 2543 784 2547 804
rect 2645 792 2655 804
rect 2645 784 2649 792
rect 2675 777 2679 841
rect 2665 771 2679 777
rect 2694 833 2698 867
rect 2771 839 2775 916
rect 2766 827 2775 839
rect 2694 776 2698 821
rect 2769 811 2775 827
rect 2791 839 2795 916
rect 2905 839 2909 916
rect 2791 827 2794 839
rect 2906 827 2909 839
rect 2791 811 2797 827
rect 2769 804 2777 811
rect 2773 784 2777 804
rect 2783 804 2797 811
rect 2903 811 2909 827
rect 2925 839 2929 916
rect 2925 827 2934 839
rect 3031 833 3035 916
rect 2925 811 2931 827
rect 3026 821 3035 833
rect 2903 804 2917 811
rect 2783 784 2787 804
rect 2913 784 2917 804
rect 2923 804 2931 811
rect 2923 784 2927 804
rect 2685 771 2698 776
rect 2665 764 2669 771
rect 2685 764 2689 771
rect 3031 764 3035 821
rect 3145 833 3149 916
rect 3265 839 3269 916
rect 3145 821 3154 833
rect 3266 827 3269 839
rect 3145 764 3149 821
rect 3263 811 3269 827
rect 3285 839 3289 916
rect 3417 853 3421 876
rect 3406 841 3421 853
rect 3425 853 3429 876
rect 3537 853 3541 876
rect 3425 841 3434 853
rect 3526 841 3541 853
rect 3545 853 3549 876
rect 3545 841 3554 853
rect 3285 827 3294 839
rect 3285 811 3291 827
rect 3263 804 3277 811
rect 3273 784 3277 804
rect 3283 804 3291 811
rect 3283 784 3287 804
rect 3405 764 3409 841
rect 3425 764 3429 841
rect 3525 764 3529 841
rect 3545 764 3549 841
rect 3645 819 3649 876
rect 3665 862 3669 876
rect 3685 862 3689 876
rect 3665 856 3680 862
rect 3685 856 3701 862
rect 3674 833 3680 856
rect 3645 807 3654 819
rect 3652 764 3656 807
rect 3674 784 3678 821
rect 3694 819 3701 856
rect 3785 833 3789 916
rect 3890 873 3894 916
rect 3887 861 3894 873
rect 3785 821 3794 833
rect 3694 794 3701 807
rect 3682 788 3701 794
rect 3682 784 3686 788
rect 3785 764 3789 821
rect 3885 784 3889 861
rect 3912 819 3916 876
rect 3920 872 3924 876
rect 3920 864 3938 872
rect 3934 853 3938 864
rect 3905 807 3914 819
rect 3905 784 3909 807
rect 3934 796 3938 841
rect 4011 839 4015 916
rect 4006 827 4015 839
rect 4009 811 4015 827
rect 4031 839 4035 916
rect 4150 873 4154 916
rect 4147 861 4154 873
rect 4031 827 4034 839
rect 4031 811 4037 827
rect 4009 804 4017 811
rect 3925 789 3938 796
rect 3925 784 3929 789
rect 4013 784 4017 804
rect 4023 804 4037 811
rect 4023 784 4027 804
rect 4145 784 4149 861
rect 4172 819 4176 876
rect 4180 872 4184 876
rect 4290 873 4294 916
rect 4180 864 4198 872
rect 4194 853 4198 864
rect 4287 861 4294 873
rect 4165 807 4174 819
rect 4165 784 4169 807
rect 4194 796 4198 841
rect 4185 789 4198 796
rect 4185 784 4189 789
rect 4285 784 4289 861
rect 4312 819 4316 876
rect 4320 872 4324 876
rect 4320 864 4338 872
rect 4334 853 4338 864
rect 4305 807 4314 819
rect 4305 784 4309 807
rect 4334 796 4338 841
rect 4431 833 4435 916
rect 4550 873 4554 916
rect 4547 861 4554 873
rect 4426 821 4435 833
rect 4325 789 4338 796
rect 4325 784 4329 789
rect 4431 764 4435 821
rect 4545 784 4549 861
rect 4572 819 4576 876
rect 4580 872 4584 876
rect 4580 864 4598 872
rect 4594 853 4598 864
rect 4671 862 4675 876
rect 4691 862 4695 876
rect 4659 856 4675 862
rect 4680 856 4695 862
rect 4565 807 4574 819
rect 4565 784 4569 807
rect 4594 796 4598 841
rect 4659 819 4666 856
rect 4680 833 4686 856
rect 4585 789 4598 796
rect 4659 794 4666 807
rect 4585 784 4589 789
rect 4659 788 4678 794
rect 4674 784 4678 788
rect 4682 784 4686 821
rect 4711 819 4715 876
rect 4823 870 4827 876
rect 4823 858 4825 870
rect 4706 807 4715 819
rect 4845 853 4849 916
rect 4950 873 4954 916
rect 4947 861 4954 873
rect 4845 841 4854 853
rect 4704 764 4708 807
rect 4823 790 4825 802
rect 4823 784 4827 790
rect 4845 764 4849 841
rect 4945 784 4949 861
rect 4972 819 4976 876
rect 4980 872 4984 876
rect 4980 864 4998 872
rect 4994 853 4998 864
rect 5071 862 5075 876
rect 5091 862 5095 876
rect 5059 856 5075 862
rect 5080 856 5095 862
rect 4965 807 4974 819
rect 4965 784 4969 807
rect 4994 796 4998 841
rect 5059 819 5066 856
rect 5080 833 5086 856
rect 4985 789 4998 796
rect 5059 794 5066 807
rect 4985 784 4989 789
rect 5059 788 5078 794
rect 5074 784 5078 788
rect 5082 784 5086 821
rect 5111 819 5115 876
rect 5235 871 5239 876
rect 5255 853 5259 876
rect 5265 872 5269 876
rect 5265 867 5278 872
rect 5106 807 5115 819
rect 5104 764 5108 807
rect 5225 792 5235 804
rect 5225 784 5229 792
rect 5255 777 5259 841
rect 5245 771 5259 777
rect 5274 833 5278 867
rect 5385 833 5389 916
rect 5485 853 5489 876
rect 5486 841 5489 853
rect 5385 821 5394 833
rect 5274 776 5278 821
rect 5265 771 5278 776
rect 5245 764 5249 771
rect 5265 764 5269 771
rect 5385 764 5389 821
rect 5480 793 5486 841
rect 5505 819 5509 876
rect 5525 854 5529 876
rect 5545 854 5549 876
rect 5656 872 5660 876
rect 5642 864 5660 872
rect 5525 848 5538 854
rect 5545 853 5565 854
rect 5642 853 5646 864
rect 5545 848 5553 853
rect 5534 819 5538 848
rect 5507 807 5509 819
rect 5505 805 5509 807
rect 5505 798 5518 805
rect 5480 789 5510 793
rect 5506 784 5510 789
rect 5514 784 5518 798
rect 5534 784 5538 807
rect 5553 799 5559 841
rect 5542 792 5559 799
rect 5642 796 5646 841
rect 5664 819 5668 876
rect 5686 873 5690 916
rect 5686 861 5693 873
rect 5666 807 5675 819
rect 5542 784 5546 792
rect 5642 789 5655 796
rect 5651 784 5655 789
rect 5671 784 5675 807
rect 5691 784 5695 861
rect 108 740 112 744
rect 116 740 120 744
rect 124 740 128 744
rect 214 740 218 744
rect 222 740 226 744
rect 244 740 248 744
rect 388 740 392 744
rect 396 740 400 744
rect 404 740 408 744
rect 512 740 516 744
rect 534 740 538 744
rect 542 740 546 744
rect 668 740 672 744
rect 676 740 680 744
rect 684 740 688 744
rect 774 740 778 744
rect 782 740 786 744
rect 804 740 808 744
rect 925 740 929 744
rect 945 740 949 744
rect 965 740 969 744
rect 1088 740 1092 744
rect 1096 740 1100 744
rect 1104 740 1108 744
rect 1191 740 1195 744
rect 1211 740 1215 744
rect 1231 740 1235 744
rect 1368 740 1372 744
rect 1376 740 1380 744
rect 1384 740 1388 744
rect 1471 740 1475 744
rect 1573 740 1577 744
rect 1583 740 1587 744
rect 1748 740 1752 744
rect 1756 740 1760 744
rect 1764 740 1768 744
rect 1888 740 1892 744
rect 1896 740 1900 744
rect 1904 740 1908 744
rect 1992 740 1996 744
rect 2000 740 2004 744
rect 2008 740 2012 744
rect 2131 740 2135 744
rect 2151 740 2155 744
rect 2171 740 2175 744
rect 2271 740 2275 744
rect 2281 740 2285 744
rect 2301 740 2305 744
rect 2411 740 2415 744
rect 2533 740 2537 744
rect 2543 740 2547 744
rect 2645 740 2649 744
rect 2665 740 2669 744
rect 2685 740 2689 744
rect 2773 740 2777 744
rect 2783 740 2787 744
rect 2913 740 2917 744
rect 2923 740 2927 744
rect 3031 740 3035 744
rect 3145 740 3149 744
rect 3273 740 3277 744
rect 3283 740 3287 744
rect 3405 740 3409 744
rect 3425 740 3429 744
rect 3525 740 3529 744
rect 3545 740 3549 744
rect 3652 740 3656 744
rect 3674 740 3678 744
rect 3682 740 3686 744
rect 3785 740 3789 744
rect 3885 740 3889 744
rect 3905 740 3909 744
rect 3925 740 3929 744
rect 4013 740 4017 744
rect 4023 740 4027 744
rect 4145 740 4149 744
rect 4165 740 4169 744
rect 4185 740 4189 744
rect 4285 740 4289 744
rect 4305 740 4309 744
rect 4325 740 4329 744
rect 4431 740 4435 744
rect 4545 740 4549 744
rect 4565 740 4569 744
rect 4585 740 4589 744
rect 4674 740 4678 744
rect 4682 740 4686 744
rect 4704 740 4708 744
rect 4823 740 4827 744
rect 4845 740 4849 744
rect 4945 740 4949 744
rect 4965 740 4969 744
rect 4985 740 4989 744
rect 5074 740 5078 744
rect 5082 740 5086 744
rect 5104 740 5108 744
rect 5225 740 5229 744
rect 5245 740 5249 744
rect 5265 740 5269 744
rect 5385 740 5389 744
rect 5506 740 5510 744
rect 5514 740 5518 744
rect 5534 740 5538 744
rect 5542 740 5546 744
rect 5651 740 5655 744
rect 5671 740 5675 744
rect 5691 740 5695 744
rect 108 716 112 720
rect 116 716 120 720
rect 124 716 128 720
rect 252 716 256 720
rect 274 716 278 720
rect 282 716 286 720
rect 408 716 412 720
rect 416 716 420 720
rect 424 716 428 720
rect 525 716 529 720
rect 545 716 549 720
rect 565 716 569 720
rect 654 716 658 720
rect 662 716 666 720
rect 684 716 688 720
rect 793 716 797 720
rect 803 716 807 720
rect 945 716 949 720
rect 965 716 969 720
rect 985 716 989 720
rect 1108 716 1112 720
rect 1116 716 1120 720
rect 1124 716 1128 720
rect 1214 716 1218 720
rect 1222 716 1226 720
rect 1244 716 1248 720
rect 1372 716 1376 720
rect 1394 716 1398 720
rect 1402 716 1406 720
rect 1512 716 1516 720
rect 1520 716 1524 720
rect 1528 716 1532 720
rect 1665 716 1669 720
rect 1685 716 1689 720
rect 1705 716 1709 720
rect 1828 716 1832 720
rect 1836 716 1840 720
rect 1844 716 1848 720
rect 1934 716 1938 720
rect 1942 716 1946 720
rect 1964 716 1968 720
rect 2085 716 2089 720
rect 2105 716 2109 720
rect 2205 716 2209 720
rect 2225 716 2229 720
rect 2245 716 2249 720
rect 2331 716 2335 720
rect 2341 716 2345 720
rect 2361 716 2365 720
rect 2473 716 2477 720
rect 2483 716 2487 720
rect 2613 716 2617 720
rect 2623 716 2627 720
rect 2725 716 2729 720
rect 2745 716 2749 720
rect 2831 716 2835 720
rect 2851 716 2855 720
rect 2871 716 2875 720
rect 2993 716 2997 720
rect 3003 716 3007 720
rect 3094 716 3098 720
rect 3102 716 3106 720
rect 3124 716 3128 720
rect 3268 716 3272 720
rect 3276 716 3280 720
rect 3284 716 3288 720
rect 3373 716 3377 720
rect 3383 716 3387 720
rect 3505 716 3509 720
rect 3525 716 3529 720
rect 3545 716 3549 720
rect 3633 716 3637 720
rect 3643 716 3647 720
rect 3765 716 3769 720
rect 3785 716 3789 720
rect 3805 716 3809 720
rect 3891 716 3895 720
rect 3911 716 3915 720
rect 3931 716 3935 720
rect 4034 716 4038 720
rect 4042 716 4046 720
rect 4064 716 4068 720
rect 4191 716 4195 720
rect 4211 716 4215 720
rect 4231 716 4235 720
rect 4345 716 4349 720
rect 4452 716 4456 720
rect 4474 716 4478 720
rect 4482 716 4486 720
rect 4585 716 4589 720
rect 4605 716 4609 720
rect 4625 716 4629 720
rect 4725 716 4729 720
rect 4745 716 4749 720
rect 4765 716 4769 720
rect 4871 716 4875 720
rect 4891 716 4895 720
rect 4911 716 4915 720
rect 5011 716 5015 720
rect 5131 716 5135 720
rect 5153 716 5157 720
rect 5265 716 5269 720
rect 5285 716 5289 720
rect 5305 716 5309 720
rect 5391 716 5395 720
rect 5411 716 5415 720
rect 5431 716 5435 720
rect 5545 716 5549 720
rect 5565 716 5569 720
rect 5585 716 5589 720
rect 5671 716 5675 720
rect 5691 716 5695 720
rect 108 599 112 656
rect 85 587 93 599
rect 105 587 112 599
rect 85 544 89 587
rect 116 579 120 656
rect 124 599 128 656
rect 252 653 256 696
rect 245 641 254 653
rect 124 587 134 599
rect 114 560 120 567
rect 105 556 120 560
rect 134 556 140 587
rect 245 584 249 641
rect 274 639 278 676
rect 282 672 286 676
rect 282 666 301 672
rect 294 653 301 666
rect 274 604 280 627
rect 294 604 301 641
rect 265 598 280 604
rect 285 598 301 604
rect 408 599 412 656
rect 265 584 269 598
rect 285 584 289 598
rect 385 587 393 599
rect 405 587 412 599
rect 105 544 109 556
rect 125 552 140 556
rect 125 544 129 552
rect 385 544 389 587
rect 416 579 420 656
rect 424 599 428 656
rect 525 599 529 676
rect 545 653 549 676
rect 565 671 569 676
rect 654 672 658 676
rect 565 664 578 671
rect 545 641 554 653
rect 424 587 434 599
rect 527 587 534 599
rect 414 560 420 567
rect 405 556 420 560
rect 434 556 440 587
rect 405 544 409 556
rect 425 552 440 556
rect 425 544 429 552
rect 530 544 534 587
rect 552 584 556 641
rect 574 619 578 664
rect 639 666 658 672
rect 639 653 646 666
rect 574 596 578 607
rect 639 604 646 641
rect 662 639 666 676
rect 684 653 688 696
rect 793 656 797 676
rect 686 641 695 653
rect 660 604 666 627
rect 639 598 655 604
rect 660 598 675 604
rect 560 588 578 596
rect 560 584 564 588
rect 651 584 655 598
rect 671 584 675 598
rect 691 584 695 641
rect 789 649 797 656
rect 803 656 807 676
rect 803 649 817 656
rect 789 633 795 649
rect 786 621 795 633
rect 791 544 795 621
rect 811 633 817 649
rect 811 621 814 633
rect 811 544 815 621
rect 945 599 949 676
rect 965 653 969 676
rect 985 671 989 676
rect 985 664 998 671
rect 965 641 974 653
rect 947 587 954 599
rect 950 544 954 587
rect 972 584 976 641
rect 994 619 998 664
rect 1214 672 1218 676
rect 1199 666 1218 672
rect 994 596 998 607
rect 1108 599 1112 656
rect 980 588 998 596
rect 980 584 984 588
rect 1085 587 1093 599
rect 1105 587 1112 599
rect 1085 544 1089 587
rect 1116 579 1120 656
rect 1124 599 1128 656
rect 1199 653 1206 666
rect 1199 604 1206 641
rect 1222 639 1226 676
rect 1244 653 1248 696
rect 1372 653 1376 696
rect 1246 641 1255 653
rect 1220 604 1226 627
rect 1124 587 1134 599
rect 1199 598 1215 604
rect 1220 598 1235 604
rect 1114 560 1120 567
rect 1105 556 1120 560
rect 1134 556 1140 587
rect 1211 584 1215 598
rect 1231 584 1235 598
rect 1251 584 1255 641
rect 1365 641 1374 653
rect 1365 584 1369 641
rect 1394 639 1398 676
rect 1402 672 1406 676
rect 1402 666 1421 672
rect 1414 653 1421 666
rect 1394 604 1400 627
rect 1414 604 1421 641
rect 1385 598 1400 604
rect 1405 598 1421 604
rect 1512 599 1516 656
rect 1385 584 1389 598
rect 1405 584 1409 598
rect 1506 587 1516 599
rect 1105 544 1109 556
rect 1125 552 1140 556
rect 1125 544 1129 552
rect 1500 556 1506 587
rect 1520 579 1524 656
rect 1528 599 1532 656
rect 1665 599 1669 676
rect 1685 653 1689 676
rect 1705 671 1709 676
rect 1705 664 1718 671
rect 1685 641 1694 653
rect 1528 587 1535 599
rect 1547 587 1555 599
rect 1667 587 1674 599
rect 1520 560 1526 567
rect 1520 556 1535 560
rect 1500 552 1515 556
rect 1511 544 1515 552
rect 1531 544 1535 556
rect 1551 544 1555 587
rect 1670 544 1674 587
rect 1692 584 1696 641
rect 1714 619 1718 664
rect 1934 672 1938 676
rect 1919 666 1938 672
rect 1714 596 1718 607
rect 1828 599 1832 656
rect 1700 588 1718 596
rect 1700 584 1704 588
rect 1805 587 1813 599
rect 1825 587 1832 599
rect 1805 544 1809 587
rect 1836 579 1840 656
rect 1844 599 1848 656
rect 1919 653 1926 666
rect 1919 604 1926 641
rect 1942 639 1946 676
rect 1964 653 1968 696
rect 1966 641 1975 653
rect 1940 604 1946 627
rect 1844 587 1854 599
rect 1919 598 1935 604
rect 1940 598 1955 604
rect 1834 560 1840 567
rect 1825 556 1840 560
rect 1854 556 1860 587
rect 1931 584 1935 598
rect 1951 584 1955 598
rect 1971 584 1975 641
rect 2085 619 2089 696
rect 2105 619 2109 696
rect 2225 689 2229 696
rect 2245 689 2249 696
rect 2225 683 2239 689
rect 2245 684 2258 689
rect 2205 668 2209 676
rect 2205 656 2215 668
rect 2235 619 2239 683
rect 2254 639 2258 684
rect 2086 607 2101 619
rect 2097 584 2101 607
rect 2105 607 2114 619
rect 2105 584 2109 607
rect 2215 584 2219 589
rect 2235 584 2239 607
rect 2254 593 2258 627
rect 2331 619 2335 676
rect 2341 633 2345 676
rect 2361 670 2365 676
rect 2367 658 2379 670
rect 2341 621 2354 633
rect 2326 607 2335 619
rect 2245 588 2258 593
rect 2245 584 2249 588
rect 1825 544 1829 556
rect 1845 552 1860 556
rect 1845 544 1849 552
rect 2331 544 2335 607
rect 2353 544 2357 621
rect 2375 584 2379 658
rect 2473 656 2477 676
rect 2469 649 2477 656
rect 2483 656 2487 676
rect 2613 656 2617 676
rect 2483 649 2497 656
rect 2469 633 2475 649
rect 2466 621 2475 633
rect 2471 544 2475 621
rect 2491 633 2497 649
rect 2603 649 2617 656
rect 2623 656 2627 676
rect 2623 649 2631 656
rect 2603 633 2609 649
rect 2491 621 2494 633
rect 2606 621 2609 633
rect 2491 544 2495 621
rect 2605 544 2609 621
rect 2625 633 2631 649
rect 2625 621 2634 633
rect 2625 544 2629 621
rect 2725 619 2729 696
rect 2745 619 2749 696
rect 2831 671 2835 676
rect 2822 664 2835 671
rect 2822 619 2826 664
rect 2851 653 2855 676
rect 2846 641 2855 653
rect 2726 607 2741 619
rect 2737 584 2741 607
rect 2745 607 2754 619
rect 2745 584 2749 607
rect 2822 596 2826 607
rect 2822 588 2840 596
rect 2836 584 2840 588
rect 2844 584 2848 641
rect 2871 599 2875 676
rect 2993 656 2997 676
rect 2983 649 2997 656
rect 3003 656 3007 676
rect 3094 672 3098 676
rect 3079 666 3098 672
rect 3003 649 3011 656
rect 3079 653 3086 666
rect 2983 633 2989 649
rect 2986 621 2989 633
rect 2866 587 2873 599
rect 2866 544 2870 587
rect 2985 544 2989 621
rect 3005 633 3011 649
rect 3005 621 3014 633
rect 3005 544 3009 621
rect 3079 604 3086 641
rect 3102 639 3106 676
rect 3124 653 3128 696
rect 3373 656 3377 676
rect 3126 641 3135 653
rect 3100 604 3106 627
rect 3079 598 3095 604
rect 3100 598 3115 604
rect 3091 584 3095 598
rect 3111 584 3115 598
rect 3131 584 3135 641
rect 3268 599 3272 656
rect 3245 587 3253 599
rect 3265 587 3272 599
rect 3245 544 3249 587
rect 3276 579 3280 656
rect 3284 599 3288 656
rect 3369 649 3377 656
rect 3383 656 3387 676
rect 3383 649 3397 656
rect 3369 633 3375 649
rect 3366 621 3375 633
rect 3284 587 3294 599
rect 3274 560 3280 567
rect 3265 556 3280 560
rect 3294 556 3300 587
rect 3265 544 3269 556
rect 3285 552 3300 556
rect 3285 544 3289 552
rect 3371 544 3375 621
rect 3391 633 3397 649
rect 3391 621 3394 633
rect 3391 544 3395 621
rect 3505 599 3509 676
rect 3525 653 3529 676
rect 3545 671 3549 676
rect 3545 664 3558 671
rect 3525 641 3534 653
rect 3507 587 3514 599
rect 3510 544 3514 587
rect 3532 584 3536 641
rect 3554 619 3558 664
rect 3633 656 3637 676
rect 3629 649 3637 656
rect 3643 656 3647 676
rect 3643 649 3657 656
rect 3629 633 3635 649
rect 3626 621 3635 633
rect 3554 596 3558 607
rect 3540 588 3558 596
rect 3540 584 3544 588
rect 3631 544 3635 621
rect 3651 633 3657 649
rect 3651 621 3654 633
rect 3651 544 3655 621
rect 3765 599 3769 676
rect 3785 653 3789 676
rect 3805 671 3809 676
rect 3891 671 3895 676
rect 3805 664 3818 671
rect 3785 641 3794 653
rect 3767 587 3774 599
rect 3770 544 3774 587
rect 3792 584 3796 641
rect 3814 619 3818 664
rect 3882 664 3895 671
rect 3882 619 3886 664
rect 3911 653 3915 676
rect 3906 641 3915 653
rect 3814 596 3818 607
rect 3800 588 3818 596
rect 3882 596 3886 607
rect 3882 588 3900 596
rect 3800 584 3804 588
rect 3896 584 3900 588
rect 3904 584 3908 641
rect 3931 599 3935 676
rect 4034 672 4038 676
rect 4019 666 4038 672
rect 4019 653 4026 666
rect 4019 604 4026 641
rect 4042 639 4046 676
rect 4064 653 4068 696
rect 4191 671 4195 676
rect 4182 664 4195 671
rect 4066 641 4075 653
rect 4040 604 4046 627
rect 3926 587 3933 599
rect 4019 598 4035 604
rect 4040 598 4055 604
rect 3926 544 3930 587
rect 4031 584 4035 598
rect 4051 584 4055 598
rect 4071 584 4075 641
rect 4182 619 4186 664
rect 4211 653 4215 676
rect 4206 641 4215 653
rect 4182 596 4186 607
rect 4182 588 4200 596
rect 4196 584 4200 588
rect 4204 584 4208 641
rect 4231 599 4235 676
rect 4345 639 4349 696
rect 4452 653 4456 696
rect 4445 641 4454 653
rect 4345 627 4354 639
rect 4226 587 4233 599
rect 4226 544 4230 587
rect 4345 544 4349 627
rect 4445 584 4449 641
rect 4474 639 4478 676
rect 4482 672 4486 676
rect 4482 666 4501 672
rect 4494 653 4501 666
rect 4474 604 4480 627
rect 4494 604 4501 641
rect 4465 598 4480 604
rect 4485 598 4501 604
rect 4585 599 4589 676
rect 4605 653 4609 676
rect 4625 671 4629 676
rect 4625 664 4638 671
rect 4605 641 4614 653
rect 4465 584 4469 598
rect 4485 584 4489 598
rect 4587 587 4594 599
rect 4590 544 4594 587
rect 4612 584 4616 641
rect 4634 619 4638 664
rect 4634 596 4638 607
rect 4725 599 4729 676
rect 4745 653 4749 676
rect 4765 671 4769 676
rect 4871 671 4875 676
rect 4765 664 4778 671
rect 4745 641 4754 653
rect 4620 588 4638 596
rect 4620 584 4624 588
rect 4727 587 4734 599
rect 4730 544 4734 587
rect 4752 584 4756 641
rect 4774 619 4778 664
rect 4862 664 4875 671
rect 4862 619 4866 664
rect 4891 653 4895 676
rect 4886 641 4895 653
rect 4774 596 4778 607
rect 4760 588 4778 596
rect 4862 596 4866 607
rect 4862 588 4880 596
rect 4760 584 4764 588
rect 4876 584 4880 588
rect 4884 584 4888 641
rect 4911 599 4915 676
rect 5011 639 5015 696
rect 5006 627 5015 639
rect 4906 587 4913 599
rect 4906 544 4910 587
rect 5011 544 5015 627
rect 5131 619 5135 696
rect 5153 670 5157 676
rect 5155 658 5157 670
rect 5126 607 5135 619
rect 5131 544 5135 607
rect 5155 590 5157 602
rect 5265 599 5269 676
rect 5285 653 5289 676
rect 5305 671 5309 676
rect 5391 671 5395 676
rect 5305 664 5318 671
rect 5285 641 5294 653
rect 5153 584 5157 590
rect 5267 587 5274 599
rect 5270 544 5274 587
rect 5292 584 5296 641
rect 5314 619 5318 664
rect 5382 664 5395 671
rect 5382 619 5386 664
rect 5411 653 5415 676
rect 5406 641 5415 653
rect 5314 596 5318 607
rect 5300 588 5318 596
rect 5382 596 5386 607
rect 5382 588 5400 596
rect 5300 584 5304 588
rect 5396 584 5400 588
rect 5404 584 5408 641
rect 5431 599 5435 676
rect 5545 599 5549 676
rect 5565 653 5569 676
rect 5585 671 5589 676
rect 5585 664 5598 671
rect 5565 641 5574 653
rect 5426 587 5433 599
rect 5547 587 5554 599
rect 5426 544 5430 587
rect 5550 544 5554 587
rect 5572 584 5576 641
rect 5594 619 5598 664
rect 5671 619 5675 696
rect 5691 619 5695 696
rect 5666 607 5675 619
rect 5594 596 5598 607
rect 5580 588 5598 596
rect 5580 584 5584 588
rect 5671 584 5675 607
rect 5679 607 5694 619
rect 5679 584 5683 607
rect 85 500 89 504
rect 105 500 109 504
rect 125 500 129 504
rect 245 500 249 504
rect 265 500 269 504
rect 285 500 289 504
rect 385 500 389 504
rect 405 500 409 504
rect 425 500 429 504
rect 530 500 534 504
rect 552 500 556 504
rect 560 500 564 504
rect 651 500 655 504
rect 671 500 675 504
rect 691 500 695 504
rect 791 500 795 504
rect 811 500 815 504
rect 950 500 954 504
rect 972 500 976 504
rect 980 500 984 504
rect 1085 500 1089 504
rect 1105 500 1109 504
rect 1125 500 1129 504
rect 1211 500 1215 504
rect 1231 500 1235 504
rect 1251 500 1255 504
rect 1365 500 1369 504
rect 1385 500 1389 504
rect 1405 500 1409 504
rect 1511 500 1515 504
rect 1531 500 1535 504
rect 1551 500 1555 504
rect 1670 500 1674 504
rect 1692 500 1696 504
rect 1700 500 1704 504
rect 1805 500 1809 504
rect 1825 500 1829 504
rect 1845 500 1849 504
rect 1931 500 1935 504
rect 1951 500 1955 504
rect 1971 500 1975 504
rect 2097 500 2101 504
rect 2105 500 2109 504
rect 2215 500 2219 504
rect 2235 500 2239 504
rect 2245 500 2249 504
rect 2331 500 2335 504
rect 2353 500 2357 504
rect 2375 500 2379 504
rect 2471 500 2475 504
rect 2491 500 2495 504
rect 2605 500 2609 504
rect 2625 500 2629 504
rect 2737 500 2741 504
rect 2745 500 2749 504
rect 2836 500 2840 504
rect 2844 500 2848 504
rect 2866 500 2870 504
rect 2985 500 2989 504
rect 3005 500 3009 504
rect 3091 500 3095 504
rect 3111 500 3115 504
rect 3131 500 3135 504
rect 3245 500 3249 504
rect 3265 500 3269 504
rect 3285 500 3289 504
rect 3371 500 3375 504
rect 3391 500 3395 504
rect 3510 500 3514 504
rect 3532 500 3536 504
rect 3540 500 3544 504
rect 3631 500 3635 504
rect 3651 500 3655 504
rect 3770 500 3774 504
rect 3792 500 3796 504
rect 3800 500 3804 504
rect 3896 500 3900 504
rect 3904 500 3908 504
rect 3926 500 3930 504
rect 4031 500 4035 504
rect 4051 500 4055 504
rect 4071 500 4075 504
rect 4196 500 4200 504
rect 4204 500 4208 504
rect 4226 500 4230 504
rect 4345 500 4349 504
rect 4445 500 4449 504
rect 4465 500 4469 504
rect 4485 500 4489 504
rect 4590 500 4594 504
rect 4612 500 4616 504
rect 4620 500 4624 504
rect 4730 500 4734 504
rect 4752 500 4756 504
rect 4760 500 4764 504
rect 4876 500 4880 504
rect 4884 500 4888 504
rect 4906 500 4910 504
rect 5011 500 5015 504
rect 5131 500 5135 504
rect 5153 500 5157 504
rect 5270 500 5274 504
rect 5292 500 5296 504
rect 5300 500 5304 504
rect 5396 500 5400 504
rect 5404 500 5408 504
rect 5426 500 5430 504
rect 5550 500 5554 504
rect 5572 500 5576 504
rect 5580 500 5584 504
rect 5671 500 5675 504
rect 5679 500 5683 504
rect 85 476 89 480
rect 105 476 109 480
rect 125 476 129 480
rect 230 476 234 480
rect 252 476 256 480
rect 260 476 264 480
rect 390 476 394 480
rect 412 476 416 480
rect 420 476 424 480
rect 525 476 529 480
rect 545 476 549 480
rect 565 476 569 480
rect 661 476 665 480
rect 683 476 687 480
rect 705 476 709 480
rect 805 476 809 480
rect 825 476 829 480
rect 845 476 849 480
rect 945 476 949 480
rect 965 476 969 480
rect 985 476 989 480
rect 1071 476 1075 480
rect 1091 476 1095 480
rect 1111 476 1115 480
rect 1235 476 1239 480
rect 1255 476 1259 480
rect 1265 476 1269 480
rect 1365 476 1369 480
rect 1385 476 1389 480
rect 1405 476 1409 480
rect 1525 476 1529 480
rect 1630 476 1634 480
rect 1652 476 1656 480
rect 1660 476 1664 480
rect 1761 476 1765 480
rect 1783 476 1787 480
rect 1805 476 1809 480
rect 1891 476 1895 480
rect 1899 476 1903 480
rect 2031 476 2035 480
rect 2150 476 2154 480
rect 2172 476 2176 480
rect 2180 476 2184 480
rect 2285 476 2289 480
rect 2305 476 2309 480
rect 2325 476 2329 480
rect 2425 476 2429 480
rect 2525 476 2529 480
rect 2545 476 2549 480
rect 2565 476 2569 480
rect 2656 476 2660 480
rect 2664 476 2668 480
rect 2686 476 2690 480
rect 2805 476 2809 480
rect 2917 476 2921 480
rect 2925 476 2929 480
rect 3011 476 3015 480
rect 3125 476 3129 480
rect 3145 476 3149 480
rect 3165 476 3169 480
rect 3271 476 3275 480
rect 3291 476 3295 480
rect 3311 476 3315 480
rect 3425 476 3429 480
rect 3536 476 3540 480
rect 3544 476 3548 480
rect 3566 476 3570 480
rect 3671 476 3675 480
rect 3691 476 3695 480
rect 3711 476 3715 480
rect 3825 476 3829 480
rect 3845 476 3849 480
rect 3865 476 3869 480
rect 3951 476 3955 480
rect 3971 476 3975 480
rect 4105 476 4109 480
rect 4125 476 4129 480
rect 4145 476 4149 480
rect 4250 476 4254 480
rect 4272 476 4276 480
rect 4280 476 4284 480
rect 4385 476 4389 480
rect 4485 476 4489 480
rect 4505 476 4509 480
rect 4610 476 4614 480
rect 4632 476 4636 480
rect 4640 476 4644 480
rect 4745 476 4749 480
rect 4850 476 4854 480
rect 4872 476 4876 480
rect 4880 476 4884 480
rect 4971 476 5005 480
rect 5021 476 5025 480
rect 5031 476 5035 480
rect 5150 476 5154 480
rect 5172 476 5176 480
rect 5180 476 5184 480
rect 5296 476 5300 480
rect 5304 476 5308 480
rect 5326 476 5330 480
rect 5465 476 5469 480
rect 5485 476 5489 480
rect 5505 476 5509 480
rect 5596 476 5600 480
rect 5604 476 5608 480
rect 5626 476 5630 480
rect 5731 476 5735 480
rect 5751 476 5755 480
rect 85 393 89 436
rect 105 424 109 436
rect 125 428 129 436
rect 125 424 140 428
rect 105 420 120 424
rect 114 413 120 420
rect 85 381 93 393
rect 105 381 112 393
rect 108 324 112 381
rect 116 324 120 401
rect 134 393 140 424
rect 230 393 234 436
rect 124 381 134 393
rect 227 381 234 393
rect 124 324 128 381
rect 225 304 229 381
rect 252 339 256 396
rect 260 392 264 396
rect 390 393 394 436
rect 260 384 278 392
rect 274 373 278 384
rect 387 381 394 393
rect 245 327 254 339
rect 245 304 249 327
rect 274 316 278 361
rect 265 309 278 316
rect 265 304 269 309
rect 385 304 389 381
rect 412 339 416 396
rect 420 392 424 396
rect 525 393 529 436
rect 545 424 549 436
rect 565 428 569 436
rect 565 424 580 428
rect 545 420 560 424
rect 554 413 560 420
rect 420 384 438 392
rect 434 373 438 384
rect 525 381 533 393
rect 545 381 552 393
rect 405 327 414 339
rect 405 304 409 327
rect 434 316 438 361
rect 548 324 552 381
rect 556 324 560 401
rect 574 393 580 424
rect 564 381 574 393
rect 564 324 568 381
rect 425 309 438 316
rect 425 304 429 309
rect 661 322 665 396
rect 683 359 687 436
rect 705 373 709 436
rect 805 393 809 436
rect 825 424 829 436
rect 845 428 849 436
rect 845 424 860 428
rect 825 420 840 424
rect 834 413 840 420
rect 805 381 813 393
rect 825 381 832 393
rect 705 361 714 373
rect 686 347 699 359
rect 661 310 673 322
rect 675 304 679 310
rect 695 304 699 347
rect 705 304 709 361
rect 828 324 832 381
rect 836 324 840 401
rect 854 393 860 424
rect 1071 428 1075 436
rect 1060 424 1075 428
rect 1091 424 1095 436
rect 844 381 854 393
rect 844 324 848 381
rect 945 339 949 396
rect 965 382 969 396
rect 985 382 989 396
rect 1060 393 1066 424
rect 1080 420 1095 424
rect 1080 413 1086 420
rect 965 376 980 382
rect 985 376 1001 382
rect 1066 381 1076 393
rect 974 353 980 376
rect 945 327 954 339
rect 952 284 956 327
rect 974 304 978 341
rect 994 339 1001 376
rect 994 314 1001 327
rect 1072 324 1076 381
rect 1080 324 1084 401
rect 1111 393 1115 436
rect 1088 381 1095 393
rect 1107 381 1115 393
rect 1235 391 1239 396
rect 1088 324 1092 381
rect 1255 373 1259 396
rect 1265 392 1269 396
rect 1365 393 1369 436
rect 1385 424 1389 436
rect 1405 428 1409 436
rect 1405 424 1420 428
rect 1385 420 1400 424
rect 1394 413 1400 420
rect 1265 387 1278 392
rect 982 308 1001 314
rect 982 304 986 308
rect 1225 312 1235 324
rect 1225 304 1229 312
rect 1255 297 1259 361
rect 1245 291 1259 297
rect 1274 353 1278 387
rect 1365 381 1373 393
rect 1385 381 1392 393
rect 1274 296 1278 341
rect 1388 324 1392 381
rect 1396 324 1400 401
rect 1414 393 1420 424
rect 1404 381 1414 393
rect 1404 324 1408 381
rect 1525 353 1529 436
rect 1630 393 1634 436
rect 1627 381 1634 393
rect 1525 341 1534 353
rect 1265 291 1278 296
rect 1245 284 1249 291
rect 1265 284 1269 291
rect 1525 284 1529 341
rect 1625 304 1629 381
rect 1652 339 1656 396
rect 1660 392 1664 396
rect 1660 384 1678 392
rect 1674 373 1678 384
rect 1645 327 1654 339
rect 1645 304 1649 327
rect 1674 316 1678 361
rect 1665 309 1678 316
rect 1761 322 1765 396
rect 1783 359 1787 436
rect 1805 373 1809 436
rect 1891 373 1895 396
rect 1805 361 1814 373
rect 1886 361 1895 373
rect 1899 373 1903 396
rect 1899 361 1914 373
rect 1786 347 1799 359
rect 1761 310 1773 322
rect 1665 304 1669 309
rect 1775 304 1779 310
rect 1795 304 1799 347
rect 1805 304 1809 361
rect 1891 284 1895 361
rect 1911 284 1915 361
rect 2031 353 2035 436
rect 2150 393 2154 436
rect 2147 381 2154 393
rect 2026 341 2035 353
rect 2031 284 2035 341
rect 2145 304 2149 381
rect 2172 339 2176 396
rect 2180 392 2184 396
rect 2180 384 2198 392
rect 2194 373 2198 384
rect 2165 327 2174 339
rect 2165 304 2169 327
rect 2194 316 2198 361
rect 2285 339 2289 396
rect 2305 382 2309 396
rect 2325 382 2329 396
rect 2305 376 2320 382
rect 2325 376 2341 382
rect 2314 353 2320 376
rect 2285 327 2294 339
rect 2185 309 2198 316
rect 2185 304 2189 309
rect 2292 284 2296 327
rect 2314 304 2318 341
rect 2334 339 2341 376
rect 2425 353 2429 436
rect 2525 393 2529 436
rect 2545 424 2549 436
rect 2565 428 2569 436
rect 2565 424 2580 428
rect 2545 420 2560 424
rect 2554 413 2560 420
rect 2525 381 2533 393
rect 2545 381 2552 393
rect 2425 341 2434 353
rect 2334 314 2341 327
rect 2322 308 2341 314
rect 2322 304 2326 308
rect 2425 284 2429 341
rect 2548 324 2552 381
rect 2556 324 2560 401
rect 2574 393 2580 424
rect 2564 381 2574 393
rect 2656 392 2660 396
rect 2642 384 2660 392
rect 2564 324 2568 381
rect 2642 373 2646 384
rect 2642 316 2646 361
rect 2664 339 2668 396
rect 2686 393 2690 436
rect 2686 381 2693 393
rect 2666 327 2675 339
rect 2642 309 2655 316
rect 2651 304 2655 309
rect 2671 304 2675 327
rect 2691 304 2695 381
rect 2805 353 2809 436
rect 2917 373 2921 396
rect 2906 361 2921 373
rect 2925 373 2929 396
rect 2925 361 2934 373
rect 2805 341 2814 353
rect 2805 284 2809 341
rect 2905 284 2909 361
rect 2925 284 2929 361
rect 3011 353 3015 436
rect 3006 341 3015 353
rect 3011 284 3015 341
rect 3125 339 3129 396
rect 3145 382 3149 396
rect 3165 382 3169 396
rect 3271 382 3275 396
rect 3291 382 3295 396
rect 3145 376 3160 382
rect 3165 376 3181 382
rect 3154 353 3160 376
rect 3125 327 3134 339
rect 3132 284 3136 327
rect 3154 304 3158 341
rect 3174 339 3181 376
rect 3259 376 3275 382
rect 3280 376 3295 382
rect 3259 339 3266 376
rect 3280 353 3286 376
rect 3174 314 3181 327
rect 3162 308 3181 314
rect 3259 314 3266 327
rect 3259 308 3278 314
rect 3162 304 3166 308
rect 3274 304 3278 308
rect 3282 304 3286 341
rect 3311 339 3315 396
rect 3306 327 3315 339
rect 3425 353 3429 436
rect 3536 392 3540 396
rect 3522 384 3540 392
rect 3522 373 3526 384
rect 3425 341 3434 353
rect 3304 284 3308 327
rect 3425 284 3429 341
rect 3522 316 3526 361
rect 3544 339 3548 396
rect 3566 393 3570 436
rect 3566 381 3573 393
rect 3671 382 3675 396
rect 3691 382 3695 396
rect 3546 327 3555 339
rect 3522 309 3535 316
rect 3531 304 3535 309
rect 3551 304 3555 327
rect 3571 304 3575 381
rect 3659 376 3675 382
rect 3680 376 3695 382
rect 3659 339 3666 376
rect 3680 353 3686 376
rect 3659 314 3666 327
rect 3659 308 3678 314
rect 3674 304 3678 308
rect 3682 304 3686 341
rect 3711 339 3715 396
rect 3825 393 3829 436
rect 3845 424 3849 436
rect 3865 428 3869 436
rect 3865 424 3880 428
rect 3845 420 3860 424
rect 3854 413 3860 420
rect 3825 381 3833 393
rect 3845 381 3852 393
rect 3706 327 3715 339
rect 3704 284 3708 327
rect 3848 324 3852 381
rect 3856 324 3860 401
rect 3874 393 3880 424
rect 3864 381 3874 393
rect 3864 324 3868 381
rect 3951 359 3955 436
rect 3946 347 3955 359
rect 3949 331 3955 347
rect 3971 359 3975 436
rect 4105 393 4109 436
rect 4125 424 4129 436
rect 4145 428 4149 436
rect 4145 424 4160 428
rect 4125 420 4140 424
rect 4134 413 4140 420
rect 4105 381 4113 393
rect 4125 381 4132 393
rect 3971 347 3974 359
rect 3971 331 3977 347
rect 3949 324 3957 331
rect 3953 304 3957 324
rect 3963 324 3977 331
rect 4128 324 4132 381
rect 4136 324 4140 401
rect 4154 393 4160 424
rect 4250 393 4254 436
rect 4144 381 4154 393
rect 4247 381 4254 393
rect 4144 324 4148 381
rect 3963 304 3967 324
rect 4245 304 4249 381
rect 4272 339 4276 396
rect 4280 392 4284 396
rect 4280 384 4298 392
rect 4294 373 4298 384
rect 4265 327 4274 339
rect 4265 304 4269 327
rect 4294 316 4298 361
rect 4285 309 4298 316
rect 4385 353 4389 436
rect 4485 359 4489 436
rect 4385 341 4394 353
rect 4486 347 4489 359
rect 4285 304 4289 309
rect 4385 284 4389 341
rect 4483 331 4489 347
rect 4505 359 4509 436
rect 4610 393 4614 436
rect 4607 381 4614 393
rect 4505 347 4514 359
rect 4505 331 4511 347
rect 4483 324 4497 331
rect 4493 304 4497 324
rect 4503 324 4511 331
rect 4503 304 4507 324
rect 4605 304 4609 381
rect 4632 339 4636 396
rect 4640 392 4644 396
rect 4640 384 4658 392
rect 4654 373 4658 384
rect 4625 327 4634 339
rect 4625 304 4629 327
rect 4654 316 4658 361
rect 4645 309 4658 316
rect 4745 353 4749 436
rect 4850 393 4854 436
rect 4971 468 4975 476
rect 4991 468 4995 472
rect 5001 468 5005 476
rect 4971 424 4975 428
rect 4963 420 4975 424
rect 4847 381 4854 393
rect 4745 341 4754 353
rect 4645 304 4649 309
rect 4745 284 4749 341
rect 4845 304 4849 381
rect 4872 339 4876 396
rect 4880 392 4884 396
rect 4880 384 4898 392
rect 4894 373 4898 384
rect 4865 327 4874 339
rect 4865 304 4869 327
rect 4894 316 4898 361
rect 4963 339 4967 420
rect 4991 383 4995 388
rect 5001 384 5005 388
rect 4982 379 4995 383
rect 4982 373 4987 379
rect 5021 374 5025 396
rect 4995 370 5025 374
rect 5031 373 5035 396
rect 5150 393 5154 436
rect 5147 381 5154 393
rect 4885 309 4898 316
rect 4885 304 4889 309
rect 4963 301 4967 327
rect 4981 330 4986 361
rect 5031 361 5034 373
rect 4981 324 4995 330
rect 4991 312 4995 324
rect 5001 312 5005 358
rect 5021 312 5025 316
rect 5031 312 5035 361
rect 4963 296 4975 301
rect 4971 292 4975 296
rect 5145 304 5149 381
rect 5172 339 5176 396
rect 5180 392 5184 396
rect 5296 392 5300 396
rect 5180 384 5198 392
rect 5194 373 5198 384
rect 5282 384 5300 392
rect 5282 373 5286 384
rect 5165 327 5174 339
rect 5165 304 5169 327
rect 5194 316 5198 361
rect 5185 309 5198 316
rect 5282 316 5286 361
rect 5304 339 5308 396
rect 5326 393 5330 436
rect 5326 381 5333 393
rect 5306 327 5315 339
rect 5282 309 5295 316
rect 5185 304 5189 309
rect 5291 304 5295 309
rect 5311 304 5315 327
rect 5331 304 5335 381
rect 5465 339 5469 396
rect 5485 382 5489 396
rect 5505 382 5509 396
rect 5596 392 5600 396
rect 5582 384 5600 392
rect 5485 376 5500 382
rect 5505 376 5521 382
rect 5494 353 5500 376
rect 5465 327 5474 339
rect 4971 264 4975 272
rect 4991 268 4995 272
rect 5001 268 5005 272
rect 5021 264 5025 272
rect 5031 268 5035 272
rect 5472 284 5476 327
rect 5494 304 5498 341
rect 5514 339 5521 376
rect 5582 373 5586 384
rect 5514 314 5521 327
rect 5502 308 5521 314
rect 5582 316 5586 361
rect 5604 339 5608 396
rect 5626 393 5630 436
rect 5626 381 5633 393
rect 5606 327 5615 339
rect 5582 309 5595 316
rect 5502 304 5506 308
rect 5591 304 5595 309
rect 5611 304 5615 327
rect 5631 304 5635 381
rect 5731 359 5735 436
rect 5726 347 5735 359
rect 5729 331 5735 347
rect 5751 359 5755 436
rect 5751 347 5754 359
rect 5751 331 5757 347
rect 5729 324 5737 331
rect 5733 304 5737 324
rect 5743 324 5757 331
rect 5743 304 5747 324
rect 108 260 112 264
rect 116 260 120 264
rect 124 260 128 264
rect 225 260 229 264
rect 245 260 249 264
rect 265 260 269 264
rect 385 260 389 264
rect 405 260 409 264
rect 425 260 429 264
rect 548 260 552 264
rect 556 260 560 264
rect 564 260 568 264
rect 675 260 679 264
rect 695 260 699 264
rect 705 260 709 264
rect 828 260 832 264
rect 836 260 840 264
rect 844 260 848 264
rect 952 260 956 264
rect 974 260 978 264
rect 982 260 986 264
rect 1072 260 1076 264
rect 1080 260 1084 264
rect 1088 260 1092 264
rect 1225 260 1229 264
rect 1245 260 1249 264
rect 1265 260 1269 264
rect 1388 260 1392 264
rect 1396 260 1400 264
rect 1404 260 1408 264
rect 1525 260 1529 264
rect 1625 260 1629 264
rect 1645 260 1649 264
rect 1665 260 1669 264
rect 1775 260 1779 264
rect 1795 260 1799 264
rect 1805 260 1809 264
rect 1891 260 1895 264
rect 1911 260 1915 264
rect 2031 260 2035 264
rect 2145 260 2149 264
rect 2165 260 2169 264
rect 2185 260 2189 264
rect 2292 260 2296 264
rect 2314 260 2318 264
rect 2322 260 2326 264
rect 2425 260 2429 264
rect 2548 260 2552 264
rect 2556 260 2560 264
rect 2564 260 2568 264
rect 2651 260 2655 264
rect 2671 260 2675 264
rect 2691 260 2695 264
rect 2805 260 2809 264
rect 2905 260 2909 264
rect 2925 260 2929 264
rect 3011 260 3015 264
rect 3132 260 3136 264
rect 3154 260 3158 264
rect 3162 260 3166 264
rect 3274 260 3278 264
rect 3282 260 3286 264
rect 3304 260 3308 264
rect 3425 260 3429 264
rect 3531 260 3535 264
rect 3551 260 3555 264
rect 3571 260 3575 264
rect 3674 260 3678 264
rect 3682 260 3686 264
rect 3704 260 3708 264
rect 3848 260 3852 264
rect 3856 260 3860 264
rect 3864 260 3868 264
rect 3953 260 3957 264
rect 3963 260 3967 264
rect 4128 260 4132 264
rect 4136 260 4140 264
rect 4144 260 4148 264
rect 4245 260 4249 264
rect 4265 260 4269 264
rect 4285 260 4289 264
rect 4385 260 4389 264
rect 4493 260 4497 264
rect 4503 260 4507 264
rect 4605 260 4609 264
rect 4625 260 4629 264
rect 4645 260 4649 264
rect 4745 260 4749 264
rect 4845 260 4849 264
rect 4865 260 4869 264
rect 4885 260 4889 264
rect 4971 260 5025 264
rect 5145 260 5149 264
rect 5165 260 5169 264
rect 5185 260 5189 264
rect 5291 260 5295 264
rect 5311 260 5315 264
rect 5331 260 5335 264
rect 5472 260 5476 264
rect 5494 260 5498 264
rect 5502 260 5506 264
rect 5591 260 5595 264
rect 5611 260 5615 264
rect 5631 260 5635 264
rect 5733 260 5737 264
rect 5743 260 5747 264
rect 108 236 112 240
rect 116 236 120 240
rect 124 236 128 240
rect 214 236 218 240
rect 222 236 226 240
rect 244 236 248 240
rect 392 236 396 240
rect 414 236 418 240
rect 422 236 426 240
rect 525 236 529 240
rect 545 236 549 240
rect 565 236 569 240
rect 651 236 655 240
rect 671 236 675 240
rect 691 236 695 240
rect 828 236 832 240
rect 836 236 840 240
rect 844 236 848 240
rect 931 236 935 240
rect 1031 236 1035 240
rect 1051 236 1055 240
rect 1071 236 1075 240
rect 1174 236 1178 240
rect 1182 236 1186 240
rect 1204 236 1208 240
rect 1311 236 1315 240
rect 1331 236 1335 240
rect 1431 236 1435 240
rect 1441 236 1445 240
rect 1461 236 1465 240
rect 1585 236 1589 240
rect 1685 236 1689 240
rect 1705 236 1709 240
rect 1725 236 1729 240
rect 1833 236 1837 240
rect 1843 236 1847 240
rect 1932 236 1936 240
rect 1940 236 1944 240
rect 1948 236 1952 240
rect 2128 236 2132 240
rect 2136 236 2140 240
rect 2144 236 2148 240
rect 2231 236 2235 240
rect 2253 236 2257 240
rect 2373 236 2377 240
rect 2383 236 2387 240
rect 2471 236 2475 240
rect 2481 236 2485 240
rect 2501 236 2505 240
rect 2632 236 2636 240
rect 2654 236 2658 240
rect 2662 236 2666 240
rect 2775 236 2779 240
rect 2795 236 2799 240
rect 2805 236 2809 240
rect 2913 236 2917 240
rect 2923 236 2927 240
rect 3053 236 3057 240
rect 3063 236 3067 240
rect 3188 236 3192 240
rect 3196 236 3200 240
rect 3204 236 3208 240
rect 3305 236 3309 240
rect 3391 236 3395 240
rect 3411 236 3415 240
rect 3431 236 3435 240
rect 3545 236 3549 240
rect 3653 236 3657 240
rect 3663 236 3667 240
rect 3763 236 3767 240
rect 3785 236 3789 240
rect 3871 236 3875 240
rect 3893 236 3897 240
rect 4013 236 4017 240
rect 4023 236 4027 240
rect 4131 236 4135 240
rect 4141 236 4145 240
rect 4161 236 4165 240
rect 4305 236 4309 240
rect 4325 236 4329 240
rect 4413 236 4417 240
rect 4423 236 4427 240
rect 4568 236 4572 240
rect 4576 236 4580 240
rect 4584 236 4588 240
rect 4705 236 4709 240
rect 4725 236 4729 240
rect 4745 236 4749 240
rect 4833 236 4837 240
rect 4843 236 4847 240
rect 4965 236 4969 240
rect 4985 236 4989 240
rect 5005 236 5009 240
rect 5091 236 5095 240
rect 5111 236 5115 240
rect 5233 236 5237 240
rect 5243 236 5247 240
rect 5331 236 5385 240
rect 5491 236 5495 240
rect 5605 236 5609 240
rect 5693 236 5697 240
rect 5703 236 5707 240
rect 214 192 218 196
rect 199 186 218 192
rect 108 119 112 176
rect 85 107 93 119
rect 105 107 112 119
rect 85 64 89 107
rect 116 99 120 176
rect 124 119 128 176
rect 199 173 206 186
rect 199 124 206 161
rect 222 159 226 196
rect 244 173 248 216
rect 392 173 396 216
rect 246 161 255 173
rect 220 124 226 147
rect 124 107 134 119
rect 199 118 215 124
rect 220 118 235 124
rect 114 80 120 87
rect 105 76 120 80
rect 134 76 140 107
rect 211 104 215 118
rect 231 104 235 118
rect 251 104 255 161
rect 385 161 394 173
rect 385 104 389 161
rect 414 159 418 196
rect 422 192 426 196
rect 422 186 441 192
rect 434 173 441 186
rect 414 124 420 147
rect 434 124 441 161
rect 405 118 420 124
rect 425 118 441 124
rect 525 119 529 196
rect 545 173 549 196
rect 565 191 569 196
rect 651 191 655 196
rect 565 184 578 191
rect 545 161 554 173
rect 405 104 409 118
rect 425 104 429 118
rect 527 107 534 119
rect 105 64 109 76
rect 125 72 140 76
rect 125 64 129 72
rect 530 64 534 107
rect 552 104 556 161
rect 574 139 578 184
rect 642 184 655 191
rect 642 139 646 184
rect 671 173 675 196
rect 666 161 675 173
rect 574 116 578 127
rect 560 108 578 116
rect 642 116 646 127
rect 642 108 660 116
rect 560 104 564 108
rect 656 104 660 108
rect 664 104 668 161
rect 691 119 695 196
rect 828 119 832 176
rect 686 107 693 119
rect 805 107 813 119
rect 825 107 832 119
rect 686 64 690 107
rect 805 64 809 107
rect 836 99 840 176
rect 844 119 848 176
rect 931 159 935 216
rect 1031 191 1035 196
rect 926 147 935 159
rect 844 107 854 119
rect 834 80 840 87
rect 825 76 840 80
rect 854 76 860 107
rect 825 64 829 76
rect 845 72 860 76
rect 845 64 849 72
rect 931 64 935 147
rect 1022 184 1035 191
rect 1022 139 1026 184
rect 1051 173 1055 196
rect 1046 161 1055 173
rect 1022 116 1026 127
rect 1022 108 1040 116
rect 1036 104 1040 108
rect 1044 104 1048 161
rect 1071 119 1075 196
rect 1174 192 1178 196
rect 1159 186 1178 192
rect 1159 173 1166 186
rect 1159 124 1166 161
rect 1182 159 1186 196
rect 1204 173 1208 216
rect 1206 161 1215 173
rect 1180 124 1186 147
rect 1066 107 1073 119
rect 1159 118 1175 124
rect 1180 118 1195 124
rect 1066 64 1070 107
rect 1171 104 1175 118
rect 1191 104 1195 118
rect 1211 104 1215 161
rect 1311 139 1315 216
rect 1331 139 1335 216
rect 1431 139 1435 196
rect 1441 153 1445 196
rect 1461 190 1465 196
rect 1467 178 1479 190
rect 1441 141 1454 153
rect 1306 127 1315 139
rect 1311 104 1315 127
rect 1319 127 1334 139
rect 1426 127 1435 139
rect 1319 104 1323 127
rect 1431 64 1435 127
rect 1453 64 1457 141
rect 1475 104 1479 178
rect 1585 159 1589 216
rect 1585 147 1594 159
rect 1585 64 1589 147
rect 1685 119 1689 196
rect 1705 173 1709 196
rect 1725 191 1729 196
rect 1725 184 1738 191
rect 1705 161 1714 173
rect 1687 107 1694 119
rect 1690 64 1694 107
rect 1712 104 1716 161
rect 1734 139 1738 184
rect 1833 176 1837 196
rect 1823 169 1837 176
rect 1843 176 1847 196
rect 1843 169 1851 176
rect 1823 153 1829 169
rect 1826 141 1829 153
rect 1734 116 1738 127
rect 1720 108 1738 116
rect 1720 104 1724 108
rect 1825 64 1829 141
rect 1845 153 1851 169
rect 1845 141 1854 153
rect 1845 64 1849 141
rect 1932 119 1936 176
rect 1926 107 1936 119
rect 1920 76 1926 107
rect 1940 99 1944 176
rect 1948 119 1952 176
rect 2128 119 2132 176
rect 1948 107 1955 119
rect 1967 107 1975 119
rect 1940 80 1946 87
rect 1940 76 1955 80
rect 1920 72 1935 76
rect 1931 64 1935 72
rect 1951 64 1955 76
rect 1971 64 1975 107
rect 2105 107 2113 119
rect 2125 107 2132 119
rect 2105 64 2109 107
rect 2136 99 2140 176
rect 2144 119 2148 176
rect 2231 139 2235 216
rect 2253 190 2257 196
rect 2255 178 2257 190
rect 2373 176 2377 196
rect 2363 169 2377 176
rect 2383 176 2387 196
rect 2383 169 2391 176
rect 2363 153 2369 169
rect 2366 141 2369 153
rect 2226 127 2235 139
rect 2144 107 2154 119
rect 2134 80 2140 87
rect 2125 76 2140 80
rect 2154 76 2160 107
rect 2125 64 2129 76
rect 2145 72 2160 76
rect 2145 64 2149 72
rect 2231 64 2235 127
rect 2255 110 2257 122
rect 2253 104 2257 110
rect 2365 64 2369 141
rect 2385 153 2391 169
rect 2385 141 2394 153
rect 2385 64 2389 141
rect 2471 139 2475 196
rect 2481 153 2485 196
rect 2501 190 2505 196
rect 2507 178 2519 190
rect 2481 141 2494 153
rect 2466 127 2475 139
rect 2471 64 2475 127
rect 2493 64 2497 141
rect 2515 104 2519 178
rect 2632 173 2636 216
rect 2625 161 2634 173
rect 2625 104 2629 161
rect 2654 159 2658 196
rect 2662 192 2666 196
rect 2662 186 2681 192
rect 2775 190 2779 196
rect 2674 173 2681 186
rect 2761 178 2773 190
rect 2654 124 2660 147
rect 2674 124 2681 161
rect 2645 118 2660 124
rect 2665 118 2681 124
rect 2645 104 2649 118
rect 2665 104 2669 118
rect 2761 104 2765 178
rect 2795 153 2799 196
rect 2786 141 2799 153
rect 2783 64 2787 141
rect 2805 139 2809 196
rect 2913 176 2917 196
rect 2909 169 2917 176
rect 2923 176 2927 196
rect 3053 176 3057 196
rect 2923 169 2937 176
rect 2909 153 2915 169
rect 2906 141 2915 153
rect 2805 127 2814 139
rect 2805 64 2809 127
rect 2911 64 2915 141
rect 2931 153 2937 169
rect 3043 169 3057 176
rect 3063 176 3067 196
rect 3063 169 3071 176
rect 3043 153 3049 169
rect 2931 141 2934 153
rect 3046 141 3049 153
rect 2931 64 2935 141
rect 3045 64 3049 141
rect 3065 153 3071 169
rect 3065 141 3074 153
rect 3065 64 3069 141
rect 3188 119 3192 176
rect 3165 107 3173 119
rect 3185 107 3192 119
rect 3165 64 3169 107
rect 3196 99 3200 176
rect 3204 119 3208 176
rect 3305 159 3309 216
rect 3391 191 3395 196
rect 3382 184 3395 191
rect 3305 147 3314 159
rect 3204 107 3214 119
rect 3194 80 3200 87
rect 3185 76 3200 80
rect 3214 76 3220 107
rect 3185 64 3189 76
rect 3205 72 3220 76
rect 3205 64 3209 72
rect 3305 64 3309 147
rect 3382 139 3386 184
rect 3411 173 3415 196
rect 3406 161 3415 173
rect 3382 116 3386 127
rect 3382 108 3400 116
rect 3396 104 3400 108
rect 3404 104 3408 161
rect 3431 119 3435 196
rect 3545 159 3549 216
rect 3653 176 3657 196
rect 3643 169 3657 176
rect 3663 176 3667 196
rect 3763 190 3767 196
rect 3763 178 3765 190
rect 3663 169 3671 176
rect 3545 147 3554 159
rect 3643 153 3649 169
rect 3426 107 3433 119
rect 3426 64 3430 107
rect 3545 64 3549 147
rect 3646 141 3649 153
rect 3645 64 3649 141
rect 3665 153 3671 169
rect 3665 141 3674 153
rect 3665 64 3669 141
rect 3785 139 3789 216
rect 3871 139 3875 216
rect 3893 190 3897 196
rect 3895 178 3897 190
rect 4013 176 4017 196
rect 4003 169 4017 176
rect 4023 176 4027 196
rect 4023 169 4031 176
rect 4003 153 4009 169
rect 4006 141 4009 153
rect 3785 127 3794 139
rect 3866 127 3875 139
rect 3763 110 3765 122
rect 3763 104 3767 110
rect 3785 64 3789 127
rect 3871 64 3875 127
rect 3895 110 3897 122
rect 3893 104 3897 110
rect 4005 64 4009 141
rect 4025 153 4031 169
rect 4025 141 4034 153
rect 4025 64 4029 141
rect 4131 139 4135 196
rect 4141 153 4145 196
rect 4161 190 4165 196
rect 4167 178 4179 190
rect 4141 141 4154 153
rect 4126 127 4135 139
rect 4131 64 4135 127
rect 4153 64 4157 141
rect 4175 104 4179 178
rect 4305 139 4309 216
rect 4325 139 4329 216
rect 4413 176 4417 196
rect 4409 169 4417 176
rect 4423 176 4427 196
rect 4423 169 4437 176
rect 4409 153 4415 169
rect 4406 141 4415 153
rect 4306 127 4321 139
rect 4317 104 4321 127
rect 4325 127 4334 139
rect 4325 104 4329 127
rect 4411 64 4415 141
rect 4431 153 4437 169
rect 4431 141 4434 153
rect 4431 64 4435 141
rect 4568 119 4572 176
rect 4545 107 4553 119
rect 4565 107 4572 119
rect 4545 64 4549 107
rect 4576 99 4580 176
rect 4584 119 4588 176
rect 4705 119 4709 196
rect 4725 173 4729 196
rect 4745 191 4749 196
rect 4745 184 4758 191
rect 4725 161 4734 173
rect 4584 107 4594 119
rect 4707 107 4714 119
rect 4574 80 4580 87
rect 4565 76 4580 80
rect 4594 76 4600 107
rect 4565 64 4569 76
rect 4585 72 4600 76
rect 4585 64 4589 72
rect 4710 64 4714 107
rect 4732 104 4736 161
rect 4754 139 4758 184
rect 4833 176 4837 196
rect 4829 169 4837 176
rect 4843 176 4847 196
rect 4843 169 4857 176
rect 4829 153 4835 169
rect 4826 141 4835 153
rect 4754 116 4758 127
rect 4740 108 4758 116
rect 4740 104 4744 108
rect 4831 64 4835 141
rect 4851 153 4857 169
rect 4851 141 4854 153
rect 4851 64 4855 141
rect 4965 119 4969 196
rect 4985 173 4989 196
rect 5005 191 5009 196
rect 5005 184 5018 191
rect 4985 161 4994 173
rect 4967 107 4974 119
rect 4970 64 4974 107
rect 4992 104 4996 161
rect 5014 139 5018 184
rect 5091 139 5095 216
rect 5111 139 5115 216
rect 5331 228 5335 236
rect 5351 228 5355 232
rect 5361 228 5365 232
rect 5381 228 5385 236
rect 5391 228 5395 232
rect 5331 204 5335 208
rect 5323 199 5335 204
rect 5233 176 5237 196
rect 5223 169 5237 176
rect 5243 176 5247 196
rect 5243 169 5251 176
rect 5323 173 5327 199
rect 5351 176 5355 188
rect 5223 153 5229 169
rect 5226 141 5229 153
rect 5086 127 5095 139
rect 5014 116 5018 127
rect 5000 108 5018 116
rect 5000 104 5004 108
rect 5091 104 5095 127
rect 5099 127 5114 139
rect 5099 104 5103 127
rect 5225 64 5229 141
rect 5245 153 5251 169
rect 5245 141 5254 153
rect 5245 64 5249 141
rect 5323 80 5327 161
rect 5341 170 5355 176
rect 5341 139 5346 170
rect 5361 142 5365 188
rect 5381 184 5385 188
rect 5342 121 5347 127
rect 5391 139 5395 188
rect 5491 159 5495 216
rect 5486 147 5495 159
rect 5355 126 5385 130
rect 5342 117 5355 121
rect 5351 112 5355 117
rect 5361 112 5365 116
rect 5323 76 5335 80
rect 5331 72 5335 76
rect 5381 104 5385 126
rect 5391 127 5394 139
rect 5391 104 5395 127
rect 5331 24 5335 32
rect 5351 28 5355 32
rect 5361 24 5365 32
rect 5491 64 5495 147
rect 5605 159 5609 216
rect 5693 176 5697 196
rect 5689 169 5697 176
rect 5703 176 5707 196
rect 5703 169 5717 176
rect 5605 147 5614 159
rect 5689 153 5695 169
rect 5605 64 5609 147
rect 5686 141 5695 153
rect 5691 64 5695 141
rect 5711 153 5717 169
rect 5711 141 5714 153
rect 5711 64 5715 141
rect 85 20 89 24
rect 105 20 109 24
rect 125 20 129 24
rect 211 20 215 24
rect 231 20 235 24
rect 251 20 255 24
rect 385 20 389 24
rect 405 20 409 24
rect 425 20 429 24
rect 530 20 534 24
rect 552 20 556 24
rect 560 20 564 24
rect 656 20 660 24
rect 664 20 668 24
rect 686 20 690 24
rect 805 20 809 24
rect 825 20 829 24
rect 845 20 849 24
rect 931 20 935 24
rect 1036 20 1040 24
rect 1044 20 1048 24
rect 1066 20 1070 24
rect 1171 20 1175 24
rect 1191 20 1195 24
rect 1211 20 1215 24
rect 1311 20 1315 24
rect 1319 20 1323 24
rect 1431 20 1435 24
rect 1453 20 1457 24
rect 1475 20 1479 24
rect 1585 20 1589 24
rect 1690 20 1694 24
rect 1712 20 1716 24
rect 1720 20 1724 24
rect 1825 20 1829 24
rect 1845 20 1849 24
rect 1931 20 1935 24
rect 1951 20 1955 24
rect 1971 20 1975 24
rect 2105 20 2109 24
rect 2125 20 2129 24
rect 2145 20 2149 24
rect 2231 20 2235 24
rect 2253 20 2257 24
rect 2365 20 2369 24
rect 2385 20 2389 24
rect 2471 20 2475 24
rect 2493 20 2497 24
rect 2515 20 2519 24
rect 2625 20 2629 24
rect 2645 20 2649 24
rect 2665 20 2669 24
rect 2761 20 2765 24
rect 2783 20 2787 24
rect 2805 20 2809 24
rect 2911 20 2915 24
rect 2931 20 2935 24
rect 3045 20 3049 24
rect 3065 20 3069 24
rect 3165 20 3169 24
rect 3185 20 3189 24
rect 3205 20 3209 24
rect 3305 20 3309 24
rect 3396 20 3400 24
rect 3404 20 3408 24
rect 3426 20 3430 24
rect 3545 20 3549 24
rect 3645 20 3649 24
rect 3665 20 3669 24
rect 3763 20 3767 24
rect 3785 20 3789 24
rect 3871 20 3875 24
rect 3893 20 3897 24
rect 4005 20 4009 24
rect 4025 20 4029 24
rect 4131 20 4135 24
rect 4153 20 4157 24
rect 4175 20 4179 24
rect 4317 20 4321 24
rect 4325 20 4329 24
rect 4411 20 4415 24
rect 4431 20 4435 24
rect 4545 20 4549 24
rect 4565 20 4569 24
rect 4585 20 4589 24
rect 4710 20 4714 24
rect 4732 20 4736 24
rect 4740 20 4744 24
rect 4831 20 4835 24
rect 4851 20 4855 24
rect 4970 20 4974 24
rect 4992 20 4996 24
rect 5000 20 5004 24
rect 5091 20 5095 24
rect 5099 20 5103 24
rect 5225 20 5229 24
rect 5245 20 5249 24
rect 5331 20 5365 24
rect 5381 20 5385 24
rect 5391 20 5395 24
rect 5491 20 5495 24
rect 5605 20 5609 24
rect 5691 20 5695 24
rect 5711 20 5715 24
<< polycontact >>
rect 75 5661 87 5673
rect 134 5641 146 5653
rect 194 5641 206 5653
rect 114 5607 126 5619
rect 253 5661 265 5673
rect 214 5607 226 5619
rect 514 5681 526 5693
rect 494 5661 506 5673
rect 414 5621 426 5633
rect 394 5607 406 5619
rect 434 5607 446 5619
rect 535 5661 547 5673
rect 655 5661 667 5673
rect 714 5641 726 5653
rect 694 5607 706 5619
rect 794 5627 806 5639
rect 834 5627 846 5639
rect 954 5621 966 5633
rect 934 5607 946 5619
rect 1054 5641 1066 5653
rect 1235 5659 1247 5671
rect 1094 5641 1106 5653
rect 1254 5641 1266 5653
rect 974 5607 986 5619
rect 1235 5592 1247 5604
rect 1274 5621 1286 5633
rect 1534 5681 1546 5693
rect 1513 5661 1525 5673
rect 1414 5641 1426 5653
rect 1374 5627 1386 5639
rect 1373 5590 1385 5602
rect 1554 5661 1566 5673
rect 1834 5681 1846 5693
rect 1813 5661 1825 5673
rect 1694 5621 1706 5633
rect 1674 5607 1686 5619
rect 1714 5607 1726 5619
rect 1854 5661 1866 5673
rect 2035 5661 2047 5673
rect 1914 5621 1926 5633
rect 2094 5641 2106 5653
rect 2154 5641 2166 5653
rect 2074 5607 2086 5619
rect 2213 5661 2225 5673
rect 2174 5607 2186 5619
rect 2314 5621 2326 5633
rect 2294 5607 2306 5619
rect 2454 5627 2466 5639
rect 2334 5607 2346 5619
rect 2614 5681 2626 5693
rect 2593 5661 2605 5673
rect 2494 5627 2506 5639
rect 2754 5681 2766 5693
rect 2634 5661 2646 5673
rect 2733 5661 2745 5673
rect 2774 5661 2786 5673
rect 2834 5627 2846 5639
rect 2874 5627 2886 5639
rect 3075 5661 3087 5673
rect 2994 5621 3006 5633
rect 3134 5641 3146 5653
rect 3114 5607 3126 5619
rect 3294 5641 3306 5653
rect 3374 5641 3386 5653
rect 3534 5681 3546 5693
rect 3513 5661 3525 5673
rect 3414 5641 3426 5653
rect 3254 5627 3266 5639
rect 3253 5590 3265 5602
rect 3554 5661 3566 5673
rect 3934 5641 3946 5653
rect 3674 5621 3686 5633
rect 3774 5621 3786 5633
rect 3834 5621 3846 5633
rect 3993 5661 4005 5673
rect 3954 5607 3966 5619
rect 4181 5684 4193 5696
rect 4233 5698 4245 5710
rect 4205 5684 4217 5696
rect 4074 5621 4086 5633
rect 4153 5652 4165 5664
rect 4167 5613 4179 5625
rect 4221 5580 4233 5592
rect 4267 5698 4279 5710
rect 4253 5678 4265 5690
rect 4285 5664 4297 5676
rect 4314 5622 4326 5634
rect 4455 5661 4467 5673
rect 4294 5608 4306 5620
rect 4269 5576 4281 5588
rect 4291 5576 4303 5588
rect 4334 5621 4346 5633
rect 4514 5641 4526 5653
rect 4494 5607 4506 5619
rect 4618 5604 4630 5616
rect 4658 5604 4670 5616
rect 4698 5604 4710 5616
rect 4734 5607 4746 5619
rect 4935 5661 4947 5673
rect 4854 5621 4866 5633
rect 4994 5641 5006 5653
rect 4974 5607 4986 5619
rect 5074 5627 5086 5639
rect 5114 5627 5126 5639
rect 5174 5627 5186 5639
rect 5294 5641 5306 5653
rect 5214 5627 5226 5639
rect 5353 5661 5365 5673
rect 5314 5607 5326 5619
rect 5434 5621 5446 5633
rect 5534 5627 5546 5639
rect 5574 5627 5586 5639
rect 5654 5621 5666 5633
rect 114 5441 126 5453
rect 75 5387 87 5399
rect 134 5407 146 5419
rect 253 5387 265 5399
rect 294 5387 306 5399
rect 393 5387 405 5399
rect 274 5367 286 5379
rect 434 5387 446 5399
rect 533 5387 545 5399
rect 414 5367 426 5379
rect 574 5387 586 5399
rect 654 5387 666 5399
rect 554 5367 566 5379
rect 814 5441 826 5453
rect 794 5407 806 5419
rect 695 5387 707 5399
rect 674 5367 686 5379
rect 853 5387 865 5399
rect 934 5387 946 5399
rect 1114 5441 1126 5453
rect 975 5387 987 5399
rect 954 5367 966 5379
rect 1154 5441 1166 5453
rect 1134 5427 1146 5439
rect 1214 5387 1226 5399
rect 1374 5407 1386 5419
rect 1255 5387 1267 5399
rect 1234 5367 1246 5379
rect 1414 5407 1426 5419
rect 1533 5387 1545 5399
rect 1654 5441 1666 5453
rect 1634 5407 1646 5419
rect 1574 5387 1586 5399
rect 1554 5367 1566 5379
rect 1693 5387 1705 5399
rect 1813 5387 1825 5399
rect 1854 5387 1866 5399
rect 1953 5387 1965 5399
rect 1834 5367 1846 5379
rect 2054 5421 2066 5433
rect 1994 5387 2006 5399
rect 1974 5367 1986 5379
rect 2333 5458 2345 5470
rect 2094 5421 2106 5433
rect 2234 5427 2246 5439
rect 2334 5421 2346 5433
rect 2454 5441 2466 5453
rect 2374 5407 2386 5419
rect 2434 5407 2446 5419
rect 2493 5387 2505 5399
rect 2633 5387 2645 5399
rect 2674 5387 2686 5399
rect 2773 5387 2785 5399
rect 2654 5367 2666 5379
rect 2894 5441 2906 5453
rect 2874 5407 2886 5419
rect 2814 5387 2826 5399
rect 2794 5367 2806 5379
rect 3014 5427 3026 5439
rect 2933 5387 2945 5399
rect 3114 5421 3126 5433
rect 3154 5421 3166 5433
rect 3254 5387 3266 5399
rect 3394 5421 3406 5433
rect 3295 5387 3307 5399
rect 3274 5367 3286 5379
rect 3434 5421 3446 5433
rect 3514 5427 3526 5439
rect 3553 5456 3565 5468
rect 3534 5407 3546 5419
rect 3553 5389 3565 5401
rect 3693 5387 3705 5399
rect 3834 5441 3846 5453
rect 3734 5387 3746 5399
rect 3714 5367 3726 5379
rect 3874 5441 3886 5453
rect 3854 5427 3866 5439
rect 3934 5421 3946 5433
rect 3974 5421 3986 5433
rect 4114 5441 4126 5453
rect 4075 5387 4087 5399
rect 4214 5421 4226 5433
rect 4134 5407 4146 5419
rect 4254 5421 4266 5433
rect 4353 5387 4365 5399
rect 4474 5441 4486 5453
rect 4514 5441 4526 5453
rect 4494 5427 4506 5439
rect 4394 5387 4406 5399
rect 4374 5367 4386 5379
rect 4614 5427 4626 5439
rect 4734 5441 4746 5453
rect 4714 5407 4726 5419
rect 4847 5435 4859 5447
rect 4773 5387 4785 5399
rect 4833 5396 4845 5408
rect 4901 5468 4913 5480
rect 4861 5364 4873 5376
rect 4885 5364 4897 5376
rect 4949 5472 4961 5484
rect 4971 5472 4983 5484
rect 4933 5370 4945 5382
rect 4913 5350 4925 5362
rect 4974 5440 4986 5452
rect 4994 5426 5006 5438
rect 5014 5427 5026 5439
rect 5094 5427 5106 5439
rect 4965 5384 4977 5396
rect 4947 5350 4959 5362
rect 5187 5435 5199 5447
rect 5173 5396 5185 5408
rect 5241 5468 5253 5480
rect 5201 5364 5213 5376
rect 5225 5364 5237 5376
rect 5289 5472 5301 5484
rect 5311 5472 5323 5484
rect 5273 5370 5285 5382
rect 5253 5350 5265 5362
rect 5314 5440 5326 5452
rect 5334 5426 5346 5438
rect 5354 5427 5366 5439
rect 5305 5384 5317 5396
rect 5287 5350 5299 5362
rect 5454 5441 5466 5453
rect 5434 5407 5446 5419
rect 5594 5421 5606 5433
rect 5493 5387 5505 5399
rect 5634 5421 5646 5433
rect 5714 5421 5726 5433
rect 5754 5421 5766 5433
rect 114 5201 126 5213
rect 93 5181 105 5193
rect 134 5181 146 5193
rect 214 5141 226 5153
rect 194 5127 206 5139
rect 494 5201 506 5213
rect 473 5181 485 5193
rect 334 5141 346 5153
rect 234 5127 246 5139
rect 514 5181 526 5193
rect 594 5141 606 5153
rect 574 5127 586 5139
rect 614 5127 626 5139
rect 874 5201 886 5213
rect 854 5181 866 5193
rect 774 5141 786 5153
rect 754 5127 766 5139
rect 794 5127 806 5139
rect 895 5181 907 5193
rect 1054 5201 1066 5213
rect 1033 5181 1045 5193
rect 1074 5181 1086 5193
rect 1294 5201 1306 5213
rect 1273 5181 1285 5193
rect 1134 5141 1146 5153
rect 1314 5181 1326 5193
rect 1415 5181 1427 5193
rect 1474 5161 1486 5173
rect 1454 5127 1466 5139
rect 1655 5181 1667 5193
rect 1574 5141 1586 5153
rect 1714 5161 1726 5173
rect 1874 5161 1886 5173
rect 1694 5127 1706 5139
rect 1894 5127 1906 5139
rect 1934 5161 1946 5173
rect 2034 5161 2046 5173
rect 2113 5161 2125 5173
rect 2055 5127 2067 5139
rect 2093 5127 2105 5139
rect 2174 5147 2186 5159
rect 2354 5201 2366 5213
rect 2333 5181 2345 5193
rect 2214 5147 2226 5159
rect 2374 5181 2386 5193
rect 2494 5141 2506 5153
rect 2474 5127 2486 5139
rect 2695 5181 2707 5193
rect 2614 5141 2626 5153
rect 2514 5127 2526 5139
rect 2855 5181 2867 5193
rect 2754 5161 2766 5173
rect 2734 5127 2746 5139
rect 2914 5161 2926 5173
rect 2894 5127 2906 5139
rect 3054 5161 3066 5173
rect 3114 5161 3126 5173
rect 3154 5161 3166 5173
rect 3014 5147 3026 5159
rect 3013 5110 3025 5122
rect 3374 5161 3386 5173
rect 3515 5181 3527 5193
rect 3414 5161 3426 5173
rect 3294 5141 3306 5153
rect 3574 5161 3586 5173
rect 3554 5127 3566 5139
rect 3634 5147 3646 5159
rect 3674 5147 3686 5159
rect 3774 5147 3786 5159
rect 3814 5147 3826 5159
rect 3914 5147 3926 5159
rect 4034 5201 4046 5213
rect 4014 5181 4026 5193
rect 3954 5147 3966 5159
rect 4055 5181 4067 5193
rect 4175 5181 4187 5193
rect 4234 5161 4246 5173
rect 4314 5161 4326 5173
rect 4214 5127 4226 5139
rect 4373 5181 4385 5193
rect 4334 5127 4346 5139
rect 4614 5201 4626 5213
rect 4593 5181 4605 5193
rect 4454 5141 4466 5153
rect 4961 5204 4973 5216
rect 5013 5218 5025 5230
rect 4985 5204 4997 5216
rect 4634 5181 4646 5193
rect 4714 5141 4726 5153
rect 4694 5127 4706 5139
rect 4834 5161 4846 5173
rect 4874 5161 4886 5173
rect 4933 5172 4945 5184
rect 4734 5127 4746 5139
rect 4947 5133 4959 5145
rect 5001 5100 5013 5112
rect 5047 5218 5059 5230
rect 5033 5198 5045 5210
rect 5065 5184 5077 5196
rect 5094 5142 5106 5154
rect 5194 5161 5206 5173
rect 5074 5128 5086 5140
rect 5049 5096 5061 5108
rect 5071 5096 5083 5108
rect 5114 5141 5126 5153
rect 5253 5181 5265 5193
rect 5214 5127 5226 5139
rect 5434 5161 5446 5173
rect 5334 5141 5346 5153
rect 5493 5181 5505 5193
rect 5454 5127 5466 5139
rect 5594 5147 5606 5159
rect 5634 5147 5646 5159
rect 5694 5147 5706 5159
rect 5734 5147 5746 5159
rect 114 4961 126 4973
rect 75 4907 87 4919
rect 134 4927 146 4939
rect 233 4907 245 4919
rect 274 4907 286 4919
rect 334 4907 346 4919
rect 254 4887 266 4899
rect 494 4961 506 4973
rect 474 4927 486 4939
rect 375 4907 387 4919
rect 354 4887 366 4899
rect 634 4941 646 4953
rect 533 4907 545 4919
rect 674 4941 686 4953
rect 794 4961 806 4973
rect 755 4907 767 4919
rect 814 4927 826 4939
rect 934 4961 946 4973
rect 895 4907 907 4919
rect 1054 4961 1066 4973
rect 954 4927 966 4939
rect 1094 4961 1106 4973
rect 1074 4947 1086 4959
rect 1214 4961 1226 4973
rect 1175 4907 1187 4919
rect 1334 4947 1346 4959
rect 1234 4927 1246 4939
rect 1414 4941 1426 4953
rect 1454 4941 1466 4953
rect 1573 4907 1585 4919
rect 1734 4961 1746 4973
rect 1614 4907 1626 4919
rect 1695 4907 1707 4919
rect 1594 4887 1606 4899
rect 1814 4961 1826 4973
rect 1754 4927 1766 4939
rect 1854 4961 1866 4973
rect 1834 4947 1846 4959
rect 1954 4941 1966 4953
rect 2114 4961 2126 4973
rect 1994 4941 2006 4953
rect 2154 4961 2166 4973
rect 2134 4947 2146 4959
rect 2274 4947 2286 4959
rect 2394 4961 2406 4973
rect 2355 4907 2367 4919
rect 2414 4927 2426 4939
rect 2513 4907 2525 4919
rect 2654 4947 2666 4959
rect 2554 4907 2566 4919
rect 2534 4887 2546 4899
rect 2754 4941 2766 4953
rect 2794 4941 2806 4953
rect 2854 4947 2866 4959
rect 2954 4907 2966 4919
rect 3154 4961 3166 4973
rect 2995 4907 3007 4919
rect 3115 4907 3127 4919
rect 2974 4887 2986 4899
rect 3174 4927 3186 4939
rect 3294 4961 3306 4973
rect 3255 4907 3267 4919
rect 3414 4961 3426 4973
rect 3314 4927 3326 4939
rect 3454 4961 3466 4973
rect 3434 4947 3446 4959
rect 3514 4947 3526 4959
rect 3553 4976 3565 4988
rect 3534 4927 3546 4939
rect 3674 4927 3686 4939
rect 3553 4909 3565 4921
rect 3714 4927 3726 4939
rect 3813 4907 3825 4919
rect 4333 4978 4345 4990
rect 3954 4947 3966 4959
rect 3854 4907 3866 4919
rect 3834 4887 3846 4899
rect 4014 4907 4026 4919
rect 4055 4907 4067 4919
rect 4154 4907 4166 4919
rect 4034 4887 4046 4899
rect 4195 4907 4207 4919
rect 4174 4887 4186 4899
rect 4334 4941 4346 4953
rect 4454 4947 4466 4959
rect 4374 4927 4386 4939
rect 4493 4976 4505 4988
rect 4474 4927 4486 4939
rect 4594 4927 4606 4939
rect 4493 4909 4505 4921
rect 4634 4927 4646 4939
rect 4774 4961 4786 4973
rect 4735 4907 4747 4919
rect 4794 4927 4806 4939
rect 4847 4955 4859 4967
rect 4833 4916 4845 4928
rect 4901 4988 4913 5000
rect 4861 4884 4873 4896
rect 4885 4884 4897 4896
rect 4949 4992 4961 5004
rect 4971 4992 4983 5004
rect 4933 4890 4945 4902
rect 4913 4870 4925 4882
rect 4974 4960 4986 4972
rect 4994 4946 5006 4958
rect 5014 4947 5026 4959
rect 4965 4904 4977 4916
rect 4947 4870 4959 4882
rect 5114 4961 5126 4973
rect 5094 4927 5106 4939
rect 5227 4955 5239 4967
rect 5153 4907 5165 4919
rect 5213 4916 5225 4928
rect 5281 4988 5293 5000
rect 5241 4884 5253 4896
rect 5265 4884 5277 4896
rect 5329 4992 5341 5004
rect 5351 4992 5363 5004
rect 5313 4890 5325 4902
rect 5293 4870 5305 4882
rect 5354 4960 5366 4972
rect 5374 4946 5386 4958
rect 5394 4947 5406 4959
rect 5345 4904 5357 4916
rect 5327 4870 5339 4882
rect 5494 4941 5506 4953
rect 5534 4941 5546 4953
rect 5594 4941 5606 4953
rect 5634 4941 5646 4953
rect 5734 4941 5746 4953
rect 5774 4941 5786 4953
rect 254 4721 266 4733
rect 233 4701 245 4713
rect 114 4661 126 4673
rect 94 4647 106 4659
rect 134 4647 146 4659
rect 274 4701 286 4713
rect 354 4661 366 4673
rect 334 4647 346 4659
rect 474 4667 486 4679
rect 374 4647 386 4659
rect 654 4721 666 4733
rect 633 4701 645 4713
rect 514 4667 526 4679
rect 814 4721 826 4733
rect 674 4701 686 4713
rect 793 4701 805 4713
rect 834 4701 846 4713
rect 894 4661 906 4673
rect 994 4661 1006 4673
rect 1215 4701 1227 4713
rect 1134 4661 1146 4673
rect 1274 4681 1286 4693
rect 1334 4681 1346 4693
rect 1254 4647 1266 4659
rect 1393 4701 1405 4713
rect 1354 4647 1366 4659
rect 1594 4721 1606 4733
rect 1574 4701 1586 4713
rect 1474 4661 1486 4673
rect 1615 4701 1627 4713
rect 1735 4701 1747 4713
rect 1794 4681 1806 4693
rect 1774 4647 1786 4659
rect 1874 4667 1886 4679
rect 1974 4681 1986 4693
rect 1914 4667 1926 4679
rect 2174 4721 2186 4733
rect 2033 4701 2045 4713
rect 2153 4701 2165 4713
rect 1994 4647 2006 4659
rect 2194 4701 2206 4713
rect 2285 4698 2297 4710
rect 2314 4681 2326 4693
rect 2285 4630 2297 4642
rect 2374 4667 2386 4679
rect 2414 4667 2426 4679
rect 2494 4667 2506 4679
rect 2645 4698 2657 4710
rect 2754 4721 2766 4733
rect 2734 4701 2746 4713
rect 2674 4681 2686 4693
rect 2534 4667 2546 4679
rect 2645 4630 2657 4642
rect 2775 4701 2787 4713
rect 2894 4681 2906 4693
rect 2934 4681 2946 4693
rect 3014 4681 3026 4693
rect 3093 4681 3105 4693
rect 3034 4647 3046 4659
rect 3070 4647 3082 4659
rect 3194 4667 3206 4679
rect 3354 4721 3366 4733
rect 3333 4701 3345 4713
rect 3234 4667 3246 4679
rect 3374 4701 3386 4713
rect 3634 4721 3646 4733
rect 3613 4701 3625 4713
rect 3494 4661 3506 4673
rect 3474 4647 3486 4659
rect 3514 4647 3526 4659
rect 3654 4701 3666 4713
rect 3874 4721 3886 4733
rect 3854 4701 3866 4713
rect 3774 4661 3786 4673
rect 3754 4647 3766 4659
rect 3794 4647 3806 4659
rect 4014 4721 4026 4733
rect 3895 4701 3907 4713
rect 3994 4701 4006 4713
rect 4035 4701 4047 4713
rect 4134 4661 4146 4673
rect 4454 4721 4466 4733
rect 4433 4701 4445 4713
rect 4314 4681 4326 4693
rect 4274 4667 4286 4679
rect 4273 4630 4285 4642
rect 4554 4721 4566 4733
rect 4474 4701 4486 4713
rect 4534 4701 4546 4713
rect 4575 4701 4587 4713
rect 4781 4724 4793 4736
rect 4833 4738 4845 4750
rect 4805 4724 4817 4736
rect 4674 4661 4686 4673
rect 4753 4692 4765 4704
rect 4767 4653 4779 4665
rect 4821 4620 4833 4632
rect 4867 4738 4879 4750
rect 4853 4718 4865 4730
rect 4885 4704 4897 4716
rect 4914 4662 4926 4674
rect 5014 4681 5026 4693
rect 4894 4648 4906 4660
rect 4869 4616 4881 4628
rect 4891 4616 4903 4628
rect 4934 4661 4946 4673
rect 5073 4701 5085 4713
rect 5034 4647 5046 4659
rect 5154 4667 5166 4679
rect 5194 4667 5206 4679
rect 5274 4667 5286 4679
rect 5314 4667 5326 4679
rect 5414 4667 5426 4679
rect 5454 4667 5466 4679
rect 5534 4667 5546 4679
rect 5714 4721 5726 4733
rect 5693 4701 5705 4713
rect 5574 4667 5586 4679
rect 5734 4701 5746 4713
rect 114 4481 126 4493
rect 75 4427 87 4439
rect 134 4447 146 4459
rect 233 4427 245 4439
rect 334 4481 346 4493
rect 374 4481 386 4493
rect 354 4467 366 4479
rect 274 4427 286 4439
rect 254 4407 266 4419
rect 554 4481 566 4493
rect 515 4427 527 4439
rect 574 4447 586 4459
rect 694 4481 706 4493
rect 655 4427 667 4439
rect 874 4481 886 4493
rect 774 4467 786 4479
rect 714 4447 726 4459
rect 914 4481 926 4493
rect 894 4467 906 4479
rect 1054 4467 1066 4479
rect 1153 4427 1165 4439
rect 1294 4481 1306 4493
rect 1194 4427 1206 4439
rect 1174 4407 1186 4419
rect 1334 4481 1346 4493
rect 1314 4467 1326 4479
rect 1434 4467 1446 4479
rect 1514 4481 1526 4493
rect 1494 4447 1506 4459
rect 1654 4461 1666 4473
rect 1553 4427 1565 4439
rect 1694 4461 1706 4473
rect 1793 4427 1805 4439
rect 1914 4447 1926 4459
rect 1834 4427 1846 4439
rect 1814 4407 1826 4419
rect 1954 4447 1966 4459
rect 2053 4427 2065 4439
rect 2094 4427 2106 4439
rect 2213 4427 2225 4439
rect 2074 4407 2086 4419
rect 2334 4461 2346 4473
rect 2254 4427 2266 4439
rect 2234 4407 2246 4419
rect 2374 4461 2386 4473
rect 2473 4427 2485 4439
rect 2514 4427 2526 4439
rect 2574 4427 2586 4439
rect 2494 4407 2506 4419
rect 2754 4467 2766 4479
rect 2615 4427 2627 4439
rect 2594 4407 2606 4419
rect 2834 4447 2846 4459
rect 2874 4447 2886 4459
rect 2973 4427 2985 4439
rect 3014 4427 3026 4439
rect 3113 4427 3125 4439
rect 2994 4407 3006 4419
rect 3214 4467 3226 4479
rect 3154 4427 3166 4439
rect 3134 4407 3146 4419
rect 3334 4481 3346 4493
rect 3314 4447 3326 4459
rect 3493 4498 3505 4510
rect 3373 4427 3385 4439
rect 3494 4461 3506 4473
rect 3775 4496 3787 4508
rect 3614 4461 3626 4473
rect 3534 4447 3546 4459
rect 3654 4461 3666 4473
rect 4025 4498 4037 4510
rect 3814 4467 3826 4479
rect 3794 4447 3806 4459
rect 3775 4429 3787 4441
rect 3874 4461 3886 4473
rect 3914 4461 3926 4473
rect 4155 4498 4167 4510
rect 4154 4461 4166 4473
rect 4054 4447 4066 4459
rect 4114 4447 4126 4459
rect 4025 4430 4037 4442
rect 4274 4461 4286 4473
rect 4314 4461 4326 4473
rect 4434 4481 4446 4493
rect 4395 4427 4407 4439
rect 4514 4461 4526 4473
rect 4454 4447 4466 4459
rect 4554 4461 4566 4473
rect 4654 4461 4666 4473
rect 4694 4461 4706 4473
rect 4754 4467 4766 4479
rect 4854 4461 4866 4473
rect 4894 4461 4906 4473
rect 4994 4481 5006 4493
rect 4974 4447 4986 4459
rect 5107 4475 5119 4487
rect 5033 4427 5045 4439
rect 5093 4436 5105 4448
rect 5161 4508 5173 4520
rect 5121 4404 5133 4416
rect 5145 4404 5157 4416
rect 5209 4512 5221 4524
rect 5231 4512 5243 4524
rect 5193 4410 5205 4422
rect 5173 4390 5185 4402
rect 5234 4480 5246 4492
rect 5254 4466 5266 4478
rect 5274 4467 5286 4479
rect 5225 4424 5237 4436
rect 5207 4390 5219 4402
rect 5374 4481 5386 4493
rect 5354 4447 5366 4459
rect 5494 4467 5506 4479
rect 5413 4427 5425 4439
rect 5533 4496 5545 4508
rect 5514 4447 5526 4459
rect 5533 4429 5545 4441
rect 5694 4481 5706 4493
rect 5655 4427 5667 4439
rect 5714 4447 5726 4459
rect 95 4221 107 4233
rect 235 4221 247 4233
rect 154 4201 166 4213
rect 134 4167 146 4179
rect 434 4241 446 4253
rect 413 4221 425 4233
rect 294 4201 306 4213
rect 274 4167 286 4179
rect 574 4241 586 4253
rect 454 4221 466 4233
rect 553 4221 565 4233
rect 594 4221 606 4233
rect 695 4219 707 4231
rect 714 4201 726 4213
rect 695 4152 707 4164
rect 815 4221 827 4233
rect 734 4181 746 4193
rect 874 4201 886 4213
rect 854 4167 866 4179
rect 934 4181 946 4193
rect 1254 4241 1266 4253
rect 1233 4221 1245 4233
rect 1094 4181 1106 4193
rect 1074 4167 1086 4179
rect 1114 4167 1126 4179
rect 1274 4221 1286 4233
rect 1354 4187 1366 4199
rect 1394 4187 1406 4199
rect 1474 4187 1486 4199
rect 1594 4201 1606 4213
rect 1754 4241 1766 4253
rect 1733 4221 1745 4233
rect 1634 4201 1646 4213
rect 1514 4187 1526 4199
rect 1894 4241 1906 4253
rect 1774 4221 1786 4233
rect 1873 4221 1885 4233
rect 1994 4241 2006 4253
rect 1914 4221 1926 4233
rect 1974 4221 1986 4233
rect 2134 4241 2146 4253
rect 2015 4221 2027 4233
rect 2114 4221 2126 4233
rect 2155 4221 2167 4233
rect 2274 4201 2286 4213
rect 2415 4221 2427 4233
rect 2314 4201 2326 4213
rect 2614 4241 2626 4253
rect 2593 4221 2605 4233
rect 2474 4201 2486 4213
rect 2454 4167 2466 4179
rect 2634 4221 2646 4233
rect 2834 4241 2846 4253
rect 2814 4221 2826 4233
rect 2694 4181 2706 4193
rect 2855 4221 2867 4233
rect 2954 4187 2966 4199
rect 2994 4187 3006 4199
rect 3094 4181 3106 4193
rect 3074 4167 3086 4179
rect 3234 4181 3246 4193
rect 3114 4167 3126 4179
rect 3214 4167 3226 4179
rect 3354 4201 3366 4213
rect 3254 4167 3266 4179
rect 3413 4221 3425 4233
rect 3374 4167 3386 4179
rect 3634 4241 3646 4253
rect 3614 4221 3626 4233
rect 3514 4181 3526 4193
rect 3774 4241 3786 4253
rect 3655 4221 3667 4233
rect 3754 4221 3766 4233
rect 3795 4221 3807 4233
rect 3914 4187 3926 4199
rect 3954 4187 3966 4199
rect 4054 4187 4066 4199
rect 4094 4187 4106 4199
rect 4174 4187 4186 4199
rect 4295 4221 4307 4233
rect 4214 4187 4226 4199
rect 4354 4201 4366 4213
rect 4334 4167 4346 4179
rect 4453 4219 4465 4231
rect 4575 4221 4587 4233
rect 4434 4201 4446 4213
rect 4414 4181 4426 4193
rect 4453 4152 4465 4164
rect 4634 4201 4646 4213
rect 4714 4201 4726 4213
rect 4614 4167 4626 4179
rect 4773 4221 4785 4233
rect 4734 4167 4746 4179
rect 4854 4201 4866 4213
rect 4894 4201 4906 4213
rect 4974 4181 4986 4193
rect 5114 4181 5126 4193
rect 5094 4167 5106 4179
rect 5234 4201 5246 4213
rect 5134 4167 5146 4179
rect 5293 4221 5305 4233
rect 5254 4167 5266 4179
rect 5474 4201 5486 4213
rect 5374 4181 5386 4193
rect 5533 4221 5545 4233
rect 5494 4167 5506 4179
rect 5661 4258 5673 4270
rect 5643 4224 5655 4236
rect 5594 4181 5606 4193
rect 5614 4182 5626 4194
rect 5634 4168 5646 4180
rect 5695 4258 5707 4270
rect 5675 4238 5687 4250
rect 5637 4136 5649 4148
rect 5659 4136 5671 4148
rect 5723 4244 5735 4256
rect 5747 4244 5759 4256
rect 5707 4140 5719 4152
rect 5775 4212 5787 4224
rect 5761 4173 5773 4185
rect 94 3987 106 3999
rect 194 4001 206 4013
rect 174 3967 186 3979
rect 434 4001 446 4013
rect 354 3987 366 3999
rect 233 3947 245 3959
rect 474 4001 486 4013
rect 454 3987 466 3999
rect 754 3987 766 3999
rect 594 3967 606 3979
rect 634 3967 646 3979
rect 834 4001 846 4013
rect 814 3967 826 3979
rect 954 3987 966 3999
rect 873 3947 885 3959
rect 1054 3947 1066 3959
rect 1215 4001 1227 4013
rect 1253 4001 1265 4013
rect 1195 3967 1207 3979
rect 1095 3947 1107 3959
rect 1074 3927 1086 3939
rect 1374 3981 1386 3993
rect 1274 3967 1286 3979
rect 1414 3981 1426 3993
rect 1534 3987 1546 3999
rect 1754 3987 1766 3999
rect 1614 3967 1626 3979
rect 1654 3967 1666 3979
rect 1814 3947 1826 3959
rect 2014 4001 2026 4013
rect 1855 3947 1867 3959
rect 1975 3947 1987 3959
rect 1834 3927 1846 3939
rect 2034 3967 2046 3979
rect 2153 3947 2165 3959
rect 2194 3947 2206 3959
rect 2254 3947 2266 3959
rect 2174 3927 2186 3939
rect 2454 4001 2466 4013
rect 2295 3947 2307 3959
rect 2415 3947 2427 3959
rect 2274 3927 2286 3939
rect 2554 3981 2566 3993
rect 2474 3967 2486 3979
rect 2594 3981 2606 3993
rect 2654 3981 2666 3993
rect 2694 3981 2706 3993
rect 2774 3947 2786 3959
rect 2815 3947 2827 3959
rect 2914 3947 2926 3959
rect 2794 3927 2806 3939
rect 3094 3987 3106 3999
rect 2955 3947 2967 3959
rect 2934 3927 2946 3939
rect 3193 3947 3205 3959
rect 3334 3987 3346 3999
rect 3234 3947 3246 3959
rect 3214 3927 3226 3939
rect 3454 4001 3466 4013
rect 3415 3947 3427 3959
rect 3695 4016 3707 4028
rect 3534 3981 3546 3993
rect 3474 3967 3486 3979
rect 3574 3981 3586 3993
rect 3734 3987 3746 3999
rect 3714 3967 3726 3979
rect 3695 3949 3707 3961
rect 3814 3981 3826 3993
rect 3854 3981 3866 3993
rect 3994 4001 4006 4013
rect 3955 3947 3967 3959
rect 4114 4001 4126 4013
rect 4014 3967 4026 3979
rect 4154 4001 4166 4013
rect 4134 3987 4146 3999
rect 4214 3981 4226 3993
rect 4254 3981 4266 3993
rect 4354 4001 4366 4013
rect 4334 3967 4346 3979
rect 4494 4001 4506 4013
rect 4474 3967 4486 3979
rect 4393 3947 4405 3959
rect 4614 3987 4626 3999
rect 4533 3947 4545 3959
rect 4653 4016 4665 4028
rect 4774 3981 4786 3993
rect 4634 3967 4646 3979
rect 4653 3949 4665 3961
rect 4814 3981 4826 3993
rect 4874 3947 4886 3959
rect 5014 3987 5026 3999
rect 4915 3947 4927 3959
rect 4894 3927 4906 3939
rect 5154 3987 5166 3999
rect 5207 3995 5219 4007
rect 5193 3956 5205 3968
rect 5261 4028 5273 4040
rect 5221 3924 5233 3936
rect 5245 3924 5257 3936
rect 5309 4032 5321 4044
rect 5331 4032 5343 4044
rect 5293 3930 5305 3942
rect 5273 3910 5285 3922
rect 5334 4000 5346 4012
rect 5354 3986 5366 3998
rect 5374 3987 5386 3999
rect 5325 3944 5337 3956
rect 5307 3910 5319 3922
rect 5447 3995 5459 4007
rect 5433 3956 5445 3968
rect 5501 4028 5513 4040
rect 5461 3924 5473 3936
rect 5485 3924 5497 3936
rect 5549 4032 5561 4044
rect 5571 4032 5583 4044
rect 5533 3930 5545 3942
rect 5513 3910 5525 3922
rect 5574 4000 5586 4012
rect 5594 3986 5606 3998
rect 5614 3987 5626 3999
rect 5565 3944 5577 3956
rect 5547 3910 5559 3922
rect 5714 4001 5726 4013
rect 5694 3967 5706 3979
rect 5753 3947 5765 3959
rect 74 3707 86 3719
rect 234 3761 246 3773
rect 213 3741 225 3753
rect 114 3707 126 3719
rect 254 3741 266 3753
rect 394 3721 406 3733
rect 414 3687 426 3699
rect 555 3741 567 3753
rect 454 3721 466 3733
rect 614 3721 626 3733
rect 594 3687 606 3699
rect 694 3707 706 3719
rect 794 3721 806 3733
rect 734 3707 746 3719
rect 853 3741 865 3753
rect 814 3687 826 3699
rect 974 3721 986 3733
rect 1053 3721 1065 3733
rect 995 3687 1007 3699
rect 1033 3687 1045 3699
rect 1114 3707 1126 3719
rect 1254 3761 1266 3773
rect 1234 3741 1246 3753
rect 1154 3707 1166 3719
rect 1275 3741 1287 3753
rect 1394 3701 1406 3713
rect 1374 3687 1386 3699
rect 1514 3721 1526 3733
rect 1414 3687 1426 3699
rect 1573 3741 1585 3753
rect 1534 3687 1546 3699
rect 1654 3701 1666 3713
rect 1774 3707 1786 3719
rect 1814 3707 1826 3719
rect 1874 3707 1886 3719
rect 1914 3707 1926 3719
rect 2033 3739 2045 3751
rect 2014 3721 2026 3733
rect 1994 3701 2006 3713
rect 2134 3707 2146 3719
rect 2274 3761 2286 3773
rect 2254 3741 2266 3753
rect 2174 3707 2186 3719
rect 2033 3672 2045 3684
rect 2295 3741 2307 3753
rect 2415 3741 2427 3753
rect 2474 3721 2486 3733
rect 2454 3687 2466 3699
rect 2534 3707 2546 3719
rect 2654 3721 2666 3733
rect 2574 3707 2586 3719
rect 2713 3741 2725 3753
rect 2674 3687 2686 3699
rect 2915 3741 2927 3753
rect 2834 3701 2846 3713
rect 2974 3721 2986 3733
rect 2954 3687 2966 3699
rect 3034 3707 3046 3719
rect 3074 3707 3086 3719
rect 3194 3707 3206 3719
rect 3234 3707 3246 3719
rect 3414 3761 3426 3773
rect 3394 3741 3406 3753
rect 3334 3701 3346 3713
rect 3435 3741 3447 3753
rect 3654 3721 3666 3733
rect 3694 3721 3706 3733
rect 3534 3701 3546 3713
rect 3774 3707 3786 3719
rect 3814 3707 3826 3719
rect 3894 3701 3906 3713
rect 4101 3764 4113 3776
rect 4153 3778 4165 3790
rect 4125 3764 4137 3776
rect 4073 3732 4085 3744
rect 4034 3701 4046 3713
rect 4087 3693 4099 3705
rect 4141 3660 4153 3672
rect 4187 3778 4199 3790
rect 4173 3758 4185 3770
rect 4205 3744 4217 3756
rect 4234 3702 4246 3714
rect 4355 3721 4367 3733
rect 4214 3688 4226 3700
rect 4189 3656 4201 3668
rect 4211 3656 4223 3668
rect 4254 3701 4266 3713
rect 4434 3721 4446 3733
rect 4378 3687 4390 3699
rect 4414 3687 4426 3699
rect 4494 3707 4506 3719
rect 4614 3721 4626 3733
rect 4654 3721 4666 3733
rect 4734 3721 4746 3733
rect 4534 3707 4546 3719
rect 4793 3741 4805 3753
rect 4754 3687 4766 3699
rect 5014 3707 5026 3719
rect 4874 3687 4886 3699
rect 5054 3707 5066 3719
rect 5461 3764 5473 3776
rect 5513 3778 5525 3790
rect 5485 3764 5497 3776
rect 5114 3701 5126 3713
rect 5258 3684 5270 3696
rect 5298 3684 5310 3696
rect 5338 3684 5350 3696
rect 5374 3687 5386 3699
rect 5433 3732 5445 3744
rect 5447 3693 5459 3705
rect 5501 3660 5513 3672
rect 5547 3778 5559 3790
rect 5533 3758 5545 3770
rect 5565 3744 5577 3756
rect 5594 3702 5606 3714
rect 5574 3688 5586 3700
rect 5549 3656 5561 3668
rect 5571 3656 5583 3668
rect 5614 3701 5626 3713
rect 5714 3707 5726 3719
rect 5754 3707 5766 3719
rect 114 3521 126 3533
rect 75 3467 87 3479
rect 194 3521 206 3533
rect 134 3487 146 3499
rect 234 3521 246 3533
rect 214 3507 226 3519
rect 334 3507 346 3519
rect 454 3521 466 3533
rect 434 3487 446 3499
rect 493 3467 505 3479
rect 574 3467 586 3479
rect 754 3501 766 3513
rect 615 3467 627 3479
rect 594 3447 606 3459
rect 794 3501 806 3513
rect 874 3501 886 3513
rect 914 3501 926 3513
rect 994 3521 1006 3533
rect 974 3487 986 3499
rect 1033 3467 1045 3479
rect 1153 3467 1165 3479
rect 1254 3501 1266 3513
rect 1194 3467 1206 3479
rect 1174 3447 1186 3459
rect 1294 3501 1306 3513
rect 1413 3467 1425 3479
rect 1534 3521 1546 3533
rect 1514 3487 1526 3499
rect 1454 3467 1466 3479
rect 1434 3447 1446 3459
rect 1694 3521 1706 3533
rect 1573 3467 1585 3479
rect 1734 3521 1746 3533
rect 1714 3507 1726 3519
rect 1833 3467 1845 3479
rect 1934 3521 1946 3533
rect 1974 3521 1986 3533
rect 1954 3507 1966 3519
rect 1874 3467 1886 3479
rect 1854 3447 1866 3459
rect 2134 3521 2146 3533
rect 2095 3467 2107 3479
rect 2254 3521 2266 3533
rect 2154 3487 2166 3499
rect 2234 3487 2246 3499
rect 2414 3521 2426 3533
rect 2293 3467 2305 3479
rect 2553 3538 2565 3550
rect 2454 3521 2466 3533
rect 2434 3507 2446 3519
rect 2554 3501 2566 3513
rect 2654 3501 2666 3513
rect 2594 3487 2606 3499
rect 2694 3501 2706 3513
rect 2834 3521 2846 3533
rect 2795 3467 2807 3479
rect 2965 3538 2977 3550
rect 3074 3501 3086 3513
rect 2854 3487 2866 3499
rect 2994 3487 3006 3499
rect 2965 3470 2977 3482
rect 3114 3501 3126 3513
rect 3174 3467 3186 3479
rect 3215 3467 3227 3479
rect 3194 3447 3206 3459
rect 3353 3467 3365 3479
rect 3514 3521 3526 3533
rect 3394 3467 3406 3479
rect 3475 3467 3487 3479
rect 3374 3447 3386 3459
rect 3534 3487 3546 3499
rect 3654 3521 3666 3533
rect 3615 3467 3627 3479
rect 3773 3538 3785 3550
rect 3674 3487 3686 3499
rect 3774 3501 3786 3513
rect 3814 3487 3826 3499
rect 3874 3487 3886 3499
rect 3914 3487 3926 3499
rect 4074 3521 4086 3533
rect 4035 3467 4047 3479
rect 4154 3507 4166 3519
rect 4094 3487 4106 3499
rect 4274 3521 4286 3533
rect 4254 3487 4266 3499
rect 4414 3501 4426 3513
rect 4313 3467 4325 3479
rect 4454 3501 4466 3513
rect 4514 3501 4526 3513
rect 4554 3501 4566 3513
rect 4627 3515 4639 3527
rect 4613 3476 4625 3488
rect 4681 3548 4693 3560
rect 4641 3444 4653 3456
rect 4665 3444 4677 3456
rect 4729 3552 4741 3564
rect 4751 3552 4763 3564
rect 4713 3450 4725 3462
rect 4693 3430 4705 3442
rect 4754 3520 4766 3532
rect 4774 3506 4786 3518
rect 4794 3507 4806 3519
rect 4745 3464 4757 3476
rect 4727 3430 4739 3442
rect 4894 3501 4906 3513
rect 4934 3501 4946 3513
rect 5054 3521 5066 3533
rect 5015 3467 5027 3479
rect 5154 3501 5166 3513
rect 5074 3487 5086 3499
rect 5194 3501 5206 3513
rect 5254 3507 5266 3519
rect 5297 3552 5309 3564
rect 5319 3552 5331 3564
rect 5294 3520 5306 3532
rect 5274 3506 5286 3518
rect 5303 3464 5315 3476
rect 5335 3450 5347 3462
rect 5321 3430 5333 3442
rect 5367 3548 5379 3560
rect 5421 3515 5433 3527
rect 5534 3501 5546 3513
rect 5435 3476 5447 3488
rect 5383 3444 5395 3456
rect 5355 3430 5367 3442
rect 5407 3444 5419 3456
rect 5574 3501 5586 3513
rect 5654 3521 5666 3533
rect 5634 3487 5646 3499
rect 5693 3467 5705 3479
rect 175 3261 187 3273
rect 94 3221 106 3233
rect 234 3241 246 3253
rect 214 3207 226 3219
rect 334 3221 346 3233
rect 394 3227 406 3239
rect 434 3227 446 3239
rect 534 3221 546 3233
rect 514 3207 526 3219
rect 654 3241 666 3253
rect 554 3207 566 3219
rect 694 3227 706 3239
rect 834 3227 846 3239
rect 994 3281 1006 3293
rect 973 3261 985 3273
rect 874 3227 886 3239
rect 695 3190 707 3202
rect 1134 3281 1146 3293
rect 1014 3261 1026 3273
rect 1113 3261 1125 3273
rect 1154 3261 1166 3273
rect 1234 3221 1246 3233
rect 1214 3207 1226 3219
rect 1254 3207 1266 3219
rect 1514 3281 1526 3293
rect 1493 3261 1505 3273
rect 1394 3221 1406 3233
rect 1654 3281 1666 3293
rect 1534 3261 1546 3273
rect 1633 3261 1645 3273
rect 1674 3261 1686 3273
rect 1794 3221 1806 3233
rect 1774 3207 1786 3219
rect 1914 3227 1926 3239
rect 1814 3207 1826 3219
rect 1954 3227 1966 3239
rect 2074 3221 2086 3233
rect 2054 3207 2066 3219
rect 2154 3227 2166 3239
rect 2094 3207 2106 3219
rect 2194 3227 2206 3239
rect 2354 3241 2366 3253
rect 2314 3227 2326 3239
rect 2313 3190 2325 3202
rect 2414 3227 2426 3239
rect 2555 3261 2567 3273
rect 2454 3227 2466 3239
rect 2614 3241 2626 3253
rect 2594 3207 2606 3219
rect 2834 3281 2846 3293
rect 2814 3261 2826 3273
rect 2734 3221 2746 3233
rect 2714 3207 2726 3219
rect 2754 3207 2766 3219
rect 2974 3281 2986 3293
rect 2855 3261 2867 3273
rect 2954 3261 2966 3273
rect 2995 3261 3007 3273
rect 3114 3227 3126 3239
rect 3154 3227 3166 3239
rect 3254 3227 3266 3239
rect 3294 3227 3306 3239
rect 3514 3281 3526 3293
rect 3493 3261 3505 3273
rect 3354 3221 3366 3233
rect 3534 3261 3546 3273
rect 3614 3221 3626 3233
rect 3594 3207 3606 3219
rect 3755 3261 3767 3273
rect 3634 3207 3646 3219
rect 3814 3241 3826 3253
rect 3794 3207 3806 3219
rect 3981 3284 3993 3296
rect 4033 3298 4045 3310
rect 4005 3284 4017 3296
rect 3874 3221 3886 3233
rect 3953 3252 3965 3264
rect 3967 3213 3979 3225
rect 4021 3180 4033 3192
rect 4067 3298 4079 3310
rect 4053 3278 4065 3290
rect 4085 3264 4097 3276
rect 4114 3222 4126 3234
rect 4214 3241 4226 3253
rect 4094 3208 4106 3220
rect 4069 3176 4081 3188
rect 4091 3176 4103 3188
rect 4134 3221 4146 3233
rect 4273 3261 4285 3273
rect 4234 3207 4246 3219
rect 4354 3241 4366 3253
rect 4501 3284 4513 3296
rect 4553 3298 4565 3310
rect 4525 3284 4537 3296
rect 4413 3261 4425 3273
rect 4374 3207 4386 3219
rect 4473 3252 4485 3264
rect 4487 3213 4499 3225
rect 4541 3180 4553 3192
rect 4587 3298 4599 3310
rect 4573 3278 4585 3290
rect 4605 3264 4617 3276
rect 4634 3222 4646 3234
rect 4734 3241 4746 3253
rect 4614 3208 4626 3220
rect 4589 3176 4601 3188
rect 4611 3176 4623 3188
rect 4654 3221 4666 3233
rect 4793 3261 4805 3273
rect 4754 3207 4766 3219
rect 4894 3227 4906 3239
rect 5015 3261 5027 3273
rect 4934 3227 4946 3239
rect 5074 3241 5086 3253
rect 5054 3207 5066 3219
rect 5174 3221 5186 3233
rect 5254 3227 5266 3239
rect 5294 3227 5306 3239
rect 5474 3241 5486 3253
rect 5354 3221 5366 3233
rect 5533 3261 5545 3273
rect 5494 3207 5506 3219
rect 5654 3227 5666 3239
rect 5694 3227 5706 3239
rect 113 3058 125 3070
rect 114 3021 126 3033
rect 154 3007 166 3019
rect 234 2987 246 2999
rect 374 3021 386 3033
rect 275 2987 287 2999
rect 254 2967 266 2979
rect 414 3021 426 3033
rect 554 3041 566 3053
rect 515 2987 527 2999
rect 654 3041 666 3053
rect 574 3007 586 3019
rect 634 3007 646 3019
rect 794 3041 806 3053
rect 774 3007 786 3019
rect 693 2987 705 2999
rect 934 3041 946 3053
rect 914 3007 926 3019
rect 833 2987 845 2999
rect 1074 3021 1086 3033
rect 973 2987 985 2999
rect 1114 3021 1126 3033
rect 1334 3041 1346 3053
rect 1214 3007 1226 3019
rect 1254 3007 1266 3019
rect 1314 3007 1326 3019
rect 1373 2987 1385 2999
rect 1493 2987 1505 2999
rect 1654 3041 1666 3053
rect 1534 2987 1546 2999
rect 1514 2967 1526 2979
rect 1694 3041 1706 3053
rect 1674 3027 1686 3039
rect 1814 3041 1826 3053
rect 1775 2987 1787 2999
rect 1914 3041 1926 3053
rect 1834 3007 1846 3019
rect 1894 3007 1906 3019
rect 2114 3041 2126 3053
rect 1953 2987 1965 2999
rect 2075 2987 2087 2999
rect 2134 3007 2146 3019
rect 2254 3041 2266 3053
rect 2215 2987 2227 2999
rect 2394 3041 2406 3053
rect 2274 3007 2286 3019
rect 2434 3041 2446 3053
rect 2534 3041 2546 3053
rect 2414 3027 2426 3039
rect 2574 3041 2586 3053
rect 2554 3027 2566 3039
rect 2675 3041 2687 3053
rect 2713 3041 2725 3053
rect 2654 3007 2666 3019
rect 2835 3056 2847 3068
rect 2874 3027 2886 3039
rect 2733 3007 2745 3019
rect 2854 3007 2866 3019
rect 2835 2989 2847 3001
rect 3233 3058 3245 3070
rect 3074 3021 3086 3033
rect 2934 3007 2946 3019
rect 2974 3007 2986 3019
rect 3114 3021 3126 3033
rect 3234 3021 3246 3033
rect 3334 3027 3346 3039
rect 3274 3007 3286 3019
rect 3373 3056 3385 3068
rect 3354 3007 3366 3019
rect 3373 2989 3385 3001
rect 3534 3041 3546 3053
rect 3495 2987 3507 2999
rect 3554 3007 3566 3019
rect 3674 3041 3686 3053
rect 3635 2987 3647 2999
rect 3795 3056 3807 3068
rect 3953 3058 3965 3070
rect 3834 3027 3846 3039
rect 3694 3007 3706 3019
rect 3814 3007 3826 3019
rect 3795 2989 3807 3001
rect 3954 3021 3966 3033
rect 3994 3007 4006 3019
rect 4054 3007 4066 3019
rect 4094 3007 4106 3019
rect 4174 2987 4186 2999
rect 4294 3027 4306 3039
rect 4337 3072 4349 3084
rect 4359 3072 4371 3084
rect 4334 3040 4346 3052
rect 4215 2987 4227 2999
rect 4194 2967 4206 2979
rect 4314 3026 4326 3038
rect 4343 2984 4355 2996
rect 4375 2970 4387 2982
rect 4361 2950 4373 2962
rect 4407 3068 4419 3080
rect 4461 3035 4473 3047
rect 4594 3041 4606 3053
rect 4475 2996 4487 3008
rect 4574 3007 4586 3019
rect 4734 3041 4746 3053
rect 4714 3007 4726 3019
rect 4633 2987 4645 2999
rect 4423 2964 4435 2976
rect 4395 2950 4407 2962
rect 4447 2964 4459 2976
rect 4874 3021 4886 3033
rect 4773 2987 4785 2999
rect 4914 3021 4926 3033
rect 4974 3021 4986 3033
rect 5014 3021 5026 3033
rect 5074 3027 5086 3039
rect 5117 3072 5129 3084
rect 5139 3072 5151 3084
rect 5114 3040 5126 3052
rect 5094 3026 5106 3038
rect 5123 2984 5135 2996
rect 5155 2970 5167 2982
rect 5141 2950 5153 2962
rect 5187 3068 5199 3080
rect 5241 3035 5253 3047
rect 5255 2996 5267 3008
rect 5378 3044 5390 3056
rect 5418 3044 5430 3056
rect 5458 3044 5470 3056
rect 5494 3041 5506 3053
rect 5567 3035 5579 3047
rect 5553 2996 5565 3008
rect 5203 2964 5215 2976
rect 5175 2950 5187 2962
rect 5227 2964 5239 2976
rect 5621 3068 5633 3080
rect 5581 2964 5593 2976
rect 5605 2964 5617 2976
rect 5669 3072 5681 3084
rect 5691 3072 5703 3084
rect 5653 2970 5665 2982
rect 5633 2950 5645 2962
rect 5694 3040 5706 3052
rect 5714 3026 5726 3038
rect 5734 3027 5746 3039
rect 5685 2984 5697 2996
rect 5667 2950 5679 2962
rect 74 2747 86 2759
rect 174 2761 186 2773
rect 114 2747 126 2759
rect 233 2781 245 2793
rect 194 2727 206 2739
rect 354 2741 366 2753
rect 434 2741 446 2753
rect 414 2727 426 2739
rect 574 2747 586 2759
rect 454 2727 466 2739
rect 674 2761 686 2773
rect 614 2747 626 2759
rect 714 2747 726 2759
rect 814 2747 826 2759
rect 854 2747 866 2759
rect 954 2741 966 2753
rect 715 2710 727 2722
rect 934 2727 946 2739
rect 1074 2747 1086 2759
rect 974 2727 986 2739
rect 1235 2781 1247 2793
rect 1114 2747 1126 2759
rect 1294 2761 1306 2773
rect 1354 2761 1366 2773
rect 1274 2727 1286 2739
rect 1413 2781 1425 2793
rect 1374 2727 1386 2739
rect 1535 2779 1547 2791
rect 1554 2761 1566 2773
rect 1535 2712 1547 2724
rect 1634 2761 1646 2773
rect 1674 2761 1686 2773
rect 1574 2741 1586 2753
rect 1834 2761 1846 2773
rect 1794 2747 1806 2759
rect 1793 2710 1805 2722
rect 1934 2747 1946 2759
rect 2034 2761 2046 2773
rect 1974 2747 1986 2759
rect 2093 2781 2105 2793
rect 2054 2727 2066 2739
rect 2254 2761 2266 2773
rect 2214 2747 2226 2759
rect 2213 2710 2225 2722
rect 2334 2747 2346 2759
rect 2454 2761 2466 2773
rect 2634 2801 2646 2813
rect 2613 2781 2625 2793
rect 2494 2761 2506 2773
rect 2374 2747 2386 2759
rect 2654 2781 2666 2793
rect 2794 2761 2806 2773
rect 2874 2761 2886 2773
rect 2754 2747 2766 2759
rect 2753 2710 2765 2722
rect 3074 2801 3086 2813
rect 2933 2781 2945 2793
rect 3053 2781 3065 2793
rect 2894 2727 2906 2739
rect 3094 2781 3106 2793
rect 3154 2747 3166 2759
rect 3295 2781 3307 2793
rect 3194 2747 3206 2759
rect 3354 2761 3366 2773
rect 3334 2727 3346 2739
rect 3494 2761 3506 2773
rect 3554 2761 3566 2773
rect 3694 2801 3706 2813
rect 3674 2781 3686 2793
rect 3594 2761 3606 2773
rect 3454 2747 3466 2759
rect 3453 2710 3465 2722
rect 3715 2781 3727 2793
rect 3814 2747 3826 2759
rect 3854 2747 3866 2759
rect 4055 2781 4067 2793
rect 3974 2727 3986 2739
rect 4114 2761 4126 2773
rect 4094 2727 4106 2739
rect 4174 2747 4186 2759
rect 4214 2747 4226 2759
rect 4501 2804 4513 2816
rect 4553 2818 4565 2830
rect 4525 2804 4537 2816
rect 4394 2741 4406 2753
rect 4294 2727 4306 2739
rect 4473 2772 4485 2784
rect 4487 2733 4499 2745
rect 4541 2700 4553 2712
rect 4587 2818 4599 2830
rect 4573 2798 4585 2810
rect 4605 2784 4617 2796
rect 4634 2742 4646 2754
rect 4781 2818 4793 2830
rect 4763 2784 4775 2796
rect 4614 2728 4626 2740
rect 4589 2696 4601 2708
rect 4611 2696 4623 2708
rect 4654 2741 4666 2753
rect 4714 2741 4726 2753
rect 4734 2742 4746 2754
rect 4754 2728 4766 2740
rect 4815 2818 4827 2830
rect 4795 2798 4807 2810
rect 4757 2696 4769 2708
rect 4779 2696 4791 2708
rect 4843 2804 4855 2816
rect 4867 2804 4879 2816
rect 4827 2700 4839 2712
rect 4895 2772 4907 2784
rect 4881 2733 4893 2745
rect 4994 2761 5006 2773
rect 5053 2781 5065 2793
rect 5014 2727 5026 2739
rect 5134 2747 5146 2759
rect 5381 2804 5393 2816
rect 5433 2818 5445 2830
rect 5405 2804 5417 2816
rect 5174 2747 5186 2759
rect 5254 2727 5266 2739
rect 5353 2772 5365 2784
rect 5367 2733 5379 2745
rect 5421 2700 5433 2712
rect 5467 2818 5479 2830
rect 5453 2798 5465 2810
rect 5485 2784 5497 2796
rect 5514 2742 5526 2754
rect 5614 2761 5626 2773
rect 5494 2728 5506 2740
rect 5469 2696 5481 2708
rect 5491 2696 5503 2708
rect 5534 2741 5546 2753
rect 5673 2781 5685 2793
rect 5634 2727 5646 2739
rect 94 2547 106 2559
rect 154 2547 166 2559
rect 294 2561 306 2573
rect 334 2561 346 2573
rect 314 2547 326 2559
rect 394 2507 406 2519
rect 534 2547 546 2559
rect 435 2507 447 2519
rect 414 2487 426 2499
rect 774 2561 786 2573
rect 634 2527 646 2539
rect 674 2527 686 2539
rect 754 2527 766 2539
rect 914 2561 926 2573
rect 954 2561 966 2573
rect 934 2547 946 2559
rect 813 2507 825 2519
rect 1114 2561 1126 2573
rect 1075 2507 1087 2519
rect 1214 2541 1226 2553
rect 1134 2527 1146 2539
rect 1254 2541 1266 2553
rect 1355 2578 1367 2590
rect 1354 2541 1366 2553
rect 1314 2527 1326 2539
rect 1493 2507 1505 2519
rect 1594 2547 1606 2559
rect 1534 2507 1546 2519
rect 1514 2487 1526 2499
rect 1714 2561 1726 2573
rect 1694 2527 1706 2539
rect 1894 2561 1906 2573
rect 1753 2507 1765 2519
rect 1855 2507 1867 2519
rect 1994 2561 2006 2573
rect 1914 2527 1926 2539
rect 1974 2527 1986 2539
rect 2033 2507 2045 2519
rect 2153 2507 2165 2519
rect 2294 2561 2306 2573
rect 2194 2507 2206 2519
rect 2174 2487 2186 2499
rect 2334 2561 2346 2573
rect 2314 2547 2326 2559
rect 2394 2541 2406 2553
rect 2434 2541 2446 2553
rect 2594 2561 2606 2573
rect 2555 2507 2567 2519
rect 2694 2561 2706 2573
rect 2614 2527 2626 2539
rect 2674 2527 2686 2539
rect 2854 2561 2866 2573
rect 2733 2507 2745 2519
rect 2894 2561 2906 2573
rect 2874 2547 2886 2559
rect 2994 2547 3006 2559
rect 3074 2561 3086 2573
rect 3054 2527 3066 2539
rect 3214 2541 3226 2553
rect 3113 2507 3125 2519
rect 3254 2541 3266 2553
rect 3373 2507 3385 2519
rect 3515 2578 3527 2590
rect 3514 2541 3526 2553
rect 3474 2527 3486 2539
rect 3414 2507 3426 2519
rect 3394 2487 3406 2499
rect 3614 2541 3626 2553
rect 3654 2541 3666 2553
rect 3755 2561 3767 2573
rect 3793 2561 3805 2573
rect 3735 2527 3747 2539
rect 4046 2560 4058 2572
rect 3814 2527 3826 2539
rect 3894 2527 3906 2539
rect 3934 2527 3946 2539
rect 4078 2560 4090 2572
rect 4045 2503 4057 2515
rect 4094 2528 4106 2540
rect 4064 2470 4076 2482
rect 4129 2578 4141 2590
rect 4258 2596 4270 2608
rect 4162 2578 4174 2590
rect 4214 2578 4226 2590
rect 4150 2533 4162 2545
rect 4109 2470 4121 2482
rect 4301 2575 4313 2587
rect 4267 2559 4279 2571
rect 4219 2545 4231 2557
rect 4194 2472 4206 2484
rect 4292 2529 4304 2541
rect 4323 2543 4335 2555
rect 4361 2519 4373 2531
rect 4378 2499 4390 2511
rect 4402 2578 4414 2590
rect 4486 2578 4498 2590
rect 4414 2541 4426 2553
rect 4400 2482 4412 2494
rect 4474 2541 4486 2553
rect 4587 2575 4599 2587
rect 4630 2596 4642 2608
rect 4565 2543 4577 2555
rect 4527 2519 4539 2531
rect 4510 2499 4522 2511
rect 4488 2482 4500 2494
rect 4621 2559 4633 2571
rect 4596 2529 4608 2541
rect 4674 2578 4686 2590
rect 4726 2578 4738 2590
rect 4669 2545 4681 2557
rect 4759 2578 4771 2590
rect 4738 2533 4750 2545
rect 4694 2472 4706 2484
rect 4810 2560 4822 2572
rect 4794 2528 4806 2540
rect 4842 2560 4854 2572
rect 4843 2503 4855 2515
rect 4779 2470 4791 2482
rect 4824 2470 4836 2482
rect 4954 2547 4966 2559
rect 4997 2592 5009 2604
rect 5019 2592 5031 2604
rect 4994 2560 5006 2572
rect 4974 2546 4986 2558
rect 5003 2504 5015 2516
rect 5035 2490 5047 2502
rect 5021 2470 5033 2482
rect 5067 2588 5079 2600
rect 5121 2555 5133 2567
rect 5135 2516 5147 2528
rect 5258 2564 5270 2576
rect 5298 2564 5310 2576
rect 5338 2564 5350 2576
rect 5374 2561 5386 2573
rect 5494 2561 5506 2573
rect 5530 2564 5542 2576
rect 5570 2564 5582 2576
rect 5610 2564 5622 2576
rect 5714 2561 5726 2573
rect 5083 2484 5095 2496
rect 5055 2470 5067 2482
rect 5107 2484 5119 2496
rect 85 2298 97 2310
rect 234 2321 246 2333
rect 213 2301 225 2313
rect 114 2281 126 2293
rect 85 2230 97 2242
rect 254 2301 266 2313
rect 314 2267 326 2279
rect 434 2281 446 2293
rect 354 2267 366 2279
rect 493 2301 505 2313
rect 595 2301 607 2313
rect 454 2247 466 2259
rect 794 2321 806 2333
rect 773 2301 785 2313
rect 654 2281 666 2293
rect 634 2247 646 2259
rect 814 2301 826 2313
rect 894 2267 906 2279
rect 1035 2299 1047 2311
rect 1054 2281 1066 2293
rect 934 2267 946 2279
rect 1035 2232 1047 2244
rect 1074 2261 1086 2273
rect 1294 2321 1306 2333
rect 1273 2301 1285 2313
rect 1134 2247 1146 2259
rect 1314 2301 1326 2313
rect 1555 2301 1567 2313
rect 1434 2261 1446 2273
rect 1414 2247 1426 2259
rect 1454 2247 1466 2259
rect 1614 2281 1626 2293
rect 1594 2247 1606 2259
rect 1874 2321 1886 2333
rect 1853 2301 1865 2313
rect 1734 2261 1746 2273
rect 1714 2247 1726 2259
rect 1754 2247 1766 2259
rect 2014 2321 2026 2333
rect 1894 2301 1906 2313
rect 1993 2301 2005 2313
rect 2034 2301 2046 2313
rect 2144 2338 2156 2350
rect 2189 2338 2201 2350
rect 2125 2305 2137 2317
rect 2126 2248 2138 2260
rect 2174 2280 2186 2292
rect 2158 2248 2170 2260
rect 2274 2336 2286 2348
rect 2230 2275 2242 2287
rect 2209 2230 2221 2242
rect 2299 2263 2311 2275
rect 2242 2230 2254 2242
rect 2294 2230 2306 2242
rect 2372 2279 2384 2291
rect 2347 2249 2359 2261
rect 2480 2326 2492 2338
rect 2458 2309 2470 2321
rect 2441 2289 2453 2301
rect 2403 2265 2415 2277
rect 2338 2212 2350 2224
rect 2381 2233 2393 2245
rect 2605 2298 2617 2310
rect 2494 2267 2506 2279
rect 2634 2281 2646 2293
rect 2714 2281 2726 2293
rect 2482 2230 2494 2242
rect 2605 2230 2617 2242
rect 2773 2301 2785 2313
rect 2734 2247 2746 2259
rect 2854 2281 2866 2293
rect 2913 2301 2925 2313
rect 2874 2247 2886 2259
rect 3014 2267 3026 2279
rect 3054 2267 3066 2279
rect 3134 2267 3146 2279
rect 3174 2267 3186 2279
rect 3314 2261 3326 2273
rect 3294 2247 3306 2259
rect 3394 2281 3406 2293
rect 3434 2281 3446 2293
rect 3534 2281 3546 2293
rect 3334 2247 3346 2259
rect 3593 2301 3605 2313
rect 3554 2247 3566 2259
rect 3674 2267 3686 2279
rect 3823 2298 3835 2310
rect 3794 2281 3806 2293
rect 3714 2267 3726 2279
rect 3964 2338 3976 2350
rect 4009 2338 4021 2350
rect 3945 2305 3957 2317
rect 3946 2248 3958 2260
rect 3823 2230 3835 2242
rect 3994 2280 4006 2292
rect 3978 2248 3990 2260
rect 4094 2336 4106 2348
rect 4050 2275 4062 2287
rect 4029 2230 4041 2242
rect 4119 2263 4131 2275
rect 4062 2230 4074 2242
rect 4114 2230 4126 2242
rect 4192 2279 4204 2291
rect 4167 2249 4179 2261
rect 4300 2326 4312 2338
rect 4278 2309 4290 2321
rect 4261 2289 4273 2301
rect 4223 2265 4235 2277
rect 4158 2212 4170 2224
rect 4201 2233 4213 2245
rect 4394 2281 4406 2293
rect 4314 2267 4326 2279
rect 4302 2230 4314 2242
rect 4434 2267 4446 2279
rect 4535 2281 4547 2293
rect 4435 2230 4447 2242
rect 4614 2281 4626 2293
rect 4555 2247 4567 2259
rect 4593 2247 4605 2259
rect 4694 2267 4706 2279
rect 4845 2298 4857 2310
rect 4874 2281 4886 2293
rect 4734 2267 4746 2279
rect 4845 2230 4857 2242
rect 5035 2281 5047 2293
rect 4934 2261 4946 2273
rect 5114 2281 5126 2293
rect 5055 2247 5067 2259
rect 5093 2247 5105 2259
rect 5194 2267 5206 2279
rect 5234 2267 5246 2279
rect 5414 2267 5426 2279
rect 5314 2247 5326 2259
rect 5454 2267 5466 2279
rect 5534 2261 5546 2273
rect 5655 2281 5667 2293
rect 5635 2247 5647 2259
rect 5675 2278 5687 2290
rect 5714 2281 5726 2293
rect 105 2098 117 2110
rect 134 2047 146 2059
rect 105 2030 117 2042
rect 253 2027 265 2039
rect 354 2081 366 2093
rect 394 2081 406 2093
rect 374 2067 386 2079
rect 294 2027 306 2039
rect 274 2007 286 2019
rect 534 2067 546 2079
rect 654 2081 666 2093
rect 615 2027 627 2039
rect 774 2081 786 2093
rect 674 2047 686 2059
rect 814 2081 826 2093
rect 794 2067 806 2079
rect 874 2027 886 2039
rect 915 2027 927 2039
rect 894 2007 906 2019
rect 1073 2027 1085 2039
rect 1234 2081 1246 2093
rect 1114 2027 1126 2039
rect 1195 2027 1207 2039
rect 1094 2007 1106 2019
rect 1254 2047 1266 2059
rect 1374 2081 1386 2093
rect 1335 2027 1347 2039
rect 1494 2081 1506 2093
rect 1394 2047 1406 2059
rect 1534 2081 1546 2093
rect 1514 2067 1526 2079
rect 1633 2027 1645 2039
rect 1754 2081 1766 2093
rect 1734 2047 1746 2059
rect 1674 2027 1686 2039
rect 1654 2007 1666 2019
rect 1874 2081 1886 2093
rect 1914 2081 1926 2093
rect 1894 2067 1906 2079
rect 1793 2027 1805 2039
rect 2114 2081 2126 2093
rect 2094 2047 2106 2059
rect 2154 2047 2166 2059
rect 2273 2027 2285 2039
rect 2406 2080 2418 2092
rect 2314 2027 2326 2039
rect 2294 2007 2306 2019
rect 2438 2080 2450 2092
rect 2405 2023 2417 2035
rect 2454 2048 2466 2060
rect 2424 1990 2436 2002
rect 2489 2098 2501 2110
rect 2618 2116 2630 2128
rect 2522 2098 2534 2110
rect 2574 2098 2586 2110
rect 2510 2053 2522 2065
rect 2469 1990 2481 2002
rect 2661 2095 2673 2107
rect 2627 2079 2639 2091
rect 2579 2065 2591 2077
rect 2554 1992 2566 2004
rect 2652 2049 2664 2061
rect 2683 2063 2695 2075
rect 2721 2039 2733 2051
rect 2738 2019 2750 2031
rect 2762 2098 2774 2110
rect 2774 2061 2786 2073
rect 2760 2002 2772 2014
rect 2874 2081 2886 2093
rect 2854 2047 2866 2059
rect 3014 2061 3026 2073
rect 2913 2027 2925 2039
rect 3054 2061 3066 2073
rect 3114 2061 3126 2073
rect 3154 2061 3166 2073
rect 3413 2098 3425 2110
rect 3254 2047 3266 2059
rect 3294 2047 3306 2059
rect 3414 2061 3426 2073
rect 3514 2081 3526 2093
rect 3454 2047 3466 2059
rect 3554 2081 3566 2093
rect 3534 2067 3546 2079
rect 3714 2081 3726 2093
rect 3794 2027 3806 2039
rect 3954 2081 3966 2093
rect 3835 2027 3847 2039
rect 3814 2007 3826 2019
rect 4113 2098 4125 2110
rect 4114 2061 4126 2073
rect 4234 2061 4246 2073
rect 4154 2047 4166 2059
rect 4274 2061 4286 2073
rect 4394 2081 4406 2093
rect 4355 2027 4367 2039
rect 4494 2081 4506 2093
rect 4414 2047 4426 2059
rect 4474 2047 4486 2059
rect 4614 2061 4626 2073
rect 4533 2027 4545 2039
rect 4654 2061 4666 2073
rect 4734 2061 4746 2073
rect 4774 2061 4786 2073
rect 4934 2081 4946 2093
rect 4895 2027 4907 2039
rect 4954 2047 4966 2059
rect 5074 2081 5086 2093
rect 5035 2027 5047 2039
rect 5154 2067 5166 2079
rect 5094 2047 5106 2059
rect 5374 2061 5386 2073
rect 5254 2047 5266 2059
rect 5294 2047 5306 2059
rect 5414 2061 5426 2073
rect 5494 2067 5506 2079
rect 5634 2067 5646 2079
rect 5714 2081 5726 2093
rect 5694 2047 5706 2059
rect 5753 2027 5765 2039
rect 114 1841 126 1853
rect 93 1821 105 1833
rect 134 1821 146 1833
rect 214 1781 226 1793
rect 194 1767 206 1779
rect 355 1821 367 1833
rect 234 1767 246 1779
rect 534 1841 546 1853
rect 513 1821 525 1833
rect 414 1801 426 1813
rect 394 1767 406 1779
rect 554 1821 566 1833
rect 654 1801 666 1813
rect 694 1801 706 1813
rect 774 1781 786 1793
rect 754 1767 766 1779
rect 794 1767 806 1779
rect 1055 1821 1067 1833
rect 954 1781 966 1793
rect 1195 1821 1207 1833
rect 1114 1801 1126 1813
rect 1094 1767 1106 1779
rect 1254 1801 1266 1813
rect 1234 1767 1246 1779
rect 1435 1821 1447 1833
rect 1354 1781 1366 1793
rect 1494 1801 1506 1813
rect 1554 1801 1566 1813
rect 1474 1767 1486 1779
rect 1613 1821 1625 1833
rect 1715 1821 1727 1833
rect 1574 1767 1586 1779
rect 1774 1801 1786 1813
rect 1754 1767 1766 1779
rect 1854 1787 1866 1799
rect 1894 1787 1906 1799
rect 1974 1787 1986 1799
rect 2014 1787 2026 1799
rect 2264 1858 2276 1870
rect 2309 1858 2321 1870
rect 2245 1825 2257 1837
rect 2154 1767 2166 1779
rect 2246 1768 2258 1780
rect 2294 1800 2306 1812
rect 2278 1768 2290 1780
rect 2394 1856 2406 1868
rect 2350 1795 2362 1807
rect 2329 1750 2341 1762
rect 2419 1783 2431 1795
rect 2362 1750 2374 1762
rect 2414 1750 2426 1762
rect 2492 1799 2504 1811
rect 2467 1769 2479 1781
rect 2600 1846 2612 1858
rect 2578 1829 2590 1841
rect 2561 1809 2573 1821
rect 2523 1785 2535 1797
rect 2458 1732 2470 1744
rect 2501 1753 2513 1765
rect 2614 1787 2626 1799
rect 2694 1787 2706 1799
rect 2602 1750 2614 1762
rect 2874 1841 2886 1853
rect 2853 1821 2865 1833
rect 2734 1787 2746 1799
rect 2894 1821 2906 1833
rect 2975 1821 2987 1833
rect 3034 1801 3046 1813
rect 3094 1801 3106 1813
rect 3134 1801 3146 1813
rect 3014 1767 3026 1779
rect 3235 1801 3247 1813
rect 3215 1767 3227 1779
rect 3255 1798 3267 1810
rect 3294 1801 3306 1813
rect 3474 1801 3486 1813
rect 3414 1781 3426 1793
rect 3655 1821 3667 1833
rect 3553 1801 3565 1813
rect 3494 1767 3506 1779
rect 3530 1767 3542 1779
rect 3815 1821 3827 1833
rect 3714 1801 3726 1813
rect 3694 1767 3706 1779
rect 3874 1801 3886 1813
rect 3934 1801 3946 1813
rect 3854 1767 3866 1779
rect 3993 1821 4005 1833
rect 3954 1767 3966 1779
rect 4094 1787 4106 1799
rect 4214 1801 4226 1813
rect 4134 1787 4146 1799
rect 4293 1801 4305 1813
rect 4235 1767 4247 1779
rect 4273 1767 4285 1779
rect 4374 1787 4386 1799
rect 4474 1801 4486 1813
rect 4414 1787 4426 1799
rect 4533 1821 4545 1833
rect 4494 1767 4506 1779
rect 4694 1801 4706 1813
rect 4774 1801 4786 1813
rect 4814 1801 4826 1813
rect 4654 1787 4666 1799
rect 4653 1750 4665 1762
rect 4894 1787 4906 1799
rect 5014 1801 5026 1813
rect 4934 1787 4946 1799
rect 5093 1801 5105 1813
rect 5035 1767 5047 1779
rect 5073 1767 5085 1779
rect 5274 1801 5286 1813
rect 5314 1801 5326 1813
rect 5374 1801 5386 1813
rect 5194 1781 5206 1793
rect 5433 1821 5445 1833
rect 5535 1821 5547 1833
rect 5394 1767 5406 1779
rect 5594 1801 5606 1813
rect 5574 1767 5586 1779
rect 5654 1767 5666 1779
rect 74 1547 86 1559
rect 115 1547 127 1559
rect 94 1527 106 1539
rect 253 1547 265 1559
rect 354 1601 366 1613
rect 394 1601 406 1613
rect 374 1587 386 1599
rect 294 1547 306 1559
rect 274 1527 286 1539
rect 534 1601 546 1613
rect 574 1601 586 1613
rect 554 1587 566 1599
rect 634 1581 646 1593
rect 674 1581 686 1593
rect 754 1587 766 1599
rect 914 1601 926 1613
rect 875 1547 887 1559
rect 934 1567 946 1579
rect 1033 1547 1045 1559
rect 1154 1581 1166 1593
rect 1074 1547 1086 1559
rect 1054 1527 1066 1539
rect 1194 1581 1206 1593
rect 1425 1618 1437 1630
rect 1574 1587 1586 1599
rect 1274 1567 1286 1579
rect 1314 1567 1326 1579
rect 1454 1567 1466 1579
rect 1425 1550 1437 1562
rect 1655 1601 1667 1613
rect 1693 1601 1705 1613
rect 1635 1567 1647 1579
rect 1826 1600 1838 1612
rect 1714 1567 1726 1579
rect 1858 1600 1870 1612
rect 1825 1543 1837 1555
rect 1874 1568 1886 1580
rect 1844 1510 1856 1522
rect 1909 1618 1921 1630
rect 2038 1636 2050 1648
rect 1942 1618 1954 1630
rect 1994 1618 2006 1630
rect 1930 1573 1942 1585
rect 1889 1510 1901 1522
rect 2081 1615 2093 1627
rect 2047 1599 2059 1611
rect 1999 1585 2011 1597
rect 1974 1512 1986 1524
rect 2072 1569 2084 1581
rect 2103 1583 2115 1595
rect 2141 1559 2153 1571
rect 2158 1539 2170 1551
rect 2182 1618 2194 1630
rect 2194 1581 2206 1593
rect 2180 1522 2192 1534
rect 2314 1601 2326 1613
rect 2294 1567 2306 1579
rect 2434 1581 2446 1593
rect 2353 1547 2365 1559
rect 2474 1581 2486 1593
rect 2614 1601 2626 1613
rect 2575 1547 2587 1559
rect 2714 1581 2726 1593
rect 2634 1567 2646 1579
rect 2754 1581 2766 1593
rect 2874 1601 2886 1613
rect 2835 1547 2847 1559
rect 2894 1567 2906 1579
rect 3014 1601 3026 1613
rect 2975 1547 2987 1559
rect 3086 1618 3098 1630
rect 3074 1581 3086 1593
rect 3034 1567 3046 1579
rect 3187 1615 3199 1627
rect 3230 1636 3242 1648
rect 3165 1583 3177 1595
rect 3127 1559 3139 1571
rect 3110 1539 3122 1551
rect 3088 1522 3100 1534
rect 3221 1599 3233 1611
rect 3196 1569 3208 1581
rect 3274 1618 3286 1630
rect 3326 1618 3338 1630
rect 3269 1585 3281 1597
rect 3359 1618 3371 1630
rect 3338 1573 3350 1585
rect 3294 1512 3306 1524
rect 3410 1600 3422 1612
rect 3394 1568 3406 1580
rect 3442 1600 3454 1612
rect 3443 1543 3455 1555
rect 3379 1510 3391 1522
rect 3424 1510 3436 1522
rect 3614 1601 3626 1613
rect 3654 1601 3666 1613
rect 3634 1587 3646 1599
rect 3734 1601 3746 1613
rect 3714 1567 3726 1579
rect 3885 1618 3897 1630
rect 4013 1618 4025 1630
rect 3914 1567 3926 1579
rect 3773 1547 3785 1559
rect 3885 1550 3897 1562
rect 4014 1581 4026 1593
rect 4114 1581 4126 1593
rect 4054 1567 4066 1579
rect 4154 1581 4166 1593
rect 4275 1601 4287 1613
rect 4313 1601 4325 1613
rect 4254 1567 4266 1579
rect 4435 1601 4447 1613
rect 4473 1601 4485 1613
rect 4333 1567 4345 1579
rect 4414 1567 4426 1579
rect 4595 1601 4607 1613
rect 4633 1601 4645 1613
rect 4493 1567 4505 1579
rect 4575 1567 4587 1579
rect 4734 1581 4746 1593
rect 4654 1567 4666 1579
rect 4774 1581 4786 1593
rect 4874 1601 4886 1613
rect 4854 1567 4866 1579
rect 5033 1618 5045 1630
rect 4913 1547 4925 1559
rect 5034 1581 5046 1593
rect 5074 1567 5086 1579
rect 5154 1547 5166 1559
rect 5315 1601 5327 1613
rect 5353 1601 5365 1613
rect 5295 1567 5307 1579
rect 5195 1547 5207 1559
rect 5174 1527 5186 1539
rect 5454 1581 5466 1593
rect 5374 1567 5386 1579
rect 5494 1581 5506 1593
rect 5574 1547 5586 1559
rect 5774 1601 5786 1613
rect 5615 1547 5627 1559
rect 5594 1527 5606 1539
rect 114 1361 126 1373
rect 93 1341 105 1353
rect 134 1341 146 1353
rect 214 1301 226 1313
rect 194 1287 206 1299
rect 394 1361 406 1373
rect 373 1341 385 1353
rect 234 1287 246 1299
rect 414 1341 426 1353
rect 495 1341 507 1353
rect 635 1341 647 1353
rect 554 1321 566 1333
rect 534 1287 546 1299
rect 694 1321 706 1333
rect 674 1287 686 1299
rect 854 1321 866 1333
rect 814 1307 826 1319
rect 813 1270 825 1282
rect 914 1307 926 1319
rect 954 1307 966 1319
rect 1154 1361 1166 1373
rect 1134 1341 1146 1353
rect 1074 1301 1086 1313
rect 1175 1341 1187 1353
rect 1274 1307 1286 1319
rect 1314 1307 1326 1319
rect 1414 1307 1426 1319
rect 1454 1307 1466 1319
rect 1534 1307 1546 1319
rect 1714 1361 1726 1373
rect 1693 1341 1705 1353
rect 1574 1307 1586 1319
rect 1734 1341 1746 1353
rect 1794 1307 1806 1319
rect 1974 1361 1986 1373
rect 1953 1341 1965 1353
rect 1834 1307 1846 1319
rect 1994 1341 2006 1353
rect 2234 1361 2246 1373
rect 2213 1341 2225 1353
rect 2094 1301 2106 1313
rect 2374 1361 2386 1373
rect 2254 1341 2266 1353
rect 2353 1341 2365 1353
rect 2394 1341 2406 1353
rect 2595 1341 2607 1353
rect 2454 1301 2466 1313
rect 2654 1321 2666 1333
rect 2634 1287 2646 1299
rect 2734 1301 2746 1313
rect 2714 1287 2726 1299
rect 2875 1341 2887 1353
rect 2754 1287 2766 1299
rect 3015 1341 3027 1353
rect 2934 1321 2946 1333
rect 2914 1287 2926 1299
rect 3155 1341 3167 1353
rect 3074 1321 3086 1333
rect 3054 1287 3066 1299
rect 3214 1321 3226 1333
rect 3194 1287 3206 1299
rect 3505 1338 3517 1350
rect 3314 1301 3326 1313
rect 3374 1301 3386 1313
rect 3534 1321 3546 1333
rect 3505 1270 3517 1282
rect 3674 1301 3686 1313
rect 3654 1287 3666 1299
rect 3754 1321 3766 1333
rect 3694 1287 3706 1299
rect 3813 1341 3825 1353
rect 3774 1287 3786 1299
rect 4015 1341 4027 1353
rect 3934 1301 3946 1313
rect 4155 1341 4167 1353
rect 4074 1321 4086 1333
rect 4054 1287 4066 1299
rect 4214 1321 4226 1333
rect 4194 1287 4206 1299
rect 4435 1341 4447 1353
rect 4334 1301 4346 1313
rect 4314 1287 4326 1299
rect 4354 1287 4366 1299
rect 4494 1321 4506 1333
rect 4574 1321 4586 1333
rect 4474 1287 4486 1299
rect 4633 1341 4645 1353
rect 4594 1287 4606 1299
rect 4714 1307 4726 1319
rect 4834 1321 4846 1333
rect 4754 1307 4766 1319
rect 4893 1341 4905 1353
rect 4854 1287 4866 1299
rect 4974 1321 4986 1333
rect 5014 1321 5026 1333
rect 5094 1307 5106 1319
rect 5134 1307 5146 1319
rect 5234 1307 5246 1319
rect 5355 1341 5367 1353
rect 5274 1307 5286 1319
rect 5414 1321 5426 1333
rect 5474 1321 5486 1333
rect 5394 1287 5406 1299
rect 5533 1341 5545 1353
rect 5494 1287 5506 1299
rect 5634 1321 5646 1333
rect 5693 1341 5705 1353
rect 5654 1287 5666 1299
rect 154 1121 166 1133
rect 94 1107 106 1119
rect 194 1121 206 1133
rect 174 1107 186 1119
rect 314 1121 326 1133
rect 294 1087 306 1099
rect 454 1121 466 1133
rect 434 1087 446 1099
rect 353 1067 365 1079
rect 493 1067 505 1079
rect 613 1067 625 1079
rect 734 1121 746 1133
rect 714 1087 726 1099
rect 654 1067 666 1079
rect 634 1047 646 1059
rect 874 1121 886 1133
rect 914 1121 926 1133
rect 894 1107 906 1119
rect 773 1067 785 1079
rect 1074 1121 1086 1133
rect 1035 1067 1047 1079
rect 1254 1121 1266 1133
rect 1194 1107 1206 1119
rect 1094 1087 1106 1099
rect 1294 1121 1306 1133
rect 1274 1107 1286 1119
rect 1434 1107 1446 1119
rect 1634 1107 1646 1119
rect 1514 1087 1526 1099
rect 1554 1087 1566 1099
rect 1773 1067 1785 1079
rect 1894 1101 1906 1113
rect 1814 1067 1826 1079
rect 1794 1047 1806 1059
rect 1934 1101 1946 1113
rect 2054 1121 2066 1133
rect 2015 1067 2027 1079
rect 2074 1087 2086 1099
rect 2173 1067 2185 1079
rect 2214 1067 2226 1079
rect 2313 1067 2325 1079
rect 2194 1047 2206 1059
rect 2474 1121 2486 1133
rect 2354 1067 2366 1079
rect 2435 1067 2447 1079
rect 2334 1047 2346 1059
rect 2494 1087 2506 1099
rect 2593 1067 2605 1079
rect 2714 1107 2726 1119
rect 2634 1067 2646 1079
rect 2614 1047 2626 1059
rect 3095 1138 3107 1150
rect 3094 1101 3106 1113
rect 2814 1087 2826 1099
rect 2854 1087 2866 1099
rect 2934 1087 2946 1099
rect 2974 1087 2986 1099
rect 3054 1087 3066 1099
rect 3494 1107 3506 1119
rect 3214 1087 3226 1099
rect 3254 1087 3266 1099
rect 3354 1087 3366 1099
rect 3394 1087 3406 1099
rect 3614 1121 3626 1133
rect 3575 1067 3587 1079
rect 3634 1087 3646 1099
rect 3754 1121 3766 1133
rect 3715 1067 3727 1079
rect 3834 1101 3846 1113
rect 3774 1087 3786 1099
rect 3874 1101 3886 1113
rect 3954 1101 3966 1113
rect 3994 1101 4006 1113
rect 4194 1107 4206 1119
rect 4074 1087 4086 1099
rect 4114 1087 4126 1099
rect 4334 1121 4346 1133
rect 4374 1121 4386 1133
rect 4354 1107 4366 1119
rect 4514 1121 4526 1133
rect 4475 1067 4487 1079
rect 4634 1121 4646 1133
rect 4534 1087 4546 1099
rect 4674 1121 4686 1133
rect 4654 1107 4666 1119
rect 4754 1121 4766 1133
rect 4734 1087 4746 1099
rect 4903 1138 4915 1150
rect 4994 1107 5006 1119
rect 5094 1107 5106 1119
rect 4874 1087 4886 1099
rect 4793 1067 4805 1079
rect 4903 1070 4915 1082
rect 5214 1101 5226 1113
rect 5254 1101 5266 1113
rect 5394 1121 5406 1133
rect 5355 1067 5367 1079
rect 5414 1087 5426 1099
rect 5474 1087 5486 1099
rect 5514 1087 5526 1099
rect 5633 1067 5645 1079
rect 5774 1107 5786 1119
rect 5674 1067 5686 1079
rect 5654 1047 5666 1059
rect 114 881 126 893
rect 93 861 105 873
rect 134 861 146 873
rect 214 821 226 833
rect 194 807 206 819
rect 394 881 406 893
rect 373 861 385 873
rect 234 807 246 819
rect 414 861 426 873
rect 674 881 686 893
rect 653 861 665 873
rect 534 821 546 833
rect 514 807 526 819
rect 554 807 566 819
rect 694 861 706 873
rect 774 821 786 833
rect 754 807 766 819
rect 915 861 927 873
rect 794 807 806 819
rect 1094 881 1106 893
rect 1073 861 1085 873
rect 974 841 986 853
rect 954 807 966 819
rect 1114 861 1126 873
rect 1174 841 1186 853
rect 1374 881 1386 893
rect 1233 861 1245 873
rect 1353 861 1365 873
rect 1194 807 1206 819
rect 1394 861 1406 873
rect 1454 821 1466 833
rect 1554 827 1566 839
rect 1754 881 1766 893
rect 1733 861 1745 873
rect 1594 827 1606 839
rect 1894 881 1906 893
rect 1774 861 1786 873
rect 1873 861 1885 873
rect 1994 881 2006 893
rect 1914 861 1926 873
rect 1974 861 1986 873
rect 2015 861 2027 873
rect 2114 841 2126 853
rect 2173 861 2185 873
rect 2134 807 2146 819
rect 2254 841 2266 853
rect 2294 827 2306 839
rect 2394 821 2406 833
rect 2514 827 2526 839
rect 2295 790 2307 802
rect 2655 859 2667 871
rect 2674 841 2686 853
rect 2554 827 2566 839
rect 2655 792 2667 804
rect 2694 821 2706 833
rect 2754 827 2766 839
rect 2794 827 2806 839
rect 2894 827 2906 839
rect 2934 827 2946 839
rect 3014 821 3026 833
rect 3154 821 3166 833
rect 3254 827 3266 839
rect 3394 841 3406 853
rect 3434 841 3446 853
rect 3514 841 3526 853
rect 3554 841 3566 853
rect 3294 827 3306 839
rect 3674 821 3686 833
rect 3654 807 3666 819
rect 3875 861 3887 873
rect 3794 821 3806 833
rect 3694 807 3706 819
rect 3934 841 3946 853
rect 3914 807 3926 819
rect 3994 827 4006 839
rect 4135 861 4147 873
rect 4034 827 4046 839
rect 4275 861 4287 873
rect 4194 841 4206 853
rect 4174 807 4186 819
rect 4334 841 4346 853
rect 4314 807 4326 819
rect 4535 861 4547 873
rect 4414 821 4426 833
rect 4594 841 4606 853
rect 4574 807 4586 819
rect 4674 821 4686 833
rect 4654 807 4666 819
rect 4825 858 4837 870
rect 4694 807 4706 819
rect 4935 861 4947 873
rect 4854 841 4866 853
rect 4825 790 4837 802
rect 4994 841 5006 853
rect 4974 807 4986 819
rect 5074 821 5086 833
rect 5054 807 5066 819
rect 5235 859 5247 871
rect 5254 841 5266 853
rect 5094 807 5106 819
rect 5235 792 5247 804
rect 5474 841 5486 853
rect 5274 821 5286 833
rect 5394 821 5406 833
rect 5553 841 5565 853
rect 5634 841 5646 853
rect 5495 807 5507 819
rect 5533 807 5545 819
rect 5693 861 5705 873
rect 5654 807 5666 819
rect 93 587 105 599
rect 254 641 266 653
rect 134 587 146 599
rect 114 567 126 579
rect 294 641 306 653
rect 274 627 286 639
rect 393 587 405 599
rect 554 641 566 653
rect 434 587 446 599
rect 515 587 527 599
rect 414 567 426 579
rect 634 641 646 653
rect 574 607 586 619
rect 674 641 686 653
rect 654 627 666 639
rect 774 621 786 633
rect 814 621 826 633
rect 974 641 986 653
rect 935 587 947 599
rect 994 607 1006 619
rect 1093 587 1105 599
rect 1194 641 1206 653
rect 1234 641 1246 653
rect 1214 627 1226 639
rect 1134 587 1146 599
rect 1114 567 1126 579
rect 1374 641 1386 653
rect 1414 641 1426 653
rect 1394 627 1406 639
rect 1494 587 1506 599
rect 1694 641 1706 653
rect 1535 587 1547 599
rect 1655 587 1667 599
rect 1514 567 1526 579
rect 1714 607 1726 619
rect 1813 587 1825 599
rect 1914 641 1926 653
rect 1954 641 1966 653
rect 1934 627 1946 639
rect 1854 587 1866 599
rect 1834 567 1846 579
rect 2215 656 2227 668
rect 2254 627 2266 639
rect 2074 607 2086 619
rect 2114 607 2126 619
rect 2234 607 2246 619
rect 2215 589 2227 601
rect 2355 658 2367 670
rect 2354 621 2366 633
rect 2314 607 2326 619
rect 2454 621 2466 633
rect 2494 621 2506 633
rect 2594 621 2606 633
rect 2634 621 2646 633
rect 2834 641 2846 653
rect 2714 607 2726 619
rect 2754 607 2766 619
rect 2814 607 2826 619
rect 2974 621 2986 633
rect 2873 587 2885 599
rect 3074 641 3086 653
rect 3014 621 3026 633
rect 3114 641 3126 653
rect 3094 627 3106 639
rect 3253 587 3265 599
rect 3354 621 3366 633
rect 3294 587 3306 599
rect 3274 567 3286 579
rect 3394 621 3406 633
rect 3534 641 3546 653
rect 3495 587 3507 599
rect 3614 621 3626 633
rect 3554 607 3566 619
rect 3654 621 3666 633
rect 3794 641 3806 653
rect 3755 587 3767 599
rect 3894 641 3906 653
rect 3814 607 3826 619
rect 3874 607 3886 619
rect 4014 641 4026 653
rect 4054 641 4066 653
rect 4034 627 4046 639
rect 3933 587 3945 599
rect 4194 641 4206 653
rect 4174 607 4186 619
rect 4454 641 4466 653
rect 4354 627 4366 639
rect 4233 587 4245 599
rect 4494 641 4506 653
rect 4474 627 4486 639
rect 4614 641 4626 653
rect 4575 587 4587 599
rect 4634 607 4646 619
rect 4754 641 4766 653
rect 4715 587 4727 599
rect 4874 641 4886 653
rect 4774 607 4786 619
rect 4854 607 4866 619
rect 4994 627 5006 639
rect 4913 587 4925 599
rect 5143 658 5155 670
rect 5114 607 5126 619
rect 5143 590 5155 602
rect 5294 641 5306 653
rect 5255 587 5267 599
rect 5394 641 5406 653
rect 5314 607 5326 619
rect 5374 607 5386 619
rect 5574 641 5586 653
rect 5433 587 5445 599
rect 5535 587 5547 599
rect 5594 607 5606 619
rect 5654 607 5666 619
rect 5694 607 5706 619
rect 114 401 126 413
rect 93 381 105 393
rect 134 381 146 393
rect 215 381 227 393
rect 375 381 387 393
rect 274 361 286 373
rect 254 327 266 339
rect 554 401 566 413
rect 533 381 545 393
rect 434 361 446 373
rect 414 327 426 339
rect 574 381 586 393
rect 834 401 846 413
rect 813 381 825 393
rect 714 361 726 373
rect 674 347 686 359
rect 673 310 685 322
rect 854 381 866 393
rect 1074 401 1086 413
rect 1054 381 1066 393
rect 974 341 986 353
rect 954 327 966 339
rect 994 327 1006 339
rect 1095 381 1107 393
rect 1235 379 1247 391
rect 1394 401 1406 413
rect 1254 361 1266 373
rect 1235 312 1247 324
rect 1373 381 1385 393
rect 1274 341 1286 353
rect 1414 381 1426 393
rect 1615 381 1627 393
rect 1534 341 1546 353
rect 1674 361 1686 373
rect 1654 327 1666 339
rect 1814 361 1826 373
rect 1874 361 1886 373
rect 1914 361 1926 373
rect 1774 347 1786 359
rect 1773 310 1785 322
rect 2135 381 2147 393
rect 2014 341 2026 353
rect 2194 361 2206 373
rect 2174 327 2186 339
rect 2314 341 2326 353
rect 2294 327 2306 339
rect 2554 401 2566 413
rect 2533 381 2545 393
rect 2434 341 2446 353
rect 2334 327 2346 339
rect 2574 381 2586 393
rect 2634 361 2646 373
rect 2693 381 2705 393
rect 2654 327 2666 339
rect 2894 361 2906 373
rect 2934 361 2946 373
rect 2814 341 2826 353
rect 2994 341 3006 353
rect 3154 341 3166 353
rect 3134 327 3146 339
rect 3274 341 3286 353
rect 3174 327 3186 339
rect 3254 327 3266 339
rect 3294 327 3306 339
rect 3514 361 3526 373
rect 3434 341 3446 353
rect 3573 381 3585 393
rect 3534 327 3546 339
rect 3674 341 3686 353
rect 3654 327 3666 339
rect 3854 401 3866 413
rect 3833 381 3845 393
rect 3694 327 3706 339
rect 3874 381 3886 393
rect 3934 347 3946 359
rect 4134 401 4146 413
rect 4113 381 4125 393
rect 3974 347 3986 359
rect 4154 381 4166 393
rect 4235 381 4247 393
rect 4294 361 4306 373
rect 4274 327 4286 339
rect 4394 341 4406 353
rect 4474 347 4486 359
rect 4595 381 4607 393
rect 4514 347 4526 359
rect 4654 361 4666 373
rect 4634 327 4646 339
rect 4835 381 4847 393
rect 4754 341 4766 353
rect 4894 361 4906 373
rect 4874 327 4886 339
rect 4975 361 4987 373
rect 5135 381 5147 393
rect 4955 327 4967 339
rect 4995 358 5007 370
rect 5034 361 5046 373
rect 5194 361 5206 373
rect 5274 361 5286 373
rect 5174 327 5186 339
rect 5333 381 5345 393
rect 5294 327 5306 339
rect 5494 341 5506 353
rect 5474 327 5486 339
rect 5574 361 5586 373
rect 5514 327 5526 339
rect 5633 381 5645 393
rect 5594 327 5606 339
rect 5714 347 5726 359
rect 5754 347 5766 359
rect 93 107 105 119
rect 194 161 206 173
rect 234 161 246 173
rect 214 147 226 159
rect 134 107 146 119
rect 114 87 126 99
rect 394 161 406 173
rect 434 161 446 173
rect 414 147 426 159
rect 554 161 566 173
rect 515 107 527 119
rect 654 161 666 173
rect 574 127 586 139
rect 634 127 646 139
rect 693 107 705 119
rect 813 107 825 119
rect 914 147 926 159
rect 854 107 866 119
rect 834 87 846 99
rect 1034 161 1046 173
rect 1014 127 1026 139
rect 1154 161 1166 173
rect 1194 161 1206 173
rect 1174 147 1186 159
rect 1073 107 1085 119
rect 1455 178 1467 190
rect 1454 141 1466 153
rect 1294 127 1306 139
rect 1334 127 1346 139
rect 1414 127 1426 139
rect 1594 147 1606 159
rect 1714 161 1726 173
rect 1675 107 1687 119
rect 1814 141 1826 153
rect 1734 127 1746 139
rect 1854 141 1866 153
rect 1914 107 1926 119
rect 1955 107 1967 119
rect 1934 87 1946 99
rect 2113 107 2125 119
rect 2243 178 2255 190
rect 2354 141 2366 153
rect 2214 127 2226 139
rect 2154 107 2166 119
rect 2134 87 2146 99
rect 2243 110 2255 122
rect 2394 141 2406 153
rect 2495 178 2507 190
rect 2494 141 2506 153
rect 2454 127 2466 139
rect 2634 161 2646 173
rect 2773 178 2785 190
rect 2674 161 2686 173
rect 2654 147 2666 159
rect 2774 141 2786 153
rect 2894 141 2906 153
rect 2814 127 2826 139
rect 2934 141 2946 153
rect 3034 141 3046 153
rect 3074 141 3086 153
rect 3173 107 3185 119
rect 3314 147 3326 159
rect 3214 107 3226 119
rect 3194 87 3206 99
rect 3394 161 3406 173
rect 3374 127 3386 139
rect 3765 178 3777 190
rect 3554 147 3566 159
rect 3433 107 3445 119
rect 3634 141 3646 153
rect 3674 141 3686 153
rect 3883 178 3895 190
rect 3994 141 4006 153
rect 3794 127 3806 139
rect 3854 127 3866 139
rect 3765 110 3777 122
rect 3883 110 3895 122
rect 4034 141 4046 153
rect 4155 178 4167 190
rect 4154 141 4166 153
rect 4114 127 4126 139
rect 4394 141 4406 153
rect 4294 127 4306 139
rect 4334 127 4346 139
rect 4434 141 4446 153
rect 4553 107 4565 119
rect 4734 161 4746 173
rect 4594 107 4606 119
rect 4695 107 4707 119
rect 4574 87 4586 99
rect 4814 141 4826 153
rect 4754 127 4766 139
rect 4854 141 4866 153
rect 4994 161 5006 173
rect 4955 107 4967 119
rect 5214 141 5226 153
rect 5014 127 5026 139
rect 5074 127 5086 139
rect 5114 127 5126 139
rect 5315 161 5327 173
rect 5254 141 5266 153
rect 5335 127 5347 139
rect 5355 130 5367 142
rect 5474 147 5486 159
rect 5394 127 5406 139
rect 5614 147 5626 159
rect 5674 141 5686 153
rect 5714 141 5726 153
<< metal1 >>
rect -62 5776 5816 5778
rect -62 5764 4 5776
rect -62 5762 5816 5764
rect -62 5298 -2 5762
rect 76 5756 88 5762
rect 126 5756 138 5762
rect 202 5756 214 5762
rect 252 5756 264 5762
rect 411 5756 423 5762
rect 497 5756 509 5762
rect 537 5756 549 5762
rect 656 5756 668 5762
rect 706 5756 718 5762
rect 518 5714 529 5716
rect 557 5714 565 5716
rect 518 5708 565 5714
rect 431 5682 443 5684
rect 403 5676 443 5682
rect 99 5641 107 5676
rect 233 5641 241 5676
rect 374 5641 382 5676
rect 558 5653 565 5708
rect 791 5756 803 5762
rect 831 5756 843 5762
rect 951 5756 963 5762
rect 1057 5756 1069 5762
rect 1241 5756 1253 5762
rect 1367 5756 1379 5762
rect 1411 5756 1423 5762
rect 1511 5756 1523 5762
rect 1551 5756 1563 5762
rect 1691 5756 1703 5762
rect 1811 5756 1823 5762
rect 1851 5756 1863 5762
rect 93 5605 101 5627
rect 679 5641 687 5676
rect 815 5661 823 5716
rect 971 5682 983 5684
rect 943 5676 983 5682
rect 239 5605 247 5627
rect 75 5598 100 5605
rect 240 5598 265 5605
rect 75 5584 83 5598
rect 91 5584 143 5587
rect 103 5578 131 5584
rect 197 5584 249 5587
rect 209 5578 237 5584
rect 257 5584 265 5598
rect 374 5584 382 5627
rect 556 5611 564 5639
rect 374 5573 400 5584
rect 111 5538 123 5544
rect 217 5538 229 5544
rect 378 5538 390 5544
rect 428 5538 440 5544
rect 534 5602 564 5611
rect 673 5605 681 5627
rect 546 5600 564 5602
rect 655 5598 680 5605
rect 815 5598 823 5647
rect 914 5641 922 5676
rect 1080 5669 1097 5676
rect 1217 5677 1221 5686
rect 655 5584 663 5598
rect 799 5592 823 5598
rect 671 5584 723 5587
rect 683 5578 711 5584
rect 799 5584 811 5592
rect 914 5584 922 5627
rect 1080 5621 1087 5669
rect 1217 5633 1226 5677
rect 1275 5668 1283 5676
rect 1247 5660 1283 5668
rect 914 5573 940 5584
rect 498 5538 510 5544
rect 691 5538 703 5544
rect 829 5538 841 5544
rect 1080 5564 1087 5607
rect 1213 5584 1220 5619
rect 1236 5604 1242 5659
rect 1351 5641 1359 5676
rect 1351 5627 1353 5641
rect 1247 5592 1257 5598
rect 918 5538 930 5544
rect 968 5538 980 5544
rect 1251 5564 1257 5592
rect 1351 5584 1359 5627
rect 1394 5602 1402 5716
rect 1495 5714 1503 5716
rect 1531 5714 1542 5716
rect 1495 5708 1542 5714
rect 1495 5653 1502 5708
rect 1711 5682 1723 5684
rect 1683 5676 1723 5682
rect 1795 5714 1803 5716
rect 1917 5756 1929 5762
rect 2036 5756 2048 5762
rect 2086 5756 2098 5762
rect 1831 5714 1842 5716
rect 1795 5708 1842 5714
rect 1654 5641 1662 5676
rect 1795 5653 1802 5708
rect 1496 5611 1504 5639
rect 1496 5602 1526 5611
rect 1385 5594 1423 5602
rect 1496 5600 1514 5602
rect 1411 5584 1423 5594
rect 1351 5574 1361 5584
rect 1654 5584 1662 5627
rect 1796 5611 1804 5639
rect 1936 5633 1944 5716
rect 2162 5756 2174 5762
rect 2212 5756 2224 5762
rect 2317 5756 2329 5762
rect 2451 5756 2463 5762
rect 2491 5756 2503 5762
rect 2591 5756 2603 5762
rect 2631 5756 2643 5762
rect 2731 5756 2743 5762
rect 2771 5756 2783 5762
rect 2297 5682 2309 5684
rect 2297 5676 2337 5682
rect 2059 5641 2067 5676
rect 2193 5641 2201 5676
rect 2358 5641 2366 5676
rect 2475 5661 2483 5716
rect 2575 5714 2583 5716
rect 2611 5714 2622 5716
rect 2575 5708 2622 5714
rect 2715 5714 2723 5716
rect 2837 5756 2849 5762
rect 2877 5756 2889 5762
rect 2991 5756 3003 5762
rect 3076 5756 3088 5762
rect 3126 5756 3138 5762
rect 3247 5756 3259 5762
rect 3291 5756 3303 5762
rect 3411 5756 3423 5762
rect 3511 5756 3523 5762
rect 3551 5756 3563 5762
rect 3671 5756 3683 5762
rect 3771 5756 3783 5762
rect 2751 5714 2762 5716
rect 2715 5708 2762 5714
rect 1796 5602 1826 5611
rect 1796 5600 1814 5602
rect 1654 5573 1680 5584
rect 1057 5538 1069 5544
rect 1097 5538 1109 5544
rect 1231 5538 1243 5544
rect 1275 5538 1283 5544
rect 1381 5538 1393 5544
rect 1550 5538 1562 5544
rect 1936 5564 1944 5619
rect 2053 5605 2061 5627
rect 2199 5605 2207 5627
rect 2575 5653 2582 5708
rect 2035 5598 2060 5605
rect 2200 5598 2225 5605
rect 2035 5584 2043 5598
rect 1658 5538 1670 5544
rect 1708 5538 1720 5544
rect 1850 5538 1862 5544
rect 2051 5584 2103 5587
rect 2063 5578 2091 5584
rect 2157 5584 2209 5587
rect 2169 5578 2197 5584
rect 2217 5584 2225 5598
rect 2358 5584 2366 5627
rect 2475 5598 2483 5647
rect 2715 5653 2722 5708
rect 2857 5661 2865 5716
rect 2576 5611 2584 5639
rect 2716 5611 2724 5639
rect 2576 5602 2606 5611
rect 2576 5600 2594 5602
rect 2340 5573 2366 5584
rect 2459 5592 2483 5598
rect 2459 5584 2471 5592
rect 2716 5602 2746 5611
rect 2716 5600 2734 5602
rect 2857 5598 2865 5647
rect 2976 5633 2984 5716
rect 3099 5641 3107 5676
rect 3231 5641 3239 5676
rect 2857 5592 2881 5598
rect 2869 5584 2881 5592
rect 1917 5538 1929 5544
rect 2071 5538 2083 5544
rect 2177 5538 2189 5544
rect 2300 5538 2312 5544
rect 2350 5538 2362 5544
rect 2489 5538 2501 5544
rect 2630 5538 2642 5544
rect 2770 5538 2782 5544
rect 2976 5564 2984 5619
rect 3093 5605 3101 5627
rect 3231 5627 3233 5641
rect 3075 5598 3100 5605
rect 3075 5584 3083 5598
rect 3091 5584 3143 5587
rect 3103 5578 3131 5584
rect 3231 5584 3239 5627
rect 3274 5602 3282 5716
rect 3495 5714 3503 5716
rect 3837 5756 3849 5762
rect 3942 5756 3954 5762
rect 3992 5756 4004 5762
rect 3531 5714 3542 5716
rect 3495 5708 3542 5714
rect 3383 5669 3400 5676
rect 3393 5621 3400 5669
rect 3495 5653 3502 5708
rect 3496 5611 3504 5639
rect 3656 5633 3664 5716
rect 3756 5633 3764 5716
rect 3856 5633 3864 5716
rect 4077 5756 4089 5762
rect 4157 5756 4169 5762
rect 4215 5756 4227 5762
rect 4261 5756 4273 5762
rect 4327 5756 4339 5762
rect 4456 5756 4468 5762
rect 4506 5756 4518 5762
rect 3973 5641 3981 5676
rect 3265 5594 3303 5602
rect 3291 5584 3303 5594
rect 3231 5574 3241 5584
rect 3393 5564 3400 5607
rect 3496 5602 3526 5611
rect 3496 5600 3514 5602
rect 3656 5564 3664 5619
rect 3756 5564 3764 5619
rect 4096 5633 4104 5716
rect 4187 5702 4199 5736
rect 4241 5710 4253 5716
rect 4295 5710 4303 5716
rect 4245 5698 4267 5710
rect 4295 5696 4313 5710
rect 4193 5678 4199 5696
rect 4217 5686 4247 5692
rect 4295 5690 4303 5696
rect 3856 5564 3864 5619
rect 3979 5605 3987 5627
rect 3980 5598 4005 5605
rect 3937 5584 3989 5587
rect 2839 5538 2851 5544
rect 2991 5538 3003 5544
rect 3111 5538 3123 5544
rect 3261 5538 3273 5544
rect 3371 5538 3383 5544
rect 3411 5538 3423 5544
rect 3550 5538 3562 5544
rect 3671 5538 3683 5544
rect 3771 5538 3783 5544
rect 3949 5578 3977 5584
rect 3997 5584 4005 5598
rect 4096 5564 4104 5619
rect 4137 5613 4145 5676
rect 4159 5664 4173 5672
rect 4193 5672 4233 5678
rect 4153 5613 4167 5627
rect 4137 5599 4153 5613
rect 4227 5600 4233 5672
rect 4241 5672 4247 5686
rect 4265 5682 4303 5690
rect 4591 5756 4603 5762
rect 4631 5756 4643 5762
rect 4671 5756 4683 5762
rect 4711 5756 4723 5762
rect 4751 5756 4763 5762
rect 4851 5756 4863 5762
rect 4936 5756 4948 5762
rect 4986 5756 4998 5762
rect 4241 5666 4285 5672
rect 4297 5668 4359 5676
rect 4287 5627 4314 5634
rect 4334 5616 4340 5621
rect 4306 5608 4340 5616
rect 4294 5600 4301 5608
rect 4137 5584 4145 5599
rect 4227 5594 4301 5600
rect 4227 5592 4233 5594
rect 4294 5588 4301 5594
rect 4187 5570 4198 5578
rect 4191 5564 4198 5570
rect 4248 5576 4269 5583
rect 4353 5584 4359 5668
rect 4479 5641 4487 5676
rect 4611 5670 4623 5676
rect 4651 5670 4663 5676
rect 4691 5670 4703 5676
rect 4731 5670 4743 5676
rect 4605 5662 4623 5670
rect 4638 5662 4663 5670
rect 4678 5662 4703 5670
rect 4717 5662 4743 5670
rect 4473 5605 4481 5627
rect 4605 5633 4612 5662
rect 4607 5619 4612 5633
rect 4455 5598 4480 5605
rect 4605 5598 4612 5619
rect 4638 5616 4646 5662
rect 4678 5616 4686 5662
rect 4717 5616 4725 5662
rect 4836 5633 4844 5716
rect 5071 5756 5083 5762
rect 5111 5756 5123 5762
rect 5177 5756 5189 5762
rect 5217 5756 5229 5762
rect 5302 5756 5314 5762
rect 5352 5756 5364 5762
rect 4959 5641 4967 5676
rect 5095 5661 5103 5716
rect 5197 5661 5205 5716
rect 5437 5756 5449 5762
rect 5537 5756 5549 5762
rect 5577 5756 5589 5762
rect 5657 5756 5669 5762
rect 4630 5604 4646 5616
rect 4670 5604 4686 5616
rect 4710 5604 4725 5616
rect 4638 5598 4646 5604
rect 4678 5598 4686 5604
rect 4717 5598 4725 5604
rect 4455 5584 4463 5598
rect 4605 5591 4624 5598
rect 4606 5590 4624 5591
rect 4638 5590 4664 5598
rect 4678 5590 4703 5598
rect 4717 5590 4744 5598
rect 4248 5564 4255 5576
rect 4313 5564 4320 5570
rect 4307 5558 4320 5564
rect 4471 5584 4523 5587
rect 4612 5584 4624 5590
rect 4652 5584 4664 5590
rect 4691 5584 4703 5590
rect 4732 5584 4744 5590
rect 4483 5578 4511 5584
rect 4836 5564 4844 5619
rect 4953 5605 4961 5627
rect 4935 5598 4960 5605
rect 5095 5598 5103 5647
rect 4935 5584 4943 5598
rect 5079 5592 5103 5598
rect 5197 5598 5205 5647
rect 5333 5641 5341 5676
rect 5456 5633 5464 5716
rect 5557 5661 5565 5716
rect 5339 5605 5347 5627
rect 5340 5598 5365 5605
rect 5197 5592 5221 5598
rect 4951 5584 5003 5587
rect 4963 5578 4991 5584
rect 5079 5584 5091 5592
rect 5209 5584 5221 5592
rect 3837 5538 3849 5544
rect 3957 5538 3969 5544
rect 4077 5538 4089 5544
rect 4159 5538 4171 5544
rect 4217 5538 4229 5544
rect 4265 5538 4277 5544
rect 4327 5538 4339 5544
rect 4491 5538 4503 5544
rect 4591 5538 4603 5544
rect 4631 5538 4643 5544
rect 4671 5538 4683 5544
rect 4711 5538 4723 5544
rect 4751 5538 4763 5544
rect 4851 5538 4863 5544
rect 4971 5538 4983 5544
rect 5109 5538 5121 5544
rect 5297 5584 5349 5587
rect 5309 5578 5337 5584
rect 5357 5584 5365 5598
rect 5456 5564 5464 5619
rect 5557 5598 5565 5647
rect 5676 5633 5684 5716
rect 5557 5592 5581 5598
rect 5569 5584 5581 5592
rect 5676 5564 5684 5619
rect 5179 5538 5191 5544
rect 5317 5538 5329 5544
rect 5437 5538 5449 5544
rect 5539 5538 5551 5544
rect 5657 5538 5669 5544
rect 5822 5538 5882 5778
rect 4 5536 5882 5538
rect 5816 5524 5882 5536
rect 4 5522 5882 5524
rect 111 5516 123 5522
rect 290 5516 302 5522
rect 430 5516 442 5522
rect 570 5516 582 5522
rect 75 5462 83 5476
rect 103 5476 131 5482
rect 91 5473 143 5476
rect 75 5455 100 5462
rect 236 5458 254 5460
rect 93 5433 101 5455
rect 236 5449 266 5458
rect 376 5458 394 5460
rect 376 5449 406 5458
rect 516 5458 534 5460
rect 516 5449 546 5458
rect 658 5516 670 5522
rect 817 5516 829 5522
rect 938 5516 950 5522
rect 1098 5516 1110 5522
rect 1148 5516 1160 5522
rect 809 5476 837 5482
rect 797 5473 849 5476
rect 857 5462 865 5476
rect 706 5458 724 5460
rect 694 5449 724 5458
rect 840 5455 865 5462
rect 1094 5476 1120 5487
rect 1218 5516 1230 5522
rect 1377 5516 1389 5522
rect 1417 5516 1429 5522
rect 1570 5516 1582 5522
rect 1657 5516 1669 5522
rect 1850 5516 1862 5522
rect 1990 5516 2002 5522
rect 986 5458 1004 5460
rect 236 5421 244 5449
rect 376 5421 384 5449
rect 516 5421 524 5449
rect 716 5421 724 5449
rect 99 5384 107 5419
rect 235 5352 242 5407
rect 375 5352 382 5407
rect 515 5352 522 5407
rect 839 5433 847 5455
rect 974 5449 1004 5458
rect 996 5421 1004 5449
rect 1094 5433 1102 5476
rect 1266 5458 1284 5460
rect 718 5352 725 5407
rect 833 5384 841 5419
rect 1254 5449 1284 5458
rect 1400 5453 1407 5496
rect 1276 5421 1284 5449
rect 235 5346 282 5352
rect 235 5344 243 5346
rect 271 5344 282 5346
rect 375 5346 422 5352
rect 375 5344 383 5346
rect 411 5344 422 5346
rect 515 5346 562 5352
rect 515 5344 523 5346
rect 551 5344 562 5346
rect 678 5346 725 5352
rect 678 5344 689 5346
rect 76 5298 88 5304
rect 126 5298 138 5304
rect 251 5298 263 5304
rect 291 5298 303 5304
rect 391 5298 403 5304
rect 431 5298 443 5304
rect 531 5298 543 5304
rect 571 5298 583 5304
rect 717 5344 725 5346
rect 998 5352 1005 5407
rect 1094 5384 1102 5419
rect 1127 5397 1193 5403
rect 958 5346 1005 5352
rect 958 5344 969 5346
rect 657 5298 669 5304
rect 697 5298 709 5304
rect 802 5298 814 5304
rect 852 5298 864 5304
rect 997 5344 1005 5346
rect 1123 5378 1163 5384
rect 1151 5376 1163 5378
rect 1278 5352 1285 5407
rect 1400 5391 1407 5439
rect 1516 5458 1534 5460
rect 1516 5449 1546 5458
rect 1649 5476 1677 5482
rect 1637 5473 1689 5476
rect 1697 5462 1705 5476
rect 1680 5455 1705 5462
rect 1796 5458 1814 5460
rect 1516 5421 1524 5449
rect 1679 5433 1687 5455
rect 1796 5449 1826 5458
rect 1936 5458 1954 5460
rect 1936 5449 1966 5458
rect 2059 5516 2071 5522
rect 2231 5516 2243 5522
rect 2341 5516 2353 5522
rect 2457 5516 2469 5522
rect 2670 5516 2682 5522
rect 2810 5516 2822 5522
rect 2897 5516 2909 5522
rect 3017 5516 3029 5522
rect 3119 5516 3131 5522
rect 3258 5516 3270 5522
rect 3399 5516 3411 5522
rect 3517 5516 3525 5522
rect 3557 5516 3569 5522
rect 3730 5516 3742 5522
rect 2089 5468 2101 5476
rect 2077 5462 2101 5468
rect 1796 5421 1804 5449
rect 1936 5421 1944 5449
rect 1400 5384 1417 5391
rect 1238 5346 1285 5352
rect 1238 5344 1249 5346
rect 1277 5344 1285 5346
rect 1515 5352 1522 5407
rect 1673 5384 1681 5419
rect 1515 5346 1562 5352
rect 1515 5344 1523 5346
rect 1551 5344 1562 5346
rect 937 5298 949 5304
rect 977 5298 989 5304
rect 1131 5298 1143 5304
rect 1217 5298 1229 5304
rect 1257 5298 1269 5304
rect 1377 5298 1389 5304
rect 1531 5298 1543 5304
rect 1571 5298 1583 5304
rect 1795 5352 1802 5407
rect 1935 5352 1942 5407
rect 2077 5413 2085 5462
rect 2216 5441 2224 5496
rect 2311 5476 2321 5486
rect 2311 5433 2319 5476
rect 2371 5466 2383 5476
rect 2449 5476 2477 5482
rect 2437 5473 2489 5476
rect 2345 5458 2383 5466
rect 2497 5462 2505 5476
rect 1795 5346 1842 5352
rect 1795 5344 1803 5346
rect 1831 5344 1842 5346
rect 1935 5346 1982 5352
rect 1935 5344 1943 5346
rect 1971 5344 1982 5346
rect 2077 5344 2085 5399
rect 2216 5344 2224 5427
rect 2311 5419 2313 5433
rect 2311 5384 2319 5419
rect 1642 5298 1654 5304
rect 1692 5298 1704 5304
rect 1811 5298 1823 5304
rect 1851 5298 1863 5304
rect 1951 5298 1963 5304
rect 1991 5298 2003 5304
rect 2354 5344 2362 5458
rect 2480 5455 2505 5462
rect 2616 5458 2634 5460
rect 2479 5433 2487 5455
rect 2616 5449 2646 5458
rect 2756 5458 2774 5460
rect 2756 5449 2786 5458
rect 2889 5476 2917 5482
rect 2877 5473 2929 5476
rect 2937 5462 2945 5476
rect 2920 5455 2945 5462
rect 2616 5421 2624 5449
rect 2756 5421 2764 5449
rect 2473 5384 2481 5419
rect 2057 5298 2069 5304
rect 2097 5298 2109 5304
rect 2231 5298 2243 5304
rect 2327 5298 2339 5304
rect 2371 5298 2383 5304
rect 2615 5352 2622 5407
rect 2919 5433 2927 5455
rect 3036 5441 3044 5496
rect 3149 5468 3161 5476
rect 3137 5462 3161 5468
rect 2755 5352 2762 5407
rect 2913 5384 2921 5419
rect 2615 5346 2662 5352
rect 2615 5344 2623 5346
rect 2651 5344 2662 5346
rect 2755 5346 2802 5352
rect 2755 5344 2763 5346
rect 2791 5344 2802 5346
rect 2442 5298 2454 5304
rect 2492 5298 2504 5304
rect 2631 5298 2643 5304
rect 2671 5298 2683 5304
rect 2771 5298 2783 5304
rect 2811 5298 2823 5304
rect 3036 5344 3044 5427
rect 3137 5413 3145 5462
rect 3429 5468 3441 5476
rect 3417 5462 3441 5468
rect 3543 5468 3549 5496
rect 3543 5462 3553 5468
rect 3306 5458 3324 5460
rect 3294 5449 3324 5458
rect 3316 5421 3324 5449
rect 3417 5413 3425 5462
rect 3137 5344 3145 5399
rect 3318 5352 3325 5407
rect 3558 5401 3564 5456
rect 3580 5441 3587 5476
rect 3676 5458 3694 5460
rect 3676 5449 3706 5458
rect 3818 5516 3830 5522
rect 3868 5516 3880 5522
rect 3814 5476 3840 5487
rect 3939 5516 3951 5522
rect 4111 5516 4123 5522
rect 4249 5516 4261 5522
rect 4390 5516 4402 5522
rect 3278 5346 3325 5352
rect 3278 5344 3289 5346
rect 2882 5298 2894 5304
rect 2932 5298 2944 5304
rect 3017 5298 3029 5304
rect 3117 5298 3129 5304
rect 3157 5298 3169 5304
rect 3317 5344 3325 5346
rect 3417 5344 3425 5399
rect 3517 5392 3553 5400
rect 3517 5384 3525 5392
rect 3574 5383 3583 5427
rect 3676 5421 3684 5449
rect 3814 5433 3822 5476
rect 3969 5468 3981 5476
rect 3957 5462 3981 5468
rect 4075 5462 4083 5476
rect 4103 5476 4131 5482
rect 4091 5473 4143 5476
rect 4219 5468 4231 5476
rect 4219 5462 4243 5468
rect 3579 5374 3583 5383
rect 3675 5352 3682 5407
rect 3814 5384 3822 5419
rect 3957 5413 3965 5462
rect 4075 5455 4100 5462
rect 4093 5433 4101 5455
rect 3675 5346 3722 5352
rect 3675 5344 3683 5346
rect 3711 5344 3722 5346
rect 3843 5378 3883 5384
rect 3871 5376 3883 5378
rect 3957 5344 3965 5399
rect 4099 5384 4107 5419
rect 4235 5413 4243 5462
rect 4336 5458 4354 5460
rect 4336 5449 4366 5458
rect 4480 5516 4492 5522
rect 4530 5516 4542 5522
rect 4617 5516 4629 5522
rect 4737 5516 4749 5522
rect 4839 5516 4851 5522
rect 4897 5516 4909 5522
rect 4945 5516 4957 5522
rect 5007 5516 5019 5522
rect 5097 5516 5109 5522
rect 5179 5516 5191 5522
rect 5237 5516 5249 5522
rect 5285 5516 5297 5522
rect 5347 5516 5359 5522
rect 5457 5516 5469 5522
rect 5599 5516 5611 5522
rect 5719 5516 5731 5522
rect 4520 5476 4546 5487
rect 4336 5421 4344 5449
rect 4538 5433 4546 5476
rect 4636 5441 4644 5496
rect 4729 5476 4757 5482
rect 4717 5473 4769 5476
rect 4987 5496 5000 5502
rect 4871 5490 4878 5496
rect 4867 5482 4878 5490
rect 4928 5484 4935 5496
rect 4993 5490 5000 5496
rect 4777 5462 4785 5476
rect 4760 5455 4785 5462
rect 4817 5461 4825 5476
rect 4928 5477 4949 5484
rect 4907 5466 4913 5468
rect 4974 5466 4981 5472
rect 3257 5298 3269 5304
rect 3297 5298 3309 5304
rect 3397 5298 3409 5304
rect 3437 5298 3449 5304
rect 3547 5298 3559 5304
rect 3691 5298 3703 5304
rect 3731 5298 3743 5304
rect 3851 5298 3863 5304
rect 3937 5298 3949 5304
rect 3977 5298 3989 5304
rect 4235 5344 4243 5399
rect 4335 5352 4342 5407
rect 4538 5384 4546 5419
rect 4477 5378 4517 5384
rect 4477 5376 4489 5378
rect 4335 5346 4382 5352
rect 4335 5344 4343 5346
rect 4076 5298 4088 5304
rect 4126 5298 4138 5304
rect 4371 5344 4382 5346
rect 4636 5344 4644 5427
rect 4759 5433 4767 5455
rect 4817 5447 4833 5461
rect 4907 5460 4981 5466
rect 4753 5384 4761 5419
rect 4817 5384 4825 5447
rect 4833 5433 4847 5447
rect 4839 5388 4853 5396
rect 4907 5388 4913 5460
rect 4974 5452 4981 5460
rect 4986 5444 5020 5452
rect 5014 5439 5020 5444
rect 4967 5426 4994 5433
rect 4873 5382 4913 5388
rect 4921 5388 4965 5394
rect 4873 5364 4879 5382
rect 4921 5374 4927 5388
rect 5033 5392 5039 5476
rect 5116 5441 5124 5496
rect 5327 5496 5340 5502
rect 5211 5490 5218 5496
rect 5207 5482 5218 5490
rect 5268 5484 5275 5496
rect 5333 5490 5340 5496
rect 5157 5461 5165 5476
rect 5268 5477 5289 5484
rect 5247 5466 5253 5468
rect 5314 5466 5321 5472
rect 5157 5447 5173 5461
rect 5247 5460 5321 5466
rect 4977 5384 5039 5392
rect 4897 5368 4927 5374
rect 4945 5370 4983 5378
rect 4975 5364 4983 5370
rect 4867 5324 4879 5358
rect 4925 5350 4947 5362
rect 4975 5350 4993 5364
rect 4921 5344 4933 5350
rect 4975 5344 4983 5350
rect 5116 5344 5124 5427
rect 5157 5384 5165 5447
rect 5173 5433 5187 5447
rect 5179 5388 5193 5396
rect 5247 5388 5253 5460
rect 5314 5452 5321 5460
rect 5326 5444 5360 5452
rect 5354 5439 5360 5444
rect 5307 5426 5334 5433
rect 5213 5382 5253 5388
rect 5261 5388 5305 5394
rect 5213 5364 5219 5382
rect 5261 5374 5267 5388
rect 5373 5392 5379 5476
rect 5449 5476 5477 5482
rect 5437 5473 5489 5476
rect 5497 5462 5505 5476
rect 5629 5468 5641 5476
rect 5749 5468 5761 5476
rect 5480 5455 5505 5462
rect 5617 5462 5641 5468
rect 5479 5433 5487 5455
rect 5317 5384 5379 5392
rect 5473 5384 5481 5419
rect 5617 5413 5625 5462
rect 5697 5457 5713 5463
rect 5237 5368 5267 5374
rect 5285 5370 5323 5378
rect 5315 5364 5323 5370
rect 5207 5324 5219 5358
rect 5265 5350 5287 5362
rect 5315 5350 5333 5364
rect 5261 5344 5273 5350
rect 5315 5344 5323 5350
rect 5617 5344 5625 5399
rect 5697 5383 5703 5457
rect 5737 5462 5761 5468
rect 5737 5413 5745 5462
rect 5697 5377 5713 5383
rect 5737 5344 5745 5399
rect 4211 5298 4223 5304
rect 4251 5298 4263 5304
rect 4351 5298 4363 5304
rect 4391 5298 4403 5304
rect 4497 5298 4509 5304
rect 4617 5298 4629 5304
rect 4722 5298 4734 5304
rect 4772 5298 4784 5304
rect 4837 5298 4849 5304
rect 4895 5298 4907 5304
rect 4941 5298 4953 5304
rect 5007 5298 5019 5304
rect 5097 5298 5109 5304
rect 5177 5298 5189 5304
rect 5235 5298 5247 5304
rect 5281 5298 5293 5304
rect 5347 5298 5359 5304
rect 5442 5298 5454 5304
rect 5492 5298 5504 5304
rect 5597 5298 5609 5304
rect 5637 5298 5649 5304
rect 5717 5298 5729 5304
rect 5757 5298 5769 5304
rect -62 5296 5816 5298
rect -62 5284 4 5296
rect -62 5282 5816 5284
rect -62 4818 -2 5282
rect 91 5276 103 5282
rect 131 5276 143 5282
rect 217 5276 229 5282
rect 337 5276 349 5282
rect 471 5276 483 5282
rect 511 5276 523 5282
rect 597 5276 609 5282
rect 771 5276 783 5282
rect 857 5276 869 5282
rect 897 5276 909 5282
rect 1031 5276 1043 5282
rect 1071 5276 1083 5282
rect 75 5234 83 5236
rect 111 5234 122 5236
rect 75 5228 122 5234
rect 75 5173 82 5228
rect 197 5202 209 5204
rect 197 5196 237 5202
rect 258 5161 266 5196
rect 76 5131 84 5159
rect 76 5122 106 5131
rect 356 5153 364 5236
rect 455 5234 463 5236
rect 491 5234 502 5236
rect 455 5228 502 5234
rect 455 5173 462 5228
rect 577 5202 589 5204
rect 577 5196 617 5202
rect 878 5234 889 5236
rect 917 5234 925 5236
rect 878 5228 925 5234
rect 791 5202 803 5204
rect 763 5196 803 5202
rect 638 5161 646 5196
rect 734 5161 742 5196
rect 918 5173 925 5228
rect 1015 5234 1023 5236
rect 1137 5276 1149 5282
rect 1271 5276 1283 5282
rect 1311 5276 1323 5282
rect 1051 5234 1062 5236
rect 1015 5228 1062 5234
rect 1015 5173 1022 5228
rect 76 5120 94 5122
rect 258 5104 266 5147
rect 130 5058 142 5064
rect 240 5093 266 5104
rect 356 5084 364 5139
rect 456 5131 464 5159
rect 456 5122 486 5131
rect 456 5120 474 5122
rect 200 5058 212 5064
rect 250 5058 262 5064
rect 638 5104 646 5147
rect 337 5058 349 5064
rect 510 5058 522 5064
rect 620 5093 646 5104
rect 734 5104 742 5147
rect 916 5131 924 5159
rect 734 5093 760 5104
rect 580 5058 592 5064
rect 630 5058 642 5064
rect 738 5058 750 5064
rect 788 5058 800 5064
rect 894 5122 924 5131
rect 906 5120 924 5122
rect 1016 5131 1024 5159
rect 1156 5153 1164 5236
rect 1255 5234 1263 5236
rect 1416 5276 1428 5282
rect 1466 5276 1478 5282
rect 1571 5276 1583 5282
rect 1291 5234 1302 5236
rect 1255 5228 1302 5234
rect 1255 5173 1262 5228
rect 1656 5276 1668 5282
rect 1706 5276 1718 5282
rect 1931 5276 1943 5282
rect 2091 5276 2103 5282
rect 2177 5276 2189 5282
rect 2217 5276 2229 5282
rect 2331 5276 2343 5282
rect 2371 5276 2383 5282
rect 2491 5276 2503 5282
rect 2611 5276 2623 5282
rect 1439 5161 1447 5196
rect 1016 5122 1046 5131
rect 1016 5120 1034 5122
rect 1156 5084 1164 5139
rect 1256 5131 1264 5159
rect 1256 5122 1286 5131
rect 1433 5125 1441 5147
rect 1556 5153 1564 5236
rect 1807 5270 1859 5276
rect 1807 5268 1819 5270
rect 1847 5268 1859 5270
rect 1831 5196 1839 5212
rect 1883 5270 1911 5276
rect 1891 5212 1903 5216
rect 1859 5208 1903 5212
rect 1847 5206 1903 5208
rect 1911 5210 1923 5216
rect 1951 5210 1963 5216
rect 1911 5204 1963 5210
rect 2043 5270 2071 5276
rect 2083 5198 2111 5204
rect 1679 5161 1687 5196
rect 1831 5188 1854 5196
rect 1256 5120 1274 5122
rect 858 5058 870 5064
rect 1070 5058 1082 5064
rect 1415 5118 1440 5125
rect 1415 5104 1423 5118
rect 1431 5104 1483 5107
rect 1443 5098 1471 5104
rect 1556 5084 1564 5139
rect 1673 5125 1681 5147
rect 1846 5153 1854 5188
rect 2052 5190 2064 5196
rect 2052 5184 2079 5190
rect 2073 5161 2079 5184
rect 2197 5181 2205 5236
rect 2315 5234 2323 5236
rect 2351 5234 2362 5236
rect 2315 5228 2362 5234
rect 1847 5139 1854 5153
rect 1655 5118 1680 5125
rect 1587 5097 1613 5103
rect 1655 5104 1663 5118
rect 1671 5104 1723 5107
rect 1683 5098 1711 5104
rect 1846 5096 1854 5139
rect 2080 5104 2087 5147
rect 2315 5173 2322 5228
rect 2696 5276 2708 5282
rect 2746 5276 2758 5282
rect 2511 5202 2523 5204
rect 2483 5196 2523 5202
rect 2197 5118 2205 5167
rect 2454 5161 2462 5196
rect 2316 5131 2324 5159
rect 2596 5153 2604 5236
rect 2856 5276 2868 5282
rect 2906 5276 2918 5282
rect 3007 5276 3019 5282
rect 3051 5276 3063 5282
rect 3117 5276 3129 5282
rect 3291 5276 3303 5282
rect 3411 5276 3423 5282
rect 2719 5161 2727 5196
rect 2879 5161 2887 5196
rect 2991 5161 2999 5196
rect 2316 5122 2346 5131
rect 2316 5120 2334 5122
rect 2197 5112 2221 5118
rect 2209 5104 2221 5112
rect 1846 5090 1918 5096
rect 1871 5084 1878 5090
rect 1911 5084 1918 5090
rect 1137 5058 1149 5064
rect 1310 5058 1322 5064
rect 1451 5058 1463 5064
rect 1571 5058 1583 5064
rect 1691 5058 1703 5064
rect 1891 5058 1903 5064
rect 1931 5058 1945 5064
rect 2052 5058 2064 5064
rect 2108 5058 2120 5064
rect 2454 5104 2462 5147
rect 2454 5093 2480 5104
rect 2179 5058 2191 5064
rect 2370 5058 2382 5064
rect 2596 5084 2604 5139
rect 2713 5125 2721 5147
rect 2873 5125 2881 5147
rect 2991 5147 2993 5161
rect 2695 5118 2720 5125
rect 2855 5118 2880 5125
rect 2695 5104 2703 5118
rect 2711 5104 2763 5107
rect 2855 5104 2863 5118
rect 2723 5098 2751 5104
rect 2871 5104 2923 5107
rect 2883 5098 2911 5104
rect 2991 5104 2999 5147
rect 3034 5122 3042 5236
rect 3140 5189 3157 5196
rect 3140 5141 3147 5189
rect 3276 5153 3284 5236
rect 3516 5276 3528 5282
rect 3566 5276 3578 5282
rect 3637 5276 3649 5282
rect 3677 5276 3689 5282
rect 3771 5276 3783 5282
rect 3811 5276 3823 5282
rect 3911 5276 3923 5282
rect 3951 5276 3963 5282
rect 4017 5276 4029 5282
rect 4057 5276 4069 5282
rect 4176 5276 4188 5282
rect 4226 5276 4238 5282
rect 3383 5189 3400 5196
rect 3393 5141 3400 5189
rect 3539 5161 3547 5196
rect 3657 5181 3665 5236
rect 3795 5181 3803 5236
rect 3935 5181 3943 5236
rect 4038 5234 4049 5236
rect 4077 5234 4085 5236
rect 4038 5228 4085 5234
rect 3967 5197 3983 5203
rect 3025 5114 3063 5122
rect 3051 5104 3063 5114
rect 2991 5094 3001 5104
rect 3140 5084 3147 5127
rect 3276 5084 3284 5139
rect 3393 5084 3400 5127
rect 3533 5125 3541 5147
rect 3515 5118 3540 5125
rect 3657 5118 3665 5167
rect 3795 5118 3803 5167
rect 3935 5118 3943 5167
rect 3977 5143 3983 5197
rect 4078 5173 4085 5228
rect 4322 5276 4334 5282
rect 4372 5276 4384 5282
rect 4457 5276 4469 5282
rect 4591 5276 4603 5282
rect 4631 5276 4643 5282
rect 4717 5276 4729 5282
rect 4837 5276 4849 5282
rect 4937 5276 4949 5282
rect 4995 5276 5007 5282
rect 5041 5276 5053 5282
rect 5107 5276 5119 5282
rect 5202 5276 5214 5282
rect 5252 5276 5264 5282
rect 4199 5161 4207 5196
rect 4353 5161 4361 5196
rect 3977 5137 4013 5143
rect 4076 5131 4084 5159
rect 3515 5104 3523 5118
rect 3657 5112 3681 5118
rect 2458 5058 2470 5064
rect 2508 5058 2520 5064
rect 2611 5058 2623 5064
rect 2731 5058 2743 5064
rect 2891 5058 2903 5064
rect 3021 5058 3033 5064
rect 3117 5058 3129 5064
rect 3157 5058 3169 5064
rect 3291 5058 3303 5064
rect 3531 5104 3583 5107
rect 3669 5104 3681 5112
rect 3543 5098 3571 5104
rect 3779 5112 3803 5118
rect 3919 5112 3943 5118
rect 3779 5104 3791 5112
rect 3919 5104 3931 5112
rect 3371 5058 3383 5064
rect 3411 5058 3423 5064
rect 3551 5058 3563 5064
rect 3639 5058 3651 5064
rect 3809 5058 3821 5064
rect 3949 5058 3961 5064
rect 4054 5122 4084 5131
rect 4193 5125 4201 5147
rect 4476 5153 4484 5236
rect 4575 5234 4583 5236
rect 4611 5234 4622 5236
rect 4575 5228 4622 5234
rect 4575 5173 4582 5228
rect 4697 5202 4709 5204
rect 4697 5196 4737 5202
rect 4758 5161 4766 5196
rect 4860 5189 4877 5196
rect 4967 5222 4979 5256
rect 5021 5230 5033 5236
rect 5075 5230 5083 5236
rect 5025 5218 5047 5230
rect 5075 5216 5093 5230
rect 4973 5198 4979 5216
rect 4997 5206 5027 5212
rect 5075 5210 5083 5216
rect 4359 5125 4367 5147
rect 4066 5120 4084 5122
rect 4175 5118 4200 5125
rect 4360 5118 4385 5125
rect 4175 5104 4183 5118
rect 4191 5104 4243 5107
rect 4203 5098 4231 5104
rect 4317 5104 4369 5107
rect 4329 5098 4357 5104
rect 4377 5104 4385 5118
rect 4476 5084 4484 5139
rect 4576 5131 4584 5159
rect 4576 5122 4606 5131
rect 4576 5120 4594 5122
rect 4758 5104 4766 5147
rect 4860 5141 4867 5189
rect 4018 5058 4030 5064
rect 4211 5058 4223 5064
rect 4337 5058 4349 5064
rect 4457 5058 4469 5064
rect 4630 5058 4642 5064
rect 4740 5093 4766 5104
rect 4860 5084 4867 5127
rect 4917 5133 4925 5196
rect 4939 5184 4953 5192
rect 4973 5192 5013 5198
rect 4933 5133 4947 5147
rect 4917 5119 4933 5133
rect 5007 5120 5013 5192
rect 5021 5192 5027 5206
rect 5045 5202 5083 5210
rect 5337 5276 5349 5282
rect 5442 5276 5454 5282
rect 5492 5276 5504 5282
rect 5021 5186 5065 5192
rect 5077 5188 5139 5196
rect 5067 5147 5094 5154
rect 5114 5136 5120 5141
rect 5086 5128 5120 5136
rect 5074 5120 5081 5128
rect 4917 5104 4925 5119
rect 5007 5114 5081 5120
rect 5007 5112 5013 5114
rect 4700 5058 4712 5064
rect 4750 5058 4762 5064
rect 5074 5108 5081 5114
rect 4967 5090 4978 5098
rect 4971 5084 4978 5090
rect 5028 5096 5049 5103
rect 5133 5104 5139 5188
rect 5233 5161 5241 5196
rect 5356 5153 5364 5236
rect 5591 5276 5603 5282
rect 5631 5276 5643 5282
rect 5697 5276 5709 5282
rect 5737 5276 5749 5282
rect 5473 5161 5481 5196
rect 5615 5181 5623 5236
rect 5717 5181 5725 5236
rect 5239 5125 5247 5147
rect 5240 5118 5265 5125
rect 5028 5084 5035 5096
rect 5093 5084 5100 5090
rect 5087 5078 5100 5084
rect 5197 5104 5249 5107
rect 5209 5098 5237 5104
rect 5257 5104 5265 5118
rect 5356 5084 5364 5139
rect 5479 5125 5487 5147
rect 5480 5118 5505 5125
rect 5615 5118 5623 5167
rect 5437 5104 5489 5107
rect 5449 5098 5477 5104
rect 5497 5104 5505 5118
rect 5599 5112 5623 5118
rect 5717 5118 5725 5167
rect 5757 5127 5763 5193
rect 5717 5112 5741 5118
rect 5599 5104 5611 5112
rect 5729 5104 5741 5112
rect 4837 5058 4849 5064
rect 4877 5058 4889 5064
rect 4939 5058 4951 5064
rect 4997 5058 5009 5064
rect 5045 5058 5057 5064
rect 5107 5058 5119 5064
rect 5217 5058 5229 5064
rect 5337 5058 5349 5064
rect 5457 5058 5469 5064
rect 5629 5058 5641 5064
rect 5699 5058 5711 5064
rect 5822 5058 5882 5522
rect 4 5056 5882 5058
rect 5816 5044 5882 5056
rect 4 5042 5882 5044
rect 111 5036 123 5042
rect 270 5036 282 5042
rect 75 4982 83 4996
rect 103 4996 131 5002
rect 91 4993 143 4996
rect 75 4975 100 4982
rect 216 4978 234 4980
rect 93 4953 101 4975
rect 216 4969 246 4978
rect 338 5036 350 5042
rect 497 5036 509 5042
rect 669 5036 681 5042
rect 791 5036 803 5042
rect 931 5036 943 5042
rect 1038 5036 1050 5042
rect 1088 5036 1100 5042
rect 1211 5036 1223 5042
rect 1331 5036 1343 5042
rect 1449 5036 1461 5042
rect 1610 5036 1622 5042
rect 1731 5036 1743 5042
rect 1820 5036 1832 5042
rect 1870 5036 1882 5042
rect 489 4996 517 5002
rect 477 4993 529 4996
rect 537 4982 545 4996
rect 639 4988 651 4996
rect 639 4982 663 4988
rect 386 4978 404 4980
rect 374 4969 404 4978
rect 520 4975 545 4982
rect 216 4941 224 4969
rect 396 4941 404 4969
rect 99 4904 107 4939
rect 215 4872 222 4927
rect 519 4953 527 4975
rect 398 4872 405 4927
rect 513 4904 521 4939
rect 655 4933 663 4982
rect 755 4982 763 4996
rect 783 4996 811 5002
rect 771 4993 823 4996
rect 895 4982 903 4996
rect 923 4996 951 5002
rect 911 4993 963 4996
rect 1034 4996 1060 5007
rect 755 4975 780 4982
rect 895 4975 920 4982
rect 773 4953 781 4975
rect 913 4953 921 4975
rect 1034 4953 1042 4996
rect 1175 4982 1183 4996
rect 1203 4996 1231 5002
rect 1191 4993 1243 4996
rect 1175 4975 1200 4982
rect 1193 4953 1201 4975
rect 1316 4961 1324 5016
rect 1419 4988 1431 4996
rect 1419 4982 1443 4988
rect 215 4866 262 4872
rect 215 4864 223 4866
rect 251 4864 262 4866
rect 358 4866 405 4872
rect 358 4864 369 4866
rect 76 4818 88 4824
rect 126 4818 138 4824
rect 231 4818 243 4824
rect 271 4818 283 4824
rect 397 4864 405 4866
rect 655 4864 663 4919
rect 779 4904 787 4939
rect 919 4904 927 4939
rect 1034 4904 1042 4939
rect 1199 4904 1207 4939
rect 337 4818 349 4824
rect 377 4818 389 4824
rect 482 4818 494 4824
rect 532 4818 544 4824
rect 631 4818 643 4824
rect 671 4818 683 4824
rect 756 4818 768 4824
rect 806 4818 818 4824
rect 1063 4898 1103 4904
rect 1091 4896 1103 4898
rect 1316 4864 1324 4947
rect 1435 4933 1443 4982
rect 1556 4978 1574 4980
rect 1556 4969 1586 4978
rect 1695 4982 1703 4996
rect 1723 4996 1751 5002
rect 1959 5036 1971 5042
rect 2098 5036 2110 5042
rect 2148 5036 2160 5042
rect 2271 5036 2283 5042
rect 2391 5036 2403 5042
rect 2550 5036 2562 5042
rect 2651 5036 2663 5042
rect 2789 5036 2801 5042
rect 1860 4996 1886 5007
rect 1711 4993 1763 4996
rect 1695 4975 1720 4982
rect 1556 4941 1564 4969
rect 1713 4953 1721 4975
rect 1878 4953 1886 4996
rect 1989 4988 2001 4996
rect 1977 4982 2001 4988
rect 2094 4996 2120 5007
rect 1435 4864 1443 4919
rect 1555 4872 1562 4927
rect 1719 4904 1727 4939
rect 1878 4904 1886 4939
rect 1977 4933 1985 4982
rect 2094 4953 2102 4996
rect 2256 4961 2264 5016
rect 2355 4982 2363 4996
rect 2383 4996 2411 5002
rect 2371 4993 2423 4996
rect 2355 4975 2380 4982
rect 2496 4978 2514 4980
rect 2373 4953 2381 4975
rect 2496 4969 2526 4978
rect 1555 4866 1602 4872
rect 1555 4864 1563 4866
rect 896 4818 908 4824
rect 946 4818 958 4824
rect 1071 4818 1083 4824
rect 1176 4818 1188 4824
rect 1226 4818 1238 4824
rect 1331 4818 1343 4824
rect 1591 4864 1602 4866
rect 1411 4818 1423 4824
rect 1451 4818 1463 4824
rect 1571 4818 1583 4824
rect 1611 4818 1623 4824
rect 1817 4898 1857 4904
rect 1817 4896 1829 4898
rect 1977 4864 1985 4919
rect 2094 4904 2102 4939
rect 2123 4898 2163 4904
rect 2151 4896 2163 4898
rect 2256 4864 2264 4947
rect 2496 4941 2504 4969
rect 2636 4961 2644 5016
rect 2857 5036 2869 5042
rect 2958 5036 2970 5042
rect 3151 5036 3163 5042
rect 3291 5036 3303 5042
rect 3398 5036 3410 5042
rect 3448 5036 3460 5042
rect 2759 4988 2771 4996
rect 2759 4982 2783 4988
rect 2379 4904 2387 4939
rect 1696 4818 1708 4824
rect 1746 4818 1758 4824
rect 1837 4818 1849 4824
rect 1957 4818 1969 4824
rect 1997 4818 2009 4824
rect 2131 4818 2143 4824
rect 2271 4818 2283 4824
rect 2495 4872 2502 4927
rect 2495 4866 2542 4872
rect 2495 4864 2503 4866
rect 2531 4864 2542 4866
rect 2636 4864 2644 4947
rect 2775 4933 2783 4982
rect 2876 4961 2884 5016
rect 3115 4982 3123 4996
rect 3143 4996 3171 5002
rect 3131 4993 3183 4996
rect 3255 4982 3263 4996
rect 3283 4996 3311 5002
rect 3271 4993 3323 4996
rect 3394 4996 3420 5007
rect 3517 5036 3525 5042
rect 3557 5036 3569 5042
rect 3671 5036 3683 5042
rect 3711 5036 3723 5042
rect 3850 5036 3862 5042
rect 3951 5036 3963 5042
rect 3006 4978 3024 4980
rect 2994 4969 3024 4978
rect 3115 4975 3140 4982
rect 3255 4975 3280 4982
rect 2775 4864 2783 4919
rect 2807 4897 2833 4903
rect 2876 4864 2884 4947
rect 3016 4941 3024 4969
rect 3133 4953 3141 4975
rect 3273 4953 3281 4975
rect 3394 4953 3402 4996
rect 3543 4988 3549 5016
rect 3543 4982 3553 4988
rect 3018 4872 3025 4927
rect 3139 4904 3147 4939
rect 3279 4904 3287 4939
rect 3394 4904 3402 4939
rect 3558 4921 3564 4976
rect 3580 4961 3587 4996
rect 3693 4973 3700 5016
rect 3796 4978 3814 4980
rect 3796 4969 3826 4978
rect 4018 5036 4030 5042
rect 4158 5036 4170 5042
rect 4341 5036 4353 5042
rect 4457 5036 4465 5042
rect 4497 5036 4509 5042
rect 4597 5036 4609 5042
rect 4637 5036 4649 5042
rect 4771 5036 4783 5042
rect 4839 5036 4851 5042
rect 4897 5036 4909 5042
rect 4945 5036 4957 5042
rect 5007 5036 5019 5042
rect 5117 5036 5129 5042
rect 5219 5036 5231 5042
rect 5277 5036 5289 5042
rect 5325 5036 5337 5042
rect 5387 5036 5399 5042
rect 5529 5036 5541 5042
rect 3517 4912 3553 4920
rect 3517 4904 3525 4912
rect 2978 4866 3025 4872
rect 2978 4864 2989 4866
rect 2356 4818 2368 4824
rect 2406 4818 2418 4824
rect 2511 4818 2523 4824
rect 2551 4818 2563 4824
rect 2651 4818 2663 4824
rect 2751 4818 2763 4824
rect 2791 4818 2803 4824
rect 3017 4864 3025 4866
rect 2857 4818 2869 4824
rect 2957 4818 2969 4824
rect 2997 4818 3009 4824
rect 3116 4818 3128 4824
rect 3166 4818 3178 4824
rect 3423 4898 3463 4904
rect 3451 4896 3463 4898
rect 3574 4903 3583 4947
rect 3693 4911 3700 4959
rect 3796 4941 3804 4969
rect 3936 4961 3944 5016
rect 4066 4978 4084 4980
rect 4054 4969 4084 4978
rect 4311 4996 4321 5006
rect 4206 4978 4224 4980
rect 4194 4969 4224 4978
rect 3579 4894 3583 4903
rect 3683 4904 3700 4911
rect 3795 4872 3802 4927
rect 3795 4866 3842 4872
rect 3795 4864 3803 4866
rect 3831 4864 3842 4866
rect 3936 4864 3944 4947
rect 4076 4941 4084 4969
rect 4127 4957 4173 4963
rect 4216 4941 4224 4969
rect 4311 4953 4319 4996
rect 4371 4986 4383 4996
rect 4345 4978 4383 4986
rect 4483 4988 4489 5016
rect 4483 4982 4493 4988
rect 4078 4872 4085 4927
rect 4311 4939 4313 4953
rect 4218 4872 4225 4927
rect 4311 4904 4319 4939
rect 4038 4866 4085 4872
rect 4038 4864 4049 4866
rect 3256 4818 3268 4824
rect 3306 4818 3318 4824
rect 3431 4818 3443 4824
rect 3547 4818 3559 4824
rect 3711 4818 3723 4824
rect 3811 4818 3823 4824
rect 3851 4818 3863 4824
rect 3951 4818 3963 4824
rect 4077 4864 4085 4866
rect 4178 4866 4225 4872
rect 4178 4864 4189 4866
rect 4217 4864 4225 4866
rect 4354 4864 4362 4978
rect 4498 4921 4504 4976
rect 4520 4961 4527 4996
rect 4620 4973 4627 5016
rect 4735 4982 4743 4996
rect 4763 4996 4791 5002
rect 4751 4993 4803 4996
rect 4987 5016 5000 5022
rect 4871 5010 4878 5016
rect 4867 5002 4878 5010
rect 4928 5004 4935 5016
rect 4993 5010 5000 5016
rect 4735 4975 4760 4982
rect 4817 4981 4825 4996
rect 4928 4997 4949 5004
rect 4907 4986 4913 4988
rect 4974 4986 4981 4992
rect 4457 4912 4493 4920
rect 4457 4904 4465 4912
rect 4514 4903 4523 4947
rect 4620 4911 4627 4959
rect 4753 4953 4761 4975
rect 4817 4967 4833 4981
rect 4907 4980 4981 4986
rect 4620 4904 4637 4911
rect 4759 4904 4767 4939
rect 4817 4904 4825 4967
rect 4833 4953 4847 4967
rect 4839 4908 4853 4916
rect 4519 4894 4523 4903
rect 4907 4908 4913 4980
rect 4974 4972 4981 4980
rect 4986 4964 5020 4972
rect 5014 4959 5020 4964
rect 4967 4946 4994 4953
rect 4873 4902 4913 4908
rect 4921 4908 4965 4914
rect 4873 4884 4879 4902
rect 4921 4894 4927 4908
rect 5033 4912 5039 4996
rect 5109 4996 5137 5002
rect 5097 4993 5149 4996
rect 5367 5016 5380 5022
rect 5251 5010 5258 5016
rect 5247 5002 5258 5010
rect 5308 5004 5315 5016
rect 5373 5010 5380 5016
rect 5157 4982 5165 4996
rect 5140 4975 5165 4982
rect 5197 4981 5205 4996
rect 5308 4997 5329 5004
rect 5287 4986 5293 4988
rect 5354 4986 5361 4992
rect 5139 4953 5147 4975
rect 5197 4967 5213 4981
rect 5287 4980 5361 4986
rect 4977 4904 5039 4912
rect 5133 4904 5141 4939
rect 5197 4904 5205 4967
rect 5213 4953 5227 4967
rect 5219 4908 5233 4916
rect 4897 4888 4927 4894
rect 4945 4890 4983 4898
rect 4975 4884 4983 4890
rect 4867 4844 4879 4878
rect 4925 4870 4947 4882
rect 4975 4870 4993 4884
rect 4921 4864 4933 4870
rect 4975 4864 4983 4870
rect 5287 4908 5293 4980
rect 5354 4972 5361 4980
rect 5366 4964 5400 4972
rect 5394 4959 5400 4964
rect 5347 4946 5374 4953
rect 5253 4902 5293 4908
rect 5301 4908 5345 4914
rect 5253 4884 5259 4902
rect 5301 4894 5307 4908
rect 5413 4912 5419 4996
rect 5599 5036 5611 5042
rect 5739 5036 5751 5042
rect 5499 4988 5511 4996
rect 5629 4988 5641 4996
rect 5769 4988 5781 4996
rect 5499 4982 5523 4988
rect 5515 4933 5523 4982
rect 5577 4977 5593 4983
rect 5357 4904 5419 4912
rect 5277 4888 5307 4894
rect 5325 4890 5363 4898
rect 5355 4884 5363 4890
rect 5247 4844 5259 4878
rect 5305 4870 5327 4882
rect 5355 4870 5373 4884
rect 5301 4864 5313 4870
rect 5355 4864 5363 4870
rect 5515 4864 5523 4919
rect 5557 4903 5563 4973
rect 5547 4897 5563 4903
rect 5577 4903 5583 4977
rect 5617 4982 5641 4988
rect 5757 4982 5781 4988
rect 5617 4933 5625 4982
rect 5757 4933 5765 4982
rect 5577 4897 5603 4903
rect 5597 4887 5603 4897
rect 5617 4864 5625 4919
rect 5757 4864 5765 4919
rect 4017 4818 4029 4824
rect 4057 4818 4069 4824
rect 4157 4818 4169 4824
rect 4197 4818 4209 4824
rect 4327 4818 4339 4824
rect 4371 4818 4383 4824
rect 4487 4818 4499 4824
rect 4597 4818 4609 4824
rect 4736 4818 4748 4824
rect 4786 4818 4798 4824
rect 4837 4818 4849 4824
rect 4895 4818 4907 4824
rect 4941 4818 4953 4824
rect 5007 4818 5019 4824
rect 5102 4818 5114 4824
rect 5152 4818 5164 4824
rect 5217 4818 5229 4824
rect 5275 4818 5287 4824
rect 5321 4818 5333 4824
rect 5387 4818 5399 4824
rect 5491 4818 5503 4824
rect 5531 4818 5543 4824
rect 5597 4818 5609 4824
rect 5637 4818 5649 4824
rect 5737 4818 5749 4824
rect 5777 4818 5789 4824
rect -62 4816 5816 4818
rect -62 4804 4 4816
rect -62 4802 5816 4804
rect -62 4338 -2 4802
rect 111 4796 123 4802
rect 231 4796 243 4802
rect 271 4796 283 4802
rect 357 4796 369 4802
rect 477 4796 489 4802
rect 517 4796 529 4802
rect 631 4796 643 4802
rect 671 4796 683 4802
rect 791 4796 803 4802
rect 831 4796 843 4802
rect 131 4722 143 4724
rect 103 4716 143 4722
rect 215 4754 223 4756
rect 251 4754 262 4756
rect 215 4748 262 4754
rect 74 4681 82 4716
rect 215 4693 222 4748
rect 337 4722 349 4724
rect 337 4716 377 4722
rect 398 4681 406 4716
rect 497 4701 505 4756
rect 615 4754 623 4756
rect 651 4754 662 4756
rect 615 4748 662 4754
rect 775 4754 783 4756
rect 897 4796 909 4802
rect 997 4796 1009 4802
rect 1131 4796 1143 4802
rect 1216 4796 1228 4802
rect 1266 4796 1278 4802
rect 811 4754 822 4756
rect 775 4748 822 4754
rect 74 4624 82 4667
rect 216 4651 224 4679
rect 216 4642 246 4651
rect 615 4693 622 4748
rect 216 4640 234 4642
rect 74 4613 100 4624
rect 398 4624 406 4667
rect 497 4638 505 4687
rect 775 4693 782 4748
rect 616 4651 624 4679
rect 776 4651 784 4679
rect 916 4673 924 4756
rect 1016 4673 1024 4756
rect 1116 4673 1124 4756
rect 1342 4796 1354 4802
rect 1392 4796 1404 4802
rect 1477 4796 1489 4802
rect 1577 4796 1589 4802
rect 1617 4796 1629 4802
rect 1736 4796 1748 4802
rect 1786 4796 1798 4802
rect 1239 4681 1247 4716
rect 1373 4681 1381 4716
rect 616 4642 646 4651
rect 616 4640 634 4642
rect 497 4632 521 4638
rect 509 4624 521 4632
rect 78 4578 90 4584
rect 128 4578 140 4584
rect 270 4578 282 4584
rect 380 4613 406 4624
rect 340 4578 352 4584
rect 390 4578 402 4584
rect 776 4642 806 4651
rect 776 4640 794 4642
rect 916 4604 924 4659
rect 1016 4604 1024 4659
rect 1116 4604 1124 4659
rect 1233 4645 1241 4667
rect 1496 4673 1504 4756
rect 1598 4754 1609 4756
rect 1637 4754 1645 4756
rect 1598 4748 1645 4754
rect 1638 4693 1645 4748
rect 1871 4796 1883 4802
rect 1911 4796 1923 4802
rect 1982 4796 1994 4802
rect 2032 4796 2044 4802
rect 2151 4796 2163 4802
rect 2191 4796 2203 4802
rect 2289 4796 2301 4802
rect 2377 4796 2389 4802
rect 2417 4796 2429 4802
rect 1759 4681 1767 4716
rect 1895 4701 1903 4756
rect 2135 4754 2143 4756
rect 2171 4754 2182 4756
rect 2135 4748 2182 4754
rect 1379 4645 1387 4667
rect 1215 4638 1240 4645
rect 1380 4638 1405 4645
rect 1215 4624 1223 4638
rect 479 4578 491 4584
rect 670 4578 682 4584
rect 830 4578 842 4584
rect 1231 4624 1283 4627
rect 1243 4618 1271 4624
rect 1337 4624 1389 4627
rect 1349 4618 1377 4624
rect 1397 4624 1405 4638
rect 1496 4604 1504 4659
rect 1636 4651 1644 4679
rect 1614 4642 1644 4651
rect 1753 4645 1761 4667
rect 1626 4640 1644 4642
rect 1735 4638 1760 4645
rect 1895 4638 1903 4687
rect 2013 4681 2021 4716
rect 2135 4693 2142 4748
rect 2497 4796 2509 4802
rect 2537 4796 2549 4802
rect 2649 4796 2661 4802
rect 2737 4796 2749 4802
rect 2777 4796 2789 4802
rect 2931 4796 2943 4802
rect 2271 4681 2279 4716
rect 2315 4710 2323 4756
rect 2297 4704 2323 4710
rect 2297 4698 2300 4704
rect 2397 4701 2405 4756
rect 2517 4701 2525 4756
rect 2019 4645 2027 4667
rect 2136 4651 2144 4679
rect 2271 4667 2273 4681
rect 2020 4638 2045 4645
rect 2136 4642 2166 4651
rect 2136 4640 2154 4642
rect 1735 4624 1743 4638
rect 1879 4632 1903 4638
rect 1751 4624 1803 4627
rect 1763 4618 1791 4624
rect 1879 4624 1891 4632
rect 1977 4624 2029 4627
rect 1989 4618 2017 4624
rect 2037 4624 2045 4638
rect 2271 4624 2279 4667
rect 2293 4642 2300 4698
rect 2297 4636 2300 4642
rect 2397 4638 2405 4687
rect 2517 4638 2525 4687
rect 2631 4681 2639 4716
rect 2675 4710 2683 4756
rect 2758 4754 2769 4756
rect 2797 4754 2805 4756
rect 2758 4748 2805 4754
rect 2657 4704 2683 4710
rect 2657 4698 2660 4704
rect 2631 4667 2633 4681
rect 2297 4630 2319 4636
rect 2397 4632 2421 4638
rect 2517 4632 2541 4638
rect 2311 4604 2319 4630
rect 2409 4624 2421 4632
rect 2529 4624 2541 4632
rect 2631 4624 2639 4667
rect 2653 4642 2660 4698
rect 2798 4693 2805 4748
rect 3017 4796 3029 4802
rect 3087 4796 3099 4802
rect 3191 4796 3203 4802
rect 3231 4796 3243 4802
rect 3331 4796 3343 4802
rect 3371 4796 3383 4802
rect 3491 4796 3503 4802
rect 3611 4796 3623 4802
rect 3651 4796 3663 4802
rect 3771 4796 3783 4802
rect 3857 4796 3869 4802
rect 3897 4796 3909 4802
rect 3997 4796 4009 4802
rect 4037 4796 4049 4802
rect 4137 4796 4149 4802
rect 4267 4796 4279 4802
rect 4311 4796 4323 4802
rect 4431 4796 4443 4802
rect 4471 4796 4483 4802
rect 2903 4709 2920 4716
rect 2796 4651 2804 4679
rect 2657 4636 2660 4642
rect 2657 4630 2679 4636
rect 2671 4604 2679 4630
rect 2774 4642 2804 4651
rect 2786 4640 2804 4642
rect 2913 4661 2920 4709
rect 3057 4681 3065 4716
rect 3215 4701 3223 4756
rect 3315 4754 3323 4756
rect 3351 4754 3362 4756
rect 3315 4748 3362 4754
rect 2913 4604 2920 4647
rect 3056 4641 3064 4667
rect 3315 4693 3322 4748
rect 3511 4722 3523 4724
rect 3483 4716 3523 4722
rect 3595 4754 3603 4756
rect 3631 4754 3642 4756
rect 3595 4748 3642 4754
rect 3056 4634 3085 4641
rect 3215 4638 3223 4687
rect 3454 4681 3462 4716
rect 3595 4693 3602 4748
rect 3878 4754 3889 4756
rect 3917 4754 3925 4756
rect 3878 4748 3925 4754
rect 4018 4754 4029 4756
rect 4057 4754 4065 4756
rect 4018 4748 4065 4754
rect 3791 4722 3803 4724
rect 3763 4716 3803 4722
rect 3316 4651 3324 4679
rect 3734 4681 3742 4716
rect 3807 4697 3823 4703
rect 3316 4642 3346 4651
rect 3316 4640 3334 4642
rect 3017 4624 3069 4626
rect 3079 4624 3085 4634
rect 3199 4632 3223 4638
rect 3199 4624 3211 4632
rect 3029 4620 3057 4624
rect 3069 4584 3097 4590
rect 3454 4624 3462 4667
rect 3596 4651 3604 4679
rect 3596 4642 3626 4651
rect 3596 4640 3614 4642
rect 3454 4613 3480 4624
rect 897 4578 909 4584
rect 997 4578 1009 4584
rect 1131 4578 1143 4584
rect 1251 4578 1263 4584
rect 1357 4578 1369 4584
rect 1477 4578 1489 4584
rect 1578 4578 1590 4584
rect 1771 4578 1783 4584
rect 1909 4578 1921 4584
rect 1997 4578 2009 4584
rect 2190 4578 2202 4584
rect 2289 4578 2301 4584
rect 2379 4578 2391 4584
rect 2499 4578 2511 4584
rect 2649 4578 2661 4584
rect 2738 4578 2750 4584
rect 2891 4578 2903 4584
rect 2931 4578 2943 4584
rect 3037 4578 3049 4584
rect 3229 4578 3241 4584
rect 3370 4578 3382 4584
rect 3734 4624 3742 4667
rect 3817 4663 3823 4697
rect 3918 4693 3925 4748
rect 4058 4693 4065 4748
rect 3817 4657 3853 4663
rect 3916 4651 3924 4679
rect 4056 4651 4064 4679
rect 4156 4673 4164 4756
rect 4251 4681 4259 4716
rect 3734 4613 3760 4624
rect 3458 4578 3470 4584
rect 3508 4578 3520 4584
rect 3650 4578 3662 4584
rect 3738 4578 3750 4584
rect 3788 4578 3800 4584
rect 3894 4642 3924 4651
rect 3906 4640 3924 4642
rect 4034 4642 4064 4651
rect 4251 4667 4253 4681
rect 4046 4640 4064 4642
rect 4156 4604 4164 4659
rect 4251 4624 4259 4667
rect 4294 4642 4302 4756
rect 4415 4754 4423 4756
rect 4537 4796 4549 4802
rect 4577 4796 4589 4802
rect 4677 4796 4689 4802
rect 4757 4796 4769 4802
rect 4815 4796 4827 4802
rect 4861 4796 4873 4802
rect 4927 4796 4939 4802
rect 5022 4796 5034 4802
rect 5072 4796 5084 4802
rect 4451 4754 4462 4756
rect 4415 4748 4462 4754
rect 4558 4754 4569 4756
rect 4597 4754 4605 4756
rect 4558 4748 4605 4754
rect 4415 4693 4422 4748
rect 4598 4693 4605 4748
rect 4416 4651 4424 4679
rect 4596 4651 4604 4679
rect 4696 4673 4704 4756
rect 4787 4742 4799 4776
rect 4841 4750 4853 4756
rect 4895 4750 4903 4756
rect 4845 4738 4867 4750
rect 4895 4736 4913 4750
rect 4793 4718 4799 4736
rect 4817 4726 4847 4732
rect 4895 4730 4903 4736
rect 4416 4642 4446 4651
rect 4285 4634 4323 4642
rect 4416 4640 4434 4642
rect 4311 4624 4323 4634
rect 4251 4614 4261 4624
rect 3858 4578 3870 4584
rect 3998 4578 4010 4584
rect 4137 4578 4149 4584
rect 4281 4578 4293 4584
rect 4470 4578 4482 4584
rect 4574 4642 4604 4651
rect 4586 4640 4604 4642
rect 4696 4604 4704 4659
rect 4737 4653 4745 4716
rect 4759 4704 4773 4712
rect 4793 4712 4833 4718
rect 4753 4653 4767 4667
rect 4737 4639 4753 4653
rect 4827 4640 4833 4712
rect 4841 4712 4847 4726
rect 4865 4722 4903 4730
rect 5157 4796 5169 4802
rect 5197 4796 5209 4802
rect 5277 4796 5289 4802
rect 5317 4796 5329 4802
rect 5417 4796 5429 4802
rect 5457 4796 5469 4802
rect 5537 4796 5549 4802
rect 5577 4796 5589 4802
rect 5691 4796 5703 4802
rect 5731 4796 5743 4802
rect 4841 4706 4885 4712
rect 4897 4708 4959 4716
rect 4887 4667 4914 4674
rect 4934 4656 4940 4661
rect 4906 4648 4940 4656
rect 4894 4640 4901 4648
rect 4737 4624 4745 4639
rect 4827 4634 4901 4640
rect 4827 4632 4833 4634
rect 4894 4628 4901 4634
rect 4787 4610 4798 4618
rect 4791 4604 4798 4610
rect 4848 4616 4869 4623
rect 4953 4624 4959 4708
rect 5053 4681 5061 4716
rect 5177 4701 5185 4756
rect 5297 4701 5305 4756
rect 5327 4717 5343 4723
rect 5337 4703 5343 4717
rect 5387 4717 5403 4723
rect 5059 4645 5067 4667
rect 5060 4638 5085 4645
rect 4848 4604 4855 4616
rect 4913 4604 4920 4610
rect 4907 4598 4920 4604
rect 5017 4624 5069 4627
rect 5029 4618 5057 4624
rect 5077 4624 5085 4638
rect 5177 4638 5185 4687
rect 5337 4697 5373 4703
rect 5297 4638 5305 4687
rect 5397 4643 5403 4717
rect 5437 4701 5445 4756
rect 5507 4717 5533 4723
rect 5557 4701 5565 4756
rect 5675 4754 5683 4756
rect 5711 4754 5722 4756
rect 5675 4748 5722 4754
rect 5607 4717 5653 4723
rect 5177 4632 5201 4638
rect 5297 4632 5321 4638
rect 5397 4637 5413 4643
rect 5437 4638 5445 4687
rect 5675 4693 5682 4748
rect 5557 4638 5565 4687
rect 5676 4651 5684 4679
rect 5676 4642 5706 4651
rect 5676 4640 5694 4642
rect 5437 4632 5461 4638
rect 5557 4632 5581 4638
rect 5189 4624 5201 4632
rect 5309 4624 5321 4632
rect 5449 4624 5461 4632
rect 5569 4624 5581 4632
rect 4538 4578 4550 4584
rect 4677 4578 4689 4584
rect 4759 4578 4771 4584
rect 4817 4578 4829 4584
rect 4865 4578 4877 4584
rect 4927 4578 4939 4584
rect 5037 4578 5049 4584
rect 5159 4578 5171 4584
rect 5279 4578 5291 4584
rect 5419 4578 5431 4584
rect 5539 4578 5551 4584
rect 5730 4578 5742 4584
rect 5822 4578 5882 5042
rect 4 4576 5882 4578
rect 5816 4564 5882 4576
rect 4 4562 5882 4564
rect 111 4556 123 4562
rect 270 4556 282 4562
rect 75 4502 83 4516
rect 103 4516 131 4522
rect 91 4513 143 4516
rect 167 4517 193 4523
rect 75 4495 100 4502
rect 216 4498 234 4500
rect 93 4473 101 4495
rect 216 4489 246 4498
rect 340 4556 352 4562
rect 390 4556 402 4562
rect 551 4556 563 4562
rect 691 4556 703 4562
rect 777 4556 789 4562
rect 880 4556 892 4562
rect 930 4556 942 4562
rect 1051 4556 1063 4562
rect 1190 4556 1202 4562
rect 380 4516 406 4527
rect 216 4461 224 4489
rect 287 4477 313 4483
rect 398 4473 406 4516
rect 515 4502 523 4516
rect 543 4516 571 4522
rect 531 4513 583 4516
rect 655 4502 663 4516
rect 683 4516 711 4522
rect 671 4513 723 4516
rect 515 4495 540 4502
rect 655 4495 680 4502
rect 533 4473 541 4495
rect 99 4424 107 4459
rect 673 4473 681 4495
rect 796 4481 804 4536
rect 920 4516 946 4527
rect 938 4473 946 4516
rect 1036 4481 1044 4536
rect 1136 4498 1154 4500
rect 215 4392 222 4447
rect 398 4424 406 4459
rect 539 4424 547 4459
rect 679 4424 687 4459
rect 337 4418 377 4424
rect 337 4416 349 4418
rect 215 4386 262 4392
rect 215 4384 223 4386
rect 251 4384 262 4386
rect 76 4338 88 4344
rect 126 4338 138 4344
rect 231 4338 243 4344
rect 271 4338 283 4344
rect 357 4338 369 4344
rect 516 4338 528 4344
rect 566 4338 578 4344
rect 796 4384 804 4467
rect 1136 4489 1166 4498
rect 1278 4556 1290 4562
rect 1328 4556 1340 4562
rect 1431 4556 1443 4562
rect 1517 4556 1529 4562
rect 1689 4556 1701 4562
rect 1830 4556 1842 4562
rect 1274 4516 1300 4527
rect 938 4424 946 4459
rect 877 4418 917 4424
rect 877 4416 889 4418
rect 656 4338 668 4344
rect 706 4338 718 4344
rect 1036 4384 1044 4467
rect 1136 4461 1144 4489
rect 1274 4473 1282 4516
rect 1416 4481 1424 4536
rect 1509 4516 1537 4522
rect 1497 4513 1549 4516
rect 1557 4502 1565 4516
rect 1659 4508 1671 4516
rect 1659 4502 1683 4508
rect 1540 4495 1565 4502
rect 1135 4392 1142 4447
rect 1274 4424 1282 4459
rect 1135 4386 1182 4392
rect 1135 4384 1143 4386
rect 1171 4384 1182 4386
rect 1303 4418 1343 4424
rect 1331 4416 1343 4418
rect 1416 4384 1424 4467
rect 1539 4473 1547 4495
rect 1533 4424 1541 4459
rect 1675 4453 1683 4502
rect 1776 4498 1794 4500
rect 1776 4489 1806 4498
rect 1911 4556 1923 4562
rect 1951 4556 1963 4562
rect 2090 4556 2102 4562
rect 2250 4556 2262 4562
rect 2369 4556 2381 4562
rect 2510 4556 2522 4562
rect 1933 4493 1940 4536
rect 1967 4497 2013 4503
rect 2036 4498 2054 4500
rect 1776 4461 1784 4489
rect 2036 4489 2066 4498
rect 2196 4498 2214 4500
rect 2196 4489 2226 4498
rect 2339 4508 2351 4516
rect 2339 4502 2363 4508
rect 777 4338 789 4344
rect 897 4338 909 4344
rect 1051 4338 1063 4344
rect 1151 4338 1163 4344
rect 1191 4338 1203 4344
rect 1311 4338 1323 4344
rect 1431 4338 1443 4344
rect 1675 4384 1683 4439
rect 1775 4392 1782 4447
rect 1933 4431 1940 4479
rect 2036 4461 2044 4489
rect 2196 4461 2204 4489
rect 1923 4424 1940 4431
rect 1775 4386 1822 4392
rect 1775 4384 1783 4386
rect 1502 4338 1514 4344
rect 1552 4338 1564 4344
rect 1811 4384 1822 4386
rect 2035 4392 2042 4447
rect 2195 4392 2202 4447
rect 2355 4453 2363 4502
rect 2456 4498 2474 4500
rect 2456 4489 2486 4498
rect 2578 4556 2590 4562
rect 2751 4556 2763 4562
rect 2831 4556 2843 4562
rect 2871 4556 2883 4562
rect 3010 4556 3022 4562
rect 3150 4556 3162 4562
rect 2626 4498 2644 4500
rect 2614 4489 2644 4498
rect 2456 4461 2464 4489
rect 2636 4461 2644 4489
rect 2736 4481 2744 4536
rect 2853 4493 2860 4536
rect 2956 4498 2974 4500
rect 2956 4489 2986 4498
rect 3096 4498 3114 4500
rect 3096 4489 3126 4498
rect 3217 4556 3229 4562
rect 3337 4556 3349 4562
rect 3501 4556 3513 4562
rect 3619 4556 3631 4562
rect 3771 4556 3783 4562
rect 3815 4556 3823 4562
rect 2035 4386 2082 4392
rect 2035 4384 2043 4386
rect 2071 4384 2082 4386
rect 2195 4386 2242 4392
rect 2195 4384 2203 4386
rect 2231 4384 2242 4386
rect 2355 4384 2363 4439
rect 2455 4392 2462 4447
rect 2638 4392 2645 4447
rect 2455 4386 2502 4392
rect 2455 4384 2463 4386
rect 1651 4338 1663 4344
rect 1691 4338 1703 4344
rect 1791 4338 1803 4344
rect 1831 4338 1843 4344
rect 1951 4338 1963 4344
rect 2051 4338 2063 4344
rect 2091 4338 2103 4344
rect 2211 4338 2223 4344
rect 2251 4338 2263 4344
rect 2491 4384 2502 4386
rect 2598 4386 2645 4392
rect 2598 4384 2609 4386
rect 2331 4338 2343 4344
rect 2371 4338 2383 4344
rect 2471 4338 2483 4344
rect 2511 4338 2523 4344
rect 2637 4384 2645 4386
rect 2736 4384 2744 4467
rect 2853 4431 2860 4479
rect 2956 4461 2964 4489
rect 3096 4461 3104 4489
rect 3236 4481 3244 4536
rect 3329 4516 3357 4522
rect 3317 4513 3369 4516
rect 3471 4516 3481 4526
rect 3879 4556 3891 4562
rect 4029 4556 4041 4562
rect 4147 4556 4159 4562
rect 4309 4556 4321 4562
rect 4431 4556 4443 4562
rect 4519 4556 4531 4562
rect 4689 4556 4701 4562
rect 3377 4502 3385 4516
rect 3360 4495 3385 4502
rect 2843 4424 2860 4431
rect 2955 4392 2962 4447
rect 3095 4392 3102 4447
rect 2955 4386 3002 4392
rect 2955 4384 2963 4386
rect 2991 4384 3002 4386
rect 3095 4386 3142 4392
rect 3095 4384 3103 4386
rect 3131 4384 3142 4386
rect 3236 4384 3244 4467
rect 3359 4473 3367 4495
rect 3471 4473 3479 4516
rect 3531 4506 3543 4516
rect 3649 4508 3661 4516
rect 3505 4498 3543 4506
rect 3637 4502 3661 4508
rect 3471 4459 3473 4473
rect 3353 4424 3361 4459
rect 3471 4424 3479 4459
rect 2577 4338 2589 4344
rect 2617 4338 2629 4344
rect 2751 4338 2763 4344
rect 2871 4338 2883 4344
rect 2971 4338 2983 4344
rect 3011 4338 3023 4344
rect 3111 4338 3123 4344
rect 3151 4338 3163 4344
rect 3514 4384 3522 4498
rect 3637 4453 3645 4502
rect 3753 4481 3760 4516
rect 3791 4508 3797 4536
rect 3909 4508 3921 4516
rect 3787 4502 3797 4508
rect 3897 4502 3921 4508
rect 3637 4384 3645 4439
rect 3757 4423 3766 4467
rect 3776 4441 3782 4496
rect 3897 4453 3905 4502
rect 4011 4473 4019 4516
rect 4051 4510 4059 4536
rect 4037 4504 4059 4510
rect 4179 4516 4189 4526
rect 4117 4506 4129 4516
rect 4037 4498 4040 4504
rect 4117 4498 4155 4506
rect 3787 4432 3823 4440
rect 4011 4459 4013 4473
rect 3815 4424 3823 4432
rect 3757 4414 3761 4423
rect 3217 4338 3229 4344
rect 3322 4338 3334 4344
rect 3372 4338 3384 4344
rect 3487 4338 3499 4344
rect 3531 4338 3543 4344
rect 3897 4384 3905 4439
rect 4011 4424 4019 4459
rect 4033 4442 4040 4498
rect 4037 4436 4040 4442
rect 4037 4430 4063 4436
rect 4055 4384 4063 4430
rect 4138 4384 4146 4498
rect 4181 4473 4189 4516
rect 4279 4508 4291 4516
rect 4279 4502 4303 4508
rect 4187 4459 4189 4473
rect 4181 4424 4189 4459
rect 4295 4453 4303 4502
rect 4395 4502 4403 4516
rect 4423 4516 4451 4522
rect 4411 4513 4463 4516
rect 4549 4508 4561 4516
rect 4537 4502 4561 4508
rect 4757 4556 4769 4562
rect 4859 4556 4871 4562
rect 4997 4556 5009 4562
rect 5099 4556 5111 4562
rect 5157 4556 5169 4562
rect 5205 4556 5217 4562
rect 5267 4556 5279 4562
rect 5377 4556 5389 4562
rect 5497 4556 5505 4562
rect 5537 4556 5549 4562
rect 5691 4556 5703 4562
rect 4659 4508 4671 4516
rect 4659 4502 4683 4508
rect 4395 4495 4420 4502
rect 4413 4473 4421 4495
rect 4295 4384 4303 4439
rect 4419 4424 4427 4459
rect 4537 4453 4545 4502
rect 4675 4453 4683 4502
rect 4776 4481 4784 4536
rect 4889 4508 4901 4516
rect 4989 4516 5017 4522
rect 4977 4513 5029 4516
rect 5247 4536 5260 4542
rect 5131 4530 5138 4536
rect 5127 4522 5138 4530
rect 5188 4524 5195 4536
rect 5253 4530 5260 4536
rect 4877 4502 4901 4508
rect 5037 4502 5045 4516
rect 3617 4338 3629 4344
rect 3657 4338 3669 4344
rect 3781 4338 3793 4344
rect 3877 4338 3889 4344
rect 3917 4338 3929 4344
rect 4029 4338 4041 4344
rect 4117 4338 4129 4344
rect 4161 4338 4173 4344
rect 4271 4338 4283 4344
rect 4311 4338 4323 4344
rect 4537 4384 4545 4439
rect 4675 4384 4683 4439
rect 4776 4384 4784 4467
rect 4877 4453 4885 4502
rect 5020 4495 5045 4502
rect 5077 4501 5085 4516
rect 5188 4517 5209 4524
rect 5167 4506 5173 4508
rect 5234 4506 5241 4512
rect 5019 4473 5027 4495
rect 5077 4487 5093 4501
rect 5167 4500 5241 4506
rect 4877 4384 4885 4439
rect 5013 4424 5021 4459
rect 5077 4424 5085 4487
rect 5093 4473 5107 4487
rect 5099 4428 5113 4436
rect 4396 4338 4408 4344
rect 4446 4338 4458 4344
rect 4517 4338 4529 4344
rect 4557 4338 4569 4344
rect 4651 4338 4663 4344
rect 4691 4338 4703 4344
rect 4757 4338 4769 4344
rect 4857 4338 4869 4344
rect 4897 4338 4909 4344
rect 5167 4428 5173 4500
rect 5234 4492 5241 4500
rect 5246 4484 5280 4492
rect 5274 4479 5280 4484
rect 5227 4466 5254 4473
rect 5133 4422 5173 4428
rect 5181 4428 5225 4434
rect 5133 4404 5139 4422
rect 5181 4414 5187 4428
rect 5293 4432 5299 4516
rect 5369 4516 5397 4522
rect 5357 4513 5409 4516
rect 5417 4502 5425 4516
rect 5523 4508 5529 4536
rect 5523 4502 5533 4508
rect 5400 4495 5425 4502
rect 5399 4473 5407 4495
rect 5237 4424 5299 4432
rect 5393 4424 5401 4459
rect 5538 4441 5544 4496
rect 5560 4481 5567 4516
rect 5655 4502 5663 4516
rect 5683 4516 5711 4522
rect 5671 4513 5723 4516
rect 5655 4495 5680 4502
rect 5673 4473 5681 4495
rect 5497 4432 5533 4440
rect 5497 4424 5505 4432
rect 5157 4408 5187 4414
rect 5205 4410 5243 4418
rect 5235 4404 5243 4410
rect 5127 4364 5139 4398
rect 5185 4390 5207 4402
rect 5235 4390 5253 4404
rect 5181 4384 5193 4390
rect 5235 4384 5243 4390
rect 5554 4423 5563 4467
rect 5679 4424 5687 4459
rect 5559 4414 5563 4423
rect 4982 4338 4994 4344
rect 5032 4338 5044 4344
rect 5097 4338 5109 4344
rect 5155 4338 5167 4344
rect 5201 4338 5213 4344
rect 5267 4338 5279 4344
rect 5362 4338 5374 4344
rect 5412 4338 5424 4344
rect 5527 4338 5539 4344
rect 5656 4338 5668 4344
rect 5706 4338 5718 4344
rect -62 4336 5816 4338
rect -62 4324 4 4336
rect -62 4322 5816 4324
rect -62 3858 -2 4322
rect 96 4316 108 4322
rect 146 4316 158 4322
rect 236 4316 248 4322
rect 286 4316 298 4322
rect 411 4316 423 4322
rect 451 4316 463 4322
rect 551 4316 563 4322
rect 591 4316 603 4322
rect 701 4316 713 4322
rect 816 4316 828 4322
rect 866 4316 878 4322
rect 395 4274 403 4276
rect 431 4274 442 4276
rect 395 4268 442 4274
rect 535 4274 543 4276
rect 571 4274 582 4276
rect 535 4268 582 4274
rect 119 4201 127 4236
rect 259 4201 267 4236
rect 395 4213 402 4268
rect 113 4165 121 4187
rect 253 4165 261 4187
rect 535 4213 542 4268
rect 677 4237 681 4246
rect 396 4171 404 4199
rect 536 4171 544 4199
rect 677 4193 686 4237
rect 937 4316 949 4322
rect 1091 4316 1103 4322
rect 1231 4316 1243 4322
rect 1271 4316 1283 4322
rect 735 4228 743 4236
rect 707 4220 743 4228
rect 95 4158 120 4165
rect 235 4158 260 4165
rect 396 4162 426 4171
rect 396 4160 414 4162
rect 95 4144 103 4158
rect 111 4144 163 4147
rect 235 4144 243 4158
rect 123 4138 151 4144
rect 251 4144 303 4147
rect 263 4138 291 4144
rect 536 4162 566 4171
rect 536 4160 554 4162
rect 507 4137 533 4143
rect 673 4144 680 4179
rect 696 4164 702 4219
rect 839 4201 847 4236
rect 833 4165 841 4187
rect 956 4193 964 4276
rect 1111 4242 1123 4244
rect 1083 4236 1123 4242
rect 1215 4274 1223 4276
rect 1351 4316 1363 4322
rect 1391 4316 1403 4322
rect 1471 4316 1483 4322
rect 1511 4316 1523 4322
rect 1631 4316 1643 4322
rect 1731 4316 1743 4322
rect 1771 4316 1783 4322
rect 1871 4316 1883 4322
rect 1911 4316 1923 4322
rect 1251 4274 1262 4276
rect 1215 4268 1262 4274
rect 1054 4201 1062 4236
rect 1215 4213 1222 4268
rect 1375 4221 1383 4276
rect 1495 4221 1503 4276
rect 1715 4274 1723 4276
rect 1751 4274 1762 4276
rect 1715 4268 1762 4274
rect 1855 4274 1863 4276
rect 1977 4316 1989 4322
rect 2017 4316 2029 4322
rect 2117 4316 2129 4322
rect 2157 4316 2169 4322
rect 2311 4316 2323 4322
rect 1891 4274 1902 4276
rect 1855 4268 1902 4274
rect 1998 4274 2009 4276
rect 2037 4274 2045 4276
rect 1998 4268 2045 4274
rect 2138 4274 2149 4276
rect 2177 4274 2185 4276
rect 2138 4268 2185 4274
rect 1603 4229 1620 4236
rect 815 4158 840 4165
rect 707 4152 717 4158
rect 711 4124 717 4152
rect 815 4144 823 4158
rect 831 4144 883 4147
rect 843 4138 871 4144
rect 956 4124 964 4179
rect 1054 4144 1062 4187
rect 1216 4171 1224 4199
rect 1216 4162 1246 4171
rect 1216 4160 1234 4162
rect 1054 4133 1080 4144
rect 1375 4158 1383 4207
rect 1495 4158 1503 4207
rect 1359 4152 1383 4158
rect 1479 4152 1503 4158
rect 1613 4181 1620 4229
rect 1715 4213 1722 4268
rect 1855 4213 1862 4268
rect 2038 4213 2045 4268
rect 2178 4213 2185 4268
rect 2416 4316 2428 4322
rect 2466 4316 2478 4322
rect 2591 4316 2603 4322
rect 2631 4316 2643 4322
rect 2575 4274 2583 4276
rect 2697 4316 2709 4322
rect 2817 4316 2829 4322
rect 2857 4316 2869 4322
rect 2957 4316 2969 4322
rect 2997 4316 3009 4322
rect 3097 4316 3109 4322
rect 3237 4316 3249 4322
rect 3362 4316 3374 4322
rect 3412 4316 3424 4322
rect 2611 4274 2622 4276
rect 2575 4268 2622 4274
rect 2283 4229 2300 4236
rect 1716 4171 1724 4199
rect 1856 4171 1864 4199
rect 2036 4171 2044 4199
rect 2176 4171 2184 4199
rect 1359 4144 1371 4152
rect 1479 4144 1491 4152
rect 1613 4124 1620 4167
rect 1716 4162 1746 4171
rect 1716 4160 1734 4162
rect 131 4098 143 4104
rect 271 4098 283 4104
rect 450 4098 462 4104
rect 590 4098 602 4104
rect 691 4098 703 4104
rect 735 4098 743 4104
rect 851 4098 863 4104
rect 937 4098 949 4104
rect 1058 4098 1070 4104
rect 1108 4098 1120 4104
rect 1270 4098 1282 4104
rect 1389 4098 1401 4104
rect 1509 4098 1521 4104
rect 1856 4162 1886 4171
rect 1856 4160 1874 4162
rect 1591 4098 1603 4104
rect 1631 4098 1643 4104
rect 1770 4098 1782 4104
rect 1910 4098 1922 4104
rect 2014 4162 2044 4171
rect 2026 4160 2044 4162
rect 2154 4162 2184 4171
rect 2166 4160 2184 4162
rect 2293 4181 2300 4229
rect 2439 4201 2447 4236
rect 2575 4213 2582 4268
rect 2293 4124 2300 4167
rect 2433 4165 2441 4187
rect 2576 4171 2584 4199
rect 2716 4193 2724 4276
rect 2838 4274 2849 4276
rect 2877 4274 2885 4276
rect 2838 4268 2885 4274
rect 2878 4213 2885 4268
rect 2977 4221 2985 4276
rect 3077 4242 3089 4244
rect 3077 4236 3117 4242
rect 3217 4242 3229 4244
rect 3217 4236 3257 4242
rect 3517 4316 3529 4322
rect 3617 4316 3629 4322
rect 3657 4316 3669 4322
rect 3757 4316 3769 4322
rect 3797 4316 3809 4322
rect 3911 4316 3923 4322
rect 3951 4316 3963 4322
rect 2415 4158 2440 4165
rect 2576 4162 2606 4171
rect 2576 4160 2594 4162
rect 2415 4144 2423 4158
rect 2431 4144 2483 4147
rect 2443 4138 2471 4144
rect 2716 4124 2724 4179
rect 2876 4171 2884 4199
rect 1978 4098 1990 4104
rect 2118 4098 2130 4104
rect 2271 4098 2283 4104
rect 2311 4098 2323 4104
rect 2451 4098 2463 4104
rect 2630 4098 2642 4104
rect 2854 4162 2884 4171
rect 2866 4160 2884 4162
rect 2977 4158 2985 4207
rect 3138 4201 3146 4236
rect 3278 4201 3286 4236
rect 3393 4201 3401 4236
rect 2977 4152 3001 4158
rect 2989 4144 3001 4152
rect 3138 4144 3146 4187
rect 3278 4144 3286 4187
rect 3536 4193 3544 4276
rect 3638 4274 3649 4276
rect 3677 4274 3685 4276
rect 3638 4268 3685 4274
rect 3778 4274 3789 4276
rect 4051 4316 4063 4322
rect 4091 4316 4103 4322
rect 4171 4316 4183 4322
rect 4211 4316 4223 4322
rect 4296 4316 4308 4322
rect 4346 4316 4358 4322
rect 4447 4316 4459 4322
rect 4576 4316 4588 4322
rect 4626 4316 4638 4322
rect 3817 4274 3825 4276
rect 3778 4268 3825 4274
rect 3678 4213 3685 4268
rect 3818 4213 3825 4268
rect 3935 4221 3943 4276
rect 4075 4221 4083 4276
rect 4195 4221 4203 4276
rect 4479 4237 4483 4246
rect 3399 4165 3407 4187
rect 3400 4158 3425 4165
rect 3120 4133 3146 4144
rect 2697 4098 2709 4104
rect 2818 4098 2830 4104
rect 2959 4098 2971 4104
rect 3080 4098 3092 4104
rect 3130 4098 3142 4104
rect 3260 4133 3286 4144
rect 3357 4144 3409 4147
rect 3369 4138 3397 4144
rect 3417 4144 3425 4158
rect 3536 4124 3544 4179
rect 3676 4171 3684 4199
rect 3816 4171 3824 4199
rect 3654 4162 3684 4171
rect 3666 4160 3684 4162
rect 3794 4162 3824 4171
rect 3806 4160 3824 4162
rect 3935 4158 3943 4207
rect 4075 4158 4083 4207
rect 4195 4158 4203 4207
rect 4319 4201 4327 4236
rect 4417 4228 4425 4236
rect 4417 4220 4453 4228
rect 4313 4165 4321 4187
rect 3919 4152 3943 4158
rect 4059 4152 4083 4158
rect 4179 4152 4203 4158
rect 4295 4158 4320 4165
rect 4458 4164 4464 4219
rect 4474 4193 4483 4237
rect 4722 4316 4734 4322
rect 4772 4316 4784 4322
rect 4857 4316 4869 4322
rect 4977 4316 4989 4322
rect 5117 4316 5129 4322
rect 5242 4316 5254 4322
rect 5292 4316 5304 4322
rect 4599 4201 4607 4236
rect 4753 4201 4761 4236
rect 4880 4229 4897 4236
rect 3919 4144 3931 4152
rect 4059 4144 4071 4152
rect 4179 4144 4191 4152
rect 4295 4144 4303 4158
rect 4443 4152 4453 4158
rect 4311 4144 4363 4147
rect 4323 4138 4351 4144
rect 4443 4124 4449 4152
rect 4480 4144 4487 4179
rect 4593 4165 4601 4187
rect 4759 4165 4767 4187
rect 4880 4181 4887 4229
rect 4996 4193 5004 4276
rect 5097 4242 5109 4244
rect 5097 4236 5137 4242
rect 5377 4316 5389 4322
rect 5482 4316 5494 4322
rect 5532 4316 5544 4322
rect 5601 4316 5613 4322
rect 5667 4316 5679 4322
rect 5713 4316 5725 4322
rect 5771 4316 5783 4322
rect 5067 4217 5133 4223
rect 5158 4201 5166 4236
rect 5273 4201 5281 4236
rect 4575 4158 4600 4165
rect 4760 4158 4785 4165
rect 4575 4144 4583 4158
rect 4591 4144 4643 4147
rect 4603 4138 4631 4144
rect 4717 4144 4769 4147
rect 4729 4138 4757 4144
rect 4777 4144 4785 4158
rect 4880 4124 4887 4167
rect 4996 4124 5004 4179
rect 5158 4144 5166 4187
rect 5396 4193 5404 4276
rect 5637 4270 5645 4276
rect 5687 4270 5699 4276
rect 5627 4256 5645 4270
rect 5673 4258 5695 4270
rect 5741 4262 5753 4296
rect 5637 4250 5645 4256
rect 5637 4242 5675 4250
rect 5693 4246 5723 4252
rect 5513 4201 5521 4236
rect 5581 4228 5643 4236
rect 5279 4165 5287 4187
rect 5280 4158 5305 4165
rect 3220 4098 3232 4104
rect 3270 4098 3282 4104
rect 3377 4098 3389 4104
rect 3517 4098 3529 4104
rect 3618 4098 3630 4104
rect 3758 4098 3770 4104
rect 3949 4098 3961 4104
rect 4089 4098 4101 4104
rect 4209 4098 4221 4104
rect 4331 4098 4343 4104
rect 4417 4098 4425 4104
rect 4457 4098 4469 4104
rect 4611 4098 4623 4104
rect 4737 4098 4749 4104
rect 4857 4098 4869 4104
rect 4897 4098 4909 4104
rect 5140 4133 5166 4144
rect 5237 4144 5289 4147
rect 5249 4138 5277 4144
rect 5297 4144 5305 4158
rect 5396 4124 5404 4179
rect 5519 4165 5527 4187
rect 5520 4158 5545 4165
rect 5477 4144 5529 4147
rect 5489 4138 5517 4144
rect 5537 4144 5545 4158
rect 5581 4144 5587 4228
rect 5693 4232 5699 4246
rect 5741 4238 5747 4256
rect 5655 4226 5699 4232
rect 5707 4232 5747 4238
rect 5626 4187 5653 4194
rect 5600 4176 5606 4181
rect 5600 4168 5634 4176
rect 5639 4160 5646 4168
rect 5707 4160 5713 4232
rect 5767 4224 5781 4232
rect 5773 4173 5787 4187
rect 5795 4173 5803 4236
rect 5639 4154 5713 4160
rect 5787 4159 5803 4173
rect 5639 4148 5646 4154
rect 5707 4152 5713 4154
rect 5671 4136 5692 4143
rect 5795 4144 5803 4159
rect 5620 4124 5627 4130
rect 5685 4124 5692 4136
rect 5742 4130 5753 4138
rect 5742 4124 5749 4130
rect 5620 4118 5633 4124
rect 4977 4098 4989 4104
rect 5100 4098 5112 4104
rect 5150 4098 5162 4104
rect 5257 4098 5269 4104
rect 5377 4098 5389 4104
rect 5497 4098 5509 4104
rect 5601 4098 5613 4104
rect 5663 4098 5675 4104
rect 5711 4098 5723 4104
rect 5769 4098 5781 4104
rect 5822 4098 5882 4562
rect 4 4096 5882 4098
rect 5816 4084 5882 4096
rect 4 4082 5882 4084
rect 91 4076 103 4082
rect 197 4076 209 4082
rect 351 4076 363 4082
rect 76 4001 84 4056
rect 189 4036 217 4042
rect 177 4033 229 4036
rect 440 4076 452 4082
rect 490 4076 502 4082
rect 237 4022 245 4036
rect 220 4015 245 4022
rect 76 3904 84 3987
rect 107 3937 133 3943
rect 157 3923 163 4013
rect 219 3993 227 4015
rect 336 4001 344 4056
rect 591 4076 603 4082
rect 631 4076 643 4082
rect 751 4076 763 4082
rect 837 4076 849 4082
rect 957 4076 969 4082
rect 1058 4076 1070 4082
rect 1200 4076 1212 4082
rect 1256 4076 1268 4082
rect 480 4036 506 4047
rect 498 3993 506 4036
rect 613 4013 620 4056
rect 736 4001 744 4056
rect 829 4036 857 4042
rect 817 4033 869 4036
rect 877 4022 885 4036
rect 860 4015 885 4022
rect 213 3944 221 3979
rect 107 3917 163 3923
rect 91 3858 103 3864
rect 336 3904 344 3987
rect 498 3944 506 3979
rect 613 3951 620 3999
rect 603 3944 620 3951
rect 437 3938 477 3944
rect 437 3936 449 3938
rect 736 3904 744 3987
rect 859 3993 867 4015
rect 976 4001 984 4056
rect 1379 4076 1391 4082
rect 1531 4076 1543 4082
rect 1611 4076 1623 4082
rect 1651 4076 1663 4082
rect 1751 4076 1763 4082
rect 1818 4076 1830 4082
rect 2011 4076 2023 4082
rect 2190 4076 2202 4082
rect 1106 4018 1124 4020
rect 1094 4009 1124 4018
rect 853 3944 861 3979
rect 182 3858 194 3864
rect 232 3858 244 3864
rect 351 3858 363 3864
rect 457 3858 469 3864
rect 631 3858 643 3864
rect 751 3858 763 3864
rect 976 3904 984 3987
rect 1116 3981 1124 4009
rect 1233 3993 1240 4036
rect 1409 4028 1421 4036
rect 1397 4022 1421 4028
rect 1118 3912 1125 3967
rect 1241 3956 1247 3979
rect 1397 3973 1405 4022
rect 1516 4001 1524 4056
rect 1633 4013 1640 4056
rect 1667 4037 1693 4043
rect 1736 4001 1744 4056
rect 1975 4022 1983 4036
rect 2003 4036 2031 4042
rect 1991 4033 2043 4036
rect 1866 4018 1884 4020
rect 1241 3950 1268 3956
rect 1256 3944 1268 3950
rect 1078 3906 1125 3912
rect 1078 3904 1089 3906
rect 822 3858 834 3864
rect 872 3858 884 3864
rect 1117 3904 1125 3906
rect 1209 3936 1237 3942
rect 1249 3864 1277 3870
rect 1397 3904 1405 3959
rect 1516 3904 1524 3987
rect 1633 3951 1640 3999
rect 1854 4009 1884 4018
rect 1975 4015 2000 4022
rect 2136 4018 2154 4020
rect 1623 3944 1640 3951
rect 1736 3904 1744 3987
rect 1876 3981 1884 4009
rect 1993 3993 2001 4015
rect 2136 4009 2166 4018
rect 2258 4076 2270 4082
rect 2451 4076 2463 4082
rect 2589 4076 2601 4082
rect 2415 4022 2423 4036
rect 2443 4036 2471 4042
rect 2431 4033 2483 4036
rect 2659 4076 2671 4082
rect 2778 4076 2790 4082
rect 2918 4076 2930 4082
rect 3091 4076 3103 4082
rect 3230 4076 3242 4082
rect 3331 4076 3343 4082
rect 3451 4076 3463 4082
rect 3539 4076 3551 4082
rect 3691 4076 3703 4082
rect 3735 4076 3743 4082
rect 2559 4028 2571 4036
rect 2689 4028 2701 4036
rect 2559 4022 2583 4028
rect 2306 4018 2324 4020
rect 2294 4009 2324 4018
rect 2415 4015 2440 4022
rect 2136 3981 2144 4009
rect 2316 3981 2324 4009
rect 2433 3993 2441 4015
rect 1878 3912 1885 3967
rect 1999 3944 2007 3979
rect 1838 3906 1885 3912
rect 1838 3904 1849 3906
rect 957 3858 969 3864
rect 1057 3858 1069 3864
rect 1097 3858 1109 3864
rect 1217 3858 1229 3864
rect 1377 3858 1389 3864
rect 1417 3858 1429 3864
rect 1531 3858 1543 3864
rect 1651 3858 1663 3864
rect 1751 3858 1763 3864
rect 1877 3904 1885 3906
rect 2135 3912 2142 3967
rect 2318 3912 2325 3967
rect 2439 3944 2447 3979
rect 2575 3973 2583 4022
rect 2607 4017 2623 4023
rect 2617 3967 2623 4017
rect 2677 4022 2701 4028
rect 2135 3906 2182 3912
rect 2135 3904 2143 3906
rect 2171 3904 2182 3906
rect 2278 3906 2325 3912
rect 2278 3904 2289 3906
rect 1817 3858 1829 3864
rect 1857 3858 1869 3864
rect 1976 3858 1988 3864
rect 2026 3858 2038 3864
rect 2151 3858 2163 3864
rect 2191 3858 2203 3864
rect 2317 3904 2325 3906
rect 2575 3904 2583 3959
rect 2637 3943 2643 3973
rect 2677 3973 2685 4022
rect 2826 4018 2844 4020
rect 2814 4009 2844 4018
rect 2966 4018 2984 4020
rect 2954 4009 2984 4018
rect 2836 3981 2844 4009
rect 2976 3981 2984 4009
rect 3076 4001 3084 4056
rect 3176 4018 3194 4020
rect 3176 4009 3206 4018
rect 2607 3937 2643 3943
rect 2677 3904 2685 3959
rect 2838 3912 2845 3967
rect 2978 3912 2985 3967
rect 2798 3906 2845 3912
rect 2798 3904 2809 3906
rect 2257 3858 2269 3864
rect 2297 3858 2309 3864
rect 2416 3858 2428 3864
rect 2466 3858 2478 3864
rect 2551 3858 2563 3864
rect 2591 3858 2603 3864
rect 2657 3858 2669 3864
rect 2697 3858 2709 3864
rect 2837 3904 2845 3906
rect 2938 3906 2985 3912
rect 2938 3904 2949 3906
rect 2977 3904 2985 3906
rect 3076 3904 3084 3987
rect 3176 3981 3184 4009
rect 3316 4001 3324 4056
rect 3415 4022 3423 4036
rect 3443 4036 3471 4042
rect 3819 4076 3831 4082
rect 3991 4076 4003 4082
rect 4098 4076 4110 4082
rect 4148 4076 4160 4082
rect 3431 4033 3483 4036
rect 3569 4028 3581 4036
rect 3557 4022 3581 4028
rect 3415 4015 3440 4022
rect 3433 3993 3441 4015
rect 3175 3912 3182 3967
rect 3175 3906 3222 3912
rect 3175 3904 3183 3906
rect 3211 3904 3222 3906
rect 3316 3904 3324 3987
rect 3439 3944 3447 3979
rect 3557 3973 3565 4022
rect 3673 4001 3680 4036
rect 3711 4028 3717 4056
rect 3849 4028 3861 4036
rect 3707 4022 3717 4028
rect 3837 4022 3861 4028
rect 3955 4022 3963 4036
rect 3983 4036 4011 4042
rect 3971 4033 4023 4036
rect 4094 4036 4120 4047
rect 4219 4076 4231 4082
rect 4357 4076 4369 4082
rect 4497 4076 4509 4082
rect 4617 4076 4625 4082
rect 4657 4076 4669 4082
rect 4809 4076 4821 4082
rect 2777 3858 2789 3864
rect 2817 3858 2829 3864
rect 2917 3858 2929 3864
rect 2957 3858 2969 3864
rect 3091 3858 3103 3864
rect 3191 3858 3203 3864
rect 3231 3858 3243 3864
rect 3331 3858 3343 3864
rect 3557 3904 3565 3959
rect 3677 3943 3686 3987
rect 3696 3961 3702 4016
rect 3837 3973 3845 4022
rect 3955 4015 3980 4022
rect 3973 3993 3981 4015
rect 3707 3952 3743 3960
rect 4094 3993 4102 4036
rect 4249 4028 4261 4036
rect 4349 4036 4377 4042
rect 4337 4033 4389 4036
rect 4489 4036 4517 4042
rect 4237 4022 4261 4028
rect 4397 4022 4405 4036
rect 4477 4033 4529 4036
rect 4537 4022 4545 4036
rect 4643 4028 4649 4056
rect 4878 4076 4890 4082
rect 5017 4076 5029 4082
rect 5151 4076 5163 4082
rect 5199 4076 5211 4082
rect 5257 4076 5269 4082
rect 5305 4076 5317 4082
rect 5367 4076 5379 4082
rect 5439 4076 5451 4082
rect 5497 4076 5509 4082
rect 5545 4076 5557 4082
rect 5607 4076 5619 4082
rect 5717 4076 5729 4082
rect 4643 4022 4653 4028
rect 3735 3944 3743 3952
rect 3677 3934 3681 3943
rect 3416 3858 3428 3864
rect 3466 3858 3478 3864
rect 3837 3904 3845 3959
rect 3979 3944 3987 3979
rect 4094 3944 4102 3979
rect 4237 3973 4245 4022
rect 4380 4015 4405 4022
rect 4520 4015 4545 4022
rect 4379 3993 4387 4015
rect 4519 3993 4527 4015
rect 3537 3858 3549 3864
rect 3577 3858 3589 3864
rect 3701 3858 3713 3864
rect 3817 3858 3829 3864
rect 3857 3858 3869 3864
rect 4123 3938 4163 3944
rect 4151 3936 4163 3938
rect 4237 3904 4245 3959
rect 4373 3944 4381 3979
rect 4513 3944 4521 3979
rect 4658 3961 4664 4016
rect 4680 4001 4687 4036
rect 4779 4028 4791 4036
rect 4779 4022 4803 4028
rect 4617 3952 4653 3960
rect 4617 3944 4625 3952
rect 3956 3858 3968 3864
rect 4006 3858 4018 3864
rect 4131 3858 4143 3864
rect 4217 3858 4229 3864
rect 4257 3858 4269 3864
rect 4342 3858 4354 3864
rect 4392 3858 4404 3864
rect 4674 3943 4683 3987
rect 4795 3973 4803 4022
rect 4926 4018 4944 4020
rect 4914 4009 4944 4018
rect 4936 3981 4944 4009
rect 5036 4001 5044 4056
rect 5136 4001 5144 4056
rect 5347 4056 5360 4062
rect 5231 4050 5238 4056
rect 5227 4042 5238 4050
rect 5288 4044 5295 4056
rect 5353 4050 5360 4056
rect 5177 4021 5185 4036
rect 5288 4037 5309 4044
rect 5267 4026 5273 4028
rect 5334 4026 5341 4032
rect 5177 4007 5193 4021
rect 5267 4020 5341 4026
rect 4679 3934 4683 3943
rect 4795 3904 4803 3959
rect 4938 3912 4945 3967
rect 4898 3906 4945 3912
rect 4898 3904 4909 3906
rect 4482 3858 4494 3864
rect 4532 3858 4544 3864
rect 4647 3858 4659 3864
rect 4771 3858 4783 3864
rect 4811 3858 4823 3864
rect 4937 3904 4945 3906
rect 5036 3904 5044 3987
rect 5136 3904 5144 3987
rect 5177 3944 5185 4007
rect 5193 3993 5207 4007
rect 5199 3948 5213 3956
rect 5267 3948 5273 4020
rect 5334 4012 5341 4020
rect 5346 4004 5380 4012
rect 5374 3999 5380 4004
rect 5327 3986 5354 3993
rect 5233 3942 5273 3948
rect 5281 3948 5325 3954
rect 5233 3924 5239 3942
rect 5281 3934 5287 3948
rect 5393 3952 5399 4036
rect 5337 3944 5399 3952
rect 5257 3928 5287 3934
rect 5305 3930 5343 3938
rect 5335 3924 5343 3930
rect 5227 3884 5239 3918
rect 5285 3910 5307 3922
rect 5335 3910 5353 3924
rect 5281 3904 5293 3910
rect 5335 3904 5343 3910
rect 5587 4056 5600 4062
rect 5471 4050 5478 4056
rect 5467 4042 5478 4050
rect 5528 4044 5535 4056
rect 5593 4050 5600 4056
rect 5417 4021 5425 4036
rect 5528 4037 5549 4044
rect 5507 4026 5513 4028
rect 5574 4026 5581 4032
rect 5417 4007 5433 4021
rect 5507 4020 5581 4026
rect 5417 3944 5425 4007
rect 5433 3993 5447 4007
rect 5439 3948 5453 3956
rect 5507 3948 5513 4020
rect 5574 4012 5581 4020
rect 5586 4004 5620 4012
rect 5614 3999 5620 4004
rect 5567 3986 5594 3993
rect 5473 3942 5513 3948
rect 5521 3948 5565 3954
rect 5473 3924 5479 3942
rect 5521 3934 5527 3948
rect 5633 3952 5639 4036
rect 5709 4036 5737 4042
rect 5697 4033 5749 4036
rect 5757 4022 5765 4036
rect 5740 4015 5765 4022
rect 5739 3993 5747 4015
rect 5577 3944 5639 3952
rect 5733 3944 5741 3979
rect 5497 3928 5527 3934
rect 5545 3930 5583 3938
rect 5575 3924 5583 3930
rect 5467 3884 5479 3918
rect 5525 3910 5547 3922
rect 5575 3910 5593 3924
rect 5521 3904 5533 3910
rect 5575 3904 5583 3910
rect 4877 3858 4889 3864
rect 4917 3858 4929 3864
rect 5017 3858 5029 3864
rect 5151 3858 5163 3864
rect 5197 3858 5209 3864
rect 5255 3858 5267 3864
rect 5301 3858 5313 3864
rect 5367 3858 5379 3864
rect 5437 3858 5449 3864
rect 5495 3858 5507 3864
rect 5541 3858 5553 3864
rect 5607 3858 5619 3864
rect 5702 3858 5714 3864
rect 5752 3858 5764 3864
rect -62 3856 5816 3858
rect -62 3844 4 3856
rect -62 3842 5816 3844
rect -62 3378 -2 3842
rect 71 3836 83 3842
rect 111 3836 123 3842
rect 211 3836 223 3842
rect 251 3836 263 3842
rect 451 3836 463 3842
rect 556 3836 568 3842
rect 606 3836 618 3842
rect 95 3741 103 3796
rect 195 3794 203 3796
rect 327 3830 379 3836
rect 327 3828 339 3830
rect 231 3794 242 3796
rect 195 3788 242 3794
rect 195 3733 202 3788
rect 367 3828 379 3830
rect 351 3756 359 3772
rect 403 3830 431 3836
rect 411 3772 423 3776
rect 379 3768 423 3772
rect 367 3766 423 3768
rect 431 3770 443 3776
rect 471 3770 483 3776
rect 431 3764 483 3770
rect 691 3836 703 3842
rect 731 3836 743 3842
rect 802 3836 814 3842
rect 852 3836 864 3842
rect 1031 3836 1043 3842
rect 1117 3836 1129 3842
rect 1157 3836 1169 3842
rect 351 3748 374 3756
rect 95 3678 103 3727
rect 196 3691 204 3719
rect 366 3713 374 3748
rect 579 3721 587 3756
rect 715 3741 723 3796
rect 983 3830 1011 3836
rect 1023 3758 1051 3764
rect 1237 3836 1249 3842
rect 1277 3836 1289 3842
rect 1397 3836 1409 3842
rect 1522 3836 1534 3842
rect 1572 3836 1584 3842
rect 367 3699 374 3713
rect 196 3682 226 3691
rect 196 3680 214 3682
rect 79 3672 103 3678
rect 79 3664 91 3672
rect 366 3656 374 3699
rect 573 3685 581 3707
rect 555 3678 580 3685
rect 715 3678 723 3727
rect 833 3721 841 3756
rect 992 3750 1004 3756
rect 992 3744 1019 3750
rect 1013 3721 1019 3744
rect 1137 3741 1145 3796
rect 1258 3794 1269 3796
rect 1297 3794 1305 3796
rect 1258 3788 1305 3794
rect 839 3685 847 3707
rect 840 3678 865 3685
rect 555 3664 563 3678
rect 699 3672 723 3678
rect 366 3650 438 3656
rect 391 3644 398 3650
rect 431 3644 438 3650
rect 571 3664 623 3667
rect 583 3658 611 3664
rect 699 3664 711 3672
rect 797 3664 849 3667
rect 809 3658 837 3664
rect 857 3664 865 3678
rect 1020 3664 1027 3707
rect 1137 3678 1145 3727
rect 1298 3733 1305 3788
rect 1377 3762 1389 3764
rect 1377 3756 1417 3762
rect 1657 3836 1669 3842
rect 1771 3836 1783 3842
rect 1811 3836 1823 3842
rect 1877 3836 1889 3842
rect 1917 3836 1929 3842
rect 2027 3836 2039 3842
rect 2137 3836 2149 3842
rect 2177 3836 2189 3842
rect 1367 3737 1413 3743
rect 1438 3721 1446 3756
rect 1553 3721 1561 3756
rect 1296 3691 1304 3719
rect 1137 3672 1161 3678
rect 1149 3664 1161 3672
rect 109 3618 121 3624
rect 250 3618 262 3624
rect 411 3618 423 3624
rect 451 3618 465 3624
rect 591 3618 603 3624
rect 729 3618 741 3624
rect 817 3618 829 3624
rect 992 3618 1004 3624
rect 1048 3618 1060 3624
rect 1274 3682 1304 3691
rect 1286 3680 1304 3682
rect 1438 3664 1446 3707
rect 1676 3713 1684 3796
rect 1795 3741 1803 3796
rect 1897 3741 1905 3796
rect 2257 3836 2269 3842
rect 2297 3836 2309 3842
rect 2416 3836 2428 3842
rect 2466 3836 2478 3842
rect 2059 3757 2063 3766
rect 1997 3748 2005 3756
rect 1559 3685 1567 3707
rect 1560 3678 1585 3685
rect 1420 3653 1446 3664
rect 1517 3664 1569 3667
rect 1529 3658 1557 3664
rect 1577 3664 1585 3678
rect 1676 3644 1684 3699
rect 1795 3678 1803 3727
rect 1997 3740 2033 3748
rect 1779 3672 1803 3678
rect 1897 3678 1905 3727
rect 2038 3684 2044 3739
rect 2054 3713 2063 3757
rect 2157 3741 2165 3796
rect 2278 3794 2289 3796
rect 2317 3794 2325 3796
rect 2278 3788 2325 3794
rect 1897 3672 1921 3678
rect 1779 3664 1791 3672
rect 1909 3664 1921 3672
rect 1119 3618 1131 3624
rect 1238 3618 1250 3624
rect 1380 3618 1392 3624
rect 1430 3618 1442 3624
rect 1537 3618 1549 3624
rect 1657 3618 1669 3624
rect 1809 3618 1821 3624
rect 2023 3672 2033 3678
rect 2023 3644 2029 3672
rect 2060 3664 2067 3699
rect 2157 3678 2165 3727
rect 2318 3733 2325 3788
rect 2537 3836 2549 3842
rect 2577 3836 2589 3842
rect 2662 3836 2674 3842
rect 2712 3836 2724 3842
rect 2831 3836 2843 3842
rect 2439 3721 2447 3756
rect 2557 3741 2565 3796
rect 2916 3836 2928 3842
rect 2966 3836 2978 3842
rect 2316 3691 2324 3719
rect 2157 3672 2181 3678
rect 2169 3664 2181 3672
rect 2294 3682 2324 3691
rect 2433 3685 2441 3707
rect 2306 3680 2324 3682
rect 2415 3678 2440 3685
rect 2557 3678 2565 3727
rect 2693 3721 2701 3756
rect 2816 3713 2824 3796
rect 3037 3836 3049 3842
rect 3077 3836 3089 3842
rect 3191 3836 3203 3842
rect 3231 3836 3243 3842
rect 3331 3836 3343 3842
rect 3397 3836 3409 3842
rect 3437 3836 3449 3842
rect 3537 3836 3549 3842
rect 3691 3836 3703 3842
rect 2939 3721 2947 3756
rect 3057 3741 3065 3796
rect 3087 3757 3193 3763
rect 3215 3741 3223 3796
rect 2699 3685 2707 3707
rect 2700 3678 2725 3685
rect 2415 3664 2423 3678
rect 2557 3672 2581 3678
rect 2431 3664 2483 3667
rect 2569 3664 2581 3672
rect 2443 3658 2471 3664
rect 2657 3664 2709 3667
rect 2669 3658 2697 3664
rect 2717 3664 2725 3678
rect 2816 3644 2824 3699
rect 2933 3685 2941 3707
rect 2915 3678 2940 3685
rect 3057 3678 3065 3727
rect 3215 3678 3223 3727
rect 3316 3713 3324 3796
rect 3418 3794 3429 3796
rect 3457 3794 3465 3796
rect 3418 3788 3465 3794
rect 3367 3777 3393 3783
rect 3458 3733 3465 3788
rect 2915 3664 2923 3678
rect 3057 3672 3081 3678
rect 2931 3664 2983 3667
rect 3069 3664 3081 3672
rect 2943 3658 2971 3664
rect 3199 3672 3223 3678
rect 3199 3664 3211 3672
rect 3316 3644 3324 3699
rect 3456 3691 3464 3719
rect 3556 3713 3564 3796
rect 3777 3836 3789 3842
rect 3817 3836 3829 3842
rect 3897 3836 3909 3842
rect 4031 3836 4043 3842
rect 4077 3836 4089 3842
rect 4135 3836 4147 3842
rect 4181 3836 4193 3842
rect 4247 3836 4259 3842
rect 4361 3836 4373 3842
rect 4431 3836 4443 3842
rect 3663 3749 3680 3756
rect 1879 3618 1891 3624
rect 1997 3618 2005 3624
rect 2037 3618 2049 3624
rect 2139 3618 2151 3624
rect 2258 3618 2270 3624
rect 2451 3618 2463 3624
rect 2539 3618 2551 3624
rect 2677 3618 2689 3624
rect 2831 3618 2843 3624
rect 2951 3618 2963 3624
rect 3039 3618 3051 3624
rect 3229 3618 3241 3624
rect 3331 3618 3343 3624
rect 3434 3682 3464 3691
rect 3673 3701 3680 3749
rect 3797 3741 3805 3796
rect 3446 3680 3464 3682
rect 3556 3644 3564 3699
rect 3673 3644 3680 3687
rect 3797 3678 3805 3727
rect 3916 3713 3924 3796
rect 4016 3713 4024 3796
rect 4107 3782 4119 3816
rect 4161 3790 4173 3796
rect 4215 3790 4223 3796
rect 4165 3778 4187 3790
rect 4215 3776 4233 3790
rect 4113 3758 4119 3776
rect 4137 3766 4167 3772
rect 4215 3770 4223 3776
rect 3797 3672 3821 3678
rect 3809 3664 3821 3672
rect 3398 3618 3410 3624
rect 3537 3618 3549 3624
rect 3651 3618 3663 3624
rect 3691 3618 3703 3624
rect 3916 3644 3924 3699
rect 4016 3644 4024 3699
rect 4057 3693 4065 3756
rect 4079 3744 4093 3752
rect 4113 3752 4153 3758
rect 4073 3693 4087 3707
rect 4057 3679 4073 3693
rect 4147 3680 4153 3752
rect 4161 3752 4167 3766
rect 4185 3762 4223 3770
rect 4497 3836 4509 3842
rect 4537 3836 4549 3842
rect 4617 3836 4629 3842
rect 4742 3836 4754 3842
rect 4792 3836 4804 3842
rect 4161 3746 4205 3752
rect 4217 3748 4279 3756
rect 4207 3707 4234 3714
rect 4254 3696 4260 3701
rect 4226 3688 4260 3696
rect 4214 3680 4221 3688
rect 4057 3664 4065 3679
rect 4147 3674 4221 3680
rect 4147 3672 4153 3674
rect 4214 3668 4221 3674
rect 4107 3650 4118 3658
rect 4111 3644 4118 3650
rect 4168 3656 4189 3663
rect 4273 3664 4279 3748
rect 4395 3721 4403 3756
rect 4517 3741 4525 3796
rect 4877 3836 4889 3842
rect 5011 3836 5023 3842
rect 5051 3836 5063 3842
rect 5117 3836 5129 3842
rect 5231 3836 5243 3842
rect 5271 3836 5283 3842
rect 5311 3836 5323 3842
rect 5351 3836 5363 3842
rect 5391 3836 5403 3842
rect 5437 3836 5449 3842
rect 5495 3836 5507 3842
rect 5541 3836 5553 3842
rect 5607 3836 5619 3842
rect 5711 3836 5723 3842
rect 5751 3836 5763 3842
rect 4640 3749 4657 3756
rect 4396 3681 4404 3707
rect 4375 3674 4404 3681
rect 4517 3678 4525 3727
rect 4640 3701 4647 3749
rect 4773 3721 4781 3756
rect 4847 3737 4873 3743
rect 4896 3721 4904 3756
rect 5035 3741 5043 3796
rect 4375 3664 4381 3674
rect 4517 3672 4541 3678
rect 4391 3664 4443 3666
rect 4529 3664 4541 3672
rect 4168 3644 4175 3656
rect 4233 3644 4240 3650
rect 4227 3638 4240 3644
rect 4363 3624 4391 3630
rect 4403 3660 4431 3664
rect 4640 3644 4647 3687
rect 4779 3685 4787 3707
rect 4780 3678 4805 3685
rect 4737 3664 4789 3667
rect 4749 3658 4777 3664
rect 4797 3664 4805 3678
rect 4896 3664 4904 3707
rect 5035 3678 5043 3727
rect 5136 3713 5144 3796
rect 5467 3782 5479 3816
rect 5521 3790 5533 3796
rect 5575 3790 5583 3796
rect 5525 3778 5547 3790
rect 5575 3776 5593 3790
rect 5473 3758 5479 3776
rect 5497 3766 5527 3772
rect 5575 3770 5583 3776
rect 5251 3750 5263 3756
rect 5291 3750 5303 3756
rect 5331 3750 5343 3756
rect 5371 3750 5383 3756
rect 5245 3742 5263 3750
rect 5278 3742 5303 3750
rect 5318 3742 5343 3750
rect 5357 3742 5383 3750
rect 5245 3713 5252 3742
rect 5247 3699 5252 3713
rect 5019 3672 5043 3678
rect 5019 3664 5031 3672
rect 5136 3644 5144 3699
rect 5245 3678 5252 3699
rect 5278 3696 5286 3742
rect 5318 3696 5326 3742
rect 5357 3696 5365 3742
rect 5270 3684 5286 3696
rect 5310 3684 5326 3696
rect 5350 3684 5365 3696
rect 5417 3693 5425 3756
rect 5439 3744 5453 3752
rect 5473 3752 5513 3758
rect 5433 3693 5447 3707
rect 5278 3678 5286 3684
rect 5318 3678 5326 3684
rect 5357 3678 5365 3684
rect 5417 3679 5433 3693
rect 5507 3680 5513 3752
rect 5521 3752 5527 3766
rect 5545 3762 5583 3770
rect 5521 3746 5565 3752
rect 5577 3748 5639 3756
rect 5567 3707 5594 3714
rect 5614 3696 5620 3701
rect 5586 3688 5620 3696
rect 5574 3680 5581 3688
rect 5245 3671 5264 3678
rect 5246 3670 5264 3671
rect 5278 3670 5304 3678
rect 5318 3670 5343 3678
rect 5357 3670 5384 3678
rect 5252 3664 5264 3670
rect 5292 3664 5304 3670
rect 5331 3664 5343 3670
rect 5372 3664 5384 3670
rect 5417 3664 5425 3679
rect 5507 3674 5581 3680
rect 5507 3672 5513 3674
rect 3779 3618 3791 3624
rect 3897 3618 3909 3624
rect 4031 3618 4043 3624
rect 4079 3618 4091 3624
rect 4137 3618 4149 3624
rect 4185 3618 4197 3624
rect 4247 3618 4259 3624
rect 4411 3618 4423 3624
rect 4499 3618 4511 3624
rect 4617 3618 4629 3624
rect 4657 3618 4669 3624
rect 4757 3618 4769 3624
rect 4877 3618 4889 3624
rect 5049 3618 5061 3624
rect 5574 3668 5581 3674
rect 5467 3650 5478 3658
rect 5471 3644 5478 3650
rect 5528 3656 5549 3663
rect 5633 3664 5639 3748
rect 5735 3741 5743 3796
rect 5735 3678 5743 3727
rect 5528 3644 5535 3656
rect 5593 3644 5600 3650
rect 5587 3638 5600 3644
rect 5719 3672 5743 3678
rect 5719 3664 5731 3672
rect 5117 3618 5129 3624
rect 5231 3618 5243 3624
rect 5271 3618 5283 3624
rect 5311 3618 5323 3624
rect 5351 3618 5363 3624
rect 5391 3618 5403 3624
rect 5439 3618 5451 3624
rect 5497 3618 5509 3624
rect 5545 3618 5557 3624
rect 5607 3618 5619 3624
rect 5749 3618 5761 3624
rect 5822 3618 5882 4082
rect 4 3616 5882 3618
rect 5816 3604 5882 3616
rect 4 3602 5882 3604
rect 111 3596 123 3602
rect 200 3596 212 3602
rect 250 3596 262 3602
rect 75 3542 83 3556
rect 103 3556 131 3562
rect 337 3596 349 3602
rect 457 3596 469 3602
rect 578 3596 590 3602
rect 789 3596 801 3602
rect 909 3596 921 3602
rect 997 3596 1009 3602
rect 1190 3596 1202 3602
rect 240 3556 266 3567
rect 91 3553 143 3556
rect 75 3535 100 3542
rect 57 3517 73 3523
rect 57 3443 63 3517
rect 93 3513 101 3535
rect 258 3513 266 3556
rect 356 3521 364 3576
rect 449 3556 477 3562
rect 437 3553 489 3556
rect 497 3542 505 3556
rect 480 3535 505 3542
rect 989 3556 1017 3562
rect 759 3548 771 3556
rect 879 3548 891 3556
rect 977 3553 1029 3556
rect 759 3542 783 3548
rect 879 3542 903 3548
rect 1037 3542 1045 3556
rect 626 3538 644 3540
rect 99 3464 107 3499
rect 258 3464 266 3499
rect 57 3437 73 3443
rect 197 3458 237 3464
rect 197 3456 209 3458
rect 356 3424 364 3507
rect 479 3513 487 3535
rect 614 3529 644 3538
rect 636 3501 644 3529
rect 473 3464 481 3499
rect 775 3493 783 3542
rect 638 3432 645 3487
rect 895 3493 903 3542
rect 1020 3535 1045 3542
rect 1136 3538 1154 3540
rect 1019 3513 1027 3535
rect 1136 3529 1166 3538
rect 1259 3596 1271 3602
rect 1450 3596 1462 3602
rect 1537 3596 1549 3602
rect 1678 3596 1690 3602
rect 1728 3596 1740 3602
rect 1870 3596 1882 3602
rect 1289 3548 1301 3556
rect 1277 3542 1301 3548
rect 1136 3501 1144 3529
rect 598 3426 645 3432
rect 598 3424 609 3426
rect 76 3378 88 3384
rect 126 3378 138 3384
rect 217 3378 229 3384
rect 337 3378 349 3384
rect 442 3378 454 3384
rect 492 3378 504 3384
rect 637 3424 645 3426
rect 775 3424 783 3479
rect 895 3424 903 3479
rect 1013 3464 1021 3499
rect 577 3378 589 3384
rect 617 3378 629 3384
rect 751 3378 763 3384
rect 791 3378 803 3384
rect 871 3378 883 3384
rect 911 3378 923 3384
rect 1135 3432 1142 3487
rect 1217 3463 1223 3513
rect 1277 3493 1285 3542
rect 1396 3538 1414 3540
rect 1396 3529 1426 3538
rect 1529 3556 1557 3562
rect 1517 3553 1569 3556
rect 1674 3556 1700 3567
rect 1577 3542 1585 3556
rect 1560 3535 1585 3542
rect 1396 3501 1404 3529
rect 1559 3513 1567 3535
rect 1674 3513 1682 3556
rect 1816 3538 1834 3540
rect 1816 3529 1846 3538
rect 1940 3596 1952 3602
rect 1990 3596 2002 3602
rect 2131 3596 2143 3602
rect 2257 3596 2269 3602
rect 2398 3596 2410 3602
rect 2448 3596 2460 3602
rect 2561 3596 2573 3602
rect 2659 3596 2671 3602
rect 2831 3596 2843 3602
rect 2969 3596 2981 3602
rect 3109 3596 3121 3602
rect 1980 3556 2006 3567
rect 1816 3501 1824 3529
rect 1998 3513 2006 3556
rect 2095 3542 2103 3556
rect 2123 3556 2151 3562
rect 2111 3553 2163 3556
rect 2249 3556 2277 3562
rect 2237 3553 2289 3556
rect 2394 3556 2420 3567
rect 2531 3556 2541 3566
rect 2095 3535 2120 3542
rect 2113 3513 2121 3535
rect 2167 3537 2193 3543
rect 2297 3542 2305 3556
rect 2280 3535 2305 3542
rect 1217 3457 1253 3463
rect 1135 3426 1182 3432
rect 1135 3424 1143 3426
rect 1171 3424 1182 3426
rect 1277 3424 1285 3479
rect 1395 3432 1402 3487
rect 1553 3464 1561 3499
rect 1674 3464 1682 3499
rect 2279 3513 2287 3535
rect 2394 3513 2402 3556
rect 2531 3513 2539 3556
rect 2591 3546 2603 3556
rect 2689 3548 2701 3556
rect 2565 3538 2603 3546
rect 2677 3542 2701 3548
rect 2795 3542 2803 3556
rect 2823 3556 2851 3562
rect 2811 3553 2863 3556
rect 2531 3499 2533 3513
rect 1395 3426 1442 3432
rect 1395 3424 1403 3426
rect 982 3378 994 3384
rect 1032 3378 1044 3384
rect 1151 3378 1163 3384
rect 1191 3378 1203 3384
rect 1431 3424 1442 3426
rect 1257 3378 1269 3384
rect 1297 3378 1309 3384
rect 1411 3378 1423 3384
rect 1451 3378 1463 3384
rect 1703 3458 1743 3464
rect 1731 3456 1743 3458
rect 1815 3432 1822 3487
rect 1998 3464 2006 3499
rect 2119 3464 2127 3499
rect 2273 3464 2281 3499
rect 2394 3464 2402 3499
rect 2531 3464 2539 3499
rect 1937 3458 1977 3464
rect 1937 3456 1949 3458
rect 1815 3426 1862 3432
rect 1815 3424 1823 3426
rect 1851 3424 1862 3426
rect 1522 3378 1534 3384
rect 1572 3378 1584 3384
rect 1711 3378 1723 3384
rect 1831 3378 1843 3384
rect 1871 3378 1883 3384
rect 1957 3378 1969 3384
rect 2096 3378 2108 3384
rect 2146 3378 2158 3384
rect 2423 3458 2463 3464
rect 2451 3456 2463 3458
rect 2574 3424 2582 3538
rect 2677 3493 2685 3542
rect 2795 3535 2820 3542
rect 2813 3513 2821 3535
rect 2951 3513 2959 3556
rect 2991 3550 2999 3576
rect 2977 3544 2999 3550
rect 3178 3596 3190 3602
rect 3390 3596 3402 3602
rect 3511 3596 3523 3602
rect 3651 3596 3663 3602
rect 3781 3596 3793 3602
rect 3877 3596 3889 3602
rect 3917 3596 3929 3602
rect 4071 3596 4083 3602
rect 4157 3596 4169 3602
rect 4277 3596 4289 3602
rect 4449 3596 4461 3602
rect 3079 3548 3091 3556
rect 2977 3538 2980 3544
rect 3079 3542 3103 3548
rect 2951 3499 2953 3513
rect 2677 3424 2685 3479
rect 2819 3464 2827 3499
rect 2951 3464 2959 3499
rect 2973 3482 2980 3538
rect 3095 3493 3103 3542
rect 3226 3538 3244 3540
rect 3214 3529 3244 3538
rect 3236 3501 3244 3529
rect 3336 3538 3354 3540
rect 3336 3529 3366 3538
rect 3475 3542 3483 3556
rect 3503 3556 3531 3562
rect 3491 3553 3543 3556
rect 3615 3542 3623 3556
rect 3643 3556 3671 3562
rect 3631 3553 3683 3556
rect 3751 3556 3761 3566
rect 3475 3535 3500 3542
rect 3615 3535 3640 3542
rect 3336 3501 3344 3529
rect 3407 3517 3433 3523
rect 3493 3513 3501 3535
rect 2977 3476 2980 3482
rect 3633 3513 3641 3535
rect 3751 3513 3759 3556
rect 3811 3546 3823 3556
rect 3785 3538 3823 3546
rect 3751 3499 3753 3513
rect 2977 3470 3003 3476
rect 2242 3378 2254 3384
rect 2292 3378 2304 3384
rect 2431 3378 2443 3384
rect 2547 3378 2559 3384
rect 2591 3378 2603 3384
rect 2657 3378 2669 3384
rect 2697 3378 2709 3384
rect 2995 3424 3003 3470
rect 3095 3424 3103 3479
rect 3238 3432 3245 3487
rect 3198 3426 3245 3432
rect 3198 3424 3209 3426
rect 2796 3378 2808 3384
rect 2846 3378 2858 3384
rect 2969 3378 2981 3384
rect 3071 3378 3083 3384
rect 3111 3378 3123 3384
rect 3237 3424 3245 3426
rect 3335 3432 3342 3487
rect 3499 3464 3507 3499
rect 3639 3464 3647 3499
rect 3751 3464 3759 3499
rect 3335 3426 3382 3432
rect 3335 3424 3343 3426
rect 3371 3424 3382 3426
rect 3177 3378 3189 3384
rect 3217 3378 3229 3384
rect 3351 3378 3363 3384
rect 3391 3378 3403 3384
rect 3476 3378 3488 3384
rect 3526 3378 3538 3384
rect 3794 3424 3802 3538
rect 3900 3533 3907 3576
rect 4035 3542 4043 3556
rect 4063 3556 4091 3562
rect 4051 3553 4103 3556
rect 4035 3535 4060 3542
rect 3900 3471 3907 3519
rect 4053 3513 4061 3535
rect 4176 3521 4184 3576
rect 4269 3556 4297 3562
rect 4257 3553 4309 3556
rect 4519 3596 4531 3602
rect 4619 3596 4631 3602
rect 4677 3596 4689 3602
rect 4725 3596 4737 3602
rect 4787 3596 4799 3602
rect 4929 3596 4941 3602
rect 5051 3596 5063 3602
rect 5159 3596 5171 3602
rect 5261 3596 5273 3602
rect 5323 3596 5335 3602
rect 5371 3596 5383 3602
rect 5429 3596 5441 3602
rect 5569 3596 5581 3602
rect 5657 3596 5669 3602
rect 4317 3542 4325 3556
rect 4419 3548 4431 3556
rect 4549 3548 4561 3556
rect 4300 3535 4325 3542
rect 3900 3464 3917 3471
rect 4059 3464 4067 3499
rect 3616 3378 3628 3384
rect 3666 3378 3678 3384
rect 3767 3378 3779 3384
rect 3811 3378 3823 3384
rect 4176 3424 4184 3507
rect 4299 3513 4307 3535
rect 4347 3537 4393 3543
rect 4419 3542 4443 3548
rect 4293 3464 4301 3499
rect 4435 3493 4443 3542
rect 4537 3542 4561 3548
rect 4767 3576 4780 3582
rect 4651 3570 4658 3576
rect 4647 3562 4658 3570
rect 4708 3564 4715 3576
rect 4773 3570 4780 3576
rect 4537 3493 4545 3542
rect 4597 3541 4605 3556
rect 4708 3557 4729 3564
rect 4687 3546 4693 3548
rect 4754 3546 4761 3552
rect 4597 3527 4613 3541
rect 4687 3540 4761 3546
rect 3877 3378 3889 3384
rect 4036 3378 4048 3384
rect 4086 3378 4098 3384
rect 4435 3424 4443 3479
rect 4537 3424 4545 3479
rect 4597 3464 4605 3527
rect 4613 3513 4627 3527
rect 4619 3468 4633 3476
rect 4157 3378 4169 3384
rect 4262 3378 4274 3384
rect 4312 3378 4324 3384
rect 4411 3378 4423 3384
rect 4451 3378 4463 3384
rect 4687 3468 4693 3540
rect 4754 3532 4761 3540
rect 4766 3524 4800 3532
rect 4794 3519 4800 3524
rect 4747 3506 4774 3513
rect 4653 3462 4693 3468
rect 4701 3468 4745 3474
rect 4653 3444 4659 3462
rect 4701 3454 4707 3468
rect 4813 3472 4819 3556
rect 4899 3548 4911 3556
rect 4899 3542 4923 3548
rect 4915 3493 4923 3542
rect 5015 3542 5023 3556
rect 5043 3556 5071 3562
rect 5031 3553 5083 3556
rect 5189 3548 5201 3556
rect 5177 3542 5201 3548
rect 5280 3576 5293 3582
rect 5280 3570 5287 3576
rect 5345 3564 5352 3576
rect 5015 3535 5040 3542
rect 5033 3513 5041 3535
rect 4757 3464 4819 3472
rect 4677 3448 4707 3454
rect 4725 3450 4763 3458
rect 4755 3444 4763 3450
rect 4647 3404 4659 3438
rect 4705 3430 4727 3442
rect 4755 3430 4773 3444
rect 4701 3424 4713 3430
rect 4755 3424 4763 3430
rect 4915 3424 4923 3479
rect 5039 3464 5047 3499
rect 5177 3493 5185 3542
rect 4517 3378 4529 3384
rect 4557 3378 4569 3384
rect 4617 3378 4629 3384
rect 4675 3378 4687 3384
rect 4721 3378 4733 3384
rect 4787 3378 4799 3384
rect 4891 3378 4903 3384
rect 4931 3378 4943 3384
rect 5177 3424 5185 3479
rect 5241 3472 5247 3556
rect 5331 3557 5352 3564
rect 5402 3570 5409 3576
rect 5402 3562 5413 3570
rect 5299 3546 5306 3552
rect 5367 3546 5373 3548
rect 5299 3540 5373 3546
rect 5455 3541 5463 3556
rect 5649 3556 5677 3562
rect 5539 3548 5551 3556
rect 5637 3553 5689 3556
rect 5539 3542 5563 3548
rect 5697 3542 5705 3556
rect 5299 3532 5306 3540
rect 5260 3524 5294 3532
rect 5260 3519 5266 3524
rect 5286 3506 5313 3513
rect 5241 3464 5303 3472
rect 5315 3468 5359 3474
rect 5016 3378 5028 3384
rect 5066 3378 5078 3384
rect 5297 3450 5335 3458
rect 5353 3454 5359 3468
rect 5367 3468 5373 3540
rect 5447 3527 5463 3541
rect 5433 3513 5447 3527
rect 5367 3462 5407 3468
rect 5427 3468 5441 3476
rect 5455 3464 5463 3527
rect 5555 3493 5563 3542
rect 5680 3535 5705 3542
rect 5679 3513 5687 3535
rect 5297 3444 5305 3450
rect 5353 3448 5383 3454
rect 5401 3444 5407 3462
rect 5287 3430 5305 3444
rect 5333 3430 5355 3442
rect 5297 3424 5305 3430
rect 5347 3424 5359 3430
rect 5401 3404 5413 3438
rect 5555 3424 5563 3479
rect 5673 3464 5681 3499
rect 5157 3378 5169 3384
rect 5197 3378 5209 3384
rect 5261 3378 5273 3384
rect 5327 3378 5339 3384
rect 5373 3378 5385 3384
rect 5431 3378 5443 3384
rect 5531 3378 5543 3384
rect 5571 3378 5583 3384
rect 5642 3378 5654 3384
rect 5692 3378 5704 3384
rect -62 3376 5816 3378
rect -62 3364 4 3376
rect -62 3362 5816 3364
rect -62 2898 -2 3362
rect 91 3356 103 3362
rect 176 3356 188 3362
rect 226 3356 238 3362
rect 331 3356 343 3362
rect 76 3233 84 3316
rect 397 3356 409 3362
rect 437 3356 449 3362
rect 537 3356 549 3362
rect 657 3356 669 3362
rect 701 3356 713 3362
rect 831 3356 843 3362
rect 871 3356 883 3362
rect 971 3356 983 3362
rect 1011 3356 1023 3362
rect 1111 3356 1123 3362
rect 1151 3356 1163 3362
rect 1237 3356 1249 3362
rect 1391 3356 1403 3362
rect 1491 3356 1503 3362
rect 1531 3356 1543 3362
rect 1631 3356 1643 3362
rect 1671 3356 1683 3362
rect 1791 3356 1803 3362
rect 1911 3356 1923 3362
rect 1951 3356 1963 3362
rect 2071 3356 2083 3362
rect 2157 3356 2169 3362
rect 2197 3356 2209 3362
rect 2307 3356 2319 3362
rect 2351 3356 2363 3362
rect 107 3257 123 3263
rect 76 3164 84 3219
rect 117 3183 123 3257
rect 199 3241 207 3276
rect 193 3205 201 3227
rect 316 3233 324 3316
rect 417 3261 425 3316
rect 517 3282 529 3284
rect 517 3276 557 3282
rect 175 3198 200 3205
rect 175 3184 183 3198
rect 107 3177 123 3183
rect 191 3184 243 3187
rect 203 3178 231 3184
rect 316 3164 324 3219
rect 417 3198 425 3247
rect 578 3241 586 3276
rect 417 3192 441 3198
rect 429 3184 441 3192
rect 578 3184 586 3227
rect 678 3202 686 3316
rect 721 3241 729 3276
rect 855 3261 863 3316
rect 955 3314 963 3316
rect 991 3314 1002 3316
rect 955 3308 1002 3314
rect 1095 3314 1103 3316
rect 1131 3314 1142 3316
rect 1095 3308 1142 3314
rect 727 3227 729 3241
rect 955 3253 962 3308
rect 91 3138 103 3144
rect 211 3138 223 3144
rect 331 3138 343 3144
rect 560 3173 586 3184
rect 657 3194 695 3202
rect 657 3184 669 3194
rect 721 3184 729 3227
rect 855 3198 863 3247
rect 1095 3253 1102 3308
rect 1217 3282 1229 3284
rect 1217 3276 1257 3282
rect 1278 3241 1286 3276
rect 956 3211 964 3239
rect 1096 3211 1104 3239
rect 956 3202 986 3211
rect 956 3200 974 3202
rect 719 3174 729 3184
rect 839 3192 863 3198
rect 839 3184 851 3192
rect 1096 3202 1126 3211
rect 1376 3233 1384 3316
rect 1475 3314 1483 3316
rect 1511 3314 1522 3316
rect 1475 3308 1522 3314
rect 1615 3314 1623 3316
rect 1651 3314 1662 3316
rect 1615 3308 1662 3314
rect 1475 3253 1482 3308
rect 1615 3253 1622 3308
rect 1867 3297 1893 3303
rect 1811 3282 1823 3284
rect 1783 3276 1823 3282
rect 1754 3241 1762 3276
rect 1935 3261 1943 3316
rect 2091 3282 2103 3284
rect 2063 3276 2103 3282
rect 1096 3200 1114 3202
rect 1278 3184 1286 3227
rect 399 3138 411 3144
rect 520 3138 532 3144
rect 570 3138 582 3144
rect 687 3138 699 3144
rect 869 3138 881 3144
rect 1010 3138 1022 3144
rect 1150 3138 1162 3144
rect 1260 3173 1286 3184
rect 1376 3164 1384 3219
rect 1476 3211 1484 3239
rect 1616 3211 1624 3239
rect 1476 3202 1506 3211
rect 1476 3200 1494 3202
rect 1616 3202 1646 3211
rect 1616 3200 1634 3202
rect 1754 3184 1762 3227
rect 1935 3198 1943 3247
rect 2034 3241 2042 3276
rect 2177 3261 2185 3316
rect 2417 3356 2429 3362
rect 2457 3356 2469 3362
rect 2556 3356 2568 3362
rect 2606 3356 2618 3362
rect 2731 3356 2743 3362
rect 2817 3356 2829 3362
rect 2857 3356 2869 3362
rect 2957 3356 2969 3362
rect 2997 3356 3009 3362
rect 3111 3356 3123 3362
rect 3151 3356 3163 3362
rect 1919 3192 1943 3198
rect 1919 3184 1931 3192
rect 2034 3184 2042 3227
rect 2177 3198 2185 3247
rect 2291 3241 2299 3276
rect 2291 3227 2293 3241
rect 2177 3192 2201 3198
rect 2189 3184 2201 3192
rect 1754 3173 1780 3184
rect 1220 3138 1232 3144
rect 1270 3138 1282 3144
rect 1391 3138 1403 3144
rect 1530 3138 1542 3144
rect 1670 3138 1682 3144
rect 2034 3173 2060 3184
rect 1758 3138 1770 3144
rect 1808 3138 1820 3144
rect 1949 3138 1961 3144
rect 2038 3138 2050 3144
rect 2088 3138 2100 3144
rect 2291 3184 2299 3227
rect 2334 3202 2342 3316
rect 2437 3261 2445 3316
rect 2838 3314 2849 3316
rect 2877 3314 2885 3316
rect 2838 3308 2885 3314
rect 2978 3314 2989 3316
rect 3251 3356 3263 3362
rect 3291 3356 3303 3362
rect 3357 3356 3369 3362
rect 3491 3356 3503 3362
rect 3531 3356 3543 3362
rect 3617 3356 3629 3362
rect 3756 3356 3768 3362
rect 3806 3356 3818 3362
rect 3017 3314 3025 3316
rect 2978 3308 3025 3314
rect 2751 3282 2763 3284
rect 2723 3276 2763 3282
rect 2325 3194 2363 3202
rect 2351 3184 2363 3194
rect 2437 3198 2445 3247
rect 2579 3241 2587 3276
rect 2694 3241 2702 3276
rect 2878 3253 2885 3308
rect 2573 3205 2581 3227
rect 3018 3253 3025 3308
rect 3135 3261 3143 3316
rect 3275 3261 3283 3316
rect 2555 3198 2580 3205
rect 2437 3192 2461 3198
rect 2449 3184 2461 3192
rect 2555 3184 2563 3198
rect 2291 3174 2301 3184
rect 2571 3184 2623 3187
rect 2583 3178 2611 3184
rect 2694 3184 2702 3227
rect 2807 3217 2833 3223
rect 2876 3211 2884 3239
rect 2947 3217 2973 3223
rect 3016 3211 3024 3239
rect 2694 3173 2720 3184
rect 2159 3138 2171 3144
rect 2321 3138 2333 3144
rect 2419 3138 2431 3144
rect 2591 3138 2603 3144
rect 2698 3138 2710 3144
rect 2748 3138 2760 3144
rect 2854 3202 2884 3211
rect 2866 3200 2884 3202
rect 2887 3177 2933 3183
rect 2994 3202 3024 3211
rect 3006 3200 3024 3202
rect 3135 3198 3143 3247
rect 3275 3198 3283 3247
rect 3376 3233 3384 3316
rect 3475 3314 3483 3316
rect 3511 3314 3522 3316
rect 3475 3308 3522 3314
rect 3475 3253 3482 3308
rect 3597 3282 3609 3284
rect 3597 3276 3637 3282
rect 3877 3356 3889 3362
rect 3957 3356 3969 3362
rect 4015 3356 4027 3362
rect 4061 3356 4073 3362
rect 4127 3356 4139 3362
rect 4222 3356 4234 3362
rect 4272 3356 4284 3362
rect 3658 3241 3666 3276
rect 3779 3241 3787 3276
rect 3119 3192 3143 3198
rect 3259 3192 3283 3198
rect 3119 3184 3131 3192
rect 3259 3184 3271 3192
rect 3376 3164 3384 3219
rect 3476 3211 3484 3239
rect 3476 3202 3506 3211
rect 3476 3200 3494 3202
rect 2818 3138 2830 3144
rect 2958 3138 2970 3144
rect 3149 3138 3161 3144
rect 3289 3138 3301 3144
rect 3658 3184 3666 3227
rect 3773 3205 3781 3227
rect 3896 3233 3904 3316
rect 3987 3302 3999 3336
rect 4041 3310 4053 3316
rect 4095 3310 4103 3316
rect 4045 3298 4067 3310
rect 4095 3296 4113 3310
rect 3993 3278 3999 3296
rect 4017 3286 4047 3292
rect 4095 3290 4103 3296
rect 3755 3198 3780 3205
rect 3755 3184 3763 3198
rect 3357 3138 3369 3144
rect 3530 3138 3542 3144
rect 3640 3173 3666 3184
rect 3771 3184 3823 3187
rect 3783 3178 3811 3184
rect 3896 3164 3904 3219
rect 3937 3213 3945 3276
rect 3959 3264 3973 3272
rect 3993 3272 4033 3278
rect 3953 3213 3967 3227
rect 3937 3199 3953 3213
rect 4027 3200 4033 3272
rect 4041 3272 4047 3286
rect 4065 3282 4103 3290
rect 4362 3356 4374 3362
rect 4412 3356 4424 3362
rect 4477 3356 4489 3362
rect 4535 3356 4547 3362
rect 4581 3356 4593 3362
rect 4647 3356 4659 3362
rect 4742 3356 4754 3362
rect 4792 3356 4804 3362
rect 4507 3302 4519 3336
rect 4561 3310 4573 3316
rect 4615 3310 4623 3316
rect 4565 3298 4587 3310
rect 4615 3296 4633 3310
rect 4513 3278 4519 3296
rect 4537 3286 4567 3292
rect 4615 3290 4623 3296
rect 4041 3266 4085 3272
rect 4097 3268 4159 3276
rect 4087 3227 4114 3234
rect 4134 3216 4140 3221
rect 4106 3208 4140 3216
rect 4094 3200 4101 3208
rect 3937 3184 3945 3199
rect 4027 3194 4101 3200
rect 4027 3192 4033 3194
rect 4094 3188 4101 3194
rect 3987 3170 3998 3178
rect 3991 3164 3998 3170
rect 4048 3176 4069 3183
rect 4153 3184 4159 3268
rect 4253 3241 4261 3276
rect 4393 3241 4401 3276
rect 4259 3205 4267 3227
rect 4399 3205 4407 3227
rect 4457 3213 4465 3276
rect 4479 3264 4493 3272
rect 4513 3272 4553 3278
rect 4473 3213 4487 3227
rect 4260 3198 4285 3205
rect 4400 3198 4425 3205
rect 4048 3164 4055 3176
rect 4113 3164 4120 3170
rect 4107 3158 4120 3164
rect 4217 3184 4269 3187
rect 4229 3178 4257 3184
rect 4277 3184 4285 3198
rect 4357 3184 4409 3187
rect 4369 3178 4397 3184
rect 4417 3184 4425 3198
rect 4457 3199 4473 3213
rect 4547 3200 4553 3272
rect 4561 3272 4567 3286
rect 4585 3282 4623 3290
rect 4891 3356 4903 3362
rect 4931 3356 4943 3362
rect 5016 3356 5028 3362
rect 5066 3356 5078 3362
rect 5171 3356 5183 3362
rect 4561 3266 4605 3272
rect 4617 3268 4679 3276
rect 4607 3227 4634 3234
rect 4654 3216 4660 3221
rect 4626 3208 4660 3216
rect 4614 3200 4621 3208
rect 4457 3184 4465 3199
rect 4547 3194 4621 3200
rect 4547 3192 4553 3194
rect 4614 3188 4621 3194
rect 4507 3170 4518 3178
rect 4511 3164 4518 3170
rect 4568 3176 4589 3183
rect 4673 3184 4679 3268
rect 4773 3241 4781 3276
rect 4915 3261 4923 3316
rect 5251 3356 5263 3362
rect 5291 3356 5303 3362
rect 5357 3356 5369 3362
rect 5482 3356 5494 3362
rect 5532 3356 5544 3362
rect 4779 3205 4787 3227
rect 4780 3198 4805 3205
rect 4915 3198 4923 3247
rect 5039 3241 5047 3276
rect 5033 3205 5041 3227
rect 5156 3233 5164 3316
rect 5275 3261 5283 3316
rect 4568 3164 4575 3176
rect 4633 3164 4640 3170
rect 4627 3158 4640 3164
rect 4737 3184 4789 3187
rect 4749 3178 4777 3184
rect 4797 3184 4805 3198
rect 4899 3192 4923 3198
rect 5015 3198 5040 3205
rect 4899 3184 4911 3192
rect 5015 3184 5023 3198
rect 5031 3184 5083 3187
rect 5043 3178 5071 3184
rect 5156 3164 5164 3219
rect 5275 3198 5283 3247
rect 5376 3233 5384 3316
rect 5651 3356 5663 3362
rect 5691 3356 5703 3362
rect 5513 3241 5521 3276
rect 5675 3261 5683 3316
rect 5259 3192 5283 3198
rect 5259 3184 5271 3192
rect 5376 3164 5384 3219
rect 5519 3205 5527 3227
rect 5520 3198 5545 3205
rect 5675 3198 5683 3247
rect 5477 3184 5529 3187
rect 3600 3138 3612 3144
rect 3650 3138 3662 3144
rect 3791 3138 3803 3144
rect 3877 3138 3889 3144
rect 3959 3138 3971 3144
rect 4017 3138 4029 3144
rect 4065 3138 4077 3144
rect 4127 3138 4139 3144
rect 4237 3138 4249 3144
rect 4377 3138 4389 3144
rect 4479 3138 4491 3144
rect 4537 3138 4549 3144
rect 4585 3138 4597 3144
rect 4647 3138 4659 3144
rect 4757 3138 4769 3144
rect 4929 3138 4941 3144
rect 5051 3138 5063 3144
rect 5171 3138 5183 3144
rect 5289 3138 5301 3144
rect 5489 3178 5517 3184
rect 5537 3184 5545 3198
rect 5659 3192 5683 3198
rect 5659 3184 5671 3192
rect 5357 3138 5369 3144
rect 5497 3138 5509 3144
rect 5689 3138 5701 3144
rect 5822 3138 5882 3602
rect 4 3136 5882 3138
rect 5816 3124 5882 3136
rect 4 3122 5882 3124
rect 121 3116 133 3122
rect 238 3116 250 3122
rect 379 3116 391 3122
rect 551 3116 563 3122
rect 657 3116 669 3122
rect 797 3116 809 3122
rect 937 3116 949 3122
rect 1109 3116 1121 3122
rect 91 3076 101 3086
rect 91 3033 99 3076
rect 151 3066 163 3076
rect 125 3058 163 3066
rect 91 3019 93 3033
rect 91 2984 99 3019
rect 134 2944 142 3058
rect 409 3068 421 3076
rect 397 3062 421 3068
rect 515 3062 523 3076
rect 543 3076 571 3082
rect 531 3073 583 3076
rect 649 3076 677 3082
rect 637 3073 689 3076
rect 789 3076 817 3082
rect 697 3062 705 3076
rect 777 3073 829 3076
rect 929 3076 957 3082
rect 837 3062 845 3076
rect 917 3073 969 3076
rect 1211 3116 1223 3122
rect 1251 3116 1263 3122
rect 1337 3116 1349 3122
rect 1530 3116 1542 3122
rect 977 3062 985 3076
rect 1079 3068 1091 3076
rect 1079 3062 1103 3068
rect 286 3058 304 3060
rect 274 3049 304 3058
rect 296 3021 304 3049
rect 397 3013 405 3062
rect 515 3055 540 3062
rect 680 3055 705 3062
rect 820 3055 845 3062
rect 960 3055 985 3062
rect 533 3033 541 3055
rect 298 2952 305 3007
rect 679 3033 687 3055
rect 819 3033 827 3055
rect 959 3033 967 3055
rect 987 3037 1013 3043
rect 258 2946 305 2952
rect 258 2944 269 2946
rect 107 2898 119 2904
rect 151 2898 163 2904
rect 297 2944 305 2946
rect 397 2944 405 2999
rect 539 2984 547 3019
rect 673 2984 681 3019
rect 813 2984 821 3019
rect 953 2984 961 3019
rect 1095 3013 1103 3062
rect 1233 3053 1240 3096
rect 1329 3076 1357 3082
rect 1317 3073 1369 3076
rect 1377 3062 1385 3076
rect 1360 3055 1385 3062
rect 1476 3058 1494 3060
rect 237 2898 249 2904
rect 277 2898 289 2904
rect 377 2898 389 2904
rect 417 2898 429 2904
rect 516 2898 528 2904
rect 566 2898 578 2904
rect 642 2898 654 2904
rect 692 2898 704 2904
rect 782 2898 794 2904
rect 832 2898 844 2904
rect 1095 2944 1103 2999
rect 1233 2991 1240 3039
rect 1359 3033 1367 3055
rect 1476 3049 1506 3058
rect 1638 3116 1650 3122
rect 1688 3116 1700 3122
rect 1811 3116 1823 3122
rect 1917 3116 1929 3122
rect 2111 3116 2123 3122
rect 2251 3116 2263 3122
rect 2378 3116 2390 3122
rect 2428 3116 2440 3122
rect 1634 3076 1660 3087
rect 1476 3021 1484 3049
rect 1634 3033 1642 3076
rect 1775 3062 1783 3076
rect 1803 3076 1831 3082
rect 1791 3073 1843 3076
rect 1909 3076 1937 3082
rect 1897 3073 1949 3076
rect 1957 3062 1965 3076
rect 1775 3055 1800 3062
rect 1940 3055 1965 3062
rect 2075 3062 2083 3076
rect 2103 3076 2131 3082
rect 2091 3073 2143 3076
rect 2215 3062 2223 3076
rect 2243 3076 2271 3082
rect 2231 3073 2283 3076
rect 2374 3076 2400 3087
rect 2518 3116 2530 3122
rect 2568 3116 2580 3122
rect 2514 3076 2540 3087
rect 2672 3116 2684 3122
rect 2728 3116 2740 3122
rect 2831 3116 2843 3122
rect 2875 3116 2883 3122
rect 2937 3116 2949 3122
rect 2977 3116 2989 3122
rect 3079 3116 3091 3122
rect 3241 3116 3253 3122
rect 3337 3116 3345 3122
rect 3377 3116 3389 3122
rect 3531 3116 3543 3122
rect 3671 3116 3683 3122
rect 3791 3116 3803 3122
rect 3835 3116 3843 3122
rect 3961 3116 3973 3122
rect 4057 3116 4069 3122
rect 4097 3116 4109 3122
rect 2075 3055 2100 3062
rect 2215 3055 2240 3062
rect 1223 2984 1240 2991
rect 1353 2984 1361 3019
rect 1793 3033 1801 3055
rect 1939 3033 1947 3055
rect 2093 3033 2101 3055
rect 2233 3033 2241 3055
rect 2374 3033 2382 3076
rect 2514 3033 2522 3076
rect 2700 3033 2707 3076
rect 2813 3041 2820 3076
rect 2851 3068 2857 3096
rect 2847 3062 2857 3068
rect 922 2898 934 2904
rect 972 2898 984 2904
rect 1071 2898 1083 2904
rect 1111 2898 1123 2904
rect 1251 2898 1263 2904
rect 1475 2952 1482 3007
rect 1634 2984 1642 3019
rect 1799 2984 1807 3019
rect 1933 2984 1941 3019
rect 2099 2984 2107 3019
rect 2239 2984 2247 3019
rect 2374 2984 2382 3019
rect 2514 2984 2522 3019
rect 2547 2997 2593 3003
rect 2693 2996 2699 3019
rect 2672 2990 2699 2996
rect 2672 2984 2684 2990
rect 1475 2946 1522 2952
rect 1475 2944 1483 2946
rect 1511 2944 1522 2946
rect 1663 2978 1703 2984
rect 1691 2976 1703 2978
rect 1322 2898 1334 2904
rect 1372 2898 1384 2904
rect 1491 2898 1503 2904
rect 1531 2898 1543 2904
rect 1671 2898 1683 2904
rect 1776 2898 1788 2904
rect 1826 2898 1838 2904
rect 1902 2898 1914 2904
rect 1952 2898 1964 2904
rect 2076 2898 2088 2904
rect 2126 2898 2138 2904
rect 2403 2978 2443 2984
rect 2431 2976 2443 2978
rect 2543 2978 2583 2984
rect 2571 2976 2583 2978
rect 2817 2983 2826 3027
rect 2836 3001 2842 3056
rect 2960 3053 2967 3096
rect 3109 3068 3121 3076
rect 2847 2992 2883 3000
rect 2875 2984 2883 2992
rect 2960 2991 2967 3039
rect 3097 3062 3121 3068
rect 3211 3076 3221 3086
rect 3097 3013 3105 3062
rect 3211 3033 3219 3076
rect 3271 3066 3283 3076
rect 3245 3058 3283 3066
rect 3363 3068 3369 3096
rect 3363 3062 3373 3068
rect 3127 3012 3153 3018
rect 3211 3019 3213 3033
rect 2960 2984 2977 2991
rect 2663 2904 2691 2910
rect 2703 2976 2731 2982
rect 2817 2974 2821 2983
rect 3097 2944 3105 2999
rect 3211 2984 3219 3019
rect 3254 2944 3262 3058
rect 3378 3001 3384 3056
rect 3400 3041 3407 3076
rect 3495 3062 3503 3076
rect 3523 3076 3551 3082
rect 3511 3073 3563 3076
rect 3635 3062 3643 3076
rect 3663 3076 3691 3082
rect 3651 3073 3703 3076
rect 3495 3055 3520 3062
rect 3635 3055 3660 3062
rect 3513 3033 3521 3055
rect 3337 2992 3373 3000
rect 3337 2984 3345 2992
rect 3394 2983 3403 3027
rect 3653 3033 3661 3055
rect 3773 3041 3780 3076
rect 3811 3068 3817 3096
rect 3807 3062 3817 3068
rect 3931 3076 3941 3086
rect 4178 3116 4190 3122
rect 4301 3116 4313 3122
rect 4363 3116 4375 3122
rect 4411 3116 4423 3122
rect 4469 3116 4481 3122
rect 4597 3116 4609 3122
rect 4737 3116 4749 3122
rect 4909 3116 4921 3122
rect 3519 2984 3527 3019
rect 3659 2984 3667 3019
rect 3399 2974 3403 2983
rect 2216 2898 2228 2904
rect 2266 2898 2278 2904
rect 2411 2898 2423 2904
rect 2551 2898 2563 2904
rect 2711 2898 2723 2904
rect 2841 2898 2853 2904
rect 2937 2898 2949 2904
rect 3077 2898 3089 2904
rect 3117 2898 3129 2904
rect 3227 2898 3239 2904
rect 3271 2898 3283 2904
rect 3367 2898 3379 2904
rect 3496 2898 3508 2904
rect 3546 2898 3558 2904
rect 3777 2983 3786 3027
rect 3796 3001 3802 3056
rect 3931 3033 3939 3076
rect 3991 3066 4003 3076
rect 3965 3058 4003 3066
rect 3931 3019 3933 3033
rect 3807 2992 3843 3000
rect 3835 2984 3843 2992
rect 3931 2984 3939 3019
rect 3777 2974 3781 2983
rect 3974 2944 3982 3058
rect 4080 3053 4087 3096
rect 4320 3096 4333 3102
rect 4320 3090 4327 3096
rect 4385 3084 4392 3096
rect 4226 3058 4244 3060
rect 4214 3049 4244 3058
rect 4080 2991 4087 3039
rect 4236 3021 4244 3049
rect 4080 2984 4097 2991
rect 3636 2898 3648 2904
rect 3686 2898 3698 2904
rect 3801 2898 3813 2904
rect 3947 2898 3959 2904
rect 3991 2898 4003 2904
rect 4238 2952 4245 3007
rect 4198 2946 4245 2952
rect 4198 2944 4209 2946
rect 4237 2944 4245 2946
rect 4281 2992 4287 3076
rect 4371 3077 4392 3084
rect 4442 3090 4449 3096
rect 4442 3082 4453 3090
rect 4339 3066 4346 3072
rect 4407 3066 4413 3068
rect 4339 3060 4413 3066
rect 4495 3061 4503 3076
rect 4589 3076 4617 3082
rect 4577 3073 4629 3076
rect 4729 3076 4757 3082
rect 4637 3062 4645 3076
rect 4717 3073 4769 3076
rect 4979 3116 4991 3122
rect 5081 3116 5093 3122
rect 5143 3116 5155 3122
rect 5191 3116 5203 3122
rect 5249 3116 5261 3122
rect 5351 3116 5363 3122
rect 5391 3116 5403 3122
rect 5431 3116 5443 3122
rect 5471 3116 5483 3122
rect 5511 3116 5523 3122
rect 5559 3116 5571 3122
rect 5617 3116 5629 3122
rect 5665 3116 5677 3122
rect 5727 3116 5739 3122
rect 4777 3062 4785 3076
rect 4879 3068 4891 3076
rect 5009 3068 5021 3076
rect 4879 3062 4903 3068
rect 4339 3052 4346 3060
rect 4300 3044 4334 3052
rect 4300 3039 4306 3044
rect 4326 3026 4353 3033
rect 4281 2984 4343 2992
rect 4355 2988 4399 2994
rect 4337 2970 4375 2978
rect 4393 2974 4399 2988
rect 4407 2988 4413 3060
rect 4487 3047 4503 3061
rect 4620 3055 4645 3062
rect 4760 3055 4785 3062
rect 4473 3033 4487 3047
rect 4407 2982 4447 2988
rect 4467 2988 4481 2996
rect 4495 2984 4503 3047
rect 4619 3033 4627 3055
rect 4759 3033 4767 3055
rect 4613 2984 4621 3019
rect 4753 2984 4761 3019
rect 4895 3013 4903 3062
rect 4997 3062 5021 3068
rect 5100 3096 5113 3102
rect 5100 3090 5107 3096
rect 5165 3084 5172 3096
rect 4997 3013 5005 3062
rect 4337 2964 4345 2970
rect 4393 2968 4423 2974
rect 4441 2964 4447 2982
rect 4327 2950 4345 2964
rect 4373 2950 4395 2962
rect 4337 2944 4345 2950
rect 4387 2944 4399 2950
rect 4441 2924 4453 2958
rect 4057 2898 4069 2904
rect 4177 2898 4189 2904
rect 4217 2898 4229 2904
rect 4301 2898 4313 2904
rect 4367 2898 4379 2904
rect 4413 2898 4425 2904
rect 4471 2898 4483 2904
rect 4582 2898 4594 2904
rect 4632 2898 4644 2904
rect 4895 2944 4903 2999
rect 4997 2944 5005 2999
rect 5061 2992 5067 3076
rect 5151 3077 5172 3084
rect 5222 3090 5229 3096
rect 5222 3082 5233 3090
rect 5119 3066 5126 3072
rect 5707 3096 5720 3102
rect 5591 3090 5598 3096
rect 5587 3082 5598 3090
rect 5648 3084 5655 3096
rect 5713 3090 5720 3096
rect 5187 3066 5193 3068
rect 5119 3060 5193 3066
rect 5275 3061 5283 3076
rect 5372 3070 5384 3076
rect 5412 3070 5424 3076
rect 5451 3070 5463 3076
rect 5492 3070 5504 3076
rect 5366 3069 5384 3070
rect 5119 3052 5126 3060
rect 5080 3044 5114 3052
rect 5080 3039 5086 3044
rect 5106 3026 5133 3033
rect 5061 2984 5123 2992
rect 5135 2988 5179 2994
rect 4722 2898 4734 2904
rect 4772 2898 4784 2904
rect 4871 2898 4883 2904
rect 4911 2898 4923 2904
rect 5117 2970 5155 2978
rect 5173 2974 5179 2988
rect 5187 2988 5193 3060
rect 5267 3047 5283 3061
rect 5253 3033 5267 3047
rect 5187 2982 5227 2988
rect 5247 2988 5261 2996
rect 5275 2984 5283 3047
rect 5365 3062 5384 3069
rect 5398 3062 5424 3070
rect 5438 3062 5463 3070
rect 5477 3062 5504 3070
rect 5365 3041 5372 3062
rect 5398 3056 5406 3062
rect 5438 3056 5446 3062
rect 5477 3056 5485 3062
rect 5390 3044 5406 3056
rect 5430 3044 5446 3056
rect 5470 3044 5485 3056
rect 5537 3061 5545 3076
rect 5648 3077 5669 3084
rect 5627 3066 5633 3068
rect 5694 3066 5701 3072
rect 5367 3027 5372 3041
rect 5365 2998 5372 3027
rect 5398 2998 5406 3044
rect 5438 2998 5446 3044
rect 5477 2998 5485 3044
rect 5537 3047 5553 3061
rect 5627 3060 5701 3066
rect 5365 2990 5383 2998
rect 5398 2990 5423 2998
rect 5438 2990 5463 2998
rect 5477 2990 5503 2998
rect 5371 2984 5383 2990
rect 5411 2984 5423 2990
rect 5451 2984 5463 2990
rect 5491 2984 5503 2990
rect 5537 2984 5545 3047
rect 5553 3033 5567 3047
rect 5559 2988 5573 2996
rect 5117 2964 5125 2970
rect 5173 2968 5203 2974
rect 5221 2964 5227 2982
rect 5107 2950 5125 2964
rect 5153 2950 5175 2962
rect 5117 2944 5125 2950
rect 5167 2944 5179 2950
rect 5221 2924 5233 2958
rect 5627 2988 5633 3060
rect 5694 3052 5701 3060
rect 5706 3044 5740 3052
rect 5734 3039 5740 3044
rect 5687 3026 5714 3033
rect 5593 2982 5633 2988
rect 5641 2988 5685 2994
rect 5593 2964 5599 2982
rect 5641 2974 5647 2988
rect 5753 2992 5759 3076
rect 5697 2984 5759 2992
rect 5617 2968 5647 2974
rect 5665 2970 5703 2978
rect 5695 2964 5703 2970
rect 5587 2924 5599 2958
rect 5645 2950 5667 2962
rect 5695 2950 5713 2964
rect 5641 2944 5653 2950
rect 5695 2944 5703 2950
rect 4977 2898 4989 2904
rect 5017 2898 5029 2904
rect 5081 2898 5093 2904
rect 5147 2898 5159 2904
rect 5193 2898 5205 2904
rect 5251 2898 5263 2904
rect 5351 2898 5363 2904
rect 5391 2898 5403 2904
rect 5431 2898 5443 2904
rect 5471 2898 5483 2904
rect 5511 2898 5523 2904
rect 5557 2898 5569 2904
rect 5615 2898 5627 2904
rect 5661 2898 5673 2904
rect 5727 2898 5739 2904
rect -62 2896 5816 2898
rect -62 2884 4 2896
rect -62 2882 4373 2884
rect -62 2418 -2 2882
rect 71 2876 83 2882
rect 111 2876 123 2882
rect 182 2876 194 2882
rect 232 2876 244 2882
rect 351 2876 363 2882
rect 437 2876 449 2882
rect 571 2876 583 2882
rect 611 2876 623 2882
rect 95 2781 103 2836
rect 95 2718 103 2767
rect 213 2761 221 2796
rect 336 2753 344 2836
rect 417 2802 429 2804
rect 417 2796 457 2802
rect 677 2876 689 2882
rect 721 2876 733 2882
rect 817 2876 829 2882
rect 857 2876 869 2882
rect 957 2876 969 2882
rect 1077 2876 1089 2882
rect 1117 2876 1129 2882
rect 478 2761 486 2796
rect 595 2781 603 2836
rect 219 2725 227 2747
rect 220 2718 245 2725
rect 79 2712 103 2718
rect 79 2704 91 2712
rect 177 2704 229 2707
rect 189 2698 217 2704
rect 237 2704 245 2718
rect 336 2684 344 2739
rect 478 2704 486 2747
rect 595 2718 603 2767
rect 698 2722 706 2836
rect 741 2761 749 2796
rect 837 2781 845 2836
rect 937 2802 949 2804
rect 937 2796 977 2802
rect 1236 2876 1248 2882
rect 1286 2876 1298 2882
rect 747 2747 749 2761
rect 109 2658 121 2664
rect 197 2658 209 2664
rect 351 2658 363 2664
rect 460 2693 486 2704
rect 579 2712 603 2718
rect 677 2714 715 2722
rect 579 2704 591 2712
rect 677 2704 689 2714
rect 741 2704 749 2747
rect 837 2718 845 2767
rect 998 2761 1006 2796
rect 1097 2781 1105 2836
rect 1362 2876 1374 2882
rect 1412 2876 1424 2882
rect 1541 2876 1553 2882
rect 1637 2876 1649 2882
rect 1787 2876 1799 2882
rect 1831 2876 1843 2882
rect 1517 2797 1521 2806
rect 837 2712 861 2718
rect 849 2704 861 2712
rect 998 2704 1006 2747
rect 1097 2718 1105 2767
rect 1259 2761 1267 2796
rect 1393 2761 1401 2796
rect 1253 2725 1261 2747
rect 1517 2753 1526 2797
rect 1931 2876 1943 2882
rect 1971 2876 1983 2882
rect 2042 2876 2054 2882
rect 2092 2876 2104 2882
rect 2207 2876 2219 2882
rect 2251 2876 2263 2882
rect 1575 2788 1583 2796
rect 1547 2780 1583 2788
rect 1660 2789 1677 2796
rect 1399 2725 1407 2747
rect 1235 2718 1260 2725
rect 1400 2718 1425 2725
rect 1097 2712 1121 2718
rect 1109 2704 1121 2712
rect 1235 2704 1243 2718
rect 739 2694 749 2704
rect 980 2693 1006 2704
rect 420 2658 432 2664
rect 470 2658 482 2664
rect 609 2658 621 2664
rect 707 2658 719 2664
rect 819 2658 831 2664
rect 940 2658 952 2664
rect 990 2658 1002 2664
rect 1251 2704 1303 2707
rect 1263 2698 1291 2704
rect 1357 2704 1409 2707
rect 1369 2698 1397 2704
rect 1417 2704 1425 2718
rect 1513 2704 1520 2739
rect 1536 2724 1542 2779
rect 1660 2741 1667 2789
rect 1771 2761 1779 2796
rect 1771 2747 1773 2761
rect 1547 2712 1557 2718
rect 1551 2684 1557 2712
rect 1607 2697 1633 2703
rect 1660 2684 1667 2727
rect 1771 2704 1779 2747
rect 1814 2722 1822 2836
rect 1955 2781 1963 2836
rect 2331 2876 2343 2882
rect 2371 2876 2383 2882
rect 2457 2876 2469 2882
rect 2611 2876 2623 2882
rect 2651 2876 2663 2882
rect 2747 2876 2759 2882
rect 2791 2876 2803 2882
rect 1805 2714 1843 2722
rect 1955 2718 1963 2767
rect 2073 2761 2081 2796
rect 2191 2761 2199 2796
rect 2079 2725 2087 2747
rect 2191 2747 2193 2761
rect 2080 2718 2105 2725
rect 1831 2704 1843 2714
rect 1771 2694 1781 2704
rect 1079 2658 1091 2664
rect 1271 2658 1283 2664
rect 1377 2658 1389 2664
rect 1531 2658 1543 2664
rect 1575 2658 1583 2664
rect 1939 2712 1963 2718
rect 1939 2704 1951 2712
rect 2037 2704 2089 2707
rect 2049 2698 2077 2704
rect 2097 2704 2105 2718
rect 2191 2704 2199 2747
rect 2234 2722 2242 2836
rect 2355 2781 2363 2836
rect 2480 2789 2497 2796
rect 2595 2834 2603 2836
rect 2631 2834 2642 2836
rect 2595 2828 2642 2834
rect 2225 2714 2263 2722
rect 2355 2718 2363 2767
rect 2480 2741 2487 2789
rect 2595 2773 2602 2828
rect 2882 2876 2894 2882
rect 2932 2876 2944 2882
rect 3051 2876 3063 2882
rect 3091 2876 3103 2882
rect 2731 2761 2739 2796
rect 2251 2704 2263 2714
rect 2191 2694 2201 2704
rect 2339 2712 2363 2718
rect 2407 2717 2453 2723
rect 2339 2704 2351 2712
rect 2480 2684 2487 2727
rect 2596 2731 2604 2759
rect 2731 2747 2733 2761
rect 2596 2722 2626 2731
rect 2596 2720 2614 2722
rect 1637 2658 1649 2664
rect 1677 2658 1689 2664
rect 1801 2658 1813 2664
rect 1969 2658 1981 2664
rect 2057 2658 2069 2664
rect 2221 2658 2233 2664
rect 2369 2658 2381 2664
rect 2731 2704 2739 2747
rect 2774 2722 2782 2836
rect 3035 2834 3043 2836
rect 3157 2876 3169 2882
rect 3197 2876 3209 2882
rect 3296 2876 3308 2882
rect 3346 2876 3358 2882
rect 3447 2876 3459 2882
rect 3491 2876 3503 2882
rect 3071 2834 3082 2836
rect 3035 2828 3082 2834
rect 2913 2761 2921 2796
rect 3035 2773 3042 2828
rect 3177 2781 3185 2836
rect 3207 2797 3233 2803
rect 3557 2876 3569 2882
rect 3677 2876 3689 2882
rect 3717 2876 3729 2882
rect 3817 2876 3829 2882
rect 3857 2876 3869 2882
rect 3971 2876 3983 2882
rect 2919 2725 2927 2747
rect 3036 2731 3044 2759
rect 2765 2714 2803 2722
rect 2920 2718 2945 2725
rect 3036 2722 3066 2731
rect 3036 2720 3054 2722
rect 2791 2704 2803 2714
rect 2731 2694 2741 2704
rect 2877 2704 2929 2707
rect 2889 2698 2917 2704
rect 2937 2704 2945 2718
rect 3177 2718 3185 2767
rect 3319 2761 3327 2796
rect 3431 2761 3439 2796
rect 3313 2725 3321 2747
rect 3431 2747 3433 2761
rect 3295 2718 3320 2725
rect 3177 2712 3201 2718
rect 3189 2704 3201 2712
rect 3295 2704 3303 2718
rect 2457 2658 2469 2664
rect 2497 2658 2509 2664
rect 2650 2658 2662 2664
rect 2761 2658 2773 2664
rect 2897 2658 2909 2664
rect 3090 2658 3102 2664
rect 3311 2704 3363 2707
rect 3323 2698 3351 2704
rect 3431 2704 3439 2747
rect 3474 2722 3482 2836
rect 3698 2834 3709 2836
rect 3737 2834 3745 2836
rect 3698 2828 3745 2834
rect 3580 2789 3597 2796
rect 3580 2741 3587 2789
rect 3738 2773 3745 2828
rect 3837 2781 3845 2836
rect 4056 2876 4068 2882
rect 4106 2876 4118 2882
rect 4177 2876 4189 2882
rect 4217 2876 4229 2882
rect 4297 2876 4309 2882
rect 3736 2731 3744 2759
rect 3465 2714 3503 2722
rect 3491 2704 3503 2714
rect 3431 2694 3441 2704
rect 3580 2684 3587 2727
rect 3159 2658 3171 2664
rect 3331 2658 3343 2664
rect 3461 2658 3473 2664
rect 3557 2658 3569 2664
rect 3597 2658 3609 2664
rect 3714 2722 3744 2731
rect 3726 2720 3744 2722
rect 3837 2718 3845 2767
rect 3956 2761 3964 2796
rect 4079 2761 4087 2796
rect 4197 2781 4205 2836
rect 4387 2882 5816 2884
rect 4397 2876 4409 2882
rect 4477 2876 4489 2882
rect 4535 2876 4547 2882
rect 4581 2876 4593 2882
rect 4647 2876 4659 2882
rect 4721 2876 4733 2882
rect 4787 2876 4799 2882
rect 4833 2876 4845 2882
rect 4891 2876 4903 2882
rect 5002 2876 5014 2882
rect 5052 2876 5064 2882
rect 3837 2712 3861 2718
rect 3849 2704 3861 2712
rect 3956 2704 3964 2747
rect 4073 2725 4081 2747
rect 4055 2718 4080 2725
rect 4197 2718 4205 2767
rect 4316 2761 4324 2796
rect 4416 2753 4424 2836
rect 4507 2822 4519 2856
rect 4561 2830 4573 2836
rect 4615 2830 4623 2836
rect 4565 2818 4587 2830
rect 4615 2816 4633 2830
rect 4513 2798 4519 2816
rect 4537 2806 4567 2812
rect 4615 2810 4623 2816
rect 4055 2704 4063 2718
rect 4197 2712 4221 2718
rect 4071 2704 4123 2707
rect 4209 2704 4221 2712
rect 4316 2704 4324 2747
rect 4083 2698 4111 2704
rect 4416 2684 4424 2739
rect 4457 2733 4465 2796
rect 4479 2784 4493 2792
rect 4513 2792 4553 2798
rect 4473 2733 4487 2747
rect 4457 2719 4473 2733
rect 4547 2720 4553 2792
rect 4561 2792 4567 2806
rect 4585 2802 4623 2810
rect 4561 2786 4605 2792
rect 4617 2788 4679 2796
rect 4607 2747 4634 2754
rect 4654 2736 4660 2741
rect 4626 2728 4660 2736
rect 4614 2720 4621 2728
rect 4457 2704 4465 2719
rect 4547 2714 4621 2720
rect 4547 2712 4553 2714
rect 4614 2708 4621 2714
rect 4507 2690 4518 2698
rect 4511 2684 4518 2690
rect 4568 2696 4589 2703
rect 4673 2704 4679 2788
rect 4568 2684 4575 2696
rect 4633 2684 4640 2690
rect 4627 2678 4640 2684
rect 4757 2830 4765 2836
rect 4807 2830 4819 2836
rect 4747 2816 4765 2830
rect 4793 2818 4815 2830
rect 4861 2822 4873 2856
rect 4757 2810 4765 2816
rect 4757 2802 4795 2810
rect 4813 2806 4843 2812
rect 4701 2788 4763 2796
rect 4701 2704 4707 2788
rect 4813 2792 4819 2806
rect 4861 2798 4867 2816
rect 4775 2786 4819 2792
rect 4827 2792 4867 2798
rect 4746 2747 4773 2754
rect 4720 2736 4726 2741
rect 4720 2728 4754 2736
rect 4759 2720 4766 2728
rect 4827 2720 4833 2792
rect 5137 2876 5149 2882
rect 5177 2876 5189 2882
rect 5257 2874 5269 2882
rect 5297 2876 5309 2882
rect 5357 2876 5369 2882
rect 5415 2876 5427 2882
rect 5461 2876 5473 2882
rect 5527 2876 5539 2882
rect 5622 2876 5634 2882
rect 5672 2876 5684 2882
rect 4887 2784 4901 2792
rect 4893 2733 4907 2747
rect 4915 2733 4923 2796
rect 5033 2761 5041 2796
rect 5157 2781 5165 2836
rect 5387 2822 5399 2856
rect 5441 2830 5453 2836
rect 5495 2830 5503 2836
rect 5445 2818 5467 2830
rect 5495 2816 5513 2830
rect 5393 2798 5399 2816
rect 5417 2806 5447 2812
rect 5495 2810 5503 2816
rect 4759 2714 4833 2720
rect 4907 2719 4923 2733
rect 5039 2725 5047 2747
rect 4759 2708 4766 2714
rect 4827 2712 4833 2714
rect 4791 2696 4812 2703
rect 4915 2704 4923 2719
rect 5040 2718 5065 2725
rect 4740 2684 4747 2690
rect 4805 2684 4812 2696
rect 4862 2690 4873 2698
rect 4862 2684 4869 2690
rect 4740 2678 4753 2684
rect 4997 2704 5049 2707
rect 5009 2698 5037 2704
rect 5057 2704 5065 2718
rect 5157 2718 5165 2767
rect 5279 2753 5288 2796
rect 5279 2739 5293 2753
rect 5157 2712 5181 2718
rect 5169 2704 5181 2712
rect 5279 2704 5288 2739
rect 5337 2733 5345 2796
rect 5359 2784 5373 2792
rect 5393 2792 5433 2798
rect 5353 2733 5367 2747
rect 5337 2719 5353 2733
rect 5427 2720 5433 2792
rect 5441 2792 5447 2806
rect 5465 2802 5503 2810
rect 5441 2786 5485 2792
rect 5497 2788 5559 2796
rect 5487 2747 5514 2754
rect 5534 2736 5540 2741
rect 5506 2728 5540 2736
rect 5494 2720 5501 2728
rect 5337 2704 5345 2719
rect 5427 2714 5501 2720
rect 5427 2712 5433 2714
rect 5494 2708 5501 2714
rect 5387 2690 5398 2698
rect 5391 2684 5398 2690
rect 5448 2696 5469 2703
rect 5553 2704 5559 2788
rect 5653 2761 5661 2796
rect 5659 2725 5667 2747
rect 5660 2718 5685 2725
rect 5448 2684 5455 2696
rect 5513 2684 5520 2690
rect 5507 2678 5520 2684
rect 5617 2704 5669 2707
rect 5629 2698 5657 2704
rect 5677 2704 5685 2718
rect 3678 2658 3690 2664
rect 3819 2658 3831 2664
rect 3971 2658 3983 2664
rect 4091 2658 4103 2664
rect 4179 2658 4191 2664
rect 4297 2658 4309 2664
rect 4397 2658 4409 2664
rect 4479 2658 4491 2664
rect 4537 2658 4549 2664
rect 4585 2658 4597 2664
rect 4647 2658 4659 2664
rect 4721 2658 4733 2664
rect 4783 2658 4795 2664
rect 4831 2658 4843 2664
rect 4889 2658 4901 2664
rect 5017 2658 5029 2664
rect 5139 2658 5151 2664
rect 5257 2658 5269 2664
rect 5297 2658 5309 2664
rect 5359 2658 5371 2664
rect 5417 2658 5429 2664
rect 5465 2658 5477 2664
rect 5527 2658 5539 2664
rect 5637 2658 5649 2664
rect 5822 2658 5882 3122
rect 4 2656 5882 2658
rect 5816 2644 5882 2656
rect 4 2642 5882 2644
rect 91 2636 103 2642
rect 157 2636 169 2642
rect 278 2636 290 2642
rect 328 2636 340 2642
rect 76 2561 84 2616
rect 176 2561 184 2616
rect 274 2596 300 2607
rect 398 2636 410 2642
rect 537 2636 549 2642
rect 637 2636 649 2642
rect 677 2636 689 2642
rect 777 2636 789 2642
rect 920 2636 932 2642
rect 970 2636 982 2642
rect 1111 2636 1123 2642
rect 1249 2636 1261 2642
rect 1347 2636 1359 2642
rect 1530 2636 1542 2642
rect 274 2553 282 2596
rect 446 2578 464 2580
rect 76 2464 84 2547
rect 176 2464 184 2547
rect 434 2569 464 2578
rect 456 2541 464 2569
rect 556 2561 564 2616
rect 660 2573 667 2616
rect 769 2596 797 2602
rect 757 2593 809 2596
rect 960 2596 986 2607
rect 817 2582 825 2596
rect 800 2575 825 2582
rect 274 2504 282 2539
rect 91 2418 103 2424
rect 303 2498 343 2504
rect 331 2496 343 2498
rect 458 2472 465 2527
rect 418 2466 465 2472
rect 418 2464 429 2466
rect 457 2464 465 2466
rect 556 2464 564 2547
rect 660 2511 667 2559
rect 799 2553 807 2575
rect 978 2553 986 2596
rect 1075 2582 1083 2596
rect 1103 2596 1131 2602
rect 1091 2593 1143 2596
rect 1379 2596 1389 2606
rect 1219 2588 1231 2596
rect 1219 2582 1243 2588
rect 1075 2575 1100 2582
rect 1093 2553 1101 2575
rect 660 2504 677 2511
rect 793 2504 801 2539
rect 978 2504 986 2539
rect 1099 2504 1107 2539
rect 1235 2533 1243 2582
rect 1317 2586 1329 2596
rect 1317 2578 1355 2586
rect 917 2498 957 2504
rect 917 2496 929 2498
rect 1235 2464 1243 2519
rect 1338 2464 1346 2578
rect 1381 2553 1389 2596
rect 1387 2539 1389 2553
rect 1476 2578 1494 2580
rect 1476 2569 1506 2578
rect 1597 2636 1609 2642
rect 1717 2636 1729 2642
rect 1891 2636 1903 2642
rect 1997 2636 2009 2642
rect 2190 2636 2202 2642
rect 1476 2541 1484 2569
rect 1616 2561 1624 2616
rect 1709 2596 1737 2602
rect 1697 2593 1749 2596
rect 1757 2582 1765 2596
rect 1740 2575 1765 2582
rect 1855 2582 1863 2596
rect 1883 2596 1911 2602
rect 1871 2593 1923 2596
rect 1989 2596 2017 2602
rect 1977 2593 2029 2596
rect 2037 2582 2045 2596
rect 1855 2575 1880 2582
rect 2020 2575 2045 2582
rect 2136 2578 2154 2580
rect 1381 2504 1389 2539
rect 157 2418 169 2424
rect 311 2418 323 2424
rect 397 2418 409 2424
rect 437 2418 449 2424
rect 537 2418 549 2424
rect 637 2418 649 2424
rect 762 2418 774 2424
rect 812 2418 824 2424
rect 937 2418 949 2424
rect 1076 2418 1088 2424
rect 1126 2418 1138 2424
rect 1211 2418 1223 2424
rect 1251 2418 1263 2424
rect 1475 2472 1482 2527
rect 1475 2466 1522 2472
rect 1475 2464 1483 2466
rect 1511 2464 1522 2466
rect 1616 2464 1624 2547
rect 1739 2553 1747 2575
rect 1873 2553 1881 2575
rect 1733 2504 1741 2539
rect 1317 2418 1329 2424
rect 1361 2418 1373 2424
rect 1491 2418 1503 2424
rect 1531 2418 1543 2424
rect 1797 2503 1803 2553
rect 2019 2553 2027 2575
rect 2136 2569 2166 2578
rect 2278 2636 2290 2642
rect 2328 2636 2340 2642
rect 2274 2596 2300 2607
rect 2399 2636 2411 2642
rect 2591 2636 2603 2642
rect 2697 2636 2709 2642
rect 2838 2636 2850 2642
rect 2888 2636 2900 2642
rect 2991 2636 3003 2642
rect 3077 2636 3089 2642
rect 3219 2636 3231 2642
rect 3410 2636 3422 2642
rect 3507 2636 3519 2642
rect 3619 2636 3631 2642
rect 3740 2636 3752 2642
rect 3796 2636 3808 2642
rect 2136 2541 2144 2569
rect 2274 2553 2282 2596
rect 2429 2588 2441 2596
rect 2417 2582 2441 2588
rect 2555 2582 2563 2596
rect 2583 2596 2611 2602
rect 2571 2593 2623 2596
rect 2689 2596 2717 2602
rect 2677 2593 2729 2596
rect 2737 2582 2745 2596
rect 2834 2596 2860 2607
rect 1879 2504 1887 2539
rect 2013 2504 2021 2539
rect 1797 2497 1843 2503
rect 1767 2477 1813 2483
rect 1837 2463 1843 2497
rect 1827 2457 1843 2463
rect 1597 2418 1609 2424
rect 1702 2418 1714 2424
rect 1752 2418 1764 2424
rect 1856 2418 1868 2424
rect 1906 2418 1918 2424
rect 2135 2472 2142 2527
rect 2274 2504 2282 2539
rect 2417 2533 2425 2582
rect 2555 2575 2580 2582
rect 2720 2575 2745 2582
rect 2573 2553 2581 2575
rect 2719 2553 2727 2575
rect 2135 2466 2182 2472
rect 2135 2464 2143 2466
rect 2171 2464 2182 2466
rect 2303 2498 2343 2504
rect 2331 2496 2343 2498
rect 2417 2464 2425 2519
rect 2579 2504 2587 2539
rect 2713 2504 2721 2539
rect 2817 2527 2823 2593
rect 2834 2553 2842 2596
rect 2976 2561 2984 2616
rect 3069 2596 3097 2602
rect 3057 2593 3109 2596
rect 3117 2582 3125 2596
rect 3249 2588 3261 2596
rect 3100 2575 3125 2582
rect 2834 2504 2842 2539
rect 1982 2418 1994 2424
rect 2032 2418 2044 2424
rect 2151 2418 2163 2424
rect 2191 2418 2203 2424
rect 2311 2418 2323 2424
rect 2397 2418 2409 2424
rect 2437 2418 2449 2424
rect 2556 2418 2568 2424
rect 2606 2418 2618 2424
rect 2863 2498 2903 2504
rect 2891 2496 2903 2498
rect 2976 2464 2984 2547
rect 3099 2553 3107 2575
rect 3187 2577 3213 2583
rect 3237 2582 3261 2588
rect 3127 2557 3143 2563
rect 3137 2543 3143 2557
rect 3093 2504 3101 2539
rect 3137 2537 3193 2543
rect 3237 2533 3245 2582
rect 3356 2578 3374 2580
rect 3356 2569 3386 2578
rect 3539 2596 3549 2606
rect 3897 2636 3909 2642
rect 3937 2636 3949 2642
rect 3985 2636 3997 2642
rect 4067 2636 4079 2642
rect 4220 2636 4232 2642
rect 4270 2636 4282 2642
rect 4394 2636 4406 2642
rect 4494 2636 4506 2642
rect 4618 2636 4630 2642
rect 4668 2636 4680 2642
rect 4821 2636 4833 2642
rect 4903 2636 4915 2642
rect 4961 2636 4973 2642
rect 5023 2636 5035 2642
rect 5071 2636 5083 2642
rect 5129 2636 5141 2642
rect 5231 2636 5243 2642
rect 5271 2636 5283 2642
rect 5311 2636 5323 2642
rect 5351 2636 5363 2642
rect 5391 2636 5403 2642
rect 3477 2586 3489 2596
rect 3477 2578 3515 2586
rect 3356 2541 3364 2569
rect 2682 2418 2694 2424
rect 2732 2418 2744 2424
rect 2871 2418 2883 2424
rect 2991 2418 3003 2424
rect 3237 2464 3245 2519
rect 3355 2472 3362 2527
rect 3355 2466 3402 2472
rect 3355 2464 3363 2466
rect 3062 2418 3074 2424
rect 3112 2418 3124 2424
rect 3391 2464 3402 2466
rect 3498 2464 3506 2578
rect 3541 2553 3549 2596
rect 3649 2588 3661 2596
rect 3637 2582 3661 2588
rect 3547 2539 3549 2553
rect 3541 2504 3549 2539
rect 3637 2533 3645 2582
rect 3717 2577 3733 2583
rect 3717 2547 3723 2577
rect 3773 2553 3780 2596
rect 3920 2573 3927 2616
rect 3217 2418 3229 2424
rect 3257 2418 3269 2424
rect 3371 2418 3383 2424
rect 3411 2418 3423 2424
rect 3637 2464 3645 2519
rect 3781 2516 3787 2539
rect 3781 2510 3808 2516
rect 3796 2504 3808 2510
rect 3920 2511 3927 2559
rect 3920 2504 3937 2511
rect 3749 2496 3777 2502
rect 3789 2424 3817 2430
rect 4007 2464 4017 2616
rect 4088 2596 4104 2604
rect 4135 2610 4147 2616
rect 4155 2610 4167 2616
rect 4175 2610 4187 2616
rect 4200 2610 4212 2616
rect 4240 2610 4252 2616
rect 4200 2598 4205 2610
rect 4247 2598 4252 2610
rect 4293 2607 4302 2616
rect 4313 2607 4322 2616
rect 4333 2607 4342 2616
rect 4270 2596 4285 2605
rect 4031 2497 4039 2596
rect 4088 2572 4098 2596
rect 4141 2578 4162 2590
rect 4180 2578 4214 2590
rect 4279 2587 4285 2596
rect 4279 2581 4301 2587
rect 4180 2572 4187 2578
rect 4313 2578 4330 2586
rect 4058 2560 4078 2572
rect 4090 2560 4098 2572
rect 4121 2565 4187 2572
rect 4121 2553 4128 2565
rect 4193 2563 4244 2572
rect 4193 2558 4199 2563
rect 4073 2546 4128 2553
rect 4135 2551 4199 2558
rect 4073 2533 4087 2546
rect 4135 2540 4141 2551
rect 4106 2528 4141 2540
rect 4237 2553 4244 2563
rect 4323 2555 4330 2578
rect 4340 2572 4347 2593
rect 4358 2590 4368 2596
rect 4358 2582 4402 2590
rect 4434 2572 4442 2596
rect 4340 2566 4442 2572
rect 4237 2547 4317 2553
rect 4150 2525 4233 2533
rect 4247 2529 4292 2537
rect 4310 2537 4317 2547
rect 4347 2553 4426 2560
rect 4347 2537 4355 2553
rect 4310 2531 4355 2537
rect 4294 2519 4361 2523
rect 4120 2517 4385 2519
rect 4120 2511 4307 2517
rect 4057 2503 4127 2511
rect 4031 2491 4133 2497
rect 4187 2496 4307 2505
rect 4050 2464 4058 2491
rect 4076 2470 4102 2478
rect 4121 2473 4153 2481
rect 4090 2464 4102 2470
rect 4136 2444 4146 2452
rect 4155 2444 4167 2467
rect 4177 2444 4186 2491
rect 4294 2489 4307 2496
rect 4327 2499 4378 2507
rect 4200 2470 4206 2472
rect 4294 2482 4400 2489
rect 4247 2470 4249 2481
rect 4200 2464 4212 2470
rect 4240 2464 4249 2470
rect 4290 2453 4293 2464
rect 4370 2464 4382 2482
rect 4434 2476 4442 2566
rect 4415 2470 4442 2476
rect 4558 2607 4567 2616
rect 4578 2607 4587 2616
rect 4598 2607 4607 2616
rect 4648 2610 4660 2616
rect 4688 2610 4700 2616
rect 4458 2572 4466 2596
rect 4532 2590 4542 2596
rect 4498 2582 4542 2590
rect 4615 2596 4630 2605
rect 4648 2598 4653 2610
rect 4695 2598 4700 2610
rect 4713 2610 4725 2616
rect 4733 2610 4745 2616
rect 4753 2610 4765 2616
rect 4796 2596 4812 2604
rect 4553 2572 4560 2593
rect 4615 2587 4621 2596
rect 4458 2566 4560 2572
rect 4570 2578 4587 2586
rect 4458 2476 4466 2566
rect 4474 2553 4553 2560
rect 4570 2555 4577 2578
rect 4599 2581 4621 2587
rect 4686 2578 4720 2590
rect 4738 2578 4759 2590
rect 4713 2572 4720 2578
rect 4802 2572 4812 2596
rect 4656 2563 4707 2572
rect 4713 2565 4779 2572
rect 4545 2537 4553 2553
rect 4656 2553 4663 2563
rect 4701 2558 4707 2563
rect 4583 2547 4663 2553
rect 4583 2537 4590 2547
rect 4701 2551 4765 2558
rect 4545 2531 4590 2537
rect 4608 2529 4653 2537
rect 4667 2525 4750 2533
rect 4759 2540 4765 2551
rect 4772 2553 4779 2565
rect 4802 2560 4810 2572
rect 4822 2560 4842 2572
rect 4772 2546 4827 2553
rect 4759 2528 4794 2540
rect 4813 2533 4827 2546
rect 4539 2519 4606 2523
rect 4515 2517 4780 2519
rect 4593 2511 4780 2517
rect 4522 2499 4573 2507
rect 4593 2496 4713 2505
rect 4593 2489 4606 2496
rect 4773 2503 4843 2511
rect 4861 2497 4869 2596
rect 4767 2491 4869 2497
rect 4500 2482 4606 2489
rect 4458 2470 4485 2476
rect 4415 2464 4422 2470
rect 4478 2464 4485 2470
rect 4518 2464 4530 2482
rect 4651 2470 4653 2481
rect 4694 2470 4700 2472
rect 4290 2444 4298 2453
rect 4313 2444 4319 2453
rect 4333 2444 4341 2453
rect 4297 2424 4298 2444
rect 4317 2424 4319 2444
rect 4337 2424 4341 2444
rect 3477 2418 3489 2424
rect 3521 2418 3533 2424
rect 3617 2418 3629 2424
rect 3657 2418 3669 2424
rect 3757 2418 3769 2424
rect 3897 2418 3909 2424
rect 3985 2418 3997 2424
rect 4030 2418 4042 2424
rect 4070 2418 4082 2424
rect 4110 2418 4122 2424
rect 4220 2418 4232 2424
rect 4265 2418 4277 2424
rect 4350 2418 4362 2424
rect 4390 2418 4402 2424
rect 4430 2418 4442 2424
rect 4651 2464 4660 2470
rect 4688 2464 4700 2470
rect 4607 2453 4610 2464
rect 4559 2444 4567 2453
rect 4581 2444 4587 2453
rect 4602 2444 4610 2453
rect 4559 2424 4563 2444
rect 4581 2424 4583 2444
rect 4602 2424 4603 2444
rect 4714 2444 4723 2491
rect 4747 2473 4779 2481
rect 4798 2470 4824 2478
rect 4733 2444 4745 2467
rect 4798 2464 4810 2470
rect 4842 2464 4850 2491
rect 4883 2464 4893 2616
rect 4980 2616 4993 2622
rect 4980 2610 4987 2616
rect 5045 2604 5052 2616
rect 4941 2512 4947 2596
rect 5031 2597 5052 2604
rect 5102 2610 5109 2616
rect 5102 2602 5113 2610
rect 4999 2586 5006 2592
rect 5477 2636 5489 2642
rect 5517 2636 5529 2642
rect 5557 2636 5569 2642
rect 5597 2636 5609 2642
rect 5637 2636 5649 2642
rect 5717 2636 5729 2642
rect 5067 2586 5073 2588
rect 4999 2580 5073 2586
rect 5155 2581 5163 2596
rect 5252 2590 5264 2596
rect 5292 2590 5304 2596
rect 5331 2590 5343 2596
rect 5372 2590 5384 2596
rect 5246 2589 5264 2590
rect 4999 2572 5006 2580
rect 4960 2564 4994 2572
rect 4960 2559 4966 2564
rect 4986 2546 5013 2553
rect 4941 2504 5003 2512
rect 5015 2508 5059 2514
rect 4754 2444 4764 2452
rect 4997 2490 5035 2498
rect 5053 2494 5059 2508
rect 5067 2508 5073 2580
rect 5147 2567 5163 2581
rect 5133 2553 5147 2567
rect 5067 2502 5107 2508
rect 5127 2508 5141 2516
rect 5155 2504 5163 2567
rect 5245 2582 5264 2589
rect 5278 2582 5304 2590
rect 5318 2582 5343 2590
rect 5357 2582 5384 2590
rect 5496 2590 5508 2596
rect 5537 2590 5549 2596
rect 5576 2590 5588 2596
rect 5616 2590 5628 2596
rect 5496 2582 5523 2590
rect 5537 2582 5562 2590
rect 5576 2582 5602 2590
rect 5616 2589 5634 2590
rect 5616 2582 5635 2589
rect 5245 2561 5252 2582
rect 5278 2576 5286 2582
rect 5318 2576 5326 2582
rect 5357 2576 5365 2582
rect 5270 2564 5286 2576
rect 5310 2564 5326 2576
rect 5350 2564 5365 2576
rect 5515 2576 5523 2582
rect 5554 2576 5562 2582
rect 5594 2576 5602 2582
rect 5247 2547 5252 2561
rect 5245 2518 5252 2547
rect 5278 2518 5286 2564
rect 5318 2518 5326 2564
rect 5357 2518 5365 2564
rect 5515 2564 5530 2576
rect 5554 2564 5570 2576
rect 5594 2564 5610 2576
rect 5515 2518 5523 2564
rect 5554 2518 5562 2564
rect 5594 2518 5602 2564
rect 5628 2561 5635 2582
rect 5628 2547 5633 2561
rect 5736 2553 5744 2596
rect 5628 2518 5635 2547
rect 5245 2510 5263 2518
rect 5278 2510 5303 2518
rect 5318 2510 5343 2518
rect 5357 2510 5383 2518
rect 5251 2504 5263 2510
rect 5291 2504 5303 2510
rect 5331 2504 5343 2510
rect 5371 2504 5383 2510
rect 5497 2510 5523 2518
rect 5537 2510 5562 2518
rect 5577 2510 5602 2518
rect 5617 2510 5635 2518
rect 5497 2504 5509 2510
rect 5537 2504 5549 2510
rect 5577 2504 5589 2510
rect 5617 2504 5629 2510
rect 5736 2504 5744 2539
rect 4997 2484 5005 2490
rect 5053 2488 5083 2494
rect 5101 2484 5107 2502
rect 4987 2470 5005 2484
rect 5033 2470 5055 2482
rect 4997 2464 5005 2470
rect 5047 2464 5059 2470
rect 5101 2444 5113 2478
rect 4458 2418 4470 2424
rect 4498 2418 4510 2424
rect 4538 2418 4550 2424
rect 4623 2418 4635 2424
rect 4668 2418 4680 2424
rect 4778 2418 4790 2424
rect 4818 2418 4830 2424
rect 4858 2418 4870 2424
rect 4903 2418 4915 2424
rect 4961 2418 4973 2424
rect 5027 2418 5039 2424
rect 5073 2418 5085 2424
rect 5131 2418 5143 2424
rect 5231 2418 5243 2424
rect 5271 2418 5283 2424
rect 5311 2418 5323 2424
rect 5351 2418 5363 2424
rect 5391 2418 5403 2424
rect 5477 2418 5489 2424
rect 5517 2418 5529 2424
rect 5557 2418 5569 2424
rect 5597 2418 5609 2424
rect 5637 2418 5649 2424
rect 5717 2418 5729 2424
rect -62 2416 5816 2418
rect -62 2404 4 2416
rect -62 2402 2533 2404
rect -62 1938 -2 2402
rect 89 2396 101 2402
rect 211 2396 223 2402
rect 251 2396 263 2402
rect 71 2281 79 2316
rect 115 2310 123 2356
rect 97 2304 123 2310
rect 195 2354 203 2356
rect 317 2396 329 2402
rect 357 2396 369 2402
rect 442 2396 454 2402
rect 492 2396 504 2402
rect 231 2354 242 2356
rect 195 2348 242 2354
rect 97 2298 100 2304
rect 71 2267 73 2281
rect 71 2224 79 2267
rect 93 2242 100 2298
rect 195 2293 202 2348
rect 337 2301 345 2356
rect 596 2396 608 2402
rect 646 2396 658 2402
rect 771 2396 783 2402
rect 811 2396 823 2402
rect 755 2354 763 2356
rect 891 2396 903 2402
rect 931 2396 943 2402
rect 1041 2396 1053 2402
rect 1137 2396 1149 2402
rect 1271 2396 1283 2402
rect 1311 2396 1323 2402
rect 1431 2396 1443 2402
rect 1556 2396 1568 2402
rect 1606 2396 1618 2402
rect 1731 2396 1743 2402
rect 1851 2396 1863 2402
rect 1891 2396 1903 2402
rect 1991 2396 2003 2402
rect 2031 2396 2043 2402
rect 791 2354 802 2356
rect 755 2348 802 2354
rect 97 2236 100 2242
rect 196 2251 204 2279
rect 196 2242 226 2251
rect 196 2240 214 2242
rect 97 2230 119 2236
rect 111 2204 119 2230
rect 337 2238 345 2287
rect 473 2281 481 2316
rect 619 2281 627 2316
rect 755 2293 762 2348
rect 915 2301 923 2356
rect 1017 2317 1021 2326
rect 479 2245 487 2267
rect 613 2245 621 2267
rect 756 2251 764 2279
rect 480 2238 505 2245
rect 337 2232 361 2238
rect 349 2224 361 2232
rect 89 2178 101 2184
rect 250 2178 262 2184
rect 437 2224 489 2227
rect 449 2218 477 2224
rect 497 2224 505 2238
rect 595 2238 620 2245
rect 756 2242 786 2251
rect 756 2240 774 2242
rect 595 2224 603 2238
rect 611 2224 663 2227
rect 623 2218 651 2224
rect 915 2238 923 2287
rect 1017 2273 1026 2317
rect 1255 2354 1263 2356
rect 1291 2354 1302 2356
rect 1255 2348 1302 2354
rect 1075 2308 1083 2316
rect 1047 2300 1083 2308
rect 899 2232 923 2238
rect 899 2224 911 2232
rect 1013 2224 1020 2259
rect 1036 2244 1042 2299
rect 1156 2281 1164 2316
rect 1255 2293 1262 2348
rect 1451 2322 1463 2324
rect 1423 2316 1463 2322
rect 1751 2322 1763 2324
rect 1723 2316 1763 2322
rect 1835 2354 1843 2356
rect 1871 2354 1882 2356
rect 1835 2348 1882 2354
rect 1975 2354 1983 2356
rect 2065 2396 2077 2402
rect 2110 2396 2122 2402
rect 2150 2396 2162 2402
rect 2190 2396 2202 2402
rect 2300 2396 2312 2402
rect 2345 2396 2357 2402
rect 2430 2396 2442 2402
rect 2470 2396 2482 2402
rect 2510 2396 2522 2402
rect 2216 2368 2226 2376
rect 2011 2354 2022 2356
rect 1975 2348 2022 2354
rect 1394 2281 1402 2316
rect 1579 2281 1587 2316
rect 1694 2281 1702 2316
rect 1835 2293 1842 2348
rect 1047 2232 1057 2238
rect 1051 2204 1057 2232
rect 1156 2224 1164 2267
rect 1256 2251 1264 2279
rect 1256 2242 1286 2251
rect 1256 2240 1274 2242
rect 319 2178 331 2184
rect 457 2178 469 2184
rect 631 2178 643 2184
rect 810 2178 822 2184
rect 929 2178 941 2184
rect 1031 2178 1043 2184
rect 1075 2178 1083 2184
rect 1394 2224 1402 2267
rect 1573 2245 1581 2267
rect 1975 2293 1982 2348
rect 1555 2238 1580 2245
rect 1555 2224 1563 2238
rect 1394 2213 1420 2224
rect 1137 2178 1149 2184
rect 1310 2178 1322 2184
rect 1571 2224 1623 2227
rect 1583 2218 1611 2224
rect 1694 2224 1702 2267
rect 1836 2251 1844 2279
rect 1976 2251 1984 2279
rect 1836 2242 1866 2251
rect 1836 2240 1854 2242
rect 1694 2213 1720 2224
rect 1976 2242 2006 2251
rect 1976 2240 1994 2242
rect 2087 2204 2097 2356
rect 2130 2329 2138 2356
rect 2170 2350 2182 2356
rect 2235 2353 2247 2376
rect 2156 2342 2182 2350
rect 2201 2339 2233 2347
rect 2257 2329 2266 2376
rect 2377 2376 2378 2396
rect 2397 2376 2399 2396
rect 2417 2376 2421 2396
rect 2370 2367 2378 2376
rect 2393 2367 2399 2376
rect 2413 2367 2421 2376
rect 2370 2356 2373 2367
rect 2280 2350 2292 2356
rect 2320 2350 2329 2356
rect 2547 2402 4353 2404
rect 2609 2396 2621 2402
rect 2722 2396 2734 2402
rect 2772 2396 2784 2402
rect 2280 2348 2286 2350
rect 2327 2339 2329 2350
rect 2450 2338 2462 2356
rect 2495 2350 2502 2356
rect 2495 2344 2522 2350
rect 2374 2331 2480 2338
rect 1398 2178 1410 2184
rect 1448 2178 1460 2184
rect 1591 2178 1603 2184
rect 1698 2178 1710 2184
rect 1748 2178 1760 2184
rect 1890 2178 1902 2184
rect 2030 2178 2042 2184
rect 2111 2323 2213 2329
rect 2111 2224 2119 2323
rect 2137 2309 2207 2317
rect 2374 2324 2387 2331
rect 2267 2315 2387 2324
rect 2407 2313 2458 2321
rect 2200 2303 2387 2309
rect 2200 2301 2465 2303
rect 2374 2297 2441 2301
rect 2153 2274 2167 2287
rect 2186 2280 2221 2292
rect 2153 2267 2208 2274
rect 2138 2248 2158 2260
rect 2170 2248 2178 2260
rect 2201 2255 2208 2267
rect 2215 2269 2221 2280
rect 2230 2287 2313 2295
rect 2327 2283 2372 2291
rect 2390 2283 2435 2289
rect 2215 2262 2279 2269
rect 2390 2273 2397 2283
rect 2317 2267 2397 2273
rect 2273 2257 2279 2262
rect 2317 2257 2324 2267
rect 2427 2267 2435 2283
rect 2201 2248 2267 2255
rect 2273 2248 2324 2257
rect 2168 2224 2178 2248
rect 2260 2242 2267 2248
rect 2221 2230 2242 2242
rect 2260 2230 2294 2242
rect 2359 2233 2381 2239
rect 2403 2242 2410 2265
rect 2427 2260 2506 2267
rect 2514 2254 2522 2344
rect 2393 2234 2410 2242
rect 2420 2248 2522 2254
rect 2359 2224 2365 2233
rect 2420 2227 2427 2248
rect 2168 2216 2184 2224
rect 2215 2204 2227 2210
rect 2235 2204 2247 2210
rect 2255 2204 2267 2210
rect 2280 2210 2285 2222
rect 2327 2210 2332 2222
rect 2350 2215 2365 2224
rect 2438 2230 2482 2238
rect 2438 2224 2448 2230
rect 2514 2224 2522 2248
rect 2591 2281 2599 2316
rect 2635 2310 2643 2356
rect 2862 2396 2874 2402
rect 2912 2396 2924 2402
rect 3011 2396 3023 2402
rect 3051 2396 3063 2402
rect 3137 2396 3149 2402
rect 3177 2396 3189 2402
rect 3311 2396 3323 2402
rect 3397 2396 3409 2402
rect 3542 2396 3554 2402
rect 3592 2396 3604 2402
rect 2617 2304 2643 2310
rect 2617 2298 2620 2304
rect 2591 2267 2593 2281
rect 2591 2224 2599 2267
rect 2613 2242 2620 2298
rect 2753 2281 2761 2316
rect 2893 2281 2901 2316
rect 3035 2301 3043 2356
rect 3157 2301 3165 2356
rect 3331 2322 3343 2324
rect 3303 2316 3343 2322
rect 2759 2245 2767 2267
rect 2899 2245 2907 2267
rect 2617 2236 2620 2242
rect 2760 2238 2785 2245
rect 2900 2238 2925 2245
rect 3035 2238 3043 2287
rect 2617 2230 2639 2236
rect 2280 2204 2292 2210
rect 2320 2204 2332 2210
rect 2373 2204 2382 2213
rect 2393 2204 2402 2213
rect 2413 2204 2422 2213
rect 2631 2204 2639 2230
rect 2717 2224 2769 2227
rect 2729 2218 2757 2224
rect 2777 2224 2785 2238
rect 2857 2224 2909 2227
rect 2869 2218 2897 2224
rect 2917 2224 2925 2238
rect 3019 2232 3043 2238
rect 3157 2238 3165 2287
rect 3157 2232 3181 2238
rect 3257 2243 3263 2293
rect 3274 2281 3282 2316
rect 3467 2377 3513 2383
rect 3677 2396 3689 2402
rect 3717 2396 3729 2402
rect 3819 2396 3831 2402
rect 3885 2396 3897 2402
rect 3930 2396 3942 2402
rect 3970 2396 3982 2402
rect 4010 2396 4022 2402
rect 4120 2396 4132 2402
rect 4165 2396 4177 2402
rect 4250 2396 4262 2402
rect 4290 2396 4302 2402
rect 4330 2396 4342 2402
rect 3377 2303 3383 2313
rect 3307 2297 3383 2303
rect 3420 2309 3437 2316
rect 3227 2237 3263 2243
rect 3019 2224 3031 2232
rect 3169 2224 3181 2232
rect 2065 2178 2077 2184
rect 2147 2178 2159 2184
rect 2300 2178 2312 2184
rect 2350 2178 2362 2184
rect 2474 2178 2486 2184
rect 2609 2178 2621 2184
rect 2737 2178 2749 2184
rect 2877 2178 2889 2184
rect 3049 2178 3061 2184
rect 3274 2224 3282 2267
rect 3420 2261 3427 2309
rect 3573 2281 3581 2316
rect 3697 2301 3705 2356
rect 3797 2310 3805 2356
rect 4036 2368 4046 2376
rect 3797 2304 3823 2310
rect 3820 2298 3823 2304
rect 3274 2213 3300 2224
rect 3420 2204 3427 2247
rect 3579 2245 3587 2267
rect 3580 2238 3605 2245
rect 3537 2224 3589 2227
rect 3139 2178 3151 2184
rect 3278 2178 3290 2184
rect 3328 2178 3340 2184
rect 3549 2218 3577 2224
rect 3597 2224 3605 2238
rect 3697 2238 3705 2287
rect 3820 2242 3827 2298
rect 3841 2281 3849 2316
rect 3847 2267 3849 2281
rect 3697 2232 3721 2238
rect 3820 2236 3823 2242
rect 3709 2224 3721 2232
rect 3801 2230 3823 2236
rect 3801 2204 3809 2230
rect 3841 2224 3849 2267
rect 3907 2204 3917 2356
rect 3950 2329 3958 2356
rect 3990 2350 4002 2356
rect 4055 2353 4067 2376
rect 3976 2342 4002 2350
rect 4021 2339 4053 2347
rect 4077 2329 4086 2376
rect 4197 2376 4198 2396
rect 4217 2376 4219 2396
rect 4237 2376 4241 2396
rect 4190 2367 4198 2376
rect 4213 2367 4219 2376
rect 4233 2367 4241 2376
rect 4190 2356 4193 2367
rect 4100 2350 4112 2356
rect 4140 2350 4149 2356
rect 4367 2402 4493 2404
rect 4397 2396 4409 2402
rect 4441 2396 4453 2402
rect 4100 2348 4106 2350
rect 4147 2339 4149 2350
rect 4270 2338 4282 2356
rect 4315 2350 4322 2356
rect 4315 2344 4342 2350
rect 4194 2331 4300 2338
rect 3931 2323 4033 2329
rect 3931 2224 3939 2323
rect 3957 2309 4027 2317
rect 4194 2324 4207 2331
rect 4087 2315 4207 2324
rect 4227 2313 4278 2321
rect 4020 2303 4207 2309
rect 4020 2301 4285 2303
rect 4194 2297 4261 2301
rect 3973 2274 3987 2287
rect 4006 2280 4041 2292
rect 3973 2267 4028 2274
rect 3958 2248 3978 2260
rect 3990 2248 3998 2260
rect 4021 2255 4028 2267
rect 4035 2269 4041 2280
rect 4050 2287 4133 2295
rect 4147 2283 4192 2291
rect 4210 2283 4255 2289
rect 4035 2262 4099 2269
rect 4210 2273 4217 2283
rect 4137 2267 4217 2273
rect 4093 2257 4099 2262
rect 4137 2257 4144 2267
rect 4247 2267 4255 2283
rect 4021 2248 4087 2255
rect 4093 2248 4144 2257
rect 3988 2224 3998 2248
rect 4080 2242 4087 2248
rect 4041 2230 4062 2242
rect 4080 2230 4114 2242
rect 4179 2233 4201 2239
rect 4223 2242 4230 2265
rect 4247 2260 4326 2267
rect 4334 2254 4342 2344
rect 4213 2234 4230 2242
rect 4240 2248 4342 2254
rect 4179 2224 4185 2233
rect 4240 2227 4247 2248
rect 3988 2216 4004 2224
rect 4035 2204 4047 2210
rect 4055 2204 4067 2210
rect 4075 2204 4087 2210
rect 4100 2210 4105 2222
rect 4147 2210 4152 2222
rect 4170 2215 4185 2224
rect 4258 2230 4302 2238
rect 4258 2224 4268 2230
rect 4334 2224 4342 2248
rect 4418 2242 4426 2356
rect 4507 2402 5816 2404
rect 4557 2396 4569 2402
rect 4697 2396 4709 2402
rect 4737 2396 4749 2402
rect 4849 2396 4861 2402
rect 4937 2396 4949 2402
rect 5057 2396 5069 2402
rect 5197 2396 5209 2402
rect 5237 2396 5249 2402
rect 4549 2318 4577 2324
rect 4589 2390 4617 2396
rect 4461 2281 4469 2316
rect 4596 2310 4608 2316
rect 4581 2304 4608 2310
rect 4581 2281 4587 2304
rect 4717 2301 4725 2356
rect 4467 2267 4469 2281
rect 4100 2204 4112 2210
rect 4140 2204 4152 2210
rect 4193 2204 4202 2213
rect 4213 2204 4222 2213
rect 4233 2204 4242 2213
rect 4397 2234 4435 2242
rect 4397 2224 4409 2234
rect 4461 2224 4469 2267
rect 4573 2224 4580 2267
rect 4717 2238 4725 2287
rect 4831 2281 4839 2316
rect 4875 2310 4883 2356
rect 4857 2304 4883 2310
rect 4857 2298 4860 2304
rect 4831 2267 4833 2281
rect 4717 2232 4741 2238
rect 4729 2224 4741 2232
rect 4831 2224 4839 2267
rect 4853 2242 4860 2298
rect 4956 2273 4964 2356
rect 5049 2318 5077 2324
rect 5089 2390 5117 2396
rect 5317 2396 5329 2402
rect 5417 2396 5429 2402
rect 5457 2396 5469 2402
rect 5096 2310 5108 2316
rect 5167 2317 5193 2323
rect 5081 2304 5108 2310
rect 5081 2281 5087 2304
rect 5217 2301 5225 2356
rect 5537 2396 5549 2402
rect 5657 2388 5669 2402
rect 5717 2396 5729 2402
rect 4857 2236 4860 2242
rect 4857 2230 4879 2236
rect 4459 2214 4469 2224
rect 3397 2178 3409 2184
rect 3437 2178 3449 2184
rect 3557 2178 3569 2184
rect 3679 2178 3691 2184
rect 3819 2178 3831 2184
rect 3885 2178 3897 2184
rect 3967 2178 3979 2184
rect 4120 2178 4132 2184
rect 4170 2178 4182 2184
rect 4294 2178 4306 2184
rect 4427 2178 4439 2184
rect 4540 2178 4552 2184
rect 4596 2178 4608 2184
rect 4871 2204 4879 2230
rect 4956 2204 4964 2259
rect 5073 2224 5080 2267
rect 5267 2297 5313 2303
rect 5217 2238 5225 2287
rect 5336 2281 5344 2316
rect 5437 2301 5445 2356
rect 5217 2232 5241 2238
rect 5229 2224 5241 2232
rect 5336 2224 5344 2267
rect 5437 2238 5445 2287
rect 5556 2273 5564 2356
rect 5643 2314 5649 2348
rect 5699 2324 5701 2326
rect 5687 2320 5701 2324
rect 5643 2308 5684 2314
rect 5675 2290 5684 2308
rect 5437 2232 5461 2238
rect 5449 2224 5461 2232
rect 4699 2178 4711 2184
rect 4849 2178 4861 2184
rect 4937 2178 4949 2184
rect 5040 2178 5052 2184
rect 5096 2178 5108 2184
rect 5556 2204 5564 2259
rect 5675 2240 5684 2278
rect 5695 2273 5701 2320
rect 5642 2234 5684 2240
rect 5642 2212 5649 2234
rect 5695 2228 5701 2259
rect 5687 2224 5701 2228
rect 5699 2222 5701 2224
rect 5199 2178 5211 2184
rect 5317 2178 5329 2184
rect 5419 2178 5431 2184
rect 5537 2178 5549 2184
rect 5657 2178 5669 2192
rect 5717 2178 5729 2192
rect 5822 2178 5882 2642
rect 4 2176 5882 2178
rect 5816 2164 5882 2176
rect 4 2162 5882 2164
rect 109 2156 121 2162
rect 290 2156 302 2162
rect 91 2073 99 2116
rect 131 2110 139 2136
rect 117 2104 139 2110
rect 117 2098 120 2104
rect 91 2059 93 2073
rect 91 2024 99 2059
rect 113 2042 120 2098
rect 236 2098 254 2100
rect 236 2089 266 2098
rect 360 2156 372 2162
rect 410 2156 422 2162
rect 531 2156 543 2162
rect 651 2156 663 2162
rect 758 2156 770 2162
rect 808 2156 820 2162
rect 400 2116 426 2127
rect 236 2061 244 2089
rect 287 2077 333 2083
rect 418 2073 426 2116
rect 516 2081 524 2136
rect 615 2102 623 2116
rect 643 2116 671 2122
rect 631 2113 683 2116
rect 754 2116 780 2127
rect 878 2156 890 2162
rect 1110 2156 1122 2162
rect 1231 2156 1243 2162
rect 1371 2156 1383 2162
rect 1478 2156 1490 2162
rect 1528 2156 1540 2162
rect 1670 2156 1682 2162
rect 1757 2156 1769 2162
rect 1880 2156 1892 2162
rect 1930 2156 1942 2162
rect 2111 2156 2123 2162
rect 2151 2156 2165 2162
rect 2310 2156 2322 2162
rect 615 2095 640 2102
rect 633 2073 641 2095
rect 117 2036 120 2042
rect 117 2030 143 2036
rect 135 1984 143 2030
rect 235 1992 242 2047
rect 418 2024 426 2059
rect 357 2018 397 2024
rect 357 2016 369 2018
rect 235 1986 282 1992
rect 235 1984 243 1986
rect 271 1984 282 1986
rect 516 1984 524 2067
rect 754 2073 762 2116
rect 926 2098 944 2100
rect 914 2089 944 2098
rect 639 2024 647 2059
rect 754 2024 762 2059
rect 857 2043 863 2073
rect 936 2061 944 2089
rect 1056 2098 1074 2100
rect 1056 2089 1086 2098
rect 1195 2102 1203 2116
rect 1223 2116 1251 2122
rect 1211 2113 1263 2116
rect 1335 2102 1343 2116
rect 1363 2116 1391 2122
rect 1351 2113 1403 2116
rect 1474 2116 1500 2127
rect 1195 2095 1220 2102
rect 1335 2095 1360 2102
rect 1056 2061 1064 2089
rect 1213 2073 1221 2095
rect 827 2037 863 2043
rect 1353 2073 1361 2095
rect 1474 2073 1482 2116
rect 1616 2098 1634 2100
rect 1616 2089 1646 2098
rect 1749 2116 1777 2122
rect 1737 2113 1789 2116
rect 2091 2130 2098 2136
rect 2131 2130 2138 2136
rect 1920 2116 1946 2127
rect 1797 2102 1805 2116
rect 1780 2095 1805 2102
rect 1616 2061 1624 2089
rect 109 1938 121 1944
rect 251 1938 263 1944
rect 291 1938 303 1944
rect 377 1938 389 1944
rect 531 1938 543 1944
rect 783 2018 823 2024
rect 811 2016 823 2018
rect 938 1992 945 2047
rect 898 1986 945 1992
rect 898 1984 909 1986
rect 937 1984 945 1986
rect 1055 1992 1062 2047
rect 1219 2024 1227 2059
rect 1359 2024 1367 2059
rect 1474 2024 1482 2059
rect 1779 2073 1787 2095
rect 1938 2073 1946 2116
rect 2066 2124 2138 2130
rect 2066 2081 2074 2124
rect 2256 2098 2274 2100
rect 2256 2089 2286 2098
rect 2345 2156 2357 2162
rect 2427 2156 2439 2162
rect 2580 2156 2592 2162
rect 2630 2156 2642 2162
rect 2754 2156 2766 2162
rect 2877 2156 2889 2162
rect 3049 2156 3061 2162
rect 2067 2067 2074 2081
rect 1055 1986 1102 1992
rect 1055 1984 1063 1986
rect 1091 1984 1102 1986
rect 616 1938 628 1944
rect 666 1938 678 1944
rect 791 1938 803 1944
rect 877 1938 889 1944
rect 917 1938 929 1944
rect 1071 1938 1083 1944
rect 1111 1938 1123 1944
rect 1196 1938 1208 1944
rect 1246 1938 1258 1944
rect 1503 2018 1543 2024
rect 1531 2016 1543 2018
rect 1615 1992 1622 2047
rect 1773 2024 1781 2059
rect 1938 2024 1946 2059
rect 2066 2032 2074 2067
rect 2256 2061 2264 2089
rect 2051 2024 2074 2032
rect 1615 1986 1662 1992
rect 1615 1984 1623 1986
rect 1651 1984 1662 1986
rect 1336 1938 1348 1944
rect 1386 1938 1398 1944
rect 1511 1938 1523 1944
rect 1631 1938 1643 1944
rect 1671 1938 1683 1944
rect 1877 2018 1917 2024
rect 1877 2016 1889 2018
rect 2051 2008 2059 2024
rect 2067 2012 2123 2014
rect 2027 1950 2039 1952
rect 2079 2008 2123 2012
rect 2111 2004 2123 2008
rect 2067 1950 2079 1952
rect 2027 1944 2079 1950
rect 2131 2010 2183 2016
rect 2131 2004 2143 2010
rect 2171 2004 2183 2010
rect 2103 1944 2131 1950
rect 2255 1992 2262 2047
rect 2255 1986 2302 1992
rect 2255 1984 2263 1986
rect 2291 1984 2302 1986
rect 2367 1984 2377 2136
rect 2448 2116 2464 2124
rect 2495 2130 2507 2136
rect 2515 2130 2527 2136
rect 2535 2130 2547 2136
rect 2560 2130 2572 2136
rect 2600 2130 2612 2136
rect 2560 2118 2565 2130
rect 2607 2118 2612 2130
rect 2653 2127 2662 2136
rect 2673 2127 2682 2136
rect 2693 2127 2702 2136
rect 2630 2116 2645 2125
rect 2391 2017 2399 2116
rect 2448 2092 2458 2116
rect 2501 2098 2522 2110
rect 2540 2098 2574 2110
rect 2639 2107 2645 2116
rect 2639 2101 2661 2107
rect 2540 2092 2547 2098
rect 2673 2098 2690 2106
rect 2418 2080 2438 2092
rect 2450 2080 2458 2092
rect 2481 2085 2547 2092
rect 2481 2073 2488 2085
rect 2553 2083 2604 2092
rect 2553 2078 2559 2083
rect 2433 2066 2488 2073
rect 2495 2071 2559 2078
rect 2433 2053 2447 2066
rect 2495 2060 2501 2071
rect 2466 2048 2501 2060
rect 2597 2073 2604 2083
rect 2683 2075 2690 2098
rect 2700 2092 2707 2113
rect 2718 2110 2728 2116
rect 2718 2102 2762 2110
rect 2794 2092 2802 2116
rect 2869 2116 2897 2122
rect 2857 2113 2909 2116
rect 3119 2156 3131 2162
rect 3257 2156 3269 2162
rect 3297 2156 3309 2162
rect 3421 2156 3433 2162
rect 3520 2156 3532 2162
rect 3570 2156 3582 2162
rect 3711 2156 3723 2162
rect 2917 2102 2925 2116
rect 3019 2108 3031 2116
rect 3149 2108 3161 2116
rect 3019 2102 3043 2108
rect 2900 2095 2925 2102
rect 2700 2086 2802 2092
rect 2597 2067 2677 2073
rect 2510 2045 2593 2053
rect 2607 2049 2652 2057
rect 2670 2057 2677 2067
rect 2707 2073 2786 2080
rect 2707 2057 2715 2073
rect 2670 2051 2715 2057
rect 2654 2039 2721 2043
rect 2480 2037 2745 2039
rect 2480 2031 2667 2037
rect 2417 2023 2487 2031
rect 2391 2011 2493 2017
rect 2547 2016 2667 2025
rect 2410 1984 2418 2011
rect 2436 1990 2462 1998
rect 2481 1993 2513 2001
rect 2450 1984 2462 1990
rect 1742 1938 1754 1944
rect 1792 1938 1804 1944
rect 1897 1938 1909 1944
rect 2151 1938 2163 1944
rect 2271 1938 2283 1944
rect 2311 1938 2323 1944
rect 2496 1964 2506 1972
rect 2515 1964 2527 1987
rect 2537 1964 2546 2011
rect 2654 2009 2667 2016
rect 2687 2019 2738 2027
rect 2560 1990 2566 1992
rect 2654 2002 2760 2009
rect 2607 1990 2609 2001
rect 2560 1984 2572 1990
rect 2600 1984 2609 1990
rect 2650 1973 2653 1984
rect 2730 1984 2742 2002
rect 2794 1996 2802 2086
rect 2899 2073 2907 2095
rect 2893 2024 2901 2059
rect 3035 2053 3043 2102
rect 3137 2102 3161 2108
rect 3137 2053 3145 2102
rect 3280 2093 3287 2136
rect 2775 1990 2802 1996
rect 2775 1984 2782 1990
rect 2650 1964 2658 1973
rect 2673 1964 2679 1973
rect 2693 1964 2701 1973
rect 2657 1944 2658 1964
rect 2677 1944 2679 1964
rect 2697 1944 2701 1964
rect 2345 1938 2357 1944
rect 2390 1938 2402 1944
rect 2430 1938 2442 1944
rect 2470 1938 2482 1944
rect 2580 1938 2592 1944
rect 2625 1938 2637 1944
rect 2710 1938 2722 1944
rect 2750 1938 2762 1944
rect 2790 1938 2802 1944
rect 2927 1997 2993 2003
rect 3035 1984 3043 2039
rect 3137 1984 3145 2039
rect 3280 2031 3287 2079
rect 3391 2116 3401 2126
rect 3560 2116 3586 2127
rect 3798 2156 3810 2162
rect 3957 2156 3969 2162
rect 4121 2156 4133 2162
rect 4269 2156 4281 2162
rect 4391 2156 4403 2162
rect 4497 2156 4509 2162
rect 4619 2156 4631 2162
rect 4739 2156 4751 2162
rect 4931 2156 4943 2162
rect 5071 2156 5083 2162
rect 5157 2156 5169 2162
rect 5257 2156 5269 2162
rect 5297 2156 5309 2162
rect 3391 2073 3399 2116
rect 3451 2106 3463 2116
rect 3425 2098 3463 2106
rect 3391 2059 3393 2073
rect 3280 2024 3297 2031
rect 3391 2024 3399 2059
rect 2862 1938 2874 1944
rect 2912 1938 2924 1944
rect 3011 1938 3023 1944
rect 3051 1938 3063 1944
rect 3117 1938 3129 1944
rect 3157 1938 3169 1944
rect 3434 1984 3442 2098
rect 3578 2073 3586 2116
rect 3696 2073 3704 2116
rect 4091 2116 4101 2126
rect 3846 2098 3864 2100
rect 3834 2089 3864 2098
rect 3856 2061 3864 2089
rect 3976 2073 3984 2116
rect 4091 2073 4099 2116
rect 4151 2106 4163 2116
rect 4125 2098 4163 2106
rect 4239 2108 4251 2116
rect 4239 2102 4263 2108
rect 3578 2024 3586 2059
rect 3696 2024 3704 2059
rect 3727 2037 3773 2043
rect 4091 2059 4093 2073
rect 3517 2018 3557 2024
rect 3517 2016 3529 2018
rect 3858 1992 3865 2047
rect 3976 2024 3984 2059
rect 4091 2024 4099 2059
rect 3818 1986 3865 1992
rect 3818 1984 3829 1986
rect 3257 1938 3269 1944
rect 3407 1938 3419 1944
rect 3451 1938 3463 1944
rect 3537 1938 3549 1944
rect 3711 1938 3723 1944
rect 3857 1984 3865 1986
rect 4134 1984 4142 2098
rect 4255 2053 4263 2102
rect 4355 2102 4363 2116
rect 4383 2116 4411 2122
rect 4371 2113 4423 2116
rect 4489 2116 4517 2122
rect 4477 2113 4529 2116
rect 4537 2102 4545 2116
rect 4649 2108 4661 2116
rect 4769 2108 4781 2116
rect 4355 2095 4380 2102
rect 4520 2095 4545 2102
rect 4637 2102 4661 2108
rect 4757 2102 4781 2108
rect 4895 2102 4903 2116
rect 4923 2116 4951 2122
rect 4911 2113 4963 2116
rect 5035 2102 5043 2116
rect 5063 2116 5091 2122
rect 5379 2156 5391 2162
rect 5497 2156 5509 2162
rect 5631 2156 5643 2162
rect 5717 2156 5729 2162
rect 5051 2113 5103 2116
rect 4373 2073 4381 2095
rect 4519 2073 4527 2095
rect 4255 1984 4263 2039
rect 4379 2024 4387 2059
rect 4513 2024 4521 2059
rect 4637 2053 4645 2102
rect 4757 2053 4765 2102
rect 4895 2095 4920 2102
rect 5035 2095 5060 2102
rect 4913 2073 4921 2095
rect 5053 2073 5061 2095
rect 5176 2081 5184 2136
rect 5280 2093 5287 2136
rect 5409 2108 5421 2116
rect 3797 1938 3809 1944
rect 3837 1938 3849 1944
rect 3957 1938 3969 1944
rect 4107 1938 4119 1944
rect 4151 1938 4163 1944
rect 4231 1938 4243 1944
rect 4271 1938 4283 1944
rect 4356 1938 4368 1944
rect 4406 1938 4418 1944
rect 4637 1984 4645 2039
rect 4757 1984 4765 2039
rect 4919 2024 4927 2059
rect 5059 2024 5067 2059
rect 4482 1938 4494 1944
rect 4532 1938 4544 1944
rect 4617 1938 4629 1944
rect 4657 1938 4669 1944
rect 4737 1938 4749 1944
rect 4777 1938 4789 1944
rect 4896 1938 4908 1944
rect 4946 1938 4958 1944
rect 5176 1984 5184 2067
rect 5280 2031 5287 2079
rect 5397 2102 5421 2108
rect 5397 2053 5405 2102
rect 5516 2081 5524 2136
rect 5616 2081 5624 2136
rect 5709 2116 5737 2122
rect 5697 2113 5749 2116
rect 5757 2102 5765 2116
rect 5740 2095 5765 2102
rect 5280 2024 5297 2031
rect 5036 1938 5048 1944
rect 5086 1938 5098 1944
rect 5397 1984 5405 2039
rect 5516 1984 5524 2067
rect 5616 1984 5624 2067
rect 5739 2073 5747 2095
rect 5733 2024 5741 2059
rect 5157 1938 5169 1944
rect 5257 1938 5269 1944
rect 5377 1938 5389 1944
rect 5417 1938 5429 1944
rect 5497 1938 5509 1944
rect 5631 1938 5643 1944
rect 5702 1938 5714 1944
rect 5752 1938 5764 1944
rect -62 1936 5816 1938
rect -62 1924 4 1936
rect -62 1922 2653 1924
rect -62 1458 -2 1922
rect 91 1916 103 1922
rect 131 1916 143 1922
rect 217 1916 229 1922
rect 356 1916 368 1922
rect 406 1916 418 1922
rect 511 1916 523 1922
rect 551 1916 563 1922
rect 691 1916 703 1922
rect 777 1916 789 1922
rect 951 1916 963 1922
rect 75 1874 83 1876
rect 111 1874 122 1876
rect 75 1868 122 1874
rect 75 1813 82 1868
rect 197 1842 209 1844
rect 197 1836 237 1842
rect 495 1874 503 1876
rect 531 1874 542 1876
rect 495 1868 542 1874
rect 258 1801 266 1836
rect 379 1801 387 1836
rect 495 1813 502 1868
rect 757 1842 769 1844
rect 757 1836 797 1842
rect 1056 1916 1068 1922
rect 1106 1916 1118 1922
rect 663 1829 680 1836
rect 76 1771 84 1799
rect 76 1762 106 1771
rect 76 1760 94 1762
rect 258 1744 266 1787
rect 373 1765 381 1787
rect 496 1771 504 1799
rect 673 1781 680 1829
rect 737 1817 793 1823
rect 355 1758 380 1765
rect 496 1762 526 1771
rect 496 1760 514 1762
rect 355 1744 363 1758
rect 130 1698 142 1704
rect 240 1733 266 1744
rect 371 1744 423 1747
rect 383 1738 411 1744
rect 673 1724 680 1767
rect 737 1763 743 1817
rect 818 1801 826 1836
rect 936 1793 944 1876
rect 1196 1916 1208 1922
rect 1246 1916 1258 1922
rect 1351 1916 1363 1922
rect 1436 1916 1448 1922
rect 1486 1916 1498 1922
rect 1079 1801 1087 1836
rect 1219 1801 1227 1836
rect 707 1757 743 1763
rect 818 1744 826 1787
rect 200 1698 212 1704
rect 250 1698 262 1704
rect 391 1698 403 1704
rect 550 1698 562 1704
rect 651 1698 663 1704
rect 691 1698 703 1704
rect 800 1733 826 1744
rect 936 1724 944 1779
rect 1073 1765 1081 1787
rect 1213 1765 1221 1787
rect 1336 1793 1344 1876
rect 1562 1916 1574 1922
rect 1612 1916 1624 1922
rect 1716 1916 1728 1922
rect 1766 1916 1778 1922
rect 1851 1916 1863 1922
rect 1891 1916 1903 1922
rect 1971 1916 1983 1922
rect 2011 1916 2023 1922
rect 2111 1916 2123 1922
rect 1459 1801 1467 1836
rect 1593 1801 1601 1836
rect 1739 1801 1747 1836
rect 1875 1821 1883 1876
rect 1995 1821 2003 1876
rect 2151 1914 2163 1922
rect 2185 1916 2197 1922
rect 2230 1916 2242 1922
rect 2270 1916 2282 1922
rect 2310 1916 2322 1922
rect 2420 1916 2432 1922
rect 2465 1916 2477 1922
rect 2550 1916 2562 1922
rect 2590 1916 2602 1922
rect 2630 1916 2642 1922
rect 2336 1888 2346 1896
rect 1055 1758 1080 1765
rect 1195 1758 1220 1765
rect 1055 1744 1063 1758
rect 1071 1744 1123 1747
rect 1195 1744 1203 1758
rect 1083 1738 1111 1744
rect 1211 1744 1263 1747
rect 1223 1738 1251 1744
rect 1336 1724 1344 1779
rect 1453 1765 1461 1787
rect 1599 1765 1607 1787
rect 1733 1765 1741 1787
rect 1435 1758 1460 1765
rect 1600 1758 1625 1765
rect 1435 1744 1443 1758
rect 1451 1744 1503 1747
rect 1463 1738 1491 1744
rect 1557 1744 1609 1747
rect 1569 1738 1597 1744
rect 1617 1744 1625 1758
rect 1715 1758 1740 1765
rect 1875 1758 1883 1807
rect 1995 1758 2003 1807
rect 2132 1793 2141 1836
rect 2127 1779 2141 1793
rect 1715 1744 1723 1758
rect 1859 1752 1883 1758
rect 1979 1752 2003 1758
rect 1731 1744 1783 1747
rect 1743 1738 1771 1744
rect 1859 1744 1871 1752
rect 1979 1744 1991 1752
rect 2132 1744 2141 1779
rect 760 1698 772 1704
rect 810 1698 822 1704
rect 951 1698 963 1704
rect 1091 1698 1103 1704
rect 1231 1698 1243 1704
rect 1351 1698 1363 1704
rect 1471 1698 1483 1704
rect 1577 1698 1589 1704
rect 1751 1698 1763 1704
rect 1889 1698 1901 1704
rect 2009 1698 2021 1704
rect 2207 1724 2217 1876
rect 2250 1849 2258 1876
rect 2290 1870 2302 1876
rect 2355 1873 2367 1896
rect 2276 1862 2302 1870
rect 2321 1859 2353 1867
rect 2377 1849 2386 1896
rect 2497 1896 2498 1916
rect 2517 1896 2519 1916
rect 2537 1896 2541 1916
rect 2490 1887 2498 1896
rect 2513 1887 2519 1896
rect 2533 1887 2541 1896
rect 2490 1876 2493 1887
rect 2400 1870 2412 1876
rect 2440 1870 2449 1876
rect 2667 1922 2773 1924
rect 2697 1916 2709 1922
rect 2737 1916 2749 1922
rect 2787 1922 5816 1924
rect 2851 1916 2863 1922
rect 2891 1916 2903 1922
rect 2400 1868 2406 1870
rect 2447 1859 2449 1870
rect 2570 1858 2582 1876
rect 2615 1870 2622 1876
rect 2615 1864 2642 1870
rect 2494 1851 2600 1858
rect 2111 1698 2123 1704
rect 2151 1698 2163 1704
rect 2231 1843 2333 1849
rect 2231 1744 2239 1843
rect 2257 1829 2327 1837
rect 2494 1844 2507 1851
rect 2387 1835 2507 1844
rect 2527 1833 2578 1841
rect 2320 1823 2507 1829
rect 2320 1821 2585 1823
rect 2494 1817 2561 1821
rect 2273 1794 2287 1807
rect 2306 1800 2341 1812
rect 2273 1787 2328 1794
rect 2258 1768 2278 1780
rect 2290 1768 2298 1780
rect 2321 1775 2328 1787
rect 2335 1789 2341 1800
rect 2350 1807 2433 1815
rect 2447 1803 2492 1811
rect 2510 1803 2555 1809
rect 2335 1782 2399 1789
rect 2510 1793 2517 1803
rect 2437 1787 2517 1793
rect 2393 1777 2399 1782
rect 2437 1777 2444 1787
rect 2547 1787 2555 1803
rect 2321 1768 2387 1775
rect 2393 1768 2444 1777
rect 2288 1744 2298 1768
rect 2380 1762 2387 1768
rect 2341 1750 2362 1762
rect 2380 1750 2414 1762
rect 2479 1753 2501 1759
rect 2523 1762 2530 1785
rect 2547 1780 2626 1787
rect 2634 1774 2642 1864
rect 2717 1821 2725 1876
rect 2835 1874 2843 1876
rect 2976 1916 2988 1922
rect 3026 1916 3038 1922
rect 2871 1874 2882 1876
rect 2835 1868 2882 1874
rect 2835 1813 2842 1868
rect 3097 1916 3109 1922
rect 3237 1908 3249 1922
rect 3297 1916 3309 1922
rect 3411 1916 3423 1922
rect 2513 1754 2530 1762
rect 2540 1768 2642 1774
rect 2479 1744 2485 1753
rect 2540 1747 2547 1768
rect 2288 1736 2304 1744
rect 2335 1724 2347 1730
rect 2355 1724 2367 1730
rect 2375 1724 2387 1730
rect 2400 1730 2405 1742
rect 2447 1730 2452 1742
rect 2470 1735 2485 1744
rect 2558 1750 2602 1758
rect 2558 1744 2568 1750
rect 2634 1744 2642 1768
rect 2717 1758 2725 1807
rect 2999 1801 3007 1836
rect 3120 1829 3137 1836
rect 3223 1834 3229 1868
rect 3279 1844 3281 1846
rect 3267 1840 3281 1844
rect 2836 1771 2844 1799
rect 2836 1762 2866 1771
rect 2993 1765 3001 1787
rect 3120 1781 3127 1829
rect 3223 1828 3264 1834
rect 3255 1810 3264 1828
rect 2836 1760 2854 1762
rect 2717 1752 2741 1758
rect 2729 1744 2741 1752
rect 2400 1724 2412 1730
rect 2440 1724 2452 1730
rect 2493 1724 2502 1733
rect 2513 1724 2522 1733
rect 2533 1724 2542 1733
rect 2975 1758 3000 1765
rect 2975 1744 2983 1758
rect 2991 1744 3043 1747
rect 3003 1738 3031 1744
rect 3120 1724 3127 1767
rect 3255 1760 3264 1798
rect 3275 1793 3281 1840
rect 3477 1916 3489 1922
rect 3547 1916 3559 1922
rect 3396 1793 3404 1876
rect 3656 1916 3668 1922
rect 3706 1916 3718 1922
rect 3816 1916 3828 1922
rect 3866 1916 3878 1922
rect 3942 1916 3954 1922
rect 3992 1916 4004 1922
rect 4091 1916 4103 1922
rect 4131 1916 4143 1922
rect 4271 1916 4283 1922
rect 4371 1916 4383 1922
rect 4411 1916 4423 1922
rect 3517 1801 3525 1836
rect 3679 1801 3687 1836
rect 3839 1801 3847 1836
rect 3222 1754 3264 1760
rect 3222 1732 3229 1754
rect 3275 1748 3281 1779
rect 3267 1744 3281 1748
rect 3279 1742 3281 1744
rect 3396 1724 3404 1779
rect 3516 1761 3524 1787
rect 3673 1765 3681 1787
rect 3833 1765 3841 1787
rect 3516 1754 3545 1761
rect 3477 1744 3529 1746
rect 3539 1744 3545 1754
rect 3655 1758 3680 1765
rect 3815 1758 3840 1765
rect 3655 1744 3663 1758
rect 2185 1698 2197 1704
rect 2267 1698 2279 1704
rect 2420 1698 2432 1704
rect 2470 1698 2482 1704
rect 2594 1698 2606 1704
rect 2699 1698 2711 1704
rect 2890 1698 2902 1704
rect 3011 1698 3023 1704
rect 3097 1698 3109 1704
rect 3137 1698 3149 1704
rect 3237 1698 3249 1712
rect 3297 1698 3309 1712
rect 3489 1740 3517 1744
rect 3529 1704 3557 1710
rect 3671 1744 3723 1747
rect 3815 1744 3823 1758
rect 3917 1763 3923 1813
rect 3973 1801 3981 1836
rect 4115 1821 4123 1876
rect 4223 1910 4251 1916
rect 4263 1838 4291 1844
rect 4482 1916 4494 1922
rect 4532 1916 4544 1922
rect 4647 1916 4659 1922
rect 4691 1916 4703 1922
rect 4811 1916 4823 1922
rect 4357 1837 4373 1843
rect 4232 1830 4244 1836
rect 4232 1824 4259 1830
rect 3979 1765 3987 1787
rect 3887 1757 3923 1763
rect 3980 1758 4005 1765
rect 4115 1758 4123 1807
rect 4253 1801 4259 1824
rect 4357 1823 4363 1837
rect 4337 1817 4363 1823
rect 4395 1821 4403 1876
rect 3683 1738 3711 1744
rect 3831 1744 3883 1747
rect 3843 1738 3871 1744
rect 3937 1744 3989 1747
rect 3949 1738 3977 1744
rect 3997 1744 4005 1758
rect 4099 1752 4123 1758
rect 4099 1744 4111 1752
rect 4260 1744 4267 1787
rect 3411 1698 3423 1704
rect 3497 1698 3509 1704
rect 3691 1698 3703 1704
rect 3851 1698 3863 1704
rect 3957 1698 3969 1704
rect 4129 1698 4141 1704
rect 4337 1727 4343 1817
rect 4395 1758 4403 1807
rect 4513 1801 4521 1836
rect 4631 1801 4639 1836
rect 4519 1765 4527 1787
rect 4631 1787 4633 1801
rect 4520 1758 4545 1765
rect 4379 1752 4403 1758
rect 4379 1744 4391 1752
rect 4477 1744 4529 1747
rect 4489 1738 4517 1744
rect 4537 1744 4545 1758
rect 4631 1744 4639 1787
rect 4674 1762 4682 1876
rect 4891 1916 4903 1922
rect 4931 1916 4943 1922
rect 5071 1916 5083 1922
rect 5191 1916 5203 1922
rect 5311 1916 5323 1922
rect 4783 1829 4800 1836
rect 4793 1781 4800 1829
rect 4915 1821 4923 1876
rect 5023 1910 5051 1916
rect 5063 1838 5091 1844
rect 5032 1830 5044 1836
rect 5032 1824 5059 1830
rect 4665 1754 4703 1762
rect 4691 1744 4703 1754
rect 4631 1734 4641 1744
rect 4793 1724 4800 1767
rect 4915 1758 4923 1807
rect 5053 1801 5059 1824
rect 4899 1752 4923 1758
rect 4899 1744 4911 1752
rect 5060 1744 5067 1787
rect 5176 1793 5184 1876
rect 5382 1916 5394 1922
rect 5432 1916 5444 1922
rect 5283 1829 5300 1836
rect 5536 1916 5548 1922
rect 5586 1916 5598 1922
rect 5657 1914 5669 1922
rect 5697 1916 5709 1922
rect 5293 1781 5300 1829
rect 4232 1698 4244 1704
rect 4288 1698 4300 1704
rect 4409 1698 4421 1704
rect 4497 1698 4509 1704
rect 4661 1698 4673 1704
rect 4771 1698 4783 1704
rect 4811 1698 4823 1704
rect 4929 1698 4941 1704
rect 5176 1724 5184 1779
rect 5293 1724 5300 1767
rect 5357 1743 5363 1833
rect 5413 1801 5421 1836
rect 5559 1801 5567 1836
rect 5419 1765 5427 1787
rect 5553 1765 5561 1787
rect 5679 1793 5688 1836
rect 5679 1779 5693 1793
rect 5420 1758 5445 1765
rect 5327 1737 5363 1743
rect 5377 1744 5429 1747
rect 5032 1698 5044 1704
rect 5088 1698 5100 1704
rect 5191 1698 5203 1704
rect 5389 1738 5417 1744
rect 5437 1744 5445 1758
rect 5535 1758 5560 1765
rect 5535 1744 5543 1758
rect 5551 1744 5603 1747
rect 5679 1744 5688 1779
rect 5563 1738 5591 1744
rect 5271 1698 5283 1704
rect 5311 1698 5323 1704
rect 5397 1698 5409 1704
rect 5571 1698 5583 1704
rect 5657 1698 5669 1704
rect 5697 1698 5709 1704
rect 5822 1698 5882 2162
rect 4 1696 5882 1698
rect 5816 1684 5882 1696
rect 4 1682 5882 1684
rect 78 1676 90 1682
rect 290 1676 302 1682
rect 126 1618 144 1620
rect 114 1609 144 1618
rect 136 1581 144 1609
rect 236 1618 254 1620
rect 236 1609 266 1618
rect 360 1676 372 1682
rect 410 1676 422 1682
rect 518 1676 530 1682
rect 568 1676 580 1682
rect 400 1636 426 1647
rect 236 1581 244 1609
rect 418 1593 426 1636
rect 514 1636 540 1647
rect 639 1676 651 1682
rect 757 1676 769 1682
rect 911 1676 923 1682
rect 1070 1676 1082 1682
rect 1189 1676 1201 1682
rect 514 1593 522 1636
rect 669 1628 681 1636
rect 657 1622 681 1628
rect 138 1512 145 1567
rect 98 1506 145 1512
rect 98 1504 109 1506
rect 137 1504 145 1506
rect 235 1512 242 1567
rect 418 1544 426 1579
rect 514 1544 522 1579
rect 657 1573 665 1622
rect 776 1601 784 1656
rect 875 1622 883 1636
rect 903 1636 931 1642
rect 891 1633 943 1636
rect 875 1615 900 1622
rect 1016 1618 1034 1620
rect 893 1593 901 1615
rect 1016 1609 1046 1618
rect 1277 1676 1289 1682
rect 1317 1676 1329 1682
rect 1429 1676 1441 1682
rect 1571 1676 1583 1682
rect 1159 1628 1171 1636
rect 1159 1622 1183 1628
rect 357 1538 397 1544
rect 357 1536 369 1538
rect 235 1506 282 1512
rect 235 1504 243 1506
rect 271 1504 282 1506
rect 543 1538 583 1544
rect 571 1536 583 1538
rect 657 1504 665 1559
rect 776 1504 784 1587
rect 1016 1581 1024 1609
rect 899 1544 907 1579
rect 77 1458 89 1464
rect 117 1458 129 1464
rect 251 1458 263 1464
rect 291 1458 303 1464
rect 377 1458 389 1464
rect 551 1458 563 1464
rect 637 1458 649 1464
rect 677 1458 689 1464
rect 1015 1512 1022 1567
rect 1175 1573 1183 1622
rect 1300 1613 1307 1656
rect 1640 1676 1652 1682
rect 1696 1676 1708 1682
rect 1015 1506 1062 1512
rect 1015 1504 1023 1506
rect 1051 1504 1062 1506
rect 1175 1504 1183 1559
rect 1300 1551 1307 1599
rect 1411 1593 1419 1636
rect 1451 1630 1459 1656
rect 1437 1624 1459 1630
rect 1437 1618 1440 1624
rect 1411 1579 1413 1593
rect 1300 1544 1317 1551
rect 1411 1544 1419 1579
rect 1433 1562 1440 1618
rect 1556 1601 1564 1656
rect 1765 1676 1777 1682
rect 1847 1676 1859 1682
rect 2000 1676 2012 1682
rect 2050 1676 2062 1682
rect 2174 1676 2186 1682
rect 2317 1676 2329 1682
rect 2439 1676 2451 1682
rect 2611 1676 2623 1682
rect 2749 1676 2761 1682
rect 2871 1676 2883 1682
rect 3011 1676 3023 1682
rect 3094 1676 3106 1682
rect 3218 1676 3230 1682
rect 3268 1676 3280 1682
rect 3421 1676 3433 1682
rect 3503 1676 3515 1682
rect 1437 1556 1440 1562
rect 1437 1550 1463 1556
rect 757 1458 769 1464
rect 876 1458 888 1464
rect 926 1458 938 1464
rect 1031 1458 1043 1464
rect 1071 1458 1083 1464
rect 1151 1458 1163 1464
rect 1191 1458 1203 1464
rect 1455 1504 1463 1550
rect 1556 1504 1564 1587
rect 1673 1593 1680 1636
rect 1681 1556 1687 1579
rect 1681 1550 1708 1556
rect 1696 1544 1708 1550
rect 1649 1536 1677 1542
rect 1689 1464 1717 1470
rect 1787 1504 1797 1656
rect 1868 1636 1884 1644
rect 1915 1650 1927 1656
rect 1935 1650 1947 1656
rect 1955 1650 1967 1656
rect 1980 1650 1992 1656
rect 2020 1650 2032 1656
rect 1980 1638 1985 1650
rect 2027 1638 2032 1650
rect 2073 1647 2082 1656
rect 2093 1647 2102 1656
rect 2113 1647 2122 1656
rect 2050 1636 2065 1645
rect 1811 1537 1819 1636
rect 1868 1612 1878 1636
rect 1921 1618 1942 1630
rect 1960 1618 1994 1630
rect 2059 1627 2065 1636
rect 2059 1621 2081 1627
rect 1960 1612 1967 1618
rect 2093 1618 2110 1626
rect 1838 1600 1858 1612
rect 1870 1600 1878 1612
rect 1901 1605 1967 1612
rect 1901 1593 1908 1605
rect 1973 1603 2024 1612
rect 1973 1598 1979 1603
rect 1853 1586 1908 1593
rect 1915 1591 1979 1598
rect 1853 1573 1867 1586
rect 1915 1580 1921 1591
rect 1886 1568 1921 1580
rect 2017 1593 2024 1603
rect 2103 1595 2110 1618
rect 2120 1612 2127 1633
rect 2138 1630 2148 1636
rect 2138 1622 2182 1630
rect 2214 1612 2222 1636
rect 2309 1636 2337 1642
rect 2297 1633 2349 1636
rect 2357 1622 2365 1636
rect 2469 1628 2481 1636
rect 2340 1615 2365 1622
rect 2457 1622 2481 1628
rect 2575 1622 2583 1636
rect 2603 1636 2631 1642
rect 2591 1633 2643 1636
rect 2719 1628 2731 1636
rect 2719 1622 2743 1628
rect 2120 1606 2222 1612
rect 2017 1587 2097 1593
rect 1930 1565 2013 1573
rect 2027 1569 2072 1577
rect 2090 1577 2097 1587
rect 2127 1593 2206 1600
rect 2127 1577 2135 1593
rect 2090 1571 2135 1577
rect 2074 1559 2141 1563
rect 1900 1557 2165 1559
rect 1900 1551 2087 1557
rect 1837 1543 1907 1551
rect 1811 1531 1913 1537
rect 1967 1536 2087 1545
rect 1830 1504 1838 1531
rect 1856 1510 1882 1518
rect 1901 1513 1933 1521
rect 1870 1504 1882 1510
rect 1916 1484 1926 1492
rect 1935 1484 1947 1507
rect 1957 1484 1966 1531
rect 2074 1529 2087 1536
rect 2107 1539 2158 1547
rect 1980 1510 1986 1512
rect 2074 1522 2180 1529
rect 2027 1510 2029 1521
rect 1980 1504 1992 1510
rect 2020 1504 2029 1510
rect 2070 1493 2073 1504
rect 2150 1504 2162 1522
rect 2214 1516 2222 1606
rect 2339 1593 2347 1615
rect 2333 1544 2341 1579
rect 2457 1573 2465 1622
rect 2575 1615 2600 1622
rect 2593 1593 2601 1615
rect 2195 1510 2222 1516
rect 2195 1504 2202 1510
rect 2070 1484 2078 1493
rect 2093 1484 2099 1493
rect 2113 1484 2121 1493
rect 2077 1464 2078 1484
rect 2097 1464 2099 1484
rect 2117 1464 2121 1484
rect 1277 1458 1289 1464
rect 1429 1458 1441 1464
rect 1571 1458 1583 1464
rect 1657 1458 1669 1464
rect 1765 1458 1777 1464
rect 1810 1458 1822 1464
rect 1850 1458 1862 1464
rect 1890 1458 1902 1464
rect 2000 1458 2012 1464
rect 2045 1458 2057 1464
rect 2130 1458 2142 1464
rect 2170 1458 2182 1464
rect 2210 1458 2222 1464
rect 2457 1504 2465 1559
rect 2599 1544 2607 1579
rect 2735 1573 2743 1622
rect 2835 1622 2843 1636
rect 2863 1636 2891 1642
rect 2851 1633 2903 1636
rect 2975 1622 2983 1636
rect 3003 1636 3031 1642
rect 2991 1633 3043 1636
rect 3158 1647 3167 1656
rect 3178 1647 3187 1656
rect 3198 1647 3207 1656
rect 3248 1650 3260 1656
rect 3288 1650 3300 1656
rect 2835 1615 2860 1622
rect 2975 1615 3000 1622
rect 2787 1597 2833 1603
rect 2853 1593 2861 1615
rect 2993 1593 3001 1615
rect 3058 1612 3066 1636
rect 3132 1630 3142 1636
rect 3098 1622 3142 1630
rect 3215 1636 3230 1645
rect 3248 1638 3253 1650
rect 3295 1638 3300 1650
rect 3313 1650 3325 1656
rect 3333 1650 3345 1656
rect 3353 1650 3365 1656
rect 3396 1636 3412 1644
rect 3153 1612 3160 1633
rect 3215 1627 3221 1636
rect 3058 1606 3160 1612
rect 3170 1618 3187 1626
rect 2302 1458 2314 1464
rect 2352 1458 2364 1464
rect 2437 1458 2449 1464
rect 2477 1458 2489 1464
rect 2735 1504 2743 1559
rect 2859 1544 2867 1579
rect 2999 1544 3007 1579
rect 2576 1458 2588 1464
rect 2626 1458 2638 1464
rect 2711 1458 2723 1464
rect 2751 1458 2763 1464
rect 2836 1458 2848 1464
rect 2886 1458 2898 1464
rect 3058 1516 3066 1606
rect 3074 1593 3153 1600
rect 3170 1595 3177 1618
rect 3199 1621 3221 1627
rect 3286 1618 3320 1630
rect 3338 1618 3359 1630
rect 3313 1612 3320 1618
rect 3402 1612 3412 1636
rect 3256 1603 3307 1612
rect 3313 1605 3379 1612
rect 3145 1577 3153 1593
rect 3256 1593 3263 1603
rect 3301 1598 3307 1603
rect 3183 1587 3263 1593
rect 3183 1577 3190 1587
rect 3301 1591 3365 1598
rect 3145 1571 3190 1577
rect 3208 1569 3253 1577
rect 3267 1565 3350 1573
rect 3359 1580 3365 1591
rect 3372 1593 3379 1605
rect 3402 1600 3410 1612
rect 3422 1600 3442 1612
rect 3372 1586 3427 1593
rect 3359 1568 3394 1580
rect 3413 1573 3427 1586
rect 3139 1559 3206 1563
rect 3115 1557 3380 1559
rect 3193 1551 3380 1557
rect 3122 1539 3173 1547
rect 3193 1536 3313 1545
rect 3193 1529 3206 1536
rect 3373 1543 3443 1551
rect 3461 1537 3469 1636
rect 3367 1531 3469 1537
rect 3598 1676 3610 1682
rect 3648 1676 3660 1682
rect 3737 1676 3749 1682
rect 3889 1676 3901 1682
rect 4021 1676 4033 1682
rect 4119 1676 4131 1682
rect 4272 1676 4284 1682
rect 4328 1676 4340 1682
rect 3100 1522 3206 1529
rect 3058 1510 3085 1516
rect 3078 1504 3085 1510
rect 3118 1504 3130 1522
rect 3251 1510 3253 1521
rect 3294 1510 3300 1512
rect 2976 1458 2988 1464
rect 3026 1458 3038 1464
rect 3251 1504 3260 1510
rect 3288 1504 3300 1510
rect 3207 1493 3210 1504
rect 3159 1484 3167 1493
rect 3181 1484 3187 1493
rect 3202 1484 3210 1493
rect 3159 1464 3163 1484
rect 3181 1464 3183 1484
rect 3202 1464 3203 1484
rect 3314 1484 3323 1531
rect 3347 1513 3379 1521
rect 3398 1510 3424 1518
rect 3333 1484 3345 1507
rect 3398 1504 3410 1510
rect 3442 1504 3450 1531
rect 3483 1504 3493 1656
rect 3594 1636 3620 1647
rect 3729 1636 3757 1642
rect 3594 1593 3602 1636
rect 3717 1633 3769 1636
rect 3777 1622 3785 1636
rect 3760 1615 3785 1622
rect 3759 1593 3767 1615
rect 3871 1593 3879 1636
rect 3911 1630 3919 1656
rect 3897 1624 3919 1630
rect 3991 1636 4001 1646
rect 4432 1676 4444 1682
rect 4488 1676 4500 1682
rect 4580 1676 4592 1682
rect 4636 1676 4648 1682
rect 4739 1676 4751 1682
rect 4877 1676 4889 1682
rect 5041 1676 5053 1682
rect 5158 1676 5170 1682
rect 5300 1676 5312 1682
rect 5356 1676 5368 1682
rect 3897 1618 3900 1624
rect 3871 1579 3873 1593
rect 3594 1544 3602 1579
rect 3753 1544 3761 1579
rect 3871 1544 3879 1579
rect 3893 1562 3900 1618
rect 3991 1593 3999 1636
rect 4051 1626 4063 1636
rect 4149 1628 4161 1636
rect 4025 1618 4063 1626
rect 4137 1622 4161 1628
rect 3991 1579 3993 1593
rect 3897 1556 3900 1562
rect 3897 1550 3923 1556
rect 3354 1484 3364 1492
rect 3623 1538 3663 1544
rect 3651 1536 3663 1538
rect 3915 1504 3923 1550
rect 3991 1544 3999 1579
rect 4034 1504 4042 1618
rect 4137 1573 4145 1622
rect 4300 1593 4307 1636
rect 4460 1593 4467 1636
rect 4507 1617 4563 1623
rect 4137 1504 4145 1559
rect 4293 1556 4299 1579
rect 4453 1556 4459 1579
rect 4557 1567 4563 1617
rect 4613 1593 4620 1636
rect 4769 1628 4781 1636
rect 4869 1636 4897 1642
rect 4857 1633 4909 1636
rect 5011 1636 5021 1646
rect 4757 1622 4781 1628
rect 4917 1622 4925 1636
rect 4272 1550 4299 1556
rect 4432 1550 4459 1556
rect 4621 1556 4627 1579
rect 4757 1573 4765 1622
rect 4900 1615 4925 1622
rect 4899 1593 4907 1615
rect 5011 1593 5019 1636
rect 5071 1626 5083 1636
rect 5045 1618 5083 1626
rect 5011 1579 5013 1593
rect 4621 1550 4648 1556
rect 4272 1544 4284 1550
rect 4432 1544 4444 1550
rect 4636 1544 4648 1550
rect 3058 1458 3070 1464
rect 3098 1458 3110 1464
rect 3138 1458 3150 1464
rect 3223 1458 3235 1464
rect 3268 1458 3280 1464
rect 3378 1458 3390 1464
rect 3418 1458 3430 1464
rect 3458 1458 3470 1464
rect 3503 1458 3515 1464
rect 3631 1458 3643 1464
rect 3722 1458 3734 1464
rect 3772 1458 3784 1464
rect 3889 1458 3901 1464
rect 4007 1458 4019 1464
rect 4051 1458 4063 1464
rect 4263 1464 4291 1470
rect 4303 1536 4331 1542
rect 4423 1464 4451 1470
rect 4463 1536 4491 1542
rect 4589 1536 4617 1542
rect 4629 1464 4657 1470
rect 4757 1504 4765 1559
rect 4893 1544 4901 1579
rect 5011 1544 5019 1579
rect 4117 1458 4129 1464
rect 4157 1458 4169 1464
rect 4311 1458 4323 1464
rect 4471 1458 4483 1464
rect 4597 1458 4609 1464
rect 4737 1458 4749 1464
rect 4777 1458 4789 1464
rect 5054 1504 5062 1618
rect 5227 1637 5253 1643
rect 5459 1676 5471 1682
rect 5578 1676 5590 1682
rect 5771 1676 5783 1682
rect 5206 1618 5224 1620
rect 5194 1609 5224 1618
rect 5137 1597 5153 1603
rect 5137 1523 5143 1597
rect 5216 1581 5224 1609
rect 5257 1617 5273 1623
rect 5137 1517 5153 1523
rect 5218 1512 5225 1567
rect 5257 1527 5263 1617
rect 5333 1593 5340 1636
rect 5489 1628 5501 1636
rect 5477 1622 5501 1628
rect 5341 1556 5347 1579
rect 5477 1573 5485 1622
rect 5517 1617 5533 1623
rect 5341 1550 5368 1556
rect 5356 1544 5368 1550
rect 5178 1506 5225 1512
rect 5178 1504 5189 1506
rect 4862 1458 4874 1464
rect 4912 1458 4924 1464
rect 5027 1458 5039 1464
rect 5071 1458 5083 1464
rect 5217 1504 5225 1506
rect 5309 1536 5337 1542
rect 5349 1464 5377 1470
rect 5477 1504 5485 1559
rect 5517 1543 5523 1617
rect 5626 1618 5644 1620
rect 5614 1609 5644 1618
rect 5636 1581 5644 1609
rect 5756 1593 5764 1636
rect 5507 1537 5523 1543
rect 5638 1512 5645 1567
rect 5756 1544 5764 1579
rect 5598 1506 5645 1512
rect 5598 1504 5609 1506
rect 5157 1458 5169 1464
rect 5197 1458 5209 1464
rect 5317 1458 5329 1464
rect 5457 1458 5469 1464
rect 5497 1458 5509 1464
rect 5637 1504 5645 1506
rect 5577 1458 5589 1464
rect 5617 1458 5629 1464
rect 5771 1458 5783 1464
rect -62 1456 5816 1458
rect -62 1444 4 1456
rect -62 1442 2133 1444
rect -62 978 -2 1442
rect 91 1436 103 1442
rect 131 1436 143 1442
rect 217 1436 229 1442
rect 371 1436 383 1442
rect 411 1436 423 1442
rect 75 1394 83 1396
rect 111 1394 122 1396
rect 75 1388 122 1394
rect 75 1333 82 1388
rect 197 1362 209 1364
rect 197 1356 237 1362
rect 355 1394 363 1396
rect 496 1436 508 1442
rect 546 1436 558 1442
rect 391 1394 402 1396
rect 355 1388 402 1394
rect 258 1321 266 1356
rect 355 1333 362 1388
rect 636 1436 648 1442
rect 686 1436 698 1442
rect 807 1436 819 1442
rect 851 1436 863 1442
rect 917 1436 929 1442
rect 957 1436 969 1442
rect 1071 1436 1083 1442
rect 1137 1436 1149 1442
rect 1177 1436 1189 1442
rect 1277 1436 1289 1442
rect 1317 1436 1329 1442
rect 76 1291 84 1319
rect 76 1282 106 1291
rect 519 1321 527 1356
rect 659 1321 667 1356
rect 791 1321 799 1356
rect 76 1280 94 1282
rect 258 1264 266 1307
rect 356 1291 364 1319
rect 356 1282 386 1291
rect 513 1285 521 1307
rect 653 1285 661 1307
rect 791 1307 793 1321
rect 356 1280 374 1282
rect 130 1218 142 1224
rect 240 1253 266 1264
rect 495 1278 520 1285
rect 635 1278 660 1285
rect 495 1264 503 1278
rect 511 1264 563 1267
rect 635 1264 643 1278
rect 523 1258 551 1264
rect 651 1264 703 1267
rect 663 1258 691 1264
rect 791 1264 799 1307
rect 834 1282 842 1396
rect 937 1341 945 1396
rect 825 1274 863 1282
rect 851 1264 863 1274
rect 937 1278 945 1327
rect 1056 1313 1064 1396
rect 1158 1394 1169 1396
rect 1411 1436 1423 1442
rect 1451 1436 1463 1442
rect 1531 1436 1543 1442
rect 1571 1436 1583 1442
rect 1691 1436 1703 1442
rect 1731 1436 1743 1442
rect 1197 1394 1205 1396
rect 1158 1388 1205 1394
rect 1198 1333 1205 1388
rect 1297 1341 1305 1396
rect 1435 1341 1443 1396
rect 1555 1341 1563 1396
rect 1675 1394 1683 1396
rect 1797 1436 1809 1442
rect 1837 1436 1849 1442
rect 1951 1436 1963 1442
rect 1991 1436 2003 1442
rect 2091 1436 2103 1442
rect 1711 1394 1722 1396
rect 1675 1388 1722 1394
rect 937 1272 961 1278
rect 949 1264 961 1272
rect 791 1254 801 1264
rect 1056 1244 1064 1299
rect 1196 1291 1204 1319
rect 200 1218 212 1224
rect 250 1218 262 1224
rect 410 1218 422 1224
rect 531 1218 543 1224
rect 671 1218 683 1224
rect 821 1218 833 1224
rect 919 1218 931 1224
rect 1071 1218 1083 1224
rect 1174 1282 1204 1291
rect 1186 1280 1204 1282
rect 1297 1278 1305 1327
rect 1435 1278 1443 1327
rect 1675 1333 1682 1388
rect 1817 1341 1825 1396
rect 1935 1394 1943 1396
rect 2147 1442 3233 1444
rect 2211 1436 2223 1442
rect 2251 1436 2263 1442
rect 2351 1436 2363 1442
rect 2391 1436 2403 1442
rect 1971 1394 1982 1396
rect 1935 1388 1982 1394
rect 1555 1278 1563 1327
rect 1935 1333 1942 1388
rect 1676 1291 1684 1319
rect 1676 1282 1706 1291
rect 1676 1280 1694 1282
rect 1297 1272 1321 1278
rect 1309 1264 1321 1272
rect 1419 1272 1443 1278
rect 1539 1272 1563 1278
rect 1419 1264 1431 1272
rect 1539 1264 1551 1272
rect 1817 1278 1825 1327
rect 1936 1291 1944 1319
rect 2076 1313 2084 1396
rect 2195 1394 2203 1396
rect 2231 1394 2242 1396
rect 2195 1388 2242 1394
rect 2335 1394 2343 1396
rect 2457 1436 2469 1442
rect 2596 1436 2608 1442
rect 2646 1436 2658 1442
rect 2737 1436 2749 1442
rect 2876 1436 2888 1442
rect 2926 1436 2938 1442
rect 2371 1394 2382 1396
rect 2335 1388 2382 1394
rect 2195 1333 2202 1388
rect 2335 1333 2342 1388
rect 1936 1282 1966 1291
rect 1936 1280 1954 1282
rect 1817 1272 1841 1278
rect 1829 1264 1841 1272
rect 1138 1218 1150 1224
rect 1279 1218 1291 1224
rect 1449 1218 1461 1224
rect 1569 1218 1581 1224
rect 1730 1218 1742 1224
rect 2076 1244 2084 1299
rect 2196 1291 2204 1319
rect 2336 1291 2344 1319
rect 2476 1313 2484 1396
rect 2717 1362 2729 1364
rect 2717 1356 2757 1362
rect 2619 1321 2627 1356
rect 2778 1321 2786 1356
rect 2196 1282 2226 1291
rect 2196 1280 2214 1282
rect 2336 1282 2366 1291
rect 2336 1280 2354 1282
rect 2476 1244 2484 1299
rect 2613 1285 2621 1307
rect 2595 1278 2620 1285
rect 2595 1264 2603 1278
rect 1799 1218 1811 1224
rect 1990 1218 2002 1224
rect 2091 1218 2103 1224
rect 2250 1218 2262 1224
rect 2390 1218 2402 1224
rect 2611 1264 2663 1267
rect 2778 1264 2786 1307
rect 2857 1283 2863 1373
rect 3016 1436 3028 1442
rect 3066 1436 3078 1442
rect 3156 1436 3168 1442
rect 3206 1436 3218 1442
rect 3247 1442 5816 1444
rect 3311 1436 3323 1442
rect 3377 1436 3389 1442
rect 3509 1436 3521 1442
rect 3671 1436 3683 1442
rect 3762 1436 3774 1442
rect 3812 1436 3824 1442
rect 3931 1436 3943 1442
rect 2899 1321 2907 1356
rect 3039 1321 3047 1356
rect 3179 1321 3187 1356
rect 2893 1285 2901 1307
rect 3033 1285 3041 1307
rect 3173 1285 3181 1307
rect 3296 1313 3304 1396
rect 3396 1313 3404 1396
rect 3491 1321 3499 1356
rect 3535 1350 3543 1396
rect 3691 1362 3703 1364
rect 3663 1356 3703 1362
rect 4016 1436 4028 1442
rect 4066 1436 4078 1442
rect 3517 1344 3543 1350
rect 3517 1338 3520 1344
rect 2847 1277 2863 1283
rect 2875 1278 2900 1285
rect 3015 1278 3040 1285
rect 3155 1278 3180 1285
rect 2875 1264 2883 1278
rect 2623 1258 2651 1264
rect 2760 1253 2786 1264
rect 2891 1264 2943 1267
rect 3015 1264 3023 1278
rect 2903 1258 2931 1264
rect 3031 1264 3083 1267
rect 3155 1264 3163 1278
rect 3043 1258 3071 1264
rect 3171 1264 3223 1267
rect 3183 1258 3211 1264
rect 3296 1244 3304 1299
rect 3491 1307 3493 1321
rect 3396 1244 3404 1299
rect 3491 1264 3499 1307
rect 3513 1282 3520 1338
rect 3634 1321 3642 1356
rect 3667 1337 3713 1343
rect 3793 1321 3801 1356
rect 3517 1276 3520 1282
rect 3517 1270 3539 1276
rect 2457 1218 2469 1224
rect 2631 1218 2643 1224
rect 2720 1218 2732 1224
rect 2770 1218 2782 1224
rect 2911 1218 2923 1224
rect 3051 1218 3063 1224
rect 3191 1218 3203 1224
rect 3311 1218 3323 1224
rect 3531 1244 3539 1270
rect 3634 1264 3642 1307
rect 3916 1313 3924 1396
rect 4156 1436 4168 1442
rect 4206 1436 4218 1442
rect 4331 1436 4343 1442
rect 4436 1436 4448 1442
rect 4486 1436 4498 1442
rect 4351 1362 4363 1364
rect 4323 1356 4363 1362
rect 4582 1436 4594 1442
rect 4632 1436 4644 1442
rect 4717 1436 4729 1442
rect 4757 1436 4769 1442
rect 4842 1436 4854 1442
rect 4892 1436 4904 1442
rect 4039 1321 4047 1356
rect 4179 1321 4187 1356
rect 4294 1321 4302 1356
rect 4459 1321 4467 1356
rect 4613 1321 4621 1356
rect 4737 1341 4745 1396
rect 4977 1436 4989 1442
rect 5097 1436 5109 1442
rect 5137 1436 5149 1442
rect 5231 1436 5243 1442
rect 5271 1436 5283 1442
rect 5356 1436 5368 1442
rect 5406 1436 5418 1442
rect 3799 1285 3807 1307
rect 3800 1278 3825 1285
rect 3757 1264 3809 1267
rect 3634 1253 3660 1264
rect 3769 1258 3797 1264
rect 3817 1264 3825 1278
rect 3916 1244 3924 1299
rect 4033 1285 4041 1307
rect 4173 1285 4181 1307
rect 4015 1278 4040 1285
rect 4155 1278 4180 1285
rect 4015 1264 4023 1278
rect 4031 1264 4083 1267
rect 4155 1264 4163 1278
rect 4043 1258 4071 1264
rect 4171 1264 4223 1267
rect 4183 1258 4211 1264
rect 4294 1264 4302 1307
rect 4453 1285 4461 1307
rect 4619 1285 4627 1307
rect 4435 1278 4460 1285
rect 4620 1278 4645 1285
rect 4435 1264 4443 1278
rect 4294 1253 4320 1264
rect 4451 1264 4503 1267
rect 4463 1258 4491 1264
rect 4577 1264 4629 1267
rect 4589 1258 4617 1264
rect 4637 1264 4645 1278
rect 4737 1278 4745 1327
rect 4873 1321 4881 1356
rect 5000 1349 5017 1356
rect 4879 1285 4887 1307
rect 5000 1301 5007 1349
rect 5117 1341 5125 1396
rect 5255 1341 5263 1396
rect 5482 1436 5494 1442
rect 5532 1436 5544 1442
rect 5642 1436 5654 1442
rect 5692 1436 5704 1442
rect 4880 1278 4905 1285
rect 4737 1272 4761 1278
rect 4749 1264 4761 1272
rect 4837 1264 4889 1267
rect 4849 1258 4877 1264
rect 4897 1264 4905 1278
rect 5000 1244 5007 1287
rect 5117 1278 5125 1327
rect 5255 1278 5263 1327
rect 5379 1321 5387 1356
rect 5513 1321 5521 1356
rect 5673 1321 5681 1356
rect 5373 1285 5381 1307
rect 5519 1285 5527 1307
rect 5679 1285 5687 1307
rect 5117 1272 5141 1278
rect 5129 1264 5141 1272
rect 3377 1218 3389 1224
rect 3509 1218 3521 1224
rect 3638 1218 3650 1224
rect 3688 1218 3700 1224
rect 3777 1218 3789 1224
rect 3931 1218 3943 1224
rect 4051 1218 4063 1224
rect 4191 1218 4203 1224
rect 4298 1218 4310 1224
rect 4348 1218 4360 1224
rect 4471 1218 4483 1224
rect 4597 1218 4609 1224
rect 4719 1218 4731 1224
rect 4857 1218 4869 1224
rect 4977 1218 4989 1224
rect 5017 1218 5029 1224
rect 5239 1272 5263 1278
rect 5355 1278 5380 1285
rect 5520 1278 5545 1285
rect 5680 1278 5705 1285
rect 5239 1264 5251 1272
rect 5355 1264 5363 1278
rect 5371 1264 5423 1267
rect 5383 1258 5411 1264
rect 5477 1264 5529 1267
rect 5489 1258 5517 1264
rect 5537 1264 5545 1278
rect 5637 1264 5689 1267
rect 5649 1258 5677 1264
rect 5697 1264 5705 1278
rect 5099 1218 5111 1224
rect 5269 1218 5281 1224
rect 5391 1218 5403 1224
rect 5497 1218 5509 1224
rect 5657 1218 5669 1224
rect 5822 1218 5882 1682
rect 4 1216 5882 1218
rect 5816 1204 5882 1216
rect 4 1202 5882 1204
rect 91 1196 103 1202
rect 160 1196 172 1202
rect 210 1196 222 1202
rect 317 1196 329 1202
rect 457 1196 469 1202
rect 650 1196 662 1202
rect 737 1196 749 1202
rect 880 1196 892 1202
rect 930 1196 942 1202
rect 1071 1196 1083 1202
rect 1191 1196 1203 1202
rect 76 1121 84 1176
rect 200 1156 226 1167
rect 218 1113 226 1156
rect 309 1156 337 1162
rect 297 1153 349 1156
rect 449 1156 477 1162
rect 357 1142 365 1156
rect 437 1153 489 1156
rect 497 1142 505 1156
rect 340 1135 365 1142
rect 480 1135 505 1142
rect 596 1138 614 1140
rect 76 1024 84 1107
rect 339 1113 347 1135
rect 479 1113 487 1135
rect 596 1129 626 1138
rect 729 1156 757 1162
rect 717 1153 769 1156
rect 920 1156 946 1167
rect 777 1142 785 1156
rect 760 1135 785 1142
rect 596 1101 604 1129
rect 218 1064 226 1099
rect 333 1064 341 1099
rect 473 1064 481 1099
rect 759 1113 767 1135
rect 938 1113 946 1156
rect 1035 1142 1043 1156
rect 1063 1156 1091 1162
rect 1260 1196 1272 1202
rect 1310 1196 1322 1202
rect 1431 1196 1443 1202
rect 1051 1153 1103 1156
rect 1035 1135 1060 1142
rect 1053 1113 1061 1135
rect 1176 1121 1184 1176
rect 1511 1196 1523 1202
rect 1551 1196 1563 1202
rect 1637 1196 1649 1202
rect 1810 1196 1822 1202
rect 1929 1196 1941 1202
rect 2051 1196 2063 1202
rect 2210 1196 2222 1202
rect 2350 1196 2362 1202
rect 2471 1196 2483 1202
rect 2630 1196 2642 1202
rect 1300 1156 1326 1167
rect 1318 1113 1326 1156
rect 1416 1121 1424 1176
rect 1533 1133 1540 1176
rect 157 1058 197 1064
rect 157 1056 169 1058
rect 91 978 103 984
rect 177 978 189 984
rect 302 978 314 984
rect 352 978 364 984
rect 595 1032 602 1087
rect 753 1064 761 1099
rect 938 1064 946 1099
rect 1059 1064 1067 1099
rect 1127 1077 1153 1083
rect 595 1026 642 1032
rect 595 1024 603 1026
rect 631 1024 642 1026
rect 442 978 454 984
rect 492 978 504 984
rect 611 978 623 984
rect 651 978 663 984
rect 877 1058 917 1064
rect 877 1056 889 1058
rect 1176 1024 1184 1107
rect 1656 1121 1664 1176
rect 1756 1138 1774 1140
rect 1756 1129 1786 1138
rect 1899 1148 1911 1156
rect 1899 1142 1923 1148
rect 1318 1064 1326 1099
rect 1257 1058 1297 1064
rect 1257 1056 1269 1058
rect 1416 1024 1424 1107
rect 1533 1071 1540 1119
rect 1523 1064 1540 1071
rect 1656 1024 1664 1107
rect 1756 1101 1764 1129
rect 1827 1117 1853 1123
rect 1755 1032 1762 1087
rect 1915 1093 1923 1142
rect 2015 1142 2023 1156
rect 2043 1156 2071 1162
rect 2031 1153 2083 1156
rect 2015 1135 2040 1142
rect 2156 1138 2174 1140
rect 2033 1113 2041 1135
rect 2156 1129 2186 1138
rect 2296 1138 2314 1140
rect 2296 1129 2326 1138
rect 2435 1142 2443 1156
rect 2463 1156 2491 1162
rect 2451 1153 2503 1156
rect 2435 1135 2460 1142
rect 2576 1138 2594 1140
rect 2156 1101 2164 1129
rect 2296 1101 2304 1129
rect 2453 1113 2461 1135
rect 2576 1129 2606 1138
rect 2717 1196 2729 1202
rect 2817 1196 2829 1202
rect 2857 1196 2869 1202
rect 2937 1196 2949 1202
rect 2977 1196 2989 1202
rect 3087 1196 3099 1202
rect 3211 1196 3223 1202
rect 3251 1196 3263 1202
rect 1755 1026 1802 1032
rect 1755 1024 1763 1026
rect 722 978 734 984
rect 772 978 784 984
rect 897 978 909 984
rect 1036 978 1048 984
rect 1086 978 1098 984
rect 1191 978 1203 984
rect 1277 978 1289 984
rect 1431 978 1443 984
rect 1551 978 1563 984
rect 1791 1024 1802 1026
rect 1915 1024 1923 1079
rect 2039 1064 2047 1099
rect 1637 978 1649 984
rect 1771 978 1783 984
rect 1811 978 1823 984
rect 1891 978 1903 984
rect 1931 978 1943 984
rect 2155 1032 2162 1087
rect 2576 1101 2584 1129
rect 2736 1121 2744 1176
rect 2840 1133 2847 1176
rect 2960 1133 2967 1176
rect 3351 1196 3363 1202
rect 3391 1196 3403 1202
rect 3491 1196 3503 1202
rect 3611 1196 3623 1202
rect 3751 1196 3763 1202
rect 3839 1196 3851 1202
rect 3959 1196 3971 1202
rect 4077 1196 4089 1202
rect 4117 1196 4129 1202
rect 3119 1156 3129 1166
rect 3057 1146 3069 1156
rect 3057 1138 3095 1146
rect 2295 1032 2302 1087
rect 2459 1064 2467 1099
rect 2155 1026 2202 1032
rect 2155 1024 2163 1026
rect 2191 1024 2202 1026
rect 2295 1026 2342 1032
rect 2295 1024 2303 1026
rect 2331 1024 2342 1026
rect 2016 978 2028 984
rect 2066 978 2078 984
rect 2171 978 2183 984
rect 2211 978 2223 984
rect 2311 978 2323 984
rect 2351 978 2363 984
rect 2575 1032 2582 1087
rect 2575 1026 2622 1032
rect 2575 1024 2583 1026
rect 2611 1024 2622 1026
rect 2736 1024 2744 1107
rect 2840 1071 2847 1119
rect 2960 1071 2967 1119
rect 2840 1064 2857 1071
rect 2960 1064 2977 1071
rect 2436 978 2448 984
rect 2486 978 2498 984
rect 2591 978 2603 984
rect 2631 978 2643 984
rect 3078 1024 3086 1138
rect 3121 1113 3129 1156
rect 3233 1133 3240 1176
rect 3373 1133 3380 1176
rect 3476 1121 3484 1176
rect 3575 1142 3583 1156
rect 3603 1156 3631 1162
rect 3591 1153 3643 1156
rect 3715 1142 3723 1156
rect 3743 1156 3771 1162
rect 4197 1196 4209 1202
rect 4318 1196 4330 1202
rect 4368 1196 4380 1202
rect 4511 1196 4523 1202
rect 4618 1196 4630 1202
rect 4668 1196 4680 1202
rect 4757 1196 4769 1202
rect 4899 1196 4911 1202
rect 4997 1196 5009 1202
rect 5097 1196 5109 1202
rect 5249 1196 5261 1202
rect 5391 1196 5403 1202
rect 5477 1196 5489 1202
rect 5517 1196 5529 1202
rect 5670 1196 5682 1202
rect 5771 1196 5783 1202
rect 3731 1153 3783 1156
rect 3869 1148 3881 1156
rect 3989 1148 4001 1156
rect 3575 1135 3600 1142
rect 3715 1135 3740 1142
rect 3127 1099 3129 1113
rect 3121 1064 3129 1099
rect 3233 1071 3240 1119
rect 3373 1071 3380 1119
rect 3593 1113 3601 1135
rect 3223 1064 3240 1071
rect 3363 1064 3380 1071
rect 3476 1024 3484 1107
rect 3733 1113 3741 1135
rect 3857 1142 3881 1148
rect 3977 1142 4001 1148
rect 3599 1064 3607 1099
rect 3739 1064 3747 1099
rect 3797 1067 3803 1133
rect 3857 1093 3865 1142
rect 3977 1093 3985 1142
rect 4100 1133 4107 1176
rect 4216 1121 4224 1176
rect 4314 1156 4340 1167
rect 2717 978 2729 984
rect 2817 978 2829 984
rect 2937 978 2949 984
rect 3057 978 3069 984
rect 3101 978 3113 984
rect 3251 978 3263 984
rect 3391 978 3403 984
rect 3491 978 3503 984
rect 3576 978 3588 984
rect 3626 978 3638 984
rect 3857 1024 3865 1079
rect 3977 1024 3985 1079
rect 4100 1071 4107 1119
rect 4314 1113 4322 1156
rect 4475 1142 4483 1156
rect 4503 1156 4531 1162
rect 4491 1153 4543 1156
rect 4614 1156 4640 1167
rect 4749 1156 4777 1162
rect 4475 1135 4500 1142
rect 4100 1064 4117 1071
rect 3716 978 3728 984
rect 3766 978 3778 984
rect 3837 978 3849 984
rect 3877 978 3889 984
rect 3957 978 3969 984
rect 3997 978 4009 984
rect 4216 1024 4224 1107
rect 4493 1113 4501 1135
rect 4614 1113 4622 1156
rect 4737 1153 4789 1156
rect 4797 1142 4805 1156
rect 4881 1150 4889 1176
rect 4881 1144 4903 1150
rect 4780 1135 4805 1142
rect 4900 1138 4903 1144
rect 4779 1113 4787 1135
rect 4314 1064 4322 1099
rect 4499 1064 4507 1099
rect 4614 1064 4622 1099
rect 4647 1077 4713 1083
rect 4773 1064 4781 1099
rect 4900 1082 4907 1138
rect 4921 1113 4929 1156
rect 5016 1121 5024 1176
rect 4927 1099 4929 1113
rect 5116 1121 5124 1176
rect 5219 1148 5231 1156
rect 5219 1142 5243 1148
rect 4900 1076 4903 1082
rect 4877 1070 4903 1076
rect 4343 1058 4383 1064
rect 4371 1056 4383 1058
rect 4643 1058 4683 1064
rect 4671 1056 4683 1058
rect 4877 1024 4885 1070
rect 4921 1064 4929 1099
rect 5016 1024 5024 1107
rect 5116 1024 5124 1107
rect 5235 1093 5243 1142
rect 5355 1142 5363 1156
rect 5383 1156 5411 1162
rect 5371 1153 5423 1156
rect 5355 1135 5380 1142
rect 5373 1113 5381 1135
rect 5500 1133 5507 1176
rect 5235 1024 5243 1079
rect 5379 1064 5387 1099
rect 5500 1071 5507 1119
rect 5616 1138 5634 1140
rect 5616 1129 5646 1138
rect 5616 1101 5624 1129
rect 5687 1117 5703 1123
rect 5756 1121 5764 1176
rect 5500 1064 5517 1071
rect 4077 978 4089 984
rect 4197 978 4209 984
rect 4351 978 4363 984
rect 4476 978 4488 984
rect 4526 978 4538 984
rect 4651 978 4663 984
rect 4742 978 4754 984
rect 4792 978 4804 984
rect 4899 978 4911 984
rect 4997 978 5009 984
rect 5097 978 5109 984
rect 5211 978 5223 984
rect 5251 978 5263 984
rect 5356 978 5368 984
rect 5406 978 5418 984
rect 5615 1032 5622 1087
rect 5697 1087 5703 1117
rect 5615 1026 5662 1032
rect 5615 1024 5623 1026
rect 5651 1024 5662 1026
rect 5756 1024 5764 1107
rect 5477 978 5489 984
rect 5631 978 5643 984
rect 5671 978 5683 984
rect 5771 978 5783 984
rect -62 976 5816 978
rect -62 964 4 976
rect -62 962 5816 964
rect -62 498 -2 962
rect 91 956 103 962
rect 131 956 143 962
rect 217 956 229 962
rect 371 956 383 962
rect 411 956 423 962
rect 531 956 543 962
rect 651 956 663 962
rect 691 956 703 962
rect 777 956 789 962
rect 916 956 928 962
rect 966 956 978 962
rect 1071 956 1083 962
rect 1111 956 1123 962
rect 75 914 83 916
rect 111 914 122 916
rect 75 908 122 914
rect 75 853 82 908
rect 197 882 209 884
rect 197 876 237 882
rect 355 914 363 916
rect 391 914 402 916
rect 355 908 402 914
rect 258 841 266 876
rect 355 853 362 908
rect 551 882 563 884
rect 523 876 563 882
rect 635 914 643 916
rect 671 914 682 916
rect 635 908 682 914
rect 76 811 84 839
rect 76 802 106 811
rect 494 841 502 876
rect 635 853 642 908
rect 757 882 769 884
rect 757 876 797 882
rect 1055 914 1063 916
rect 1182 956 1194 962
rect 1232 956 1244 962
rect 1351 956 1363 962
rect 1391 956 1403 962
rect 1091 914 1102 916
rect 1055 908 1102 914
rect 76 800 94 802
rect 258 784 266 827
rect 356 811 364 839
rect 818 841 826 876
rect 939 841 947 876
rect 1055 853 1062 908
rect 1335 914 1343 916
rect 1457 956 1469 962
rect 1557 956 1569 962
rect 1597 956 1609 962
rect 1731 956 1743 962
rect 1771 956 1783 962
rect 1871 956 1883 962
rect 1911 956 1923 962
rect 1371 914 1382 916
rect 1335 908 1382 914
rect 356 802 386 811
rect 356 800 374 802
rect 130 738 142 744
rect 240 773 266 784
rect 494 784 502 827
rect 636 811 644 839
rect 636 802 666 811
rect 636 800 654 802
rect 494 773 520 784
rect 200 738 212 744
rect 250 738 262 744
rect 410 738 422 744
rect 818 784 826 827
rect 933 805 941 827
rect 1213 841 1221 876
rect 1335 853 1342 908
rect 1056 811 1064 839
rect 915 798 940 805
rect 1056 802 1086 811
rect 1056 800 1074 802
rect 915 784 923 798
rect 498 738 510 744
rect 548 738 560 744
rect 690 738 702 744
rect 800 773 826 784
rect 931 784 983 787
rect 943 778 971 784
rect 1147 797 1173 803
rect 1219 805 1227 827
rect 1336 811 1344 839
rect 1476 833 1484 916
rect 1577 861 1585 916
rect 1715 914 1723 916
rect 1751 914 1762 916
rect 1715 908 1762 914
rect 1855 914 1863 916
rect 1977 956 1989 962
rect 2017 956 2029 962
rect 2122 956 2134 962
rect 2172 956 2184 962
rect 1891 914 1902 916
rect 1855 908 1902 914
rect 1998 914 2009 916
rect 2037 914 2045 916
rect 1998 908 2045 914
rect 1607 877 1653 883
rect 1715 853 1722 908
rect 1220 798 1245 805
rect 1336 802 1366 811
rect 1336 800 1354 802
rect 1177 784 1229 787
rect 1189 778 1217 784
rect 1237 784 1245 798
rect 1476 764 1484 819
rect 1577 798 1585 847
rect 1855 853 1862 908
rect 2038 853 2045 908
rect 2257 956 2269 962
rect 2301 956 2313 962
rect 2397 956 2409 962
rect 2511 956 2523 962
rect 2551 956 2563 962
rect 2661 956 2673 962
rect 2757 956 2769 962
rect 2797 956 2809 962
rect 2153 841 2161 876
rect 1716 811 1724 839
rect 1856 811 1864 839
rect 2036 811 2044 839
rect 1716 802 1746 811
rect 1716 800 1734 802
rect 1577 792 1601 798
rect 1589 784 1601 792
rect 760 738 772 744
rect 810 738 822 744
rect 951 738 963 744
rect 1110 738 1122 744
rect 1197 738 1209 744
rect 1390 738 1402 744
rect 1856 802 1886 811
rect 1856 800 1874 802
rect 1457 738 1469 744
rect 1559 738 1571 744
rect 1770 738 1782 744
rect 1910 738 1922 744
rect 2014 802 2044 811
rect 2159 805 2167 827
rect 2026 800 2044 802
rect 2160 798 2185 805
rect 2278 802 2286 916
rect 2321 841 2329 876
rect 2327 827 2329 841
rect 2416 833 2424 916
rect 2535 861 2543 916
rect 2637 877 2641 886
rect 2117 784 2169 787
rect 2129 778 2157 784
rect 2177 784 2185 798
rect 2257 794 2295 802
rect 2257 784 2269 794
rect 2321 784 2329 827
rect 2319 774 2329 784
rect 2416 764 2424 819
rect 2535 798 2543 847
rect 2637 833 2646 877
rect 2891 956 2903 962
rect 2931 956 2943 962
rect 3017 956 3029 962
rect 3151 956 3163 962
rect 3251 956 3263 962
rect 3291 956 3303 962
rect 3431 956 3443 962
rect 3551 956 3563 962
rect 3671 956 3683 962
rect 3791 956 3803 962
rect 2695 868 2703 876
rect 2667 860 2703 868
rect 2777 861 2785 916
rect 2915 861 2923 916
rect 2519 792 2543 798
rect 2519 784 2531 792
rect 2633 784 2640 819
rect 2656 804 2662 859
rect 2777 798 2785 847
rect 2915 798 2923 847
rect 3036 833 3044 916
rect 3136 833 3144 916
rect 3275 861 3283 916
rect 3876 956 3888 962
rect 3926 956 3938 962
rect 3691 882 3703 884
rect 3663 876 3703 882
rect 3403 869 3420 876
rect 3523 869 3540 876
rect 2667 792 2677 798
rect 2777 792 2801 798
rect 2671 764 2677 792
rect 2789 784 2801 792
rect 1978 738 1990 744
rect 2137 738 2149 744
rect 2287 738 2299 744
rect 2397 738 2409 744
rect 2549 738 2561 744
rect 2651 738 2663 744
rect 2695 738 2703 744
rect 2899 792 2923 798
rect 2899 784 2911 792
rect 3036 764 3044 819
rect 3136 764 3144 819
rect 3275 798 3283 847
rect 3259 792 3283 798
rect 3413 821 3420 869
rect 3533 821 3540 869
rect 3634 841 3642 876
rect 3776 833 3784 916
rect 3817 877 3853 883
rect 3259 784 3271 792
rect 2759 738 2771 744
rect 2929 738 2941 744
rect 3413 764 3420 807
rect 3533 764 3540 807
rect 3634 784 3642 827
rect 3634 773 3660 784
rect 3017 738 3029 744
rect 3151 738 3163 744
rect 3289 738 3301 744
rect 3391 738 3403 744
rect 3431 738 3443 744
rect 3511 738 3523 744
rect 3551 738 3563 744
rect 3776 764 3784 819
rect 3817 783 3823 877
rect 3997 956 4009 962
rect 4037 956 4049 962
rect 4136 956 4148 962
rect 4186 956 4198 962
rect 3899 841 3907 876
rect 4017 861 4025 916
rect 4276 956 4288 962
rect 4326 956 4338 962
rect 4417 956 4429 962
rect 4536 956 4548 962
rect 4586 956 4598 962
rect 4677 956 4689 962
rect 4829 956 4841 962
rect 4936 956 4948 962
rect 4986 956 4998 962
rect 5077 956 5089 962
rect 5241 956 5253 962
rect 5391 956 5403 962
rect 5531 956 5543 962
rect 5642 956 5654 962
rect 5692 956 5704 962
rect 3893 805 3901 827
rect 3875 798 3900 805
rect 4017 798 4025 847
rect 4159 841 4167 876
rect 4299 841 4307 876
rect 4153 805 4161 827
rect 4293 805 4301 827
rect 4436 833 4444 916
rect 4657 882 4669 884
rect 4657 876 4697 882
rect 4559 841 4567 876
rect 4718 841 4726 876
rect 4811 841 4819 876
rect 4855 870 4863 916
rect 5057 882 5069 884
rect 5057 876 5097 882
rect 5217 877 5221 886
rect 4837 864 4863 870
rect 4837 858 4840 864
rect 4135 798 4160 805
rect 4275 798 4300 805
rect 3875 784 3883 798
rect 4017 792 4041 798
rect 3807 777 3823 783
rect 3891 784 3943 787
rect 4029 784 4041 792
rect 4135 784 4143 798
rect 3903 778 3931 784
rect 4151 784 4203 787
rect 4275 784 4283 798
rect 4163 778 4191 784
rect 4291 784 4343 787
rect 4303 778 4331 784
rect 4436 764 4444 819
rect 4553 805 4561 827
rect 4811 827 4813 841
rect 4535 798 4560 805
rect 4535 784 4543 798
rect 4551 784 4603 787
rect 4718 784 4726 827
rect 4811 784 4819 827
rect 4833 802 4840 858
rect 4959 841 4967 876
rect 5047 857 5093 863
rect 5118 841 5126 876
rect 4953 805 4961 827
rect 5217 833 5226 877
rect 5275 868 5283 876
rect 5247 860 5283 868
rect 4837 796 4840 802
rect 4935 798 4960 805
rect 4837 790 4859 796
rect 4563 778 4591 784
rect 4700 773 4726 784
rect 4851 764 4859 790
rect 4935 784 4943 798
rect 4951 784 5003 787
rect 5118 784 5126 827
rect 5213 784 5220 819
rect 5236 804 5242 859
rect 5376 833 5384 916
rect 5483 950 5511 956
rect 5523 878 5551 884
rect 5492 870 5504 876
rect 5492 864 5519 870
rect 5513 841 5519 864
rect 5673 841 5681 876
rect 5247 792 5257 798
rect 4963 778 4991 784
rect 5100 773 5126 784
rect 5251 764 5257 792
rect 5376 764 5384 819
rect 5520 784 5527 827
rect 5679 805 5687 827
rect 5680 798 5705 805
rect 5637 784 5689 787
rect 3638 738 3650 744
rect 3688 738 3700 744
rect 3791 738 3803 744
rect 3911 738 3923 744
rect 3999 738 4011 744
rect 4171 738 4183 744
rect 4311 738 4323 744
rect 4417 738 4429 744
rect 4571 738 4583 744
rect 4660 738 4672 744
rect 4710 738 4722 744
rect 4829 738 4841 744
rect 4971 738 4983 744
rect 5060 738 5072 744
rect 5110 738 5122 744
rect 5231 738 5243 744
rect 5275 738 5283 744
rect 5391 738 5403 744
rect 5649 778 5677 784
rect 5697 784 5705 798
rect 5492 738 5504 744
rect 5548 738 5560 744
rect 5657 738 5669 744
rect 5822 738 5882 1202
rect 4 736 5882 738
rect 5816 724 5882 736
rect 4 722 5882 724
rect 130 716 142 722
rect 76 658 94 660
rect 76 649 106 658
rect 238 716 250 722
rect 288 716 300 722
rect 430 716 442 722
rect 551 716 563 722
rect 640 716 652 722
rect 690 716 702 722
rect 234 676 260 687
rect 76 621 84 649
rect 234 633 242 676
rect 376 658 394 660
rect 376 649 406 658
rect 515 662 523 676
rect 543 676 571 682
rect 779 716 791 722
rect 971 716 983 722
rect 1130 716 1142 722
rect 680 676 706 687
rect 531 673 583 676
rect 515 655 540 662
rect 376 621 384 649
rect 533 633 541 655
rect 75 552 82 607
rect 234 584 242 619
rect 698 633 706 676
rect 809 668 821 676
rect 797 662 821 668
rect 935 662 943 676
rect 963 676 991 682
rect 951 673 1003 676
rect 75 546 122 552
rect 75 544 83 546
rect 111 544 122 546
rect 263 578 303 584
rect 291 576 303 578
rect 375 552 382 607
rect 539 584 547 619
rect 698 584 706 619
rect 797 613 805 662
rect 935 655 960 662
rect 1076 658 1094 660
rect 953 633 961 655
rect 1076 649 1106 658
rect 1200 716 1212 722
rect 1250 716 1262 722
rect 1358 716 1370 722
rect 1408 716 1420 722
rect 1240 676 1266 687
rect 1076 621 1084 649
rect 1258 633 1266 676
rect 1354 676 1380 687
rect 1498 716 1510 722
rect 1691 716 1703 722
rect 1850 716 1862 722
rect 1354 633 1362 676
rect 1655 662 1663 676
rect 1683 676 1711 682
rect 1671 673 1723 676
rect 1546 658 1564 660
rect 375 546 422 552
rect 375 544 383 546
rect 411 544 422 546
rect 91 498 103 504
rect 131 498 143 504
rect 271 498 283 504
rect 391 498 403 504
rect 431 498 443 504
rect 637 578 677 584
rect 637 576 649 578
rect 797 544 805 599
rect 959 584 967 619
rect 1534 649 1564 658
rect 1655 655 1680 662
rect 1796 658 1814 660
rect 1556 621 1564 649
rect 1673 633 1681 655
rect 1796 649 1826 658
rect 1920 716 1932 722
rect 1970 716 1982 722
rect 2071 716 2083 722
rect 2111 716 2123 722
rect 2211 716 2223 722
rect 2255 716 2263 722
rect 2347 716 2359 722
rect 2459 716 2471 722
rect 2629 716 2641 722
rect 1960 676 1986 687
rect 516 498 528 504
rect 566 498 578 504
rect 657 498 669 504
rect 777 498 789 504
rect 817 498 829 504
rect 1075 552 1082 607
rect 1258 584 1266 619
rect 1354 584 1362 619
rect 1796 621 1804 649
rect 1978 633 1986 676
rect 2093 653 2100 696
rect 2193 641 2200 676
rect 2231 668 2237 696
rect 2227 662 2237 668
rect 2379 676 2389 686
rect 2317 666 2329 676
rect 2317 658 2355 666
rect 1197 578 1237 584
rect 1197 576 1209 578
rect 1075 546 1122 552
rect 1075 544 1083 546
rect 1111 544 1122 546
rect 1383 578 1423 584
rect 1411 576 1423 578
rect 1558 552 1565 607
rect 1679 584 1687 619
rect 1518 546 1565 552
rect 1518 544 1529 546
rect 1557 544 1565 546
rect 1795 552 1802 607
rect 1978 584 1986 619
rect 2093 591 2100 639
rect 2083 584 2100 591
rect 1917 578 1957 584
rect 1917 576 1929 578
rect 1795 546 1842 552
rect 1795 544 1803 546
rect 1831 544 1842 546
rect 2197 583 2206 627
rect 2216 601 2222 656
rect 2227 592 2263 600
rect 2255 584 2263 592
rect 2197 574 2201 583
rect 2338 544 2346 658
rect 2381 633 2389 676
rect 2489 668 2501 676
rect 2477 662 2501 668
rect 2711 716 2723 722
rect 2751 716 2763 722
rect 2837 716 2849 722
rect 3009 716 3021 722
rect 2599 668 2611 676
rect 2599 662 2623 668
rect 2387 619 2389 633
rect 2381 584 2389 619
rect 2477 613 2485 662
rect 2615 613 2623 662
rect 2733 653 2740 696
rect 2829 676 2857 682
rect 2817 673 2869 676
rect 3080 716 3092 722
rect 3130 716 3142 722
rect 3290 716 3302 722
rect 3120 676 3146 687
rect 2877 662 2885 676
rect 2979 668 2991 676
rect 2979 662 3003 668
rect 2860 655 2885 662
rect 2477 544 2485 599
rect 2615 544 2623 599
rect 2733 591 2740 639
rect 2859 633 2867 655
rect 2723 584 2740 591
rect 2853 584 2861 619
rect 2995 613 3003 662
rect 3138 633 3146 676
rect 3236 658 3254 660
rect 3236 649 3266 658
rect 3359 716 3371 722
rect 3531 716 3543 722
rect 3619 716 3631 722
rect 3791 716 3803 722
rect 3897 716 3909 722
rect 4020 716 4032 722
rect 4070 716 4082 722
rect 4197 716 4209 722
rect 4351 716 4363 722
rect 3389 668 3401 676
rect 3377 662 3401 668
rect 3495 662 3503 676
rect 3523 676 3551 682
rect 3511 673 3563 676
rect 3649 668 3661 676
rect 3637 662 3661 668
rect 3755 662 3763 676
rect 3783 676 3811 682
rect 3771 673 3823 676
rect 3889 676 3917 682
rect 3877 673 3929 676
rect 4060 676 4086 687
rect 3236 621 3244 649
rect 3287 637 3313 643
rect 936 498 948 504
rect 986 498 998 504
rect 1091 498 1103 504
rect 1131 498 1143 504
rect 1217 498 1229 504
rect 1391 498 1403 504
rect 1497 498 1509 504
rect 1537 498 1549 504
rect 1656 498 1668 504
rect 1706 498 1718 504
rect 1811 498 1823 504
rect 1851 498 1863 504
rect 1937 498 1949 504
rect 2111 498 2123 504
rect 2221 498 2233 504
rect 2317 498 2329 504
rect 2361 498 2373 504
rect 2457 498 2469 504
rect 2497 498 2509 504
rect 2591 498 2603 504
rect 2631 498 2643 504
rect 2751 498 2763 504
rect 2995 544 3003 599
rect 3138 584 3146 619
rect 3077 578 3117 584
rect 3077 576 3089 578
rect 2822 498 2834 504
rect 2872 498 2884 504
rect 3235 552 3242 607
rect 3377 613 3385 662
rect 3495 655 3520 662
rect 3513 633 3521 655
rect 3235 546 3282 552
rect 3235 544 3243 546
rect 3271 544 3282 546
rect 3377 544 3385 599
rect 3519 584 3527 619
rect 3637 613 3645 662
rect 3755 655 3780 662
rect 3857 657 3873 663
rect 3707 637 3733 643
rect 3773 633 3781 655
rect 3857 627 3863 657
rect 3937 662 3945 676
rect 3920 655 3945 662
rect 2971 498 2983 504
rect 3011 498 3023 504
rect 3097 498 3109 504
rect 3251 498 3263 504
rect 3291 498 3303 504
rect 3357 498 3369 504
rect 3397 498 3409 504
rect 3637 544 3645 599
rect 3779 584 3787 619
rect 3919 633 3927 655
rect 4078 633 4086 676
rect 4189 676 4217 682
rect 4177 673 4229 676
rect 4438 716 4450 722
rect 4488 716 4500 722
rect 4611 716 4623 722
rect 4751 716 4763 722
rect 4877 716 4889 722
rect 4997 716 5009 722
rect 5139 716 5151 722
rect 5291 716 5303 722
rect 5397 716 5409 722
rect 5571 716 5583 722
rect 5657 716 5669 722
rect 5697 716 5709 722
rect 4237 662 4245 676
rect 4220 655 4245 662
rect 4219 633 4227 655
rect 4336 641 4344 696
rect 4434 676 4460 687
rect 4434 633 4442 676
rect 4575 662 4583 676
rect 4603 676 4631 682
rect 4591 673 4643 676
rect 4715 662 4723 676
rect 4743 676 4771 682
rect 4731 673 4783 676
rect 4869 676 4897 682
rect 4857 673 4909 676
rect 4917 662 4925 676
rect 4575 655 4600 662
rect 4715 655 4740 662
rect 4900 655 4925 662
rect 3913 584 3921 619
rect 4078 584 4086 619
rect 4213 584 4221 619
rect 3496 498 3508 504
rect 3546 498 3558 504
rect 3617 498 3629 504
rect 3657 498 3669 504
rect 3756 498 3768 504
rect 3806 498 3818 504
rect 4017 578 4057 584
rect 4017 576 4029 578
rect 4336 544 4344 627
rect 4593 633 4601 655
rect 4733 633 4741 655
rect 4899 633 4907 655
rect 5016 641 5024 696
rect 5121 670 5129 696
rect 5121 664 5143 670
rect 5140 658 5143 664
rect 4434 584 4442 619
rect 4599 584 4607 619
rect 4739 584 4747 619
rect 4893 584 4901 619
rect 4463 578 4503 584
rect 4491 576 4503 578
rect 3882 498 3894 504
rect 3932 498 3944 504
rect 4037 498 4049 504
rect 4182 498 4194 504
rect 4232 498 4244 504
rect 4351 498 4363 504
rect 4471 498 4483 504
rect 4576 498 4588 504
rect 4626 498 4638 504
rect 4716 498 4728 504
rect 4766 498 4778 504
rect 5016 544 5024 627
rect 5140 602 5147 658
rect 5161 633 5169 676
rect 5255 662 5263 676
rect 5283 676 5311 682
rect 5271 673 5323 676
rect 5389 676 5417 682
rect 5377 673 5429 676
rect 5437 662 5445 676
rect 5255 655 5280 662
rect 5420 655 5445 662
rect 5535 662 5543 676
rect 5563 676 5591 682
rect 5551 673 5603 676
rect 5535 655 5560 662
rect 5167 619 5169 633
rect 5273 633 5281 655
rect 5419 633 5427 655
rect 5553 633 5561 655
rect 5680 653 5687 696
rect 5140 596 5143 602
rect 5117 590 5143 596
rect 5117 544 5125 590
rect 5161 584 5169 619
rect 5279 584 5287 619
rect 5413 584 5421 619
rect 5559 584 5567 619
rect 5680 591 5687 639
rect 5680 584 5697 591
rect 4862 498 4874 504
rect 4912 498 4924 504
rect 4997 498 5009 504
rect 5139 498 5151 504
rect 5256 498 5268 504
rect 5306 498 5318 504
rect 5382 498 5394 504
rect 5432 498 5444 504
rect 5536 498 5548 504
rect 5586 498 5598 504
rect 5657 498 5669 504
rect -62 496 5816 498
rect -62 484 4 496
rect -62 482 5816 484
rect -62 18 -2 482
rect 91 476 103 482
rect 131 476 143 482
rect 75 434 83 436
rect 216 476 228 482
rect 266 476 278 482
rect 111 434 122 436
rect 75 428 122 434
rect 75 373 82 428
rect 376 476 388 482
rect 426 476 438 482
rect 531 476 543 482
rect 571 476 583 482
rect 667 476 679 482
rect 711 476 723 482
rect 811 476 823 482
rect 851 476 863 482
rect 971 476 983 482
rect 1057 476 1069 482
rect 1097 476 1109 482
rect 1241 476 1253 482
rect 1371 476 1383 482
rect 1411 476 1423 482
rect 1531 476 1543 482
rect 515 434 523 436
rect 551 434 562 436
rect 515 428 562 434
rect 239 361 247 396
rect 399 361 407 396
rect 515 373 522 428
rect 76 331 84 359
rect 76 322 106 331
rect 233 325 241 347
rect 393 325 401 347
rect 651 361 659 396
rect 516 331 524 359
rect 651 347 653 361
rect 76 320 94 322
rect 215 318 240 325
rect 375 318 400 325
rect 516 322 546 331
rect 516 320 534 322
rect 215 304 223 318
rect 231 304 283 307
rect 375 304 383 318
rect 243 298 271 304
rect 391 304 443 307
rect 403 298 431 304
rect 651 304 659 347
rect 694 322 702 436
rect 795 434 803 436
rect 831 434 842 436
rect 795 428 842 434
rect 795 373 802 428
rect 1078 434 1089 436
rect 1117 434 1125 436
rect 1078 428 1125 434
rect 991 402 1003 404
rect 963 396 1003 402
rect 934 361 942 396
rect 1118 373 1125 428
rect 1217 397 1221 406
rect 796 331 804 359
rect 796 322 826 331
rect 685 314 723 322
rect 796 320 814 322
rect 711 304 723 314
rect 651 294 661 304
rect 934 304 942 347
rect 1116 331 1124 359
rect 1217 353 1226 397
rect 1275 388 1283 396
rect 1247 380 1283 388
rect 1355 434 1363 436
rect 1616 476 1628 482
rect 1666 476 1678 482
rect 1767 476 1779 482
rect 1811 476 1823 482
rect 1391 434 1402 436
rect 1355 428 1402 434
rect 934 293 960 304
rect 130 258 142 264
rect 251 258 263 264
rect 411 258 423 264
rect 570 258 582 264
rect 681 258 693 264
rect 850 258 862 264
rect 938 258 950 264
rect 988 258 1000 264
rect 1094 322 1124 331
rect 1106 320 1124 322
rect 1213 304 1220 339
rect 1236 324 1242 379
rect 1355 373 1362 428
rect 1356 331 1364 359
rect 1516 353 1524 436
rect 1877 476 1889 482
rect 2017 476 2029 482
rect 2136 476 2148 482
rect 2186 476 2198 482
rect 2311 476 2323 482
rect 2431 476 2443 482
rect 2531 476 2543 482
rect 2571 476 2583 482
rect 1639 361 1647 396
rect 1751 361 1759 396
rect 1427 337 1473 343
rect 1356 322 1386 331
rect 1356 320 1374 322
rect 1247 312 1257 318
rect 1251 284 1257 312
rect 1516 284 1524 339
rect 1633 325 1641 347
rect 1751 347 1753 361
rect 1615 318 1640 325
rect 1615 304 1623 318
rect 1631 304 1683 307
rect 1643 298 1671 304
rect 1751 304 1759 347
rect 1794 322 1802 436
rect 1900 389 1917 396
rect 1900 341 1907 389
rect 2036 353 2044 436
rect 2331 402 2343 404
rect 2303 396 2343 402
rect 2159 361 2167 396
rect 2274 361 2282 396
rect 1785 314 1823 322
rect 1811 304 1823 314
rect 1751 294 1761 304
rect 1900 284 1907 327
rect 2036 284 2044 339
rect 2153 325 2161 347
rect 2416 353 2424 436
rect 2515 434 2523 436
rect 2642 476 2654 482
rect 2692 476 2704 482
rect 2811 476 2823 482
rect 2931 476 2943 482
rect 2551 434 2562 436
rect 2515 428 2562 434
rect 2515 373 2522 428
rect 2673 361 2681 396
rect 2135 318 2160 325
rect 2135 304 2143 318
rect 1058 258 1070 264
rect 1231 258 1243 264
rect 1275 258 1283 264
rect 1410 258 1422 264
rect 1531 258 1543 264
rect 1651 258 1663 264
rect 1781 258 1793 264
rect 1877 258 1889 264
rect 1917 258 1929 264
rect 2151 304 2203 307
rect 2163 298 2191 304
rect 2274 304 2282 347
rect 2274 293 2300 304
rect 2416 284 2424 339
rect 2516 331 2524 359
rect 2796 353 2804 436
rect 2997 476 3009 482
rect 3151 476 3163 482
rect 3277 476 3289 482
rect 3431 476 3443 482
rect 2903 389 2920 396
rect 2516 322 2546 331
rect 2679 325 2687 347
rect 2913 341 2920 389
rect 3016 353 3024 436
rect 3171 402 3183 404
rect 3143 396 3183 402
rect 3257 402 3269 404
rect 3257 396 3297 402
rect 3522 476 3534 482
rect 3572 476 3584 482
rect 3677 476 3689 482
rect 3831 476 3843 482
rect 3871 476 3883 482
rect 3114 361 3122 396
rect 3167 377 3293 383
rect 3318 361 3326 396
rect 2516 320 2534 322
rect 2680 318 2705 325
rect 2637 304 2689 307
rect 2649 298 2677 304
rect 2697 304 2705 318
rect 2796 284 2804 339
rect 2913 284 2920 327
rect 3016 284 3024 339
rect 3114 304 3122 347
rect 3416 353 3424 436
rect 3657 402 3669 404
rect 3657 396 3697 402
rect 3815 434 3823 436
rect 3937 476 3949 482
rect 3977 476 3989 482
rect 4111 476 4123 482
rect 4151 476 4163 482
rect 3851 434 3862 436
rect 3815 428 3862 434
rect 3553 361 3561 396
rect 3718 361 3726 396
rect 3815 373 3822 428
rect 3957 381 3965 436
rect 4095 434 4103 436
rect 4236 476 4248 482
rect 4286 476 4298 482
rect 4391 476 4403 482
rect 4131 434 4142 436
rect 4095 428 4142 434
rect 3318 304 3326 347
rect 3114 293 3140 304
rect 2017 258 2029 264
rect 2171 258 2183 264
rect 2278 258 2290 264
rect 2328 258 2340 264
rect 2431 258 2443 264
rect 2570 258 2582 264
rect 2657 258 2669 264
rect 2811 258 2823 264
rect 2891 258 2903 264
rect 2931 258 2943 264
rect 2997 258 3009 264
rect 3118 258 3130 264
rect 3168 258 3180 264
rect 3300 293 3326 304
rect 3416 284 3424 339
rect 3559 325 3567 347
rect 4095 373 4102 428
rect 4471 476 4483 482
rect 4511 476 4523 482
rect 4596 476 4608 482
rect 4646 476 4658 482
rect 4751 476 4763 482
rect 3560 318 3585 325
rect 3517 304 3569 307
rect 3529 298 3557 304
rect 3577 304 3585 318
rect 3718 304 3726 347
rect 3816 331 3824 359
rect 3816 322 3846 331
rect 3816 320 3834 322
rect 3700 293 3726 304
rect 3957 318 3965 367
rect 4259 361 4267 396
rect 4096 331 4104 359
rect 4096 322 4126 331
rect 4253 325 4261 347
rect 4376 353 4384 436
rect 4495 381 4503 436
rect 4836 476 4848 482
rect 4886 476 4898 482
rect 4096 320 4114 322
rect 3957 312 3981 318
rect 3969 304 3981 312
rect 3260 258 3272 264
rect 3310 258 3322 264
rect 3431 258 3443 264
rect 3537 258 3549 264
rect 3660 258 3672 264
rect 3710 258 3722 264
rect 3870 258 3882 264
rect 4235 318 4260 325
rect 4235 304 4243 318
rect 4251 304 4303 307
rect 4263 298 4291 304
rect 4376 284 4384 339
rect 4495 318 4503 367
rect 4619 361 4627 396
rect 4613 325 4621 347
rect 4736 353 4744 436
rect 4977 468 4989 482
rect 5037 476 5049 482
rect 4859 361 4867 396
rect 4963 394 4969 428
rect 5019 404 5021 406
rect 5007 400 5021 404
rect 4963 388 5004 394
rect 4479 312 4503 318
rect 4595 318 4620 325
rect 4479 304 4491 312
rect 4595 304 4603 318
rect 4611 304 4663 307
rect 4623 298 4651 304
rect 4736 284 4744 339
rect 4853 325 4861 347
rect 4995 370 5004 388
rect 4835 318 4860 325
rect 4995 320 5004 358
rect 5015 353 5021 400
rect 5136 476 5148 482
rect 5186 476 5198 482
rect 5282 476 5294 482
rect 5332 476 5344 482
rect 5491 476 5503 482
rect 5582 476 5594 482
rect 5632 476 5644 482
rect 5511 402 5523 404
rect 5483 396 5523 402
rect 5717 476 5729 482
rect 5757 476 5769 482
rect 5159 361 5167 396
rect 5313 361 5321 396
rect 5454 361 5462 396
rect 5613 361 5621 396
rect 5737 381 5745 436
rect 4835 304 4843 318
rect 4962 314 5004 320
rect 4851 304 4903 307
rect 4863 298 4891 304
rect 4962 292 4969 314
rect 5015 308 5021 339
rect 5153 325 5161 347
rect 5319 325 5327 347
rect 5135 318 5160 325
rect 5320 318 5345 325
rect 5007 304 5021 308
rect 5019 302 5021 304
rect 5135 304 5143 318
rect 3939 258 3951 264
rect 4150 258 4162 264
rect 4271 258 4283 264
rect 4391 258 4403 264
rect 4509 258 4521 264
rect 4631 258 4643 264
rect 4751 258 4763 264
rect 4871 258 4883 264
rect 4977 258 4989 272
rect 5037 258 5049 272
rect 5151 304 5203 307
rect 5163 298 5191 304
rect 5277 304 5329 307
rect 5289 298 5317 304
rect 5337 304 5345 318
rect 5454 304 5462 347
rect 5619 325 5627 347
rect 5620 318 5645 325
rect 5577 304 5629 307
rect 5454 293 5480 304
rect 5589 298 5617 304
rect 5637 304 5645 318
rect 5737 318 5745 367
rect 5737 312 5761 318
rect 5749 304 5761 312
rect 5171 258 5183 264
rect 5297 258 5309 264
rect 5458 258 5470 264
rect 5508 258 5520 264
rect 5597 258 5609 264
rect 5719 258 5731 264
rect 5822 258 5882 722
rect 4 256 5882 258
rect 5816 244 5882 256
rect 4 242 5882 244
rect 130 236 142 242
rect 76 178 94 180
rect 76 169 106 178
rect 200 236 212 242
rect 250 236 262 242
rect 378 236 390 242
rect 428 236 440 242
rect 551 236 563 242
rect 657 236 669 242
rect 850 236 862 242
rect 240 196 266 207
rect 76 141 84 169
rect 258 153 266 196
rect 374 196 400 207
rect 374 153 382 196
rect 515 182 523 196
rect 543 196 571 202
rect 531 193 583 196
rect 649 196 677 202
rect 637 193 689 196
rect 697 182 705 196
rect 515 175 540 182
rect 680 175 705 182
rect 796 178 814 180
rect 533 153 541 175
rect 679 153 687 175
rect 796 169 826 178
rect 917 236 929 242
rect 1037 236 1049 242
rect 1160 236 1172 242
rect 1210 236 1222 242
rect 796 141 804 169
rect 936 161 944 216
rect 1029 196 1057 202
rect 1017 193 1069 196
rect 1297 236 1309 242
rect 1337 236 1349 242
rect 1447 236 1459 242
rect 1591 236 1603 242
rect 1711 236 1723 242
rect 1849 236 1861 242
rect 1200 196 1226 207
rect 1077 182 1085 196
rect 1060 175 1085 182
rect 75 72 82 127
rect 258 104 266 139
rect 374 104 382 139
rect 539 104 547 139
rect 673 104 681 139
rect 197 98 237 104
rect 197 96 209 98
rect 75 66 122 72
rect 75 64 83 66
rect 111 64 122 66
rect 403 98 443 104
rect 431 96 443 98
rect 91 18 103 24
rect 131 18 143 24
rect 217 18 229 24
rect 411 18 423 24
rect 516 18 528 24
rect 566 18 578 24
rect 795 72 802 127
rect 795 66 842 72
rect 795 64 803 66
rect 831 64 842 66
rect 936 64 944 147
rect 1059 153 1067 175
rect 1218 153 1226 196
rect 1320 173 1327 216
rect 1479 196 1489 206
rect 1417 186 1429 196
rect 1417 178 1455 186
rect 1053 104 1061 139
rect 1218 104 1226 139
rect 1320 111 1327 159
rect 1320 104 1337 111
rect 642 18 654 24
rect 692 18 704 24
rect 811 18 823 24
rect 851 18 863 24
rect 1157 98 1197 104
rect 1157 96 1169 98
rect 1438 64 1446 178
rect 1481 153 1489 196
rect 1576 161 1584 216
rect 1675 182 1683 196
rect 1703 196 1731 202
rect 1691 193 1743 196
rect 1918 236 1930 242
rect 2150 236 2162 242
rect 2239 236 2251 242
rect 2389 236 2401 242
rect 2487 236 2499 242
rect 2618 236 2630 242
rect 2668 236 2680 242
rect 2781 236 2793 242
rect 2899 236 2911 242
rect 3069 236 3081 242
rect 3210 236 3222 242
rect 3311 236 3323 242
rect 3397 236 3409 242
rect 3551 236 3563 242
rect 3669 236 3681 242
rect 3769 236 3781 242
rect 3879 236 3891 242
rect 4029 236 4041 242
rect 4147 236 4159 242
rect 4291 236 4303 242
rect 4331 236 4343 242
rect 1819 188 1831 196
rect 1819 182 1843 188
rect 1675 175 1700 182
rect 1487 139 1489 153
rect 1693 153 1701 175
rect 1481 104 1489 139
rect 1576 64 1584 147
rect 1699 104 1707 139
rect 1835 133 1843 182
rect 1966 178 1984 180
rect 1954 169 1984 178
rect 1976 141 1984 169
rect 2096 178 2114 180
rect 2096 169 2126 178
rect 2221 190 2229 216
rect 2519 196 2529 206
rect 2221 184 2243 190
rect 2240 178 2243 184
rect 2096 141 2104 169
rect 917 18 929 24
rect 1022 18 1034 24
rect 1072 18 1084 24
rect 1177 18 1189 24
rect 1297 18 1309 24
rect 1417 18 1429 24
rect 1461 18 1473 24
rect 1591 18 1603 24
rect 1835 64 1843 119
rect 1978 72 1985 127
rect 1938 66 1985 72
rect 1938 64 1949 66
rect 1676 18 1688 24
rect 1726 18 1738 24
rect 1811 18 1823 24
rect 1851 18 1863 24
rect 1977 64 1985 66
rect 2095 72 2102 127
rect 2240 122 2247 178
rect 2261 153 2269 196
rect 2359 188 2371 196
rect 2359 182 2383 188
rect 2267 139 2269 153
rect 2240 116 2243 122
rect 2217 110 2243 116
rect 2095 66 2142 72
rect 2095 64 2103 66
rect 2131 64 2142 66
rect 2217 64 2225 110
rect 2261 104 2269 139
rect 2375 133 2383 182
rect 2457 186 2469 196
rect 2457 178 2495 186
rect 2375 64 2383 119
rect 2478 64 2486 178
rect 2521 153 2529 196
rect 2614 196 2640 207
rect 2751 196 2761 206
rect 2614 153 2622 196
rect 2527 139 2529 153
rect 2751 153 2759 196
rect 2811 186 2823 196
rect 2929 188 2941 196
rect 2785 178 2823 186
rect 2917 182 2941 188
rect 3039 188 3051 196
rect 3039 182 3063 188
rect 2751 139 2753 153
rect 2521 104 2529 139
rect 2614 104 2622 139
rect 2751 104 2759 139
rect 1917 18 1929 24
rect 1957 18 1969 24
rect 2111 18 2123 24
rect 2151 18 2163 24
rect 2239 18 2251 24
rect 2351 18 2363 24
rect 2391 18 2403 24
rect 2643 98 2683 104
rect 2671 96 2683 98
rect 2794 64 2802 178
rect 2917 133 2925 182
rect 3055 133 3063 182
rect 3156 178 3174 180
rect 3156 169 3186 178
rect 3156 141 3164 169
rect 3296 161 3304 216
rect 3389 196 3417 202
rect 3377 193 3429 196
rect 3437 182 3445 196
rect 3420 175 3445 182
rect 2917 64 2925 119
rect 2987 97 3033 103
rect 3055 64 3063 119
rect 3155 72 3162 127
rect 3155 66 3202 72
rect 3155 64 3163 66
rect 2457 18 2469 24
rect 2501 18 2513 24
rect 2651 18 2663 24
rect 2767 18 2779 24
rect 2811 18 2823 24
rect 2897 18 2909 24
rect 2937 18 2949 24
rect 3191 64 3202 66
rect 3296 64 3304 147
rect 3419 153 3427 175
rect 3536 161 3544 216
rect 3639 188 3651 196
rect 3639 182 3663 188
rect 3413 104 3421 139
rect 3031 18 3043 24
rect 3071 18 3083 24
rect 3171 18 3183 24
rect 3211 18 3223 24
rect 3311 18 3323 24
rect 3536 64 3544 147
rect 3655 133 3663 182
rect 3751 153 3759 196
rect 3791 190 3799 216
rect 3777 184 3799 190
rect 3861 190 3869 216
rect 4399 236 4411 242
rect 4590 236 4602 242
rect 4731 236 4743 242
rect 4819 236 4831 242
rect 4991 236 5003 242
rect 5077 236 5089 242
rect 5117 236 5129 242
rect 5249 236 5261 242
rect 4179 196 4189 206
rect 3861 184 3883 190
rect 3777 178 3780 184
rect 3751 139 3753 153
rect 3655 64 3663 119
rect 3751 104 3759 139
rect 3773 122 3780 178
rect 3880 178 3883 184
rect 3777 116 3780 122
rect 3880 122 3887 178
rect 3901 153 3909 196
rect 3999 188 4011 196
rect 3999 182 4023 188
rect 3907 139 3909 153
rect 3880 116 3883 122
rect 3777 110 3803 116
rect 3382 18 3394 24
rect 3432 18 3444 24
rect 3551 18 3563 24
rect 3795 64 3803 110
rect 3857 110 3883 116
rect 3857 64 3865 110
rect 3901 104 3909 139
rect 4015 133 4023 182
rect 4117 186 4129 196
rect 4117 178 4155 186
rect 4015 64 4023 119
rect 4138 64 4146 178
rect 4181 153 4189 196
rect 4313 173 4320 216
rect 4429 188 4441 196
rect 4417 182 4441 188
rect 4187 139 4189 153
rect 4181 104 4189 139
rect 4313 111 4320 159
rect 4417 133 4425 182
rect 4536 178 4554 180
rect 4536 169 4566 178
rect 4695 182 4703 196
rect 4723 196 4751 202
rect 4711 193 4763 196
rect 4849 188 4861 196
rect 4837 182 4861 188
rect 4955 182 4963 196
rect 4983 196 5011 202
rect 4971 193 5023 196
rect 4695 175 4720 182
rect 4536 141 4544 169
rect 4587 157 4613 163
rect 4713 153 4721 175
rect 4303 104 4320 111
rect 3631 18 3643 24
rect 3671 18 3683 24
rect 3769 18 3781 24
rect 3879 18 3891 24
rect 3991 18 4003 24
rect 4031 18 4043 24
rect 4417 64 4425 119
rect 4535 72 4542 127
rect 4719 104 4727 139
rect 4837 133 4845 182
rect 4955 175 4980 182
rect 4973 153 4981 175
rect 5100 173 5107 216
rect 5337 228 5349 242
rect 5397 228 5409 242
rect 5219 188 5231 196
rect 5219 182 5243 188
rect 4535 66 4582 72
rect 4535 64 4543 66
rect 4117 18 4129 24
rect 4161 18 4173 24
rect 4331 18 4343 24
rect 4571 64 4582 66
rect 4397 18 4409 24
rect 4437 18 4449 24
rect 4551 18 4563 24
rect 4591 18 4603 24
rect 4837 64 4845 119
rect 4979 104 4987 139
rect 5100 111 5107 159
rect 5235 133 5243 182
rect 5322 186 5329 208
rect 5379 196 5381 198
rect 5367 192 5381 196
rect 5322 180 5364 186
rect 5355 142 5364 180
rect 5375 161 5381 192
rect 5477 236 5489 242
rect 5611 236 5623 242
rect 5679 236 5691 242
rect 5496 161 5504 216
rect 5596 161 5604 216
rect 5709 188 5721 196
rect 5697 182 5721 188
rect 5100 104 5117 111
rect 4696 18 4708 24
rect 4746 18 4758 24
rect 4817 18 4829 24
rect 4857 18 4869 24
rect 4956 18 4968 24
rect 5006 18 5018 24
rect 5235 64 5243 119
rect 5355 112 5364 130
rect 5323 106 5364 112
rect 5323 72 5329 106
rect 5375 100 5381 147
rect 5367 96 5381 100
rect 5379 94 5381 96
rect 5077 18 5089 24
rect 5211 18 5223 24
rect 5251 18 5263 24
rect 5337 18 5349 32
rect 5496 64 5504 147
rect 5596 64 5604 147
rect 5697 133 5705 182
rect 5697 64 5705 119
rect 5397 18 5409 24
rect 5477 18 5489 24
rect 5611 18 5623 24
rect 5677 18 5689 24
rect 5717 18 5729 24
rect -62 16 5816 18
rect -62 4 4 16
rect -62 2 5816 4
rect 5822 2 5882 242
<< m2contact >>
rect 73 5647 87 5661
rect 253 5647 267 5661
rect 513 5667 527 5681
rect 493 5647 507 5661
rect 533 5647 547 5661
rect 93 5627 107 5641
rect 113 5619 127 5633
rect 133 5627 147 5641
rect 193 5627 207 5641
rect 213 5619 227 5633
rect 233 5627 247 5641
rect 373 5627 387 5641
rect 553 5639 567 5653
rect 653 5647 667 5661
rect 393 5619 407 5633
rect 413 5607 427 5621
rect 433 5619 447 5633
rect 673 5627 687 5641
rect 693 5619 707 5633
rect 713 5627 727 5641
rect 793 5639 807 5653
rect 813 5647 827 5661
rect 833 5639 847 5653
rect 913 5627 927 5641
rect 933 5619 947 5633
rect 953 5607 967 5621
rect 973 5619 987 5633
rect 1053 5627 1067 5641
rect 1093 5627 1107 5641
rect 1073 5607 1087 5621
rect 1213 5619 1227 5633
rect 1253 5627 1267 5641
rect 1353 5627 1367 5641
rect 1373 5639 1387 5653
rect 1273 5607 1287 5621
rect 1533 5667 1547 5681
rect 1413 5627 1427 5641
rect 1493 5639 1507 5653
rect 1513 5647 1527 5661
rect 1553 5647 1567 5661
rect 1833 5667 1847 5681
rect 1653 5627 1667 5641
rect 1793 5639 1807 5653
rect 1813 5647 1827 5661
rect 1853 5647 1867 5661
rect 1673 5619 1687 5633
rect 1693 5607 1707 5621
rect 1713 5619 1727 5633
rect 2033 5647 2047 5661
rect 2213 5647 2227 5661
rect 1913 5607 1927 5621
rect 1933 5619 1947 5633
rect 2053 5627 2067 5641
rect 2073 5619 2087 5633
rect 2093 5627 2107 5641
rect 2153 5627 2167 5641
rect 2173 5619 2187 5633
rect 2193 5627 2207 5641
rect 2293 5619 2307 5633
rect 2313 5607 2327 5621
rect 2333 5619 2347 5633
rect 2353 5627 2367 5641
rect 2453 5639 2467 5653
rect 2473 5647 2487 5661
rect 2613 5667 2627 5681
rect 2493 5639 2507 5653
rect 2573 5639 2587 5653
rect 2593 5647 2607 5661
rect 2633 5647 2647 5661
rect 2753 5667 2767 5681
rect 2713 5639 2727 5653
rect 2733 5647 2747 5661
rect 2773 5647 2787 5661
rect 2833 5639 2847 5653
rect 2853 5647 2867 5661
rect 2873 5639 2887 5653
rect 3073 5647 3087 5661
rect 2973 5619 2987 5633
rect 3093 5627 3107 5641
rect 2993 5607 3007 5621
rect 3113 5619 3127 5633
rect 3133 5627 3147 5641
rect 3233 5627 3247 5641
rect 3253 5639 3267 5653
rect 3293 5627 3307 5641
rect 3373 5627 3387 5641
rect 3533 5667 3547 5681
rect 3413 5627 3427 5641
rect 3493 5639 3507 5653
rect 3513 5647 3527 5661
rect 3553 5647 3567 5661
rect 3393 5607 3407 5621
rect 3993 5647 4007 5661
rect 3653 5619 3667 5633
rect 3673 5607 3687 5621
rect 3753 5619 3767 5633
rect 3773 5607 3787 5621
rect 3833 5607 3847 5621
rect 3853 5619 3867 5633
rect 3933 5627 3947 5641
rect 3953 5619 3967 5633
rect 3973 5627 3987 5641
rect 4173 5702 4187 5716
rect 4313 5696 4327 5710
rect 4073 5607 4087 5621
rect 4093 5619 4107 5633
rect 4173 5664 4187 5678
rect 4153 5599 4167 5613
rect 4233 5627 4247 5641
rect 4273 5627 4287 5641
rect 4173 5570 4187 5584
rect 4453 5647 4467 5661
rect 4473 5627 4487 5641
rect 4493 5619 4507 5633
rect 4513 5627 4527 5641
rect 4593 5619 4607 5633
rect 4933 5647 4947 5661
rect 4733 5619 4747 5633
rect 4833 5619 4847 5633
rect 4953 5627 4967 5641
rect 4313 5570 4327 5584
rect 4853 5607 4867 5621
rect 4973 5619 4987 5633
rect 4993 5627 5007 5641
rect 5073 5639 5087 5653
rect 5093 5647 5107 5661
rect 5113 5639 5127 5653
rect 5173 5639 5187 5653
rect 5193 5647 5207 5661
rect 5213 5639 5227 5653
rect 5353 5647 5367 5661
rect 5293 5627 5307 5641
rect 5313 5619 5327 5633
rect 5333 5627 5347 5641
rect 5533 5639 5547 5653
rect 5553 5647 5567 5661
rect 5433 5607 5447 5621
rect 5453 5619 5467 5633
rect 5573 5639 5587 5653
rect 5653 5607 5667 5621
rect 5673 5619 5687 5633
rect 93 5419 107 5433
rect 113 5427 127 5441
rect 133 5419 147 5433
rect 73 5399 87 5413
rect 233 5407 247 5421
rect 253 5399 267 5413
rect 293 5399 307 5413
rect 373 5407 387 5421
rect 273 5379 287 5393
rect 393 5399 407 5413
rect 433 5399 447 5413
rect 513 5407 527 5421
rect 413 5379 427 5393
rect 533 5399 547 5413
rect 573 5399 587 5413
rect 653 5399 667 5413
rect 693 5399 707 5413
rect 713 5407 727 5421
rect 793 5419 807 5433
rect 813 5427 827 5441
rect 833 5419 847 5433
rect 553 5379 567 5393
rect 673 5379 687 5393
rect 853 5399 867 5413
rect 933 5399 947 5413
rect 973 5399 987 5413
rect 993 5407 1007 5421
rect 1093 5419 1107 5433
rect 1113 5427 1127 5441
rect 1133 5439 1147 5453
rect 1153 5427 1167 5441
rect 1393 5439 1407 5453
rect 953 5379 967 5393
rect 1113 5393 1127 5407
rect 1193 5393 1207 5407
rect 1213 5399 1227 5413
rect 1253 5399 1267 5413
rect 1273 5407 1287 5421
rect 1373 5419 1387 5433
rect 1233 5379 1247 5393
rect 1413 5419 1427 5433
rect 1513 5407 1527 5421
rect 1633 5419 1647 5433
rect 1653 5427 1667 5441
rect 1673 5419 1687 5433
rect 1533 5399 1547 5413
rect 1573 5399 1587 5413
rect 1553 5379 1567 5393
rect 1693 5399 1707 5413
rect 1793 5407 1807 5421
rect 1813 5399 1827 5413
rect 1853 5399 1867 5413
rect 1933 5407 1947 5421
rect 1833 5379 1847 5393
rect 1953 5399 1967 5413
rect 1993 5399 2007 5413
rect 2053 5407 2067 5421
rect 2213 5427 2227 5441
rect 2233 5439 2247 5453
rect 2073 5399 2087 5413
rect 2093 5407 2107 5421
rect 1973 5379 1987 5393
rect 2313 5419 2327 5433
rect 2333 5407 2347 5421
rect 2373 5419 2387 5433
rect 2433 5419 2447 5433
rect 2453 5427 2467 5441
rect 2473 5419 2487 5433
rect 2493 5399 2507 5413
rect 2613 5407 2627 5421
rect 2633 5399 2647 5413
rect 2673 5399 2687 5413
rect 2753 5407 2767 5421
rect 2873 5419 2887 5433
rect 2893 5427 2907 5441
rect 3013 5439 3027 5453
rect 2913 5419 2927 5433
rect 3033 5427 3047 5441
rect 2653 5379 2667 5393
rect 2773 5399 2787 5413
rect 2813 5399 2827 5413
rect 2793 5379 2807 5393
rect 2933 5399 2947 5413
rect 3113 5407 3127 5421
rect 3133 5399 3147 5413
rect 3153 5407 3167 5421
rect 3253 5399 3267 5413
rect 3293 5399 3307 5413
rect 3313 5407 3327 5421
rect 3393 5407 3407 5421
rect 3513 5439 3527 5453
rect 3273 5379 3287 5393
rect 3413 5399 3427 5413
rect 3433 5407 3447 5421
rect 3533 5419 3547 5433
rect 3573 5427 3587 5441
rect 3673 5407 3687 5421
rect 3813 5419 3827 5433
rect 3833 5427 3847 5441
rect 3853 5439 3867 5453
rect 3873 5427 3887 5441
rect 3693 5399 3707 5413
rect 3733 5399 3747 5413
rect 3713 5379 3727 5393
rect 3933 5407 3947 5421
rect 3953 5399 3967 5413
rect 3973 5407 3987 5421
rect 4093 5419 4107 5433
rect 4113 5427 4127 5441
rect 4133 5419 4147 5433
rect 4073 5399 4087 5413
rect 4213 5407 4227 5421
rect 4473 5427 4487 5441
rect 4493 5439 4507 5453
rect 4513 5427 4527 5441
rect 4613 5439 4627 5453
rect 4853 5476 4867 5490
rect 4993 5476 5007 5490
rect 4233 5399 4247 5413
rect 4253 5407 4267 5421
rect 4333 5407 4347 5421
rect 4533 5419 4547 5433
rect 4633 5427 4647 5441
rect 4353 5399 4367 5413
rect 4393 5399 4407 5413
rect 4373 5379 4387 5393
rect 4713 5419 4727 5433
rect 4733 5427 4747 5441
rect 4753 5419 4767 5433
rect 4833 5447 4847 5461
rect 4773 5399 4787 5413
rect 4853 5382 4867 5396
rect 4913 5419 4927 5433
rect 4953 5419 4967 5433
rect 5093 5439 5107 5453
rect 5193 5476 5207 5490
rect 5333 5476 5347 5490
rect 5173 5447 5187 5461
rect 5113 5427 5127 5441
rect 4853 5344 4867 5358
rect 4993 5350 5007 5364
rect 5193 5382 5207 5396
rect 5253 5419 5267 5433
rect 5293 5419 5307 5433
rect 5433 5419 5447 5433
rect 5453 5427 5467 5441
rect 5473 5419 5487 5433
rect 5493 5399 5507 5413
rect 5593 5407 5607 5421
rect 5613 5399 5627 5413
rect 5633 5407 5647 5421
rect 5193 5344 5207 5358
rect 5333 5350 5347 5364
rect 5713 5453 5727 5467
rect 5713 5407 5727 5421
rect 5733 5399 5747 5413
rect 5753 5407 5767 5421
rect 5713 5373 5727 5387
rect 113 5187 127 5201
rect 73 5159 87 5173
rect 93 5167 107 5181
rect 133 5167 147 5181
rect 193 5139 207 5153
rect 213 5127 227 5141
rect 233 5139 247 5153
rect 253 5147 267 5161
rect 493 5187 507 5201
rect 453 5159 467 5173
rect 473 5167 487 5181
rect 513 5167 527 5181
rect 873 5187 887 5201
rect 853 5167 867 5181
rect 893 5167 907 5181
rect 1053 5187 1067 5201
rect 333 5127 347 5141
rect 353 5139 367 5153
rect 573 5139 587 5153
rect 593 5127 607 5141
rect 613 5139 627 5153
rect 633 5147 647 5161
rect 733 5147 747 5161
rect 913 5159 927 5173
rect 1013 5159 1027 5173
rect 1033 5167 1047 5181
rect 1073 5167 1087 5181
rect 753 5139 767 5153
rect 773 5127 787 5141
rect 793 5139 807 5153
rect 1293 5187 1307 5201
rect 1253 5159 1267 5173
rect 1273 5167 1287 5181
rect 1313 5167 1327 5181
rect 1413 5167 1427 5181
rect 1133 5127 1147 5141
rect 1153 5139 1167 5153
rect 1433 5147 1447 5161
rect 1453 5139 1467 5153
rect 1473 5147 1487 5161
rect 1653 5167 1667 5181
rect 1553 5139 1567 5153
rect 1673 5147 1687 5161
rect 1573 5127 1587 5141
rect 1693 5139 1707 5153
rect 1713 5147 1727 5161
rect 1833 5139 1847 5153
rect 1873 5147 1887 5161
rect 1893 5139 1907 5153
rect 1933 5147 1947 5161
rect 2033 5147 2047 5161
rect 2053 5139 2067 5153
rect 2073 5147 2087 5161
rect 1573 5093 1587 5107
rect 1613 5093 1627 5107
rect 2093 5139 2107 5153
rect 2113 5147 2127 5161
rect 2173 5159 2187 5173
rect 2193 5167 2207 5181
rect 2353 5187 2367 5201
rect 2213 5159 2227 5173
rect 2313 5159 2327 5173
rect 2333 5167 2347 5181
rect 2373 5167 2387 5181
rect 2453 5147 2467 5161
rect 2693 5167 2707 5181
rect 2853 5167 2867 5181
rect 2473 5139 2487 5153
rect 2493 5127 2507 5141
rect 2513 5139 2527 5153
rect 2593 5139 2607 5153
rect 2713 5147 2727 5161
rect 2613 5127 2627 5141
rect 2733 5139 2747 5153
rect 2753 5147 2767 5161
rect 2873 5147 2887 5161
rect 2893 5139 2907 5153
rect 2913 5147 2927 5161
rect 2993 5147 3007 5161
rect 3013 5159 3027 5173
rect 3053 5147 3067 5161
rect 3113 5147 3127 5161
rect 3153 5147 3167 5161
rect 3133 5127 3147 5141
rect 3273 5139 3287 5153
rect 3373 5147 3387 5161
rect 3513 5167 3527 5181
rect 3953 5193 3967 5207
rect 3413 5147 3427 5161
rect 3533 5147 3547 5161
rect 3293 5127 3307 5141
rect 3393 5127 3407 5141
rect 3553 5139 3567 5153
rect 3573 5147 3587 5161
rect 3633 5159 3647 5173
rect 3653 5167 3667 5181
rect 3673 5159 3687 5173
rect 3773 5159 3787 5173
rect 3793 5167 3807 5181
rect 3813 5159 3827 5173
rect 3913 5159 3927 5173
rect 3933 5167 3947 5181
rect 3953 5159 3967 5173
rect 4033 5187 4047 5201
rect 4013 5167 4027 5181
rect 4053 5167 4067 5181
rect 4073 5159 4087 5173
rect 4173 5167 4187 5181
rect 4373 5167 4387 5181
rect 4013 5133 4027 5147
rect 4193 5147 4207 5161
rect 4213 5139 4227 5153
rect 4233 5147 4247 5161
rect 4313 5147 4327 5161
rect 4333 5139 4347 5153
rect 4353 5147 4367 5161
rect 4613 5187 4627 5201
rect 4573 5159 4587 5173
rect 4593 5167 4607 5181
rect 4633 5167 4647 5181
rect 4953 5222 4967 5236
rect 5093 5216 5107 5230
rect 4453 5127 4467 5141
rect 4473 5139 4487 5153
rect 4693 5139 4707 5153
rect 4713 5127 4727 5141
rect 4733 5139 4747 5153
rect 4753 5147 4767 5161
rect 4833 5147 4847 5161
rect 4873 5147 4887 5161
rect 4853 5127 4867 5141
rect 4953 5184 4967 5198
rect 4933 5119 4947 5133
rect 5013 5147 5027 5161
rect 5053 5147 5067 5161
rect 4953 5090 4967 5104
rect 5253 5167 5267 5181
rect 5193 5147 5207 5161
rect 5213 5139 5227 5153
rect 5233 5147 5247 5161
rect 5753 5193 5767 5207
rect 5493 5167 5507 5181
rect 5333 5127 5347 5141
rect 5353 5139 5367 5153
rect 5433 5147 5447 5161
rect 5453 5139 5467 5153
rect 5473 5147 5487 5161
rect 5593 5159 5607 5173
rect 5613 5167 5627 5181
rect 5093 5090 5107 5104
rect 5633 5159 5647 5173
rect 5693 5159 5707 5173
rect 5713 5167 5727 5181
rect 5733 5159 5747 5173
rect 5753 5113 5767 5127
rect 93 4939 107 4953
rect 113 4947 127 4961
rect 133 4939 147 4953
rect 73 4919 87 4933
rect 213 4927 227 4941
rect 233 4919 247 4933
rect 273 4919 287 4933
rect 333 4919 347 4933
rect 373 4919 387 4933
rect 393 4927 407 4941
rect 473 4939 487 4953
rect 493 4947 507 4961
rect 513 4939 527 4953
rect 253 4899 267 4913
rect 353 4899 367 4913
rect 533 4919 547 4933
rect 633 4927 647 4941
rect 653 4919 667 4933
rect 673 4927 687 4941
rect 773 4939 787 4953
rect 793 4947 807 4961
rect 813 4939 827 4953
rect 913 4939 927 4953
rect 933 4947 947 4961
rect 953 4939 967 4953
rect 1033 4939 1047 4953
rect 1053 4947 1067 4961
rect 1073 4959 1087 4973
rect 1093 4947 1107 4961
rect 1193 4939 1207 4953
rect 1213 4947 1227 4961
rect 1233 4939 1247 4953
rect 1313 4947 1327 4961
rect 1333 4959 1347 4973
rect 753 4919 767 4933
rect 893 4919 907 4933
rect 1173 4919 1187 4933
rect 1413 4927 1427 4941
rect 1433 4919 1447 4933
rect 1453 4927 1467 4941
rect 1553 4927 1567 4941
rect 1713 4939 1727 4953
rect 1733 4947 1747 4961
rect 1753 4939 1767 4953
rect 1813 4947 1827 4961
rect 1833 4959 1847 4973
rect 1853 4947 1867 4961
rect 1873 4939 1887 4953
rect 1573 4919 1587 4933
rect 1613 4919 1627 4933
rect 1693 4919 1707 4933
rect 1593 4899 1607 4913
rect 1953 4927 1967 4941
rect 1973 4919 1987 4933
rect 1993 4927 2007 4941
rect 2093 4939 2107 4953
rect 2113 4947 2127 4961
rect 2133 4959 2147 4973
rect 2153 4947 2167 4961
rect 2253 4947 2267 4961
rect 2273 4959 2287 4973
rect 2373 4939 2387 4953
rect 2393 4947 2407 4961
rect 2413 4939 2427 4953
rect 2633 4947 2647 4961
rect 2653 4959 2667 4973
rect 2353 4919 2367 4933
rect 2493 4927 2507 4941
rect 2513 4919 2527 4933
rect 2553 4919 2567 4933
rect 2533 4899 2547 4913
rect 2753 4927 2767 4941
rect 2853 4959 2867 4973
rect 2873 4947 2887 4961
rect 2773 4919 2787 4933
rect 2793 4927 2807 4941
rect 2793 4893 2807 4907
rect 2833 4893 2847 4907
rect 2953 4919 2967 4933
rect 2993 4919 3007 4933
rect 3013 4927 3027 4941
rect 3133 4939 3147 4953
rect 3153 4947 3167 4961
rect 3173 4939 3187 4953
rect 3273 4939 3287 4953
rect 3293 4947 3307 4961
rect 3313 4939 3327 4953
rect 3393 4939 3407 4953
rect 3413 4947 3427 4961
rect 3433 4959 3447 4973
rect 3453 4947 3467 4961
rect 3513 4959 3527 4973
rect 3533 4939 3547 4953
rect 2973 4899 2987 4913
rect 3113 4919 3127 4933
rect 3253 4919 3267 4933
rect 3573 4947 3587 4961
rect 3693 4959 3707 4973
rect 3673 4939 3687 4953
rect 3713 4939 3727 4953
rect 3933 4947 3947 4961
rect 3953 4959 3967 4973
rect 3793 4927 3807 4941
rect 3813 4919 3827 4933
rect 3853 4919 3867 4933
rect 3833 4899 3847 4913
rect 4113 4953 4127 4967
rect 4173 4953 4187 4967
rect 4013 4919 4027 4933
rect 4053 4919 4067 4933
rect 4073 4927 4087 4941
rect 4033 4899 4047 4913
rect 4153 4919 4167 4933
rect 4193 4919 4207 4933
rect 4213 4927 4227 4941
rect 4313 4939 4327 4953
rect 4173 4899 4187 4913
rect 4333 4927 4347 4941
rect 4453 4959 4467 4973
rect 4373 4939 4387 4953
rect 4473 4939 4487 4953
rect 4853 4996 4867 5010
rect 4993 4996 5007 5010
rect 4513 4947 4527 4961
rect 4613 4959 4627 4973
rect 4593 4939 4607 4953
rect 4833 4967 4847 4981
rect 4633 4939 4647 4953
rect 4753 4939 4767 4953
rect 4773 4947 4787 4961
rect 4793 4939 4807 4953
rect 4733 4919 4747 4933
rect 4853 4902 4867 4916
rect 4913 4939 4927 4953
rect 4953 4939 4967 4953
rect 5233 4996 5247 5010
rect 5373 4996 5387 5010
rect 5093 4939 5107 4953
rect 5113 4947 5127 4961
rect 5133 4939 5147 4953
rect 5213 4967 5227 4981
rect 5153 4919 5167 4933
rect 4853 4864 4867 4878
rect 4993 4870 5007 4884
rect 5233 4902 5247 4916
rect 5293 4939 5307 4953
rect 5333 4939 5347 4953
rect 5493 4927 5507 4941
rect 5553 4973 5567 4987
rect 5513 4919 5527 4933
rect 5533 4927 5547 4941
rect 5233 4864 5247 4878
rect 5373 4870 5387 4884
rect 5533 4893 5547 4907
rect 5593 4973 5607 4987
rect 5593 4927 5607 4941
rect 5613 4919 5627 4933
rect 5633 4927 5647 4941
rect 5733 4927 5747 4941
rect 5753 4919 5767 4933
rect 5773 4927 5787 4941
rect 5593 4873 5607 4887
rect 253 4707 267 4721
rect 73 4667 87 4681
rect 213 4679 227 4693
rect 233 4687 247 4701
rect 273 4687 287 4701
rect 93 4659 107 4673
rect 113 4647 127 4661
rect 133 4659 147 4673
rect 333 4659 347 4673
rect 353 4647 367 4661
rect 373 4659 387 4673
rect 393 4667 407 4681
rect 473 4679 487 4693
rect 493 4687 507 4701
rect 653 4707 667 4721
rect 513 4679 527 4693
rect 613 4679 627 4693
rect 633 4687 647 4701
rect 673 4687 687 4701
rect 813 4707 827 4721
rect 773 4679 787 4693
rect 793 4687 807 4701
rect 833 4687 847 4701
rect 1213 4687 1227 4701
rect 1393 4687 1407 4701
rect 893 4647 907 4661
rect 913 4659 927 4673
rect 993 4647 1007 4661
rect 1013 4659 1027 4673
rect 1113 4659 1127 4673
rect 1233 4667 1247 4681
rect 1133 4647 1147 4661
rect 1253 4659 1267 4673
rect 1273 4667 1287 4681
rect 1333 4667 1347 4681
rect 1353 4659 1367 4673
rect 1373 4667 1387 4681
rect 1593 4707 1607 4721
rect 1573 4687 1587 4701
rect 1613 4687 1627 4701
rect 1633 4679 1647 4693
rect 1733 4687 1747 4701
rect 1473 4647 1487 4661
rect 1493 4659 1507 4673
rect 1753 4667 1767 4681
rect 1773 4659 1787 4673
rect 1793 4667 1807 4681
rect 1873 4679 1887 4693
rect 1893 4687 1907 4701
rect 1913 4679 1927 4693
rect 2033 4687 2047 4701
rect 2173 4707 2187 4721
rect 1973 4667 1987 4681
rect 1993 4659 2007 4673
rect 2013 4667 2027 4681
rect 2133 4679 2147 4693
rect 2153 4687 2167 4701
rect 2193 4687 2207 4701
rect 2273 4667 2287 4681
rect 2313 4667 2327 4681
rect 2373 4679 2387 4693
rect 2393 4687 2407 4701
rect 2413 4679 2427 4693
rect 2493 4679 2507 4693
rect 2513 4687 2527 4701
rect 2533 4679 2547 4693
rect 2753 4707 2767 4721
rect 2633 4667 2647 4681
rect 2733 4687 2747 4701
rect 2773 4687 2787 4701
rect 2673 4667 2687 4681
rect 2793 4679 2807 4693
rect 2893 4667 2907 4681
rect 2933 4667 2947 4681
rect 3013 4667 3027 4681
rect 2913 4647 2927 4661
rect 3033 4659 3047 4673
rect 3053 4667 3067 4681
rect 3073 4659 3087 4673
rect 3093 4667 3107 4681
rect 3193 4679 3207 4693
rect 3213 4687 3227 4701
rect 3353 4707 3367 4721
rect 3233 4679 3247 4693
rect 3313 4679 3327 4693
rect 3333 4687 3347 4701
rect 3373 4687 3387 4701
rect 3633 4707 3647 4721
rect 3453 4667 3467 4681
rect 3593 4679 3607 4693
rect 3613 4687 3627 4701
rect 3653 4687 3667 4701
rect 3793 4693 3807 4707
rect 3873 4707 3887 4721
rect 3473 4659 3487 4673
rect 3493 4647 3507 4661
rect 3513 4659 3527 4673
rect 3733 4667 3747 4681
rect 3753 4659 3767 4673
rect 3773 4647 3787 4661
rect 3793 4659 3807 4673
rect 3853 4687 3867 4701
rect 3893 4687 3907 4701
rect 4013 4707 4027 4721
rect 3913 4679 3927 4693
rect 3993 4687 4007 4701
rect 4033 4687 4047 4701
rect 4053 4679 4067 4693
rect 3853 4653 3867 4667
rect 4133 4647 4147 4661
rect 4153 4659 4167 4673
rect 4253 4667 4267 4681
rect 4273 4679 4287 4693
rect 4453 4707 4467 4721
rect 4553 4707 4567 4721
rect 4313 4667 4327 4681
rect 4413 4679 4427 4693
rect 4433 4687 4447 4701
rect 4473 4687 4487 4701
rect 4533 4687 4547 4701
rect 4573 4687 4587 4701
rect 4593 4679 4607 4693
rect 4773 4742 4787 4756
rect 4913 4736 4927 4750
rect 4673 4647 4687 4661
rect 4693 4659 4707 4673
rect 4773 4704 4787 4718
rect 4753 4639 4767 4653
rect 4833 4667 4847 4681
rect 4873 4667 4887 4681
rect 4773 4610 4787 4624
rect 5313 4713 5327 4727
rect 5373 4713 5387 4727
rect 5073 4687 5087 4701
rect 5013 4667 5027 4681
rect 5033 4659 5047 4673
rect 5053 4667 5067 4681
rect 5153 4679 5167 4693
rect 5173 4687 5187 4701
rect 4913 4610 4927 4624
rect 5193 4679 5207 4693
rect 5273 4679 5287 4693
rect 5293 4687 5307 4701
rect 5373 4693 5387 4707
rect 5313 4679 5327 4693
rect 5493 4713 5507 4727
rect 5533 4713 5547 4727
rect 5593 4713 5607 4727
rect 5653 4713 5667 4727
rect 5413 4679 5427 4693
rect 5433 4687 5447 4701
rect 5413 4633 5427 4647
rect 5453 4679 5467 4693
rect 5533 4679 5547 4693
rect 5553 4687 5567 4701
rect 5713 4707 5727 4721
rect 5573 4679 5587 4693
rect 5673 4679 5687 4693
rect 5693 4687 5707 4701
rect 5733 4687 5747 4701
rect 153 4513 167 4527
rect 193 4513 207 4527
rect 93 4459 107 4473
rect 113 4467 127 4481
rect 133 4459 147 4473
rect 273 4473 287 4487
rect 313 4473 327 4487
rect 333 4467 347 4481
rect 353 4479 367 4493
rect 373 4467 387 4481
rect 73 4439 87 4453
rect 213 4447 227 4461
rect 393 4459 407 4473
rect 533 4459 547 4473
rect 553 4467 567 4481
rect 573 4459 587 4473
rect 673 4459 687 4473
rect 693 4467 707 4481
rect 773 4479 787 4493
rect 713 4459 727 4473
rect 793 4467 807 4481
rect 873 4467 887 4481
rect 893 4479 907 4493
rect 913 4467 927 4481
rect 233 4439 247 4453
rect 273 4439 287 4453
rect 253 4419 267 4433
rect 513 4439 527 4453
rect 653 4439 667 4453
rect 933 4459 947 4473
rect 1033 4467 1047 4481
rect 1053 4479 1067 4493
rect 1133 4447 1147 4461
rect 1273 4459 1287 4473
rect 1293 4467 1307 4481
rect 1313 4479 1327 4493
rect 1333 4467 1347 4481
rect 1413 4467 1427 4481
rect 1433 4479 1447 4493
rect 1153 4439 1167 4453
rect 1193 4439 1207 4453
rect 1173 4419 1187 4433
rect 1493 4459 1507 4473
rect 1513 4467 1527 4481
rect 1533 4459 1547 4473
rect 1553 4439 1567 4453
rect 1653 4447 1667 4461
rect 1953 4493 1967 4507
rect 2013 4493 2027 4507
rect 1933 4479 1947 4493
rect 1673 4439 1687 4453
rect 1693 4447 1707 4461
rect 1773 4447 1787 4461
rect 1913 4459 1927 4473
rect 1793 4439 1807 4453
rect 1833 4439 1847 4453
rect 1813 4419 1827 4433
rect 1953 4459 1967 4473
rect 2033 4447 2047 4461
rect 2053 4439 2067 4453
rect 2093 4439 2107 4453
rect 2193 4447 2207 4461
rect 2073 4419 2087 4433
rect 2213 4439 2227 4453
rect 2253 4439 2267 4453
rect 2333 4447 2347 4461
rect 2733 4467 2747 4481
rect 2753 4479 2767 4493
rect 2853 4479 2867 4493
rect 2353 4439 2367 4453
rect 2373 4447 2387 4461
rect 2453 4447 2467 4461
rect 2233 4419 2247 4433
rect 2473 4439 2487 4453
rect 2513 4439 2527 4453
rect 2573 4439 2587 4453
rect 2613 4439 2627 4453
rect 2633 4447 2647 4461
rect 2493 4419 2507 4433
rect 2593 4419 2607 4433
rect 2833 4459 2847 4473
rect 2873 4459 2887 4473
rect 3213 4479 3227 4493
rect 3233 4467 3247 4481
rect 2953 4447 2967 4461
rect 2973 4439 2987 4453
rect 3013 4439 3027 4453
rect 3093 4447 3107 4461
rect 2993 4419 3007 4433
rect 3113 4439 3127 4453
rect 3153 4439 3167 4453
rect 3133 4419 3147 4433
rect 3313 4459 3327 4473
rect 3333 4467 3347 4481
rect 3353 4459 3367 4473
rect 3473 4459 3487 4473
rect 3373 4439 3387 4453
rect 3493 4447 3507 4461
rect 3533 4459 3547 4473
rect 3613 4447 3627 4461
rect 3753 4467 3767 4481
rect 3633 4439 3647 4453
rect 3653 4447 3667 4461
rect 3813 4479 3827 4493
rect 3793 4459 3807 4473
rect 3873 4447 3887 4461
rect 3893 4439 3907 4453
rect 3913 4447 3927 4461
rect 4013 4459 4027 4473
rect 4053 4459 4067 4473
rect 4113 4459 4127 4473
rect 4153 4447 4167 4461
rect 4173 4459 4187 4473
rect 4273 4447 4287 4461
rect 4293 4439 4307 4453
rect 4313 4447 4327 4461
rect 4413 4459 4427 4473
rect 4433 4467 4447 4481
rect 4453 4459 4467 4473
rect 4393 4439 4407 4453
rect 4513 4447 4527 4461
rect 4533 4439 4547 4453
rect 4553 4447 4567 4461
rect 4653 4447 4667 4461
rect 4753 4479 4767 4493
rect 5113 4516 5127 4530
rect 4773 4467 4787 4481
rect 4673 4439 4687 4453
rect 4693 4447 4707 4461
rect 4853 4447 4867 4461
rect 5253 4516 5267 4530
rect 4873 4439 4887 4453
rect 4893 4447 4907 4461
rect 4973 4459 4987 4473
rect 4993 4467 5007 4481
rect 5013 4459 5027 4473
rect 5093 4487 5107 4501
rect 5033 4439 5047 4453
rect 5113 4422 5127 4436
rect 5173 4459 5187 4473
rect 5213 4459 5227 4473
rect 5353 4459 5367 4473
rect 5373 4467 5387 4481
rect 5493 4479 5507 4493
rect 5393 4459 5407 4473
rect 5513 4459 5527 4473
rect 5413 4439 5427 4453
rect 5553 4467 5567 4481
rect 5113 4384 5127 4398
rect 5253 4390 5267 4404
rect 5673 4459 5687 4473
rect 5693 4467 5707 4481
rect 5713 4459 5727 4473
rect 5653 4439 5667 4453
rect 93 4207 107 4221
rect 233 4207 247 4221
rect 433 4227 447 4241
rect 113 4187 127 4201
rect 133 4179 147 4193
rect 153 4187 167 4201
rect 253 4187 267 4201
rect 273 4179 287 4193
rect 293 4187 307 4201
rect 393 4199 407 4213
rect 413 4207 427 4221
rect 453 4207 467 4221
rect 573 4227 587 4241
rect 533 4199 547 4213
rect 553 4207 567 4221
rect 593 4207 607 4221
rect 673 4179 687 4193
rect 493 4133 507 4147
rect 533 4133 547 4147
rect 813 4207 827 4221
rect 713 4187 727 4201
rect 833 4187 847 4201
rect 733 4167 747 4181
rect 853 4179 867 4193
rect 873 4187 887 4201
rect 1253 4227 1267 4241
rect 933 4167 947 4181
rect 953 4179 967 4193
rect 1053 4187 1067 4201
rect 1213 4199 1227 4213
rect 1233 4207 1247 4221
rect 1273 4207 1287 4221
rect 1353 4199 1367 4213
rect 1373 4207 1387 4221
rect 1073 4179 1087 4193
rect 1093 4167 1107 4181
rect 1113 4179 1127 4193
rect 1393 4199 1407 4213
rect 1473 4199 1487 4213
rect 1493 4207 1507 4221
rect 1513 4199 1527 4213
rect 1593 4187 1607 4201
rect 1753 4227 1767 4241
rect 1633 4187 1647 4201
rect 1713 4199 1727 4213
rect 1733 4207 1747 4221
rect 1773 4207 1787 4221
rect 1893 4227 1907 4241
rect 1993 4227 2007 4241
rect 1853 4199 1867 4213
rect 1873 4207 1887 4221
rect 1913 4207 1927 4221
rect 1973 4207 1987 4221
rect 2013 4207 2027 4221
rect 2133 4227 2147 4241
rect 2033 4199 2047 4213
rect 2113 4207 2127 4221
rect 2153 4207 2167 4221
rect 2173 4199 2187 4213
rect 1613 4167 1627 4181
rect 2273 4187 2287 4201
rect 2413 4207 2427 4221
rect 2613 4227 2627 4241
rect 2313 4187 2327 4201
rect 2433 4187 2447 4201
rect 2293 4167 2307 4181
rect 2453 4179 2467 4193
rect 2473 4187 2487 4201
rect 2573 4199 2587 4213
rect 2593 4207 2607 4221
rect 2633 4207 2647 4221
rect 2833 4227 2847 4241
rect 2813 4207 2827 4221
rect 2853 4207 2867 4221
rect 2873 4199 2887 4213
rect 2953 4199 2967 4213
rect 2973 4207 2987 4221
rect 2693 4167 2707 4181
rect 2713 4179 2727 4193
rect 2993 4199 3007 4213
rect 3413 4207 3427 4221
rect 3073 4179 3087 4193
rect 3093 4167 3107 4181
rect 3113 4179 3127 4193
rect 3133 4187 3147 4201
rect 3213 4179 3227 4193
rect 3233 4167 3247 4181
rect 3253 4179 3267 4193
rect 3273 4187 3287 4201
rect 3353 4187 3367 4201
rect 3373 4179 3387 4193
rect 3393 4187 3407 4201
rect 3633 4227 3647 4241
rect 3613 4207 3627 4221
rect 3653 4207 3667 4221
rect 3773 4227 3787 4241
rect 3673 4199 3687 4213
rect 3753 4207 3767 4221
rect 3793 4207 3807 4221
rect 3813 4199 3827 4213
rect 3913 4199 3927 4213
rect 3933 4207 3947 4221
rect 3513 4167 3527 4181
rect 3533 4179 3547 4193
rect 3953 4199 3967 4213
rect 4053 4199 4067 4213
rect 4073 4207 4087 4221
rect 4093 4199 4107 4213
rect 4173 4199 4187 4213
rect 4193 4207 4207 4221
rect 4213 4199 4227 4213
rect 4293 4207 4307 4221
rect 4313 4187 4327 4201
rect 4333 4179 4347 4193
rect 4353 4187 4367 4201
rect 4433 4187 4447 4201
rect 4413 4167 4427 4181
rect 4573 4207 4587 4221
rect 4773 4207 4787 4221
rect 4473 4179 4487 4193
rect 4593 4187 4607 4201
rect 4613 4179 4627 4193
rect 4633 4187 4647 4201
rect 4713 4187 4727 4201
rect 4733 4179 4747 4193
rect 4753 4187 4767 4201
rect 4853 4187 4867 4201
rect 4893 4187 4907 4201
rect 5053 4213 5067 4227
rect 5133 4213 5147 4227
rect 5293 4207 5307 4221
rect 4873 4167 4887 4181
rect 4973 4167 4987 4181
rect 4993 4179 5007 4193
rect 5093 4179 5107 4193
rect 5113 4167 5127 4181
rect 5133 4179 5147 4193
rect 5153 4187 5167 4201
rect 5233 4187 5247 4201
rect 5253 4179 5267 4193
rect 5273 4187 5287 4201
rect 5613 4256 5627 4270
rect 5753 4262 5767 4276
rect 5533 4207 5547 4221
rect 5373 4167 5387 4181
rect 5393 4179 5407 4193
rect 5473 4187 5487 4201
rect 5493 4179 5507 4193
rect 5513 4187 5527 4201
rect 5653 4187 5667 4201
rect 5693 4187 5707 4201
rect 5753 4224 5767 4238
rect 5773 4159 5787 4173
rect 5613 4130 5627 4144
rect 5753 4130 5767 4144
rect 153 4013 167 4027
rect 73 3987 87 4001
rect 93 3999 107 4013
rect 93 3933 107 3947
rect 133 3933 147 3947
rect 93 3913 107 3927
rect 173 3979 187 3993
rect 193 3987 207 4001
rect 213 3979 227 3993
rect 333 3987 347 4001
rect 353 3999 367 4013
rect 433 3987 447 4001
rect 453 3999 467 4013
rect 473 3987 487 4001
rect 613 3999 627 4013
rect 233 3959 247 3973
rect 493 3979 507 3993
rect 593 3979 607 3993
rect 633 3979 647 3993
rect 733 3987 747 4001
rect 753 3999 767 4013
rect 813 3979 827 3993
rect 833 3987 847 4001
rect 953 3999 967 4013
rect 853 3979 867 3993
rect 973 3987 987 4001
rect 873 3959 887 3973
rect 1053 3959 1067 3973
rect 1093 3959 1107 3973
rect 1113 3967 1127 3981
rect 1193 3979 1207 3993
rect 1213 3987 1227 4001
rect 1233 3979 1247 3993
rect 1253 3987 1267 4001
rect 1273 3979 1287 3993
rect 1073 3939 1087 3953
rect 1373 3967 1387 3981
rect 1653 4033 1667 4047
rect 1693 4033 1707 4047
rect 1513 3987 1527 4001
rect 1533 3999 1547 4013
rect 1633 3999 1647 4013
rect 1393 3959 1407 3973
rect 1413 3967 1427 3981
rect 1613 3979 1627 3993
rect 1653 3979 1667 3993
rect 1733 3987 1747 4001
rect 1753 3999 1767 4013
rect 1813 3959 1827 3973
rect 1853 3959 1867 3973
rect 1873 3967 1887 3981
rect 1993 3979 2007 3993
rect 2013 3987 2027 4001
rect 2033 3979 2047 3993
rect 1833 3939 1847 3953
rect 1973 3959 1987 3973
rect 2133 3967 2147 3981
rect 2153 3959 2167 3973
rect 2193 3959 2207 3973
rect 2253 3959 2267 3973
rect 2293 3959 2307 3973
rect 2313 3967 2327 3981
rect 2433 3979 2447 3993
rect 2453 3987 2467 4001
rect 2473 3979 2487 3993
rect 2173 3939 2187 3953
rect 2273 3939 2287 3953
rect 2413 3959 2427 3973
rect 2553 3967 2567 3981
rect 2593 4013 2607 4027
rect 2573 3959 2587 3973
rect 2593 3967 2607 3981
rect 2633 3973 2647 3987
rect 2613 3953 2627 3967
rect 2593 3933 2607 3947
rect 2653 3967 2667 3981
rect 3073 3987 3087 4001
rect 3093 3999 3107 4013
rect 2673 3959 2687 3973
rect 2693 3967 2707 3981
rect 2773 3959 2787 3973
rect 2813 3959 2827 3973
rect 2833 3967 2847 3981
rect 2793 3939 2807 3953
rect 2913 3959 2927 3973
rect 2953 3959 2967 3973
rect 2973 3967 2987 3981
rect 2933 3939 2947 3953
rect 3313 3987 3327 4001
rect 3333 3999 3347 4013
rect 3173 3967 3187 3981
rect 3193 3959 3207 3973
rect 3233 3959 3247 3973
rect 3213 3939 3227 3953
rect 3433 3979 3447 3993
rect 3453 3987 3467 4001
rect 3473 3979 3487 3993
rect 3413 3959 3427 3973
rect 3533 3967 3547 3981
rect 3673 3987 3687 4001
rect 3553 3959 3567 3973
rect 3573 3967 3587 3981
rect 3733 3999 3747 4013
rect 3713 3979 3727 3993
rect 3813 3967 3827 3981
rect 3833 3959 3847 3973
rect 3853 3967 3867 3981
rect 3973 3979 3987 3993
rect 3993 3987 4007 4001
rect 4013 3979 4027 3993
rect 4093 3979 4107 3993
rect 4113 3987 4127 4001
rect 4133 3999 4147 4013
rect 4153 3987 4167 4001
rect 3953 3959 3967 3973
rect 4213 3967 4227 3981
rect 4233 3959 4247 3973
rect 4253 3967 4267 3981
rect 4333 3979 4347 3993
rect 4353 3987 4367 4001
rect 4373 3979 4387 3993
rect 4473 3979 4487 3993
rect 4493 3987 4507 4001
rect 4613 3999 4627 4013
rect 4513 3979 4527 3993
rect 4633 3979 4647 3993
rect 4393 3959 4407 3973
rect 4533 3959 4547 3973
rect 4673 3987 4687 4001
rect 4773 3967 4787 3981
rect 5013 3999 5027 4013
rect 5213 4036 5227 4050
rect 5353 4036 5367 4050
rect 5033 3987 5047 4001
rect 5133 3987 5147 4001
rect 5153 3999 5167 4013
rect 5193 4007 5207 4021
rect 4793 3959 4807 3973
rect 4813 3967 4827 3981
rect 4873 3959 4887 3973
rect 4913 3959 4927 3973
rect 4933 3967 4947 3981
rect 4893 3939 4907 3953
rect 5213 3942 5227 3956
rect 5273 3979 5287 3993
rect 5313 3979 5327 3993
rect 5213 3904 5227 3918
rect 5353 3910 5367 3924
rect 5453 4036 5467 4050
rect 5593 4036 5607 4050
rect 5433 4007 5447 4021
rect 5453 3942 5467 3956
rect 5513 3979 5527 3993
rect 5553 3979 5567 3993
rect 5693 3979 5707 3993
rect 5713 3987 5727 4001
rect 5733 3979 5747 3993
rect 5753 3959 5767 3973
rect 5453 3904 5467 3918
rect 5593 3910 5607 3924
rect 73 3719 87 3733
rect 93 3727 107 3741
rect 233 3747 247 3761
rect 113 3719 127 3733
rect 193 3719 207 3733
rect 213 3727 227 3741
rect 253 3727 267 3741
rect 553 3727 567 3741
rect 353 3699 367 3713
rect 393 3707 407 3721
rect 413 3699 427 3713
rect 453 3707 467 3721
rect 573 3707 587 3721
rect 593 3699 607 3713
rect 613 3707 627 3721
rect 693 3719 707 3733
rect 713 3727 727 3741
rect 733 3719 747 3733
rect 853 3727 867 3741
rect 1253 3747 1267 3761
rect 793 3707 807 3721
rect 813 3699 827 3713
rect 833 3707 847 3721
rect 973 3707 987 3721
rect 993 3699 1007 3713
rect 1013 3707 1027 3721
rect 1033 3699 1047 3713
rect 1053 3707 1067 3721
rect 1113 3719 1127 3733
rect 1133 3727 1147 3741
rect 1153 3719 1167 3733
rect 1233 3727 1247 3741
rect 1273 3727 1287 3741
rect 1353 3733 1367 3747
rect 1413 3733 1427 3747
rect 1293 3719 1307 3733
rect 1573 3727 1587 3741
rect 1373 3699 1387 3713
rect 1393 3687 1407 3701
rect 1413 3699 1427 3713
rect 1433 3707 1447 3721
rect 1513 3707 1527 3721
rect 1533 3699 1547 3713
rect 1553 3707 1567 3721
rect 1773 3719 1787 3733
rect 1793 3727 1807 3741
rect 1653 3687 1667 3701
rect 1673 3699 1687 3713
rect 1813 3719 1827 3733
rect 1873 3719 1887 3733
rect 1893 3727 1907 3741
rect 1913 3719 1927 3733
rect 2013 3707 2027 3721
rect 1993 3687 2007 3701
rect 2273 3747 2287 3761
rect 2133 3719 2147 3733
rect 2153 3727 2167 3741
rect 2053 3699 2067 3713
rect 2173 3719 2187 3733
rect 2253 3727 2267 3741
rect 2293 3727 2307 3741
rect 2313 3719 2327 3733
rect 2413 3727 2427 3741
rect 2433 3707 2447 3721
rect 2453 3699 2467 3713
rect 2473 3707 2487 3721
rect 2533 3719 2547 3733
rect 2553 3727 2567 3741
rect 2573 3719 2587 3733
rect 2713 3727 2727 3741
rect 2653 3707 2667 3721
rect 2673 3699 2687 3713
rect 2693 3707 2707 3721
rect 2913 3727 2927 3741
rect 3073 3753 3087 3767
rect 3193 3753 3207 3767
rect 2813 3699 2827 3713
rect 2933 3707 2947 3721
rect 2833 3687 2847 3701
rect 2953 3699 2967 3713
rect 2973 3707 2987 3721
rect 3033 3719 3047 3733
rect 3053 3727 3067 3741
rect 3073 3719 3087 3733
rect 3193 3719 3207 3733
rect 3213 3727 3227 3741
rect 3233 3719 3247 3733
rect 3353 3773 3367 3787
rect 3393 3773 3407 3787
rect 3413 3747 3427 3761
rect 3393 3727 3407 3741
rect 3433 3727 3447 3741
rect 3453 3719 3467 3733
rect 3313 3699 3327 3713
rect 3333 3687 3347 3701
rect 3533 3687 3547 3701
rect 3553 3699 3567 3713
rect 3653 3707 3667 3721
rect 3693 3707 3707 3721
rect 3773 3719 3787 3733
rect 3793 3727 3807 3741
rect 3673 3687 3687 3701
rect 3813 3719 3827 3733
rect 4093 3782 4107 3796
rect 4233 3776 4247 3790
rect 3893 3687 3907 3701
rect 3913 3699 3927 3713
rect 4013 3699 4027 3713
rect 4033 3687 4047 3701
rect 4093 3744 4107 3758
rect 4073 3679 4087 3693
rect 4153 3707 4167 3721
rect 4193 3707 4207 3721
rect 4093 3650 4107 3664
rect 4353 3707 4367 3721
rect 4373 3699 4387 3713
rect 4393 3707 4407 3721
rect 4413 3699 4427 3713
rect 4433 3707 4447 3721
rect 4493 3719 4507 3733
rect 4513 3727 4527 3741
rect 4533 3719 4547 3733
rect 4613 3707 4627 3721
rect 4793 3727 4807 3741
rect 4833 3733 4847 3747
rect 4873 3733 4887 3747
rect 4653 3707 4667 3721
rect 4733 3707 4747 3721
rect 4633 3687 4647 3701
rect 4753 3699 4767 3713
rect 4773 3707 4787 3721
rect 4233 3650 4247 3664
rect 4873 3699 4887 3713
rect 4893 3707 4907 3721
rect 5013 3719 5027 3733
rect 5033 3727 5047 3741
rect 5053 3719 5067 3733
rect 5453 3782 5467 3796
rect 5593 3776 5607 3790
rect 5113 3687 5127 3701
rect 5133 3699 5147 3713
rect 5233 3699 5247 3713
rect 5373 3699 5387 3713
rect 5453 3744 5467 3758
rect 5433 3679 5447 3693
rect 5513 3707 5527 3721
rect 5553 3707 5567 3721
rect 5453 3650 5467 3664
rect 5713 3719 5727 3733
rect 5733 3727 5747 3741
rect 5753 3719 5767 3733
rect 5593 3650 5607 3664
rect 73 3513 87 3527
rect 93 3499 107 3513
rect 113 3507 127 3521
rect 133 3499 147 3513
rect 193 3507 207 3521
rect 213 3519 227 3533
rect 233 3507 247 3521
rect 333 3519 347 3533
rect 253 3499 267 3513
rect 353 3507 367 3521
rect 73 3479 87 3493
rect 73 3433 87 3447
rect 433 3499 447 3513
rect 453 3507 467 3521
rect 473 3499 487 3513
rect 493 3479 507 3493
rect 573 3479 587 3493
rect 613 3479 627 3493
rect 633 3487 647 3501
rect 753 3487 767 3501
rect 593 3459 607 3473
rect 773 3479 787 3493
rect 793 3487 807 3501
rect 873 3487 887 3501
rect 893 3479 907 3493
rect 913 3487 927 3501
rect 973 3499 987 3513
rect 993 3507 1007 3521
rect 1013 3499 1027 3513
rect 1213 3513 1227 3527
rect 1033 3479 1047 3493
rect 1133 3487 1147 3501
rect 1153 3479 1167 3493
rect 1193 3479 1207 3493
rect 1173 3459 1187 3473
rect 1253 3487 1267 3501
rect 1273 3479 1287 3493
rect 1293 3487 1307 3501
rect 1393 3487 1407 3501
rect 1513 3499 1527 3513
rect 1533 3507 1547 3521
rect 1553 3499 1567 3513
rect 1673 3499 1687 3513
rect 1693 3507 1707 3521
rect 1713 3519 1727 3533
rect 1733 3507 1747 3521
rect 1933 3507 1947 3521
rect 1953 3519 1967 3533
rect 1973 3507 1987 3521
rect 2153 3533 2167 3547
rect 2193 3533 2207 3547
rect 1253 3453 1267 3467
rect 1413 3479 1427 3493
rect 1453 3479 1467 3493
rect 1433 3459 1447 3473
rect 1573 3479 1587 3493
rect 1813 3487 1827 3501
rect 1993 3499 2007 3513
rect 2113 3499 2127 3513
rect 2133 3507 2147 3521
rect 2153 3499 2167 3513
rect 2233 3499 2247 3513
rect 2253 3507 2267 3521
rect 2273 3499 2287 3513
rect 2393 3499 2407 3513
rect 2413 3507 2427 3521
rect 2433 3519 2447 3533
rect 2453 3507 2467 3521
rect 2533 3499 2547 3513
rect 1833 3479 1847 3493
rect 1873 3479 1887 3493
rect 1853 3459 1867 3473
rect 2093 3479 2107 3493
rect 2293 3479 2307 3493
rect 2553 3487 2567 3501
rect 2593 3499 2607 3513
rect 2653 3487 2667 3501
rect 2673 3479 2687 3493
rect 2693 3487 2707 3501
rect 2813 3499 2827 3513
rect 2833 3507 2847 3521
rect 2853 3499 2867 3513
rect 2953 3499 2967 3513
rect 2793 3479 2807 3493
rect 2993 3499 3007 3513
rect 3073 3487 3087 3501
rect 3393 3513 3407 3527
rect 3433 3513 3447 3527
rect 3093 3479 3107 3493
rect 3113 3487 3127 3501
rect 3173 3479 3187 3493
rect 3213 3479 3227 3493
rect 3233 3487 3247 3501
rect 3333 3487 3347 3501
rect 3493 3499 3507 3513
rect 3513 3507 3527 3521
rect 3533 3499 3547 3513
rect 3633 3499 3647 3513
rect 3653 3507 3667 3521
rect 3673 3499 3687 3513
rect 3753 3499 3767 3513
rect 3193 3459 3207 3473
rect 3353 3479 3367 3493
rect 3393 3479 3407 3493
rect 3473 3479 3487 3493
rect 3373 3459 3387 3473
rect 3613 3479 3627 3493
rect 3773 3487 3787 3501
rect 3893 3519 3907 3533
rect 3813 3499 3827 3513
rect 3873 3499 3887 3513
rect 3913 3499 3927 3513
rect 4053 3499 4067 3513
rect 4073 3507 4087 3521
rect 4153 3519 4167 3533
rect 4093 3499 4107 3513
rect 4173 3507 4187 3521
rect 4033 3479 4047 3493
rect 4253 3499 4267 3513
rect 4273 3507 4287 3521
rect 4333 3533 4347 3547
rect 4393 3533 4407 3547
rect 4293 3499 4307 3513
rect 4313 3479 4327 3493
rect 4413 3487 4427 3501
rect 4633 3556 4647 3570
rect 4433 3479 4447 3493
rect 4453 3487 4467 3501
rect 4513 3487 4527 3501
rect 4773 3556 4787 3570
rect 4613 3527 4627 3541
rect 4533 3479 4547 3493
rect 4553 3487 4567 3501
rect 4633 3462 4647 3476
rect 4693 3499 4707 3513
rect 4733 3499 4747 3513
rect 4893 3487 4907 3501
rect 5273 3556 5287 3570
rect 4913 3479 4927 3493
rect 4933 3487 4947 3501
rect 5033 3499 5047 3513
rect 5053 3507 5067 3521
rect 5073 3499 5087 3513
rect 5013 3479 5027 3493
rect 4633 3424 4647 3438
rect 4773 3430 4787 3444
rect 5153 3487 5167 3501
rect 5173 3479 5187 3493
rect 5193 3487 5207 3501
rect 5413 3556 5427 3570
rect 5313 3499 5327 3513
rect 5353 3499 5367 3513
rect 5433 3527 5447 3541
rect 5413 3462 5427 3476
rect 5533 3487 5547 3501
rect 5553 3479 5567 3493
rect 5573 3487 5587 3501
rect 5633 3499 5647 3513
rect 5653 3507 5667 3521
rect 5673 3499 5687 3513
rect 5273 3430 5287 3444
rect 5413 3424 5427 3438
rect 5693 3479 5707 3493
rect 93 3253 107 3267
rect 73 3219 87 3233
rect 93 3207 107 3221
rect 93 3173 107 3187
rect 173 3247 187 3261
rect 193 3227 207 3241
rect 213 3219 227 3233
rect 233 3227 247 3241
rect 393 3239 407 3253
rect 413 3247 427 3261
rect 313 3219 327 3233
rect 333 3207 347 3221
rect 433 3239 447 3253
rect 513 3219 527 3233
rect 533 3207 547 3221
rect 553 3219 567 3233
rect 573 3227 587 3241
rect 653 3227 667 3241
rect 693 3239 707 3253
rect 713 3227 727 3241
rect 833 3239 847 3253
rect 853 3247 867 3261
rect 993 3267 1007 3281
rect 873 3239 887 3253
rect 953 3239 967 3253
rect 973 3247 987 3261
rect 1013 3247 1027 3261
rect 1133 3267 1147 3281
rect 1093 3239 1107 3253
rect 1113 3247 1127 3261
rect 1153 3247 1167 3261
rect 1213 3219 1227 3233
rect 1233 3207 1247 3221
rect 1253 3219 1267 3233
rect 1273 3227 1287 3241
rect 1513 3267 1527 3281
rect 1473 3239 1487 3253
rect 1493 3247 1507 3261
rect 1533 3247 1547 3261
rect 1653 3267 1667 3281
rect 1853 3293 1867 3307
rect 1893 3293 1907 3307
rect 1613 3239 1627 3253
rect 1633 3247 1647 3261
rect 1673 3247 1687 3261
rect 1373 3219 1387 3233
rect 1393 3207 1407 3221
rect 1753 3227 1767 3241
rect 1913 3239 1927 3253
rect 1933 3247 1947 3261
rect 1773 3219 1787 3233
rect 1793 3207 1807 3221
rect 1813 3219 1827 3233
rect 1953 3239 1967 3253
rect 2033 3227 2047 3241
rect 2153 3239 2167 3253
rect 2173 3247 2187 3261
rect 2053 3219 2067 3233
rect 2073 3207 2087 3221
rect 2093 3219 2107 3233
rect 2193 3239 2207 3253
rect 2293 3227 2307 3241
rect 2313 3239 2327 3253
rect 2353 3227 2367 3241
rect 2413 3239 2427 3253
rect 2433 3247 2447 3261
rect 2453 3239 2467 3253
rect 2553 3247 2567 3261
rect 2833 3267 2847 3281
rect 2813 3247 2827 3261
rect 2853 3247 2867 3261
rect 2973 3267 2987 3281
rect 2573 3227 2587 3241
rect 2593 3219 2607 3233
rect 2613 3227 2627 3241
rect 2693 3227 2707 3241
rect 2873 3239 2887 3253
rect 2953 3247 2967 3261
rect 2993 3247 3007 3261
rect 3013 3239 3027 3253
rect 3113 3239 3127 3253
rect 3133 3247 3147 3261
rect 2713 3219 2727 3233
rect 2733 3207 2747 3221
rect 2753 3219 2767 3233
rect 2793 3213 2807 3227
rect 2833 3213 2847 3227
rect 2933 3213 2947 3227
rect 2973 3213 2987 3227
rect 2873 3173 2887 3187
rect 2933 3173 2947 3187
rect 3153 3239 3167 3253
rect 3253 3239 3267 3253
rect 3273 3247 3287 3261
rect 3293 3239 3307 3253
rect 3513 3267 3527 3281
rect 3473 3239 3487 3253
rect 3493 3247 3507 3261
rect 3533 3247 3547 3261
rect 3753 3247 3767 3261
rect 3353 3207 3367 3221
rect 3373 3219 3387 3233
rect 3593 3219 3607 3233
rect 3613 3207 3627 3221
rect 3633 3219 3647 3233
rect 3653 3227 3667 3241
rect 3773 3227 3787 3241
rect 3793 3219 3807 3233
rect 3813 3227 3827 3241
rect 3973 3302 3987 3316
rect 4113 3296 4127 3310
rect 3873 3207 3887 3221
rect 3893 3219 3907 3233
rect 3973 3264 3987 3278
rect 3953 3199 3967 3213
rect 4493 3302 4507 3316
rect 4633 3296 4647 3310
rect 4033 3227 4047 3241
rect 4073 3227 4087 3241
rect 3973 3170 3987 3184
rect 4273 3247 4287 3261
rect 4413 3247 4427 3261
rect 4213 3227 4227 3241
rect 4233 3219 4247 3233
rect 4253 3227 4267 3241
rect 4353 3227 4367 3241
rect 4373 3219 4387 3233
rect 4393 3227 4407 3241
rect 4493 3264 4507 3278
rect 4113 3170 4127 3184
rect 4473 3199 4487 3213
rect 4553 3227 4567 3241
rect 4593 3227 4607 3241
rect 4493 3170 4507 3184
rect 4793 3247 4807 3261
rect 4733 3227 4747 3241
rect 4753 3219 4767 3233
rect 4773 3227 4787 3241
rect 4893 3239 4907 3253
rect 4913 3247 4927 3261
rect 4933 3239 4947 3253
rect 5013 3247 5027 3261
rect 5033 3227 5047 3241
rect 5053 3219 5067 3233
rect 5073 3227 5087 3241
rect 5253 3239 5267 3253
rect 5273 3247 5287 3261
rect 5153 3219 5167 3233
rect 4633 3170 4647 3184
rect 5173 3207 5187 3221
rect 5293 3239 5307 3253
rect 5533 3247 5547 3261
rect 5353 3207 5367 3221
rect 5373 3219 5387 3233
rect 5473 3227 5487 3241
rect 5493 3219 5507 3233
rect 5513 3227 5527 3241
rect 5653 3239 5667 3253
rect 5673 3247 5687 3261
rect 5693 3239 5707 3253
rect 93 3019 107 3033
rect 113 3007 127 3021
rect 153 3019 167 3033
rect 233 2999 247 3013
rect 273 2999 287 3013
rect 293 3007 307 3021
rect 373 3007 387 3021
rect 253 2979 267 2993
rect 393 2999 407 3013
rect 413 3007 427 3021
rect 533 3019 547 3033
rect 553 3027 567 3041
rect 573 3019 587 3033
rect 633 3019 647 3033
rect 653 3027 667 3041
rect 673 3019 687 3033
rect 773 3019 787 3033
rect 793 3027 807 3041
rect 813 3019 827 3033
rect 913 3019 927 3033
rect 933 3027 947 3041
rect 973 3033 987 3047
rect 1013 3033 1027 3047
rect 953 3019 967 3033
rect 513 2999 527 3013
rect 693 2999 707 3013
rect 833 2999 847 3013
rect 973 2999 987 3013
rect 1073 3007 1087 3021
rect 1233 3039 1247 3053
rect 1093 2999 1107 3013
rect 1113 3007 1127 3021
rect 1213 3019 1227 3033
rect 1253 3019 1267 3033
rect 1313 3019 1327 3033
rect 1333 3027 1347 3041
rect 1353 3019 1367 3033
rect 1373 2999 1387 3013
rect 1473 3007 1487 3021
rect 1633 3019 1647 3033
rect 1653 3027 1667 3041
rect 1673 3039 1687 3053
rect 1693 3027 1707 3041
rect 1793 3019 1807 3033
rect 1813 3027 1827 3041
rect 1833 3019 1847 3033
rect 1893 3019 1907 3033
rect 1913 3027 1927 3041
rect 1933 3019 1947 3033
rect 2093 3019 2107 3033
rect 2113 3027 2127 3041
rect 2133 3019 2147 3033
rect 2233 3019 2247 3033
rect 2253 3027 2267 3041
rect 2273 3019 2287 3033
rect 2373 3019 2387 3033
rect 2393 3027 2407 3041
rect 2413 3039 2427 3053
rect 2433 3027 2447 3041
rect 2513 3019 2527 3033
rect 2533 3027 2547 3041
rect 2553 3039 2567 3053
rect 2573 3027 2587 3041
rect 2653 3019 2667 3033
rect 2673 3027 2687 3041
rect 2693 3019 2707 3033
rect 2713 3027 2727 3041
rect 2733 3019 2747 3033
rect 2813 3027 2827 3041
rect 1493 2999 1507 3013
rect 1533 2999 1547 3013
rect 1513 2979 1527 2993
rect 1773 2999 1787 3013
rect 1953 2999 1967 3013
rect 2073 2999 2087 3013
rect 2213 2999 2227 3013
rect 2533 2993 2547 3007
rect 2593 2993 2607 3007
rect 2873 3039 2887 3053
rect 2953 3039 2967 3053
rect 2853 3019 2867 3033
rect 2933 3019 2947 3033
rect 2973 3019 2987 3033
rect 3073 3007 3087 3021
rect 3093 2999 3107 3013
rect 3113 3007 3127 3021
rect 3153 3009 3167 3023
rect 3213 3019 3227 3033
rect 3233 3007 3247 3021
rect 3333 3039 3347 3053
rect 3273 3019 3287 3033
rect 3353 3019 3367 3033
rect 3393 3027 3407 3041
rect 3513 3019 3527 3033
rect 3533 3027 3547 3041
rect 3553 3019 3567 3033
rect 3653 3019 3667 3033
rect 3673 3027 3687 3041
rect 3693 3019 3707 3033
rect 3773 3027 3787 3041
rect 3493 2999 3507 3013
rect 3633 2999 3647 3013
rect 3833 3039 3847 3053
rect 3813 3019 3827 3033
rect 3933 3019 3947 3033
rect 3953 3007 3967 3021
rect 4313 3076 4327 3090
rect 4073 3039 4087 3053
rect 3993 3019 4007 3033
rect 4053 3019 4067 3033
rect 4093 3019 4107 3033
rect 4173 2999 4187 3013
rect 4213 2999 4227 3013
rect 4233 3007 4247 3021
rect 4193 2979 4207 2993
rect 4453 3076 4467 3090
rect 4353 3019 4367 3033
rect 4393 3019 4407 3033
rect 4473 3047 4487 3061
rect 4453 2982 4467 2996
rect 4573 3019 4587 3033
rect 4593 3027 4607 3041
rect 4613 3019 4627 3033
rect 4713 3019 4727 3033
rect 4733 3027 4747 3041
rect 4753 3019 4767 3033
rect 4633 2999 4647 3013
rect 4773 2999 4787 3013
rect 4873 3007 4887 3021
rect 5093 3076 5107 3090
rect 4893 2999 4907 3013
rect 4913 3007 4927 3021
rect 4973 3007 4987 3021
rect 4993 2999 5007 3013
rect 5013 3007 5027 3021
rect 4313 2950 4327 2964
rect 4453 2944 4467 2958
rect 5233 3076 5247 3090
rect 5573 3076 5587 3090
rect 5133 3019 5147 3033
rect 5173 3019 5187 3033
rect 5253 3047 5267 3061
rect 5233 2982 5247 2996
rect 5713 3076 5727 3090
rect 5353 3027 5367 3041
rect 5553 3047 5567 3061
rect 5493 3027 5507 3041
rect 5093 2950 5107 2964
rect 5233 2944 5247 2958
rect 5573 2982 5587 2996
rect 5633 3019 5647 3033
rect 5673 3019 5687 3033
rect 5573 2944 5587 2958
rect 5713 2950 5727 2964
rect 4373 2884 4387 2887
rect 73 2759 87 2773
rect 93 2767 107 2781
rect 113 2759 127 2773
rect 233 2767 247 2781
rect 173 2747 187 2761
rect 193 2739 207 2753
rect 213 2747 227 2761
rect 333 2739 347 2753
rect 353 2727 367 2741
rect 413 2739 427 2753
rect 433 2727 447 2741
rect 453 2739 467 2753
rect 473 2747 487 2761
rect 573 2759 587 2773
rect 593 2767 607 2781
rect 613 2759 627 2773
rect 673 2747 687 2761
rect 713 2759 727 2773
rect 733 2747 747 2761
rect 813 2759 827 2773
rect 833 2767 847 2781
rect 853 2759 867 2773
rect 933 2739 947 2753
rect 953 2727 967 2741
rect 973 2739 987 2753
rect 993 2747 1007 2761
rect 1073 2759 1087 2773
rect 1093 2767 1107 2781
rect 1113 2759 1127 2773
rect 1233 2767 1247 2781
rect 1413 2767 1427 2781
rect 1253 2747 1267 2761
rect 1273 2739 1287 2753
rect 1293 2747 1307 2761
rect 1353 2747 1367 2761
rect 1373 2739 1387 2753
rect 1393 2747 1407 2761
rect 1513 2739 1527 2753
rect 1553 2747 1567 2761
rect 1633 2747 1647 2761
rect 1673 2747 1687 2761
rect 1773 2747 1787 2761
rect 1793 2759 1807 2773
rect 1573 2727 1587 2741
rect 1653 2727 1667 2741
rect 1593 2693 1607 2707
rect 1633 2693 1647 2707
rect 1833 2747 1847 2761
rect 1933 2759 1947 2773
rect 1953 2767 1967 2781
rect 1973 2759 1987 2773
rect 2093 2767 2107 2781
rect 2033 2747 2047 2761
rect 2053 2739 2067 2753
rect 2073 2747 2087 2761
rect 2193 2747 2207 2761
rect 2213 2759 2227 2773
rect 2253 2747 2267 2761
rect 2333 2759 2347 2773
rect 2353 2767 2367 2781
rect 2373 2759 2387 2773
rect 2453 2747 2467 2761
rect 2633 2787 2647 2801
rect 2493 2747 2507 2761
rect 2593 2759 2607 2773
rect 2613 2767 2627 2781
rect 2653 2767 2667 2781
rect 2473 2727 2487 2741
rect 2393 2713 2407 2727
rect 2453 2713 2467 2727
rect 2733 2747 2747 2761
rect 2753 2759 2767 2773
rect 2933 2767 2947 2781
rect 3073 2787 3087 2801
rect 3193 2793 3207 2807
rect 3233 2793 3247 2807
rect 2793 2747 2807 2761
rect 2873 2747 2887 2761
rect 2893 2739 2907 2753
rect 2913 2747 2927 2761
rect 3033 2759 3047 2773
rect 3053 2767 3067 2781
rect 3093 2767 3107 2781
rect 3153 2759 3167 2773
rect 3173 2767 3187 2781
rect 3193 2759 3207 2773
rect 3293 2767 3307 2781
rect 3313 2747 3327 2761
rect 3333 2739 3347 2753
rect 3353 2747 3367 2761
rect 3433 2747 3447 2761
rect 3453 2759 3467 2773
rect 3493 2747 3507 2761
rect 3553 2747 3567 2761
rect 3693 2787 3707 2801
rect 3673 2767 3687 2781
rect 3713 2767 3727 2781
rect 3593 2747 3607 2761
rect 3733 2759 3747 2773
rect 3813 2759 3827 2773
rect 3833 2767 3847 2781
rect 3573 2727 3587 2741
rect 3853 2759 3867 2773
rect 4053 2767 4067 2781
rect 4373 2873 4387 2884
rect 3953 2747 3967 2761
rect 3973 2739 3987 2753
rect 4073 2747 4087 2761
rect 4093 2739 4107 2753
rect 4113 2747 4127 2761
rect 4173 2759 4187 2773
rect 4193 2767 4207 2781
rect 4213 2759 4227 2773
rect 4293 2739 4307 2753
rect 4313 2747 4327 2761
rect 4493 2822 4507 2836
rect 4633 2816 4647 2830
rect 4393 2727 4407 2741
rect 4413 2739 4427 2753
rect 4493 2784 4507 2798
rect 4473 2719 4487 2733
rect 4553 2747 4567 2761
rect 4593 2747 4607 2761
rect 4493 2690 4507 2704
rect 4633 2690 4647 2704
rect 4733 2816 4747 2830
rect 4873 2822 4887 2836
rect 4773 2747 4787 2761
rect 4813 2747 4827 2761
rect 4873 2784 4887 2798
rect 5373 2822 5387 2836
rect 5513 2816 5527 2830
rect 5053 2767 5067 2781
rect 4993 2747 5007 2761
rect 5013 2739 5027 2753
rect 5033 2747 5047 2761
rect 5133 2759 5147 2773
rect 5153 2767 5167 2781
rect 4893 2719 4907 2733
rect 4733 2690 4747 2704
rect 4873 2690 4887 2704
rect 5173 2759 5187 2773
rect 5253 2739 5267 2753
rect 5293 2739 5307 2753
rect 5373 2784 5387 2798
rect 5353 2719 5367 2733
rect 5433 2747 5447 2761
rect 5473 2747 5487 2761
rect 5373 2690 5387 2704
rect 5673 2767 5687 2781
rect 5613 2747 5627 2761
rect 5633 2739 5647 2753
rect 5653 2747 5667 2761
rect 5513 2690 5527 2704
rect 73 2547 87 2561
rect 93 2559 107 2573
rect 153 2559 167 2573
rect 173 2547 187 2561
rect 273 2539 287 2553
rect 293 2547 307 2561
rect 313 2559 327 2573
rect 333 2547 347 2561
rect 533 2559 547 2573
rect 553 2547 567 2561
rect 653 2559 667 2573
rect 393 2519 407 2533
rect 433 2519 447 2533
rect 453 2527 467 2541
rect 413 2499 427 2513
rect 633 2539 647 2553
rect 673 2539 687 2553
rect 753 2539 767 2553
rect 773 2547 787 2561
rect 793 2539 807 2553
rect 913 2547 927 2561
rect 933 2559 947 2573
rect 953 2547 967 2561
rect 973 2539 987 2553
rect 1093 2539 1107 2553
rect 1113 2547 1127 2561
rect 1133 2539 1147 2553
rect 813 2519 827 2533
rect 1073 2519 1087 2533
rect 1213 2527 1227 2541
rect 1233 2519 1247 2533
rect 1253 2527 1267 2541
rect 1313 2539 1327 2553
rect 1353 2527 1367 2541
rect 1373 2539 1387 2553
rect 1593 2559 1607 2573
rect 1613 2547 1627 2561
rect 1473 2527 1487 2541
rect 1493 2519 1507 2533
rect 1533 2519 1547 2533
rect 1513 2499 1527 2513
rect 1693 2539 1707 2553
rect 1713 2547 1727 2561
rect 1793 2553 1807 2567
rect 1733 2539 1747 2553
rect 1753 2519 1767 2533
rect 1873 2539 1887 2553
rect 1893 2547 1907 2561
rect 1913 2539 1927 2553
rect 1973 2539 1987 2553
rect 1993 2547 2007 2561
rect 2013 2539 2027 2553
rect 2813 2593 2827 2607
rect 1853 2519 1867 2533
rect 2033 2519 2047 2533
rect 2133 2527 2147 2541
rect 2273 2539 2287 2553
rect 2293 2547 2307 2561
rect 2313 2559 2327 2573
rect 2333 2547 2347 2561
rect 1753 2473 1767 2487
rect 1813 2473 1827 2487
rect 1813 2453 1827 2467
rect 2153 2519 2167 2533
rect 2193 2519 2207 2533
rect 2173 2499 2187 2513
rect 2393 2527 2407 2541
rect 2413 2519 2427 2533
rect 2433 2527 2447 2541
rect 2573 2539 2587 2553
rect 2593 2547 2607 2561
rect 2613 2539 2627 2553
rect 2673 2539 2687 2553
rect 2693 2547 2707 2561
rect 2713 2539 2727 2553
rect 2553 2519 2567 2533
rect 2733 2519 2747 2533
rect 2833 2539 2847 2553
rect 2853 2547 2867 2561
rect 2873 2559 2887 2573
rect 2893 2547 2907 2561
rect 2973 2547 2987 2561
rect 2993 2559 3007 2573
rect 2813 2513 2827 2527
rect 3053 2539 3067 2553
rect 3073 2547 3087 2561
rect 3173 2573 3187 2587
rect 3213 2573 3227 2587
rect 3113 2553 3127 2567
rect 3093 2539 3107 2553
rect 3193 2533 3207 2547
rect 3113 2519 3127 2533
rect 3213 2527 3227 2541
rect 3233 2519 3247 2533
rect 3253 2527 3267 2541
rect 3353 2527 3367 2541
rect 3473 2539 3487 2553
rect 3373 2519 3387 2533
rect 3413 2519 3427 2533
rect 3393 2499 3407 2513
rect 3513 2527 3527 2541
rect 3533 2539 3547 2553
rect 3613 2527 3627 2541
rect 3733 2573 3747 2587
rect 3633 2519 3647 2533
rect 3653 2527 3667 2541
rect 3713 2533 3727 2547
rect 3733 2539 3747 2553
rect 3753 2547 3767 2561
rect 3773 2539 3787 2553
rect 3793 2547 3807 2561
rect 3913 2559 3927 2573
rect 3813 2539 3827 2553
rect 3893 2539 3907 2553
rect 3933 2539 3947 2553
rect 3993 2547 4007 2561
rect 4133 2596 4147 2610
rect 4153 2596 4167 2610
rect 4173 2596 4187 2610
rect 4205 2596 4219 2610
rect 4233 2596 4247 2610
rect 4293 2593 4307 2607
rect 4313 2593 4327 2607
rect 4333 2593 4347 2607
rect 4073 2519 4087 2533
rect 4205 2543 4219 2557
rect 4253 2559 4267 2573
rect 4233 2525 4247 2539
rect 4373 2519 4387 2533
rect 4413 2527 4427 2541
rect 4133 2491 4147 2505
rect 4173 2491 4187 2505
rect 4153 2467 4167 2481
rect 4132 2452 4146 2466
rect 4313 2495 4327 2509
rect 4206 2470 4220 2484
rect 4233 2470 4247 2484
rect 4293 2453 4307 2467
rect 4313 2453 4327 2467
rect 4333 2453 4347 2467
rect 4553 2593 4567 2607
rect 4573 2593 4587 2607
rect 4593 2593 4607 2607
rect 4653 2596 4667 2610
rect 4681 2596 4695 2610
rect 4713 2596 4727 2610
rect 4733 2596 4747 2610
rect 4753 2596 4767 2610
rect 4633 2559 4647 2573
rect 4473 2527 4487 2541
rect 4681 2543 4695 2557
rect 4513 2519 4527 2533
rect 4653 2525 4667 2539
rect 4813 2519 4827 2533
rect 4573 2495 4587 2509
rect 4713 2491 4727 2505
rect 4753 2491 4767 2505
rect 4653 2470 4667 2484
rect 4680 2470 4694 2484
rect 4553 2453 4567 2467
rect 4573 2453 4587 2467
rect 4593 2453 4607 2467
rect 4733 2467 4747 2481
rect 4754 2452 4768 2466
rect 4973 2596 4987 2610
rect 4893 2547 4907 2561
rect 5113 2596 5127 2610
rect 5013 2539 5027 2553
rect 5053 2539 5067 2553
rect 5133 2567 5147 2581
rect 5113 2502 5127 2516
rect 5233 2547 5247 2561
rect 5373 2547 5387 2561
rect 5493 2547 5507 2561
rect 5633 2547 5647 2561
rect 5713 2547 5727 2561
rect 5733 2539 5747 2553
rect 4973 2470 4987 2484
rect 5113 2464 5127 2478
rect 2533 2404 2547 2407
rect 4353 2404 4367 2407
rect 4493 2404 4507 2407
rect 73 2267 87 2281
rect 233 2307 247 2321
rect 113 2267 127 2281
rect 193 2279 207 2293
rect 213 2287 227 2301
rect 253 2287 267 2301
rect 313 2279 327 2293
rect 333 2287 347 2301
rect 353 2279 367 2293
rect 493 2287 507 2301
rect 593 2287 607 2301
rect 793 2307 807 2321
rect 433 2267 447 2281
rect 453 2259 467 2273
rect 473 2267 487 2281
rect 613 2267 627 2281
rect 633 2259 647 2273
rect 653 2267 667 2281
rect 753 2279 767 2293
rect 773 2287 787 2301
rect 813 2287 827 2301
rect 893 2279 907 2293
rect 913 2287 927 2301
rect 933 2279 947 2293
rect 1013 2259 1027 2273
rect 1293 2307 1307 2321
rect 1053 2267 1067 2281
rect 1073 2247 1087 2261
rect 1133 2259 1147 2273
rect 1153 2267 1167 2281
rect 1253 2279 1267 2293
rect 1273 2287 1287 2301
rect 1313 2287 1327 2301
rect 1553 2287 1567 2301
rect 1873 2307 1887 2321
rect 1393 2267 1407 2281
rect 1413 2259 1427 2273
rect 1433 2247 1447 2261
rect 1453 2259 1467 2273
rect 1573 2267 1587 2281
rect 1593 2259 1607 2273
rect 1613 2267 1627 2281
rect 1693 2267 1707 2281
rect 1833 2279 1847 2293
rect 1853 2287 1867 2301
rect 1893 2287 1907 2301
rect 2013 2307 2027 2321
rect 1973 2279 1987 2293
rect 1993 2287 2007 2301
rect 2033 2287 2047 2301
rect 1713 2259 1727 2273
rect 1733 2247 1747 2261
rect 1753 2259 1767 2273
rect 2073 2259 2087 2273
rect 2212 2354 2226 2368
rect 2233 2339 2247 2353
rect 2373 2353 2387 2367
rect 2393 2353 2407 2367
rect 2413 2353 2427 2367
rect 2533 2393 2547 2404
rect 2286 2336 2300 2350
rect 2313 2336 2327 2350
rect 2213 2315 2227 2329
rect 2253 2315 2267 2329
rect 2393 2311 2407 2325
rect 2153 2287 2167 2301
rect 2313 2281 2327 2295
rect 2453 2287 2467 2301
rect 2285 2263 2299 2277
rect 2493 2279 2507 2293
rect 2333 2247 2347 2261
rect 2213 2210 2227 2224
rect 2233 2210 2247 2224
rect 2253 2210 2267 2224
rect 2285 2210 2299 2224
rect 2313 2210 2327 2224
rect 2373 2213 2387 2227
rect 2393 2213 2407 2227
rect 2413 2213 2427 2227
rect 2593 2267 2607 2281
rect 2773 2287 2787 2301
rect 2913 2287 2927 2301
rect 2633 2267 2647 2281
rect 2713 2267 2727 2281
rect 2733 2259 2747 2273
rect 2753 2267 2767 2281
rect 2853 2267 2867 2281
rect 2873 2259 2887 2273
rect 2893 2267 2907 2281
rect 3013 2279 3027 2293
rect 3033 2287 3047 2301
rect 3053 2279 3067 2293
rect 3133 2279 3147 2293
rect 3153 2287 3167 2301
rect 3253 2293 3267 2307
rect 3173 2279 3187 2293
rect 3213 2233 3227 2247
rect 3373 2313 3387 2327
rect 3453 2373 3467 2387
rect 3513 2373 3527 2387
rect 3293 2293 3307 2307
rect 3273 2267 3287 2281
rect 3293 2259 3307 2273
rect 3313 2247 3327 2261
rect 3333 2259 3347 2273
rect 3393 2267 3407 2281
rect 3593 2287 3607 2301
rect 3433 2267 3447 2281
rect 3533 2267 3547 2281
rect 3413 2247 3427 2261
rect 3553 2259 3567 2273
rect 3573 2267 3587 2281
rect 3673 2279 3687 2293
rect 3693 2287 3707 2301
rect 3713 2279 3727 2293
rect 3793 2267 3807 2281
rect 3833 2267 3847 2281
rect 3893 2259 3907 2273
rect 4032 2354 4046 2368
rect 4053 2339 4067 2353
rect 4193 2353 4207 2367
rect 4213 2353 4227 2367
rect 4233 2353 4247 2367
rect 4353 2393 4367 2404
rect 4106 2336 4120 2350
rect 4133 2336 4147 2350
rect 4033 2315 4047 2329
rect 4073 2315 4087 2329
rect 4213 2311 4227 2325
rect 3973 2287 3987 2301
rect 4133 2281 4147 2295
rect 4273 2287 4287 2301
rect 4105 2263 4119 2277
rect 4313 2279 4327 2293
rect 4153 2247 4167 2261
rect 4393 2267 4407 2281
rect 4033 2210 4047 2224
rect 4053 2210 4067 2224
rect 4073 2210 4087 2224
rect 4105 2210 4119 2224
rect 4133 2210 4147 2224
rect 4193 2213 4207 2227
rect 4213 2213 4227 2227
rect 4233 2213 4247 2227
rect 4493 2393 4507 2404
rect 4433 2279 4447 2293
rect 4453 2267 4467 2281
rect 4533 2267 4547 2281
rect 4553 2259 4567 2273
rect 4573 2267 4587 2281
rect 4593 2259 4607 2273
rect 4613 2267 4627 2281
rect 4693 2279 4707 2293
rect 4713 2287 4727 2301
rect 4733 2279 4747 2293
rect 4833 2267 4847 2281
rect 4873 2267 4887 2281
rect 5153 2313 5167 2327
rect 5193 2313 5207 2327
rect 4933 2247 4947 2261
rect 4953 2259 4967 2273
rect 5033 2267 5047 2281
rect 5053 2259 5067 2273
rect 5073 2267 5087 2281
rect 5093 2259 5107 2273
rect 5113 2267 5127 2281
rect 5193 2279 5207 2293
rect 5213 2287 5227 2301
rect 5253 2293 5267 2307
rect 5313 2293 5327 2307
rect 5233 2279 5247 2293
rect 5313 2259 5327 2273
rect 5333 2267 5347 2281
rect 5413 2279 5427 2293
rect 5433 2287 5447 2301
rect 5453 2279 5467 2293
rect 5533 2247 5547 2261
rect 5553 2259 5567 2273
rect 5633 2259 5647 2273
rect 5653 2267 5667 2281
rect 5693 2259 5707 2273
rect 5713 2267 5727 2281
rect 93 2059 107 2073
rect 133 2059 147 2073
rect 273 2073 287 2087
rect 333 2073 347 2087
rect 353 2067 367 2081
rect 373 2079 387 2093
rect 393 2067 407 2081
rect 233 2047 247 2061
rect 413 2059 427 2073
rect 513 2067 527 2081
rect 533 2079 547 2093
rect 253 2039 267 2053
rect 293 2039 307 2053
rect 273 2019 287 2033
rect 633 2059 647 2073
rect 653 2067 667 2081
rect 673 2059 687 2073
rect 753 2059 767 2073
rect 773 2067 787 2081
rect 793 2079 807 2093
rect 813 2067 827 2081
rect 853 2073 867 2087
rect 613 2039 627 2053
rect 813 2033 827 2047
rect 873 2039 887 2053
rect 913 2039 927 2053
rect 933 2047 947 2061
rect 1053 2047 1067 2061
rect 1213 2059 1227 2073
rect 1233 2067 1247 2081
rect 1253 2059 1267 2073
rect 1353 2059 1367 2073
rect 1373 2067 1387 2081
rect 1393 2059 1407 2073
rect 1473 2059 1487 2073
rect 1493 2067 1507 2081
rect 1513 2079 1527 2093
rect 1533 2067 1547 2081
rect 893 2019 907 2033
rect 1073 2039 1087 2053
rect 1113 2039 1127 2053
rect 1193 2039 1207 2053
rect 1093 2019 1107 2033
rect 1333 2039 1347 2053
rect 1613 2047 1627 2061
rect 1733 2059 1747 2073
rect 1753 2067 1767 2081
rect 1773 2059 1787 2073
rect 1873 2067 1887 2081
rect 1893 2079 1907 2093
rect 1913 2067 1927 2081
rect 1933 2059 1947 2073
rect 2053 2067 2067 2081
rect 1633 2039 1647 2053
rect 1673 2039 1687 2053
rect 1653 2019 1667 2033
rect 1793 2039 1807 2053
rect 2093 2059 2107 2073
rect 2113 2067 2127 2081
rect 2153 2059 2167 2073
rect 2353 2067 2367 2081
rect 2253 2047 2267 2061
rect 2273 2039 2287 2053
rect 2313 2039 2327 2053
rect 2293 2019 2307 2033
rect 2493 2116 2507 2130
rect 2513 2116 2527 2130
rect 2533 2116 2547 2130
rect 2565 2116 2579 2130
rect 2593 2116 2607 2130
rect 2653 2113 2667 2127
rect 2673 2113 2687 2127
rect 2693 2113 2707 2127
rect 2433 2039 2447 2053
rect 2565 2063 2579 2077
rect 2613 2079 2627 2093
rect 2593 2045 2607 2059
rect 2733 2039 2747 2053
rect 2773 2047 2787 2061
rect 2493 2011 2507 2025
rect 2533 2011 2547 2025
rect 2513 1987 2527 2001
rect 2492 1972 2506 1986
rect 2673 2015 2687 2029
rect 2566 1990 2580 2004
rect 2593 1990 2607 2004
rect 2653 1973 2667 1987
rect 2673 1973 2687 1987
rect 2693 1973 2707 1987
rect 2853 2059 2867 2073
rect 2873 2067 2887 2081
rect 2893 2059 2907 2073
rect 2913 2039 2927 2053
rect 3013 2047 3027 2061
rect 3033 2039 3047 2053
rect 3053 2047 3067 2061
rect 3113 2047 3127 2061
rect 3273 2079 3287 2093
rect 3133 2039 3147 2053
rect 3153 2047 3167 2061
rect 3253 2059 3267 2073
rect 2913 1993 2927 2007
rect 2993 1993 3007 2007
rect 3293 2059 3307 2073
rect 3393 2059 3407 2073
rect 3413 2047 3427 2061
rect 3453 2059 3467 2073
rect 3513 2067 3527 2081
rect 3533 2079 3547 2093
rect 3553 2067 3567 2081
rect 3573 2059 3587 2073
rect 3693 2059 3707 2073
rect 3713 2067 3727 2081
rect 3953 2067 3967 2081
rect 3713 2033 3727 2047
rect 3773 2033 3787 2047
rect 3793 2039 3807 2053
rect 3833 2039 3847 2053
rect 3853 2047 3867 2061
rect 3973 2059 3987 2073
rect 4093 2059 4107 2073
rect 3813 2019 3827 2033
rect 4113 2047 4127 2061
rect 4153 2059 4167 2073
rect 4233 2047 4247 2061
rect 4253 2039 4267 2053
rect 4273 2047 4287 2061
rect 4373 2059 4387 2073
rect 4393 2067 4407 2081
rect 4413 2059 4427 2073
rect 4473 2059 4487 2073
rect 4493 2067 4507 2081
rect 4513 2059 4527 2073
rect 4353 2039 4367 2053
rect 4533 2039 4547 2053
rect 4613 2047 4627 2061
rect 4633 2039 4647 2053
rect 4653 2047 4667 2061
rect 4733 2047 4747 2061
rect 4753 2039 4767 2053
rect 4773 2047 4787 2061
rect 4913 2059 4927 2073
rect 4933 2067 4947 2081
rect 4953 2059 4967 2073
rect 5053 2059 5067 2073
rect 5073 2067 5087 2081
rect 5153 2079 5167 2093
rect 5093 2059 5107 2073
rect 5173 2067 5187 2081
rect 5273 2079 5287 2093
rect 4893 2039 4907 2053
rect 5033 2039 5047 2053
rect 5253 2059 5267 2073
rect 5293 2059 5307 2073
rect 5373 2047 5387 2061
rect 5493 2079 5507 2093
rect 5513 2067 5527 2081
rect 5613 2067 5627 2081
rect 5633 2079 5647 2093
rect 5393 2039 5407 2053
rect 5413 2047 5427 2061
rect 5693 2059 5707 2073
rect 5713 2067 5727 2081
rect 5733 2059 5747 2073
rect 5753 2039 5767 2053
rect 2653 1924 2667 1927
rect 2773 1924 2787 1927
rect 113 1827 127 1841
rect 73 1799 87 1813
rect 93 1807 107 1821
rect 133 1807 147 1821
rect 353 1807 367 1821
rect 533 1827 547 1841
rect 193 1779 207 1793
rect 213 1767 227 1781
rect 233 1779 247 1793
rect 253 1787 267 1801
rect 373 1787 387 1801
rect 393 1779 407 1793
rect 413 1787 427 1801
rect 493 1799 507 1813
rect 513 1807 527 1821
rect 553 1807 567 1821
rect 653 1787 667 1801
rect 693 1787 707 1801
rect 673 1767 687 1781
rect 693 1753 707 1767
rect 793 1813 807 1827
rect 753 1779 767 1793
rect 773 1767 787 1781
rect 793 1779 807 1793
rect 813 1787 827 1801
rect 1053 1807 1067 1821
rect 1193 1807 1207 1821
rect 933 1779 947 1793
rect 1073 1787 1087 1801
rect 953 1767 967 1781
rect 1093 1779 1107 1793
rect 1113 1787 1127 1801
rect 1213 1787 1227 1801
rect 1233 1779 1247 1793
rect 1253 1787 1267 1801
rect 1433 1807 1447 1821
rect 1613 1807 1627 1821
rect 1713 1807 1727 1821
rect 1333 1779 1347 1793
rect 1453 1787 1467 1801
rect 1353 1767 1367 1781
rect 1473 1779 1487 1793
rect 1493 1787 1507 1801
rect 1553 1787 1567 1801
rect 1573 1779 1587 1793
rect 1593 1787 1607 1801
rect 1733 1787 1747 1801
rect 1753 1779 1767 1793
rect 1773 1787 1787 1801
rect 1853 1799 1867 1813
rect 1873 1807 1887 1821
rect 1893 1799 1907 1813
rect 1973 1799 1987 1813
rect 1993 1807 2007 1821
rect 2013 1799 2027 1813
rect 2113 1779 2127 1793
rect 2153 1779 2167 1793
rect 2193 1779 2207 1793
rect 2332 1874 2346 1888
rect 2353 1859 2367 1873
rect 2493 1873 2507 1887
rect 2513 1873 2527 1887
rect 2533 1873 2547 1887
rect 2653 1913 2667 1924
rect 2773 1913 2787 1924
rect 2406 1856 2420 1870
rect 2433 1856 2447 1870
rect 2333 1835 2347 1849
rect 2373 1835 2387 1849
rect 2513 1831 2527 1845
rect 2273 1807 2287 1821
rect 2433 1801 2447 1815
rect 2573 1807 2587 1821
rect 2405 1783 2419 1797
rect 2613 1799 2627 1813
rect 2453 1767 2467 1781
rect 2693 1799 2707 1813
rect 2713 1807 2727 1821
rect 2873 1827 2887 1841
rect 2333 1730 2347 1744
rect 2353 1730 2367 1744
rect 2373 1730 2387 1744
rect 2405 1730 2419 1744
rect 2433 1730 2447 1744
rect 2493 1733 2507 1747
rect 2513 1733 2527 1747
rect 2533 1733 2547 1747
rect 2733 1799 2747 1813
rect 2833 1799 2847 1813
rect 2853 1807 2867 1821
rect 2893 1807 2907 1821
rect 2973 1807 2987 1821
rect 2993 1787 3007 1801
rect 3013 1779 3027 1793
rect 3033 1787 3047 1801
rect 3093 1787 3107 1801
rect 3133 1787 3147 1801
rect 3113 1767 3127 1781
rect 3213 1779 3227 1793
rect 3233 1787 3247 1801
rect 3273 1779 3287 1793
rect 3293 1787 3307 1801
rect 3653 1807 3667 1821
rect 3813 1807 3827 1821
rect 3913 1813 3927 1827
rect 3393 1779 3407 1793
rect 3473 1787 3487 1801
rect 3413 1767 3427 1781
rect 3493 1779 3507 1793
rect 3513 1787 3527 1801
rect 3533 1779 3547 1793
rect 3553 1787 3567 1801
rect 3673 1787 3687 1801
rect 3693 1779 3707 1793
rect 3713 1787 3727 1801
rect 3833 1787 3847 1801
rect 3853 1779 3867 1793
rect 3873 1787 3887 1801
rect 3873 1753 3887 1767
rect 3993 1807 4007 1821
rect 3933 1787 3947 1801
rect 3953 1779 3967 1793
rect 3973 1787 3987 1801
rect 4093 1799 4107 1813
rect 4113 1807 4127 1821
rect 4133 1799 4147 1813
rect 4373 1833 4387 1847
rect 4213 1787 4227 1801
rect 4233 1779 4247 1793
rect 4253 1787 4267 1801
rect 4273 1779 4287 1793
rect 4293 1787 4307 1801
rect 4373 1799 4387 1813
rect 4393 1807 4407 1821
rect 4413 1799 4427 1813
rect 4533 1807 4547 1821
rect 4473 1787 4487 1801
rect 4493 1779 4507 1793
rect 4513 1787 4527 1801
rect 4633 1787 4647 1801
rect 4653 1799 4667 1813
rect 4333 1713 4347 1727
rect 4693 1787 4707 1801
rect 4773 1787 4787 1801
rect 4813 1787 4827 1801
rect 4893 1799 4907 1813
rect 4913 1807 4927 1821
rect 4793 1767 4807 1781
rect 4933 1799 4947 1813
rect 5013 1787 5027 1801
rect 5033 1779 5047 1793
rect 5053 1787 5067 1801
rect 5073 1779 5087 1793
rect 5093 1787 5107 1801
rect 5353 1833 5367 1847
rect 5173 1779 5187 1793
rect 5273 1787 5287 1801
rect 5313 1787 5327 1801
rect 5193 1767 5207 1781
rect 5293 1767 5307 1781
rect 5313 1733 5327 1747
rect 5433 1807 5447 1821
rect 5533 1807 5547 1821
rect 5373 1787 5387 1801
rect 5393 1779 5407 1793
rect 5413 1787 5427 1801
rect 5553 1787 5567 1801
rect 5573 1779 5587 1793
rect 5593 1787 5607 1801
rect 5653 1779 5667 1793
rect 5693 1779 5707 1793
rect 353 1587 367 1601
rect 373 1599 387 1613
rect 393 1587 407 1601
rect 73 1559 87 1573
rect 113 1559 127 1573
rect 133 1567 147 1581
rect 233 1567 247 1581
rect 413 1579 427 1593
rect 513 1579 527 1593
rect 533 1587 547 1601
rect 553 1599 567 1613
rect 573 1587 587 1601
rect 93 1539 107 1553
rect 253 1559 267 1573
rect 293 1559 307 1573
rect 273 1539 287 1553
rect 633 1567 647 1581
rect 753 1599 767 1613
rect 773 1587 787 1601
rect 653 1559 667 1573
rect 673 1567 687 1581
rect 893 1579 907 1593
rect 913 1587 927 1601
rect 933 1579 947 1593
rect 873 1559 887 1573
rect 1013 1567 1027 1581
rect 1033 1559 1047 1573
rect 1073 1559 1087 1573
rect 1153 1567 1167 1581
rect 1293 1599 1307 1613
rect 1173 1559 1187 1573
rect 1193 1567 1207 1581
rect 1273 1579 1287 1593
rect 1053 1539 1067 1553
rect 1313 1579 1327 1593
rect 1413 1579 1427 1593
rect 1453 1579 1467 1593
rect 1553 1587 1567 1601
rect 1573 1599 1587 1613
rect 1633 1579 1647 1593
rect 1653 1587 1667 1601
rect 1673 1579 1687 1593
rect 1693 1587 1707 1601
rect 1713 1579 1727 1593
rect 1773 1587 1787 1601
rect 1913 1636 1927 1650
rect 1933 1636 1947 1650
rect 1953 1636 1967 1650
rect 1985 1636 1999 1650
rect 2013 1636 2027 1650
rect 2073 1633 2087 1647
rect 2093 1633 2107 1647
rect 2113 1633 2127 1647
rect 1853 1559 1867 1573
rect 1985 1583 1999 1597
rect 2033 1599 2047 1613
rect 2013 1565 2027 1579
rect 2153 1559 2167 1573
rect 2193 1567 2207 1581
rect 1913 1531 1927 1545
rect 1953 1531 1967 1545
rect 1933 1507 1947 1521
rect 1912 1492 1926 1506
rect 2093 1535 2107 1549
rect 1986 1510 2000 1524
rect 2013 1510 2027 1524
rect 2073 1493 2087 1507
rect 2093 1493 2107 1507
rect 2113 1493 2127 1507
rect 2293 1579 2307 1593
rect 2313 1587 2327 1601
rect 2333 1579 2347 1593
rect 2353 1559 2367 1573
rect 2433 1567 2447 1581
rect 2453 1559 2467 1573
rect 2473 1567 2487 1581
rect 2593 1579 2607 1593
rect 2613 1587 2627 1601
rect 2633 1579 2647 1593
rect 2573 1559 2587 1573
rect 2713 1567 2727 1581
rect 2773 1593 2787 1607
rect 2833 1593 2847 1607
rect 2733 1559 2747 1573
rect 2753 1567 2767 1581
rect 2853 1579 2867 1593
rect 2873 1587 2887 1601
rect 3153 1633 3167 1647
rect 3173 1633 3187 1647
rect 3193 1633 3207 1647
rect 3253 1636 3267 1650
rect 3281 1636 3295 1650
rect 3313 1636 3327 1650
rect 3333 1636 3347 1650
rect 3353 1636 3367 1650
rect 2893 1579 2907 1593
rect 2993 1579 3007 1593
rect 3013 1587 3027 1601
rect 3033 1579 3047 1593
rect 2833 1559 2847 1573
rect 2973 1559 2987 1573
rect 3233 1599 3247 1613
rect 3073 1567 3087 1581
rect 3281 1583 3295 1597
rect 3113 1559 3127 1573
rect 3253 1565 3267 1579
rect 3413 1559 3427 1573
rect 3173 1535 3187 1549
rect 3313 1531 3327 1545
rect 3353 1531 3367 1545
rect 3253 1510 3267 1524
rect 3280 1510 3294 1524
rect 3153 1493 3167 1507
rect 3173 1493 3187 1507
rect 3193 1493 3207 1507
rect 3333 1507 3347 1521
rect 3354 1492 3368 1506
rect 3493 1587 3507 1601
rect 3593 1579 3607 1593
rect 3613 1587 3627 1601
rect 3633 1599 3647 1613
rect 3653 1587 3667 1601
rect 3713 1579 3727 1593
rect 3733 1587 3747 1601
rect 3753 1579 3767 1593
rect 3873 1579 3887 1593
rect 3773 1559 3787 1573
rect 3913 1579 3927 1593
rect 3993 1579 4007 1593
rect 4013 1567 4027 1581
rect 4053 1579 4067 1593
rect 4113 1567 4127 1581
rect 4133 1559 4147 1573
rect 4153 1567 4167 1581
rect 4253 1579 4267 1593
rect 4273 1587 4287 1601
rect 4293 1579 4307 1593
rect 4313 1587 4327 1601
rect 4333 1579 4347 1593
rect 4413 1579 4427 1593
rect 4433 1587 4447 1601
rect 4493 1613 4507 1627
rect 4453 1579 4467 1593
rect 4473 1587 4487 1601
rect 4493 1579 4507 1593
rect 4573 1579 4587 1593
rect 4593 1587 4607 1601
rect 4613 1579 4627 1593
rect 4633 1587 4647 1601
rect 4653 1579 4667 1593
rect 4553 1553 4567 1567
rect 4733 1567 4747 1581
rect 4753 1559 4767 1573
rect 4773 1567 4787 1581
rect 4853 1579 4867 1593
rect 4873 1587 4887 1601
rect 4893 1579 4907 1593
rect 5013 1579 5027 1593
rect 4913 1559 4927 1573
rect 5033 1567 5047 1581
rect 5213 1633 5227 1647
rect 5253 1633 5267 1647
rect 5073 1579 5087 1593
rect 5153 1593 5167 1607
rect 5153 1559 5167 1573
rect 5193 1559 5207 1573
rect 5213 1567 5227 1581
rect 5173 1539 5187 1553
rect 5153 1513 5167 1527
rect 5273 1613 5287 1627
rect 5293 1579 5307 1593
rect 5313 1587 5327 1601
rect 5333 1579 5347 1593
rect 5353 1587 5367 1601
rect 5373 1579 5387 1593
rect 5453 1567 5467 1581
rect 5473 1559 5487 1573
rect 5493 1567 5507 1581
rect 5253 1513 5267 1527
rect 5493 1533 5507 1547
rect 5533 1613 5547 1627
rect 5573 1559 5587 1573
rect 5613 1559 5627 1573
rect 5633 1567 5647 1581
rect 5753 1579 5767 1593
rect 5773 1587 5787 1601
rect 5593 1539 5607 1553
rect 2133 1444 2147 1447
rect 3233 1444 3247 1447
rect 113 1347 127 1361
rect 73 1319 87 1333
rect 93 1327 107 1341
rect 133 1327 147 1341
rect 393 1347 407 1361
rect 193 1299 207 1313
rect 213 1287 227 1301
rect 233 1299 247 1313
rect 253 1307 267 1321
rect 353 1319 367 1333
rect 373 1327 387 1341
rect 413 1327 427 1341
rect 493 1327 507 1341
rect 633 1327 647 1341
rect 513 1307 527 1321
rect 533 1299 547 1313
rect 553 1307 567 1321
rect 653 1307 667 1321
rect 673 1299 687 1313
rect 693 1307 707 1321
rect 793 1307 807 1321
rect 813 1319 827 1333
rect 853 1307 867 1321
rect 913 1319 927 1333
rect 933 1327 947 1341
rect 953 1319 967 1333
rect 1153 1347 1167 1361
rect 1133 1327 1147 1341
rect 1173 1327 1187 1341
rect 1193 1319 1207 1333
rect 1273 1319 1287 1333
rect 1293 1327 1307 1341
rect 1053 1299 1067 1313
rect 1073 1287 1087 1301
rect 1313 1319 1327 1333
rect 1413 1319 1427 1333
rect 1433 1327 1447 1341
rect 1453 1319 1467 1333
rect 1533 1319 1547 1333
rect 1553 1327 1567 1341
rect 1713 1347 1727 1361
rect 2133 1433 2147 1444
rect 1573 1319 1587 1333
rect 1673 1319 1687 1333
rect 1693 1327 1707 1341
rect 1733 1327 1747 1341
rect 1793 1319 1807 1333
rect 1813 1327 1827 1341
rect 1973 1347 1987 1361
rect 1833 1319 1847 1333
rect 1933 1319 1947 1333
rect 1953 1327 1967 1341
rect 1993 1327 2007 1341
rect 2233 1347 2247 1361
rect 2193 1319 2207 1333
rect 2213 1327 2227 1341
rect 2253 1327 2267 1341
rect 2373 1347 2387 1361
rect 2333 1319 2347 1333
rect 2353 1327 2367 1341
rect 2393 1327 2407 1341
rect 2073 1299 2087 1313
rect 2093 1287 2107 1301
rect 2853 1373 2867 1387
rect 2593 1327 2607 1341
rect 2453 1287 2467 1301
rect 2473 1299 2487 1313
rect 2613 1307 2627 1321
rect 2633 1299 2647 1313
rect 2653 1307 2667 1321
rect 2713 1299 2727 1313
rect 2733 1287 2747 1301
rect 2753 1299 2767 1313
rect 2773 1307 2787 1321
rect 2833 1273 2847 1287
rect 3233 1433 3247 1444
rect 2873 1327 2887 1341
rect 3013 1327 3027 1341
rect 3153 1327 3167 1341
rect 2893 1307 2907 1321
rect 2913 1299 2927 1313
rect 2933 1307 2947 1321
rect 3033 1307 3047 1321
rect 3053 1299 3067 1313
rect 3073 1307 3087 1321
rect 3173 1307 3187 1321
rect 3193 1299 3207 1313
rect 3213 1307 3227 1321
rect 3293 1299 3307 1313
rect 3313 1287 3327 1301
rect 3373 1287 3387 1301
rect 3393 1299 3407 1313
rect 3493 1307 3507 1321
rect 3653 1333 3667 1347
rect 3713 1333 3727 1347
rect 3813 1327 3827 1341
rect 3533 1307 3547 1321
rect 3633 1307 3647 1321
rect 3653 1299 3667 1313
rect 3673 1287 3687 1301
rect 3693 1299 3707 1313
rect 3753 1307 3767 1321
rect 3773 1299 3787 1313
rect 3793 1307 3807 1321
rect 4013 1327 4027 1341
rect 4153 1327 4167 1341
rect 4433 1327 4447 1341
rect 4633 1327 4647 1341
rect 3913 1299 3927 1313
rect 4033 1307 4047 1321
rect 3933 1287 3947 1301
rect 4053 1299 4067 1313
rect 4073 1307 4087 1321
rect 4173 1307 4187 1321
rect 4193 1299 4207 1313
rect 4213 1307 4227 1321
rect 4293 1307 4307 1321
rect 4313 1299 4327 1313
rect 4333 1287 4347 1301
rect 4353 1299 4367 1313
rect 4453 1307 4467 1321
rect 4473 1299 4487 1313
rect 4493 1307 4507 1321
rect 4573 1307 4587 1321
rect 4593 1299 4607 1313
rect 4613 1307 4627 1321
rect 4713 1319 4727 1333
rect 4733 1327 4747 1341
rect 4753 1319 4767 1333
rect 4893 1327 4907 1341
rect 4833 1307 4847 1321
rect 4853 1299 4867 1313
rect 4873 1307 4887 1321
rect 4973 1307 4987 1321
rect 5013 1307 5027 1321
rect 5093 1319 5107 1333
rect 5113 1327 5127 1341
rect 4993 1287 5007 1301
rect 5133 1319 5147 1333
rect 5233 1319 5247 1333
rect 5253 1327 5267 1341
rect 5273 1319 5287 1333
rect 5353 1327 5367 1341
rect 5533 1327 5547 1341
rect 5693 1327 5707 1341
rect 5373 1307 5387 1321
rect 5393 1299 5407 1313
rect 5413 1307 5427 1321
rect 5473 1307 5487 1321
rect 5493 1299 5507 1313
rect 5513 1307 5527 1321
rect 5633 1307 5647 1321
rect 5653 1299 5667 1313
rect 5673 1307 5687 1321
rect 73 1107 87 1121
rect 93 1119 107 1133
rect 153 1107 167 1121
rect 173 1119 187 1133
rect 193 1107 207 1121
rect 213 1099 227 1113
rect 293 1099 307 1113
rect 313 1107 327 1121
rect 333 1099 347 1113
rect 433 1099 447 1113
rect 453 1107 467 1121
rect 473 1099 487 1113
rect 353 1079 367 1093
rect 493 1079 507 1093
rect 593 1087 607 1101
rect 713 1099 727 1113
rect 733 1107 747 1121
rect 753 1099 767 1113
rect 873 1107 887 1121
rect 893 1119 907 1133
rect 913 1107 927 1121
rect 933 1099 947 1113
rect 1053 1099 1067 1113
rect 1073 1107 1087 1121
rect 1093 1099 1107 1113
rect 1173 1107 1187 1121
rect 1193 1119 1207 1133
rect 1253 1107 1267 1121
rect 1273 1119 1287 1133
rect 1293 1107 1307 1121
rect 613 1079 627 1093
rect 653 1079 667 1093
rect 633 1059 647 1073
rect 773 1079 787 1093
rect 1033 1079 1047 1093
rect 1113 1073 1127 1087
rect 1153 1073 1167 1087
rect 1313 1099 1327 1113
rect 1413 1107 1427 1121
rect 1433 1119 1447 1133
rect 1533 1119 1547 1133
rect 1633 1119 1647 1133
rect 1513 1099 1527 1113
rect 1553 1099 1567 1113
rect 1653 1107 1667 1121
rect 1813 1113 1827 1127
rect 1853 1113 1867 1127
rect 1753 1087 1767 1101
rect 1773 1079 1787 1093
rect 1813 1079 1827 1093
rect 1893 1087 1907 1101
rect 1913 1079 1927 1093
rect 1933 1087 1947 1101
rect 2033 1099 2047 1113
rect 2053 1107 2067 1121
rect 2073 1099 2087 1113
rect 2013 1079 2027 1093
rect 1793 1059 1807 1073
rect 2153 1087 2167 1101
rect 2173 1079 2187 1093
rect 2213 1079 2227 1093
rect 2293 1087 2307 1101
rect 2453 1099 2467 1113
rect 2473 1107 2487 1121
rect 2493 1099 2507 1113
rect 2713 1119 2727 1133
rect 2733 1107 2747 1121
rect 2833 1119 2847 1133
rect 2953 1119 2967 1133
rect 2193 1059 2207 1073
rect 2313 1079 2327 1093
rect 2353 1079 2367 1093
rect 2433 1079 2447 1093
rect 2333 1059 2347 1073
rect 2573 1087 2587 1101
rect 2593 1079 2607 1093
rect 2633 1079 2647 1093
rect 2613 1059 2627 1073
rect 2813 1099 2827 1113
rect 2853 1099 2867 1113
rect 2933 1099 2947 1113
rect 2973 1099 2987 1113
rect 3053 1099 3067 1113
rect 3233 1119 3247 1133
rect 3373 1119 3387 1133
rect 3093 1087 3107 1101
rect 3113 1099 3127 1113
rect 3213 1099 3227 1113
rect 3253 1099 3267 1113
rect 3353 1099 3367 1113
rect 3393 1099 3407 1113
rect 3473 1107 3487 1121
rect 3493 1119 3507 1133
rect 3593 1099 3607 1113
rect 3613 1107 3627 1121
rect 3793 1133 3807 1147
rect 3633 1099 3647 1113
rect 3733 1099 3747 1113
rect 3753 1107 3767 1121
rect 3773 1099 3787 1113
rect 3573 1079 3587 1093
rect 3713 1079 3727 1093
rect 3833 1087 3847 1101
rect 3853 1079 3867 1093
rect 3873 1087 3887 1101
rect 3953 1087 3967 1101
rect 4093 1119 4107 1133
rect 4193 1119 4207 1133
rect 3973 1079 3987 1093
rect 3993 1087 4007 1101
rect 4073 1099 4087 1113
rect 3793 1053 3807 1067
rect 4113 1099 4127 1113
rect 4213 1107 4227 1121
rect 4313 1099 4327 1113
rect 4333 1107 4347 1121
rect 4353 1119 4367 1133
rect 4373 1107 4387 1121
rect 4493 1099 4507 1113
rect 4513 1107 4527 1121
rect 4533 1099 4547 1113
rect 4613 1099 4627 1113
rect 4633 1107 4647 1121
rect 4653 1119 4667 1133
rect 4673 1107 4687 1121
rect 4733 1099 4747 1113
rect 4753 1107 4767 1121
rect 4773 1099 4787 1113
rect 4873 1099 4887 1113
rect 4473 1079 4487 1093
rect 4633 1073 4647 1087
rect 4713 1073 4727 1087
rect 4793 1079 4807 1093
rect 4993 1119 5007 1133
rect 4913 1099 4927 1113
rect 5013 1107 5027 1121
rect 5093 1119 5107 1133
rect 5113 1107 5127 1121
rect 5213 1087 5227 1101
rect 5233 1079 5247 1093
rect 5253 1087 5267 1101
rect 5373 1099 5387 1113
rect 5393 1107 5407 1121
rect 5493 1119 5507 1133
rect 5413 1099 5427 1113
rect 5473 1099 5487 1113
rect 5353 1079 5367 1093
rect 5513 1099 5527 1113
rect 5673 1113 5687 1127
rect 5613 1087 5627 1101
rect 5633 1079 5647 1093
rect 5673 1079 5687 1093
rect 5753 1107 5767 1121
rect 5773 1119 5787 1133
rect 5653 1059 5667 1073
rect 5693 1073 5707 1087
rect 113 867 127 881
rect 73 839 87 853
rect 93 847 107 861
rect 133 847 147 861
rect 393 867 407 881
rect 193 819 207 833
rect 213 807 227 821
rect 233 819 247 833
rect 253 827 267 841
rect 353 839 367 853
rect 373 847 387 861
rect 413 847 427 861
rect 673 867 687 881
rect 493 827 507 841
rect 633 839 647 853
rect 653 847 667 861
rect 693 847 707 861
rect 913 847 927 861
rect 1093 867 1107 881
rect 513 819 527 833
rect 533 807 547 821
rect 553 819 567 833
rect 753 819 767 833
rect 773 807 787 821
rect 793 819 807 833
rect 813 827 827 841
rect 933 827 947 841
rect 953 819 967 833
rect 973 827 987 841
rect 1053 839 1067 853
rect 1073 847 1087 861
rect 1113 847 1127 861
rect 1233 847 1247 861
rect 1373 867 1387 881
rect 1173 827 1187 841
rect 1193 819 1207 833
rect 1213 827 1227 841
rect 1333 839 1347 853
rect 1353 847 1367 861
rect 1393 847 1407 861
rect 1133 793 1147 807
rect 1173 793 1187 807
rect 1593 873 1607 887
rect 1653 873 1667 887
rect 1553 839 1567 853
rect 1573 847 1587 861
rect 1753 867 1767 881
rect 1453 807 1467 821
rect 1473 819 1487 833
rect 1593 839 1607 853
rect 1713 839 1727 853
rect 1733 847 1747 861
rect 1773 847 1787 861
rect 1893 867 1907 881
rect 1993 867 2007 881
rect 1853 839 1867 853
rect 1873 847 1887 861
rect 1913 847 1927 861
rect 1973 847 1987 861
rect 2013 847 2027 861
rect 2033 839 2047 853
rect 2173 847 2187 861
rect 2113 827 2127 841
rect 2133 819 2147 833
rect 2153 827 2167 841
rect 2253 827 2267 841
rect 2293 839 2307 853
rect 2313 827 2327 841
rect 2513 839 2527 853
rect 2533 847 2547 861
rect 2393 807 2407 821
rect 2413 819 2427 833
rect 2553 839 2567 853
rect 2633 819 2647 833
rect 2673 827 2687 841
rect 2753 839 2767 853
rect 2773 847 2787 861
rect 2693 807 2707 821
rect 2793 839 2807 853
rect 2893 839 2907 853
rect 2913 847 2927 861
rect 2933 839 2947 853
rect 3253 839 3267 853
rect 3273 847 3287 861
rect 3013 807 3027 821
rect 3033 819 3047 833
rect 3133 819 3147 833
rect 3153 807 3167 821
rect 3293 839 3307 853
rect 3393 827 3407 841
rect 3433 827 3447 841
rect 3513 827 3527 841
rect 3553 827 3567 841
rect 3633 827 3647 841
rect 3413 807 3427 821
rect 3533 807 3547 821
rect 3653 819 3667 833
rect 3673 807 3687 821
rect 3693 819 3707 833
rect 3773 819 3787 833
rect 3793 807 3807 821
rect 3793 773 3807 787
rect 3853 873 3867 887
rect 3873 847 3887 861
rect 3893 827 3907 841
rect 3913 819 3927 833
rect 3933 827 3947 841
rect 3993 839 4007 853
rect 4013 847 4027 861
rect 4033 839 4047 853
rect 4133 847 4147 861
rect 4273 847 4287 861
rect 4153 827 4167 841
rect 4173 819 4187 833
rect 4193 827 4207 841
rect 4293 827 4307 841
rect 4313 819 4327 833
rect 4333 827 4347 841
rect 4533 847 4547 861
rect 4413 807 4427 821
rect 4433 819 4447 833
rect 4553 827 4567 841
rect 4573 819 4587 833
rect 4593 827 4607 841
rect 4653 819 4667 833
rect 4673 807 4687 821
rect 4693 819 4707 833
rect 4713 827 4727 841
rect 4813 827 4827 841
rect 4933 847 4947 861
rect 5033 853 5047 867
rect 5093 853 5107 867
rect 4853 827 4867 841
rect 4953 827 4967 841
rect 4973 819 4987 833
rect 4993 827 5007 841
rect 5053 819 5067 833
rect 5073 807 5087 821
rect 5093 819 5107 833
rect 5113 827 5127 841
rect 5213 819 5227 833
rect 5253 827 5267 841
rect 5693 847 5707 861
rect 5273 807 5287 821
rect 5373 819 5387 833
rect 5473 827 5487 841
rect 5393 807 5407 821
rect 5493 819 5507 833
rect 5513 827 5527 841
rect 5533 819 5547 833
rect 5553 827 5567 841
rect 5633 827 5647 841
rect 5653 819 5667 833
rect 5673 827 5687 841
rect 73 607 87 621
rect 233 619 247 633
rect 253 627 267 641
rect 273 639 287 653
rect 293 627 307 641
rect 93 599 107 613
rect 133 599 147 613
rect 113 579 127 593
rect 373 607 387 621
rect 533 619 547 633
rect 553 627 567 641
rect 573 619 587 633
rect 633 627 647 641
rect 653 639 667 653
rect 673 627 687 641
rect 693 619 707 633
rect 393 599 407 613
rect 433 599 447 613
rect 513 599 527 613
rect 413 579 427 593
rect 773 607 787 621
rect 793 599 807 613
rect 813 607 827 621
rect 953 619 967 633
rect 973 627 987 641
rect 993 619 1007 633
rect 1193 627 1207 641
rect 1213 639 1227 653
rect 1233 627 1247 641
rect 933 599 947 613
rect 1073 607 1087 621
rect 1253 619 1267 633
rect 1353 619 1367 633
rect 1373 627 1387 641
rect 1393 639 1407 653
rect 1413 627 1427 641
rect 1093 599 1107 613
rect 1133 599 1147 613
rect 1113 579 1127 593
rect 1493 599 1507 613
rect 1533 599 1547 613
rect 1553 607 1567 621
rect 1673 619 1687 633
rect 1693 627 1707 641
rect 1713 619 1727 633
rect 1913 627 1927 641
rect 1933 639 1947 653
rect 1953 627 1967 641
rect 2093 639 2107 653
rect 1513 579 1527 593
rect 1653 599 1667 613
rect 1793 607 1807 621
rect 1973 619 1987 633
rect 2073 619 2087 633
rect 1813 599 1827 613
rect 1853 599 1867 613
rect 1833 579 1847 593
rect 2113 619 2127 633
rect 2193 627 2207 641
rect 2253 639 2267 653
rect 2233 619 2247 633
rect 2313 619 2327 633
rect 2353 607 2367 621
rect 2373 619 2387 633
rect 2453 607 2467 621
rect 2473 599 2487 613
rect 2493 607 2507 621
rect 2593 607 2607 621
rect 2733 639 2747 653
rect 2613 599 2627 613
rect 2633 607 2647 621
rect 2713 619 2727 633
rect 2753 619 2767 633
rect 2813 619 2827 633
rect 2833 627 2847 641
rect 2853 619 2867 633
rect 2873 599 2887 613
rect 2973 607 2987 621
rect 3073 627 3087 641
rect 3093 639 3107 653
rect 3113 627 3127 641
rect 2993 599 3007 613
rect 3013 607 3027 621
rect 3133 619 3147 633
rect 3273 633 3287 647
rect 3313 633 3327 647
rect 3233 607 3247 621
rect 3253 599 3267 613
rect 3293 599 3307 613
rect 3353 607 3367 621
rect 3373 599 3387 613
rect 3393 607 3407 621
rect 3513 619 3527 633
rect 3533 627 3547 641
rect 3553 619 3567 633
rect 3493 599 3507 613
rect 3273 579 3287 593
rect 3613 607 3627 621
rect 3693 633 3707 647
rect 3733 633 3747 647
rect 3633 599 3647 613
rect 3653 607 3667 621
rect 3773 619 3787 633
rect 3793 627 3807 641
rect 3813 619 3827 633
rect 3873 653 3887 667
rect 3753 599 3767 613
rect 3853 613 3867 627
rect 3873 619 3887 633
rect 3893 627 3907 641
rect 3913 619 3927 633
rect 4013 627 4027 641
rect 4033 639 4047 653
rect 4053 627 4067 641
rect 4073 619 4087 633
rect 4173 619 4187 633
rect 4193 627 4207 641
rect 4213 619 4227 633
rect 4333 627 4347 641
rect 4353 639 4367 653
rect 3933 599 3947 613
rect 4233 599 4247 613
rect 4433 619 4447 633
rect 4453 627 4467 641
rect 4473 639 4487 653
rect 4493 627 4507 641
rect 4593 619 4607 633
rect 4613 627 4627 641
rect 4633 619 4647 633
rect 4733 619 4747 633
rect 4753 627 4767 641
rect 4773 619 4787 633
rect 4853 619 4867 633
rect 4873 627 4887 641
rect 4993 639 5007 653
rect 4893 619 4907 633
rect 5013 627 5027 641
rect 4573 599 4587 613
rect 4713 599 4727 613
rect 4913 599 4927 613
rect 5113 619 5127 633
rect 5153 619 5167 633
rect 5273 619 5287 633
rect 5293 627 5307 641
rect 5313 619 5327 633
rect 5373 619 5387 633
rect 5393 627 5407 641
rect 5413 619 5427 633
rect 5553 619 5567 633
rect 5573 627 5587 641
rect 5673 639 5687 653
rect 5593 619 5607 633
rect 5653 619 5667 633
rect 5253 599 5267 613
rect 5433 599 5447 613
rect 5533 599 5547 613
rect 5693 619 5707 633
rect 113 387 127 401
rect 73 359 87 373
rect 93 367 107 381
rect 133 367 147 381
rect 213 367 227 381
rect 373 367 387 381
rect 553 387 567 401
rect 233 347 247 361
rect 253 339 267 353
rect 273 347 287 361
rect 393 347 407 361
rect 413 339 427 353
rect 433 347 447 361
rect 513 359 527 373
rect 533 367 547 381
rect 573 367 587 381
rect 653 347 667 361
rect 673 359 687 373
rect 833 387 847 401
rect 713 347 727 361
rect 793 359 807 373
rect 813 367 827 381
rect 853 367 867 381
rect 1073 387 1087 401
rect 1053 367 1067 381
rect 1093 367 1107 381
rect 933 347 947 361
rect 1113 359 1127 373
rect 953 339 967 353
rect 973 327 987 341
rect 993 339 1007 353
rect 1213 339 1227 353
rect 1393 387 1407 401
rect 1253 347 1267 361
rect 1353 359 1367 373
rect 1373 367 1387 381
rect 1413 367 1427 381
rect 1273 327 1287 341
rect 1613 367 1627 381
rect 1413 333 1427 347
rect 1473 333 1487 347
rect 1513 339 1527 353
rect 1633 347 1647 361
rect 1533 327 1547 341
rect 1653 339 1667 353
rect 1673 347 1687 361
rect 1753 347 1767 361
rect 1773 359 1787 373
rect 1813 347 1827 361
rect 1873 347 1887 361
rect 1913 347 1927 361
rect 2133 367 2147 381
rect 1893 327 1907 341
rect 2013 327 2027 341
rect 2033 339 2047 353
rect 2153 347 2167 361
rect 2173 339 2187 353
rect 2193 347 2207 361
rect 2273 347 2287 361
rect 2553 387 2567 401
rect 2513 359 2527 373
rect 2533 367 2547 381
rect 2573 367 2587 381
rect 2693 367 2707 381
rect 2293 339 2307 353
rect 2313 327 2327 341
rect 2333 339 2347 353
rect 2413 339 2427 353
rect 2433 327 2447 341
rect 2633 347 2647 361
rect 2653 339 2667 353
rect 2673 347 2687 361
rect 2793 339 2807 353
rect 2893 347 2907 361
rect 2933 347 2947 361
rect 3153 373 3167 387
rect 3293 373 3307 387
rect 2813 327 2827 341
rect 2913 327 2927 341
rect 2993 327 3007 341
rect 3013 339 3027 353
rect 3113 347 3127 361
rect 3133 339 3147 353
rect 3153 327 3167 341
rect 3173 339 3187 353
rect 3253 339 3267 353
rect 3273 327 3287 341
rect 3293 339 3307 353
rect 3313 347 3327 361
rect 3573 367 3587 381
rect 3853 387 3867 401
rect 3413 339 3427 353
rect 3513 347 3527 361
rect 3433 327 3447 341
rect 3533 339 3547 353
rect 3553 347 3567 361
rect 3653 339 3667 353
rect 3673 327 3687 341
rect 3693 339 3707 353
rect 3713 347 3727 361
rect 3813 359 3827 373
rect 3833 367 3847 381
rect 3873 367 3887 381
rect 3933 359 3947 373
rect 3953 367 3967 381
rect 4133 387 4147 401
rect 3973 359 3987 373
rect 4093 359 4107 373
rect 4113 367 4127 381
rect 4153 367 4167 381
rect 4233 367 4247 381
rect 4253 347 4267 361
rect 4273 339 4287 353
rect 4293 347 4307 361
rect 4473 359 4487 373
rect 4493 367 4507 381
rect 4373 339 4387 353
rect 4393 327 4407 341
rect 4513 359 4527 373
rect 4593 367 4607 381
rect 4613 347 4627 361
rect 4633 339 4647 353
rect 4653 347 4667 361
rect 4833 367 4847 381
rect 4733 339 4747 353
rect 4853 347 4867 361
rect 4753 327 4767 341
rect 4873 339 4887 353
rect 4893 347 4907 361
rect 4953 339 4967 353
rect 4973 347 4987 361
rect 5133 367 5147 381
rect 5333 367 5347 381
rect 5633 367 5647 381
rect 5013 339 5027 353
rect 5033 347 5047 361
rect 5153 347 5167 361
rect 5173 339 5187 353
rect 5193 347 5207 361
rect 5273 347 5287 361
rect 5293 339 5307 353
rect 5313 347 5327 361
rect 5453 347 5467 361
rect 5473 339 5487 353
rect 5493 327 5507 341
rect 5513 339 5527 353
rect 5573 347 5587 361
rect 5593 339 5607 353
rect 5613 347 5627 361
rect 5713 359 5727 373
rect 5733 367 5747 381
rect 5753 359 5767 373
rect 193 147 207 161
rect 213 159 227 173
rect 233 147 247 161
rect 73 127 87 141
rect 253 139 267 153
rect 373 139 387 153
rect 393 147 407 161
rect 413 159 427 173
rect 433 147 447 161
rect 533 139 547 153
rect 553 147 567 161
rect 573 139 587 153
rect 633 139 647 153
rect 653 147 667 161
rect 673 139 687 153
rect 913 159 927 173
rect 933 147 947 161
rect 93 119 107 133
rect 133 119 147 133
rect 113 99 127 113
rect 513 119 527 133
rect 693 119 707 133
rect 793 127 807 141
rect 813 119 827 133
rect 853 119 867 133
rect 833 99 847 113
rect 1013 139 1027 153
rect 1033 147 1047 161
rect 1053 139 1067 153
rect 1153 147 1167 161
rect 1173 159 1187 173
rect 1193 147 1207 161
rect 1313 159 1327 173
rect 1213 139 1227 153
rect 1293 139 1307 153
rect 1073 119 1087 133
rect 1333 139 1347 153
rect 1413 139 1427 153
rect 1453 127 1467 141
rect 1473 139 1487 153
rect 1573 147 1587 161
rect 1593 159 1607 173
rect 1693 139 1707 153
rect 1713 147 1727 161
rect 1733 139 1747 153
rect 1673 119 1687 133
rect 1813 127 1827 141
rect 1833 119 1847 133
rect 1853 127 1867 141
rect 1913 119 1927 133
rect 1953 119 1967 133
rect 1973 127 1987 141
rect 2093 127 2107 141
rect 2213 139 2227 153
rect 1933 99 1947 113
rect 2113 119 2127 133
rect 2153 119 2167 133
rect 2253 139 2267 153
rect 2133 99 2147 113
rect 2353 127 2367 141
rect 2373 119 2387 133
rect 2393 127 2407 141
rect 2453 139 2467 153
rect 2493 127 2507 141
rect 2513 139 2527 153
rect 2613 139 2627 153
rect 2633 147 2647 161
rect 2653 159 2667 173
rect 2673 147 2687 161
rect 2753 139 2767 153
rect 2773 127 2787 141
rect 2813 139 2827 153
rect 2893 127 2907 141
rect 2913 119 2927 133
rect 2933 127 2947 141
rect 3033 127 3047 141
rect 3293 147 3307 161
rect 3313 159 3327 173
rect 3053 119 3067 133
rect 3073 127 3087 141
rect 3153 127 3167 141
rect 2973 93 2987 107
rect 3033 93 3047 107
rect 3173 119 3187 133
rect 3213 119 3227 133
rect 3193 99 3207 113
rect 3373 139 3387 153
rect 3393 147 3407 161
rect 3413 139 3427 153
rect 3533 147 3547 161
rect 3553 159 3567 173
rect 3433 119 3447 133
rect 3633 127 3647 141
rect 3653 119 3667 133
rect 3673 127 3687 141
rect 3753 139 3767 153
rect 3793 139 3807 153
rect 3853 139 3867 153
rect 3893 139 3907 153
rect 3993 127 4007 141
rect 4013 119 4027 133
rect 4033 127 4047 141
rect 4113 139 4127 153
rect 4313 159 4327 173
rect 4153 127 4167 141
rect 4173 139 4187 153
rect 4293 139 4307 153
rect 4333 139 4347 153
rect 4393 127 4407 141
rect 4573 153 4587 167
rect 4613 153 4627 167
rect 4413 119 4427 133
rect 4433 127 4447 141
rect 4533 127 4547 141
rect 4713 139 4727 153
rect 4733 147 4747 161
rect 4753 139 4767 153
rect 4553 119 4567 133
rect 4593 119 4607 133
rect 4693 119 4707 133
rect 4573 99 4587 113
rect 4813 127 4827 141
rect 4833 119 4847 133
rect 4853 127 4867 141
rect 4973 139 4987 153
rect 4993 147 5007 161
rect 5093 159 5107 173
rect 5013 139 5027 153
rect 5073 139 5087 153
rect 4953 119 4967 133
rect 5113 139 5127 153
rect 5213 127 5227 141
rect 5313 147 5327 161
rect 5233 119 5247 133
rect 5253 127 5267 141
rect 5333 139 5347 153
rect 5373 147 5387 161
rect 5473 159 5487 173
rect 5393 139 5407 153
rect 5493 147 5507 161
rect 5593 147 5607 161
rect 5613 159 5627 173
rect 5673 127 5687 141
rect 5693 119 5707 133
rect 5713 127 5727 141
<< metal2 >>
rect 4177 5678 4185 5702
rect 73 5633 87 5647
rect 76 5467 83 5633
rect 93 5613 107 5627
rect 253 5633 267 5647
rect 233 5613 247 5627
rect 96 5487 103 5613
rect 136 5447 143 5453
rect 73 5423 87 5427
rect 56 5416 87 5423
rect 56 5387 63 5416
rect 73 5413 87 5416
rect 133 5433 147 5447
rect 196 5427 203 5613
rect 236 5443 243 5613
rect 256 5547 263 5633
rect 433 5643 447 5647
rect 456 5643 463 5653
rect 433 5636 463 5643
rect 433 5633 447 5636
rect 236 5436 263 5443
rect 256 5427 263 5436
rect 36 4787 43 5013
rect 36 4187 43 4673
rect 56 4507 63 5313
rect 76 5187 83 5373
rect 96 5327 103 5393
rect 156 5187 163 5213
rect 73 5173 87 5187
rect 113 5173 127 5187
rect 116 5167 123 5173
rect 133 5153 147 5167
rect 116 4983 123 5153
rect 136 5127 143 5153
rect 96 4976 123 4983
rect 76 4947 83 4973
rect 96 4967 103 4976
rect 93 4953 107 4967
rect 133 4963 147 4967
rect 73 4933 87 4947
rect 113 4933 127 4947
rect 133 4956 163 4963
rect 133 4953 147 4956
rect 116 4887 123 4933
rect 96 4687 103 4753
rect 116 4707 123 4773
rect 136 4687 143 4833
rect 156 4767 163 4956
rect 176 4803 183 5233
rect 196 5187 203 5413
rect 233 5393 247 5407
rect 253 5413 267 5427
rect 276 5407 283 5433
rect 396 5427 403 5473
rect 293 5423 307 5427
rect 293 5416 323 5423
rect 293 5413 307 5416
rect 273 5393 287 5407
rect 236 5247 243 5393
rect 236 5167 243 5213
rect 316 5187 323 5416
rect 373 5393 387 5407
rect 393 5413 407 5427
rect 233 5153 247 5167
rect 253 5143 267 5147
rect 276 5143 283 5173
rect 253 5136 283 5143
rect 253 5133 267 5136
rect 316 5123 323 5173
rect 356 5167 363 5393
rect 333 5123 347 5127
rect 316 5116 347 5123
rect 333 5113 347 5116
rect 216 4967 223 5113
rect 376 5027 383 5393
rect 456 5367 463 5636
rect 553 5663 567 5667
rect 793 5663 807 5667
rect 493 5633 507 5647
rect 553 5656 583 5663
rect 553 5653 567 5656
rect 496 5607 503 5633
rect 536 5607 543 5633
rect 496 5443 503 5593
rect 576 5487 583 5656
rect 776 5656 807 5663
rect 653 5633 667 5647
rect 656 5567 663 5633
rect 673 5613 687 5627
rect 713 5613 727 5627
rect 476 5436 503 5443
rect 376 4947 383 4973
rect 396 4967 403 5333
rect 416 5147 423 5353
rect 476 5347 483 5436
rect 536 5427 543 5473
rect 576 5427 583 5453
rect 496 5367 503 5413
rect 533 5413 547 5427
rect 573 5413 587 5427
rect 196 4847 203 4933
rect 273 4943 287 4947
rect 273 4936 293 4943
rect 273 4933 287 4936
rect 296 4907 303 4933
rect 373 4933 387 4947
rect 176 4796 203 4803
rect 73 4653 87 4667
rect 93 4673 107 4687
rect 133 4673 147 4687
rect 76 4483 83 4653
rect 96 4487 103 4493
rect 136 4487 143 4573
rect 156 4527 163 4713
rect 56 4476 83 4483
rect 56 4127 63 4476
rect 93 4473 107 4487
rect 133 4473 147 4487
rect 156 4423 163 4493
rect 176 4447 183 4773
rect 196 4727 203 4796
rect 216 4707 223 4893
rect 213 4703 227 4707
rect 196 4696 227 4703
rect 196 4647 203 4696
rect 213 4693 227 4696
rect 253 4693 267 4707
rect 236 4647 243 4673
rect 256 4627 263 4693
rect 156 4416 183 4423
rect 56 3983 63 4093
rect 76 4027 83 4413
rect 93 4193 107 4207
rect 96 4107 103 4193
rect 176 4187 183 4416
rect 153 4173 167 4187
rect 73 3983 87 3987
rect 56 3976 87 3983
rect 73 3973 87 3976
rect 96 3947 103 3973
rect 16 3027 23 3133
rect 16 1507 23 1553
rect 36 1147 43 1573
rect 36 607 43 1133
rect 56 627 63 3773
rect 96 3763 103 3913
rect 116 3787 123 4113
rect 136 3967 143 4153
rect 156 4087 163 4173
rect 156 4027 163 4033
rect 176 4027 183 4153
rect 196 4047 203 4513
rect 236 4467 243 4553
rect 233 4453 247 4467
rect 256 4447 263 4493
rect 276 4487 283 4653
rect 296 4487 303 4873
rect 316 4787 323 4913
rect 416 4783 423 4973
rect 396 4776 423 4783
rect 376 4687 383 4713
rect 396 4707 403 4776
rect 333 4683 347 4687
rect 316 4676 347 4683
rect 316 4647 323 4676
rect 333 4673 347 4676
rect 393 4663 407 4667
rect 416 4663 423 4753
rect 393 4656 423 4663
rect 393 4653 407 4656
rect 356 4627 363 4633
rect 233 4193 247 4207
rect 216 4147 223 4193
rect 236 4167 243 4193
rect 293 4173 307 4187
rect 176 4007 183 4013
rect 173 3993 187 4007
rect 76 3756 103 3763
rect 76 3747 83 3756
rect 116 3747 123 3753
rect 93 3713 107 3727
rect 113 3733 127 3747
rect 76 3527 83 3693
rect 96 3607 103 3713
rect 136 3707 143 3933
rect 96 3527 103 3573
rect 136 3527 143 3553
rect 93 3513 107 3527
rect 87 3436 93 3443
rect 76 3247 83 3253
rect 96 3247 103 3253
rect 73 3233 87 3247
rect 116 3187 123 3433
rect 136 3227 143 3453
rect 76 2987 83 3173
rect 96 3047 103 3173
rect 156 3063 163 3993
rect 236 3987 243 4113
rect 256 3987 263 4133
rect 296 4087 303 4173
rect 296 4047 303 4073
rect 233 3973 247 3987
rect 176 3467 183 3953
rect 316 3747 323 4473
rect 416 4467 423 4553
rect 336 4447 343 4453
rect 336 4187 343 4413
rect 356 4027 363 4053
rect 353 4013 367 4027
rect 213 3713 227 3727
rect 253 3713 267 3727
rect 216 3707 223 3713
rect 256 3707 263 3713
rect 216 3547 223 3593
rect 296 3587 303 3713
rect 276 3507 283 3573
rect 193 3213 207 3227
rect 136 3056 163 3063
rect 93 3033 107 3047
rect 76 2787 83 2793
rect 116 2787 123 2973
rect 73 2773 87 2787
rect 96 2587 103 2733
rect 93 2573 107 2587
rect 73 2533 87 2547
rect 76 2307 83 2533
rect 116 2527 123 2733
rect 76 1827 83 2113
rect 96 2087 103 2273
rect 113 2253 127 2267
rect 116 2167 123 2253
rect 136 2103 143 3056
rect 176 3003 183 3213
rect 156 2996 183 3003
rect 156 2747 163 2996
rect 196 2767 203 3213
rect 256 3207 263 3273
rect 276 3227 283 3253
rect 233 3023 247 3027
rect 216 3016 247 3023
rect 216 3007 223 3016
rect 233 3013 247 3016
rect 256 3007 263 3033
rect 276 3027 283 3213
rect 296 3047 303 3513
rect 316 3287 323 3733
rect 353 3723 367 3727
rect 336 3716 367 3723
rect 336 3707 343 3716
rect 353 3713 367 3716
rect 376 3703 383 4253
rect 396 4227 403 4433
rect 436 4267 443 5153
rect 496 5107 503 5173
rect 513 5163 527 5167
rect 536 5163 543 5193
rect 513 5156 543 5163
rect 513 5153 527 5156
rect 516 4967 523 5133
rect 536 5127 543 5156
rect 596 5163 603 5413
rect 616 5227 623 5433
rect 656 5427 663 5533
rect 676 5427 683 5613
rect 716 5587 723 5613
rect 696 5427 703 5473
rect 736 5427 743 5633
rect 776 5627 783 5656
rect 793 5653 807 5656
rect 813 5633 827 5647
rect 1373 5663 1387 5667
rect 1373 5656 1403 5663
rect 1373 5653 1387 5656
rect 776 5467 783 5613
rect 816 5567 823 5633
rect 896 5587 903 5633
rect 913 5613 927 5627
rect 973 5643 987 5647
rect 973 5636 1003 5643
rect 973 5633 987 5636
rect 916 5607 923 5613
rect 996 5607 1003 5636
rect 1053 5613 1067 5627
rect 953 5593 967 5607
rect 796 5447 803 5553
rect 956 5447 963 5593
rect 1056 5547 1063 5613
rect 1093 5613 1107 5627
rect 1096 5603 1103 5613
rect 1096 5596 1123 5603
rect 793 5433 807 5447
rect 653 5413 667 5427
rect 693 5413 707 5427
rect 713 5393 727 5407
rect 716 5367 723 5393
rect 616 5167 623 5173
rect 796 5167 803 5173
rect 587 5156 603 5163
rect 613 5153 627 5167
rect 633 5133 647 5147
rect 793 5153 807 5167
rect 636 4967 643 5133
rect 816 5147 823 5413
rect 916 5187 923 5413
rect 956 5407 963 5433
rect 1076 5427 1083 5593
rect 1116 5587 1123 5596
rect 1096 5447 1103 5573
rect 1093 5433 1107 5447
rect 953 5393 967 5407
rect 1113 5413 1127 5427
rect 1116 5407 1123 5413
rect 993 5393 1007 5407
rect 996 5207 1003 5393
rect 873 5173 887 5187
rect 876 5167 883 5173
rect 853 5153 867 5167
rect 913 5173 927 5187
rect 1033 5153 1047 5167
rect 856 5147 863 5153
rect 856 5127 863 5133
rect 473 4963 487 4967
rect 456 4956 487 4963
rect 456 4767 463 4956
rect 473 4953 487 4956
rect 493 4933 507 4947
rect 513 4953 527 4967
rect 533 4943 547 4947
rect 533 4936 553 4943
rect 533 4933 547 4936
rect 496 4887 503 4933
rect 556 4847 563 4933
rect 473 4703 487 4707
rect 456 4696 487 4703
rect 456 4667 463 4696
rect 473 4693 487 4696
rect 456 4447 463 4633
rect 496 4587 503 4673
rect 393 4213 407 4227
rect 433 4213 447 4227
rect 413 4193 427 4207
rect 416 4127 423 4193
rect 436 4107 443 4213
rect 496 4147 503 4533
rect 516 4467 523 4593
rect 536 4487 543 4653
rect 576 4547 583 4953
rect 633 4913 647 4927
rect 636 4907 643 4913
rect 576 4487 583 4513
rect 596 4487 603 4893
rect 653 4693 667 4707
rect 656 4687 663 4693
rect 633 4673 647 4687
rect 673 4673 687 4687
rect 636 4547 643 4673
rect 533 4473 547 4487
rect 513 4453 527 4467
rect 573 4473 587 4487
rect 656 4467 663 4533
rect 676 4507 683 4673
rect 696 4567 703 4953
rect 716 4487 723 4513
rect 653 4453 667 4467
rect 536 4227 543 4433
rect 533 4213 547 4227
rect 573 4213 587 4227
rect 553 4193 567 4207
rect 416 3983 423 4053
rect 456 4027 463 4093
rect 453 4013 467 4027
rect 493 4003 507 4007
rect 433 3983 447 3987
rect 416 3976 447 3983
rect 433 3973 447 3976
rect 493 3996 523 4003
rect 493 3993 507 3996
rect 393 3703 407 3707
rect 376 3696 407 3703
rect 393 3693 407 3696
rect 336 3547 343 3693
rect 376 3547 383 3553
rect 333 3533 347 3547
rect 353 3503 367 3507
rect 376 3503 383 3533
rect 396 3507 403 3693
rect 353 3496 383 3503
rect 353 3493 367 3496
rect 416 3307 423 3573
rect 436 3527 443 3693
rect 496 3567 503 3713
rect 433 3513 447 3527
rect 496 3507 503 3553
rect 493 3493 507 3507
rect 516 3463 523 3996
rect 536 3707 543 4133
rect 556 4127 563 4193
rect 576 4167 583 4213
rect 736 4207 743 5093
rect 756 4947 763 5093
rect 753 4933 767 4947
rect 776 4707 783 4913
rect 773 4693 787 4707
rect 813 4693 827 4707
rect 816 4507 823 4693
rect 833 4673 847 4687
rect 836 4607 843 4673
rect 876 4667 883 5153
rect 896 4967 903 5113
rect 916 4967 923 5133
rect 1036 5107 1043 5153
rect 1056 4983 1063 5173
rect 1116 5087 1123 5393
rect 1156 5387 1163 5413
rect 1176 5407 1183 5453
rect 1213 5423 1227 5427
rect 1196 5416 1227 5423
rect 1196 5407 1203 5416
rect 1213 5413 1227 5416
rect 1273 5403 1287 5407
rect 1296 5403 1303 5433
rect 1273 5396 1303 5403
rect 1273 5393 1287 5396
rect 1176 5383 1183 5393
rect 1176 5376 1203 5383
rect 1167 5156 1183 5163
rect 1073 4983 1087 4987
rect 1056 4976 1087 4983
rect 1073 4973 1087 4976
rect 956 4967 963 4973
rect 913 4953 927 4967
rect 896 4947 903 4953
rect 893 4933 907 4947
rect 953 4953 967 4967
rect 996 4947 1003 4973
rect 1033 4963 1047 4967
rect 1016 4956 1047 4963
rect 1016 4727 1023 4956
rect 1033 4953 1047 4956
rect 1093 4943 1107 4947
rect 1116 4943 1123 4953
rect 1093 4936 1123 4943
rect 1093 4933 1107 4936
rect 913 4683 927 4687
rect 913 4676 943 4683
rect 913 4673 927 4676
rect 893 4633 907 4647
rect 896 4607 903 4633
rect 936 4547 943 4676
rect 1056 4647 1063 4933
rect 993 4633 1007 4647
rect 996 4567 1003 4633
rect 856 4463 863 4533
rect 896 4507 903 4513
rect 873 4463 887 4467
rect 856 4456 887 4463
rect 873 4453 887 4456
rect 996 4467 1003 4553
rect 1053 4503 1067 4507
rect 1053 4496 1083 4503
rect 1053 4493 1067 4496
rect 673 4203 687 4207
rect 656 4196 687 4203
rect 576 4147 583 4153
rect 596 4067 603 4193
rect 656 4127 663 4196
rect 673 4193 687 4196
rect 713 4173 727 4187
rect 556 3987 563 4033
rect 616 4027 623 4033
rect 613 4013 627 4027
rect 636 4007 643 4093
rect 716 4007 723 4173
rect 733 4153 747 4167
rect 736 4107 743 4153
rect 756 4027 763 4193
rect 873 4173 887 4187
rect 753 4013 767 4027
rect 633 3993 647 4007
rect 716 3967 723 3993
rect 816 4007 823 4153
rect 876 4047 883 4173
rect 813 3993 827 4007
rect 876 3987 883 4033
rect 873 3973 887 3987
rect 693 3743 707 3747
rect 676 3736 707 3743
rect 553 3713 567 3727
rect 556 3707 563 3713
rect 573 3693 587 3707
rect 613 3693 627 3707
rect 576 3667 583 3693
rect 616 3687 623 3693
rect 573 3503 587 3507
rect 556 3496 587 3503
rect 556 3487 563 3496
rect 573 3493 587 3496
rect 596 3487 603 3513
rect 616 3507 623 3533
rect 613 3493 627 3507
rect 593 3473 607 3487
rect 633 3473 647 3487
rect 496 3456 523 3463
rect 316 3247 323 3253
rect 333 3203 347 3207
rect 356 3203 363 3293
rect 396 3267 403 3273
rect 393 3253 407 3267
rect 433 3263 447 3267
rect 433 3256 463 3263
rect 433 3253 447 3256
rect 456 3227 463 3256
rect 333 3196 363 3203
rect 333 3193 347 3196
rect 356 3067 363 3196
rect 396 3087 403 3213
rect 396 3027 403 3073
rect 273 3013 287 3027
rect 293 3003 307 3007
rect 316 3003 323 3013
rect 293 2996 323 3003
rect 293 2993 307 2996
rect 373 2993 387 3007
rect 393 3013 407 3027
rect 216 2987 223 2993
rect 376 2987 383 2993
rect 173 2733 187 2747
rect 193 2753 207 2767
rect 233 2753 247 2767
rect 176 2667 183 2733
rect 156 2587 163 2593
rect 153 2573 167 2587
rect 156 2267 163 2433
rect 136 2096 163 2103
rect 93 2073 107 2087
rect 133 2083 147 2087
rect 116 2076 147 2083
rect 116 2007 123 2076
rect 133 2073 147 2076
rect 73 1813 87 1827
rect 116 1767 123 1813
rect 133 1793 147 1807
rect 136 1787 143 1793
rect 136 1707 143 1773
rect 76 1587 83 1633
rect 73 1573 87 1587
rect 76 1347 83 1513
rect 116 1427 123 1533
rect 73 1333 87 1347
rect 113 1333 127 1347
rect 116 1247 123 1333
rect 133 1313 147 1327
rect 136 1227 143 1313
rect 96 1147 103 1173
rect 93 1133 107 1147
rect 156 1143 163 2096
rect 176 1267 183 2513
rect 196 2307 203 2713
rect 236 2587 243 2753
rect 256 2447 263 2793
rect 376 2787 383 2973
rect 416 2863 423 2993
rect 476 2907 483 3033
rect 496 2883 503 3456
rect 556 3447 563 3473
rect 556 3247 563 3253
rect 553 3233 567 3247
rect 573 3213 587 3227
rect 533 3203 547 3207
rect 516 3196 547 3203
rect 516 3027 523 3196
rect 533 3193 547 3196
rect 576 3127 583 3213
rect 576 3047 583 3053
rect 573 3033 587 3047
rect 596 2947 603 3433
rect 636 3187 643 3473
rect 656 3307 663 3733
rect 676 3587 683 3736
rect 693 3733 707 3736
rect 713 3713 727 3727
rect 716 3707 723 3713
rect 793 3703 807 3707
rect 776 3696 807 3703
rect 896 3707 903 4293
rect 953 4203 967 4207
rect 953 4196 983 4203
rect 953 4193 967 4196
rect 916 4167 923 4193
rect 956 4027 963 4033
rect 976 4027 983 4196
rect 953 4013 967 4027
rect 716 3647 723 3693
rect 653 3223 667 3227
rect 676 3223 683 3293
rect 653 3216 683 3223
rect 653 3213 667 3216
rect 636 3047 643 3053
rect 676 3047 683 3053
rect 633 3033 647 3047
rect 496 2876 523 2883
rect 396 2856 423 2863
rect 353 2713 367 2727
rect 356 2667 363 2713
rect 276 2567 283 2653
rect 376 2607 383 2773
rect 396 2727 403 2856
rect 496 2747 503 2813
rect 473 2733 487 2747
rect 476 2727 483 2733
rect 433 2713 447 2727
rect 436 2707 443 2713
rect 313 2583 327 2587
rect 313 2576 363 2583
rect 313 2573 327 2576
rect 273 2553 287 2567
rect 356 2527 363 2576
rect 396 2547 403 2553
rect 393 2533 407 2547
rect 193 2293 207 2307
rect 236 2263 243 2293
rect 253 2273 267 2287
rect 256 2267 263 2273
rect 216 2256 243 2263
rect 196 2047 203 2093
rect 216 2023 223 2256
rect 276 2107 283 2513
rect 296 2267 303 2313
rect 356 2307 363 2313
rect 353 2293 367 2307
rect 276 2047 283 2073
rect 296 2067 303 2093
rect 273 2033 287 2047
rect 216 2016 243 2023
rect 196 1807 203 1833
rect 216 1827 223 1853
rect 236 1827 243 2016
rect 253 1773 267 1787
rect 196 1547 203 1673
rect 216 1567 223 1733
rect 256 1727 263 1773
rect 276 1607 283 1953
rect 296 1687 303 2013
rect 316 1783 323 2253
rect 376 2247 383 2533
rect 453 2523 467 2527
rect 476 2523 483 2573
rect 453 2516 483 2523
rect 453 2513 467 2516
rect 336 2087 343 2193
rect 416 2187 423 2273
rect 493 2273 507 2287
rect 473 2253 487 2267
rect 336 1967 343 2073
rect 353 2053 367 2067
rect 356 2027 363 2053
rect 336 1803 343 1833
rect 376 1827 383 1933
rect 396 1807 403 1873
rect 416 1827 423 2013
rect 353 1803 367 1807
rect 336 1796 367 1803
rect 353 1793 367 1796
rect 316 1776 343 1783
rect 233 1553 247 1567
rect 293 1583 307 1587
rect 316 1583 323 1613
rect 293 1576 323 1583
rect 293 1573 307 1576
rect 276 1567 283 1573
rect 273 1553 287 1567
rect 236 1547 243 1553
rect 196 1327 203 1333
rect 213 1273 227 1287
rect 216 1227 223 1273
rect 136 1136 163 1143
rect 76 867 83 1073
rect 136 887 143 1136
rect 216 1127 223 1153
rect 213 1113 227 1127
rect 73 853 87 867
rect 113 853 127 867
rect 116 807 123 853
rect 136 727 143 833
rect 116 607 123 633
rect 133 623 147 627
rect 156 623 163 653
rect 133 616 163 623
rect 133 613 147 616
rect 113 593 127 607
rect 156 587 163 616
rect 76 387 83 573
rect 73 373 87 387
rect 113 373 127 387
rect 116 347 123 373
rect 133 363 147 367
rect 156 363 163 533
rect 133 356 163 363
rect 133 353 147 356
rect 96 147 103 153
rect 116 147 123 333
rect 93 133 107 147
rect 156 127 163 173
rect 176 167 183 873
rect 236 867 243 1253
rect 276 1247 283 1313
rect 296 1167 303 1473
rect 316 1467 323 1576
rect 316 1267 323 1413
rect 336 1127 343 1776
rect 393 1793 407 1807
rect 413 1773 427 1787
rect 356 1727 363 1773
rect 416 1767 423 1773
rect 416 1607 423 1733
rect 393 1573 407 1587
rect 413 1593 427 1607
rect 356 1547 363 1573
rect 376 1527 383 1573
rect 396 1567 403 1573
rect 396 1487 403 1553
rect 356 1347 363 1453
rect 353 1333 367 1347
rect 393 1333 407 1347
rect 396 1327 403 1333
rect 373 1313 387 1327
rect 413 1313 427 1327
rect 376 1287 383 1313
rect 293 1123 307 1127
rect 276 1116 307 1123
rect 276 1107 283 1116
rect 293 1113 307 1116
rect 313 1093 327 1107
rect 333 1113 347 1127
rect 356 1107 363 1113
rect 376 1107 383 1253
rect 396 1127 403 1313
rect 353 1093 367 1107
rect 236 847 243 853
rect 233 833 247 847
rect 276 807 283 1093
rect 316 1087 323 1093
rect 316 827 323 1073
rect 396 1027 403 1113
rect 416 1027 423 1313
rect 436 1307 443 2253
rect 476 2247 483 2253
rect 496 2247 503 2273
rect 516 2227 523 2876
rect 616 2803 623 3033
rect 673 3033 687 3047
rect 736 3027 743 3693
rect 776 3687 783 3696
rect 793 3693 807 3696
rect 776 3507 783 3673
rect 896 3507 903 3573
rect 916 3527 923 3993
rect 973 3973 987 3987
rect 976 3967 983 3973
rect 1016 3767 1023 4473
rect 1076 4447 1083 4496
rect 1096 4427 1103 4873
rect 1113 4683 1127 4687
rect 1136 4683 1143 5093
rect 1156 4903 1163 5073
rect 1176 4967 1183 5156
rect 1196 4967 1203 5376
rect 1256 5187 1263 5373
rect 1253 5173 1267 5187
rect 1273 5153 1287 5167
rect 1276 5107 1283 5153
rect 1296 4987 1303 5173
rect 1313 5153 1327 5167
rect 1316 5127 1323 5153
rect 1336 5147 1343 5653
rect 1396 5627 1403 5656
rect 1533 5653 1547 5667
rect 1353 5613 1367 5627
rect 1413 5613 1427 5627
rect 1356 5587 1363 5613
rect 1376 5507 1383 5613
rect 1416 5607 1423 5613
rect 1536 5607 1543 5653
rect 1793 5663 1807 5667
rect 1776 5656 1807 5663
rect 1553 5633 1567 5647
rect 1556 5627 1563 5633
rect 1376 5447 1383 5493
rect 1396 5467 1403 5533
rect 1393 5453 1407 5467
rect 1373 5433 1387 5447
rect 1416 5447 1423 5593
rect 1636 5487 1643 5653
rect 1653 5613 1667 5627
rect 1713 5643 1727 5647
rect 1713 5636 1743 5643
rect 1713 5633 1727 5636
rect 1356 5167 1363 5433
rect 1513 5393 1527 5407
rect 1556 5407 1563 5433
rect 1573 5423 1587 5427
rect 1596 5423 1603 5433
rect 1573 5416 1603 5423
rect 1573 5413 1587 5416
rect 1553 5393 1567 5407
rect 1516 5183 1523 5393
rect 1496 5176 1523 5183
rect 1236 4967 1243 4973
rect 1193 4953 1207 4967
rect 1176 4947 1183 4953
rect 1173 4933 1187 4947
rect 1233 4953 1247 4967
rect 1156 4896 1183 4903
rect 1113 4676 1143 4683
rect 1113 4673 1127 4676
rect 1156 4467 1163 4673
rect 1176 4507 1183 4896
rect 1296 4787 1303 4973
rect 1356 4747 1363 5113
rect 1416 5027 1423 5153
rect 1473 5133 1487 5147
rect 1396 4723 1403 4933
rect 1413 4913 1427 4927
rect 1416 4907 1423 4913
rect 1476 4887 1483 5133
rect 1496 4927 1503 5176
rect 1396 4716 1423 4723
rect 1273 4653 1287 4667
rect 1333 4653 1347 4667
rect 1393 4673 1407 4687
rect 1373 4653 1387 4667
rect 1133 4433 1147 4447
rect 1176 4447 1183 4473
rect 1173 4433 1187 4447
rect 1036 3983 1043 4213
rect 1136 4207 1143 4433
rect 1053 4173 1067 4187
rect 1113 4203 1127 4207
rect 1113 4196 1133 4203
rect 1113 4193 1127 4196
rect 1056 4167 1063 4173
rect 1093 4153 1107 4167
rect 1096 4127 1103 4153
rect 1096 3987 1103 4013
rect 1053 3983 1067 3987
rect 1036 3976 1067 3983
rect 1053 3973 1067 3976
rect 1093 3973 1107 3987
rect 1113 3953 1127 3967
rect 956 3547 963 3753
rect 996 3727 1003 3733
rect 1036 3727 1043 3793
rect 973 3693 987 3707
rect 993 3713 1007 3727
rect 1033 3713 1047 3727
rect 1053 3703 1067 3707
rect 1076 3703 1083 3813
rect 1053 3696 1083 3703
rect 1053 3693 1067 3696
rect 976 3587 983 3693
rect 1096 3687 1103 3853
rect 1116 3767 1123 3953
rect 1156 3947 1163 4413
rect 1216 4243 1223 4633
rect 1256 4267 1263 4633
rect 1276 4547 1283 4653
rect 1336 4643 1343 4653
rect 1376 4647 1383 4653
rect 1336 4636 1363 4643
rect 1316 4507 1323 4613
rect 1276 4487 1283 4493
rect 1273 4473 1287 4487
rect 1293 4453 1307 4467
rect 1296 4447 1303 4453
rect 1356 4447 1363 4636
rect 1356 4367 1363 4433
rect 1196 4236 1223 4243
rect 1176 4003 1183 4233
rect 1196 4167 1203 4236
rect 1296 4227 1303 4253
rect 1256 4127 1263 4213
rect 1273 4203 1287 4207
rect 1273 4196 1303 4203
rect 1273 4193 1287 4196
rect 1276 4187 1283 4193
rect 1236 4007 1243 4073
rect 1276 4007 1283 4013
rect 1193 4003 1207 4007
rect 1176 3996 1207 4003
rect 1176 3827 1183 3996
rect 1193 3993 1207 3996
rect 1213 3973 1227 3987
rect 1233 3993 1247 4007
rect 1253 3973 1267 3987
rect 1273 3993 1287 4007
rect 1216 3967 1223 3973
rect 1216 3807 1223 3953
rect 1256 3867 1263 3973
rect 1296 3907 1303 4196
rect 1316 3967 1323 4253
rect 1376 4247 1383 4573
rect 1396 4547 1403 4673
rect 1416 4503 1423 4716
rect 1436 4587 1443 4713
rect 1516 4647 1523 5153
rect 1536 5147 1543 5373
rect 1596 5287 1603 5416
rect 1556 5167 1563 5273
rect 1553 5153 1567 5167
rect 1616 5163 1623 5473
rect 1656 5467 1663 5613
rect 1736 5627 1743 5636
rect 1696 5427 1703 5473
rect 1736 5467 1743 5613
rect 1693 5413 1707 5427
rect 1596 5156 1623 5163
rect 1696 5167 1703 5173
rect 1756 5167 1763 5633
rect 1776 5607 1783 5656
rect 1793 5653 1807 5656
rect 1833 5653 1847 5667
rect 1813 5633 1827 5647
rect 1816 5567 1823 5633
rect 1836 5623 1843 5653
rect 1936 5647 1943 5653
rect 2076 5647 2083 5653
rect 1853 5643 1867 5647
rect 1853 5636 1883 5643
rect 1853 5633 1867 5636
rect 1876 5627 1883 5636
rect 1933 5633 1947 5647
rect 1836 5616 1863 5623
rect 1856 5607 1863 5616
rect 2053 5613 2067 5627
rect 2073 5633 2087 5647
rect 2093 5613 2107 5627
rect 1573 5113 1587 5127
rect 1576 5107 1583 5113
rect 1576 4947 1583 4973
rect 1553 4913 1567 4927
rect 1573 4933 1587 4947
rect 1596 4927 1603 5156
rect 1616 4947 1623 5093
rect 1613 4943 1627 4947
rect 1613 4936 1643 4943
rect 1613 4933 1627 4936
rect 1593 4913 1607 4927
rect 1636 4927 1643 4936
rect 1536 4687 1543 4913
rect 1556 4907 1563 4913
rect 1556 4707 1563 4893
rect 1613 4683 1627 4687
rect 1596 4676 1627 4683
rect 1596 4663 1603 4676
rect 1613 4673 1627 4676
rect 1576 4656 1603 4663
rect 1473 4633 1487 4647
rect 1476 4627 1483 4633
rect 1436 4507 1443 4533
rect 1396 4496 1423 4503
rect 1396 4263 1403 4496
rect 1433 4493 1447 4507
rect 1396 4256 1423 4263
rect 1387 4236 1403 4243
rect 1396 4227 1403 4236
rect 1393 4213 1407 4227
rect 1133 3713 1147 3727
rect 1136 3707 1143 3713
rect 1016 3527 1023 3673
rect 973 3523 987 3527
rect 956 3516 987 3523
rect 753 3473 767 3487
rect 773 3493 787 3507
rect 793 3473 807 3487
rect 873 3473 887 3487
rect 893 3493 907 3507
rect 756 3227 763 3473
rect 796 3467 803 3473
rect 876 3447 883 3473
rect 816 3223 823 3433
rect 836 3267 843 3293
rect 833 3253 847 3267
rect 853 3233 867 3247
rect 816 3216 843 3223
rect 693 3023 707 3027
rect 693 3016 723 3023
rect 693 3013 707 3016
rect 656 2967 663 2993
rect 616 2796 643 2803
rect 573 2783 587 2787
rect 556 2776 587 2783
rect 536 2687 543 2753
rect 556 2747 563 2776
rect 573 2773 587 2776
rect 456 1267 463 2213
rect 476 2067 483 2173
rect 536 2107 543 2233
rect 576 2227 583 2733
rect 636 2707 643 2796
rect 656 2767 663 2953
rect 716 2947 723 3016
rect 836 3027 843 3216
rect 856 3167 863 3233
rect 756 2987 763 3013
rect 756 2727 763 2973
rect 776 2747 783 2793
rect 796 2787 803 2993
rect 856 2827 863 3093
rect 816 2787 823 2793
rect 856 2787 863 2813
rect 813 2773 827 2787
rect 853 2773 867 2787
rect 636 2567 643 2653
rect 633 2553 647 2567
rect 676 2567 683 2673
rect 593 2273 607 2287
rect 596 2207 603 2273
rect 613 2253 627 2267
rect 653 2263 667 2267
rect 676 2263 683 2293
rect 653 2256 683 2263
rect 653 2253 667 2256
rect 616 2207 623 2253
rect 656 2247 663 2253
rect 533 2093 547 2107
rect 513 2053 527 2067
rect 476 1747 483 2053
rect 516 2047 523 2053
rect 516 1847 523 1873
rect 496 1827 503 1833
rect 493 1813 507 1827
rect 513 1793 527 1807
rect 516 1747 523 1793
rect 496 1736 513 1743
rect 496 1587 503 1736
rect 516 1607 523 1713
rect 536 1623 543 1813
rect 556 1727 563 1773
rect 576 1647 583 2133
rect 636 2087 643 2213
rect 633 2073 647 2087
rect 616 2067 623 2073
rect 613 2053 627 2067
rect 653 2053 667 2067
rect 656 1947 663 2053
rect 716 2027 723 2673
rect 736 2547 743 2693
rect 876 2687 883 3193
rect 896 2807 903 3453
rect 916 3267 923 3473
rect 916 3047 923 3213
rect 936 3167 943 3493
rect 956 3447 963 3516
rect 973 3513 987 3516
rect 1013 3513 1027 3527
rect 973 3233 987 3247
rect 1013 3233 1027 3247
rect 976 3207 983 3233
rect 976 3047 983 3173
rect 913 3033 927 3047
rect 996 2883 1003 3153
rect 1016 3087 1023 3233
rect 1036 3147 1043 3353
rect 976 2876 1003 2883
rect 896 2727 903 2773
rect 936 2767 943 2773
rect 976 2767 983 2876
rect 973 2753 987 2767
rect 756 2567 763 2573
rect 796 2567 803 2593
rect 753 2553 767 2567
rect 793 2553 807 2567
rect 816 2547 823 2553
rect 876 2547 883 2573
rect 813 2533 827 2547
rect 896 2447 903 2713
rect 936 2587 943 2693
rect 933 2573 947 2587
rect 953 2533 967 2547
rect 756 2307 763 2433
rect 936 2307 943 2533
rect 753 2293 767 2307
rect 793 2293 807 2307
rect 773 2273 787 2287
rect 776 2207 783 2273
rect 796 2127 803 2293
rect 913 2273 927 2287
rect 933 2293 947 2307
rect 856 2087 863 2273
rect 916 2147 923 2273
rect 956 2267 963 2533
rect 773 2053 787 2067
rect 776 2047 783 2053
rect 816 2027 823 2033
rect 716 1847 723 1853
rect 536 1616 553 1623
rect 513 1593 527 1607
rect 573 1583 587 1587
rect 596 1583 603 1793
rect 653 1773 667 1787
rect 573 1576 603 1583
rect 573 1573 587 1576
rect 536 1347 543 1573
rect 596 1567 603 1576
rect 476 1303 483 1333
rect 476 1296 503 1303
rect 496 1283 503 1296
rect 556 1287 563 1293
rect 496 1276 543 1283
rect 536 1267 543 1276
rect 436 1147 443 1173
rect 436 1127 443 1133
rect 476 1127 483 1233
rect 433 1113 447 1127
rect 453 1093 467 1107
rect 473 1113 487 1127
rect 456 1087 463 1093
rect 356 867 363 1013
rect 516 967 523 1253
rect 536 1087 543 1213
rect 353 853 367 867
rect 393 853 407 867
rect 376 807 383 833
rect 396 807 403 853
rect 413 843 427 847
rect 436 843 443 853
rect 413 836 443 843
rect 413 833 427 836
rect 216 463 223 793
rect 236 647 243 793
rect 233 633 247 647
rect 196 456 223 463
rect 196 343 203 456
rect 296 367 303 413
rect 233 343 247 347
rect 196 336 247 343
rect 233 333 247 336
rect 273 333 287 347
rect 176 127 183 153
rect 256 167 263 313
rect 276 267 283 333
rect 296 327 303 353
rect 316 347 323 613
rect 336 307 343 793
rect 356 603 363 713
rect 373 603 387 607
rect 356 596 387 603
rect 433 623 447 627
rect 456 623 463 653
rect 433 616 463 623
rect 433 613 447 616
rect 373 593 387 596
rect 456 547 463 616
rect 416 367 423 373
rect 373 353 387 367
rect 376 347 383 353
rect 393 333 407 347
rect 433 333 447 347
rect 396 307 403 333
rect 436 327 443 333
rect 376 167 383 253
rect 416 187 423 193
rect 413 173 427 187
rect 233 133 247 147
rect 253 153 267 167
rect 373 153 387 167
rect 433 143 447 147
rect 456 143 463 353
rect 476 247 483 953
rect 576 907 583 1313
rect 616 1147 623 1633
rect 656 1587 663 1773
rect 716 1767 723 1833
rect 796 1807 803 1813
rect 836 1807 843 2073
rect 873 2063 887 2067
rect 856 2056 887 2063
rect 856 2047 863 2056
rect 873 2053 887 2056
rect 896 2047 903 2093
rect 916 2067 923 2113
rect 933 2033 947 2047
rect 753 1803 767 1807
rect 736 1796 767 1803
rect 673 1763 687 1767
rect 673 1756 693 1763
rect 673 1753 687 1756
rect 736 1707 743 1796
rect 753 1793 767 1796
rect 793 1793 807 1807
rect 856 1747 863 2033
rect 936 2027 943 2033
rect 956 1827 963 2013
rect 976 1787 983 2513
rect 996 2427 1003 2593
rect 1016 2323 1023 3033
rect 1036 3027 1043 3133
rect 1036 2527 1043 2913
rect 1056 2543 1063 3533
rect 1096 3467 1103 3513
rect 1116 3483 1123 3553
rect 1156 3507 1163 3513
rect 1133 3483 1147 3487
rect 1116 3476 1147 3483
rect 1153 3493 1167 3507
rect 1176 3487 1183 3753
rect 1296 3747 1303 3833
rect 1196 3627 1203 3733
rect 1273 3713 1287 3727
rect 1293 3733 1307 3747
rect 1216 3527 1223 3613
rect 1193 3503 1207 3507
rect 1193 3496 1223 3503
rect 1193 3493 1207 3496
rect 1133 3473 1147 3476
rect 1216 3463 1223 3496
rect 1196 3456 1223 3463
rect 1076 3107 1083 3313
rect 1133 3253 1147 3267
rect 1136 3187 1143 3253
rect 1153 3243 1167 3247
rect 1176 3243 1183 3273
rect 1153 3236 1183 3243
rect 1153 3233 1167 3236
rect 1176 3147 1183 3213
rect 1073 2993 1087 3007
rect 1113 2993 1127 3007
rect 1076 2987 1083 2993
rect 1096 2803 1103 2973
rect 1116 2967 1123 2993
rect 1096 2796 1123 2803
rect 1116 2787 1123 2796
rect 1093 2753 1107 2767
rect 1113 2773 1127 2787
rect 1096 2587 1103 2753
rect 1136 2567 1143 3113
rect 1156 3007 1163 3073
rect 1156 2847 1163 2933
rect 1073 2543 1087 2547
rect 1056 2536 1087 2543
rect 996 2316 1023 2323
rect 996 2083 1003 2316
rect 1056 2303 1063 2536
rect 1073 2533 1087 2536
rect 1133 2553 1147 2567
rect 1156 2523 1163 2833
rect 1176 2607 1183 3053
rect 1196 2687 1203 3456
rect 1236 3327 1243 3713
rect 1276 3627 1283 3713
rect 1316 3647 1323 3933
rect 1336 3767 1343 4013
rect 1356 3747 1363 4173
rect 1416 4003 1423 4256
rect 1436 4207 1443 4453
rect 1456 4183 1463 4473
rect 1476 4347 1483 4613
rect 1536 4487 1543 4513
rect 1513 4453 1527 4467
rect 1533 4473 1547 4487
rect 1556 4467 1563 4473
rect 1553 4453 1567 4467
rect 1516 4427 1523 4453
rect 1516 4227 1523 4233
rect 1493 4193 1507 4207
rect 1513 4213 1527 4227
rect 1456 4176 1483 4183
rect 1416 3996 1443 4003
rect 1396 3987 1403 3993
rect 1373 3953 1387 3967
rect 1393 3973 1407 3987
rect 1413 3953 1427 3967
rect 1376 3947 1383 3953
rect 1336 3527 1343 3733
rect 1293 3473 1307 3487
rect 1296 3467 1303 3473
rect 1256 3303 1263 3453
rect 1236 3296 1263 3303
rect 1216 3247 1223 3253
rect 1236 3247 1243 3296
rect 1256 3247 1263 3273
rect 1273 3213 1287 3227
rect 1233 3193 1247 3207
rect 1236 3187 1243 3193
rect 1216 3047 1223 3153
rect 1236 3067 1243 3133
rect 1276 3067 1283 3213
rect 1296 3127 1303 3433
rect 1336 3147 1343 3493
rect 1356 3487 1363 3733
rect 1396 3727 1403 3753
rect 1416 3747 1423 3953
rect 1436 3747 1443 3996
rect 1456 3727 1463 3993
rect 1393 3673 1407 3687
rect 1396 3667 1403 3673
rect 1376 3607 1383 3633
rect 1376 3447 1383 3593
rect 1416 3507 1423 3513
rect 1413 3493 1427 3507
rect 1233 3053 1247 3067
rect 1213 3033 1227 3047
rect 1316 3047 1323 3053
rect 1356 3047 1363 3293
rect 1393 3193 1407 3207
rect 1396 3127 1403 3193
rect 1253 3043 1267 3047
rect 1253 3036 1283 3043
rect 1253 3033 1267 3036
rect 1276 2967 1283 3036
rect 1313 3033 1327 3047
rect 1296 2827 1303 3033
rect 1353 3033 1367 3047
rect 1373 3023 1387 3027
rect 1373 3016 1403 3023
rect 1373 3013 1387 3016
rect 1396 2927 1403 3016
rect 1416 3007 1423 3453
rect 1476 3407 1483 4176
rect 1496 4047 1503 4193
rect 1536 4047 1543 4193
rect 1556 4127 1563 4413
rect 1576 4163 1583 4656
rect 1596 4627 1603 4633
rect 1596 4427 1603 4613
rect 1616 4207 1623 4653
rect 1656 4527 1663 5153
rect 1693 5153 1707 5167
rect 1696 4947 1703 5113
rect 1716 4967 1723 4973
rect 1756 4967 1763 5133
rect 1776 5127 1783 5413
rect 1836 5407 1843 5593
rect 1916 5587 1923 5593
rect 1856 5427 1863 5453
rect 1853 5413 1867 5427
rect 1833 5393 1847 5407
rect 1916 5187 1923 5573
rect 1956 5427 1963 5433
rect 1933 5393 1947 5407
rect 1953 5413 1967 5427
rect 1976 5407 1983 5473
rect 2056 5467 2063 5613
rect 2096 5467 2103 5613
rect 2116 5607 2123 5653
rect 2493 5663 2507 5667
rect 2573 5663 2587 5667
rect 1993 5423 2007 5427
rect 1993 5416 2023 5423
rect 1993 5413 2007 5416
rect 1936 5183 1943 5393
rect 2016 5387 2023 5416
rect 1936 5176 1963 5183
rect 1896 5167 1903 5173
rect 1893 5163 1907 5167
rect 1713 4953 1727 4967
rect 1693 4943 1707 4947
rect 1676 4936 1707 4943
rect 1676 4907 1683 4936
rect 1693 4933 1707 4936
rect 1753 4953 1767 4967
rect 1776 4947 1783 5033
rect 1796 4947 1803 5153
rect 1873 5133 1887 5147
rect 1893 5156 1923 5163
rect 1893 5153 1907 5156
rect 1876 5127 1883 5133
rect 1916 5047 1923 5156
rect 1813 4933 1827 4947
rect 1956 4963 1963 5176
rect 1996 4983 2003 5193
rect 2016 5143 2023 5213
rect 2036 5207 2043 5413
rect 2096 5387 2103 5393
rect 2056 5167 2063 5173
rect 2096 5167 2103 5193
rect 2136 5167 2143 5633
rect 2153 5613 2167 5627
rect 2213 5633 2227 5647
rect 2293 5643 2307 5647
rect 2276 5636 2307 5643
rect 2216 5627 2223 5633
rect 2193 5613 2207 5627
rect 2156 5607 2163 5613
rect 2196 5607 2203 5613
rect 2216 5563 2223 5613
rect 2276 5567 2283 5636
rect 2293 5633 2307 5636
rect 2353 5623 2367 5627
rect 2376 5623 2383 5653
rect 2493 5656 2523 5663
rect 2493 5653 2507 5656
rect 2353 5616 2383 5623
rect 2353 5613 2367 5616
rect 2313 5593 2327 5607
rect 2316 5587 2323 5593
rect 2196 5556 2223 5563
rect 2196 5423 2203 5556
rect 2316 5447 2323 5553
rect 2376 5547 2383 5616
rect 2416 5467 2423 5633
rect 2516 5467 2523 5656
rect 2556 5656 2587 5663
rect 2556 5487 2563 5656
rect 2573 5653 2587 5656
rect 2733 5633 2747 5647
rect 2833 5663 2847 5667
rect 2816 5656 2847 5663
rect 2773 5633 2787 5647
rect 2213 5423 2227 5427
rect 2196 5416 2227 5423
rect 2313 5433 2327 5447
rect 2373 5443 2387 5447
rect 2416 5443 2423 5453
rect 2433 5443 2447 5447
rect 2373 5436 2403 5443
rect 2373 5433 2387 5436
rect 2176 5187 2183 5293
rect 2196 5227 2203 5416
rect 2213 5413 2227 5416
rect 2333 5393 2347 5407
rect 2336 5307 2343 5393
rect 2396 5207 2403 5436
rect 2416 5436 2447 5443
rect 2216 5187 2223 5193
rect 2173 5183 2187 5187
rect 2156 5176 2187 5183
rect 2033 5143 2047 5147
rect 2016 5136 2047 5143
rect 2053 5153 2067 5167
rect 2033 5133 2047 5136
rect 2093 5153 2107 5167
rect 2113 5133 2127 5147
rect 2116 5107 2123 5133
rect 2156 5107 2163 5176
rect 2173 5173 2187 5176
rect 2213 5173 2227 5187
rect 1996 4976 2023 4983
rect 1936 4956 1963 4963
rect 1816 4927 1823 4933
rect 1816 4807 1823 4913
rect 1716 4683 1723 4693
rect 1733 4683 1747 4687
rect 1716 4676 1747 4683
rect 1716 4667 1723 4676
rect 1733 4673 1747 4676
rect 1753 4653 1767 4667
rect 1676 4467 1683 4593
rect 1716 4467 1723 4633
rect 1756 4563 1763 4653
rect 1736 4556 1763 4563
rect 1653 4433 1667 4447
rect 1673 4453 1687 4467
rect 1693 4433 1707 4447
rect 1656 4227 1663 4433
rect 1696 4407 1703 4433
rect 1633 4173 1647 4187
rect 1576 4156 1603 4163
rect 1536 4027 1543 4033
rect 1533 4013 1547 4027
rect 1513 3973 1527 3987
rect 1516 3747 1523 3973
rect 1556 3947 1563 4033
rect 1536 3727 1543 3753
rect 1496 3687 1503 3713
rect 1533 3713 1547 3727
rect 1596 3647 1603 4156
rect 1636 4127 1643 4173
rect 1656 4163 1663 4213
rect 1676 4187 1683 4273
rect 1736 4267 1743 4556
rect 1756 4443 1763 4533
rect 1796 4467 1803 4493
rect 1773 4443 1787 4447
rect 1756 4436 1787 4443
rect 1793 4453 1807 4467
rect 1816 4447 1823 4533
rect 1836 4467 1843 4573
rect 1773 4433 1787 4436
rect 1796 4227 1803 4413
rect 1856 4387 1863 4893
rect 1896 4723 1903 4933
rect 1916 4927 1923 4953
rect 1887 4716 1903 4723
rect 1876 4707 1883 4713
rect 1873 4693 1887 4707
rect 1913 4703 1927 4707
rect 1936 4703 1943 4956
rect 1993 4923 2007 4927
rect 2016 4923 2023 4976
rect 2096 4967 2103 5033
rect 2093 4953 2107 4967
rect 2196 4947 2203 5153
rect 2276 4987 2283 5153
rect 2356 5067 2363 5173
rect 2373 5153 2387 5167
rect 2376 5127 2383 5153
rect 2416 5147 2423 5436
rect 2433 5433 2447 5436
rect 2453 5413 2467 5427
rect 2496 5427 2503 5453
rect 2493 5413 2507 5427
rect 2456 5403 2463 5413
rect 2436 5396 2463 5403
rect 2273 4973 2287 4987
rect 2356 4947 2363 5053
rect 2436 5047 2443 5396
rect 2556 5387 2563 5433
rect 2476 5167 2483 5173
rect 2473 5153 2487 5167
rect 2527 5156 2543 5163
rect 2376 4967 2383 4973
rect 2373 4953 2387 4967
rect 2153 4933 2167 4947
rect 2353 4933 2367 4947
rect 2156 4927 2163 4933
rect 1993 4916 2023 4923
rect 1993 4913 2007 4916
rect 1893 4673 1907 4687
rect 1913 4696 1943 4703
rect 1913 4693 1927 4696
rect 1713 4223 1727 4227
rect 1696 4216 1727 4223
rect 1656 4156 1683 4163
rect 1616 4103 1623 4113
rect 1616 4096 1663 4103
rect 1656 4047 1663 4096
rect 1656 4007 1663 4013
rect 1653 3993 1667 4007
rect 1556 3527 1563 3633
rect 1513 3523 1527 3527
rect 1496 3516 1527 3523
rect 1496 3287 1503 3516
rect 1513 3513 1527 3516
rect 1553 3513 1567 3527
rect 1513 3253 1527 3267
rect 1493 3233 1507 3247
rect 1233 2753 1247 2767
rect 1236 2667 1243 2753
rect 1253 2733 1267 2747
rect 1316 2747 1323 2773
rect 1293 2733 1307 2747
rect 1136 2516 1163 2523
rect 1036 2296 1063 2303
rect 1016 2287 1023 2293
rect 1013 2273 1027 2287
rect 1036 2247 1043 2296
rect 1053 2253 1067 2267
rect 1056 2227 1063 2253
rect 1096 2227 1103 2393
rect 1116 2087 1123 2293
rect 1136 2287 1143 2516
rect 1133 2273 1147 2287
rect 996 2076 1023 2083
rect 996 1767 1003 2053
rect 1016 1887 1023 2076
rect 1116 2067 1123 2073
rect 1113 2053 1127 2067
rect 1136 1847 1143 2073
rect 1053 1793 1067 1807
rect 1036 1767 1043 1793
rect 953 1753 967 1767
rect 956 1747 963 1753
rect 736 1627 743 1693
rect 653 1573 667 1587
rect 673 1563 687 1567
rect 696 1563 703 1613
rect 856 1587 863 1733
rect 896 1607 903 1613
rect 936 1607 943 1653
rect 893 1593 907 1607
rect 876 1587 883 1593
rect 873 1573 887 1587
rect 933 1593 947 1607
rect 673 1556 703 1563
rect 673 1553 687 1556
rect 633 1313 647 1327
rect 636 1307 643 1313
rect 653 1293 667 1307
rect 693 1293 707 1307
rect 656 1267 663 1293
rect 616 1107 623 1113
rect 656 1107 663 1153
rect 613 1093 627 1107
rect 653 1093 667 1107
rect 676 1087 683 1133
rect 696 1123 703 1293
rect 756 1127 763 1533
rect 956 1527 963 1733
rect 976 1587 983 1613
rect 816 1347 823 1353
rect 916 1347 923 1353
rect 813 1333 827 1347
rect 913 1333 927 1347
rect 853 1303 867 1307
rect 876 1303 883 1333
rect 933 1313 947 1327
rect 853 1296 883 1303
rect 853 1293 867 1296
rect 936 1167 943 1313
rect 713 1123 727 1127
rect 696 1116 727 1123
rect 696 1087 703 1116
rect 713 1113 727 1116
rect 733 1093 747 1107
rect 753 1113 767 1127
rect 776 1107 783 1153
rect 996 1147 1003 1753
rect 1056 1747 1063 1793
rect 1073 1773 1087 1787
rect 1076 1603 1083 1773
rect 1136 1687 1143 1753
rect 1056 1596 1083 1603
rect 1036 1587 1043 1593
rect 1013 1553 1027 1567
rect 1056 1567 1063 1596
rect 1073 1583 1087 1587
rect 1096 1583 1103 1653
rect 1073 1576 1103 1583
rect 1073 1573 1087 1576
rect 1053 1553 1067 1567
rect 1016 1367 1023 1553
rect 1073 1283 1087 1287
rect 1096 1283 1103 1576
rect 1136 1563 1143 1673
rect 1156 1607 1163 2253
rect 1176 2227 1183 2573
rect 1256 2563 1263 2733
rect 1296 2707 1303 2733
rect 1336 2727 1343 2753
rect 1353 2733 1367 2747
rect 1356 2667 1363 2733
rect 1313 2563 1327 2567
rect 1373 2563 1387 2567
rect 1256 2556 1283 2563
rect 1196 2447 1203 2533
rect 1213 2513 1227 2527
rect 1276 2527 1283 2556
rect 1313 2556 1343 2563
rect 1313 2553 1327 2556
rect 1253 2523 1267 2527
rect 1253 2516 1273 2523
rect 1253 2513 1267 2516
rect 1216 2507 1223 2513
rect 1336 2507 1343 2556
rect 1373 2556 1403 2563
rect 1373 2553 1387 2556
rect 1196 2203 1203 2433
rect 1396 2347 1403 2556
rect 1416 2547 1423 2553
rect 1416 2307 1423 2533
rect 1436 2307 1443 3233
rect 1496 3207 1503 3233
rect 1516 3227 1523 3253
rect 1533 3243 1547 3247
rect 1556 3243 1563 3273
rect 1533 3236 1563 3243
rect 1533 3233 1547 3236
rect 1496 3027 1503 3073
rect 1493 3013 1507 3027
rect 1516 3007 1523 3053
rect 1536 3027 1543 3113
rect 1513 2993 1527 3007
rect 1556 2987 1563 3193
rect 1576 3067 1583 3253
rect 1596 3247 1603 3613
rect 1616 3487 1623 3493
rect 1616 3267 1623 3473
rect 1636 3467 1643 3973
rect 1676 3867 1683 4156
rect 1696 4147 1703 4216
rect 1713 4213 1727 4216
rect 1733 4193 1747 4207
rect 1736 4187 1743 4193
rect 1816 4167 1823 4373
rect 1696 3987 1703 4033
rect 1676 3727 1683 3733
rect 1673 3713 1687 3727
rect 1716 3567 1723 4153
rect 1816 3987 1823 4033
rect 1836 4027 1843 4253
rect 1856 4227 1863 4273
rect 1896 4267 1903 4673
rect 1956 4667 1963 4913
rect 1996 4687 2003 4913
rect 1973 4663 1987 4667
rect 1967 4656 1987 4663
rect 2033 4673 2047 4687
rect 1973 4653 1987 4656
rect 2013 4653 2027 4667
rect 1936 4507 1943 4553
rect 2016 4527 2023 4653
rect 2036 4647 2043 4673
rect 1933 4493 1947 4507
rect 1956 4487 1963 4493
rect 1953 4473 1967 4487
rect 1936 4267 1943 4453
rect 1976 4363 1983 4513
rect 2027 4496 2043 4503
rect 2036 4487 2043 4496
rect 2016 4443 2023 4473
rect 2033 4443 2047 4447
rect 2016 4436 2047 4443
rect 2076 4447 2083 4673
rect 2096 4587 2103 4653
rect 2096 4467 2103 4573
rect 2093 4453 2107 4467
rect 2033 4433 2047 4436
rect 1956 4356 1983 4363
rect 1853 4213 1867 4227
rect 1893 4213 1907 4227
rect 1873 4193 1887 4207
rect 1876 4187 1883 4193
rect 1733 3973 1747 3987
rect 1813 3973 1827 3987
rect 1736 3727 1743 3973
rect 1836 3967 1843 4013
rect 1876 4007 1883 4173
rect 1896 4167 1903 4213
rect 1936 4207 1943 4253
rect 1913 4203 1927 4207
rect 1913 4196 1933 4203
rect 1913 4193 1927 4196
rect 1833 3953 1847 3967
rect 1873 3953 1887 3967
rect 1876 3767 1883 3953
rect 1896 3767 1903 3973
rect 1816 3747 1823 3753
rect 1773 3743 1787 3747
rect 1756 3736 1787 3743
rect 1756 3707 1763 3736
rect 1773 3733 1787 3736
rect 1793 3713 1807 3727
rect 1813 3733 1827 3747
rect 1913 3743 1927 3747
rect 1913 3736 1943 3743
rect 1913 3733 1927 3736
rect 1656 3487 1663 3533
rect 1693 3503 1707 3507
rect 1733 3503 1747 3507
rect 1756 3503 1763 3573
rect 1693 3496 1723 3503
rect 1693 3493 1707 3496
rect 1673 3243 1687 3247
rect 1696 3243 1703 3473
rect 1716 3247 1723 3496
rect 1733 3496 1763 3503
rect 1733 3493 1747 3496
rect 1736 3287 1743 3493
rect 1756 3263 1763 3453
rect 1776 3307 1783 3493
rect 1736 3256 1763 3263
rect 1673 3236 1703 3243
rect 1673 3233 1687 3236
rect 1676 3227 1683 3233
rect 1476 2563 1483 2753
rect 1496 2747 1503 2953
rect 1573 2713 1587 2727
rect 1576 2647 1583 2713
rect 1596 2707 1603 3093
rect 1616 2887 1623 3133
rect 1716 3027 1723 3233
rect 1736 3123 1743 3256
rect 1776 3247 1783 3293
rect 1796 3247 1803 3713
rect 1936 3667 1943 3736
rect 1956 3707 1963 4356
rect 2056 4247 2063 4413
rect 2116 4267 2123 4773
rect 2136 4707 2143 4733
rect 2133 4693 2147 4707
rect 2173 4693 2187 4707
rect 2153 4673 2167 4687
rect 2156 4467 2163 4673
rect 2176 4647 2183 4693
rect 2193 4673 2207 4687
rect 2196 4667 2203 4673
rect 2176 4547 2183 4633
rect 2216 4487 2223 4493
rect 2156 4287 2163 4453
rect 2176 4443 2183 4473
rect 2216 4467 2223 4473
rect 2193 4443 2207 4447
rect 2176 4436 2207 4443
rect 2213 4453 2227 4467
rect 2236 4447 2243 4713
rect 2416 4707 2423 4733
rect 2373 4703 2387 4707
rect 2356 4696 2387 4703
rect 2356 4687 2363 4696
rect 2373 4693 2387 4696
rect 2413 4693 2427 4707
rect 2436 4687 2443 5013
rect 2313 4653 2327 4667
rect 2256 4467 2263 4653
rect 2316 4627 2323 4653
rect 2253 4453 2267 4467
rect 2193 4433 2207 4436
rect 2233 4433 2247 4447
rect 1993 4213 2007 4227
rect 1996 4167 2003 4213
rect 2056 4187 2063 4233
rect 1976 3987 1983 4093
rect 1996 4007 2003 4053
rect 2036 4007 2043 4053
rect 1993 3993 2007 4007
rect 2013 3973 2027 3987
rect 2033 3993 2047 4007
rect 2016 3947 2023 3973
rect 1976 3687 1983 3933
rect 2056 3807 2063 4093
rect 2076 3987 2083 4213
rect 2096 4203 2103 4253
rect 2176 4227 2183 4233
rect 2113 4203 2127 4207
rect 2096 4196 2127 4203
rect 2113 4193 2127 4196
rect 1996 3727 2003 3753
rect 2013 3703 2027 3707
rect 2036 3703 2043 3733
rect 2056 3727 2063 3733
rect 2013 3696 2043 3703
rect 2053 3713 2067 3727
rect 2013 3693 2027 3696
rect 1993 3673 2007 3687
rect 1996 3667 2003 3673
rect 1836 3507 1843 3513
rect 1833 3493 1847 3507
rect 1856 3487 1863 3493
rect 1853 3473 1867 3487
rect 1896 3307 1903 3633
rect 1916 3507 1923 3533
rect 1996 3527 2003 3553
rect 1933 3493 1947 3507
rect 1973 3493 1987 3507
rect 1993 3513 2007 3527
rect 2016 3507 2023 3513
rect 1816 3247 1823 3273
rect 1753 3213 1767 3227
rect 1773 3233 1787 3247
rect 1813 3233 1827 3247
rect 1756 3167 1763 3213
rect 1736 3116 1763 3123
rect 1693 3013 1707 3027
rect 1656 2967 1663 3013
rect 1696 3007 1703 3013
rect 1716 2983 1723 3013
rect 1736 3007 1743 3073
rect 1716 2976 1743 2983
rect 1673 2733 1687 2747
rect 1676 2727 1683 2733
rect 1653 2713 1667 2727
rect 1656 2707 1663 2713
rect 1476 2556 1503 2563
rect 1496 2547 1503 2556
rect 1473 2513 1487 2527
rect 1493 2533 1507 2547
rect 1476 2507 1483 2513
rect 1293 2293 1307 2307
rect 1296 2247 1303 2293
rect 1313 2283 1327 2287
rect 1336 2283 1343 2293
rect 1416 2287 1423 2293
rect 1456 2287 1463 2373
rect 1313 2276 1343 2283
rect 1313 2273 1327 2276
rect 1393 2253 1407 2267
rect 1413 2273 1427 2287
rect 1176 2196 1203 2203
rect 1176 1807 1183 2196
rect 1276 2067 1283 2093
rect 1236 1807 1243 1833
rect 1193 1793 1207 1807
rect 1196 1767 1203 1793
rect 1213 1773 1227 1787
rect 1153 1563 1167 1567
rect 1136 1556 1167 1563
rect 1153 1553 1167 1556
rect 1153 1333 1167 1347
rect 1156 1307 1163 1333
rect 1216 1327 1223 1773
rect 1276 1607 1283 1793
rect 1296 1647 1303 2213
rect 1356 2087 1363 2113
rect 1396 2107 1403 2253
rect 1353 2073 1367 2087
rect 1333 2063 1347 2067
rect 1316 2056 1347 2063
rect 1316 1727 1323 2056
rect 1333 2053 1347 2056
rect 1396 1787 1403 1933
rect 1353 1763 1367 1767
rect 1353 1756 1383 1763
rect 1353 1753 1367 1756
rect 1273 1603 1287 1607
rect 1256 1596 1287 1603
rect 1316 1607 1323 1673
rect 1256 1567 1263 1596
rect 1273 1593 1287 1596
rect 1313 1593 1327 1607
rect 1256 1343 1263 1513
rect 1316 1347 1323 1553
rect 1273 1343 1287 1347
rect 1256 1336 1287 1343
rect 1256 1287 1263 1336
rect 1273 1333 1287 1336
rect 1293 1313 1307 1327
rect 1313 1333 1327 1347
rect 1296 1307 1303 1313
rect 1073 1276 1103 1283
rect 1073 1273 1087 1276
rect 676 1027 683 1073
rect 556 847 563 853
rect 616 827 623 893
rect 636 867 643 1013
rect 736 907 743 1093
rect 633 853 647 867
rect 653 833 667 847
rect 693 843 707 847
rect 676 836 707 843
rect 656 787 663 833
rect 676 767 683 836
rect 693 833 707 836
rect 716 823 723 853
rect 796 847 803 853
rect 753 843 767 847
rect 696 816 723 823
rect 736 836 767 843
rect 573 643 587 647
rect 553 613 567 627
rect 573 636 603 643
rect 573 633 587 636
rect 596 627 603 636
rect 696 647 703 816
rect 736 787 743 836
rect 753 833 767 836
rect 793 833 807 847
rect 773 793 787 807
rect 776 767 783 793
rect 633 613 647 627
rect 693 633 707 647
rect 516 387 523 533
rect 556 427 563 613
rect 513 373 527 387
rect 553 373 567 387
rect 476 147 483 233
rect 516 147 523 213
rect 556 207 563 373
rect 573 353 587 367
rect 576 247 583 353
rect 596 267 603 613
rect 636 607 643 613
rect 773 593 787 607
rect 813 603 827 607
rect 836 603 843 1113
rect 936 1127 943 1133
rect 913 1103 927 1107
rect 896 1096 927 1103
rect 933 1113 947 1127
rect 1093 1123 1107 1127
rect 896 1087 903 1096
rect 913 1093 927 1096
rect 1073 1093 1087 1107
rect 1093 1116 1123 1123
rect 1093 1113 1107 1116
rect 1116 1107 1123 1116
rect 1076 1083 1083 1093
rect 1076 1076 1113 1083
rect 856 607 863 833
rect 813 596 843 603
rect 813 593 827 596
rect 776 587 783 593
rect 676 387 683 573
rect 816 407 823 593
rect 673 373 687 387
rect 713 343 727 347
rect 736 343 743 393
rect 833 373 847 387
rect 813 353 827 367
rect 713 336 743 343
rect 713 333 727 336
rect 816 287 823 353
rect 536 167 543 173
rect 576 167 583 173
rect 636 167 643 173
rect 676 167 683 193
rect 533 153 547 167
rect 433 136 463 143
rect 433 133 447 136
rect 513 133 527 147
rect 573 153 587 167
rect 633 153 647 167
rect 673 153 687 167
rect 816 147 823 273
rect 836 227 843 373
rect 853 363 867 367
rect 876 363 883 873
rect 896 827 903 1073
rect 1136 867 1143 1153
rect 1173 1093 1187 1107
rect 1176 1083 1183 1093
rect 1167 1076 1183 1083
rect 1216 887 1223 1113
rect 1316 1127 1323 1273
rect 1336 1147 1343 1613
rect 1253 1093 1267 1107
rect 1313 1113 1327 1127
rect 1256 1087 1263 1093
rect 1053 863 1067 867
rect 1036 856 1067 863
rect 933 813 947 827
rect 1016 827 1023 833
rect 973 813 987 827
rect 936 807 943 813
rect 936 627 943 673
rect 956 647 963 773
rect 976 667 983 813
rect 996 647 1003 653
rect 953 633 967 647
rect 933 613 947 627
rect 993 633 1007 647
rect 1016 627 1023 813
rect 1036 767 1043 856
rect 1053 853 1067 856
rect 1093 853 1107 867
rect 1096 807 1103 853
rect 1136 847 1143 853
rect 1113 833 1127 847
rect 1096 647 1103 793
rect 1116 783 1123 833
rect 1136 807 1143 833
rect 1173 813 1187 827
rect 1233 833 1247 847
rect 1176 807 1183 813
rect 1236 807 1243 833
rect 1116 776 1143 783
rect 1096 627 1103 633
rect 956 367 963 373
rect 976 367 983 613
rect 1093 613 1107 627
rect 1116 607 1123 673
rect 1136 627 1143 776
rect 1216 667 1223 673
rect 1213 653 1227 667
rect 1113 593 1127 607
rect 1156 547 1163 633
rect 1256 647 1263 1053
rect 1296 827 1303 1033
rect 1336 887 1343 1133
rect 1356 1047 1363 1733
rect 1376 1727 1383 1756
rect 1416 1747 1423 2213
rect 1476 2147 1483 2293
rect 1496 2267 1503 2453
rect 1516 2227 1523 2273
rect 1536 2263 1543 2493
rect 1556 2487 1563 2513
rect 1576 2507 1583 2613
rect 1596 2587 1603 2653
rect 1593 2573 1607 2587
rect 1636 2527 1643 2693
rect 1676 2643 1683 2713
rect 1667 2636 1683 2643
rect 1696 2607 1703 2973
rect 1656 2563 1663 2593
rect 1736 2567 1743 2976
rect 1756 2707 1763 3116
rect 1796 3047 1803 3173
rect 1836 3047 1843 3133
rect 1793 3033 1807 3047
rect 1793 2783 1807 2787
rect 1793 2776 1823 2783
rect 1793 2773 1807 2776
rect 1816 2767 1823 2776
rect 1833 2733 1847 2747
rect 1836 2727 1843 2733
rect 1656 2556 1683 2563
rect 1596 2287 1603 2313
rect 1536 2256 1563 2263
rect 1476 1807 1483 1973
rect 1556 1943 1563 2256
rect 1573 2253 1587 2267
rect 1593 2273 1607 2287
rect 1613 2253 1627 2267
rect 1576 2247 1583 2253
rect 1616 2227 1623 2253
rect 1576 1947 1583 2113
rect 1536 1936 1563 1943
rect 1433 1793 1447 1807
rect 1436 1767 1443 1793
rect 1453 1773 1467 1787
rect 1473 1793 1487 1807
rect 1536 1787 1543 1936
rect 1596 1823 1603 2133
rect 1636 2067 1643 2353
rect 1656 2087 1663 2333
rect 1676 2087 1683 2556
rect 1713 2533 1727 2547
rect 1733 2553 1747 2567
rect 1716 2523 1723 2533
rect 1696 2516 1723 2523
rect 1696 2467 1703 2516
rect 1716 2347 1723 2493
rect 1747 2476 1753 2483
rect 1716 2287 1723 2293
rect 1736 2287 1743 2453
rect 1756 2287 1763 2353
rect 1753 2273 1767 2287
rect 1756 2227 1763 2233
rect 1613 2033 1627 2047
rect 1656 2063 1663 2073
rect 1656 2056 1673 2063
rect 1696 2047 1703 2093
rect 1616 2027 1623 2033
rect 1576 1816 1603 1823
rect 1576 1807 1583 1816
rect 1573 1793 1587 1807
rect 1613 1793 1627 1807
rect 1616 1787 1623 1793
rect 1593 1773 1607 1787
rect 1413 1603 1427 1607
rect 1396 1596 1427 1603
rect 1376 1427 1383 1593
rect 1396 1507 1403 1596
rect 1413 1593 1427 1596
rect 1436 1363 1443 1673
rect 1456 1627 1463 1773
rect 1453 1603 1467 1607
rect 1453 1596 1483 1603
rect 1453 1593 1467 1596
rect 1476 1567 1483 1596
rect 1416 1356 1443 1363
rect 1416 1347 1423 1356
rect 1413 1333 1427 1347
rect 1433 1313 1447 1327
rect 1436 1167 1443 1313
rect 1433 1143 1447 1147
rect 1433 1136 1463 1143
rect 1433 1133 1447 1136
rect 1376 1107 1383 1133
rect 1413 1093 1427 1107
rect 1416 1087 1423 1093
rect 1456 1087 1463 1136
rect 1333 863 1347 867
rect 1316 856 1347 863
rect 1253 633 1267 647
rect 1196 607 1203 613
rect 1316 587 1323 856
rect 1333 853 1347 856
rect 1393 843 1407 847
rect 1416 843 1423 853
rect 1393 836 1423 843
rect 1393 833 1407 836
rect 853 356 883 363
rect 853 353 867 356
rect 856 207 863 353
rect 953 353 967 367
rect 973 313 987 327
rect 976 307 983 313
rect 1016 227 1023 413
rect 1116 387 1123 533
rect 1036 283 1043 373
rect 1053 353 1067 367
rect 1113 373 1127 387
rect 1213 363 1227 367
rect 1196 356 1227 363
rect 1056 307 1063 353
rect 1196 287 1203 356
rect 1213 353 1227 356
rect 1236 323 1243 553
rect 1336 347 1343 733
rect 1373 613 1387 627
rect 1376 567 1383 613
rect 1416 587 1423 613
rect 1413 353 1427 367
rect 1416 347 1423 353
rect 1216 316 1243 323
rect 1036 276 1063 283
rect 856 147 863 193
rect 916 187 923 213
rect 913 173 927 187
rect 876 147 883 173
rect 196 107 203 133
rect 236 127 243 133
rect 793 113 807 127
rect 813 133 827 147
rect 853 133 867 147
rect 836 127 843 133
rect 896 127 903 173
rect 1016 167 1023 213
rect 1056 167 1063 276
rect 1013 153 1027 167
rect 933 133 947 147
rect 936 127 943 133
rect 956 127 963 153
rect 1033 133 1047 147
rect 1053 153 1067 167
rect 1076 147 1083 273
rect 1073 133 1087 147
rect 1136 143 1143 193
rect 1216 167 1223 316
rect 1273 313 1287 327
rect 1153 143 1167 147
rect 1136 136 1167 143
rect 1153 133 1167 136
rect 1213 153 1227 167
rect 1236 147 1243 173
rect 1276 167 1283 313
rect 1336 187 1343 333
rect 1436 203 1443 873
rect 1456 867 1463 1073
rect 1496 1067 1503 1733
rect 1516 1167 1523 1753
rect 1596 1687 1603 1773
rect 1636 1627 1643 1793
rect 1676 1607 1683 2013
rect 1716 1987 1723 2193
rect 1756 2103 1763 2213
rect 1776 2127 1783 2653
rect 1796 2567 1803 2693
rect 1796 2507 1803 2533
rect 1816 2487 1823 2553
rect 1836 2543 1843 2713
rect 1856 2607 1863 3293
rect 1916 3283 1923 3493
rect 1936 3467 1943 3493
rect 1976 3487 1983 3493
rect 1936 3307 1943 3453
rect 1896 3276 1923 3283
rect 1896 3207 1903 3276
rect 1953 3263 1967 3267
rect 1933 3233 1947 3247
rect 1953 3256 1983 3263
rect 1953 3253 1967 3256
rect 1936 3207 1943 3233
rect 1896 3047 1903 3153
rect 1936 3047 1943 3073
rect 1976 3067 1983 3256
rect 1893 3043 1907 3047
rect 1876 3036 1907 3043
rect 1876 3027 1883 3036
rect 1893 3033 1907 3036
rect 1933 3033 1947 3047
rect 1953 3023 1967 3027
rect 1953 3016 1983 3023
rect 1953 3013 1967 3016
rect 1976 2987 1983 3016
rect 1916 2667 1923 2853
rect 1936 2787 1943 2793
rect 1976 2787 1983 2933
rect 1996 2807 2003 3373
rect 2016 3287 2023 3493
rect 2036 3447 2043 3673
rect 2016 3047 2023 3273
rect 2056 3247 2063 3513
rect 2076 3307 2083 3793
rect 2096 3727 2103 4173
rect 2116 3707 2123 4173
rect 2136 4167 2143 4213
rect 2173 4213 2187 4227
rect 2196 4207 2203 4273
rect 2156 4047 2163 4193
rect 2176 3967 2183 4013
rect 2173 3953 2187 3967
rect 2136 3747 2143 3753
rect 2133 3733 2147 3747
rect 2153 3713 2167 3727
rect 2096 3683 2103 3693
rect 2096 3676 2123 3683
rect 2116 3527 2123 3676
rect 2156 3547 2163 3713
rect 2216 3627 2223 4313
rect 2236 4187 2243 4233
rect 2276 4223 2283 4553
rect 2333 4433 2347 4447
rect 2373 4443 2387 4447
rect 2396 4443 2403 4653
rect 2456 4587 2463 4953
rect 2536 4927 2543 5156
rect 2556 5147 2563 5193
rect 2596 5167 2603 5433
rect 2676 5427 2683 5433
rect 2673 5413 2687 5427
rect 2696 5363 2703 5633
rect 2736 5607 2743 5633
rect 2776 5567 2783 5633
rect 2776 5427 2783 5533
rect 2773 5413 2787 5427
rect 2796 5407 2803 5653
rect 2816 5567 2823 5656
rect 2833 5653 2847 5656
rect 2853 5633 2867 5647
rect 2816 5427 2823 5553
rect 2856 5467 2863 5633
rect 3093 5613 3107 5627
rect 3133 5613 3147 5627
rect 3413 5623 3427 5627
rect 3436 5623 3443 5653
rect 4096 5647 4103 5653
rect 3553 5633 3567 5647
rect 3753 5643 3767 5647
rect 2993 5593 3007 5607
rect 2996 5547 3003 5593
rect 2856 5427 2863 5453
rect 2876 5447 2883 5533
rect 2916 5447 2923 5453
rect 2873 5433 2887 5447
rect 2813 5413 2827 5427
rect 2913 5433 2927 5447
rect 2936 5427 2943 5473
rect 3096 5447 3103 5613
rect 3136 5607 3143 5613
rect 3413 5616 3443 5623
rect 3413 5613 3427 5616
rect 3396 5527 3403 5593
rect 3256 5427 3263 5453
rect 3436 5447 3443 5616
rect 3496 5463 3503 5613
rect 3513 5463 3527 5467
rect 3496 5456 3527 5463
rect 2933 5413 2947 5427
rect 3033 5413 3047 5427
rect 2793 5393 2807 5407
rect 3036 5407 3043 5413
rect 3253 5413 3267 5427
rect 3153 5393 3167 5407
rect 3156 5387 3163 5393
rect 2676 5356 2703 5363
rect 2593 5153 2607 5167
rect 2676 5127 2683 5356
rect 3013 5183 3027 5187
rect 2693 5153 2707 5167
rect 2556 4947 2563 5113
rect 2656 4987 2663 5053
rect 2696 5027 2703 5153
rect 2713 5133 2727 5147
rect 2753 5133 2767 5147
rect 2716 5127 2723 5133
rect 2756 4987 2763 5133
rect 2653 4973 2667 4987
rect 2776 4947 2783 4973
rect 2553 4943 2567 4947
rect 2553 4936 2583 4943
rect 2553 4933 2567 4936
rect 2576 4903 2583 4936
rect 2773 4933 2787 4947
rect 2793 4913 2807 4927
rect 2556 4896 2583 4903
rect 2536 4727 2543 4873
rect 2536 4707 2543 4713
rect 2533 4693 2547 4707
rect 2516 4607 2523 4673
rect 2476 4467 2483 4493
rect 2373 4436 2403 4443
rect 2373 4433 2387 4436
rect 2336 4427 2343 4433
rect 2336 4407 2343 4413
rect 2256 4216 2283 4223
rect 2256 4107 2263 4216
rect 2313 4173 2327 4187
rect 2316 4107 2323 4173
rect 2336 4167 2343 4353
rect 2356 4187 2363 4253
rect 2253 3983 2267 3987
rect 2247 3976 2267 3983
rect 2253 3973 2267 3976
rect 2236 3723 2243 3973
rect 2276 3967 2283 4013
rect 2376 4007 2383 4333
rect 2396 4227 2403 4436
rect 2416 4327 2423 4453
rect 2436 4307 2443 4453
rect 2453 4433 2467 4447
rect 2496 4447 2503 4513
rect 2556 4463 2563 4896
rect 2596 4867 2603 4913
rect 2796 4907 2803 4913
rect 2576 4667 2583 4693
rect 2596 4567 2603 4853
rect 2576 4467 2583 4513
rect 2616 4467 2623 4493
rect 2493 4433 2507 4447
rect 2536 4456 2563 4463
rect 2456 4347 2463 4433
rect 2456 4207 2463 4253
rect 2413 4193 2427 4207
rect 2416 4147 2423 4193
rect 2453 4193 2467 4207
rect 2473 4173 2487 4187
rect 2476 4167 2483 4173
rect 2296 3987 2303 3993
rect 2293 3973 2307 3987
rect 2273 3953 2287 3967
rect 2336 3767 2343 3993
rect 2396 3887 2403 4113
rect 2416 3987 2423 4093
rect 2496 4083 2503 4233
rect 2516 4127 2523 4253
rect 2496 4076 2523 4083
rect 2453 3973 2467 3987
rect 2496 3987 2503 4013
rect 2456 3927 2463 3973
rect 2516 3967 2523 4076
rect 2273 3733 2287 3747
rect 2276 3727 2283 3733
rect 2253 3723 2267 3727
rect 2236 3716 2267 3723
rect 2253 3713 2267 3716
rect 2293 3713 2307 3727
rect 2256 3667 2263 3713
rect 2256 3543 2263 3573
rect 2276 3567 2283 3713
rect 2296 3707 2303 3713
rect 2336 3703 2343 3753
rect 2316 3696 2343 3703
rect 2256 3536 2283 3543
rect 2113 3513 2127 3527
rect 2176 3507 2183 3533
rect 2033 3213 2047 3227
rect 2053 3233 2067 3247
rect 2036 3147 2043 3213
rect 2073 3203 2087 3207
rect 2073 3196 2103 3203
rect 2073 3193 2087 3196
rect 2036 2867 2043 3073
rect 2076 3027 2083 3053
rect 2096 3047 2103 3196
rect 2116 3087 2123 3393
rect 2196 3287 2203 3533
rect 2276 3527 2283 3536
rect 2233 3523 2247 3527
rect 2216 3516 2247 3523
rect 2216 3487 2223 3516
rect 2233 3513 2247 3516
rect 2273 3513 2287 3527
rect 2296 3507 2303 3513
rect 2293 3493 2307 3507
rect 2316 3483 2323 3696
rect 2336 3507 2343 3533
rect 2316 3476 2343 3483
rect 2153 3263 2167 3267
rect 2147 3256 2167 3263
rect 2153 3253 2167 3256
rect 2136 3107 2143 3253
rect 2093 3033 2107 3047
rect 2133 3043 2147 3047
rect 2073 3013 2087 3027
rect 2133 3036 2163 3043
rect 2133 3033 2147 3036
rect 2156 3007 2163 3036
rect 1933 2773 1947 2787
rect 1973 2773 1987 2787
rect 1996 2747 2003 2793
rect 2016 2743 2023 2773
rect 2056 2767 2063 2813
rect 2033 2743 2047 2747
rect 2016 2736 2047 2743
rect 2053 2753 2067 2767
rect 2093 2753 2107 2767
rect 2033 2733 2047 2736
rect 2073 2733 2087 2747
rect 1916 2567 1923 2613
rect 1853 2543 1867 2547
rect 1836 2536 1867 2543
rect 1836 2487 1843 2536
rect 1853 2533 1867 2536
rect 1893 2533 1907 2547
rect 1913 2553 1927 2567
rect 1896 2523 1903 2533
rect 1876 2516 1903 2523
rect 1796 2267 1803 2473
rect 1876 2467 1883 2516
rect 1816 2227 1823 2453
rect 1876 2447 1883 2453
rect 1836 2307 1843 2333
rect 1896 2323 1903 2473
rect 1896 2316 1923 2323
rect 1916 2307 1923 2316
rect 1833 2293 1847 2307
rect 1893 2283 1907 2287
rect 1893 2276 1923 2283
rect 1893 2273 1907 2276
rect 1736 2096 1763 2103
rect 1736 2087 1743 2096
rect 1776 2087 1783 2093
rect 1733 2073 1747 2087
rect 1753 2053 1767 2067
rect 1773 2073 1787 2087
rect 1793 2063 1807 2067
rect 1816 2063 1823 2193
rect 1793 2056 1823 2063
rect 1793 2053 1807 2056
rect 1756 2047 1763 2053
rect 1696 1803 1703 1853
rect 1756 1807 1763 1933
rect 1713 1803 1727 1807
rect 1696 1796 1727 1803
rect 1713 1793 1727 1796
rect 1716 1607 1723 1793
rect 1773 1773 1787 1787
rect 1736 1627 1743 1773
rect 1776 1767 1783 1773
rect 1816 1747 1823 2056
rect 1836 2027 1843 2173
rect 1876 2167 1883 2273
rect 1916 2267 1923 2276
rect 1896 2187 1903 2253
rect 1936 2127 1943 2593
rect 1836 1767 1843 1953
rect 1856 1867 1863 2113
rect 1893 1823 1907 1827
rect 1916 1823 1923 1913
rect 1873 1793 1887 1807
rect 1893 1816 1923 1823
rect 1893 1813 1907 1816
rect 1876 1727 1883 1793
rect 1556 1363 1563 1573
rect 1536 1356 1563 1363
rect 1536 1347 1543 1356
rect 1533 1333 1547 1347
rect 1573 1343 1587 1347
rect 1596 1343 1603 1593
rect 1673 1593 1687 1607
rect 1713 1603 1727 1607
rect 1693 1573 1707 1587
rect 1713 1596 1743 1603
rect 1713 1593 1727 1596
rect 1696 1387 1703 1573
rect 1736 1367 1743 1596
rect 1773 1573 1787 1587
rect 1776 1567 1783 1573
rect 1796 1523 1803 1673
rect 1776 1516 1803 1523
rect 1573 1336 1603 1343
rect 1573 1333 1587 1336
rect 1516 1127 1523 1153
rect 1513 1113 1527 1127
rect 1556 1127 1563 1173
rect 1553 1113 1567 1127
rect 1476 847 1483 853
rect 1473 833 1487 847
rect 1456 367 1463 693
rect 1536 687 1543 1093
rect 1596 887 1603 1336
rect 1733 1323 1747 1327
rect 1756 1323 1763 1373
rect 1733 1316 1763 1323
rect 1733 1313 1747 1316
rect 1596 867 1603 873
rect 1593 853 1607 867
rect 1616 807 1623 1173
rect 1636 1147 1643 1153
rect 1633 1133 1647 1147
rect 1776 1107 1783 1516
rect 1796 1347 1803 1373
rect 1836 1347 1843 1613
rect 1856 1587 1863 1693
rect 1916 1687 1923 1816
rect 1936 1747 1943 1873
rect 1956 1827 1963 2733
rect 1976 2567 1983 2573
rect 1973 2553 1987 2567
rect 1993 2533 2007 2547
rect 1996 2527 2003 2533
rect 1976 2307 1983 2373
rect 2056 2327 2063 2573
rect 1973 2293 1987 2307
rect 1993 2273 2007 2287
rect 2033 2273 2047 2287
rect 1996 2207 2003 2273
rect 2036 2267 2043 2273
rect 1976 1947 1983 2113
rect 1996 2087 2003 2193
rect 2056 2103 2063 2313
rect 2076 2303 2083 2733
rect 2096 2667 2103 2753
rect 2116 2547 2123 2813
rect 2136 2567 2143 2893
rect 2156 2747 2163 2993
rect 2176 2827 2183 3113
rect 2196 2967 2203 3213
rect 2216 3207 2223 3473
rect 2236 3227 2243 3253
rect 2236 3063 2243 3213
rect 2256 3127 2263 3273
rect 2276 3203 2283 3433
rect 2316 3267 2323 3293
rect 2313 3253 2327 3267
rect 2276 3196 2303 3203
rect 2216 3056 2243 3063
rect 2216 3027 2223 3056
rect 2213 3013 2227 3027
rect 2256 2943 2263 3013
rect 2256 2936 2283 2943
rect 2096 2427 2103 2533
rect 2133 2513 2147 2527
rect 2176 2527 2183 2793
rect 2196 2787 2203 2893
rect 2196 2547 2203 2593
rect 2193 2533 2207 2547
rect 2116 2347 2123 2513
rect 2136 2367 2143 2513
rect 2136 2323 2143 2353
rect 2156 2327 2163 2493
rect 2216 2467 2223 2733
rect 2236 2603 2243 2913
rect 2253 2733 2267 2747
rect 2256 2707 2263 2733
rect 2236 2596 2263 2603
rect 2236 2467 2243 2553
rect 2256 2487 2263 2596
rect 2276 2587 2283 2936
rect 2296 2727 2303 3196
rect 2316 2807 2323 3153
rect 2336 3147 2343 3476
rect 2356 3467 2363 3513
rect 2376 3507 2383 3813
rect 2396 3587 2403 3793
rect 2456 3727 2463 3873
rect 2476 3807 2483 3873
rect 2433 3693 2447 3707
rect 2436 3647 2443 3693
rect 2436 3547 2443 3573
rect 2433 3533 2447 3547
rect 2396 3527 2403 3533
rect 2393 3513 2407 3527
rect 2413 3493 2427 3507
rect 2353 3223 2367 3227
rect 2376 3223 2383 3493
rect 2416 3383 2423 3493
rect 2396 3376 2423 3383
rect 2396 3227 2403 3376
rect 2416 3267 2423 3293
rect 2456 3267 2463 3493
rect 2413 3253 2427 3267
rect 2433 3233 2447 3247
rect 2453 3253 2467 3267
rect 2353 3216 2383 3223
rect 2353 3213 2367 3216
rect 2356 3067 2363 3113
rect 2356 3027 2363 3053
rect 2376 3047 2383 3193
rect 2436 3127 2443 3233
rect 2476 3223 2483 3253
rect 2456 3216 2483 3223
rect 2373 3033 2387 3047
rect 2433 3013 2447 3027
rect 2333 2783 2347 2787
rect 2316 2776 2347 2783
rect 2316 2707 2323 2776
rect 2333 2773 2347 2776
rect 2387 2776 2403 2783
rect 2396 2727 2403 2776
rect 2416 2767 2423 3013
rect 2436 2927 2443 3013
rect 2316 2587 2323 2593
rect 2313 2573 2327 2587
rect 2276 2567 2283 2573
rect 2273 2553 2287 2567
rect 2293 2533 2307 2547
rect 2296 2527 2303 2533
rect 2336 2487 2343 2533
rect 2356 2527 2363 2573
rect 2116 2316 2143 2323
rect 2076 2296 2103 2303
rect 2096 2227 2103 2296
rect 2116 2267 2123 2316
rect 2056 2096 2083 2103
rect 2076 2067 2083 2096
rect 2076 2047 2083 2053
rect 1976 1827 1983 1873
rect 2016 1827 2023 1973
rect 1973 1813 1987 1827
rect 1993 1793 2007 1807
rect 2013 1813 2027 1827
rect 1996 1687 2003 1793
rect 1853 1573 1867 1587
rect 1917 1545 1925 1636
rect 1917 1506 1925 1531
rect 1935 1521 1943 1636
rect 1956 1545 1964 1636
rect 1989 1597 1997 1636
rect 1989 1524 1997 1583
rect 2017 1579 2025 1636
rect 2017 1524 2025 1565
rect 2036 1487 2043 1573
rect 1793 1333 1807 1347
rect 1813 1313 1827 1327
rect 1833 1333 1847 1347
rect 1653 1093 1667 1107
rect 1656 887 1663 1093
rect 1773 1093 1787 1107
rect 1796 1087 1803 1233
rect 1816 1127 1823 1313
rect 1813 1103 1827 1107
rect 1836 1103 1843 1133
rect 1813 1096 1843 1103
rect 1813 1093 1827 1096
rect 1793 1073 1807 1087
rect 1516 647 1523 653
rect 1493 623 1507 627
rect 1476 616 1507 623
rect 1476 567 1483 616
rect 1493 613 1507 616
rect 1516 607 1523 633
rect 1513 593 1527 607
rect 1476 347 1483 393
rect 1596 387 1603 613
rect 1636 427 1643 853
rect 1753 853 1767 867
rect 1733 833 1747 847
rect 1736 827 1743 833
rect 1756 787 1763 853
rect 1816 827 1823 993
rect 1836 847 1843 1096
rect 1856 1067 1863 1113
rect 1876 1087 1883 1333
rect 1993 1313 2007 1327
rect 1996 1287 2003 1313
rect 2016 1187 2023 1333
rect 2056 1327 2063 1933
rect 2116 1807 2123 1833
rect 2113 1793 2127 1807
rect 2075 1507 2083 1633
rect 2095 1549 2103 1633
rect 2095 1507 2103 1535
rect 2115 1507 2123 1633
rect 2136 1607 2143 2293
rect 2153 2273 2167 2287
rect 2156 2167 2163 2273
rect 2176 2247 2183 2373
rect 2217 2329 2225 2354
rect 2153 2083 2167 2087
rect 2176 2083 2183 2233
rect 2196 2087 2203 2313
rect 2217 2224 2225 2315
rect 2235 2224 2243 2339
rect 2256 2224 2264 2315
rect 2289 2277 2297 2336
rect 2317 2295 2325 2336
rect 2289 2224 2297 2263
rect 2317 2224 2325 2281
rect 2153 2076 2183 2083
rect 2153 2073 2167 2076
rect 2156 1807 2163 1813
rect 2196 1807 2203 1813
rect 2153 1793 2167 1807
rect 2193 1793 2207 1807
rect 2153 1583 2167 1587
rect 2136 1576 2167 1583
rect 2076 1327 2083 1373
rect 2073 1313 2087 1327
rect 2076 1127 2083 1173
rect 1893 1073 1907 1087
rect 2073 1113 2087 1127
rect 1896 1067 1903 1073
rect 1856 867 1863 873
rect 1853 853 1867 867
rect 1873 833 1887 847
rect 1876 827 1883 833
rect 1656 627 1663 653
rect 1696 387 1703 613
rect 1516 367 1523 373
rect 1656 367 1663 373
rect 1716 367 1723 593
rect 1513 353 1527 367
rect 1616 327 1623 353
rect 1633 333 1647 347
rect 1653 353 1667 367
rect 1736 347 1743 633
rect 1776 627 1783 793
rect 1956 747 1963 1073
rect 1993 853 2007 867
rect 1996 787 2003 853
rect 2013 833 2027 847
rect 2016 827 2023 833
rect 1816 687 1823 693
rect 1816 627 1823 673
rect 1856 627 1863 693
rect 1976 647 1983 753
rect 1996 747 2003 773
rect 1996 647 2003 653
rect 1793 593 1807 607
rect 1813 613 1827 627
rect 1973 633 1987 647
rect 1996 627 2003 633
rect 1796 587 1803 593
rect 1753 333 1767 347
rect 1636 307 1643 333
rect 1416 196 1443 203
rect 1336 167 1343 173
rect 1416 167 1423 196
rect 1596 187 1603 193
rect 1593 173 1607 187
rect 1333 153 1347 167
rect 1036 127 1043 133
rect 1436 123 1443 173
rect 1473 163 1487 167
rect 1473 156 1503 163
rect 1473 153 1487 156
rect 1496 127 1503 156
rect 1736 167 1743 173
rect 1733 153 1747 167
rect 1756 147 1763 333
rect 1453 123 1467 127
rect 1436 116 1467 123
rect 1453 113 1467 116
rect 1796 123 1803 153
rect 1836 147 1843 553
rect 1916 407 1923 613
rect 2056 607 2063 853
rect 2076 827 2083 1053
rect 2096 767 2103 1253
rect 2116 1107 2123 1473
rect 2136 1447 2143 1576
rect 2153 1573 2167 1576
rect 2136 907 2143 1373
rect 2176 1303 2183 1773
rect 2193 1563 2207 1567
rect 2216 1563 2223 1833
rect 2236 1807 2243 2153
rect 2276 2067 2283 2173
rect 2253 2033 2267 2047
rect 2273 2053 2287 2067
rect 2313 2063 2327 2067
rect 2336 2063 2343 2213
rect 2356 2203 2363 2513
rect 2376 2387 2383 2553
rect 2416 2547 2423 2593
rect 2436 2567 2443 2793
rect 2456 2787 2463 3216
rect 2476 3007 2483 3053
rect 2496 3003 2503 3953
rect 2516 3887 2523 3953
rect 2536 3887 2543 4456
rect 2573 4453 2587 4467
rect 2613 4453 2627 4467
rect 2633 4433 2647 4447
rect 2636 4387 2643 4433
rect 2656 4407 2663 4733
rect 2673 4653 2687 4667
rect 2676 4627 2683 4653
rect 2676 4607 2683 4613
rect 2573 4223 2587 4227
rect 2556 4216 2587 4223
rect 2556 4147 2563 4216
rect 2573 4213 2587 4216
rect 2613 4213 2627 4227
rect 2596 4187 2603 4193
rect 2596 4003 2603 4013
rect 2576 3996 2603 4003
rect 2576 3987 2583 3996
rect 2616 3987 2623 4213
rect 2676 4147 2683 4573
rect 2696 4307 2703 4693
rect 2733 4673 2747 4687
rect 2773 4673 2787 4687
rect 2816 4687 2823 5173
rect 3013 5176 3043 5183
rect 3013 5173 3027 5176
rect 2853 5153 2867 5167
rect 2836 4907 2843 5033
rect 2856 4987 2863 5153
rect 2913 5133 2927 5147
rect 3036 5147 3043 5176
rect 3053 5133 3067 5147
rect 2916 5127 2923 5133
rect 2976 4927 2983 4953
rect 2996 4947 3003 5013
rect 2993 4933 3007 4947
rect 2973 4913 2987 4927
rect 3013 4923 3027 4927
rect 3036 4923 3043 5093
rect 3056 5007 3063 5133
rect 3153 5133 3167 5147
rect 3156 5007 3163 5133
rect 3116 4947 3123 4993
rect 3176 4987 3183 5413
rect 3276 5407 3283 5433
rect 3273 5393 3287 5407
rect 3313 5393 3327 5407
rect 3273 5163 3287 5167
rect 3256 5156 3287 5163
rect 3173 4963 3187 4967
rect 3013 4916 3043 4923
rect 3113 4933 3127 4947
rect 3153 4933 3167 4947
rect 3173 4956 3203 4963
rect 3173 4953 3187 4956
rect 3156 4923 3163 4933
rect 3136 4916 3163 4923
rect 3013 4913 3027 4916
rect 2736 4667 2743 4673
rect 2776 4667 2783 4673
rect 2776 4647 2783 4653
rect 2756 4507 2763 4553
rect 2753 4493 2767 4507
rect 2716 4447 2723 4493
rect 2836 4487 2843 4553
rect 2876 4527 2883 4913
rect 3136 4847 3143 4916
rect 3176 4903 3183 4913
rect 3156 4896 3183 4903
rect 2893 4653 2907 4667
rect 2933 4663 2947 4667
rect 2956 4663 2963 4693
rect 3036 4687 3043 4693
rect 2896 4587 2903 4653
rect 2933 4656 2963 4663
rect 2933 4653 2947 4656
rect 3013 4653 3027 4667
rect 3033 4673 3047 4687
rect 3053 4653 3067 4667
rect 2913 4633 2927 4647
rect 2916 4627 2923 4633
rect 3016 4587 3023 4653
rect 3056 4643 3063 4653
rect 3036 4636 3063 4643
rect 2833 4483 2847 4487
rect 2816 4476 2847 4483
rect 2716 4227 2723 4253
rect 2693 4153 2707 4167
rect 2696 4127 2703 4153
rect 2636 3987 2643 3993
rect 2676 3987 2683 3993
rect 2573 3973 2587 3987
rect 2653 3963 2667 3967
rect 2647 3956 2667 3963
rect 2673 3973 2687 3987
rect 2653 3953 2667 3956
rect 2576 3747 2583 3753
rect 2533 3743 2547 3747
rect 2516 3736 2547 3743
rect 2516 3667 2523 3736
rect 2533 3733 2547 3736
rect 2573 3733 2587 3747
rect 2596 3687 2603 3933
rect 2616 3927 2623 3953
rect 2516 3127 2523 3633
rect 2596 3527 2603 3613
rect 2593 3513 2607 3527
rect 2556 3367 2563 3413
rect 2576 3287 2583 3513
rect 2616 3327 2623 3873
rect 2636 3667 2643 3953
rect 2656 3807 2663 3873
rect 2676 3727 2683 3913
rect 2716 3803 2723 4133
rect 2736 3827 2743 4353
rect 2756 4127 2763 4453
rect 2816 4243 2823 4476
rect 2833 4473 2847 4476
rect 2796 4236 2823 4243
rect 2776 3987 2783 4213
rect 2796 4203 2803 4236
rect 2813 4203 2827 4207
rect 2853 4203 2867 4207
rect 2796 4196 2827 4203
rect 2813 4193 2827 4196
rect 2836 4196 2867 4203
rect 2836 4107 2843 4196
rect 2853 4193 2867 4196
rect 2896 4167 2903 4233
rect 2916 4207 2923 4513
rect 2936 4347 2943 4453
rect 2953 4433 2967 4447
rect 2996 4447 3003 4473
rect 3016 4467 3023 4493
rect 3013 4453 3027 4467
rect 2956 4287 2963 4433
rect 3036 4367 3043 4636
rect 3116 4467 3123 4513
rect 3136 4507 3143 4713
rect 3156 4707 3163 4896
rect 3093 4433 3107 4447
rect 3113 4453 3127 4467
rect 3136 4447 3143 4493
rect 3156 4467 3163 4693
rect 3176 4667 3183 4873
rect 3196 4747 3203 4956
rect 3236 4727 3243 4973
rect 3256 4947 3263 5156
rect 3273 5153 3287 5156
rect 3276 4967 3283 5013
rect 3316 4987 3323 5393
rect 3336 5387 3343 5413
rect 3376 5403 3383 5433
rect 3393 5403 3407 5407
rect 3376 5396 3407 5403
rect 3393 5393 3407 5396
rect 3496 5267 3503 5456
rect 3513 5453 3527 5456
rect 3536 5447 3543 5473
rect 3556 5467 3563 5633
rect 3736 5636 3767 5643
rect 3556 5187 3563 5213
rect 3556 5167 3563 5173
rect 3373 5133 3387 5147
rect 3513 5153 3527 5167
rect 3376 5127 3383 5133
rect 3413 5133 3427 5147
rect 3393 5113 3407 5127
rect 3396 5023 3403 5113
rect 3376 5016 3403 5023
rect 3376 4967 3383 5016
rect 3416 5007 3423 5133
rect 3516 5127 3523 5153
rect 3533 5133 3547 5147
rect 3553 5153 3567 5167
rect 3573 5143 3587 5147
rect 3596 5143 3603 5433
rect 3573 5136 3603 5143
rect 3573 5133 3587 5136
rect 3396 4967 3403 4993
rect 3516 4987 3523 4993
rect 3536 4987 3543 5133
rect 3513 4973 3527 4987
rect 3273 4953 3287 4967
rect 3253 4933 3267 4947
rect 3293 4933 3307 4947
rect 3393 4953 3407 4967
rect 3376 4947 3383 4953
rect 3453 4933 3467 4947
rect 3296 4887 3303 4933
rect 3436 4907 3443 4933
rect 3236 4707 3243 4713
rect 3316 4707 3323 4853
rect 3213 4673 3227 4687
rect 3233 4693 3247 4707
rect 3313 4693 3327 4707
rect 3353 4693 3367 4707
rect 3153 4453 3167 4467
rect 3133 4433 3147 4447
rect 2996 4227 3003 4333
rect 2973 4193 2987 4207
rect 2993 4213 3007 4227
rect 2836 4087 2843 4093
rect 2816 4007 2823 4033
rect 2816 3987 2823 3993
rect 2756 3967 2763 3973
rect 2813 3973 2827 3987
rect 2833 3953 2847 3967
rect 2756 3943 2763 3953
rect 2756 3936 2783 3943
rect 2716 3796 2743 3803
rect 2696 3747 2703 3773
rect 2653 3693 2667 3707
rect 2693 3693 2707 3707
rect 2656 3643 2663 3693
rect 2696 3687 2703 3693
rect 2636 3636 2663 3643
rect 2553 3233 2567 3247
rect 2556 3187 2563 3233
rect 2613 3213 2627 3227
rect 2616 3167 2623 3213
rect 2516 3047 2523 3093
rect 2576 3067 2583 3113
rect 2513 3033 2527 3047
rect 2573 3013 2587 3027
rect 2496 2996 2523 3003
rect 2493 2733 2507 2747
rect 2473 2713 2487 2727
rect 2413 2533 2427 2547
rect 2456 2507 2463 2713
rect 2476 2707 2483 2713
rect 2496 2707 2503 2733
rect 2476 2527 2483 2693
rect 2496 2547 2503 2693
rect 2516 2627 2523 2996
rect 2536 2603 2543 2993
rect 2576 2827 2583 3013
rect 2596 3007 2603 3133
rect 2636 3107 2643 3636
rect 2716 3487 2723 3693
rect 2736 3647 2743 3796
rect 2736 3507 2743 3613
rect 2656 3367 2663 3473
rect 2756 3347 2763 3853
rect 2656 3207 2663 3273
rect 2636 3087 2643 3093
rect 2656 3047 2663 3173
rect 2676 3087 2683 3293
rect 2716 3247 2723 3253
rect 2756 3247 2763 3313
rect 2776 3287 2783 3936
rect 2796 3687 2803 3733
rect 2816 3727 2823 3793
rect 2836 3767 2843 3953
rect 2836 3727 2843 3753
rect 2813 3713 2827 3727
rect 2856 3527 2863 4133
rect 2876 4047 2883 4153
rect 2876 3947 2883 4013
rect 2916 4003 2923 4193
rect 2896 3996 2923 4003
rect 2896 3843 2903 3996
rect 2956 3987 2963 4113
rect 2976 4067 2983 4193
rect 3016 4043 3023 4233
rect 3036 4187 3043 4333
rect 3073 4203 3087 4207
rect 3056 4196 3087 4203
rect 3096 4203 3103 4433
rect 3113 4203 3127 4207
rect 3096 4196 3127 4203
rect 3056 4107 3063 4196
rect 3073 4193 3087 4196
rect 3113 4193 3127 4196
rect 3133 4173 3147 4187
rect 3093 4163 3107 4167
rect 3093 4156 3113 4163
rect 3093 4153 3107 4156
rect 2996 4036 3023 4043
rect 2996 4027 3003 4036
rect 3076 4023 3083 4113
rect 3056 4016 3083 4023
rect 2956 3887 2963 3933
rect 2996 3927 3003 3973
rect 3036 3967 3043 4013
rect 3056 3947 3063 4016
rect 3073 3973 3087 3987
rect 2876 3836 2903 3843
rect 2876 3527 2883 3836
rect 2956 3727 2963 3793
rect 2953 3713 2967 3727
rect 2996 3707 3003 3893
rect 2973 3693 2987 3707
rect 2976 3687 2983 3693
rect 2833 3493 2847 3507
rect 2853 3513 2867 3527
rect 2836 3487 2843 3493
rect 2856 3387 2863 3473
rect 2796 3263 2803 3333
rect 2876 3307 2883 3493
rect 2776 3256 2803 3263
rect 2876 3267 2883 3293
rect 2713 3233 2727 3247
rect 2776 3203 2783 3256
rect 2833 3253 2847 3267
rect 2836 3247 2843 3253
rect 2853 3233 2867 3247
rect 2873 3253 2887 3267
rect 2796 3227 2803 3233
rect 2776 3196 2803 3203
rect 2696 3047 2703 3113
rect 2673 3013 2687 3027
rect 2693 3033 2707 3047
rect 2713 3013 2727 3027
rect 2676 3007 2683 3013
rect 2576 2743 2583 2813
rect 2596 2787 2603 2913
rect 2676 2787 2683 2993
rect 2593 2773 2607 2787
rect 2613 2753 2627 2767
rect 2616 2743 2623 2753
rect 2576 2736 2623 2743
rect 2636 2623 2643 2773
rect 2696 2747 2703 2993
rect 2716 2987 2723 3013
rect 2616 2616 2643 2623
rect 2616 2607 2623 2616
rect 2516 2596 2543 2603
rect 2375 2227 2383 2353
rect 2395 2325 2403 2353
rect 2395 2227 2403 2311
rect 2415 2227 2423 2353
rect 2436 2263 2443 2493
rect 2496 2487 2503 2513
rect 2516 2367 2523 2596
rect 2556 2547 2563 2573
rect 2576 2567 2583 2593
rect 2573 2553 2587 2567
rect 2553 2533 2567 2547
rect 2596 2487 2603 2533
rect 2493 2303 2507 2307
rect 2476 2296 2507 2303
rect 2436 2256 2463 2263
rect 2356 2196 2383 2203
rect 2313 2056 2343 2063
rect 2313 2053 2327 2056
rect 2256 1967 2263 2033
rect 2236 1707 2243 1793
rect 2256 1663 2263 1813
rect 2296 1763 2303 1993
rect 2336 1947 2343 2056
rect 2353 2053 2367 2067
rect 2356 2027 2363 2053
rect 2376 2007 2383 2196
rect 2416 1907 2423 2093
rect 2436 2067 2443 2153
rect 2433 2053 2447 2067
rect 2456 1963 2463 2256
rect 2476 2067 2483 2296
rect 2493 2293 2507 2296
rect 2516 2187 2523 2353
rect 2536 2287 2543 2393
rect 2556 2187 2563 2413
rect 2636 2403 2643 2593
rect 2616 2396 2643 2403
rect 2593 2253 2607 2267
rect 2596 2227 2603 2253
rect 2616 2243 2623 2396
rect 2656 2307 2663 2713
rect 2696 2583 2703 2733
rect 2716 2587 2723 2953
rect 2756 2807 2763 3113
rect 2776 3047 2783 3073
rect 2796 3003 2803 3196
rect 2813 3023 2827 3027
rect 2836 3023 2843 3213
rect 2856 3207 2863 3233
rect 2856 3176 2873 3183
rect 2856 3147 2863 3176
rect 2876 3067 2883 3073
rect 2873 3053 2887 3067
rect 2813 3016 2843 3023
rect 2813 3013 2827 3016
rect 2796 2996 2823 3003
rect 2733 2733 2747 2747
rect 2776 2743 2783 2853
rect 2793 2743 2807 2747
rect 2776 2736 2807 2743
rect 2793 2733 2807 2736
rect 2736 2707 2743 2733
rect 2816 2723 2823 2996
rect 2836 2767 2843 2793
rect 2796 2716 2823 2723
rect 2676 2576 2703 2583
rect 2676 2567 2683 2576
rect 2693 2533 2707 2547
rect 2733 2543 2747 2547
rect 2733 2536 2763 2543
rect 2733 2533 2747 2536
rect 2696 2487 2703 2533
rect 2716 2303 2723 2513
rect 2756 2507 2763 2536
rect 2776 2447 2783 2573
rect 2796 2307 2803 2716
rect 2816 2607 2823 2693
rect 2836 2583 2843 2733
rect 2816 2576 2843 2583
rect 2856 2583 2863 2873
rect 2876 2867 2883 3013
rect 2896 2967 2903 3573
rect 2936 3523 2943 3653
rect 2996 3527 3003 3533
rect 2953 3523 2967 3527
rect 2936 3516 2967 3523
rect 2916 3387 2923 3413
rect 2916 3247 2923 3293
rect 2936 3267 2943 3516
rect 2953 3513 2967 3516
rect 2993 3513 3007 3527
rect 3016 3467 3023 3893
rect 3076 3767 3083 3973
rect 3116 3847 3123 4153
rect 3136 4127 3143 4173
rect 3156 4127 3163 4373
rect 3136 3847 3143 4033
rect 3053 3713 3067 3727
rect 3036 3547 3043 3693
rect 3056 3547 3063 3713
rect 3116 3707 3123 3793
rect 3076 3607 3083 3653
rect 3036 3327 3043 3533
rect 3056 3507 3063 3513
rect 3096 3507 3103 3593
rect 3056 3483 3063 3493
rect 3073 3483 3087 3487
rect 3056 3476 3087 3483
rect 3093 3493 3107 3507
rect 3073 3473 3087 3476
rect 3113 3473 3127 3487
rect 3116 3467 3123 3473
rect 2936 3243 2943 3253
rect 2973 3253 2987 3267
rect 3013 3263 3027 3267
rect 2953 3243 2967 3247
rect 2936 3236 2967 3243
rect 2953 3233 2967 3236
rect 2976 3227 2983 3253
rect 2993 3233 3007 3247
rect 3013 3256 3043 3263
rect 3013 3253 3027 3256
rect 2936 3187 2943 3213
rect 2996 3203 3003 3233
rect 2976 3196 3003 3203
rect 2896 2767 2903 2873
rect 2916 2807 2923 3173
rect 2936 3047 2943 3073
rect 2976 3067 2983 3196
rect 2933 3033 2947 3047
rect 2987 3036 3003 3043
rect 2873 2733 2887 2747
rect 2893 2753 2907 2767
rect 2933 2763 2947 2767
rect 2956 2763 2963 2833
rect 2933 2756 2963 2763
rect 2933 2753 2947 2756
rect 2876 2727 2883 2733
rect 2873 2583 2887 2587
rect 2856 2576 2887 2583
rect 2816 2547 2823 2576
rect 2873 2573 2887 2576
rect 2893 2543 2907 2547
rect 2916 2543 2923 2713
rect 2936 2547 2943 2673
rect 2893 2536 2923 2543
rect 2893 2533 2907 2536
rect 2716 2296 2743 2303
rect 2736 2287 2743 2296
rect 2713 2253 2727 2267
rect 2733 2273 2747 2287
rect 2753 2253 2767 2267
rect 2716 2247 2723 2253
rect 2616 2236 2643 2243
rect 2497 2025 2505 2116
rect 2497 1986 2505 2011
rect 2515 2001 2523 2116
rect 2536 2025 2544 2116
rect 2569 2077 2577 2116
rect 2569 2004 2577 2063
rect 2597 2059 2605 2116
rect 2616 2107 2623 2113
rect 2613 2093 2627 2107
rect 2597 2004 2605 2045
rect 2616 1967 2623 2053
rect 2456 1956 2483 1963
rect 2337 1849 2345 1874
rect 2193 1556 2223 1563
rect 2236 1656 2263 1663
rect 2276 1756 2303 1763
rect 2193 1553 2207 1556
rect 2236 1387 2243 1656
rect 2256 1587 2263 1633
rect 2213 1313 2227 1327
rect 2216 1307 2223 1313
rect 2176 1296 2203 1303
rect 2176 1107 2183 1113
rect 2173 1093 2187 1107
rect 2196 1087 2203 1296
rect 2256 1147 2263 1313
rect 2276 1267 2283 1756
rect 2337 1744 2345 1835
rect 2355 1744 2363 1859
rect 2376 1744 2384 1835
rect 2409 1797 2417 1856
rect 2437 1815 2445 1856
rect 2409 1744 2417 1783
rect 2437 1744 2445 1801
rect 2476 1707 2483 1956
rect 2495 1747 2503 1873
rect 2515 1845 2523 1873
rect 2515 1747 2523 1831
rect 2535 1747 2543 1873
rect 2556 1767 2563 1893
rect 2336 1607 2343 1613
rect 2333 1593 2347 1607
rect 2396 1543 2403 1693
rect 2416 1563 2423 1593
rect 2433 1563 2447 1567
rect 2416 1556 2447 1563
rect 2473 1563 2487 1567
rect 2496 1563 2503 1633
rect 2433 1553 2447 1556
rect 2473 1556 2503 1563
rect 2473 1553 2487 1556
rect 2436 1547 2443 1553
rect 2396 1536 2423 1543
rect 2296 1347 2303 1433
rect 2333 1343 2347 1347
rect 2316 1336 2347 1343
rect 2316 1287 2323 1336
rect 2333 1333 2347 1336
rect 2353 1313 2367 1327
rect 2356 1307 2363 1313
rect 2216 1107 2223 1133
rect 2316 1127 2323 1193
rect 2316 1107 2323 1113
rect 2336 1107 2343 1273
rect 2356 1267 2363 1293
rect 2376 1247 2383 1333
rect 2213 1093 2227 1107
rect 2136 847 2143 853
rect 2113 813 2127 827
rect 2133 833 2147 847
rect 2173 833 2187 847
rect 2116 807 2123 813
rect 2176 687 2183 833
rect 2116 647 2123 653
rect 2113 633 2127 647
rect 2176 623 2183 673
rect 2193 623 2207 627
rect 2176 616 2207 623
rect 2193 613 2207 616
rect 1856 343 1863 373
rect 1873 343 1887 347
rect 1856 336 1887 343
rect 1873 333 1887 336
rect 1893 313 1907 327
rect 1996 323 2003 373
rect 2013 323 2027 327
rect 1996 316 2027 323
rect 2013 313 2027 316
rect 1896 187 1903 313
rect 1916 147 1923 153
rect 1813 123 1827 127
rect 1796 116 1827 123
rect 1833 133 1847 147
rect 1813 113 1827 116
rect 1853 113 1867 127
rect 1913 133 1927 147
rect 2076 127 2083 493
rect 2176 367 2183 573
rect 2216 383 2223 893
rect 2236 823 2243 913
rect 2276 887 2283 1093
rect 2293 1073 2307 1087
rect 2313 1093 2327 1107
rect 2336 1087 2343 1093
rect 2333 1073 2347 1087
rect 2296 927 2303 1073
rect 2296 867 2303 893
rect 2293 863 2307 867
rect 2276 856 2307 863
rect 2253 823 2267 827
rect 2236 816 2267 823
rect 2253 813 2267 816
rect 2256 667 2263 813
rect 2276 647 2283 856
rect 2293 853 2307 856
rect 2313 813 2327 827
rect 2316 807 2323 813
rect 2376 707 2383 1113
rect 2396 1107 2403 1313
rect 2416 1063 2423 1536
rect 2516 1543 2523 1673
rect 2496 1536 2523 1543
rect 2473 1323 2487 1327
rect 2496 1323 2503 1536
rect 2536 1483 2543 1613
rect 2576 1587 2583 1733
rect 2596 1727 2603 1933
rect 2616 1847 2623 1953
rect 2616 1827 2623 1833
rect 2613 1813 2627 1827
rect 2636 1787 2643 2236
rect 2655 1987 2663 2113
rect 2675 2029 2683 2113
rect 2675 1987 2683 2015
rect 2695 1987 2703 2113
rect 2716 1947 2723 2213
rect 2756 2107 2763 2253
rect 2776 2207 2783 2253
rect 2733 2063 2747 2067
rect 2733 2056 2763 2063
rect 2733 2053 2747 2056
rect 2756 1923 2763 2056
rect 2773 2033 2787 2047
rect 2776 1967 2783 2033
rect 2756 1916 2773 1923
rect 2656 1807 2663 1913
rect 2696 1827 2703 1893
rect 2796 1887 2803 2293
rect 2816 1887 2823 2513
rect 2836 2287 2843 2393
rect 2876 2287 2883 2533
rect 2853 2253 2867 2267
rect 2873 2273 2887 2287
rect 2913 2273 2927 2287
rect 2856 2227 2863 2253
rect 2916 2247 2923 2273
rect 2856 2087 2863 2093
rect 2896 2087 2903 2113
rect 2916 2107 2923 2233
rect 2853 2083 2867 2087
rect 2836 2076 2867 2083
rect 2836 2027 2843 2076
rect 2853 2073 2867 2076
rect 2893 2073 2907 2087
rect 2693 1823 2707 1827
rect 2676 1816 2707 1823
rect 2733 1823 2747 1827
rect 2756 1823 2763 1833
rect 2633 1603 2647 1607
rect 2573 1573 2587 1587
rect 2613 1573 2627 1587
rect 2633 1596 2663 1603
rect 2633 1593 2647 1596
rect 2473 1316 2503 1323
rect 2473 1313 2487 1316
rect 2496 1187 2503 1316
rect 2516 1476 2543 1483
rect 2516 1243 2523 1476
rect 2536 1287 2543 1453
rect 2556 1307 2563 1393
rect 2596 1363 2603 1413
rect 2616 1407 2623 1573
rect 2656 1527 2663 1596
rect 2576 1356 2603 1363
rect 2576 1323 2583 1356
rect 2636 1327 2643 1353
rect 2676 1327 2683 1816
rect 2693 1813 2707 1816
rect 2713 1793 2727 1807
rect 2733 1816 2763 1823
rect 2733 1813 2747 1816
rect 2593 1323 2607 1327
rect 2576 1316 2607 1323
rect 2593 1313 2607 1316
rect 2633 1313 2647 1327
rect 2653 1293 2667 1307
rect 2516 1236 2543 1243
rect 2436 1107 2443 1133
rect 2496 1127 2503 1173
rect 2433 1093 2447 1107
rect 2493 1113 2507 1127
rect 2416 1056 2443 1063
rect 2416 847 2423 1033
rect 2413 833 2427 847
rect 2436 827 2443 1056
rect 2516 1047 2523 1213
rect 2536 1107 2543 1236
rect 2556 1083 2563 1133
rect 2596 1107 2603 1113
rect 2573 1083 2587 1087
rect 2556 1076 2587 1083
rect 2593 1093 2607 1107
rect 2556 907 2563 1076
rect 2573 1073 2587 1076
rect 2553 863 2567 867
rect 2533 833 2547 847
rect 2553 856 2583 863
rect 2553 853 2567 856
rect 2576 847 2583 856
rect 2636 847 2643 853
rect 2633 833 2647 847
rect 2393 793 2407 807
rect 2313 643 2327 647
rect 2296 636 2327 643
rect 2296 507 2303 636
rect 2313 633 2327 636
rect 2373 643 2387 647
rect 2396 643 2403 793
rect 2373 636 2403 643
rect 2373 633 2387 636
rect 2436 603 2443 753
rect 2453 603 2467 607
rect 2436 596 2467 603
rect 2453 593 2467 596
rect 2493 593 2507 607
rect 2216 376 2243 383
rect 2153 333 2167 347
rect 2173 353 2187 367
rect 2193 343 2207 347
rect 2216 343 2223 353
rect 2193 336 2223 343
rect 2193 333 2207 336
rect 2156 167 2163 333
rect 2176 187 2183 193
rect 2116 147 2123 153
rect 2093 113 2107 127
rect 2113 133 2127 147
rect 2153 143 2167 147
rect 2176 143 2183 173
rect 2153 136 2183 143
rect 2213 163 2227 167
rect 2236 163 2243 376
rect 2256 187 2263 413
rect 2336 367 2343 533
rect 2333 353 2347 367
rect 2356 327 2363 393
rect 2456 347 2463 593
rect 2496 567 2503 593
rect 2536 427 2543 833
rect 2656 767 2663 1293
rect 2676 1107 2683 1313
rect 2696 1207 2703 1753
rect 2716 1747 2723 1793
rect 2756 1767 2763 1816
rect 2716 1627 2723 1733
rect 2776 1607 2783 1813
rect 2796 1807 2803 1873
rect 2816 1767 2823 1853
rect 2893 1793 2907 1807
rect 2896 1787 2903 1793
rect 2916 1747 2923 1993
rect 2753 1553 2767 1567
rect 2756 1547 2763 1553
rect 2796 1547 2803 1613
rect 2736 1327 2743 1413
rect 2756 1336 2803 1343
rect 2756 1327 2763 1336
rect 2753 1313 2767 1327
rect 2733 1273 2747 1287
rect 2716 1187 2723 1273
rect 2736 1227 2743 1273
rect 2716 1147 2723 1173
rect 2713 1133 2727 1147
rect 2756 1127 2763 1193
rect 2756 867 2763 1113
rect 2776 1107 2783 1273
rect 2796 1227 2803 1336
rect 2816 1307 2823 1713
rect 2856 1607 2863 1633
rect 2896 1607 2903 1653
rect 2853 1593 2867 1607
rect 2836 1587 2843 1593
rect 2833 1573 2847 1587
rect 2873 1573 2887 1587
rect 2893 1593 2907 1607
rect 2836 1307 2843 1393
rect 2856 1387 2863 1513
rect 2876 1407 2883 1573
rect 2916 1547 2923 1713
rect 2936 1427 2943 2213
rect 2956 2127 2963 2756
rect 2976 2607 2983 2913
rect 2996 2787 3003 3036
rect 2996 2607 3003 2713
rect 2996 2587 3003 2593
rect 2993 2573 3007 2587
rect 3016 2543 3023 3213
rect 3036 3207 3043 3256
rect 3056 3227 3063 3453
rect 3036 2827 3043 3113
rect 3076 3047 3083 3273
rect 3096 3187 3103 3393
rect 3136 3347 3143 3673
rect 3156 3407 3163 4053
rect 3176 4027 3183 4633
rect 3216 4567 3223 4673
rect 3256 4647 3263 4673
rect 3356 4627 3363 4693
rect 3373 4683 3387 4687
rect 3396 4683 3403 4773
rect 3416 4687 3423 4713
rect 3373 4676 3403 4683
rect 3373 4673 3387 4676
rect 3216 4547 3223 4553
rect 3233 4453 3247 4467
rect 3236 4207 3243 4453
rect 3256 4207 3263 4533
rect 3213 4203 3227 4207
rect 3196 4196 3227 4203
rect 3196 4107 3203 4196
rect 3213 4193 3227 4196
rect 3253 4193 3267 4207
rect 3216 4083 3223 4113
rect 3196 4076 3223 4083
rect 3196 3987 3203 4076
rect 3173 3953 3187 3967
rect 3193 3973 3207 3987
rect 3216 3967 3223 4053
rect 3236 3987 3243 4113
rect 3276 4003 3283 4093
rect 3296 4047 3303 4593
rect 3316 4487 3323 4493
rect 3313 4473 3327 4487
rect 3333 4453 3347 4467
rect 3376 4467 3383 4473
rect 3373 4453 3387 4467
rect 3336 4447 3343 4453
rect 3316 4103 3323 4273
rect 3336 4167 3343 4393
rect 3393 4173 3407 4187
rect 3316 4096 3343 4103
rect 3336 4087 3343 4096
rect 3316 4027 3323 4073
rect 3336 4027 3343 4053
rect 3333 4013 3347 4027
rect 3276 3996 3303 4003
rect 3233 3973 3247 3987
rect 3213 3953 3227 3967
rect 3256 3967 3263 3993
rect 3176 3587 3183 3953
rect 3236 3847 3243 3873
rect 3196 3747 3203 3753
rect 3193 3733 3207 3747
rect 3256 3647 3263 3833
rect 3276 3663 3283 3973
rect 3296 3827 3303 3996
rect 3296 3687 3303 3753
rect 3316 3727 3323 3733
rect 3336 3727 3343 3813
rect 3356 3807 3363 4033
rect 3376 3847 3383 4153
rect 3396 4107 3403 4173
rect 3436 4107 3443 4793
rect 3456 4767 3463 4933
rect 3476 4707 3483 4753
rect 3476 4687 3483 4693
rect 3496 4687 3503 4973
rect 3533 4963 3547 4967
rect 3556 4963 3563 5113
rect 3533 4956 3563 4963
rect 3533 4953 3547 4956
rect 3516 4687 3523 4913
rect 3556 4867 3563 4956
rect 3573 4933 3587 4947
rect 3576 4927 3583 4933
rect 3616 4907 3623 5573
rect 3736 5547 3743 5636
rect 3753 5633 3767 5636
rect 3773 5593 3787 5607
rect 3933 5613 3947 5627
rect 3993 5633 4007 5647
rect 4093 5633 4107 5647
rect 3973 5613 3987 5627
rect 3936 5607 3943 5613
rect 3833 5593 3847 5607
rect 3947 5596 3963 5603
rect 3776 5587 3783 5593
rect 3716 5427 3723 5533
rect 3736 5447 3743 5533
rect 3636 5187 3643 5193
rect 3633 5173 3647 5187
rect 3673 5183 3687 5187
rect 3653 5153 3667 5167
rect 3673 5176 3693 5183
rect 3673 5173 3687 5176
rect 3656 5147 3663 5153
rect 3696 4987 3703 5173
rect 3693 4973 3707 4987
rect 3673 4963 3687 4967
rect 3656 4956 3687 4963
rect 3716 4967 3723 5093
rect 3453 4653 3467 4667
rect 3473 4673 3487 4687
rect 3513 4683 3527 4687
rect 3513 4676 3543 4683
rect 3513 4673 3527 4676
rect 3456 4647 3463 4653
rect 3536 4667 3543 4676
rect 3456 4207 3463 4513
rect 3476 4487 3483 4513
rect 3473 4473 3487 4487
rect 3493 4443 3507 4447
rect 3516 4443 3523 4493
rect 3493 4436 3523 4443
rect 3493 4433 3507 4436
rect 3516 4407 3523 4436
rect 3396 3787 3403 4073
rect 3476 4007 3483 4153
rect 3496 4127 3503 4193
rect 3556 4167 3563 4453
rect 3576 4247 3583 4893
rect 3656 4747 3663 4956
rect 3673 4953 3687 4956
rect 3713 4953 3727 4967
rect 3596 4707 3603 4713
rect 3593 4693 3607 4707
rect 3633 4693 3647 4707
rect 3636 4687 3643 4693
rect 3613 4673 3627 4687
rect 3616 4667 3623 4673
rect 3636 4647 3643 4673
rect 3656 4527 3663 4593
rect 3596 4447 3603 4473
rect 3636 4467 3643 4473
rect 3613 4433 3627 4447
rect 3633 4453 3647 4467
rect 3616 4407 3623 4433
rect 3636 4387 3643 4413
rect 3453 3973 3467 3987
rect 3473 3993 3487 4007
rect 3456 3947 3463 3973
rect 3496 3963 3503 4093
rect 3556 3987 3563 4053
rect 3576 4047 3583 4233
rect 3596 4203 3603 4253
rect 3676 4227 3683 4853
rect 3696 4487 3703 4813
rect 3716 4663 3723 4873
rect 3756 4707 3763 5493
rect 3776 5387 3783 5493
rect 3796 5427 3803 5513
rect 3836 5467 3843 5593
rect 3956 5527 3963 5596
rect 3976 5567 3983 5613
rect 3996 5607 4003 5633
rect 4153 5623 4167 5627
rect 4136 5616 4167 5623
rect 3976 5507 3983 5533
rect 3856 5467 3863 5493
rect 3853 5453 3867 5467
rect 3873 5423 3887 5427
rect 3896 5423 3903 5433
rect 3873 5416 3903 5423
rect 3873 5413 3887 5416
rect 3813 5183 3827 5187
rect 3813 5176 3843 5183
rect 3813 5173 3827 5176
rect 3836 5047 3843 5176
rect 3836 5007 3843 5033
rect 3856 5003 3863 5413
rect 3876 5407 3883 5413
rect 3916 5403 3923 5473
rect 3956 5427 3963 5493
rect 3933 5403 3947 5407
rect 3916 5396 3947 5403
rect 3953 5413 3967 5427
rect 3933 5393 3947 5396
rect 3973 5393 3987 5407
rect 3896 5167 3903 5393
rect 3976 5267 3983 5393
rect 3996 5387 4003 5593
rect 4136 5587 4143 5616
rect 4153 5613 4167 5616
rect 4177 5584 4185 5664
rect 4233 5613 4247 5627
rect 4236 5607 4243 5613
rect 4316 5584 4324 5696
rect 4716 5667 4723 5823
rect 5196 5816 5223 5823
rect 4736 5647 4743 5653
rect 4836 5647 4843 5673
rect 4593 5643 4607 5647
rect 4576 5636 4607 5643
rect 4513 5613 4527 5627
rect 4516 5567 4523 5613
rect 4133 5443 4147 5447
rect 4073 5423 4087 5427
rect 4056 5416 4087 5423
rect 4056 5367 4063 5416
rect 4073 5413 4087 5416
rect 4133 5436 4153 5443
rect 4133 5433 4147 5436
rect 4156 5407 4163 5433
rect 4213 5393 4227 5407
rect 4316 5403 4323 5453
rect 4333 5403 4347 5407
rect 4316 5396 4347 5403
rect 4376 5407 4383 5453
rect 4393 5423 4407 5427
rect 4393 5416 4423 5423
rect 4393 5413 4407 5416
rect 4333 5393 4347 5396
rect 4416 5407 4423 5416
rect 3956 5187 3963 5193
rect 3933 5153 3947 5167
rect 3953 5173 3967 5187
rect 3856 4996 3883 5003
rect 3776 4923 3783 4993
rect 3856 4947 3863 4973
rect 3793 4923 3807 4927
rect 3776 4916 3807 4923
rect 3853 4933 3867 4947
rect 3793 4913 3807 4916
rect 3796 4807 3803 4913
rect 3876 4827 3883 4996
rect 3916 4943 3923 5093
rect 3936 5067 3943 5153
rect 3933 4943 3947 4947
rect 3916 4936 3947 4943
rect 3933 4933 3947 4936
rect 3796 4687 3803 4693
rect 3733 4663 3747 4667
rect 3716 4656 3747 4663
rect 3793 4673 3807 4687
rect 3733 4653 3747 4656
rect 3816 4647 3823 4713
rect 3916 4707 3923 4773
rect 3773 4633 3787 4647
rect 3696 4447 3703 4473
rect 3633 4213 3647 4227
rect 3613 4203 3627 4207
rect 3596 4196 3627 4203
rect 3613 4193 3627 4196
rect 3636 4187 3643 4213
rect 3653 4193 3667 4207
rect 3476 3956 3503 3963
rect 3356 3747 3363 3773
rect 3313 3713 3327 3727
rect 3276 3656 3303 3663
rect 3196 3487 3203 3513
rect 3256 3467 3263 3493
rect 3276 3443 3283 3633
rect 3256 3436 3283 3443
rect 3116 3267 3123 3333
rect 3156 3283 3163 3313
rect 3156 3276 3183 3283
rect 3113 3253 3127 3267
rect 3133 3233 3147 3247
rect 3136 3167 3143 3233
rect 3096 3027 3103 3153
rect 3093 3013 3107 3027
rect 3113 2993 3127 3007
rect 3116 2987 3123 2993
rect 3136 2927 3143 3033
rect 3156 3023 3163 3073
rect 3116 2787 3123 2813
rect 3053 2753 3067 2767
rect 3093 2753 3107 2767
rect 3036 2547 3043 2733
rect 3056 2687 3063 2753
rect 3096 2747 3103 2753
rect 3136 2747 3143 2873
rect 3176 2807 3183 3276
rect 3196 3167 3203 3333
rect 3236 3267 3243 3333
rect 3256 3267 3263 3436
rect 3296 3347 3303 3656
rect 3316 3407 3323 3573
rect 3376 3503 3383 3753
rect 3393 3713 3407 3727
rect 3396 3587 3403 3713
rect 3396 3527 3403 3533
rect 3393 3503 3407 3507
rect 3376 3496 3407 3503
rect 3393 3493 3407 3496
rect 3416 3467 3423 3533
rect 3476 3523 3483 3956
rect 3553 3973 3567 3987
rect 3496 3547 3503 3913
rect 3516 3547 3523 3813
rect 3556 3727 3563 3753
rect 3553 3713 3567 3727
rect 3533 3673 3547 3687
rect 3536 3587 3543 3673
rect 3536 3527 3543 3573
rect 3556 3567 3563 3673
rect 3493 3523 3507 3527
rect 3476 3516 3507 3523
rect 3493 3513 3507 3516
rect 3296 3267 3303 3273
rect 3253 3253 3267 3267
rect 3273 3233 3287 3247
rect 3293 3253 3307 3267
rect 3276 3147 3283 3233
rect 3216 3047 3223 3113
rect 3213 3033 3227 3047
rect 3256 3003 3263 3053
rect 3276 3047 3283 3073
rect 3273 3033 3287 3047
rect 3247 2996 3263 3003
rect 3296 2847 3303 2933
rect 3196 2787 3203 2793
rect 3173 2753 3187 2767
rect 3193 2773 3207 2787
rect 3176 2667 3183 2753
rect 3056 2576 3123 2583
rect 3056 2567 3063 2576
rect 3116 2567 3123 2576
rect 3053 2553 3067 2567
rect 2996 2536 3023 2543
rect 2976 2327 2983 2533
rect 2956 2007 2963 2113
rect 2996 2007 3003 2536
rect 3073 2533 3087 2547
rect 3113 2543 3127 2547
rect 3113 2536 3143 2543
rect 3113 2533 3127 2536
rect 3076 2467 3083 2533
rect 3016 2307 3023 2413
rect 3056 2307 3063 2313
rect 3053 2293 3067 2307
rect 3036 2147 3043 2253
rect 3013 2033 3027 2047
rect 3053 2033 3067 2047
rect 3016 1983 3023 2033
rect 3056 2027 3063 2033
rect 3056 2007 3063 2013
rect 2996 1976 3023 1983
rect 2996 1867 3003 1976
rect 3016 1807 3023 1933
rect 3036 1827 3043 1993
rect 2993 1773 3007 1787
rect 3013 1793 3027 1807
rect 3033 1773 3047 1787
rect 2916 1367 2923 1373
rect 2856 1287 2863 1353
rect 2916 1327 2923 1353
rect 2913 1313 2927 1327
rect 2933 1293 2947 1307
rect 2816 1127 2823 1173
rect 2836 1147 2843 1273
rect 2833 1133 2847 1147
rect 2936 1143 2943 1293
rect 2956 1187 2963 1773
rect 2996 1767 3003 1773
rect 3036 1767 3043 1773
rect 2996 1607 3003 1633
rect 3056 1627 3063 1993
rect 3076 1763 3083 1953
rect 3096 1827 3103 2373
rect 3136 2307 3143 2536
rect 3156 2527 3163 2553
rect 3176 2507 3183 2573
rect 3196 2567 3203 2593
rect 3216 2587 3223 2773
rect 3236 2747 3243 2793
rect 3256 2727 3263 2793
rect 3276 2763 3283 2833
rect 3316 2787 3323 3313
rect 3336 3227 3343 3453
rect 3356 3367 3363 3453
rect 3416 3367 3423 3433
rect 3336 3067 3343 3113
rect 3333 3053 3347 3067
rect 3356 3047 3363 3153
rect 3396 3087 3403 3253
rect 3353 3033 3367 3047
rect 3376 2947 3383 3033
rect 3293 2763 3307 2767
rect 3276 2756 3307 2763
rect 3293 2753 3307 2756
rect 3353 2733 3367 2747
rect 3356 2727 3363 2733
rect 3236 2547 3243 2593
rect 3196 2487 3203 2533
rect 3233 2533 3247 2547
rect 3276 2527 3283 2553
rect 3196 2367 3203 2413
rect 3176 2307 3183 2333
rect 3133 2303 3147 2307
rect 3116 2296 3147 2303
rect 3116 2247 3123 2296
rect 3133 2293 3147 2296
rect 3153 2273 3167 2287
rect 3173 2293 3187 2307
rect 3156 2247 3163 2273
rect 3196 2267 3203 2333
rect 3216 2267 3223 2493
rect 3296 2467 3303 2673
rect 3207 2236 3213 2243
rect 3136 2067 3143 2173
rect 3113 2033 3127 2047
rect 3133 2053 3147 2067
rect 3153 2043 3167 2047
rect 3176 2043 3183 2093
rect 3153 2036 3183 2043
rect 3153 2033 3167 2036
rect 3116 1827 3123 2033
rect 3133 1773 3147 1787
rect 3076 1756 3103 1763
rect 3036 1607 3043 1613
rect 2993 1593 3007 1607
rect 3013 1573 3027 1587
rect 3033 1593 3047 1607
rect 3076 1603 3083 1733
rect 3056 1596 3083 1603
rect 2976 1307 2983 1533
rect 3016 1527 3023 1573
rect 2996 1203 3003 1353
rect 3036 1343 3043 1373
rect 3056 1367 3063 1596
rect 3073 1563 3087 1567
rect 3096 1563 3103 1756
rect 3136 1683 3143 1773
rect 3116 1676 3143 1683
rect 3116 1607 3123 1676
rect 3156 1663 3163 1873
rect 3176 1727 3183 1933
rect 3196 1687 3203 2033
rect 3216 1807 3223 2073
rect 3236 2067 3243 2353
rect 3256 2307 3263 2393
rect 3316 2307 3323 2673
rect 3376 2667 3383 2773
rect 3396 2687 3403 2993
rect 3416 2787 3423 3353
rect 3436 3187 3443 3513
rect 3533 3513 3547 3527
rect 3456 3427 3463 3473
rect 3496 3447 3503 3473
rect 3556 3387 3563 3553
rect 3576 3327 3583 3733
rect 3596 3463 3603 4173
rect 3656 4167 3663 4193
rect 3616 3687 3623 4153
rect 3716 4087 3723 4593
rect 3736 4187 3743 4633
rect 3776 4627 3783 4633
rect 3816 4507 3823 4553
rect 3813 4493 3827 4507
rect 3816 4227 3823 4453
rect 3753 4203 3767 4207
rect 3753 4196 3783 4203
rect 3753 4193 3767 4196
rect 3636 3807 3643 4073
rect 3716 4007 3723 4053
rect 3736 4027 3743 4073
rect 3776 4047 3783 4196
rect 3813 4213 3827 4227
rect 3836 4207 3843 4693
rect 3873 4693 3887 4707
rect 3876 4663 3883 4693
rect 3893 4673 3907 4687
rect 3913 4693 3927 4707
rect 3867 4656 3883 4663
rect 3856 4467 3863 4653
rect 3896 4647 3903 4673
rect 3896 4627 3903 4633
rect 3936 4607 3943 4933
rect 3976 4867 3983 5193
rect 4076 5187 4083 5353
rect 4013 5163 4027 5167
rect 4013 5156 4043 5163
rect 4013 5153 4027 5156
rect 3996 5087 4003 5153
rect 4016 5127 4023 5133
rect 4016 4947 4023 4973
rect 4013 4933 4027 4947
rect 4036 4927 4043 5156
rect 4073 5173 4087 5187
rect 4056 4947 4063 4953
rect 4053 4933 4067 4947
rect 3956 4707 3963 4793
rect 3896 4467 3903 4493
rect 3893 4453 3907 4467
rect 3913 4443 3927 4447
rect 3936 4443 3943 4553
rect 3913 4436 3943 4443
rect 3913 4433 3927 4436
rect 3916 4227 3923 4253
rect 3976 4247 3983 4853
rect 4053 4703 4067 4707
rect 3993 4673 4007 4687
rect 4033 4673 4047 4687
rect 4053 4696 4083 4703
rect 4053 4693 4067 4696
rect 3996 4667 4003 4673
rect 3953 4223 3967 4227
rect 3953 4216 3983 4223
rect 3953 4213 3967 4216
rect 3976 4187 3983 4216
rect 3996 4167 4003 4653
rect 4036 4607 4043 4673
rect 4076 4647 4083 4696
rect 4016 4487 4023 4493
rect 4013 4473 4027 4487
rect 4036 4447 4043 4593
rect 4096 4527 4103 5053
rect 4136 5027 4143 5373
rect 4216 5367 4223 5393
rect 4173 5153 4187 5167
rect 4176 5127 4183 5153
rect 4256 5147 4263 5173
rect 4233 5133 4247 5147
rect 4116 4927 4123 4953
rect 4136 4943 4143 4973
rect 4176 4967 4183 5113
rect 4236 5047 4243 5133
rect 4153 4943 4167 4947
rect 4136 4936 4167 4943
rect 4136 4903 4143 4936
rect 4153 4933 4167 4936
rect 4116 4896 4143 4903
rect 4116 4547 4123 4896
rect 4156 4687 4163 4753
rect 4176 4687 4183 4693
rect 4153 4673 4167 4687
rect 4176 4647 4183 4673
rect 4236 4607 4243 5013
rect 4276 4967 4283 5333
rect 4296 5103 4303 5153
rect 4313 5133 4327 5147
rect 4373 5153 4387 5167
rect 4376 5147 4383 5153
rect 4316 5127 4323 5133
rect 4296 5096 4323 5103
rect 4316 4967 4323 5096
rect 4376 4967 4383 4973
rect 4313 4953 4327 4967
rect 4373 4963 4387 4967
rect 4276 4887 4283 4893
rect 4276 4727 4283 4873
rect 4276 4707 4283 4713
rect 4273 4693 4287 4707
rect 4296 4687 4303 4953
rect 4356 4956 4387 4963
rect 4356 4927 4363 4956
rect 4373 4953 4387 4956
rect 4333 4913 4347 4927
rect 4336 4827 4343 4913
rect 4253 4653 4267 4667
rect 4313 4653 4327 4667
rect 4256 4627 4263 4653
rect 4056 4487 4063 4513
rect 4116 4507 4123 4533
rect 4116 4487 4123 4493
rect 4053 4473 4067 4487
rect 4113 4473 4127 4487
rect 4173 4483 4187 4487
rect 4173 4476 4203 4483
rect 4173 4473 4187 4476
rect 4153 4433 4167 4447
rect 4036 4263 4043 4433
rect 4156 4427 4163 4433
rect 4036 4256 4063 4263
rect 3733 4013 3747 4027
rect 3673 3973 3687 3987
rect 3713 3993 3727 4007
rect 3676 3967 3683 3973
rect 3636 3707 3643 3793
rect 3716 3747 3723 3933
rect 3653 3693 3667 3707
rect 3616 3507 3623 3573
rect 3636 3527 3643 3613
rect 3656 3567 3663 3693
rect 3673 3673 3687 3687
rect 3676 3647 3683 3673
rect 3676 3527 3683 3613
rect 3633 3513 3647 3527
rect 3613 3493 3627 3507
rect 3673 3513 3687 3527
rect 3596 3456 3623 3463
rect 3596 3303 3603 3393
rect 3576 3296 3603 3303
rect 3436 3127 3443 3173
rect 3456 3007 3463 3273
rect 3513 3253 3527 3267
rect 3493 3233 3507 3247
rect 3436 2787 3443 2953
rect 3476 2807 3483 3133
rect 3496 3047 3503 3233
rect 3516 3167 3523 3253
rect 3536 3143 3543 3213
rect 3516 3136 3543 3143
rect 3516 3047 3523 3136
rect 3556 3047 3563 3193
rect 3576 3147 3583 3296
rect 3616 3287 3623 3456
rect 3676 3267 3683 3453
rect 3696 3427 3703 3533
rect 3696 3227 3703 3393
rect 3613 3193 3627 3207
rect 3616 3167 3623 3193
rect 3513 3033 3527 3047
rect 3496 3027 3503 3033
rect 3493 3013 3507 3027
rect 3533 3013 3547 3027
rect 3536 3007 3543 3013
rect 3516 2823 3523 2993
rect 3516 2816 3543 2823
rect 3453 2783 3467 2787
rect 3453 2776 3483 2783
rect 3453 2773 3467 2776
rect 3336 2487 3343 2653
rect 3376 2547 3383 2553
rect 3416 2547 3423 2713
rect 3373 2533 3387 2547
rect 3413 2533 3427 2547
rect 3287 2296 3293 2303
rect 3336 2287 3343 2353
rect 3256 2187 3263 2273
rect 3333 2273 3347 2287
rect 3313 2233 3327 2247
rect 3316 2227 3323 2233
rect 3356 2187 3363 2493
rect 3436 2467 3443 2513
rect 3376 2327 3383 2353
rect 3396 2307 3403 2433
rect 3296 2087 3303 2113
rect 3293 2073 3307 2087
rect 3233 1773 3247 1787
rect 3236 1667 3243 1773
rect 3256 1727 3263 1973
rect 3276 1807 3283 2053
rect 3316 2047 3323 2113
rect 3336 2047 3343 2173
rect 3273 1793 3287 1807
rect 3296 1747 3303 1773
rect 3316 1687 3323 1813
rect 3356 1787 3363 2093
rect 3376 1847 3383 2293
rect 3416 2287 3423 2433
rect 3456 2387 3463 2693
rect 3476 2687 3483 2776
rect 3516 2747 3523 2793
rect 3493 2743 3507 2747
rect 3493 2736 3513 2743
rect 3493 2733 3507 2736
rect 3476 2567 3483 2653
rect 3393 2253 3407 2267
rect 3433 2263 3447 2267
rect 3456 2263 3463 2353
rect 3476 2327 3483 2473
rect 3396 2227 3403 2253
rect 3433 2256 3463 2263
rect 3433 2253 3447 2256
rect 3413 2233 3427 2247
rect 3416 2187 3423 2233
rect 3396 2087 3403 2173
rect 3393 2073 3407 2087
rect 3413 2033 3427 2047
rect 3416 1827 3423 2033
rect 3136 1656 3163 1663
rect 3073 1556 3103 1563
rect 3073 1553 3087 1556
rect 3116 1407 3123 1533
rect 3136 1527 3143 1656
rect 3157 1507 3165 1633
rect 3177 1549 3185 1633
rect 3177 1507 3185 1535
rect 3197 1507 3205 1633
rect 3216 1423 3223 1653
rect 3236 1627 3243 1633
rect 3233 1613 3247 1627
rect 3255 1579 3263 1636
rect 3283 1597 3291 1636
rect 3236 1447 3243 1573
rect 3255 1524 3263 1565
rect 3283 1524 3291 1583
rect 3316 1545 3324 1636
rect 3337 1521 3345 1636
rect 3355 1545 3363 1636
rect 3355 1506 3363 1531
rect 3376 1523 3383 1813
rect 3413 1753 3427 1767
rect 3396 1543 3403 1753
rect 3416 1707 3423 1753
rect 3413 1583 3427 1587
rect 3436 1583 3443 2153
rect 3476 2127 3483 2313
rect 3496 2267 3503 2713
rect 3536 2667 3543 2816
rect 3553 2733 3567 2747
rect 3616 2747 3623 3133
rect 3696 3127 3703 3193
rect 3656 3047 3663 3053
rect 3696 3047 3703 3113
rect 3653 3033 3667 3047
rect 3636 3027 3643 3033
rect 3633 3013 3647 3027
rect 3673 3013 3687 3027
rect 3693 3033 3707 3047
rect 3676 3007 3683 3013
rect 3716 2847 3723 3733
rect 3736 3667 3743 3713
rect 3756 3543 3763 3993
rect 3776 3927 3783 4033
rect 3796 3963 3803 4053
rect 3813 3963 3827 3967
rect 3796 3956 3827 3963
rect 3853 3963 3867 3967
rect 3876 3963 3883 4073
rect 3813 3953 3827 3956
rect 3853 3956 3883 3963
rect 3853 3953 3867 3956
rect 3816 3747 3823 3833
rect 3793 3713 3807 3727
rect 3813 3733 3827 3747
rect 3796 3683 3803 3713
rect 3776 3676 3803 3683
rect 3776 3587 3783 3676
rect 3836 3667 3843 3753
rect 3736 3536 3763 3543
rect 3736 2823 3743 3536
rect 3796 3467 3803 3653
rect 3813 3523 3827 3527
rect 3813 3516 3843 3523
rect 3813 3513 3827 3516
rect 3836 3507 3843 3516
rect 3796 3247 3803 3453
rect 3836 3407 3843 3493
rect 3753 3233 3767 3247
rect 3756 3067 3763 3233
rect 3773 3213 3787 3227
rect 3793 3233 3807 3247
rect 3836 3227 3843 3233
rect 3813 3223 3827 3227
rect 3813 3216 3833 3223
rect 3813 3213 3827 3216
rect 3776 3167 3783 3213
rect 3736 2816 3763 2823
rect 3556 2687 3563 2733
rect 3533 2563 3547 2567
rect 3533 2556 3563 2563
rect 3533 2553 3547 2556
rect 3513 2513 3527 2527
rect 3516 2507 3523 2513
rect 3413 1576 3443 1583
rect 3413 1573 3427 1576
rect 3396 1536 3423 1543
rect 3376 1516 3403 1523
rect 3216 1416 3243 1423
rect 3036 1336 3063 1343
rect 3056 1327 3063 1336
rect 3196 1327 3203 1353
rect 3053 1313 3067 1327
rect 3073 1293 3087 1307
rect 3173 1293 3187 1307
rect 3193 1313 3207 1327
rect 3213 1293 3227 1307
rect 2976 1196 3023 1203
rect 2813 1113 2827 1127
rect 2916 1136 2943 1143
rect 2853 1123 2867 1127
rect 2853 1116 2883 1123
rect 2853 1113 2867 1116
rect 2876 1047 2883 1116
rect 2896 867 2903 1113
rect 2916 987 2923 1136
rect 2976 1127 2983 1196
rect 2973 1113 2987 1127
rect 2976 947 2983 1073
rect 2936 867 2943 873
rect 2753 863 2767 867
rect 2736 856 2767 863
rect 2793 863 2807 867
rect 2736 827 2743 856
rect 2753 853 2767 856
rect 2793 856 2823 863
rect 2793 853 2807 856
rect 2693 793 2707 807
rect 2696 787 2703 793
rect 2816 787 2823 856
rect 2713 643 2727 647
rect 2696 636 2727 643
rect 2856 647 2863 853
rect 2913 833 2927 847
rect 2933 853 2947 867
rect 2753 643 2767 647
rect 2813 643 2827 647
rect 2593 593 2607 607
rect 2633 593 2647 607
rect 2596 547 2603 593
rect 2636 527 2643 593
rect 2696 547 2703 636
rect 2713 633 2727 636
rect 2753 636 2783 643
rect 2753 633 2767 636
rect 2513 383 2527 387
rect 2496 376 2527 383
rect 2213 156 2243 163
rect 2253 163 2267 167
rect 2253 156 2283 163
rect 2213 153 2227 156
rect 2253 153 2267 156
rect 2153 133 2167 136
rect 796 107 803 113
rect 1856 107 1863 113
rect 2096 107 2103 113
rect 2276 47 2283 156
rect 2336 123 2343 153
rect 2376 147 2383 293
rect 2496 163 2503 376
rect 2513 373 2527 376
rect 2573 363 2587 367
rect 2596 363 2603 433
rect 2636 407 2643 513
rect 2656 367 2663 453
rect 2573 356 2603 363
rect 2573 353 2587 356
rect 2576 327 2583 353
rect 2633 333 2647 347
rect 2653 353 2667 367
rect 2693 353 2707 367
rect 2696 347 2703 353
rect 2636 307 2643 333
rect 2716 207 2723 393
rect 2736 367 2743 613
rect 2776 527 2783 636
rect 2796 636 2827 643
rect 2796 587 2803 636
rect 2813 633 2827 636
rect 2853 633 2867 647
rect 2876 627 2883 653
rect 2873 613 2887 627
rect 2796 367 2803 513
rect 2916 467 2923 833
rect 2996 807 3003 1173
rect 3016 847 3023 1196
rect 3036 847 3043 1273
rect 3056 1127 3063 1133
rect 3076 1127 3083 1293
rect 3053 1113 3067 1127
rect 3136 1067 3143 1293
rect 3176 1227 3183 1293
rect 3156 1087 3163 1153
rect 3033 833 3047 847
rect 3013 793 3027 807
rect 2793 353 2807 367
rect 2516 167 2523 193
rect 2353 123 2367 127
rect 2336 116 2367 123
rect 2373 133 2387 147
rect 2476 156 2503 163
rect 2476 127 2483 156
rect 2513 153 2527 167
rect 2716 147 2723 193
rect 2756 167 2763 333
rect 2836 327 2843 413
rect 2876 347 2883 373
rect 2893 333 2907 347
rect 2896 327 2903 333
rect 2813 323 2827 327
rect 2813 316 2833 323
rect 2813 313 2827 316
rect 2753 153 2767 167
rect 2813 163 2827 167
rect 2813 156 2843 163
rect 2813 153 2827 156
rect 2353 113 2367 116
rect 2493 123 2507 127
rect 2487 116 2507 123
rect 2493 113 2507 116
rect 2836 147 2843 156
rect 2916 147 2923 153
rect 2773 113 2787 127
rect 2893 113 2907 127
rect 2913 133 2927 147
rect 2776 107 2783 113
rect 2896 107 2903 113
rect 2636 -24 2643 13
rect 2676 -24 2683 33
rect 2956 27 2963 793
rect 3016 783 3023 793
rect 2996 776 3023 783
rect 2996 627 3003 776
rect 2976 107 2983 533
rect 2996 127 3003 313
rect 3036 187 3043 633
rect 3056 407 3063 833
rect 3116 807 3123 873
rect 3096 343 3103 573
rect 3156 547 3163 633
rect 3176 627 3183 833
rect 3196 667 3203 1233
rect 3216 1187 3223 1293
rect 3216 1127 3223 1173
rect 3236 1147 3243 1416
rect 3256 1147 3263 1473
rect 3276 1287 3283 1473
rect 3296 1327 3303 1393
rect 3396 1327 3403 1516
rect 3293 1313 3307 1327
rect 3393 1313 3407 1327
rect 3416 1307 3423 1536
rect 3436 1507 3443 1553
rect 3373 1273 3387 1287
rect 3376 1247 3383 1273
rect 3376 1147 3383 1153
rect 3233 1133 3247 1147
rect 3373 1133 3387 1147
rect 3213 1113 3227 1127
rect 3253 1123 3267 1127
rect 3253 1116 3283 1123
rect 3253 1113 3267 1116
rect 3236 643 3243 1093
rect 3276 1067 3283 1116
rect 3353 1123 3367 1127
rect 3336 1116 3367 1123
rect 3396 1127 3403 1133
rect 3256 867 3263 913
rect 3253 853 3267 867
rect 3273 833 3287 847
rect 3276 787 3283 833
rect 3316 647 3323 1113
rect 3336 1047 3343 1116
rect 3353 1113 3367 1116
rect 3393 1113 3407 1127
rect 3336 807 3343 1033
rect 3416 847 3423 1213
rect 3436 1207 3443 1493
rect 3456 1467 3463 1973
rect 3496 1927 3503 2233
rect 3516 2207 3523 2373
rect 3556 2287 3563 2556
rect 3576 2487 3583 2653
rect 3596 2503 3603 2693
rect 3636 2547 3643 2673
rect 3656 2567 3663 2793
rect 3736 2787 3743 2793
rect 3673 2753 3687 2767
rect 3733 2773 3747 2787
rect 3756 2767 3763 2816
rect 3676 2747 3683 2753
rect 3633 2533 3647 2547
rect 3653 2513 3667 2527
rect 3596 2496 3623 2503
rect 3576 2307 3583 2473
rect 3553 2273 3567 2287
rect 3593 2273 3607 2287
rect 3596 2187 3603 2273
rect 3576 2087 3583 2093
rect 3573 2073 3587 2087
rect 3556 2047 3563 2053
rect 3616 2047 3623 2496
rect 3656 2487 3663 2513
rect 3676 2507 3683 2713
rect 3636 2267 3643 2373
rect 3656 2247 3663 2373
rect 3676 2307 3683 2393
rect 3696 2387 3703 2673
rect 3736 2587 3743 2733
rect 3756 2587 3763 2753
rect 3716 2563 3723 2573
rect 3776 2567 3783 2733
rect 3796 2707 3803 3153
rect 3836 3003 3843 3013
rect 3816 2996 3843 3003
rect 3816 2947 3823 2996
rect 3836 2803 3843 2893
rect 3856 2827 3863 3933
rect 3896 3827 3903 4033
rect 3916 3727 3923 3773
rect 3913 3713 3927 3727
rect 3893 3673 3907 3687
rect 3896 3647 3903 3673
rect 3876 3527 3883 3593
rect 3896 3547 3903 3613
rect 3893 3533 3907 3547
rect 3916 3207 3923 3373
rect 3876 3087 3883 3193
rect 3876 2987 3883 3033
rect 3896 3007 3903 3033
rect 3836 2796 3863 2803
rect 3856 2787 3863 2796
rect 3833 2753 3847 2767
rect 3853 2773 3867 2787
rect 3836 2647 3843 2753
rect 3816 2567 3823 2573
rect 3733 2563 3747 2567
rect 3716 2556 3747 2563
rect 3733 2553 3747 2556
rect 3753 2533 3767 2547
rect 3773 2553 3787 2567
rect 3813 2553 3827 2567
rect 3716 2447 3723 2533
rect 3756 2527 3763 2533
rect 3673 2293 3687 2307
rect 3713 2303 3727 2307
rect 3736 2303 3743 2513
rect 3693 2273 3707 2287
rect 3713 2296 3743 2303
rect 3713 2293 3727 2296
rect 3696 2267 3703 2273
rect 3496 1867 3503 1913
rect 3536 1807 3543 1913
rect 3473 1773 3487 1787
rect 3513 1773 3527 1787
rect 3533 1793 3547 1807
rect 3553 1773 3567 1787
rect 3476 1747 3483 1773
rect 3476 1567 3483 1693
rect 3493 1573 3507 1587
rect 3456 1307 3463 1373
rect 3436 1027 3443 1133
rect 3433 813 3447 827
rect 3436 787 3443 813
rect 3216 636 3243 643
rect 3176 467 3183 613
rect 3136 367 3143 413
rect 3216 407 3223 636
rect 3276 607 3283 633
rect 3273 593 3287 607
rect 3156 367 3163 373
rect 3256 367 3263 553
rect 3316 427 3323 633
rect 3376 627 3383 653
rect 3296 367 3303 373
rect 3113 343 3127 347
rect 3096 336 3127 343
rect 3133 353 3147 367
rect 3113 333 3127 336
rect 3293 353 3307 367
rect 3313 333 3327 347
rect 3316 223 3323 333
rect 3336 327 3343 613
rect 3373 613 3387 627
rect 3393 603 3407 607
rect 3416 603 3423 653
rect 3393 596 3423 603
rect 3393 593 3407 596
rect 3356 567 3363 593
rect 3416 367 3423 393
rect 3456 367 3463 1273
rect 3476 1207 3483 1533
rect 3496 1387 3503 1573
rect 3516 1547 3523 1773
rect 3556 1687 3563 1773
rect 3536 1547 3543 1593
rect 3493 1293 3507 1307
rect 3496 1227 3503 1293
rect 3496 1147 3503 1173
rect 3493 1133 3507 1147
rect 3473 1093 3487 1107
rect 3476 867 3483 1093
rect 3516 1007 3523 1513
rect 3536 1447 3543 1473
rect 3556 1167 3563 1613
rect 3576 1267 3583 1813
rect 3596 1627 3603 2013
rect 3636 1963 3643 2073
rect 3656 2027 3663 2213
rect 3676 2107 3683 2253
rect 3693 2083 3707 2087
rect 3676 2076 3707 2083
rect 3676 2007 3683 2076
rect 3693 2073 3707 2076
rect 3716 1987 3723 2033
rect 3616 1956 3643 1963
rect 3616 1907 3623 1956
rect 3616 1787 3623 1833
rect 3636 1767 3643 1933
rect 3696 1807 3703 1893
rect 3653 1793 3667 1807
rect 3656 1767 3663 1793
rect 3673 1773 3687 1787
rect 3693 1793 3707 1807
rect 3656 1747 3663 1753
rect 3636 1627 3643 1713
rect 3676 1687 3683 1773
rect 3633 1613 3647 1627
rect 3613 1573 3627 1587
rect 3616 1567 3623 1573
rect 3596 1187 3603 1533
rect 3656 1407 3663 1573
rect 3676 1567 3683 1613
rect 3696 1587 3703 1713
rect 3736 1667 3743 2273
rect 3756 1647 3763 2353
rect 3776 2247 3783 2473
rect 3796 2307 3803 2513
rect 3816 2427 3823 2493
rect 3793 2253 3807 2267
rect 3796 2207 3803 2253
rect 3816 2187 3823 2413
rect 3836 2307 3843 2613
rect 3856 2547 3863 2573
rect 3856 2347 3863 2513
rect 3833 2253 3847 2267
rect 3836 2247 3843 2253
rect 3776 2047 3783 2173
rect 3836 2087 3843 2233
rect 3856 2223 3863 2333
rect 3876 2243 3883 2813
rect 3916 2707 3923 3173
rect 3936 3147 3943 3993
rect 4036 3967 4043 4233
rect 4056 4227 4063 4256
rect 4096 4227 4103 4233
rect 4073 4193 4087 4207
rect 4093 4213 4107 4227
rect 3996 3683 4003 3953
rect 4033 3683 4047 3687
rect 4056 3683 4063 4173
rect 4076 4007 4083 4193
rect 4136 4067 4143 4213
rect 4156 4107 4163 4413
rect 4196 4267 4203 4476
rect 4236 4307 4243 4573
rect 4316 4547 4323 4653
rect 4176 4227 4183 4253
rect 4173 4213 4187 4227
rect 4213 4223 4227 4227
rect 4236 4223 4243 4293
rect 4213 4216 4243 4223
rect 4213 4213 4227 4216
rect 4236 4187 4243 4216
rect 4096 4007 4103 4053
rect 4136 4027 4143 4033
rect 4133 4013 4147 4027
rect 4093 3993 4107 4007
rect 4153 3983 4167 3987
rect 4176 3983 4183 4053
rect 4153 3976 4183 3983
rect 4153 3973 4167 3976
rect 4196 3947 4203 4173
rect 4256 4047 4263 4473
rect 4313 4433 4327 4447
rect 4316 4407 4323 4433
rect 4336 4407 4343 4673
rect 4276 4387 4283 4393
rect 4213 3953 4227 3967
rect 4253 3953 4267 3967
rect 4216 3947 4223 3953
rect 4256 3847 4263 3953
rect 4097 3758 4105 3782
rect 3996 3676 4023 3683
rect 3976 3487 3983 3613
rect 3996 3527 4003 3633
rect 3977 3278 3985 3302
rect 3956 3247 3963 3253
rect 3956 3227 3963 3233
rect 3953 3213 3967 3227
rect 3977 3184 3985 3264
rect 3996 3167 4003 3373
rect 4016 3367 4023 3676
rect 4033 3676 4063 3683
rect 4033 3673 4047 3676
rect 4036 3627 4043 3673
rect 4097 3664 4105 3744
rect 4136 3667 4143 3713
rect 4153 3693 4167 3707
rect 4193 3693 4207 3707
rect 4156 3607 4163 3693
rect 4196 3587 4203 3693
rect 4056 3527 4063 3533
rect 4053 3513 4067 3527
rect 4093 3523 4107 3527
rect 4073 3493 4087 3507
rect 4093 3516 4123 3523
rect 4093 3513 4107 3516
rect 4116 3507 4123 3516
rect 4076 3483 4083 3493
rect 4056 3476 4083 3483
rect 3953 2993 3967 3007
rect 3956 2987 3963 2993
rect 3976 2807 3983 3133
rect 3996 3047 4003 3053
rect 4016 2907 4023 3253
rect 4033 3213 4047 3227
rect 4036 3167 4043 3213
rect 4056 3067 4063 3476
rect 4076 3467 4083 3476
rect 4073 3213 4087 3227
rect 4076 3187 4083 3213
rect 4076 3067 4083 3113
rect 4096 3067 4103 3233
rect 4116 3184 4124 3296
rect 4073 3053 4087 3067
rect 4053 3043 4067 3047
rect 4047 3036 4067 3043
rect 4093 3043 4107 3047
rect 4053 3033 4067 3036
rect 3936 2567 3943 2793
rect 3996 2787 4003 2793
rect 4016 2787 4023 2873
rect 3953 2733 3967 2747
rect 3956 2647 3963 2733
rect 3996 2687 4003 2773
rect 3933 2553 3947 2567
rect 3876 2236 3903 2243
rect 3856 2216 3883 2223
rect 3796 2067 3803 2073
rect 3793 2053 3807 2067
rect 3853 2043 3867 2047
rect 3876 2043 3883 2216
rect 3853 2036 3883 2043
rect 3853 2033 3867 2036
rect 3776 1787 3783 2013
rect 3776 1747 3783 1773
rect 3756 1607 3763 1613
rect 3753 1593 3767 1607
rect 3736 1547 3743 1573
rect 3796 1427 3803 1873
rect 3856 1807 3863 1833
rect 3813 1793 3827 1807
rect 3816 1767 3823 1793
rect 3853 1793 3867 1807
rect 3873 1773 3887 1787
rect 3876 1767 3883 1773
rect 3856 1756 3873 1763
rect 3836 1443 3843 1593
rect 3856 1527 3863 1756
rect 3896 1707 3903 2236
rect 3916 2007 3923 2533
rect 3936 2063 3943 2493
rect 3976 2343 3983 2653
rect 3993 2533 4007 2547
rect 3996 2367 4003 2533
rect 4016 2487 4023 2773
rect 4036 2527 4043 3033
rect 4093 3036 4123 3043
rect 4093 3033 4107 3036
rect 4116 2987 4123 3036
rect 4053 2753 4067 2767
rect 4056 2707 4063 2753
rect 4073 2733 4087 2747
rect 4113 2733 4127 2747
rect 4076 2727 4083 2733
rect 4116 2727 4123 2733
rect 4136 2707 4143 3313
rect 4156 3047 4163 3333
rect 4176 3127 4183 3473
rect 4196 3247 4203 3553
rect 4216 3547 4223 3693
rect 4236 3664 4244 3776
rect 4256 3563 4263 3833
rect 4276 3567 4283 4373
rect 4356 4223 4363 4453
rect 4376 4427 4383 4913
rect 4396 4487 4403 5073
rect 4416 4947 4423 5213
rect 4416 4727 4423 4933
rect 4436 4887 4443 5473
rect 4536 5447 4543 5513
rect 4556 5507 4563 5633
rect 4576 5607 4583 5636
rect 4593 5633 4607 5636
rect 4733 5633 4747 5647
rect 4833 5633 4847 5647
rect 4576 5527 4583 5593
rect 4613 5463 4627 5467
rect 4596 5456 4627 5463
rect 4596 5447 4603 5456
rect 4613 5453 4627 5456
rect 4533 5433 4547 5447
rect 4716 5447 4723 5493
rect 4756 5447 4763 5453
rect 4713 5433 4727 5447
rect 4733 5413 4747 5427
rect 4753 5433 4767 5447
rect 4816 5443 4823 5593
rect 4833 5443 4847 5447
rect 4816 5436 4847 5443
rect 4833 5433 4847 5436
rect 4773 5423 4787 5427
rect 4773 5416 4803 5423
rect 4773 5413 4787 5416
rect 4476 5367 4483 5413
rect 4516 5407 4523 5413
rect 4736 5407 4743 5413
rect 4473 4963 4487 4967
rect 4473 4956 4493 4963
rect 4473 4953 4487 4956
rect 4496 4827 4503 4953
rect 4513 4943 4527 4947
rect 4536 4943 4543 5133
rect 4513 4936 4543 4943
rect 4513 4933 4527 4936
rect 4556 4927 4563 5393
rect 4796 5383 4803 5416
rect 4776 5376 4803 5383
rect 4576 5187 4583 5193
rect 4573 5173 4587 5187
rect 4613 5173 4627 5187
rect 4593 5153 4607 5167
rect 4596 5147 4603 5153
rect 4616 5127 4623 5173
rect 4656 5047 4663 5133
rect 4616 4987 4623 5033
rect 4613 4973 4627 4987
rect 4596 4967 4603 4973
rect 4593 4953 4607 4967
rect 4676 4943 4683 5253
rect 4753 5143 4767 5147
rect 4776 5143 4783 5376
rect 4753 5136 4783 5143
rect 4753 5133 4767 5136
rect 4656 4936 4683 4943
rect 4616 4847 4623 4913
rect 4453 4693 4467 4707
rect 4456 4647 4463 4693
rect 4476 4547 4483 4673
rect 4453 4483 4467 4487
rect 4476 4483 4483 4513
rect 4433 4453 4447 4467
rect 4453 4476 4483 4483
rect 4453 4473 4467 4476
rect 4436 4447 4443 4453
rect 4476 4323 4483 4476
rect 4496 4447 4503 4713
rect 4596 4707 4603 4813
rect 4553 4693 4567 4707
rect 4536 4467 4543 4593
rect 4556 4587 4563 4693
rect 4573 4673 4587 4687
rect 4593 4693 4607 4707
rect 4576 4667 4583 4673
rect 4533 4453 4547 4467
rect 4553 4433 4567 4447
rect 4476 4316 4503 4323
rect 4356 4216 4383 4223
rect 4293 4193 4307 4207
rect 4296 4127 4303 4193
rect 4353 4183 4367 4187
rect 4376 4183 4383 4216
rect 4353 4176 4383 4183
rect 4353 4173 4367 4176
rect 4376 4167 4383 4176
rect 4396 4127 4403 4173
rect 4496 4147 4503 4316
rect 4556 4307 4563 4433
rect 4596 4347 4603 4633
rect 4616 4367 4623 4833
rect 4656 4623 4663 4936
rect 4696 4687 4703 4733
rect 4656 4616 4683 4623
rect 4676 4467 4683 4616
rect 4653 4433 4667 4447
rect 4673 4453 4687 4467
rect 4693 4433 4707 4447
rect 4656 4403 4663 4433
rect 4696 4407 4703 4433
rect 4656 4396 4683 4403
rect 4596 4227 4603 4333
rect 4296 3603 4303 4093
rect 4336 4007 4343 4113
rect 4376 4007 4383 4033
rect 4373 3993 4387 4007
rect 4473 4003 4487 4007
rect 4456 3996 4487 4003
rect 4296 3596 4323 3603
rect 4236 3556 4263 3563
rect 4216 3327 4223 3533
rect 4236 3267 4243 3556
rect 4256 3527 4263 3533
rect 4296 3527 4303 3573
rect 4316 3527 4323 3596
rect 4336 3563 4343 3873
rect 4376 3727 4383 3873
rect 4416 3727 4423 3893
rect 4436 3747 4443 3973
rect 4353 3693 4367 3707
rect 4413 3713 4427 3727
rect 4456 3707 4463 3996
rect 4473 3993 4487 3996
rect 4493 3973 4507 3987
rect 4536 3987 4543 3993
rect 4533 3973 4547 3987
rect 4476 3743 4483 3913
rect 4496 3767 4503 3973
rect 4556 3923 4563 4213
rect 4616 4207 4623 4293
rect 4573 4193 4587 4207
rect 4576 4127 4583 4193
rect 4593 4173 4607 4187
rect 4633 4173 4647 4187
rect 4596 4023 4603 4173
rect 4636 4167 4643 4173
rect 4656 4167 4663 4353
rect 4676 4187 4683 4396
rect 4716 4243 4723 5033
rect 4756 4967 4763 5113
rect 4796 4967 4803 5353
rect 4836 5347 4843 5433
rect 4857 5396 4865 5476
rect 4857 5358 4865 5382
rect 4876 5347 4883 5653
rect 4836 5107 4843 5133
rect 4853 5113 4867 5127
rect 4856 5087 4863 5113
rect 4896 5047 4903 5653
rect 4976 5647 4983 5673
rect 5076 5667 5083 5773
rect 5073 5663 5087 5667
rect 5056 5656 5087 5663
rect 5113 5663 5127 5667
rect 5136 5663 5143 5673
rect 4933 5633 4947 5647
rect 4936 5607 4943 5633
rect 4953 5613 4967 5627
rect 4973 5633 4987 5647
rect 5056 5627 5063 5656
rect 5073 5653 5087 5656
rect 5093 5633 5107 5647
rect 5113 5656 5143 5663
rect 5113 5653 5127 5656
rect 4916 5447 4923 5513
rect 4956 5447 4963 5613
rect 4996 5603 5003 5613
rect 5096 5607 5103 5633
rect 5136 5627 5143 5656
rect 4976 5596 5003 5603
rect 4913 5433 4927 5447
rect 4953 5433 4967 5447
rect 4957 5198 4965 5222
rect 4933 5143 4947 5147
rect 4916 5136 4947 5143
rect 4916 5067 4923 5136
rect 4933 5133 4947 5136
rect 4957 5104 4965 5184
rect 4753 4953 4767 4967
rect 4736 4947 4743 4953
rect 4733 4933 4747 4947
rect 4793 4953 4807 4967
rect 4833 4963 4847 4967
rect 4816 4956 4847 4963
rect 4777 4718 4785 4742
rect 4753 4663 4767 4667
rect 4736 4656 4767 4663
rect 4736 4647 4743 4656
rect 4753 4653 4767 4656
rect 4777 4624 4785 4704
rect 4816 4643 4823 4956
rect 4833 4953 4847 4956
rect 4857 4916 4865 4996
rect 4857 4878 4865 4902
rect 4833 4663 4847 4667
rect 4833 4656 4863 4663
rect 4833 4653 4847 4656
rect 4816 4636 4843 4643
rect 4753 4503 4767 4507
rect 4736 4496 4767 4503
rect 4736 4327 4743 4496
rect 4753 4493 4767 4496
rect 4773 4453 4787 4467
rect 4776 4447 4783 4453
rect 4696 4236 4723 4243
rect 4613 4023 4627 4027
rect 4596 4016 4627 4023
rect 4596 4007 4603 4016
rect 4613 4013 4627 4016
rect 4633 4003 4647 4007
rect 4633 3996 4653 4003
rect 4633 3993 4647 3996
rect 4556 3916 4583 3923
rect 4536 3747 4543 3833
rect 4493 3743 4507 3747
rect 4476 3736 4507 3743
rect 4533 3743 4547 3747
rect 4356 3587 4363 3693
rect 4476 3687 4483 3736
rect 4493 3733 4507 3736
rect 4533 3736 4563 3743
rect 4533 3733 4547 3736
rect 4556 3687 4563 3736
rect 4576 3683 4583 3916
rect 4656 3823 4663 3993
rect 4673 3973 4687 3987
rect 4676 3967 4683 3973
rect 4696 3827 4703 4236
rect 4736 4207 4743 4313
rect 4713 4173 4727 4187
rect 4733 4193 4747 4207
rect 4773 4203 4787 4207
rect 4796 4203 4803 4413
rect 4773 4196 4803 4203
rect 4773 4193 4787 4196
rect 4716 4147 4723 4173
rect 4716 4103 4723 4133
rect 4716 4096 4743 4103
rect 4716 3927 4723 4013
rect 4736 3907 4743 4096
rect 4756 3967 4763 4013
rect 4796 3987 4803 4196
rect 4816 4147 4823 4613
rect 4836 4587 4843 4636
rect 4836 4443 4843 4573
rect 4856 4507 4863 4656
rect 4873 4653 4887 4667
rect 4876 4647 4883 4653
rect 4896 4607 4903 4993
rect 4916 4624 4924 4736
rect 4936 4627 4943 5093
rect 4956 4967 4963 4973
rect 4953 4953 4967 4967
rect 4976 4927 4983 5596
rect 4996 5364 5004 5476
rect 5013 5143 5027 5147
rect 5036 5143 5043 5513
rect 5096 5467 5103 5473
rect 5093 5453 5107 5467
rect 5136 5447 5143 5473
rect 5113 5413 5127 5427
rect 5156 5423 5163 5753
rect 5176 5667 5183 5673
rect 5216 5667 5223 5816
rect 5236 5787 5243 5823
rect 5173 5653 5187 5667
rect 5213 5663 5227 5667
rect 5213 5656 5243 5663
rect 5213 5653 5227 5656
rect 5136 5416 5163 5423
rect 5116 5367 5123 5413
rect 5013 5136 5043 5143
rect 5013 5133 5027 5136
rect 5053 5133 5067 5147
rect 5016 5007 5023 5133
rect 5056 5087 5063 5133
rect 5076 5127 5083 5173
rect 4996 4884 5004 4996
rect 5016 4967 5023 4993
rect 5056 4887 5063 4953
rect 5056 4727 5063 4873
rect 5076 4807 5083 5113
rect 5096 5104 5104 5216
rect 5136 5107 5143 5416
rect 5197 5396 5205 5476
rect 5136 4967 5143 4973
rect 5156 4967 5163 5393
rect 5197 5358 5205 5382
rect 5113 4933 5127 4947
rect 5133 4953 5147 4967
rect 5116 4823 5123 4933
rect 5096 4816 5123 4823
rect 4956 4667 4963 4713
rect 5053 4653 5067 4667
rect 4876 4467 4883 4473
rect 4853 4443 4867 4447
rect 4836 4436 4867 4443
rect 4873 4453 4887 4467
rect 4936 4447 4943 4473
rect 4793 3973 4807 3987
rect 4636 3816 4663 3823
rect 4596 3703 4603 3793
rect 4636 3727 4643 3816
rect 4613 3703 4627 3707
rect 4596 3696 4627 3703
rect 4613 3693 4627 3696
rect 4676 3703 4683 3793
rect 4756 3727 4763 3773
rect 4667 3696 4683 3703
rect 4753 3713 4767 3727
rect 4773 3693 4787 3707
rect 4576 3676 4603 3683
rect 4336 3556 4363 3563
rect 4253 3513 4267 3527
rect 4293 3513 4307 3527
rect 4196 3107 4203 3233
rect 4213 3213 4227 3227
rect 4273 3243 4287 3247
rect 4296 3243 4303 3253
rect 4273 3236 4303 3243
rect 4273 3233 4287 3236
rect 4253 3213 4267 3227
rect 4216 3207 4223 3213
rect 4256 3187 4263 3213
rect 4336 3187 4343 3533
rect 4356 3427 4363 3556
rect 4376 3467 4383 3673
rect 4416 3603 4423 3673
rect 4396 3596 4423 3603
rect 4396 3547 4403 3596
rect 4396 3516 4503 3523
rect 4396 3507 4403 3516
rect 4496 3507 4503 3516
rect 4413 3473 4427 3487
rect 4416 3363 4423 3473
rect 4416 3356 4443 3363
rect 4353 3213 4367 3227
rect 4393 3213 4407 3227
rect 4216 3047 4223 3073
rect 4216 3027 4223 3033
rect 4173 3023 4187 3027
rect 4156 3016 4187 3023
rect 4156 2787 4163 3016
rect 4173 3013 4187 3016
rect 4213 3013 4227 3027
rect 4233 2993 4247 3007
rect 4236 2987 4243 2993
rect 4256 2827 4263 3113
rect 4256 2787 4263 2813
rect 4236 2727 4243 2753
rect 4096 2407 4103 2693
rect 4137 2505 4145 2596
rect 4137 2466 4145 2491
rect 4155 2481 4163 2596
rect 4176 2505 4184 2596
rect 4209 2557 4217 2596
rect 4209 2484 4217 2543
rect 4237 2539 4245 2596
rect 4256 2587 4263 2733
rect 4253 2573 4267 2587
rect 4237 2484 4245 2525
rect 3976 2336 4003 2343
rect 3956 2283 3963 2333
rect 3973 2283 3987 2287
rect 3956 2276 3987 2283
rect 3956 2167 3963 2276
rect 3973 2273 3987 2276
rect 3953 2063 3967 2067
rect 3936 2056 3967 2063
rect 3996 2067 4003 2336
rect 4037 2329 4045 2354
rect 4016 2087 4023 2293
rect 4037 2224 4045 2315
rect 4055 2224 4063 2339
rect 4076 2224 4084 2315
rect 4109 2277 4117 2336
rect 4137 2295 4145 2336
rect 4109 2224 4117 2263
rect 4137 2224 4145 2281
rect 3953 2053 3967 2056
rect 3936 2007 3943 2033
rect 3936 1983 3943 1993
rect 3916 1976 3943 1983
rect 3916 1827 3923 1976
rect 3956 1827 3963 2053
rect 4016 1863 4023 2053
rect 4036 1887 4043 2153
rect 4056 2047 4063 2113
rect 4016 1856 4043 1863
rect 3973 1773 3987 1787
rect 3916 1607 3923 1653
rect 3913 1593 3927 1607
rect 3836 1436 3863 1443
rect 3656 1327 3663 1333
rect 3696 1327 3703 1393
rect 3633 1293 3647 1307
rect 3653 1313 3667 1327
rect 3636 1223 3643 1293
rect 3716 1267 3723 1333
rect 3736 1287 3743 1373
rect 3776 1327 3783 1373
rect 3773 1313 3787 1327
rect 3813 1313 3827 1327
rect 3793 1293 3807 1307
rect 3796 1267 3803 1293
rect 3816 1227 3823 1313
rect 3636 1216 3663 1223
rect 3413 353 3427 367
rect 3433 313 3447 327
rect 3436 307 3443 313
rect 3316 216 3343 223
rect 3316 187 3323 193
rect 3313 173 3327 187
rect 3033 113 3047 127
rect 3153 113 3167 127
rect 3196 127 3203 173
rect 3336 147 3343 216
rect 3376 167 3383 193
rect 3373 153 3387 167
rect 3193 113 3207 127
rect 3036 107 3043 113
rect 3156 107 3163 113
rect 3476 -17 3483 833
rect 3496 823 3503 973
rect 3536 927 3543 1133
rect 3636 1127 3643 1193
rect 3633 1113 3647 1127
rect 3656 1107 3663 1216
rect 3496 816 3513 823
rect 3553 813 3567 827
rect 3556 807 3563 813
rect 3556 647 3563 673
rect 3596 663 3603 1073
rect 3656 1047 3663 1093
rect 3656 847 3663 913
rect 3676 847 3683 1173
rect 3696 1087 3703 1113
rect 3716 1107 3723 1193
rect 3776 1127 3783 1193
rect 3796 1147 3803 1173
rect 3773 1123 3787 1127
rect 3836 1123 3843 1413
rect 3856 1187 3863 1436
rect 3896 1227 3903 1573
rect 3956 1427 3963 1733
rect 3976 1707 3983 1773
rect 3996 1667 4003 1773
rect 3916 1327 3923 1353
rect 3913 1313 3927 1327
rect 3933 1273 3947 1287
rect 3713 1093 3727 1107
rect 3753 1093 3767 1107
rect 3773 1116 3803 1123
rect 3773 1113 3787 1116
rect 3756 1047 3763 1093
rect 3796 1087 3803 1116
rect 3816 1116 3843 1123
rect 3696 847 3703 973
rect 3796 947 3803 1053
rect 3816 923 3823 1116
rect 3856 1107 3863 1133
rect 3853 1093 3867 1107
rect 3796 916 3823 923
rect 3633 813 3647 827
rect 3653 833 3667 847
rect 3693 833 3707 847
rect 3636 683 3643 813
rect 3576 656 3603 663
rect 3616 676 3643 683
rect 3496 407 3503 433
rect 3576 407 3583 656
rect 3616 647 3623 676
rect 3596 603 3603 633
rect 3636 627 3643 653
rect 3613 603 3627 607
rect 3596 596 3627 603
rect 3633 613 3647 627
rect 3613 593 3627 596
rect 3496 343 3503 393
rect 3536 367 3543 373
rect 3513 343 3527 347
rect 3496 336 3527 343
rect 3533 353 3547 367
rect 3573 363 3587 367
rect 3596 363 3603 393
rect 3676 387 3683 633
rect 3696 627 3703 633
rect 3696 367 3703 453
rect 3716 383 3723 853
rect 3796 847 3803 916
rect 3773 843 3787 847
rect 3756 836 3787 843
rect 3736 647 3743 833
rect 3756 807 3763 836
rect 3773 833 3787 836
rect 3796 727 3803 773
rect 3816 667 3823 893
rect 3836 863 3843 1073
rect 3856 887 3863 933
rect 3876 907 3883 1073
rect 3896 867 3903 1113
rect 3916 1027 3923 1093
rect 3936 1083 3943 1273
rect 3976 1127 3983 1613
rect 4016 1607 4023 1833
rect 4013 1563 4027 1567
rect 4036 1563 4043 1856
rect 4056 1607 4063 1873
rect 4076 1687 4083 2093
rect 4153 2083 4167 2087
rect 4176 2083 4183 2253
rect 4195 2227 4203 2353
rect 4215 2325 4223 2353
rect 4215 2227 4223 2311
rect 4235 2227 4243 2353
rect 4256 2347 4263 2533
rect 4276 2323 4283 3133
rect 4356 3107 4363 3213
rect 4296 2807 4303 3053
rect 4316 2964 4324 3076
rect 4296 2767 4303 2793
rect 4293 2753 4307 2767
rect 4313 2743 4327 2747
rect 4336 2743 4343 3093
rect 4356 3047 4363 3053
rect 4353 3033 4367 3047
rect 4376 3007 4383 3173
rect 4396 3067 4403 3213
rect 4416 3167 4423 3173
rect 4393 3043 4407 3047
rect 4416 3043 4423 3153
rect 4436 3107 4443 3356
rect 4476 3243 4483 3493
rect 4553 3483 4567 3487
rect 4576 3483 4583 3533
rect 4553 3476 4583 3483
rect 4553 3473 4567 3476
rect 4497 3278 4505 3302
rect 4467 3236 4483 3243
rect 4473 3223 4487 3227
rect 4456 3216 4487 3223
rect 4456 3127 4463 3216
rect 4473 3213 4487 3216
rect 4497 3184 4505 3264
rect 4393 3036 4423 3043
rect 4393 3033 4407 3036
rect 4313 2736 4343 2743
rect 4313 2733 4327 2736
rect 4295 2467 4303 2593
rect 4315 2509 4323 2593
rect 4315 2467 4323 2495
rect 4335 2467 4343 2593
rect 4356 2443 4363 2993
rect 4376 2547 4383 2873
rect 4416 2767 4423 2933
rect 4373 2533 4387 2547
rect 4413 2513 4427 2527
rect 4416 2447 4423 2513
rect 4336 2436 4363 2443
rect 4256 2316 4283 2323
rect 4256 2107 4263 2316
rect 4316 2307 4323 2433
rect 4313 2303 4327 2307
rect 4296 2296 4327 2303
rect 4153 2076 4183 2083
rect 4153 2073 4167 2076
rect 4096 1827 4103 1933
rect 4116 1847 4123 2033
rect 4136 1907 4143 2073
rect 4093 1813 4107 1827
rect 4156 1787 4163 1913
rect 4176 1887 4183 2076
rect 4053 1593 4067 1607
rect 4013 1556 4043 1563
rect 4013 1553 4027 1556
rect 4016 1487 4023 1553
rect 4076 1367 4083 1633
rect 4096 1327 4103 1693
rect 4136 1587 4143 1593
rect 4113 1553 4127 1567
rect 4133 1573 4147 1587
rect 4116 1527 4123 1553
rect 4176 1387 4183 1833
rect 4196 1783 4203 2053
rect 4216 2043 4223 2073
rect 4233 2043 4247 2047
rect 4216 2036 4247 2043
rect 4233 2033 4247 2036
rect 4273 2033 4287 2047
rect 4276 2027 4283 2033
rect 4296 1987 4303 2296
rect 4313 2293 4327 2296
rect 4336 2163 4343 2436
rect 4356 2287 4363 2393
rect 4376 2227 4383 2313
rect 4316 2156 4343 2163
rect 4296 1967 4303 1973
rect 4316 1927 4323 2156
rect 4416 2087 4423 2393
rect 4436 2327 4443 3033
rect 4455 2996 4463 3076
rect 4455 2958 4463 2982
rect 4456 2743 4463 2833
rect 4497 2798 4505 2822
rect 4473 2743 4487 2747
rect 4456 2736 4487 2743
rect 4456 2507 4463 2736
rect 4473 2733 4487 2736
rect 4497 2704 4505 2784
rect 4516 2667 4523 3453
rect 4556 3287 4563 3473
rect 4596 3387 4603 3676
rect 4616 3467 4623 3513
rect 4637 3476 4645 3556
rect 4637 3438 4645 3462
rect 4553 3213 4567 3227
rect 4556 3187 4563 3213
rect 4576 3207 4583 3273
rect 4576 3047 4583 3193
rect 4636 3184 4644 3296
rect 4656 3207 4663 3553
rect 4676 3547 4683 3593
rect 4676 3187 4683 3533
rect 4696 3527 4703 3533
rect 4736 3527 4743 3593
rect 4693 3513 4707 3527
rect 4733 3513 4747 3527
rect 4716 3223 4723 3273
rect 4756 3247 4763 3653
rect 4776 3607 4783 3693
rect 4776 3444 4784 3556
rect 4816 3447 4823 3853
rect 4836 3747 4843 4436
rect 4853 4433 4867 4436
rect 4853 4173 4867 4187
rect 4893 4183 4907 4187
rect 4916 4183 4923 4293
rect 4856 4167 4863 4173
rect 4893 4176 4923 4183
rect 4893 4173 4907 4176
rect 4856 3887 4863 4153
rect 4936 4107 4943 4393
rect 4916 3987 4923 4013
rect 4913 3973 4927 3987
rect 4896 3967 4903 3973
rect 4893 3953 4907 3967
rect 4836 3427 4843 3453
rect 4733 3223 4747 3227
rect 4716 3216 4747 3223
rect 4753 3233 4767 3247
rect 4793 3233 4807 3247
rect 4796 3227 4803 3233
rect 4733 3213 4747 3216
rect 4716 3067 4723 3093
rect 4716 3047 4723 3053
rect 4573 3033 4587 3047
rect 4593 3013 4607 3027
rect 4713 3033 4727 3047
rect 4536 2727 4543 3013
rect 4596 3003 4603 3013
rect 4576 2996 4603 3003
rect 4553 2733 4567 2747
rect 4556 2687 4563 2733
rect 4576 2627 4583 2996
rect 4616 2843 4623 2993
rect 4596 2836 4623 2843
rect 4596 2787 4603 2836
rect 4513 2543 4527 2547
rect 4473 2513 4487 2527
rect 4496 2536 4527 2543
rect 4456 2487 4463 2493
rect 4476 2447 4483 2513
rect 4496 2407 4503 2536
rect 4513 2533 4527 2536
rect 4557 2467 4565 2593
rect 4577 2509 4585 2593
rect 4577 2467 4585 2495
rect 4597 2467 4605 2593
rect 4436 2307 4443 2313
rect 4433 2293 4447 2307
rect 4453 2263 4467 2267
rect 4476 2263 4483 2293
rect 4453 2256 4483 2263
rect 4453 2253 4467 2256
rect 4456 2143 4463 2253
rect 4516 2147 4523 2453
rect 4616 2387 4623 2813
rect 4636 2704 4644 2816
rect 4696 2747 4703 3033
rect 4733 3013 4747 3027
rect 4776 3027 4783 3033
rect 4773 3013 4787 3027
rect 4736 2947 4743 3013
rect 4796 2967 4803 3193
rect 4816 3007 4823 3273
rect 4736 2704 4744 2816
rect 4636 2587 4643 2593
rect 4633 2573 4647 2587
rect 4655 2539 4663 2596
rect 4683 2557 4691 2596
rect 4655 2484 4663 2525
rect 4683 2484 4691 2543
rect 4716 2505 4724 2596
rect 4737 2481 4745 2596
rect 4755 2505 4763 2596
rect 4755 2466 4763 2491
rect 4796 2443 4803 2953
rect 4813 2733 4827 2747
rect 4816 2687 4823 2733
rect 4816 2547 4823 2673
rect 4813 2533 4827 2547
rect 4836 2467 4843 3413
rect 4776 2436 4803 2443
rect 4556 2287 4563 2313
rect 4533 2253 4547 2267
rect 4553 2273 4567 2287
rect 4573 2253 4587 2267
rect 4536 2207 4543 2253
rect 4576 2223 4583 2253
rect 4556 2216 4583 2223
rect 4436 2136 4463 2143
rect 4353 2063 4367 2067
rect 4336 2056 4367 2063
rect 4216 1867 4223 1893
rect 4276 1807 4283 1833
rect 4213 1783 4227 1787
rect 4196 1776 4227 1783
rect 4213 1773 4227 1776
rect 4273 1793 4287 1807
rect 4293 1773 4307 1787
rect 4296 1723 4303 1773
rect 4336 1767 4343 2056
rect 4353 2053 4367 2056
rect 4413 2073 4427 2087
rect 4436 2067 4443 2136
rect 4336 1747 4343 1753
rect 4296 1716 4323 1723
rect 4316 1683 4323 1716
rect 4336 1707 4343 1713
rect 4356 1683 4363 1833
rect 4376 1827 4383 1833
rect 4416 1827 4423 1913
rect 4456 1847 4463 2093
rect 4516 2087 4523 2093
rect 4556 2087 4563 2216
rect 4513 2073 4527 2087
rect 4373 1813 4387 1827
rect 4413 1823 4427 1827
rect 4393 1793 4407 1807
rect 4413 1816 4443 1823
rect 4413 1813 4427 1816
rect 4316 1676 4343 1683
rect 4356 1676 4383 1683
rect 4013 1313 4027 1327
rect 4016 1287 4023 1313
rect 4033 1293 4047 1307
rect 4073 1303 4087 1307
rect 4096 1303 4103 1313
rect 4073 1296 4103 1303
rect 4073 1293 4087 1296
rect 3953 1083 3967 1087
rect 3936 1076 3967 1083
rect 3993 1083 4007 1087
rect 4016 1083 4023 1133
rect 3953 1073 3967 1076
rect 3993 1076 4023 1083
rect 3993 1073 4007 1076
rect 3836 856 3863 863
rect 3816 647 3823 653
rect 3753 623 3767 627
rect 3736 616 3767 623
rect 3736 607 3743 616
rect 3753 613 3767 616
rect 3813 633 3827 647
rect 3736 407 3743 593
rect 3716 376 3743 383
rect 3573 356 3603 363
rect 3573 353 3587 356
rect 3653 363 3667 367
rect 3647 356 3667 363
rect 3653 353 3667 356
rect 3513 333 3527 336
rect 3553 333 3567 347
rect 3556 207 3563 333
rect 3636 323 3643 353
rect 3693 353 3707 367
rect 3636 316 3663 323
rect 3656 147 3663 316
rect 3673 313 3687 327
rect 3676 307 3683 313
rect 3736 187 3743 376
rect 3796 167 3803 393
rect 3816 387 3823 513
rect 3836 407 3843 833
rect 3856 767 3863 856
rect 3873 833 3887 847
rect 3856 643 3863 753
rect 3876 707 3883 833
rect 3933 823 3947 827
rect 3956 823 3963 1073
rect 3996 867 4003 893
rect 4036 883 4043 1293
rect 4073 1123 4087 1127
rect 4056 1116 4087 1123
rect 4056 1067 4063 1116
rect 4073 1113 4087 1116
rect 4136 887 4143 1353
rect 4173 1293 4187 1307
rect 4213 1293 4227 1307
rect 4176 1287 4183 1293
rect 4176 1143 4183 1273
rect 4216 1247 4223 1293
rect 4216 1207 4223 1233
rect 4193 1143 4207 1147
rect 4176 1136 4207 1143
rect 4193 1133 4207 1136
rect 4036 876 4063 883
rect 3993 853 4007 867
rect 3933 816 3963 823
rect 3933 813 3947 816
rect 3896 663 3903 713
rect 3887 656 3903 663
rect 3873 643 3887 647
rect 3856 636 3887 643
rect 3873 633 3887 636
rect 3936 627 3943 653
rect 3933 613 3947 627
rect 3856 427 3863 613
rect 3956 547 3963 816
rect 4056 807 4063 876
rect 3996 627 4003 793
rect 4036 667 4043 693
rect 4033 653 4047 667
rect 4076 647 4083 773
rect 4013 613 4027 627
rect 3813 373 3827 387
rect 3833 353 3847 367
rect 3873 353 3887 367
rect 3836 347 3843 353
rect 3876 347 3883 353
rect 3896 183 3903 413
rect 3916 367 3923 533
rect 4016 527 4023 613
rect 4096 403 4103 873
rect 4156 867 4163 1113
rect 4116 447 4123 853
rect 4176 847 4183 1113
rect 4213 1093 4227 1107
rect 4216 927 4223 1093
rect 4133 833 4147 847
rect 4136 807 4143 833
rect 4153 813 4167 827
rect 4156 407 4163 813
rect 4216 667 4223 913
rect 4236 907 4243 1673
rect 4296 1607 4303 1653
rect 4336 1607 4343 1676
rect 4293 1593 4307 1607
rect 4313 1573 4327 1587
rect 4316 1487 4323 1573
rect 4276 1287 4283 1473
rect 4356 1407 4363 1653
rect 4356 1327 4363 1393
rect 4353 1313 4367 1327
rect 4376 1187 4383 1676
rect 4396 1643 4403 1793
rect 4436 1787 4443 1816
rect 4496 1807 4503 1833
rect 4456 1707 4463 1793
rect 4493 1793 4507 1807
rect 4533 1793 4547 1807
rect 4513 1773 4527 1787
rect 4396 1636 4423 1643
rect 4416 1607 4423 1636
rect 4487 1616 4493 1623
rect 4456 1607 4463 1613
rect 4413 1593 4427 1607
rect 4453 1593 4467 1607
rect 4473 1573 4487 1587
rect 4476 1563 4483 1573
rect 4476 1556 4503 1563
rect 4476 1327 4483 1473
rect 4496 1347 4503 1556
rect 4433 1313 4447 1327
rect 4436 1267 4443 1313
rect 4473 1313 4487 1327
rect 4516 1307 4523 1773
rect 4536 1747 4543 1793
rect 4556 1787 4563 1833
rect 4556 1727 4563 1773
rect 4536 1387 4543 1613
rect 4556 1587 4563 1693
rect 4576 1607 4583 2193
rect 4596 1807 4603 2233
rect 4636 2167 4643 2313
rect 4653 2033 4667 2047
rect 4616 1707 4623 2013
rect 4656 2007 4663 2033
rect 4676 1847 4683 2353
rect 4696 2307 4703 2393
rect 4693 2293 4707 2307
rect 4713 2273 4727 2287
rect 4716 2267 4723 2273
rect 4653 1823 4667 1827
rect 4696 1823 4703 2093
rect 4716 2027 4723 2173
rect 4776 2107 4783 2436
rect 4773 2043 4787 2047
rect 4796 2043 4803 2393
rect 4856 2367 4863 3813
rect 4876 3727 4883 3733
rect 4873 3713 4887 3727
rect 4893 3703 4907 3707
rect 4916 3703 4923 3893
rect 4893 3696 4923 3703
rect 4893 3693 4907 3696
rect 4876 3227 4883 3673
rect 4896 3587 4903 3693
rect 4933 3473 4947 3487
rect 4936 3367 4943 3473
rect 4956 3287 4963 4653
rect 5056 4647 5063 4653
rect 5016 4487 5023 4613
rect 4993 4453 5007 4467
rect 5013 4473 5027 4487
rect 5076 4483 5083 4593
rect 5096 4527 5103 4816
rect 5116 4667 5123 4693
rect 5136 4547 5143 4913
rect 5176 4847 5183 5333
rect 5216 5327 5223 5613
rect 5236 5567 5243 5656
rect 5316 5647 5323 5653
rect 5313 5633 5327 5647
rect 5353 5633 5367 5647
rect 5333 5613 5347 5627
rect 5236 5487 5243 5553
rect 5236 5407 5243 5473
rect 5256 5447 5263 5513
rect 5253 5433 5267 5447
rect 5236 5387 5243 5393
rect 5193 5133 5207 5147
rect 5253 5163 5267 5167
rect 5276 5163 5283 5413
rect 5253 5156 5283 5163
rect 5253 5153 5267 5156
rect 5233 5133 5247 5147
rect 5196 5127 5203 5133
rect 5196 4963 5203 5093
rect 5236 5087 5243 5133
rect 5296 5023 5303 5193
rect 5276 5016 5303 5023
rect 5213 4963 5227 4967
rect 5196 4956 5227 4963
rect 5213 4953 5227 4956
rect 5216 4867 5223 4953
rect 5237 4916 5245 4996
rect 5237 4878 5245 4902
rect 5196 4707 5203 4713
rect 5193 4693 5207 4707
rect 5093 4483 5107 4487
rect 5076 4476 5107 4483
rect 5033 4463 5047 4467
rect 5033 4456 5063 4463
rect 5033 4453 5047 4456
rect 4996 4427 5003 4453
rect 4973 4153 4987 4167
rect 4976 4007 4983 4153
rect 4976 3383 4983 3493
rect 4996 3487 5003 4133
rect 5016 4027 5023 4433
rect 5056 4427 5063 4456
rect 5056 4167 5063 4213
rect 5013 4013 5027 4027
rect 5033 3983 5047 3987
rect 5027 3976 5047 3983
rect 5033 3973 5047 3976
rect 5016 3747 5023 3753
rect 5013 3733 5027 3747
rect 5076 3687 5083 4476
rect 5093 4473 5107 4476
rect 5117 4436 5125 4516
rect 5117 4398 5125 4422
rect 5136 4407 5143 4453
rect 5156 4227 5163 4513
rect 5176 4487 5183 4493
rect 5173 4473 5187 4487
rect 5196 4443 5203 4633
rect 5216 4527 5223 4733
rect 5236 4443 5243 4833
rect 5276 4747 5283 5016
rect 5296 4967 5303 4993
rect 5293 4953 5307 4967
rect 5316 4727 5323 5593
rect 5336 5523 5343 5613
rect 5356 5607 5363 5633
rect 5336 5516 5363 5523
rect 5336 5364 5344 5476
rect 5356 5207 5363 5516
rect 5333 5113 5347 5127
rect 5376 5123 5383 5613
rect 5356 5116 5383 5123
rect 5336 5107 5343 5113
rect 5336 4967 5343 5053
rect 5333 4953 5347 4967
rect 5256 4563 5263 4713
rect 5276 4707 5283 4713
rect 5273 4693 5287 4707
rect 5293 4673 5307 4687
rect 5296 4567 5303 4673
rect 5316 4607 5323 4653
rect 5336 4647 5343 4693
rect 5356 4647 5363 5116
rect 5376 4884 5384 4996
rect 5376 4727 5383 4773
rect 5376 4667 5383 4693
rect 5396 4607 5403 5773
rect 5456 5647 5463 5693
rect 5516 5663 5523 5823
rect 5556 5767 5563 5823
rect 5596 5787 5603 5823
rect 5636 5687 5643 5823
rect 5533 5663 5547 5667
rect 5516 5656 5547 5663
rect 5453 5633 5467 5647
rect 5516 5627 5523 5656
rect 5533 5653 5547 5656
rect 5553 5633 5567 5647
rect 5416 4707 5423 5573
rect 5436 5447 5443 5473
rect 5433 5433 5447 5447
rect 5453 5413 5467 5427
rect 5496 5427 5503 5433
rect 5493 5413 5507 5427
rect 5456 5367 5463 5413
rect 5433 5133 5447 5147
rect 5493 5153 5507 5167
rect 5436 4927 5443 5133
rect 5456 5067 5463 5113
rect 5436 4907 5443 4913
rect 5456 4787 5463 4973
rect 5256 4556 5283 4563
rect 5176 4436 5203 4443
rect 5216 4436 5243 4443
rect 5136 4207 5143 4213
rect 5133 4193 5147 4207
rect 5153 4183 5167 4187
rect 5176 4183 5183 4436
rect 5196 4407 5203 4413
rect 5196 4207 5203 4393
rect 5153 4176 5183 4183
rect 5153 4173 5167 4176
rect 5113 4153 5127 4167
rect 5116 4127 5123 4153
rect 5116 3987 5123 4093
rect 5176 4003 5183 4153
rect 5196 4047 5203 4193
rect 5216 4147 5223 4436
rect 5256 4404 5264 4516
rect 5276 4227 5283 4556
rect 5296 4527 5303 4533
rect 5296 4247 5303 4513
rect 5233 4173 5247 4187
rect 5273 4173 5287 4187
rect 5316 4183 5323 4593
rect 5296 4176 5323 4183
rect 5236 4107 5243 4173
rect 5276 4087 5283 4173
rect 5296 4067 5303 4176
rect 5193 4003 5207 4007
rect 5133 3973 5147 3987
rect 5176 3996 5207 4003
rect 5136 3967 5143 3973
rect 5036 3527 5043 3553
rect 5033 3513 5047 3527
rect 5053 3493 5067 3507
rect 5056 3467 5063 3493
rect 4976 3376 5003 3383
rect 4896 3267 4903 3273
rect 4893 3253 4907 3267
rect 4976 3227 4983 3353
rect 4996 3243 5003 3376
rect 5013 3243 5027 3247
rect 4996 3236 5027 3243
rect 5013 3233 5027 3236
rect 5033 3213 5047 3227
rect 4913 2993 4927 3007
rect 4916 2987 4923 2993
rect 4875 2798 4883 2822
rect 4875 2704 4883 2784
rect 4893 2743 4907 2747
rect 4893 2736 4923 2743
rect 4893 2733 4907 2736
rect 4916 2727 4923 2736
rect 4893 2533 4907 2547
rect 4816 2107 4823 2273
rect 4833 2253 4847 2267
rect 4836 2247 4843 2253
rect 4773 2036 4803 2043
rect 4773 2033 4787 2036
rect 4716 1867 4723 1873
rect 4653 1816 4703 1823
rect 4653 1813 4667 1816
rect 4616 1607 4623 1613
rect 4593 1573 4607 1587
rect 4613 1593 4627 1607
rect 4556 1327 4563 1553
rect 4596 1547 4603 1573
rect 4676 1347 4683 1816
rect 4693 1783 4707 1787
rect 4716 1783 4723 1853
rect 4736 1827 4743 2033
rect 4816 2027 4823 2093
rect 4693 1776 4723 1783
rect 4693 1773 4707 1776
rect 4493 1293 4507 1307
rect 4613 1293 4627 1307
rect 4436 1227 4443 1253
rect 4256 843 4263 1173
rect 4356 1147 4363 1153
rect 4373 1103 4387 1107
rect 4396 1103 4403 1153
rect 4373 1096 4403 1103
rect 4373 1093 4387 1096
rect 4416 1087 4423 1193
rect 4456 1107 4463 1133
rect 4476 1107 4483 1253
rect 4496 1167 4503 1293
rect 4536 1127 4543 1153
rect 4473 1093 4487 1107
rect 4533 1113 4547 1127
rect 4576 847 4583 1273
rect 4616 1147 4623 1293
rect 4656 1187 4663 1333
rect 4696 1287 4703 1753
rect 4736 1703 4743 1813
rect 4756 1767 4763 2013
rect 4796 1807 4803 1873
rect 4773 1773 4787 1787
rect 4776 1747 4783 1773
rect 4793 1753 4807 1767
rect 4716 1696 4743 1703
rect 4716 1347 4723 1696
rect 4776 1607 4783 1673
rect 4796 1647 4803 1753
rect 4756 1587 4763 1593
rect 4753 1573 4767 1587
rect 4773 1553 4787 1567
rect 4736 1507 4743 1553
rect 4776 1527 4783 1553
rect 4756 1347 4763 1413
rect 4753 1333 4767 1347
rect 4796 1287 4803 1613
rect 4816 1547 4823 1693
rect 4836 1667 4843 2233
rect 4856 2047 4863 2333
rect 4896 2327 4903 2533
rect 4896 2187 4903 2293
rect 4916 2287 4923 2713
rect 4936 2307 4943 3213
rect 4956 2787 4963 3213
rect 5036 3047 5043 3213
rect 5096 3203 5103 3933
rect 5136 3927 5143 3953
rect 5136 3727 5143 3793
rect 5133 3713 5147 3727
rect 5156 3707 5163 3753
rect 5156 3527 5163 3693
rect 5176 3587 5183 3996
rect 5193 3993 5207 3996
rect 5217 3956 5225 4036
rect 5217 3918 5225 3942
rect 5136 3467 5143 3513
rect 5193 3473 5207 3487
rect 5076 3196 5103 3203
rect 4996 3027 5003 3033
rect 4973 2993 4987 3007
rect 4993 3013 5007 3027
rect 4976 2987 4983 2993
rect 4956 2747 4963 2773
rect 4976 2723 4983 2753
rect 5033 2733 5047 2747
rect 4996 2727 5003 2733
rect 4956 2716 4983 2723
rect 4956 2287 4963 2716
rect 4976 2484 4984 2596
rect 5013 2563 5027 2567
rect 5036 2563 5043 2733
rect 5056 2567 5063 2673
rect 5013 2556 5043 2563
rect 5013 2553 5027 2556
rect 5053 2553 5067 2567
rect 4953 2273 4967 2287
rect 4976 2267 4983 2433
rect 5076 2347 5083 3196
rect 5096 2964 5104 3076
rect 5116 3067 5123 3453
rect 5156 3267 5163 3473
rect 5196 3467 5203 3473
rect 5173 3193 5187 3207
rect 5176 3067 5183 3193
rect 5116 3007 5123 3053
rect 5173 3043 5187 3047
rect 5173 3036 5203 3043
rect 5173 3033 5187 3036
rect 5196 3027 5203 3036
rect 5176 2787 5183 2973
rect 5115 2516 5123 2596
rect 5133 2553 5147 2567
rect 5115 2478 5123 2502
rect 5136 2447 5143 2553
rect 5033 2253 5047 2267
rect 5073 2253 5087 2267
rect 4956 2087 4963 2133
rect 4856 1627 4863 1833
rect 4876 1627 4883 2073
rect 4953 2073 4967 2087
rect 4976 1883 4983 2253
rect 5036 2207 5043 2253
rect 5036 2187 5043 2193
rect 4956 1876 4983 1883
rect 4896 1827 4903 1853
rect 4893 1813 4907 1827
rect 4853 1603 4867 1607
rect 4836 1596 4867 1603
rect 4836 1567 4843 1596
rect 4853 1593 4867 1596
rect 4873 1573 4887 1587
rect 4916 1587 4923 1733
rect 4913 1573 4927 1587
rect 4856 1407 4863 1553
rect 4876 1527 4883 1573
rect 4816 1303 4823 1393
rect 4856 1327 4863 1373
rect 4833 1303 4847 1307
rect 4816 1296 4847 1303
rect 4853 1313 4867 1327
rect 4833 1293 4847 1296
rect 4873 1293 4887 1307
rect 4796 1267 4803 1273
rect 4656 1147 4663 1173
rect 4653 1133 4667 1147
rect 4613 1123 4627 1127
rect 4596 1116 4627 1123
rect 4596 887 4603 1116
rect 4613 1113 4627 1116
rect 4633 1093 4647 1107
rect 4636 1087 4643 1093
rect 4656 883 4663 1093
rect 4696 1087 4703 1173
rect 4716 1147 4723 1153
rect 4716 1107 4723 1133
rect 4736 1127 4743 1133
rect 4733 1113 4747 1127
rect 4753 1093 4767 1107
rect 4796 1107 4803 1253
rect 4876 1207 4883 1293
rect 4873 1123 4887 1127
rect 4856 1116 4887 1123
rect 4793 1093 4807 1107
rect 4756 1087 4763 1093
rect 4727 1076 4743 1083
rect 4736 1063 4743 1076
rect 4816 1087 4823 1113
rect 4856 1087 4863 1116
rect 4873 1113 4887 1116
rect 4776 1063 4783 1073
rect 4736 1056 4783 1063
rect 4636 876 4663 883
rect 4273 843 4287 847
rect 4256 836 4287 843
rect 4256 827 4263 836
rect 4273 833 4287 836
rect 4293 813 4307 827
rect 4533 833 4547 847
rect 4333 813 4347 827
rect 4296 807 4303 813
rect 4336 767 4343 813
rect 4356 667 4363 673
rect 4353 653 4367 667
rect 4176 647 4183 653
rect 4173 633 4187 647
rect 4216 567 4223 593
rect 4076 396 4103 403
rect 3973 383 3987 387
rect 3973 376 4003 383
rect 3973 373 3987 376
rect 3996 347 4003 376
rect 4016 267 4023 353
rect 3876 176 3903 183
rect 3753 163 3767 167
rect 3753 156 3783 163
rect 3753 153 3767 156
rect 3633 113 3647 127
rect 3653 133 3667 147
rect 3636 107 3643 113
rect 3776 -17 3783 156
rect 3793 153 3807 167
rect 3876 -17 3883 176
rect 3893 163 3907 167
rect 3893 156 3923 163
rect 3893 153 3907 156
rect 3916 -17 3923 156
rect 4016 147 4023 253
rect 4033 123 4047 127
rect 4056 123 4063 193
rect 4076 167 4083 396
rect 4153 363 4167 367
rect 4176 363 4183 393
rect 4196 367 4203 433
rect 4216 396 4323 403
rect 4153 356 4183 363
rect 4153 353 4167 356
rect 4216 347 4223 396
rect 4233 353 4247 367
rect 4176 287 4183 313
rect 4236 307 4243 353
rect 4293 333 4307 347
rect 4296 303 4303 333
rect 4316 327 4323 396
rect 4376 367 4383 653
rect 4396 627 4403 833
rect 4516 747 4523 833
rect 4536 827 4543 833
rect 4553 813 4567 827
rect 4593 823 4607 827
rect 4616 823 4623 853
rect 4593 816 4623 823
rect 4593 813 4607 816
rect 4556 807 4563 813
rect 4436 647 4443 693
rect 4433 633 4447 647
rect 4596 647 4603 673
rect 4636 647 4643 876
rect 4656 847 4663 853
rect 4653 833 4667 847
rect 4713 813 4727 827
rect 4673 793 4687 807
rect 4676 747 4683 793
rect 4716 687 4723 813
rect 4736 807 4743 833
rect 4776 807 4783 853
rect 4593 633 4607 647
rect 4493 613 4507 627
rect 4656 627 4663 653
rect 4776 647 4783 753
rect 4796 667 4803 873
rect 4813 813 4827 827
rect 4853 813 4867 827
rect 4816 807 4823 813
rect 4856 787 4863 813
rect 4716 627 4723 633
rect 4713 613 4727 627
rect 4796 627 4803 653
rect 4836 627 4843 673
rect 4856 647 4863 693
rect 4876 667 4883 873
rect 4896 867 4903 1273
rect 4916 1127 4923 1133
rect 4913 1113 4927 1127
rect 4896 847 4903 853
rect 4916 787 4923 1073
rect 4936 887 4943 1613
rect 4956 1087 4963 1876
rect 4976 1807 4983 1833
rect 4996 1827 5003 2153
rect 5016 2087 5023 2113
rect 5056 2087 5063 2133
rect 5076 2127 5083 2253
rect 5136 2247 5143 2273
rect 5096 2087 5103 2113
rect 5053 2073 5067 2087
rect 5033 2063 5047 2067
rect 5016 2056 5047 2063
rect 5016 2027 5023 2056
rect 5033 2053 5047 2056
rect 5073 2053 5087 2067
rect 5093 2073 5107 2087
rect 5076 2047 5083 2053
rect 4996 1767 5003 1813
rect 5036 1807 5043 1833
rect 5076 1807 5083 1913
rect 5033 1793 5047 1807
rect 5073 1793 5087 1807
rect 5093 1773 5107 1787
rect 5016 1687 5023 1773
rect 5096 1767 5103 1773
rect 5016 1627 5023 1673
rect 5013 1603 5027 1607
rect 4996 1596 5027 1603
rect 4996 1527 5003 1596
rect 5013 1593 5027 1596
rect 5033 1553 5047 1567
rect 5036 1547 5043 1553
rect 4973 1293 4987 1307
rect 4976 1147 4983 1293
rect 5016 1287 5023 1293
rect 4993 1273 5007 1287
rect 4996 1247 5003 1273
rect 5013 1093 5027 1107
rect 5016 1067 5023 1093
rect 4993 823 5007 827
rect 5016 823 5023 953
rect 5036 907 5043 1453
rect 5056 967 5063 1753
rect 5116 1663 5123 2113
rect 5136 1807 5143 2233
rect 5156 2127 5163 2313
rect 5176 2107 5183 2733
rect 5196 2687 5203 3013
rect 5216 2707 5223 3873
rect 5236 3747 5243 4053
rect 5256 3807 5263 4033
rect 5316 4007 5323 4053
rect 5336 4007 5343 4493
rect 5356 4487 5363 4513
rect 5353 4473 5367 4487
rect 5373 4453 5387 4467
rect 5416 4467 5423 4633
rect 5413 4453 5427 4467
rect 5356 4127 5363 4433
rect 5376 4427 5383 4453
rect 5273 4003 5287 4007
rect 5273 3996 5293 4003
rect 5273 3993 5287 3996
rect 5313 3993 5327 4007
rect 5296 3727 5303 3993
rect 5356 3924 5364 4036
rect 5376 3727 5383 4133
rect 5396 3887 5403 4153
rect 5416 4047 5423 4413
rect 5436 4167 5443 4653
rect 5456 4087 5463 4633
rect 5476 4447 5483 5113
rect 5496 5107 5503 5153
rect 5516 5127 5523 5593
rect 5556 4987 5563 5633
rect 5576 5367 5583 5613
rect 5636 5483 5643 5653
rect 5653 5593 5667 5607
rect 5656 5587 5663 5593
rect 5636 5476 5663 5483
rect 5593 5393 5607 5407
rect 5596 5367 5603 5393
rect 5576 4967 5583 5193
rect 5596 5187 5603 5313
rect 5636 5187 5643 5353
rect 5593 5173 5607 5187
rect 5613 5153 5627 5167
rect 5616 4983 5623 5153
rect 5607 4976 5623 4983
rect 5556 4956 5573 4963
rect 5493 4913 5507 4927
rect 5533 4923 5547 4927
rect 5556 4923 5563 4956
rect 5533 4916 5563 4923
rect 5533 4913 5547 4916
rect 5496 4887 5503 4913
rect 5536 4727 5543 4893
rect 5576 4747 5583 4933
rect 5593 4913 5607 4927
rect 5596 4903 5603 4913
rect 5596 4896 5623 4903
rect 5596 4727 5603 4873
rect 5616 4807 5623 4896
rect 5656 4743 5663 5476
rect 5676 5407 5683 5533
rect 5696 5403 5703 5823
rect 5716 5467 5723 5633
rect 5736 5547 5743 5823
rect 5736 5427 5743 5433
rect 5713 5403 5727 5407
rect 5696 5396 5727 5403
rect 5733 5413 5747 5427
rect 5676 5207 5683 5393
rect 5696 5187 5703 5396
rect 5713 5393 5727 5396
rect 5753 5393 5767 5407
rect 5756 5387 5763 5393
rect 5716 5207 5723 5373
rect 5747 5196 5753 5203
rect 5693 5183 5707 5187
rect 5676 5176 5707 5183
rect 5733 5183 5747 5187
rect 5676 4927 5683 5176
rect 5693 5173 5707 5176
rect 5733 5176 5763 5183
rect 5733 5173 5747 5176
rect 5756 5147 5763 5176
rect 5636 4736 5663 4743
rect 5496 4527 5503 4713
rect 5533 4703 5547 4707
rect 5516 4696 5547 4703
rect 5573 4703 5587 4707
rect 5516 4627 5523 4696
rect 5533 4693 5547 4696
rect 5573 4696 5603 4703
rect 5573 4693 5587 4696
rect 5596 4667 5603 4696
rect 5513 4483 5527 4487
rect 5513 4476 5543 4483
rect 5513 4473 5527 4476
rect 5536 4407 5543 4476
rect 5553 4463 5567 4467
rect 5576 4463 5583 4653
rect 5553 4456 5583 4463
rect 5553 4453 5567 4456
rect 5533 4203 5547 4207
rect 5556 4203 5563 4293
rect 5533 4196 5563 4203
rect 5533 4193 5547 4196
rect 5576 4187 5583 4413
rect 5513 4173 5527 4187
rect 5416 4003 5423 4013
rect 5433 4003 5447 4007
rect 5416 3996 5447 4003
rect 5433 3993 5447 3996
rect 5416 3763 5423 3973
rect 5436 3827 5443 3993
rect 5457 3956 5465 4036
rect 5457 3918 5465 3942
rect 5396 3756 5423 3763
rect 5457 3758 5465 3782
rect 5373 3723 5387 3727
rect 5356 3716 5387 3723
rect 5356 3627 5363 3716
rect 5373 3713 5387 3716
rect 5236 3147 5243 3573
rect 5276 3444 5284 3556
rect 5316 3527 5323 3553
rect 5313 3513 5327 3527
rect 5296 3283 5303 3513
rect 5336 3523 5343 3533
rect 5353 3523 5367 3527
rect 5336 3516 5367 3523
rect 5296 3276 5323 3283
rect 5256 3267 5263 3273
rect 5253 3253 5267 3267
rect 5273 3233 5287 3247
rect 5276 3207 5283 3233
rect 5235 2996 5243 3076
rect 5235 2958 5243 2982
rect 5256 2767 5263 3033
rect 5316 2767 5323 3276
rect 5336 3023 5343 3516
rect 5353 3513 5367 3516
rect 5376 3487 5383 3533
rect 5353 3193 5367 3207
rect 5356 3067 5363 3193
rect 5353 3023 5367 3027
rect 5336 3016 5367 3023
rect 5353 3013 5367 3016
rect 5377 2798 5385 2822
rect 5253 2753 5267 2767
rect 5293 2763 5307 2767
rect 5276 2756 5307 2763
rect 5196 2327 5203 2473
rect 5276 2367 5283 2756
rect 5293 2753 5307 2756
rect 5316 2347 5323 2733
rect 5377 2704 5385 2784
rect 5196 2307 5203 2313
rect 5316 2307 5323 2333
rect 5193 2293 5207 2307
rect 5213 2273 5227 2287
rect 5216 2267 5223 2273
rect 5096 1656 5123 1663
rect 5076 1607 5083 1653
rect 5073 1593 5087 1607
rect 5076 1467 5083 1553
rect 5096 1427 5103 1656
rect 5116 1527 5123 1633
rect 5136 1387 5143 1773
rect 5156 1607 5163 2053
rect 5196 2047 5203 2093
rect 5193 1753 5207 1767
rect 5153 1583 5167 1587
rect 5176 1583 5183 1713
rect 5196 1687 5203 1753
rect 5196 1587 5203 1653
rect 5216 1647 5223 2193
rect 5236 2043 5243 2113
rect 5256 2087 5263 2293
rect 5276 2107 5283 2293
rect 5316 2287 5323 2293
rect 5313 2273 5327 2287
rect 5333 2253 5347 2267
rect 5293 2083 5307 2087
rect 5293 2076 5323 2083
rect 5293 2073 5307 2076
rect 5316 2067 5323 2076
rect 5236 2036 5263 2043
rect 5236 1747 5243 2013
rect 5256 1927 5263 2036
rect 5153 1576 5183 1583
rect 5153 1573 5167 1576
rect 5193 1573 5207 1587
rect 5213 1553 5227 1567
rect 5136 1347 5143 1353
rect 5133 1333 5147 1347
rect 5093 1143 5107 1147
rect 5076 1136 5107 1143
rect 5036 827 5043 853
rect 5056 847 5063 953
rect 5076 847 5083 1136
rect 5093 1133 5107 1136
rect 5113 1103 5127 1107
rect 5136 1103 5143 1173
rect 5113 1096 5143 1103
rect 5113 1093 5127 1096
rect 5096 847 5103 853
rect 5053 833 5067 847
rect 5093 833 5107 847
rect 4993 816 5023 823
rect 4993 813 5007 816
rect 5113 813 5127 827
rect 5116 807 5123 813
rect 4996 667 5003 673
rect 4993 653 5007 667
rect 4916 627 4923 653
rect 4913 613 4927 627
rect 4496 467 4503 613
rect 4516 387 4523 393
rect 4473 383 4487 387
rect 4456 376 4487 383
rect 4393 323 4407 327
rect 4416 323 4423 373
rect 4393 316 4423 323
rect 4393 313 4407 316
rect 4296 296 4323 303
rect 4096 127 4103 153
rect 4033 116 4063 123
rect 4033 113 4047 116
rect 4136 123 4143 193
rect 4176 167 4183 273
rect 4316 187 4323 296
rect 4313 173 4327 187
rect 4173 153 4187 167
rect 4336 167 4343 193
rect 4333 153 4347 167
rect 4416 147 4423 293
rect 4456 267 4463 376
rect 4473 373 4487 376
rect 4536 367 4543 453
rect 4593 353 4607 367
rect 4576 287 4583 353
rect 4596 347 4603 353
rect 4613 333 4627 347
rect 4653 343 4667 347
rect 4676 343 4683 353
rect 4653 336 4683 343
rect 4653 333 4667 336
rect 4616 327 4623 333
rect 4516 156 4573 163
rect 4153 123 4167 127
rect 4136 116 4167 123
rect 4153 113 4167 116
rect 4413 133 4427 147
rect 4433 123 4447 127
rect 4456 123 4463 133
rect 4516 127 4523 156
rect 4596 147 4603 213
rect 4616 147 4623 153
rect 4433 116 4463 123
rect 4433 113 4447 116
rect 4533 113 4547 127
rect 4593 133 4607 147
rect 4536 107 4543 113
rect 4636 107 4643 233
rect 4696 147 4703 213
rect 4756 167 4763 173
rect 4693 133 4707 147
rect 4733 133 4747 147
rect 4753 153 4767 167
rect 4736 123 4743 133
rect 4796 123 4803 493
rect 4816 387 4823 593
rect 4816 363 4823 373
rect 4876 367 4883 613
rect 4956 367 4963 653
rect 5013 613 5027 627
rect 5016 387 5023 613
rect 5096 487 5103 653
rect 5116 647 5123 773
rect 5136 667 5143 893
rect 5156 687 5163 1513
rect 5156 647 5163 653
rect 5113 633 5127 647
rect 5153 633 5167 647
rect 5136 427 5143 633
rect 4833 363 4847 367
rect 4816 356 4847 363
rect 4816 327 4823 356
rect 4833 353 4847 356
rect 4853 333 4867 347
rect 4873 353 4887 367
rect 5013 363 5027 367
rect 4973 333 4987 347
rect 4996 356 5027 363
rect 4856 247 4863 333
rect 4976 327 4983 333
rect 4813 123 4827 127
rect 4736 116 4827 123
rect 4853 123 4867 127
rect 4876 123 4883 153
rect 4956 147 4963 213
rect 4996 207 5003 356
rect 5013 353 5027 356
rect 5076 187 5083 393
rect 5156 387 5163 433
rect 5176 387 5183 1433
rect 5196 403 5203 1533
rect 5216 1527 5223 1553
rect 5236 1447 5243 1713
rect 5256 1667 5263 1853
rect 5296 1807 5303 1893
rect 5336 1867 5343 2253
rect 5356 2207 5363 2693
rect 5376 2107 5383 2313
rect 5396 2267 5403 3756
rect 5436 3707 5443 3713
rect 5433 3693 5447 3707
rect 5457 3664 5465 3744
rect 5415 3476 5423 3556
rect 5433 3513 5447 3527
rect 5415 3438 5423 3462
rect 5436 3447 5443 3513
rect 5436 3403 5443 3433
rect 5416 3396 5443 3403
rect 5416 2427 5423 3396
rect 5436 2847 5443 3373
rect 5456 2927 5463 3613
rect 5476 3387 5483 4113
rect 5496 3987 5503 4073
rect 5516 4067 5523 4173
rect 5516 4007 5523 4033
rect 5496 3487 5503 3733
rect 5536 3527 5543 4153
rect 5553 3693 5567 3707
rect 5556 3667 5563 3693
rect 5576 3527 5583 4173
rect 5596 4083 5603 4513
rect 5616 4307 5623 4733
rect 5616 4144 5624 4256
rect 5596 4076 5623 4083
rect 5596 3924 5604 4036
rect 5616 3787 5623 4076
rect 5596 3664 5604 3776
rect 5516 3287 5523 3493
rect 5573 3483 5587 3487
rect 5596 3483 5603 3513
rect 5573 3476 5603 3483
rect 5573 3473 5587 3476
rect 5576 3447 5583 3473
rect 5533 3243 5547 3247
rect 5556 3243 5563 3273
rect 5533 3236 5563 3243
rect 5533 3233 5547 3236
rect 5513 3213 5527 3227
rect 5516 3047 5523 3213
rect 5536 3043 5543 3053
rect 5553 3043 5567 3047
rect 5536 3036 5567 3043
rect 5553 3033 5567 3036
rect 5493 3013 5507 3027
rect 5496 2927 5503 3013
rect 5433 2733 5447 2747
rect 5436 2687 5443 2733
rect 5456 2547 5463 2913
rect 5496 2723 5503 2833
rect 5476 2716 5503 2723
rect 5416 2307 5423 2373
rect 5413 2293 5427 2307
rect 5433 2273 5447 2287
rect 5356 2043 5363 2073
rect 5396 2067 5403 2233
rect 5436 2127 5443 2273
rect 5373 2043 5387 2047
rect 5356 2036 5387 2043
rect 5393 2053 5407 2067
rect 5373 2033 5387 2036
rect 5413 2033 5427 2047
rect 5356 1847 5363 1853
rect 5313 1773 5327 1787
rect 5316 1767 5323 1773
rect 5293 1753 5307 1767
rect 5296 1743 5303 1753
rect 5296 1736 5313 1743
rect 5336 1687 5343 1833
rect 5376 1823 5383 2033
rect 5416 2027 5423 2033
rect 5356 1816 5383 1823
rect 5356 1767 5363 1816
rect 5396 1807 5403 1853
rect 5436 1847 5443 2093
rect 5393 1793 5407 1807
rect 5433 1793 5447 1807
rect 5376 1727 5383 1773
rect 5256 1547 5263 1633
rect 5276 1627 5283 1673
rect 5296 1607 5303 1653
rect 5376 1607 5383 1633
rect 5293 1593 5307 1607
rect 5216 1287 5223 1373
rect 5236 1347 5243 1413
rect 5256 1367 5263 1513
rect 5276 1363 5283 1593
rect 5373 1593 5387 1607
rect 5276 1356 5303 1363
rect 5233 1333 5247 1347
rect 5296 1267 5303 1356
rect 5316 1347 5323 1513
rect 5336 1467 5343 1553
rect 5396 1547 5403 1713
rect 5416 1507 5423 1753
rect 5436 1747 5443 1793
rect 5456 1727 5463 2253
rect 5476 2047 5483 2716
rect 5516 2704 5524 2816
rect 5536 2707 5543 2733
rect 5496 2107 5503 2373
rect 5556 2327 5563 3033
rect 5577 2996 5585 3076
rect 5577 2958 5585 2982
rect 5576 2523 5583 2913
rect 5596 2547 5603 3453
rect 5616 3267 5623 3733
rect 5636 3547 5643 4736
rect 5696 4727 5703 5133
rect 5716 4907 5723 5133
rect 5756 5107 5763 5113
rect 5756 4947 5763 4973
rect 5753 4933 5767 4947
rect 5773 4913 5787 4927
rect 5776 4907 5783 4913
rect 5656 4467 5663 4713
rect 5676 4707 5683 4713
rect 5673 4693 5687 4707
rect 5713 4693 5727 4707
rect 5693 4673 5707 4687
rect 5696 4667 5703 4673
rect 5716 4627 5723 4693
rect 5733 4683 5747 4687
rect 5756 4683 5763 4713
rect 5733 4676 5763 4683
rect 5733 4673 5747 4676
rect 5776 4667 5783 4793
rect 5713 4483 5727 4487
rect 5736 4483 5743 4653
rect 5653 4453 5667 4467
rect 5693 4453 5707 4467
rect 5713 4476 5743 4483
rect 5713 4473 5727 4476
rect 5696 4443 5703 4453
rect 5696 4436 5723 4443
rect 5676 4227 5683 4433
rect 5656 3947 5663 4153
rect 5676 4003 5683 4193
rect 5693 4173 5707 4187
rect 5696 4047 5703 4173
rect 5716 4147 5723 4436
rect 5736 4427 5743 4476
rect 5755 4238 5763 4262
rect 5755 4144 5763 4224
rect 5693 4003 5707 4007
rect 5676 3996 5707 4003
rect 5676 3927 5683 3996
rect 5693 3993 5707 3996
rect 5713 3973 5727 3987
rect 5716 3967 5723 3973
rect 5676 3527 5683 3653
rect 5673 3513 5687 3527
rect 5696 3507 5703 3773
rect 5716 3767 5723 3913
rect 5736 3767 5743 3953
rect 5716 3747 5723 3753
rect 5756 3747 5763 3933
rect 5713 3733 5727 3747
rect 5693 3493 5707 3507
rect 5716 3467 5723 3693
rect 5656 3267 5663 3433
rect 5653 3263 5667 3267
rect 5636 3256 5667 3263
rect 5636 3227 5643 3256
rect 5653 3253 5667 3256
rect 5673 3233 5687 3247
rect 5676 3063 5683 3233
rect 5676 3056 5703 3063
rect 5633 3043 5647 3047
rect 5616 3036 5647 3043
rect 5616 3027 5623 3036
rect 5633 3033 5647 3036
rect 5613 2733 5627 2747
rect 5673 2763 5687 2767
rect 5696 2763 5703 3056
rect 5716 2964 5724 3076
rect 5736 2927 5743 3493
rect 5673 2756 5703 2763
rect 5673 2753 5687 2756
rect 5653 2733 5667 2747
rect 5616 2727 5623 2733
rect 5656 2707 5663 2733
rect 5616 2543 5623 2673
rect 5633 2543 5647 2547
rect 5616 2536 5647 2543
rect 5633 2533 5647 2536
rect 5576 2516 5603 2523
rect 5516 2247 5523 2293
rect 5533 2233 5547 2247
rect 5536 2167 5543 2233
rect 5536 2147 5543 2153
rect 5493 2093 5507 2107
rect 5496 2056 5513 2063
rect 5436 1567 5443 1693
rect 5476 1667 5483 2013
rect 5496 1887 5503 2056
rect 5496 1807 5503 1873
rect 5476 1587 5483 1593
rect 5473 1573 5487 1587
rect 5316 1147 5323 1333
rect 5396 1327 5403 1333
rect 5373 1293 5387 1307
rect 5393 1313 5407 1327
rect 5413 1293 5427 1307
rect 5376 1167 5383 1293
rect 5416 1267 5423 1293
rect 5236 1107 5243 1133
rect 5213 1073 5227 1087
rect 5233 1093 5247 1107
rect 5253 1083 5267 1087
rect 5276 1083 5283 1113
rect 5253 1076 5283 1083
rect 5253 1073 5267 1076
rect 5216 847 5223 1073
rect 5213 833 5227 847
rect 5216 527 5223 673
rect 5196 396 5223 403
rect 5136 327 5143 353
rect 5096 187 5103 193
rect 5093 173 5107 187
rect 4813 113 4827 116
rect 4853 116 4883 123
rect 4953 133 4967 147
rect 5036 147 5043 173
rect 5076 167 5083 173
rect 5073 153 5087 167
rect 5196 123 5203 233
rect 5216 207 5223 396
rect 5236 367 5243 873
rect 5256 747 5263 793
rect 5276 687 5283 793
rect 5296 787 5303 1133
rect 5336 1123 5343 1153
rect 5416 1127 5423 1133
rect 5316 1116 5343 1123
rect 5316 887 5323 1116
rect 5353 1103 5367 1107
rect 5336 1096 5367 1103
rect 5316 827 5323 833
rect 5316 647 5323 813
rect 5336 807 5343 1096
rect 5353 1093 5367 1096
rect 5413 1113 5427 1127
rect 5416 827 5423 893
rect 5436 747 5443 1473
rect 5293 613 5307 627
rect 5313 633 5327 647
rect 5296 607 5303 613
rect 5336 607 5343 713
rect 5356 467 5363 693
rect 5376 647 5383 693
rect 5373 633 5387 647
rect 5436 627 5443 693
rect 5456 667 5463 1533
rect 5496 1347 5503 1533
rect 5516 1487 5523 2033
rect 5576 1807 5583 2273
rect 5596 2063 5603 2516
rect 5636 2287 5643 2333
rect 5633 2273 5647 2287
rect 5676 2243 5683 2733
rect 5733 2563 5747 2567
rect 5733 2556 5763 2563
rect 5733 2553 5747 2556
rect 5716 2307 5723 2533
rect 5713 2253 5727 2267
rect 5716 2247 5723 2253
rect 5656 2236 5683 2243
rect 5636 2107 5643 2233
rect 5633 2093 5647 2107
rect 5613 2063 5627 2067
rect 5596 2056 5627 2063
rect 5613 2053 5627 2056
rect 5553 1773 5567 1787
rect 5573 1793 5587 1807
rect 5593 1773 5607 1787
rect 5536 1627 5543 1773
rect 5536 1387 5543 1593
rect 5556 1567 5563 1773
rect 5596 1767 5603 1773
rect 5576 1647 5583 1733
rect 5576 1587 5583 1633
rect 5636 1627 5643 2053
rect 5656 2023 5663 2236
rect 5736 2207 5743 2273
rect 5676 2107 5683 2193
rect 5736 2163 5743 2173
rect 5756 2163 5763 2556
rect 5736 2156 5763 2163
rect 5736 2107 5743 2156
rect 5693 2083 5707 2087
rect 5676 2076 5707 2083
rect 5676 2047 5683 2076
rect 5693 2073 5707 2076
rect 5756 2067 5763 2133
rect 5753 2053 5767 2067
rect 5656 2016 5683 2023
rect 5633 1553 5647 1567
rect 5473 1293 5487 1307
rect 5533 1323 5547 1327
rect 5556 1323 5563 1353
rect 5533 1316 5563 1323
rect 5533 1313 5547 1316
rect 5513 1293 5527 1307
rect 5476 1187 5483 1293
rect 5476 1127 5483 1133
rect 5473 1113 5487 1127
rect 5516 1127 5523 1293
rect 5536 927 5543 1133
rect 5576 1087 5583 1393
rect 5596 1207 5603 1333
rect 5496 847 5503 913
rect 5536 847 5543 873
rect 5576 847 5583 1073
rect 5513 813 5527 827
rect 5533 833 5547 847
rect 5596 827 5603 1173
rect 5616 1127 5623 1533
rect 5636 1347 5643 1553
rect 5656 1407 5663 1593
rect 5676 1547 5683 2016
rect 5696 2003 5703 2033
rect 5716 2027 5723 2053
rect 5776 2047 5783 4133
rect 5696 1996 5723 2003
rect 5696 1807 5703 1973
rect 5693 1793 5707 1807
rect 5716 1643 5723 1996
rect 5696 1636 5723 1643
rect 5656 1327 5663 1373
rect 5696 1367 5703 1636
rect 5633 1293 5647 1307
rect 5653 1313 5667 1327
rect 5693 1313 5707 1327
rect 5673 1293 5687 1307
rect 5636 1287 5643 1293
rect 5636 1107 5643 1193
rect 5676 1187 5683 1293
rect 5676 1127 5683 1153
rect 5696 1107 5703 1313
rect 5716 1147 5723 1613
rect 5613 1073 5627 1087
rect 5633 1093 5647 1107
rect 5616 907 5623 1073
rect 5696 887 5703 1073
rect 5476 627 5483 733
rect 5433 613 5447 627
rect 5496 547 5503 773
rect 5236 167 5243 353
rect 5256 343 5263 453
rect 5296 367 5303 393
rect 5273 343 5287 347
rect 5256 336 5287 343
rect 5293 353 5307 367
rect 5273 333 5287 336
rect 5313 333 5327 347
rect 5316 227 5323 333
rect 5356 247 5363 413
rect 5376 347 5383 393
rect 5336 167 5343 193
rect 5396 167 5403 513
rect 5516 507 5523 813
rect 5596 707 5603 813
rect 5556 647 5563 673
rect 5596 647 5603 693
rect 5553 633 5567 647
rect 5536 627 5543 633
rect 5533 613 5547 627
rect 5416 327 5423 473
rect 5333 163 5347 167
rect 5213 123 5227 127
rect 5196 116 5227 123
rect 5296 143 5303 153
rect 5313 143 5327 147
rect 5296 136 5327 143
rect 5333 156 5363 163
rect 5333 153 5347 156
rect 5356 147 5363 156
rect 5313 133 5327 136
rect 5373 133 5387 147
rect 5393 153 5407 167
rect 5376 127 5383 133
rect 5436 127 5443 373
rect 5516 367 5523 393
rect 5453 333 5467 347
rect 5513 353 5527 367
rect 5456 187 5463 333
rect 5556 343 5563 393
rect 5596 367 5603 473
rect 5616 447 5623 853
rect 5656 847 5663 853
rect 5633 813 5647 827
rect 5653 833 5667 847
rect 5636 667 5643 813
rect 5616 387 5623 433
rect 5636 407 5643 653
rect 5656 647 5663 733
rect 5676 667 5683 713
rect 5673 653 5687 667
rect 5653 633 5667 647
rect 5716 603 5723 1093
rect 5736 607 5743 2033
rect 5756 1607 5763 1633
rect 5796 1607 5803 5693
rect 5816 3947 5823 5673
rect 5816 2147 5823 3813
rect 5753 1593 5767 1607
rect 5773 1573 5787 1587
rect 5776 1527 5783 1573
rect 5756 1167 5763 1353
rect 5776 1147 5783 1493
rect 5773 1133 5787 1147
rect 5696 596 5723 603
rect 5573 343 5587 347
rect 5556 336 5587 343
rect 5593 353 5607 367
rect 5573 333 5587 336
rect 5473 183 5487 187
rect 5467 176 5487 183
rect 5473 173 5487 176
rect 5656 147 5663 593
rect 5676 187 5683 533
rect 5696 147 5703 596
rect 5756 407 5763 873
rect 5716 387 5723 393
rect 5713 373 5727 387
rect 5753 383 5767 387
rect 5776 383 5783 1093
rect 5753 376 5783 383
rect 5753 373 5767 376
rect 5796 367 5803 1573
rect 4853 113 4867 116
rect 5213 113 5227 116
rect 5693 133 5707 147
rect 5713 123 5727 127
rect 5736 123 5743 173
rect 5713 116 5743 123
rect 5713 113 5727 116
rect 3476 -24 3503 -17
rect 3756 -24 3783 -17
rect 3856 -24 3883 -17
rect 3896 -24 3923 -17
<< m3contact >>
rect 453 5653 467 5667
rect 113 5633 127 5647
rect 133 5613 147 5627
rect 193 5613 207 5627
rect 213 5633 227 5647
rect 93 5473 107 5487
rect 73 5453 87 5467
rect 133 5453 147 5467
rect 93 5433 107 5447
rect 113 5413 127 5427
rect 373 5613 387 5627
rect 393 5633 407 5647
rect 413 5593 427 5607
rect 253 5533 267 5547
rect 393 5473 407 5487
rect 273 5433 287 5447
rect 193 5413 207 5427
rect 93 5393 107 5407
rect 53 5373 67 5387
rect 73 5373 87 5387
rect 53 5313 67 5327
rect 33 5013 47 5027
rect 33 4773 47 4787
rect 33 4673 47 4687
rect 93 5313 107 5327
rect 173 5233 187 5247
rect 153 5213 167 5227
rect 153 5173 167 5187
rect 93 5153 107 5167
rect 113 5153 127 5167
rect 73 4973 87 4987
rect 133 5113 147 5127
rect 113 4873 127 4887
rect 133 4833 147 4847
rect 113 4773 127 4787
rect 93 4753 107 4767
rect 113 4693 127 4707
rect 233 5233 247 5247
rect 233 5213 247 5227
rect 193 5173 207 5187
rect 353 5393 367 5407
rect 433 5413 447 5427
rect 413 5393 427 5407
rect 273 5173 287 5187
rect 313 5173 327 5187
rect 193 5153 207 5167
rect 213 5113 227 5127
rect 353 5153 367 5167
rect 513 5653 527 5667
rect 533 5633 547 5647
rect 493 5593 507 5607
rect 533 5593 547 5607
rect 693 5633 707 5647
rect 733 5633 747 5647
rect 653 5553 667 5567
rect 653 5533 667 5547
rect 533 5473 547 5487
rect 573 5473 587 5487
rect 413 5353 427 5367
rect 453 5353 467 5367
rect 393 5333 407 5347
rect 373 5013 387 5027
rect 373 4973 387 4987
rect 213 4953 227 4967
rect 573 5453 587 5467
rect 613 5433 627 5447
rect 493 5413 507 5427
rect 513 5393 527 5407
rect 593 5413 607 5427
rect 553 5393 567 5407
rect 493 5353 507 5367
rect 473 5333 487 5347
rect 533 5193 547 5207
rect 453 5173 467 5187
rect 433 5153 447 5167
rect 493 5173 507 5187
rect 473 5153 487 5167
rect 413 5133 427 5147
rect 413 4973 427 4987
rect 393 4953 407 4967
rect 193 4933 207 4947
rect 213 4913 227 4927
rect 233 4933 247 4947
rect 293 4933 307 4947
rect 333 4933 347 4947
rect 253 4913 267 4927
rect 213 4893 227 4907
rect 313 4913 327 4927
rect 353 4913 367 4927
rect 393 4913 407 4927
rect 293 4893 307 4907
rect 193 4833 207 4847
rect 173 4773 187 4787
rect 153 4753 167 4767
rect 153 4713 167 4727
rect 53 4493 67 4507
rect 113 4633 127 4647
rect 133 4573 147 4587
rect 93 4493 107 4507
rect 153 4493 167 4507
rect 33 4173 47 4187
rect 73 4453 87 4467
rect 113 4453 127 4467
rect 73 4413 87 4427
rect 193 4713 207 4727
rect 293 4873 307 4887
rect 233 4673 247 4687
rect 193 4633 207 4647
rect 233 4633 247 4647
rect 273 4673 287 4687
rect 273 4653 287 4667
rect 253 4613 267 4627
rect 233 4553 247 4567
rect 173 4433 187 4447
rect 53 4113 67 4127
rect 53 4093 67 4107
rect 113 4173 127 4187
rect 133 4193 147 4207
rect 173 4173 187 4187
rect 133 4153 147 4167
rect 113 4113 127 4127
rect 93 4093 107 4107
rect 73 4013 87 4027
rect 93 4013 107 4027
rect 93 3973 107 3987
rect 53 3773 67 3787
rect 13 3133 27 3147
rect 13 3013 27 3027
rect 33 1573 47 1587
rect 13 1553 27 1567
rect 13 1493 27 1507
rect 33 1133 47 1147
rect 173 4153 187 4167
rect 153 4073 167 4087
rect 153 4033 167 4047
rect 253 4493 267 4507
rect 213 4433 227 4447
rect 313 4773 327 4787
rect 373 4713 387 4727
rect 413 4753 427 4767
rect 393 4693 407 4707
rect 373 4673 387 4687
rect 313 4633 327 4647
rect 353 4633 367 4647
rect 353 4613 367 4627
rect 413 4553 427 4567
rect 353 4493 367 4507
rect 293 4473 307 4487
rect 273 4453 287 4467
rect 253 4433 267 4447
rect 213 4193 227 4207
rect 253 4173 267 4187
rect 273 4193 287 4207
rect 233 4153 247 4167
rect 213 4133 227 4147
rect 253 4133 267 4147
rect 233 4113 247 4127
rect 193 4033 207 4047
rect 173 4013 187 4027
rect 153 3993 167 4007
rect 133 3953 147 3967
rect 113 3773 127 3787
rect 113 3753 127 3767
rect 73 3733 87 3747
rect 73 3693 87 3707
rect 133 3693 147 3707
rect 93 3593 107 3607
rect 93 3573 107 3587
rect 133 3553 147 3567
rect 73 3493 87 3507
rect 113 3493 127 3507
rect 133 3513 147 3527
rect 133 3453 147 3467
rect 93 3433 107 3447
rect 113 3433 127 3447
rect 73 3253 87 3267
rect 93 3233 107 3247
rect 93 3193 107 3207
rect 133 3213 147 3227
rect 73 3173 87 3187
rect 113 3173 127 3187
rect 193 3973 207 3987
rect 213 3993 227 4007
rect 293 4073 307 4087
rect 293 4033 307 4047
rect 253 3973 267 3987
rect 173 3953 187 3967
rect 333 4453 347 4467
rect 373 4453 387 4467
rect 393 4473 407 4487
rect 413 4453 427 4467
rect 333 4433 347 4447
rect 393 4433 407 4447
rect 333 4413 347 4427
rect 373 4253 387 4267
rect 333 4173 347 4187
rect 353 4053 367 4067
rect 333 3973 347 3987
rect 193 3733 207 3747
rect 233 3733 247 3747
rect 313 3733 327 3747
rect 293 3713 307 3727
rect 213 3693 227 3707
rect 253 3693 267 3707
rect 213 3593 227 3607
rect 273 3573 287 3587
rect 293 3573 307 3587
rect 213 3533 227 3547
rect 193 3493 207 3507
rect 233 3493 247 3507
rect 253 3513 267 3527
rect 293 3513 307 3527
rect 273 3493 287 3507
rect 173 3453 187 3467
rect 253 3273 267 3287
rect 173 3233 187 3247
rect 173 3213 187 3227
rect 213 3233 227 3247
rect 233 3213 247 3227
rect 113 2993 127 3007
rect 73 2973 87 2987
rect 113 2973 127 2987
rect 73 2793 87 2807
rect 93 2753 107 2767
rect 113 2773 127 2787
rect 93 2733 107 2747
rect 113 2733 127 2747
rect 113 2513 127 2527
rect 73 2293 87 2307
rect 93 2273 107 2287
rect 73 2253 87 2267
rect 73 2113 87 2127
rect 113 2153 127 2167
rect 153 3033 167 3047
rect 273 3253 287 3267
rect 273 3213 287 3227
rect 253 3193 267 3207
rect 253 3033 267 3047
rect 213 2993 227 3007
rect 333 3693 347 3707
rect 513 5133 527 5147
rect 493 5093 507 5107
rect 573 5153 587 5167
rect 713 5573 727 5587
rect 693 5473 707 5487
rect 833 5653 847 5667
rect 1333 5653 1347 5667
rect 893 5633 907 5647
rect 773 5613 787 5627
rect 933 5633 947 5647
rect 913 5593 927 5607
rect 993 5593 1007 5607
rect 893 5573 907 5587
rect 793 5553 807 5567
rect 813 5553 827 5567
rect 773 5453 787 5467
rect 1213 5633 1227 5647
rect 1253 5613 1267 5627
rect 1073 5593 1087 5607
rect 1053 5533 1067 5547
rect 673 5413 687 5427
rect 673 5393 687 5407
rect 733 5413 747 5427
rect 813 5413 827 5427
rect 833 5433 847 5447
rect 953 5433 967 5447
rect 853 5413 867 5427
rect 913 5413 927 5427
rect 933 5413 947 5427
rect 713 5353 727 5367
rect 613 5213 627 5227
rect 613 5173 627 5187
rect 793 5173 807 5187
rect 733 5133 747 5147
rect 753 5153 767 5167
rect 533 5113 547 5127
rect 593 5113 607 5127
rect 1273 5593 1287 5607
rect 1093 5573 1107 5587
rect 1113 5573 1127 5587
rect 1133 5453 1147 5467
rect 1173 5453 1187 5467
rect 973 5413 987 5427
rect 1073 5413 1087 5427
rect 1153 5413 1167 5427
rect 993 5193 1007 5207
rect 873 5153 887 5167
rect 893 5153 907 5167
rect 1013 5173 1027 5187
rect 1053 5173 1067 5187
rect 813 5133 827 5147
rect 853 5133 867 5147
rect 773 5113 787 5127
rect 853 5113 867 5127
rect 733 5093 747 5107
rect 753 5093 767 5107
rect 573 4953 587 4967
rect 633 4953 647 4967
rect 693 4953 707 4967
rect 553 4933 567 4947
rect 493 4873 507 4887
rect 553 4833 567 4847
rect 453 4753 467 4767
rect 493 4673 507 4687
rect 513 4693 527 4707
rect 453 4653 467 4667
rect 453 4633 467 4647
rect 533 4653 547 4667
rect 513 4593 527 4607
rect 493 4573 507 4587
rect 493 4533 507 4547
rect 453 4433 467 4447
rect 433 4253 447 4267
rect 413 4113 427 4127
rect 453 4193 467 4207
rect 653 4933 667 4947
rect 673 4913 687 4927
rect 593 4893 607 4907
rect 633 4893 647 4907
rect 573 4533 587 4547
rect 573 4513 587 4527
rect 613 4693 627 4707
rect 653 4673 667 4687
rect 633 4533 647 4547
rect 653 4533 667 4547
rect 553 4453 567 4467
rect 593 4473 607 4487
rect 693 4553 707 4567
rect 713 4513 727 4527
rect 673 4493 687 4507
rect 673 4473 687 4487
rect 693 4453 707 4467
rect 713 4473 727 4487
rect 533 4433 547 4447
rect 433 4093 447 4107
rect 453 4093 467 4107
rect 413 4053 427 4067
rect 473 3973 487 3987
rect 413 3713 427 3727
rect 493 3713 507 3727
rect 433 3693 447 3707
rect 453 3693 467 3707
rect 373 3553 387 3567
rect 373 3533 387 3547
rect 413 3573 427 3587
rect 393 3493 407 3507
rect 493 3553 507 3567
rect 453 3493 467 3507
rect 473 3513 487 3527
rect 773 4953 787 4967
rect 793 4933 807 4947
rect 813 4953 827 4967
rect 773 4913 787 4927
rect 793 4673 807 4687
rect 913 5133 927 5147
rect 893 5113 907 5127
rect 1033 5093 1047 5107
rect 953 4973 967 4987
rect 993 4973 1007 4987
rect 1073 5153 1087 5167
rect 1293 5433 1307 5447
rect 1173 5393 1187 5407
rect 1253 5413 1267 5427
rect 1233 5393 1247 5407
rect 1153 5373 1167 5387
rect 1153 5153 1167 5167
rect 1133 5113 1147 5127
rect 1133 5093 1147 5107
rect 1113 5073 1127 5087
rect 893 4953 907 4967
rect 933 4933 947 4947
rect 993 4933 1007 4947
rect 1053 4933 1067 4947
rect 1113 4953 1127 4967
rect 1013 4713 1027 4727
rect 873 4653 887 4667
rect 833 4593 847 4607
rect 893 4593 907 4607
rect 1013 4673 1027 4687
rect 1093 4873 1107 4887
rect 1053 4633 1067 4647
rect 993 4553 1007 4567
rect 853 4533 867 4547
rect 933 4533 947 4547
rect 773 4493 787 4507
rect 813 4493 827 4507
rect 793 4453 807 4467
rect 893 4513 907 4527
rect 893 4493 907 4507
rect 913 4453 927 4467
rect 933 4473 947 4487
rect 1013 4473 1027 4487
rect 993 4453 1007 4467
rect 893 4293 907 4307
rect 593 4193 607 4207
rect 573 4153 587 4167
rect 573 4133 587 4147
rect 553 4113 567 4127
rect 733 4193 747 4207
rect 753 4193 767 4207
rect 813 4193 827 4207
rect 653 4113 667 4127
rect 633 4093 647 4107
rect 593 4053 607 4067
rect 553 4033 567 4047
rect 613 4033 627 4047
rect 593 3993 607 4007
rect 733 4093 747 4107
rect 833 4173 847 4187
rect 853 4193 867 4207
rect 813 4153 827 4167
rect 553 3973 567 3987
rect 713 3993 727 4007
rect 873 4033 887 4047
rect 733 3973 747 3987
rect 833 3973 847 3987
rect 853 3993 867 4007
rect 713 3953 727 3967
rect 653 3733 667 3747
rect 533 3693 547 3707
rect 553 3693 567 3707
rect 593 3713 607 3727
rect 613 3673 627 3687
rect 573 3653 587 3667
rect 613 3533 627 3547
rect 593 3513 607 3527
rect 553 3473 567 3487
rect 353 3293 367 3307
rect 413 3293 427 3307
rect 313 3273 327 3287
rect 313 3253 327 3267
rect 313 3233 327 3247
rect 393 3273 407 3287
rect 413 3233 427 3247
rect 393 3213 407 3227
rect 453 3213 467 3227
rect 393 3073 407 3087
rect 353 3053 367 3067
rect 293 3033 307 3047
rect 473 3033 487 3047
rect 253 2993 267 3007
rect 313 3013 327 3027
rect 413 2993 427 3007
rect 213 2973 227 2987
rect 373 2973 387 2987
rect 253 2793 267 2807
rect 153 2733 167 2747
rect 213 2733 227 2747
rect 193 2713 207 2727
rect 173 2653 187 2667
rect 153 2593 167 2607
rect 173 2533 187 2547
rect 173 2513 187 2527
rect 153 2433 167 2447
rect 153 2253 167 2267
rect 113 1993 127 2007
rect 113 1813 127 1827
rect 93 1793 107 1807
rect 133 1773 147 1787
rect 113 1753 127 1767
rect 133 1693 147 1707
rect 73 1633 87 1647
rect 113 1573 127 1587
rect 93 1553 107 1567
rect 133 1553 147 1567
rect 113 1533 127 1547
rect 73 1513 87 1527
rect 113 1413 127 1427
rect 93 1313 107 1327
rect 113 1233 127 1247
rect 133 1213 147 1227
rect 93 1173 107 1187
rect 233 2573 247 2587
rect 473 2893 487 2907
rect 553 3433 567 3447
rect 593 3433 607 3447
rect 553 3253 567 3267
rect 513 3233 527 3247
rect 573 3113 587 3127
rect 573 3053 587 3067
rect 533 3033 547 3047
rect 513 3013 527 3027
rect 553 3013 567 3027
rect 733 3733 747 3747
rect 713 3693 727 3707
rect 733 3693 747 3707
rect 813 3713 827 3727
rect 853 3713 867 3727
rect 913 4193 927 4207
rect 913 4153 927 4167
rect 933 4153 947 4167
rect 953 4033 967 4047
rect 973 4013 987 4027
rect 913 3993 927 4007
rect 713 3633 727 3647
rect 673 3573 687 3587
rect 653 3293 667 3307
rect 673 3293 687 3307
rect 693 3253 707 3267
rect 713 3213 727 3227
rect 633 3173 647 3187
rect 633 3053 647 3067
rect 673 3053 687 3067
rect 613 3033 627 3047
rect 593 2933 607 2947
rect 373 2773 387 2787
rect 333 2753 347 2767
rect 273 2653 287 2667
rect 353 2653 367 2667
rect 493 2813 507 2827
rect 413 2753 427 2767
rect 453 2753 467 2767
rect 493 2733 507 2747
rect 393 2713 407 2727
rect 473 2713 487 2727
rect 433 2693 447 2707
rect 373 2593 387 2607
rect 293 2533 307 2547
rect 333 2533 347 2547
rect 473 2573 487 2587
rect 393 2553 407 2567
rect 373 2533 387 2547
rect 273 2513 287 2527
rect 353 2513 367 2527
rect 253 2433 267 2447
rect 233 2293 247 2307
rect 213 2273 227 2287
rect 193 2093 207 2107
rect 193 2033 207 2047
rect 253 2253 267 2267
rect 293 2313 307 2327
rect 353 2313 367 2327
rect 313 2293 327 2307
rect 333 2273 347 2287
rect 293 2253 307 2267
rect 313 2253 327 2267
rect 273 2093 287 2107
rect 293 2093 307 2107
rect 233 2033 247 2047
rect 253 2053 267 2067
rect 293 2053 307 2067
rect 213 1853 227 1867
rect 193 1833 207 1847
rect 293 2013 307 2027
rect 273 1953 287 1967
rect 213 1813 227 1827
rect 233 1813 247 1827
rect 193 1793 207 1807
rect 233 1793 247 1807
rect 213 1753 227 1767
rect 213 1733 227 1747
rect 193 1673 207 1687
rect 253 1713 267 1727
rect 433 2533 447 2547
rect 413 2513 427 2527
rect 413 2273 427 2287
rect 373 2233 387 2247
rect 333 2193 347 2207
rect 433 2253 447 2267
rect 453 2273 467 2287
rect 413 2173 427 2187
rect 373 2093 387 2107
rect 393 2053 407 2067
rect 413 2073 427 2087
rect 353 2013 367 2027
rect 413 2013 427 2027
rect 333 1953 347 1967
rect 373 1933 387 1947
rect 333 1833 347 1847
rect 393 1873 407 1887
rect 373 1813 387 1827
rect 413 1813 427 1827
rect 293 1673 307 1687
rect 313 1613 327 1627
rect 273 1593 287 1607
rect 213 1553 227 1567
rect 253 1573 267 1587
rect 273 1573 287 1587
rect 193 1533 207 1547
rect 233 1533 247 1547
rect 293 1473 307 1487
rect 193 1333 207 1347
rect 193 1313 207 1327
rect 233 1313 247 1327
rect 273 1313 287 1327
rect 253 1293 267 1307
rect 173 1253 187 1267
rect 233 1253 247 1267
rect 213 1213 227 1227
rect 213 1153 227 1167
rect 73 1093 87 1107
rect 73 1073 87 1087
rect 173 1133 187 1147
rect 153 1093 167 1107
rect 193 1093 207 1107
rect 133 873 147 887
rect 173 873 187 887
rect 93 833 107 847
rect 133 833 147 847
rect 113 793 127 807
rect 133 713 147 727
rect 153 653 167 667
rect 113 633 127 647
rect 53 613 67 627
rect 33 593 47 607
rect 73 593 87 607
rect 93 613 107 627
rect 73 573 87 587
rect 153 573 167 587
rect 153 533 167 547
rect 93 353 107 367
rect 113 333 127 347
rect 93 153 107 167
rect 153 173 167 187
rect 73 113 87 127
rect 113 133 127 147
rect 133 133 147 147
rect 113 113 127 127
rect 273 1233 287 1247
rect 313 1453 327 1467
rect 313 1413 327 1427
rect 313 1253 327 1267
rect 293 1153 307 1167
rect 353 1773 367 1787
rect 373 1773 387 1787
rect 413 1753 427 1767
rect 413 1733 427 1747
rect 353 1713 367 1727
rect 373 1613 387 1627
rect 353 1573 367 1587
rect 373 1573 387 1587
rect 353 1533 367 1547
rect 393 1553 407 1567
rect 373 1513 387 1527
rect 393 1473 407 1487
rect 353 1453 367 1467
rect 393 1313 407 1327
rect 373 1273 387 1287
rect 373 1253 387 1267
rect 273 1093 287 1107
rect 353 1113 367 1127
rect 393 1113 407 1127
rect 373 1093 387 1107
rect 233 853 247 867
rect 193 833 207 847
rect 253 813 267 827
rect 313 1073 327 1087
rect 473 2233 487 2247
rect 493 2233 507 2247
rect 653 3013 667 3027
rect 833 3693 847 3707
rect 893 3693 907 3707
rect 773 3673 787 3687
rect 893 3573 907 3587
rect 973 3953 987 3967
rect 1033 4453 1047 4467
rect 1073 4433 1087 4447
rect 1153 5073 1167 5087
rect 1253 5373 1267 5387
rect 1293 5173 1307 5187
rect 1273 5093 1287 5107
rect 1493 5653 1507 5667
rect 1513 5633 1527 5647
rect 1373 5613 1387 5627
rect 1393 5613 1407 5627
rect 1353 5573 1367 5587
rect 1633 5653 1647 5667
rect 1553 5613 1567 5627
rect 1413 5593 1427 5607
rect 1533 5593 1547 5607
rect 1393 5533 1407 5547
rect 1373 5493 1387 5507
rect 1353 5433 1367 5447
rect 1673 5633 1687 5647
rect 1613 5473 1627 5487
rect 1633 5473 1647 5487
rect 1413 5433 1427 5447
rect 1553 5433 1567 5447
rect 1593 5433 1607 5447
rect 1533 5413 1547 5427
rect 1533 5373 1547 5387
rect 1353 5153 1367 5167
rect 1413 5153 1427 5167
rect 1333 5133 1347 5147
rect 1313 5113 1327 5127
rect 1353 5113 1367 5127
rect 1233 4973 1247 4987
rect 1293 4973 1307 4987
rect 1333 4973 1347 4987
rect 1173 4953 1187 4967
rect 1213 4933 1227 4947
rect 1153 4673 1167 4687
rect 1133 4633 1147 4647
rect 1313 4933 1327 4947
rect 1293 4773 1307 4787
rect 1433 5133 1447 5147
rect 1453 5153 1467 5167
rect 1413 5013 1427 5027
rect 1393 4933 1407 4947
rect 1353 4733 1367 4747
rect 1433 4933 1447 4947
rect 1453 4913 1467 4927
rect 1413 4893 1427 4907
rect 1513 5153 1527 5167
rect 1493 4913 1507 4927
rect 1473 4873 1487 4887
rect 1213 4673 1227 4687
rect 1233 4653 1247 4667
rect 1253 4673 1267 4687
rect 1353 4673 1367 4687
rect 1213 4633 1227 4647
rect 1253 4633 1267 4647
rect 1173 4493 1187 4507
rect 1173 4473 1187 4487
rect 1153 4453 1167 4467
rect 1193 4453 1207 4467
rect 1093 4413 1107 4427
rect 1033 4213 1047 4227
rect 1153 4413 1167 4427
rect 1073 4193 1087 4207
rect 1133 4193 1147 4207
rect 1053 4153 1067 4167
rect 1093 4113 1107 4127
rect 1093 4013 1107 4027
rect 1073 3953 1087 3967
rect 1093 3853 1107 3867
rect 1073 3813 1087 3827
rect 1033 3793 1047 3807
rect 953 3753 967 3767
rect 1013 3753 1027 3767
rect 993 3733 1007 3747
rect 1013 3693 1027 3707
rect 1173 4233 1187 4247
rect 1313 4613 1327 4627
rect 1273 4533 1287 4547
rect 1273 4493 1287 4507
rect 1313 4493 1327 4507
rect 1333 4453 1347 4467
rect 1373 4633 1387 4647
rect 1373 4573 1387 4587
rect 1293 4433 1307 4447
rect 1353 4433 1367 4447
rect 1353 4353 1367 4367
rect 1253 4253 1267 4267
rect 1293 4253 1307 4267
rect 1313 4253 1327 4267
rect 1213 4213 1227 4227
rect 1253 4213 1267 4227
rect 1233 4193 1247 4207
rect 1193 4153 1207 4167
rect 1293 4213 1307 4227
rect 1273 4173 1287 4187
rect 1253 4113 1267 4127
rect 1233 4073 1247 4087
rect 1273 4013 1287 4027
rect 1153 3933 1167 3947
rect 1213 3953 1227 3967
rect 1173 3813 1187 3827
rect 1393 4533 1407 4547
rect 1433 4713 1447 4727
rect 1493 4673 1507 4687
rect 1553 5273 1567 5287
rect 1593 5273 1607 5287
rect 1753 5633 1767 5647
rect 1733 5613 1747 5627
rect 1693 5593 1707 5607
rect 1693 5473 1707 5487
rect 1653 5453 1667 5467
rect 1633 5433 1647 5447
rect 1653 5413 1667 5427
rect 1673 5433 1687 5447
rect 1733 5453 1747 5467
rect 1533 5133 1547 5147
rect 1693 5173 1707 5187
rect 1773 5593 1787 5607
rect 1933 5653 1947 5667
rect 2073 5653 2087 5667
rect 2113 5653 2127 5667
rect 2033 5633 2047 5647
rect 1873 5613 1887 5627
rect 1833 5593 1847 5607
rect 1853 5593 1867 5607
rect 1913 5593 1927 5607
rect 1813 5553 1827 5567
rect 1773 5413 1787 5427
rect 1573 4973 1587 4987
rect 1533 4913 1547 4927
rect 1653 5153 1667 5167
rect 1633 4913 1647 4927
rect 1553 4893 1567 4907
rect 1553 4693 1567 4707
rect 1593 4693 1607 4707
rect 1533 4673 1547 4687
rect 1573 4673 1587 4687
rect 1633 4693 1647 4707
rect 1513 4633 1527 4647
rect 1473 4613 1487 4627
rect 1433 4573 1447 4587
rect 1433 4533 1447 4547
rect 1453 4473 1467 4487
rect 1413 4453 1427 4467
rect 1433 4453 1447 4467
rect 1373 4233 1387 4247
rect 1353 4213 1367 4227
rect 1373 4193 1387 4207
rect 1353 4173 1367 4187
rect 1333 4013 1347 4027
rect 1313 3953 1327 3967
rect 1313 3933 1327 3947
rect 1293 3893 1307 3907
rect 1253 3853 1267 3867
rect 1293 3833 1307 3847
rect 1213 3793 1227 3807
rect 1113 3753 1127 3767
rect 1173 3753 1187 3767
rect 1113 3733 1127 3747
rect 1153 3733 1167 3747
rect 1133 3693 1147 3707
rect 1013 3673 1027 3687
rect 1093 3673 1107 3687
rect 973 3573 987 3587
rect 953 3533 967 3547
rect 1113 3553 1127 3567
rect 1053 3533 1067 3547
rect 913 3513 927 3527
rect 933 3493 947 3507
rect 913 3473 927 3487
rect 793 3453 807 3467
rect 893 3453 907 3467
rect 813 3433 827 3447
rect 873 3433 887 3447
rect 753 3213 767 3227
rect 833 3293 847 3307
rect 873 3253 887 3267
rect 773 3033 787 3047
rect 653 2993 667 3007
rect 653 2953 667 2967
rect 533 2753 547 2767
rect 593 2753 607 2767
rect 613 2773 627 2787
rect 553 2733 567 2747
rect 573 2733 587 2747
rect 533 2673 547 2687
rect 533 2573 547 2587
rect 553 2533 567 2547
rect 533 2233 547 2247
rect 453 2213 467 2227
rect 513 2213 527 2227
rect 433 1293 447 1307
rect 473 2173 487 2187
rect 733 3013 747 3027
rect 753 3013 767 3027
rect 793 3013 807 3027
rect 813 3033 827 3047
rect 873 3193 887 3207
rect 853 3153 867 3167
rect 853 3093 867 3107
rect 833 3013 847 3027
rect 793 2993 807 3007
rect 753 2973 767 2987
rect 713 2933 727 2947
rect 713 2773 727 2787
rect 653 2753 667 2767
rect 673 2733 687 2747
rect 733 2733 747 2747
rect 773 2793 787 2807
rect 853 2813 867 2827
rect 813 2793 827 2807
rect 793 2773 807 2787
rect 833 2753 847 2767
rect 773 2733 787 2747
rect 753 2713 767 2727
rect 633 2693 647 2707
rect 733 2693 747 2707
rect 673 2673 687 2687
rect 713 2673 727 2687
rect 633 2653 647 2667
rect 653 2573 667 2587
rect 673 2553 687 2567
rect 673 2293 687 2307
rect 573 2213 587 2227
rect 633 2273 647 2287
rect 653 2233 667 2247
rect 633 2213 647 2227
rect 593 2193 607 2207
rect 613 2193 627 2207
rect 573 2133 587 2147
rect 473 2053 487 2067
rect 513 2033 527 2047
rect 513 1873 527 1887
rect 493 1833 507 1847
rect 513 1833 527 1847
rect 533 1813 547 1827
rect 473 1733 487 1747
rect 513 1733 527 1747
rect 513 1713 527 1727
rect 553 1793 567 1807
rect 553 1773 567 1787
rect 553 1713 567 1727
rect 613 2073 627 2087
rect 673 2073 687 2087
rect 913 3253 927 3267
rect 913 3213 927 3227
rect 993 3493 1007 3507
rect 1033 3493 1047 3507
rect 953 3433 967 3447
rect 1033 3353 1047 3367
rect 953 3253 967 3267
rect 993 3253 1007 3267
rect 973 3193 987 3207
rect 973 3173 987 3187
rect 933 3153 947 3167
rect 993 3153 1007 3167
rect 933 3013 947 3027
rect 953 3033 967 3047
rect 973 3013 987 3027
rect 1033 3133 1047 3147
rect 1013 3073 1027 3087
rect 893 2793 907 2807
rect 893 2773 907 2787
rect 933 2773 947 2787
rect 933 2753 947 2767
rect 993 2733 1007 2747
rect 893 2713 907 2727
rect 953 2713 967 2727
rect 873 2673 887 2687
rect 793 2593 807 2607
rect 753 2573 767 2587
rect 873 2573 887 2587
rect 733 2533 747 2547
rect 773 2533 787 2547
rect 813 2553 827 2567
rect 873 2533 887 2547
rect 933 2693 947 2707
rect 993 2593 1007 2607
rect 913 2533 927 2547
rect 933 2533 947 2547
rect 973 2553 987 2567
rect 753 2433 767 2447
rect 893 2433 907 2447
rect 773 2193 787 2207
rect 893 2293 907 2307
rect 813 2273 827 2287
rect 853 2273 867 2287
rect 793 2113 807 2127
rect 793 2093 807 2107
rect 753 2073 767 2087
rect 973 2513 987 2527
rect 953 2253 967 2267
rect 913 2133 927 2147
rect 913 2113 927 2127
rect 893 2093 907 2107
rect 833 2073 847 2087
rect 813 2053 827 2067
rect 773 2033 787 2047
rect 713 2013 727 2027
rect 813 2013 827 2027
rect 653 1933 667 1947
rect 713 1853 727 1867
rect 713 1833 727 1847
rect 593 1793 607 1807
rect 573 1633 587 1647
rect 553 1613 567 1627
rect 493 1573 507 1587
rect 533 1573 547 1587
rect 613 1633 627 1647
rect 593 1553 607 1567
rect 473 1333 487 1347
rect 533 1333 547 1347
rect 493 1313 507 1327
rect 513 1293 527 1307
rect 533 1313 547 1327
rect 573 1313 587 1327
rect 553 1293 567 1307
rect 553 1273 567 1287
rect 453 1253 467 1267
rect 513 1253 527 1267
rect 533 1253 547 1267
rect 473 1233 487 1247
rect 433 1173 447 1187
rect 433 1133 447 1147
rect 493 1093 507 1107
rect 453 1073 467 1087
rect 353 1013 367 1027
rect 393 1013 407 1027
rect 413 1013 427 1027
rect 533 1213 547 1227
rect 533 1073 547 1087
rect 473 953 487 967
rect 513 953 527 967
rect 373 833 387 847
rect 313 813 327 827
rect 433 853 447 867
rect 213 793 227 807
rect 233 793 247 807
rect 273 793 287 807
rect 333 793 347 807
rect 373 793 387 807
rect 393 793 407 807
rect 273 653 287 667
rect 253 613 267 627
rect 293 613 307 627
rect 313 613 327 627
rect 293 413 307 427
rect 213 353 227 367
rect 253 353 267 367
rect 293 353 307 367
rect 253 313 267 327
rect 213 173 227 187
rect 173 153 187 167
rect 313 333 327 347
rect 293 313 307 327
rect 353 713 367 727
rect 453 653 467 667
rect 393 613 407 627
rect 413 593 427 607
rect 453 533 467 547
rect 413 373 427 387
rect 373 333 387 347
rect 413 353 427 367
rect 453 353 467 367
rect 433 313 447 327
rect 333 293 347 307
rect 393 293 407 307
rect 273 253 287 267
rect 373 253 387 267
rect 413 193 427 207
rect 193 133 207 147
rect 393 133 407 147
rect 693 1773 707 1787
rect 853 2033 867 2047
rect 913 2053 927 2067
rect 893 2033 907 2047
rect 713 1753 727 1767
rect 833 1793 847 1807
rect 813 1773 827 1787
rect 773 1753 787 1767
rect 933 2013 947 2027
rect 953 2013 967 2027
rect 953 1813 967 1827
rect 933 1793 947 1807
rect 993 2413 1007 2427
rect 1033 3013 1047 3027
rect 1033 2913 1047 2927
rect 1093 3513 1107 3527
rect 1153 3513 1167 3527
rect 1193 3733 1207 3747
rect 1253 3733 1267 3747
rect 1233 3713 1247 3727
rect 1193 3613 1207 3627
rect 1213 3613 1227 3627
rect 1173 3473 1187 3487
rect 1093 3453 1107 3467
rect 1073 3313 1087 3327
rect 1173 3273 1187 3287
rect 1093 3253 1107 3267
rect 1113 3233 1127 3247
rect 1173 3213 1187 3227
rect 1133 3173 1147 3187
rect 1173 3133 1187 3147
rect 1133 3113 1147 3127
rect 1073 3093 1087 3107
rect 1093 3013 1107 3027
rect 1073 2973 1087 2987
rect 1093 2973 1107 2987
rect 1113 2953 1127 2967
rect 1073 2773 1087 2787
rect 1093 2573 1107 2587
rect 1153 3073 1167 3087
rect 1173 3053 1187 3067
rect 1153 2993 1167 3007
rect 1153 2933 1167 2947
rect 1153 2833 1167 2847
rect 1093 2553 1107 2567
rect 1033 2513 1047 2527
rect 1013 2293 1027 2307
rect 1113 2533 1127 2547
rect 1333 3753 1347 3767
rect 1393 3993 1407 4007
rect 1433 4193 1447 4207
rect 1533 4513 1547 4527
rect 1493 4473 1507 4487
rect 1553 4473 1567 4487
rect 1513 4413 1527 4427
rect 1553 4413 1567 4427
rect 1473 4333 1487 4347
rect 1513 4233 1527 4247
rect 1473 4213 1487 4227
rect 1533 4193 1547 4207
rect 1373 3933 1387 3947
rect 1393 3753 1407 3767
rect 1333 3733 1347 3747
rect 1313 3633 1327 3647
rect 1273 3613 1287 3627
rect 1333 3513 1347 3527
rect 1253 3473 1267 3487
rect 1273 3493 1287 3507
rect 1333 3493 1347 3507
rect 1293 3453 1307 3467
rect 1233 3313 1247 3327
rect 1293 3433 1307 3447
rect 1213 3253 1227 3267
rect 1253 3273 1267 3287
rect 1213 3233 1227 3247
rect 1233 3233 1247 3247
rect 1253 3233 1267 3247
rect 1233 3173 1247 3187
rect 1213 3153 1227 3167
rect 1233 3133 1247 3147
rect 1453 3993 1467 4007
rect 1433 3733 1447 3747
rect 1373 3713 1387 3727
rect 1393 3713 1407 3727
rect 1413 3713 1427 3727
rect 1453 3713 1467 3727
rect 1433 3693 1447 3707
rect 1393 3653 1407 3667
rect 1373 3633 1387 3647
rect 1373 3593 1387 3607
rect 1353 3473 1367 3487
rect 1413 3513 1427 3527
rect 1393 3473 1407 3487
rect 1453 3493 1467 3507
rect 1433 3473 1447 3487
rect 1413 3453 1427 3467
rect 1373 3433 1387 3447
rect 1353 3293 1367 3307
rect 1333 3133 1347 3147
rect 1293 3113 1307 3127
rect 1273 3053 1287 3067
rect 1313 3053 1327 3067
rect 1373 3233 1387 3247
rect 1393 3113 1407 3127
rect 1293 3033 1307 3047
rect 1273 2953 1287 2967
rect 1333 3013 1347 3027
rect 1613 4653 1627 4667
rect 1593 4633 1607 4647
rect 1593 4613 1607 4627
rect 1593 4413 1607 4427
rect 1673 5133 1687 5147
rect 1753 5153 1767 5167
rect 1713 5133 1727 5147
rect 1753 5133 1767 5147
rect 1693 5113 1707 5127
rect 1713 4973 1727 4987
rect 1793 5393 1807 5407
rect 1813 5413 1827 5427
rect 1913 5573 1927 5587
rect 1853 5453 1867 5467
rect 1973 5473 1987 5487
rect 1953 5433 1967 5447
rect 2373 5653 2387 5667
rect 2453 5653 2467 5667
rect 2133 5633 2147 5647
rect 2113 5593 2127 5607
rect 2053 5453 2067 5467
rect 2093 5453 2107 5467
rect 1973 5393 1987 5407
rect 1893 5173 1907 5187
rect 1913 5173 1927 5187
rect 2033 5413 2047 5427
rect 2013 5373 2027 5387
rect 2013 5213 2027 5227
rect 1993 5193 2007 5207
rect 1793 5153 1807 5167
rect 1833 5153 1847 5167
rect 1773 5113 1787 5127
rect 1773 5033 1787 5047
rect 1733 4933 1747 4947
rect 1873 5113 1887 5127
rect 1933 5133 1947 5147
rect 1913 5033 1927 5047
rect 1833 4973 1847 4987
rect 1773 4933 1787 4947
rect 1793 4933 1807 4947
rect 1853 4933 1867 4947
rect 1873 4953 1887 4967
rect 1913 4953 1927 4967
rect 2053 5393 2067 5407
rect 2073 5413 2087 5427
rect 2093 5393 2107 5407
rect 2093 5373 2107 5387
rect 2033 5193 2047 5207
rect 2093 5193 2107 5207
rect 2053 5173 2067 5187
rect 2173 5633 2187 5647
rect 2213 5613 2227 5627
rect 2153 5593 2167 5607
rect 2193 5593 2207 5607
rect 2333 5633 2347 5647
rect 2413 5633 2427 5647
rect 2473 5633 2487 5647
rect 2313 5573 2327 5587
rect 2273 5553 2287 5567
rect 2313 5553 2327 5567
rect 2233 5453 2247 5467
rect 2373 5533 2387 5547
rect 2613 5653 2627 5667
rect 2593 5633 2607 5647
rect 2713 5653 2727 5667
rect 2633 5633 2647 5647
rect 2693 5633 2707 5647
rect 2753 5653 2767 5667
rect 2793 5653 2807 5667
rect 2553 5473 2567 5487
rect 2413 5453 2427 5467
rect 2493 5453 2507 5467
rect 2513 5453 2527 5467
rect 2173 5293 2187 5307
rect 2333 5293 2347 5307
rect 2193 5213 2207 5227
rect 2213 5193 2227 5207
rect 2393 5193 2407 5207
rect 2073 5133 2087 5147
rect 2133 5153 2147 5167
rect 2193 5153 2207 5167
rect 2313 5173 2327 5187
rect 2273 5153 2287 5167
rect 2353 5173 2367 5187
rect 2333 5153 2347 5167
rect 2113 5093 2127 5107
rect 2153 5093 2167 5107
rect 2093 5033 2107 5047
rect 1893 4933 1907 4947
rect 1813 4913 1827 4927
rect 1673 4893 1687 4907
rect 1853 4893 1867 4907
rect 1813 4793 1827 4807
rect 1713 4693 1727 4707
rect 1713 4653 1727 4667
rect 1773 4673 1787 4687
rect 1793 4653 1807 4667
rect 1713 4633 1727 4647
rect 1673 4593 1687 4607
rect 1653 4513 1667 4527
rect 1833 4573 1847 4587
rect 1713 4453 1727 4467
rect 1693 4393 1707 4407
rect 1673 4273 1687 4287
rect 1653 4213 1667 4227
rect 1613 4193 1627 4207
rect 1593 4173 1607 4187
rect 1553 4113 1567 4127
rect 1493 4033 1507 4047
rect 1533 4033 1547 4047
rect 1553 4033 1567 4047
rect 1553 3933 1567 3947
rect 1533 3753 1547 3767
rect 1513 3733 1527 3747
rect 1493 3713 1507 3727
rect 1513 3693 1527 3707
rect 1573 3713 1587 3727
rect 1553 3693 1567 3707
rect 1493 3673 1507 3687
rect 1613 4153 1627 4167
rect 1753 4533 1767 4547
rect 1813 4533 1827 4547
rect 1793 4493 1807 4507
rect 1833 4453 1847 4467
rect 1813 4433 1827 4447
rect 1793 4413 1807 4427
rect 1733 4253 1747 4267
rect 1873 4713 1887 4727
rect 1913 4913 1927 4927
rect 1953 4913 1967 4927
rect 1973 4933 1987 4947
rect 2133 4973 2147 4987
rect 2113 4933 2127 4947
rect 2473 5433 2487 5447
rect 2553 5433 2567 5447
rect 2593 5433 2607 5447
rect 2673 5433 2687 5447
rect 2413 5133 2427 5147
rect 2373 5113 2387 5127
rect 2353 5053 2367 5067
rect 2553 5373 2567 5387
rect 2553 5193 2567 5207
rect 2473 5173 2487 5187
rect 2453 5133 2467 5147
rect 2513 5153 2527 5167
rect 2493 5113 2507 5127
rect 2433 5033 2447 5047
rect 2433 5013 2447 5027
rect 2373 4973 2387 4987
rect 2193 4933 2207 4947
rect 2253 4933 2267 4947
rect 2393 4933 2407 4947
rect 2413 4953 2427 4967
rect 2153 4913 2167 4927
rect 1813 4373 1827 4387
rect 1853 4373 1867 4387
rect 1673 4173 1687 4187
rect 1613 4113 1627 4127
rect 1633 4113 1647 4127
rect 1633 4013 1647 4027
rect 1653 4013 1667 4027
rect 1613 3993 1627 4007
rect 1633 3973 1647 3987
rect 1553 3633 1567 3647
rect 1593 3633 1607 3647
rect 1593 3613 1607 3627
rect 1473 3393 1487 3407
rect 1533 3493 1547 3507
rect 1573 3493 1587 3507
rect 1493 3273 1507 3287
rect 1553 3273 1567 3287
rect 1473 3253 1487 3267
rect 1433 3233 1447 3247
rect 1413 2993 1427 3007
rect 1393 2913 1407 2927
rect 1293 2813 1307 2827
rect 1313 2773 1327 2787
rect 1193 2673 1207 2687
rect 1273 2753 1287 2767
rect 1333 2753 1347 2767
rect 1313 2733 1327 2747
rect 1233 2653 1247 2667
rect 1173 2593 1187 2607
rect 1173 2573 1187 2587
rect 1093 2393 1107 2407
rect 1033 2233 1047 2247
rect 1073 2233 1087 2247
rect 1113 2293 1127 2307
rect 1053 2213 1067 2227
rect 1093 2213 1107 2227
rect 1153 2253 1167 2267
rect 993 2053 1007 2067
rect 973 1773 987 1787
rect 1113 2073 1127 2087
rect 1133 2073 1147 2087
rect 1053 2033 1067 2047
rect 1073 2053 1087 2067
rect 1093 2033 1107 2047
rect 1013 1873 1027 1887
rect 1133 1833 1147 1847
rect 1033 1793 1047 1807
rect 993 1753 1007 1767
rect 1033 1753 1047 1767
rect 853 1733 867 1747
rect 953 1733 967 1747
rect 733 1693 747 1707
rect 693 1613 707 1627
rect 733 1613 747 1627
rect 753 1613 767 1627
rect 633 1553 647 1567
rect 933 1653 947 1667
rect 893 1613 907 1627
rect 873 1593 887 1607
rect 773 1573 787 1587
rect 853 1573 867 1587
rect 913 1573 927 1587
rect 753 1533 767 1547
rect 633 1293 647 1307
rect 673 1313 687 1327
rect 653 1253 667 1267
rect 653 1153 667 1167
rect 613 1133 627 1147
rect 613 1113 627 1127
rect 673 1133 687 1147
rect 593 1073 607 1087
rect 633 1073 647 1087
rect 973 1613 987 1627
rect 973 1573 987 1587
rect 953 1513 967 1527
rect 813 1353 827 1367
rect 913 1353 927 1367
rect 873 1333 887 1347
rect 793 1293 807 1307
rect 953 1333 967 1347
rect 773 1153 787 1167
rect 933 1153 947 1167
rect 1093 1793 1107 1807
rect 1113 1773 1127 1787
rect 1053 1733 1067 1747
rect 1033 1593 1047 1607
rect 1133 1753 1147 1767
rect 1133 1673 1147 1687
rect 1093 1653 1107 1667
rect 1033 1573 1047 1587
rect 1013 1353 1027 1367
rect 1053 1313 1067 1327
rect 1373 2753 1387 2767
rect 1413 2753 1427 2767
rect 1393 2733 1407 2747
rect 1333 2713 1347 2727
rect 1293 2693 1307 2707
rect 1353 2653 1367 2667
rect 1193 2533 1207 2547
rect 1233 2533 1247 2547
rect 1273 2513 1287 2527
rect 1353 2513 1367 2527
rect 1213 2493 1227 2507
rect 1333 2493 1347 2507
rect 1193 2433 1207 2447
rect 1173 2213 1187 2227
rect 1413 2553 1427 2567
rect 1413 2533 1427 2547
rect 1393 2333 1407 2347
rect 1573 3253 1587 3267
rect 1513 3213 1527 3227
rect 1493 3193 1507 3207
rect 1553 3193 1567 3207
rect 1533 3113 1547 3127
rect 1493 3073 1507 3087
rect 1513 3053 1527 3067
rect 1473 2993 1487 3007
rect 1533 3013 1547 3027
rect 1613 3493 1627 3507
rect 1613 3473 1627 3487
rect 1753 4213 1767 4227
rect 1793 4213 1807 4227
rect 1773 4193 1787 4207
rect 1733 4173 1747 4187
rect 1853 4273 1867 4287
rect 1833 4253 1847 4267
rect 1713 4153 1727 4167
rect 1813 4153 1827 4167
rect 1693 4133 1707 4147
rect 1693 3973 1707 3987
rect 1673 3853 1687 3867
rect 1673 3733 1687 3747
rect 1653 3673 1667 3687
rect 1813 4033 1827 4047
rect 1753 4013 1767 4027
rect 2113 4773 2127 4787
rect 1953 4653 1967 4667
rect 1993 4673 2007 4687
rect 2073 4673 2087 4687
rect 1933 4553 1947 4567
rect 2033 4633 2047 4647
rect 1973 4513 1987 4527
rect 2013 4513 2027 4527
rect 1913 4473 1927 4487
rect 1933 4453 1947 4467
rect 2013 4473 2027 4487
rect 2033 4473 2047 4487
rect 2053 4453 2067 4467
rect 2093 4653 2107 4667
rect 2093 4573 2107 4587
rect 2073 4433 2087 4447
rect 2053 4413 2067 4427
rect 1893 4253 1907 4267
rect 1933 4253 1947 4267
rect 1873 4173 1887 4187
rect 1833 4013 1847 4027
rect 1933 4193 1947 4207
rect 1893 4153 1907 4167
rect 1873 3993 1887 4007
rect 1853 3973 1867 3987
rect 1893 3973 1907 3987
rect 1813 3753 1827 3767
rect 1873 3753 1887 3767
rect 1893 3753 1907 3767
rect 1733 3713 1747 3727
rect 1873 3733 1887 3747
rect 1893 3713 1907 3727
rect 1753 3693 1767 3707
rect 1753 3573 1767 3587
rect 1713 3553 1727 3567
rect 1653 3533 1667 3547
rect 1713 3533 1727 3547
rect 1673 3513 1687 3527
rect 1653 3473 1667 3487
rect 1693 3473 1707 3487
rect 1633 3453 1647 3467
rect 1613 3253 1627 3267
rect 1593 3233 1607 3247
rect 1653 3253 1667 3267
rect 1633 3233 1647 3247
rect 1773 3493 1787 3507
rect 1753 3453 1767 3467
rect 1733 3273 1747 3287
rect 1773 3293 1787 3307
rect 1713 3233 1727 3247
rect 1673 3213 1687 3227
rect 1613 3133 1627 3147
rect 1593 3093 1607 3107
rect 1573 3053 1587 3067
rect 1553 2973 1567 2987
rect 1493 2953 1507 2967
rect 1473 2753 1487 2767
rect 1513 2753 1527 2767
rect 1493 2733 1507 2747
rect 1553 2733 1567 2747
rect 1673 3053 1687 3067
rect 1633 3033 1647 3047
rect 1653 3013 1667 3027
rect 2133 4733 2147 4747
rect 2413 4733 2427 4747
rect 2233 4713 2247 4727
rect 2193 4653 2207 4667
rect 2173 4633 2187 4647
rect 2173 4533 2187 4547
rect 2213 4493 2227 4507
rect 2173 4473 2187 4487
rect 2213 4473 2227 4487
rect 2153 4453 2167 4467
rect 2253 4653 2267 4667
rect 2273 4653 2287 4667
rect 2353 4673 2367 4687
rect 2393 4673 2407 4687
rect 2453 4953 2467 4967
rect 2433 4673 2447 4687
rect 2393 4653 2407 4667
rect 2313 4613 2327 4627
rect 2273 4553 2287 4567
rect 2213 4313 2227 4327
rect 2153 4273 2167 4287
rect 2193 4273 2207 4287
rect 2093 4253 2107 4267
rect 2113 4253 2127 4267
rect 2053 4233 2067 4247
rect 1973 4193 1987 4207
rect 2013 4193 2027 4207
rect 2033 4213 2047 4227
rect 2073 4213 2087 4227
rect 2053 4173 2067 4187
rect 1993 4153 2007 4167
rect 1973 4093 1987 4107
rect 2053 4093 2067 4107
rect 1993 4053 2007 4067
rect 2033 4053 2047 4067
rect 1973 3973 1987 3987
rect 1973 3933 1987 3947
rect 2013 3933 2027 3947
rect 1953 3693 1967 3707
rect 2173 4233 2187 4247
rect 2133 4213 2147 4227
rect 2093 4173 2107 4187
rect 2113 4173 2127 4187
rect 2073 3973 2087 3987
rect 2053 3793 2067 3807
rect 2073 3793 2087 3807
rect 1993 3753 2007 3767
rect 2033 3733 2047 3747
rect 2053 3733 2067 3747
rect 1993 3713 2007 3727
rect 1973 3673 1987 3687
rect 2033 3673 2047 3687
rect 1933 3653 1947 3667
rect 1993 3653 2007 3667
rect 1893 3633 1907 3647
rect 1833 3513 1847 3527
rect 1813 3473 1827 3487
rect 1853 3493 1867 3507
rect 1873 3493 1887 3507
rect 1993 3553 2007 3567
rect 1913 3533 1927 3547
rect 1953 3533 1967 3547
rect 1913 3493 1927 3507
rect 2013 3513 2027 3527
rect 2013 3493 2027 3507
rect 1813 3273 1827 3287
rect 1793 3233 1807 3247
rect 1793 3193 1807 3207
rect 1793 3173 1807 3187
rect 1753 3153 1767 3167
rect 1733 3073 1747 3087
rect 1713 3013 1727 3027
rect 1693 2993 1707 3007
rect 1693 2973 1707 2987
rect 1733 2993 1747 3007
rect 1653 2953 1667 2967
rect 1613 2873 1627 2887
rect 1633 2733 1647 2747
rect 1673 2713 1687 2727
rect 1653 2693 1667 2707
rect 1593 2653 1607 2667
rect 1573 2633 1587 2647
rect 1573 2613 1587 2627
rect 1533 2533 1547 2547
rect 1513 2513 1527 2527
rect 1553 2513 1567 2527
rect 1473 2493 1487 2507
rect 1533 2493 1547 2507
rect 1493 2453 1507 2467
rect 1453 2373 1467 2387
rect 1253 2293 1267 2307
rect 1273 2273 1287 2287
rect 1333 2293 1347 2307
rect 1413 2293 1427 2307
rect 1433 2293 1447 2307
rect 1473 2293 1487 2307
rect 1453 2273 1467 2287
rect 1293 2233 1307 2247
rect 1293 2213 1307 2227
rect 1273 2093 1287 2107
rect 1213 2073 1227 2087
rect 1193 2053 1207 2067
rect 1233 2053 1247 2067
rect 1253 2073 1267 2087
rect 1273 2053 1287 2067
rect 1233 1833 1247 1847
rect 1173 1793 1187 1807
rect 1233 1793 1247 1807
rect 1273 1793 1287 1807
rect 1253 1773 1267 1787
rect 1193 1753 1207 1767
rect 1153 1593 1167 1607
rect 1173 1573 1187 1587
rect 1193 1553 1207 1567
rect 1133 1313 1147 1327
rect 1173 1313 1187 1327
rect 1193 1333 1207 1347
rect 1353 2113 1367 2127
rect 1433 2233 1447 2247
rect 1413 2213 1427 2227
rect 1393 2093 1407 2107
rect 1373 2053 1387 2067
rect 1393 2073 1407 2087
rect 1393 1933 1407 1947
rect 1333 1793 1347 1807
rect 1393 1773 1407 1787
rect 1353 1733 1367 1747
rect 1313 1713 1327 1727
rect 1313 1673 1327 1687
rect 1293 1633 1307 1647
rect 1293 1613 1307 1627
rect 1333 1613 1347 1627
rect 1253 1553 1267 1567
rect 1313 1553 1327 1567
rect 1253 1513 1267 1527
rect 1213 1313 1227 1327
rect 1153 1293 1167 1307
rect 1293 1293 1307 1307
rect 1253 1273 1267 1287
rect 1313 1273 1327 1287
rect 1133 1153 1147 1167
rect 893 1133 907 1147
rect 933 1133 947 1147
rect 993 1133 1007 1147
rect 833 1113 847 1127
rect 773 1093 787 1107
rect 673 1073 687 1087
rect 693 1073 707 1087
rect 633 1013 647 1027
rect 673 1013 687 1027
rect 573 893 587 907
rect 613 893 627 907
rect 553 853 567 867
rect 493 813 507 827
rect 513 833 527 847
rect 553 833 567 847
rect 733 893 747 907
rect 673 853 687 867
rect 713 853 727 867
rect 793 853 807 867
rect 613 813 627 827
rect 533 793 547 807
rect 653 773 667 787
rect 673 753 687 767
rect 653 653 667 667
rect 533 633 547 647
rect 513 613 527 627
rect 813 813 827 827
rect 733 773 747 787
rect 773 753 787 767
rect 593 613 607 627
rect 673 613 687 627
rect 513 533 527 547
rect 553 413 567 427
rect 533 353 547 367
rect 473 233 487 247
rect 513 213 527 227
rect 633 593 647 607
rect 793 613 807 627
rect 873 1093 887 1107
rect 1053 1113 1067 1127
rect 1033 1093 1047 1107
rect 1113 1093 1127 1107
rect 893 1073 907 1087
rect 873 873 887 887
rect 853 833 867 847
rect 853 593 867 607
rect 673 573 687 587
rect 773 573 787 587
rect 733 393 747 407
rect 813 393 827 407
rect 653 333 667 347
rect 793 373 807 387
rect 813 273 827 287
rect 593 253 607 267
rect 573 233 587 247
rect 553 193 567 207
rect 673 193 687 207
rect 533 173 547 187
rect 573 173 587 187
rect 633 173 647 187
rect 473 133 487 147
rect 553 133 567 147
rect 653 133 667 147
rect 1193 1133 1207 1147
rect 1273 1133 1287 1147
rect 1213 1113 1227 1127
rect 1333 1133 1347 1147
rect 1293 1093 1307 1107
rect 1253 1073 1267 1087
rect 1253 1053 1267 1067
rect 1213 873 1227 887
rect 913 833 927 847
rect 893 813 907 827
rect 953 833 967 847
rect 1013 833 1027 847
rect 1013 813 1027 827
rect 933 793 947 807
rect 953 773 967 787
rect 933 673 947 687
rect 973 653 987 667
rect 993 653 1007 667
rect 973 613 987 627
rect 1073 833 1087 847
rect 1133 853 1147 867
rect 1133 833 1147 847
rect 1093 793 1107 807
rect 1033 753 1047 767
rect 1193 833 1207 847
rect 1213 813 1227 827
rect 1233 793 1247 807
rect 1113 673 1127 687
rect 1093 633 1107 647
rect 1013 613 1027 627
rect 953 373 967 387
rect 1073 593 1087 607
rect 1213 673 1227 687
rect 1153 633 1167 647
rect 1133 613 1147 627
rect 1293 1033 1307 1047
rect 1513 2273 1527 2287
rect 1493 2253 1507 2267
rect 1613 2533 1627 2547
rect 1653 2633 1667 2647
rect 1653 2593 1667 2607
rect 1693 2593 1707 2607
rect 1833 3133 1847 3147
rect 1773 3013 1787 3027
rect 1813 3013 1827 3027
rect 1833 3033 1847 3047
rect 1813 2753 1827 2767
rect 1773 2733 1787 2747
rect 1833 2713 1847 2727
rect 1753 2693 1767 2707
rect 1793 2693 1807 2707
rect 1773 2653 1787 2667
rect 1633 2513 1647 2527
rect 1573 2493 1587 2507
rect 1553 2473 1567 2487
rect 1633 2353 1647 2367
rect 1593 2313 1607 2327
rect 1553 2273 1567 2287
rect 1513 2213 1527 2227
rect 1473 2133 1487 2147
rect 1513 2093 1527 2107
rect 1473 2073 1487 2087
rect 1493 2053 1507 2067
rect 1533 2053 1547 2067
rect 1473 1973 1487 1987
rect 1573 2233 1587 2247
rect 1613 2213 1627 2227
rect 1593 2133 1607 2147
rect 1573 2113 1587 2127
rect 1573 1933 1587 1947
rect 1653 2333 1667 2347
rect 1693 2553 1707 2567
rect 1753 2533 1767 2547
rect 1713 2493 1727 2507
rect 1693 2453 1707 2467
rect 1733 2473 1747 2487
rect 1733 2453 1747 2467
rect 1713 2333 1727 2347
rect 1713 2293 1727 2307
rect 1753 2353 1767 2367
rect 1693 2253 1707 2267
rect 1713 2273 1727 2287
rect 1733 2273 1747 2287
rect 1733 2233 1747 2247
rect 1753 2233 1767 2247
rect 1753 2213 1767 2227
rect 1713 2193 1727 2207
rect 1693 2093 1707 2107
rect 1653 2073 1667 2087
rect 1673 2073 1687 2087
rect 1633 2053 1647 2067
rect 1673 2053 1687 2067
rect 1653 2033 1667 2047
rect 1693 2033 1707 2047
rect 1613 2013 1627 2027
rect 1673 2013 1687 2027
rect 1493 1773 1507 1787
rect 1533 1773 1547 1787
rect 1553 1773 1567 1787
rect 1633 1793 1647 1807
rect 1613 1773 1627 1787
rect 1433 1753 1447 1767
rect 1413 1733 1427 1747
rect 1373 1713 1387 1727
rect 1433 1673 1447 1687
rect 1373 1593 1387 1607
rect 1393 1493 1407 1507
rect 1373 1413 1387 1427
rect 1513 1753 1527 1767
rect 1493 1733 1507 1747
rect 1453 1613 1467 1627
rect 1473 1553 1487 1567
rect 1453 1333 1467 1347
rect 1433 1153 1447 1167
rect 1373 1133 1387 1147
rect 1373 1093 1387 1107
rect 1413 1073 1427 1087
rect 1453 1073 1467 1087
rect 1353 1033 1367 1047
rect 1333 873 1347 887
rect 1433 873 1447 887
rect 1293 813 1307 827
rect 1193 613 1207 627
rect 1233 613 1247 627
rect 1193 593 1207 607
rect 1373 853 1387 867
rect 1353 833 1367 847
rect 1413 853 1427 867
rect 1333 733 1347 747
rect 1313 573 1327 587
rect 1233 553 1247 567
rect 1113 533 1127 547
rect 1153 533 1167 547
rect 1013 413 1027 427
rect 833 213 847 227
rect 933 333 947 347
rect 973 353 987 367
rect 993 353 1007 367
rect 973 293 987 307
rect 1033 373 1047 387
rect 1073 373 1087 387
rect 1093 353 1107 367
rect 1053 293 1067 307
rect 1393 653 1407 667
rect 1353 633 1367 647
rect 1413 613 1427 627
rect 1413 573 1427 587
rect 1373 553 1387 567
rect 1353 373 1367 387
rect 1393 373 1407 387
rect 1373 353 1387 367
rect 1253 333 1267 347
rect 1333 333 1347 347
rect 913 213 927 227
rect 1013 213 1027 227
rect 853 193 867 207
rect 873 173 887 187
rect 893 173 907 187
rect 693 133 707 147
rect 153 113 167 127
rect 173 113 187 127
rect 233 113 247 127
rect 833 133 847 147
rect 873 133 887 147
rect 833 113 847 127
rect 1073 273 1087 287
rect 1193 273 1207 287
rect 953 153 967 167
rect 1133 193 1147 207
rect 1173 173 1187 187
rect 1233 173 1247 187
rect 1193 133 1207 147
rect 1593 1673 1607 1687
rect 1573 1613 1587 1627
rect 1633 1613 1647 1627
rect 1813 2553 1827 2567
rect 1793 2533 1807 2547
rect 1793 2493 1807 2507
rect 1973 3473 1987 3487
rect 1933 3453 1947 3467
rect 1993 3373 2007 3387
rect 1933 3293 1947 3307
rect 1913 3253 1927 3267
rect 1893 3193 1907 3207
rect 1933 3193 1947 3207
rect 1893 3153 1907 3167
rect 1933 3073 1947 3087
rect 1973 3053 1987 3067
rect 1873 3013 1887 3027
rect 1913 3013 1927 3027
rect 1973 2973 1987 2987
rect 1973 2933 1987 2947
rect 1913 2853 1927 2867
rect 1933 2793 1947 2807
rect 2053 3513 2067 3527
rect 2033 3433 2047 3447
rect 2013 3273 2027 3287
rect 2093 3713 2107 3727
rect 2153 4193 2167 4207
rect 2193 4193 2207 4207
rect 2133 4153 2147 4167
rect 2153 4033 2167 4047
rect 2173 4013 2187 4027
rect 2133 3953 2147 3967
rect 2153 3973 2167 3987
rect 2193 3973 2207 3987
rect 2133 3753 2147 3767
rect 2173 3733 2187 3747
rect 2093 3693 2107 3707
rect 2113 3693 2127 3707
rect 2233 4233 2247 4247
rect 2353 4453 2367 4467
rect 2493 4913 2507 4927
rect 2513 4933 2527 4947
rect 2613 5393 2627 5407
rect 2633 5413 2647 5427
rect 2653 5393 2667 5407
rect 2733 5593 2747 5607
rect 2773 5553 2787 5567
rect 2773 5533 2787 5547
rect 2753 5393 2767 5407
rect 2873 5653 2887 5667
rect 3253 5653 3267 5667
rect 3433 5653 3447 5667
rect 3493 5653 3507 5667
rect 2973 5633 2987 5647
rect 3073 5633 3087 5647
rect 2813 5553 2827 5567
rect 3113 5633 3127 5647
rect 3233 5613 3247 5627
rect 3293 5613 3307 5627
rect 3373 5613 3387 5627
rect 3533 5653 3547 5667
rect 3513 5633 3527 5647
rect 4093 5653 4107 5667
rect 3653 5633 3667 5647
rect 2873 5533 2887 5547
rect 2993 5533 3007 5547
rect 2853 5453 2867 5467
rect 2933 5473 2947 5487
rect 2913 5453 2927 5467
rect 2853 5413 2867 5427
rect 2893 5413 2907 5427
rect 3013 5453 3027 5467
rect 3133 5593 3147 5607
rect 3393 5593 3407 5607
rect 3393 5513 3407 5527
rect 3253 5453 3267 5467
rect 3093 5433 3107 5447
rect 3493 5613 3507 5627
rect 3533 5473 3547 5487
rect 3273 5433 3287 5447
rect 3373 5433 3387 5447
rect 3433 5433 3447 5447
rect 3033 5393 3047 5407
rect 3113 5393 3127 5407
rect 3133 5413 3147 5427
rect 3173 5413 3187 5427
rect 3153 5373 3167 5387
rect 2553 5133 2567 5147
rect 2813 5173 2827 5187
rect 2553 5113 2567 5127
rect 2613 5113 2627 5127
rect 2673 5113 2687 5127
rect 2653 5053 2667 5067
rect 2733 5153 2747 5167
rect 2713 5113 2727 5127
rect 2693 5013 2707 5027
rect 2753 4973 2767 4987
rect 2773 4973 2787 4987
rect 2533 4913 2547 4927
rect 2633 4933 2647 4947
rect 2593 4913 2607 4927
rect 2753 4913 2767 4927
rect 2533 4873 2547 4887
rect 2533 4713 2547 4727
rect 2493 4693 2507 4707
rect 2513 4673 2527 4687
rect 2513 4593 2527 4607
rect 2453 4573 2467 4587
rect 2493 4513 2507 4527
rect 2473 4493 2487 4507
rect 2413 4453 2427 4467
rect 2433 4453 2447 4467
rect 2333 4413 2347 4427
rect 2333 4393 2347 4407
rect 2333 4353 2347 4367
rect 2233 4173 2247 4187
rect 2273 4173 2287 4187
rect 2293 4153 2307 4167
rect 2373 4333 2387 4347
rect 2353 4253 2367 4267
rect 2353 4173 2367 4187
rect 2333 4153 2347 4167
rect 2253 4093 2267 4107
rect 2313 4093 2327 4107
rect 2273 4013 2287 4027
rect 2233 3973 2247 3987
rect 2413 4313 2427 4327
rect 2473 4453 2487 4467
rect 2513 4453 2527 4467
rect 2593 4853 2607 4867
rect 2573 4693 2587 4707
rect 2573 4653 2587 4667
rect 2653 4733 2667 4747
rect 2633 4653 2647 4667
rect 2593 4553 2607 4567
rect 2573 4513 2587 4527
rect 2613 4493 2627 4507
rect 2453 4333 2467 4347
rect 2433 4293 2447 4307
rect 2453 4253 2467 4267
rect 2513 4253 2527 4267
rect 2393 4213 2407 4227
rect 2493 4233 2507 4247
rect 2433 4173 2447 4187
rect 2473 4153 2487 4167
rect 2413 4133 2427 4147
rect 2393 4113 2407 4127
rect 2293 3993 2307 4007
rect 2333 3993 2347 4007
rect 2373 3993 2387 4007
rect 2313 3953 2327 3967
rect 2413 4093 2427 4107
rect 2513 4113 2527 4127
rect 2493 4013 2507 4027
rect 2433 3993 2447 4007
rect 2413 3973 2427 3987
rect 2473 3993 2487 4007
rect 2493 3973 2507 3987
rect 2493 3953 2507 3967
rect 2513 3953 2527 3967
rect 2453 3913 2467 3927
rect 2393 3873 2407 3887
rect 2453 3873 2467 3887
rect 2473 3873 2487 3887
rect 2373 3813 2387 3827
rect 2333 3753 2347 3767
rect 2273 3713 2287 3727
rect 2313 3733 2327 3747
rect 2253 3653 2267 3667
rect 2213 3613 2227 3627
rect 2253 3573 2267 3587
rect 2173 3533 2187 3547
rect 2293 3693 2307 3707
rect 2273 3553 2287 3567
rect 2093 3493 2107 3507
rect 2133 3493 2147 3507
rect 2153 3513 2167 3527
rect 2173 3493 2187 3507
rect 2113 3393 2127 3407
rect 2073 3293 2087 3307
rect 2093 3233 2107 3247
rect 2033 3133 2047 3147
rect 2033 3073 2047 3087
rect 2013 3033 2027 3047
rect 2073 3053 2087 3067
rect 2253 3493 2267 3507
rect 2293 3513 2307 3527
rect 2213 3473 2227 3487
rect 2333 3533 2347 3547
rect 2353 3513 2367 3527
rect 2333 3493 2347 3507
rect 2193 3273 2207 3287
rect 2133 3253 2147 3267
rect 2173 3233 2187 3247
rect 2193 3253 2207 3267
rect 2193 3213 2207 3227
rect 2173 3113 2187 3127
rect 2133 3093 2147 3107
rect 2113 3073 2127 3087
rect 2113 3013 2127 3027
rect 2153 2993 2167 3007
rect 2133 2893 2147 2907
rect 2033 2853 2047 2867
rect 2053 2813 2067 2827
rect 2113 2813 2127 2827
rect 1993 2793 2007 2807
rect 1953 2753 1967 2767
rect 2013 2773 2027 2787
rect 1953 2733 1967 2747
rect 1993 2733 2007 2747
rect 1913 2653 1927 2667
rect 1913 2613 1927 2627
rect 1853 2593 1867 2607
rect 1933 2593 1947 2607
rect 1873 2553 1887 2567
rect 1793 2473 1807 2487
rect 1833 2473 1847 2487
rect 1893 2473 1907 2487
rect 1873 2453 1887 2467
rect 1793 2253 1807 2267
rect 1873 2433 1887 2447
rect 1833 2333 1847 2347
rect 1873 2293 1887 2307
rect 1913 2293 1927 2307
rect 1853 2273 1867 2287
rect 1873 2273 1887 2287
rect 1813 2213 1827 2227
rect 1813 2193 1827 2207
rect 1773 2113 1787 2127
rect 1773 2093 1787 2107
rect 1833 2173 1847 2187
rect 1753 2033 1767 2047
rect 1713 1973 1727 1987
rect 1753 1933 1767 1947
rect 1693 1853 1707 1867
rect 1733 1773 1747 1787
rect 1753 1793 1767 1807
rect 1773 1753 1787 1767
rect 1893 2253 1907 2267
rect 1913 2253 1927 2267
rect 1893 2173 1907 2187
rect 1873 2153 1887 2167
rect 1853 2113 1867 2127
rect 1933 2113 1947 2127
rect 1833 2013 1847 2027
rect 1833 1953 1847 1967
rect 1893 2093 1907 2107
rect 1873 2053 1887 2067
rect 1913 2053 1927 2067
rect 1933 2073 1947 2087
rect 1913 1913 1927 1927
rect 1853 1853 1867 1867
rect 1853 1813 1867 1827
rect 1933 1873 1947 1887
rect 1833 1753 1847 1767
rect 1813 1733 1827 1747
rect 1873 1713 1887 1727
rect 1853 1693 1867 1707
rect 1793 1673 1807 1687
rect 1733 1613 1747 1627
rect 1593 1593 1607 1607
rect 1633 1593 1647 1607
rect 1553 1573 1567 1587
rect 1653 1573 1667 1587
rect 1693 1373 1707 1387
rect 1773 1553 1787 1567
rect 1833 1613 1847 1627
rect 1753 1373 1767 1387
rect 1733 1353 1747 1367
rect 1553 1313 1567 1327
rect 1553 1173 1567 1187
rect 1513 1153 1527 1167
rect 1533 1133 1547 1147
rect 1533 1093 1547 1107
rect 1493 1053 1507 1067
rect 1453 853 1467 867
rect 1473 853 1487 867
rect 1453 793 1467 807
rect 1453 693 1467 707
rect 1673 1333 1687 1347
rect 1713 1333 1727 1347
rect 1693 1313 1707 1327
rect 1613 1173 1627 1187
rect 1553 853 1567 867
rect 1573 833 1587 847
rect 1633 1153 1647 1167
rect 1793 1373 1807 1387
rect 1973 2573 1987 2587
rect 2053 2573 2067 2587
rect 2013 2553 2027 2567
rect 2033 2533 2047 2547
rect 1993 2513 2007 2527
rect 1973 2373 1987 2387
rect 2053 2313 2067 2327
rect 2013 2293 2027 2307
rect 2033 2253 2047 2267
rect 1993 2193 2007 2207
rect 1973 2113 1987 2127
rect 2093 2653 2107 2667
rect 2273 3433 2287 3447
rect 2253 3273 2267 3287
rect 2233 3253 2247 3267
rect 2233 3213 2247 3227
rect 2213 3193 2227 3207
rect 2313 3293 2327 3307
rect 2293 3213 2307 3227
rect 2253 3113 2267 3127
rect 2233 3033 2247 3047
rect 2253 3013 2267 3027
rect 2273 3033 2287 3047
rect 2193 2953 2207 2967
rect 2233 2913 2247 2927
rect 2193 2893 2207 2907
rect 2173 2813 2187 2827
rect 2173 2793 2187 2807
rect 2153 2733 2167 2747
rect 2133 2553 2147 2567
rect 2093 2533 2107 2547
rect 2113 2533 2127 2547
rect 2113 2513 2127 2527
rect 2153 2533 2167 2547
rect 2193 2773 2207 2787
rect 2213 2773 2227 2787
rect 2193 2733 2207 2747
rect 2213 2733 2227 2747
rect 2193 2593 2207 2607
rect 2173 2513 2187 2527
rect 2093 2413 2107 2427
rect 2153 2493 2167 2507
rect 2133 2353 2147 2367
rect 2113 2333 2127 2347
rect 2253 2693 2267 2707
rect 2233 2553 2247 2567
rect 2313 3153 2327 3167
rect 2393 3793 2407 3807
rect 2473 3793 2487 3807
rect 2413 3713 2427 3727
rect 2453 3713 2467 3727
rect 2473 3693 2487 3707
rect 2433 3633 2447 3647
rect 2393 3573 2407 3587
rect 2433 3573 2447 3587
rect 2393 3533 2407 3547
rect 2373 3493 2387 3507
rect 2453 3493 2467 3507
rect 2353 3453 2367 3467
rect 2413 3293 2427 3307
rect 2473 3253 2487 3267
rect 2393 3213 2407 3227
rect 2373 3193 2387 3207
rect 2333 3133 2347 3147
rect 2353 3113 2367 3127
rect 2353 3053 2367 3067
rect 2433 3113 2447 3127
rect 2413 3053 2427 3067
rect 2353 3013 2367 3027
rect 2393 3013 2407 3027
rect 2413 3013 2427 3027
rect 2313 2793 2327 2807
rect 2293 2713 2307 2727
rect 2353 2753 2367 2767
rect 2373 2773 2387 2787
rect 2433 2913 2447 2927
rect 2433 2793 2447 2807
rect 2413 2753 2427 2767
rect 2313 2693 2327 2707
rect 2313 2593 2327 2607
rect 2413 2593 2427 2607
rect 2273 2573 2287 2587
rect 2353 2573 2367 2587
rect 2333 2533 2347 2547
rect 2293 2513 2307 2527
rect 2373 2553 2387 2567
rect 2353 2513 2367 2527
rect 2253 2473 2267 2487
rect 2333 2473 2347 2487
rect 2213 2453 2227 2467
rect 2233 2453 2247 2467
rect 2173 2373 2187 2387
rect 2073 2273 2087 2287
rect 2153 2313 2167 2327
rect 2133 2293 2147 2307
rect 2113 2253 2127 2267
rect 2093 2213 2107 2227
rect 1993 2073 2007 2087
rect 2093 2073 2107 2087
rect 2053 2053 2067 2067
rect 2073 2053 2087 2067
rect 2113 2053 2127 2067
rect 2073 2033 2087 2047
rect 2013 1973 2027 1987
rect 1973 1933 1987 1947
rect 1973 1873 1987 1887
rect 2053 1933 2067 1947
rect 1953 1813 1967 1827
rect 1933 1733 1947 1747
rect 1913 1673 1927 1687
rect 1993 1673 2007 1687
rect 2033 1613 2047 1627
rect 2033 1573 2047 1587
rect 2033 1473 2047 1487
rect 1873 1333 1887 1347
rect 1933 1333 1947 1347
rect 1793 1233 1807 1247
rect 1753 1073 1767 1087
rect 1833 1133 1847 1147
rect 1813 993 1827 1007
rect 1633 853 1647 867
rect 1713 853 1727 867
rect 1613 793 1627 807
rect 1533 673 1547 687
rect 1513 653 1527 667
rect 1513 633 1527 647
rect 1533 613 1547 627
rect 1593 613 1607 627
rect 1553 593 1567 607
rect 1473 553 1487 567
rect 1473 393 1487 407
rect 1453 353 1467 367
rect 1733 813 1747 827
rect 1773 833 1787 847
rect 1973 1333 1987 1347
rect 1953 1313 1967 1327
rect 2013 1333 2027 1347
rect 1993 1273 2007 1287
rect 2113 1833 2127 1847
rect 2193 2313 2207 2327
rect 2173 2233 2187 2247
rect 2153 2153 2167 2167
rect 2333 2233 2347 2247
rect 2333 2213 2347 2227
rect 2273 2173 2287 2187
rect 2233 2153 2247 2167
rect 2193 2073 2207 2087
rect 2213 1833 2227 1847
rect 2153 1813 2167 1827
rect 2193 1813 2207 1827
rect 2173 1773 2187 1787
rect 2133 1593 2147 1607
rect 2113 1473 2127 1487
rect 2073 1373 2087 1387
rect 2053 1313 2067 1327
rect 2093 1273 2107 1287
rect 2093 1253 2107 1267
rect 2013 1173 2027 1187
rect 2073 1173 2087 1187
rect 2033 1113 2047 1127
rect 1873 1073 1887 1087
rect 1913 1093 1927 1107
rect 2013 1093 2027 1107
rect 2053 1093 2067 1107
rect 1933 1073 1947 1087
rect 1953 1073 1967 1087
rect 1853 1053 1867 1067
rect 1893 1053 1907 1067
rect 1853 873 1867 887
rect 1833 833 1847 847
rect 1893 853 1907 867
rect 1913 833 1927 847
rect 1813 813 1827 827
rect 1873 813 1887 827
rect 1773 793 1787 807
rect 1753 773 1767 787
rect 1653 653 1667 667
rect 1673 633 1687 647
rect 1653 613 1667 627
rect 1693 613 1707 627
rect 1713 633 1727 647
rect 1733 633 1747 647
rect 1633 413 1647 427
rect 1713 593 1727 607
rect 1513 373 1527 387
rect 1593 373 1607 387
rect 1653 373 1667 387
rect 1693 373 1707 387
rect 1613 353 1627 367
rect 1713 353 1727 367
rect 2073 1053 2087 1067
rect 1973 833 1987 847
rect 2033 853 2047 867
rect 2053 853 2067 867
rect 2013 813 2027 827
rect 1993 773 2007 787
rect 1973 753 1987 767
rect 1953 733 1967 747
rect 1813 693 1827 707
rect 1853 693 1867 707
rect 1813 673 1827 687
rect 1933 653 1947 667
rect 1993 733 2007 747
rect 1993 653 2007 667
rect 1773 613 1787 627
rect 1853 613 1867 627
rect 1913 613 1927 627
rect 1953 613 1967 627
rect 1993 633 2007 647
rect 1993 613 2007 627
rect 1833 593 1847 607
rect 1793 573 1807 587
rect 1833 553 1847 567
rect 1773 373 1787 387
rect 1673 333 1687 347
rect 1733 333 1747 347
rect 1813 333 1827 347
rect 1533 313 1547 327
rect 1613 313 1627 327
rect 1633 293 1647 307
rect 1313 173 1327 187
rect 1333 173 1347 187
rect 1273 153 1287 167
rect 1293 153 1307 167
rect 1593 193 1607 207
rect 1433 173 1447 187
rect 1733 173 1747 187
rect 1233 133 1247 147
rect 1413 153 1427 167
rect 893 113 907 127
rect 933 113 947 127
rect 953 113 967 127
rect 1033 113 1047 127
rect 1693 153 1707 167
rect 1573 133 1587 147
rect 1673 133 1687 147
rect 1713 133 1727 147
rect 1793 153 1807 167
rect 1753 133 1767 147
rect 1493 113 1507 127
rect 2073 813 2087 827
rect 2133 1373 2147 1387
rect 2113 1093 2127 1107
rect 2473 3053 2487 3067
rect 2473 2993 2487 3007
rect 2593 4433 2607 4447
rect 2693 4693 2707 4707
rect 2673 4613 2687 4627
rect 2673 4593 2687 4607
rect 2673 4573 2687 4587
rect 2653 4393 2667 4407
rect 2633 4373 2647 4387
rect 2593 4193 2607 4207
rect 2593 4173 2607 4187
rect 2553 4133 2567 4147
rect 2633 4193 2647 4207
rect 2753 4693 2767 4707
rect 2793 4693 2807 4707
rect 2833 5033 2847 5047
rect 2873 5133 2887 5147
rect 2893 5153 2907 5167
rect 2993 5133 3007 5147
rect 3033 5133 3047 5147
rect 3113 5133 3127 5147
rect 2913 5113 2927 5127
rect 3033 5093 3047 5107
rect 2993 5013 3007 5027
rect 2853 4973 2867 4987
rect 2973 4953 2987 4967
rect 2873 4933 2887 4947
rect 2953 4933 2967 4947
rect 2873 4913 2887 4927
rect 3133 5113 3147 5127
rect 3053 4993 3067 5007
rect 3113 4993 3127 5007
rect 3153 4993 3167 5007
rect 3293 5413 3307 5427
rect 3333 5413 3347 5427
rect 3173 4973 3187 4987
rect 3233 4973 3247 4987
rect 3133 4953 3147 4967
rect 2813 4673 2827 4687
rect 2733 4653 2747 4667
rect 2773 4653 2787 4667
rect 2773 4633 2787 4647
rect 2753 4553 2767 4567
rect 2833 4553 2847 4567
rect 2713 4493 2727 4507
rect 3173 4913 3187 4927
rect 3133 4833 3147 4847
rect 3133 4713 3147 4727
rect 2953 4693 2967 4707
rect 3033 4693 3047 4707
rect 3073 4673 3087 4687
rect 3093 4653 3107 4667
rect 2913 4613 2927 4627
rect 2893 4573 2907 4587
rect 3013 4573 3027 4587
rect 2873 4513 2887 4527
rect 2913 4513 2927 4527
rect 2853 4493 2867 4507
rect 2733 4453 2747 4467
rect 2753 4453 2767 4467
rect 2713 4433 2727 4447
rect 2733 4353 2747 4367
rect 2693 4293 2707 4307
rect 2713 4253 2727 4267
rect 2713 4213 2727 4227
rect 2713 4193 2727 4207
rect 2673 4133 2687 4147
rect 2713 4133 2727 4147
rect 2693 4113 2707 4127
rect 2633 3993 2647 4007
rect 2673 3993 2687 4007
rect 2553 3953 2567 3967
rect 2613 3973 2627 3987
rect 2593 3953 2607 3967
rect 2633 3953 2647 3967
rect 2693 3953 2707 3967
rect 2513 3873 2527 3887
rect 2533 3873 2547 3887
rect 2573 3753 2587 3767
rect 2553 3713 2567 3727
rect 2613 3913 2627 3927
rect 2613 3873 2627 3887
rect 2593 3673 2607 3687
rect 2513 3653 2527 3667
rect 2513 3633 2527 3647
rect 2593 3613 2607 3627
rect 2533 3513 2547 3527
rect 2573 3513 2587 3527
rect 2553 3473 2567 3487
rect 2553 3413 2567 3427
rect 2553 3353 2567 3367
rect 2673 3913 2687 3927
rect 2653 3873 2667 3887
rect 2653 3793 2667 3807
rect 2873 4473 2887 4487
rect 2773 4213 2787 4227
rect 2753 4113 2767 4127
rect 2893 4233 2907 4247
rect 2833 4213 2847 4227
rect 2873 4213 2887 4227
rect 3013 4493 3027 4507
rect 2993 4473 3007 4487
rect 2933 4453 2947 4467
rect 2973 4453 2987 4467
rect 2993 4433 3007 4447
rect 2933 4333 2947 4347
rect 3113 4513 3127 4527
rect 3173 4873 3187 4887
rect 3153 4693 3167 4707
rect 3133 4493 3147 4507
rect 3193 4733 3207 4747
rect 3293 5113 3307 5127
rect 3273 5013 3287 5027
rect 3413 5413 3427 5427
rect 3433 5393 3447 5407
rect 3333 5373 3347 5387
rect 3673 5593 3687 5607
rect 3613 5573 3627 5587
rect 3553 5453 3567 5467
rect 3533 5433 3547 5447
rect 3593 5433 3607 5447
rect 3573 5413 3587 5427
rect 3493 5253 3507 5267
rect 3553 5213 3567 5227
rect 3553 5173 3567 5187
rect 3373 5113 3387 5127
rect 3313 4973 3327 4987
rect 3513 5113 3527 5127
rect 3393 4993 3407 5007
rect 3413 4993 3427 5007
rect 3513 4993 3527 5007
rect 3553 5113 3567 5127
rect 3433 4973 3447 4987
rect 3493 4973 3507 4987
rect 3533 4973 3547 4987
rect 3313 4953 3327 4967
rect 3373 4953 3387 4967
rect 3373 4933 3387 4947
rect 3413 4933 3427 4947
rect 3433 4933 3447 4947
rect 3433 4893 3447 4907
rect 3293 4873 3307 4887
rect 3313 4853 3327 4867
rect 3233 4713 3247 4727
rect 3433 4793 3447 4807
rect 3393 4773 3407 4787
rect 3193 4693 3207 4707
rect 3253 4673 3267 4687
rect 3333 4673 3347 4687
rect 3173 4653 3187 4667
rect 3173 4633 3187 4647
rect 3033 4353 3047 4367
rect 2993 4333 3007 4347
rect 3033 4333 3047 4347
rect 2953 4273 2967 4287
rect 3013 4233 3027 4247
rect 2953 4213 2967 4227
rect 2913 4193 2927 4207
rect 2873 4153 2887 4167
rect 2893 4153 2907 4167
rect 2853 4133 2867 4147
rect 2833 4093 2847 4107
rect 2833 4073 2847 4087
rect 2813 4033 2827 4047
rect 2813 3993 2827 4007
rect 2753 3973 2767 3987
rect 2773 3973 2787 3987
rect 2753 3953 2767 3967
rect 2793 3953 2807 3967
rect 2753 3853 2767 3867
rect 2733 3813 2747 3827
rect 2693 3773 2707 3787
rect 2693 3733 2707 3747
rect 2673 3713 2687 3727
rect 2713 3713 2727 3727
rect 2713 3693 2727 3707
rect 2633 3653 2647 3667
rect 2693 3673 2707 3687
rect 2613 3313 2627 3327
rect 2573 3273 2587 3287
rect 2573 3213 2587 3227
rect 2593 3233 2607 3247
rect 2553 3173 2567 3187
rect 2613 3153 2627 3167
rect 2593 3133 2607 3147
rect 2513 3113 2527 3127
rect 2573 3113 2587 3127
rect 2513 3093 2527 3107
rect 2553 3053 2567 3067
rect 2573 3053 2587 3067
rect 2533 3013 2547 3027
rect 2453 2773 2467 2787
rect 2453 2733 2467 2747
rect 2433 2553 2447 2567
rect 2393 2513 2407 2527
rect 2433 2513 2447 2527
rect 2473 2693 2487 2707
rect 2493 2693 2507 2707
rect 2513 2613 2527 2627
rect 2653 3473 2667 3487
rect 2673 3493 2687 3507
rect 2733 3633 2747 3647
rect 2733 3613 2747 3627
rect 2733 3493 2747 3507
rect 2693 3473 2707 3487
rect 2713 3473 2727 3487
rect 2653 3353 2667 3367
rect 2753 3333 2767 3347
rect 2753 3313 2767 3327
rect 2673 3293 2687 3307
rect 2653 3273 2667 3287
rect 2653 3193 2667 3207
rect 2653 3173 2667 3187
rect 2633 3093 2647 3107
rect 2633 3073 2647 3087
rect 2713 3253 2727 3267
rect 2813 3793 2827 3807
rect 2793 3733 2807 3747
rect 2833 3753 2847 3767
rect 2833 3713 2847 3727
rect 2793 3673 2807 3687
rect 2833 3673 2847 3687
rect 2873 4033 2887 4047
rect 2873 4013 2887 4027
rect 2953 4113 2967 4127
rect 2873 3933 2887 3947
rect 2973 4053 2987 4067
rect 3153 4373 3167 4387
rect 3033 4173 3047 4187
rect 3113 4153 3127 4167
rect 3073 4113 3087 4127
rect 3053 4093 3067 4107
rect 2993 4013 3007 4027
rect 3033 4013 3047 4027
rect 2913 3973 2927 3987
rect 2953 3973 2967 3987
rect 2933 3953 2947 3967
rect 2993 3973 3007 3987
rect 2973 3953 2987 3967
rect 2953 3933 2967 3947
rect 3033 3953 3047 3967
rect 3093 4013 3107 4027
rect 3053 3933 3067 3947
rect 2993 3913 3007 3927
rect 2993 3893 3007 3907
rect 3013 3893 3027 3907
rect 2953 3873 2967 3887
rect 2953 3793 2967 3807
rect 2913 3713 2927 3727
rect 2933 3693 2947 3707
rect 2993 3693 3007 3707
rect 2973 3673 2987 3687
rect 2933 3653 2947 3667
rect 2893 3573 2907 3587
rect 2813 3513 2827 3527
rect 2793 3493 2807 3507
rect 2873 3513 2887 3527
rect 2873 3493 2887 3507
rect 2833 3473 2847 3487
rect 2853 3473 2867 3487
rect 2853 3373 2867 3387
rect 2793 3333 2807 3347
rect 2773 3273 2787 3287
rect 2873 3293 2887 3307
rect 2693 3213 2707 3227
rect 2753 3233 2767 3247
rect 2733 3193 2747 3207
rect 2793 3233 2807 3247
rect 2813 3233 2827 3247
rect 2833 3233 2847 3247
rect 2693 3113 2707 3127
rect 2753 3113 2767 3127
rect 2673 3073 2687 3087
rect 2653 3033 2667 3047
rect 2733 3033 2747 3047
rect 2673 2993 2687 3007
rect 2693 2993 2707 3007
rect 2593 2913 2607 2927
rect 2573 2813 2587 2827
rect 2633 2773 2647 2787
rect 2673 2773 2687 2787
rect 2653 2753 2667 2767
rect 2713 2973 2727 2987
rect 2713 2953 2727 2967
rect 2693 2733 2707 2747
rect 2653 2713 2667 2727
rect 2493 2533 2507 2547
rect 2473 2513 2487 2527
rect 2493 2513 2507 2527
rect 2433 2493 2447 2507
rect 2453 2493 2467 2507
rect 2373 2373 2387 2387
rect 2493 2473 2507 2487
rect 2573 2593 2587 2607
rect 2613 2593 2627 2607
rect 2633 2593 2647 2607
rect 2553 2573 2567 2587
rect 2593 2533 2607 2547
rect 2613 2553 2627 2567
rect 2593 2473 2607 2487
rect 2553 2413 2567 2427
rect 2513 2353 2527 2367
rect 2453 2273 2467 2287
rect 2293 2033 2307 2047
rect 2293 1993 2307 2007
rect 2253 1953 2267 1967
rect 2253 1813 2267 1827
rect 2233 1793 2247 1807
rect 2233 1693 2247 1707
rect 2273 1793 2287 1807
rect 2353 2013 2367 2027
rect 2433 2153 2447 2167
rect 2413 2093 2427 2107
rect 2373 1993 2387 2007
rect 2333 1933 2347 1947
rect 2533 2273 2547 2287
rect 2773 3073 2787 3087
rect 2773 3033 2787 3047
rect 2853 3193 2867 3207
rect 2853 3133 2867 3147
rect 2873 3073 2887 3087
rect 2853 3033 2867 3047
rect 2873 3013 2887 3027
rect 2773 2853 2787 2867
rect 2753 2793 2767 2807
rect 2753 2773 2767 2787
rect 2853 2873 2867 2887
rect 2833 2793 2847 2807
rect 2833 2753 2847 2767
rect 2833 2733 2847 2747
rect 2733 2693 2747 2707
rect 2713 2573 2727 2587
rect 2773 2573 2787 2587
rect 2673 2553 2687 2567
rect 2713 2553 2727 2567
rect 2713 2513 2727 2527
rect 2693 2473 2707 2487
rect 2653 2293 2667 2307
rect 2753 2493 2767 2507
rect 2773 2433 2787 2447
rect 2813 2693 2827 2707
rect 2993 3533 3007 3547
rect 2913 3413 2927 3427
rect 2913 3373 2927 3387
rect 2913 3293 2927 3307
rect 3133 4113 3147 4127
rect 3153 4113 3167 4127
rect 3153 4053 3167 4067
rect 3133 4033 3147 4047
rect 3113 3833 3127 3847
rect 3133 3833 3147 3847
rect 3113 3793 3127 3807
rect 3033 3733 3047 3747
rect 3073 3733 3087 3747
rect 3033 3693 3047 3707
rect 3113 3693 3127 3707
rect 3133 3673 3147 3687
rect 3073 3653 3087 3667
rect 3073 3593 3087 3607
rect 3093 3593 3107 3607
rect 3033 3533 3047 3547
rect 3053 3533 3067 3547
rect 3013 3453 3027 3467
rect 3053 3513 3067 3527
rect 3053 3493 3067 3507
rect 3053 3453 3067 3467
rect 3113 3453 3127 3467
rect 3033 3313 3047 3327
rect 2933 3253 2947 3267
rect 2913 3233 2927 3247
rect 3013 3213 3027 3227
rect 2913 3173 2927 3187
rect 2893 2953 2907 2967
rect 2893 2873 2907 2887
rect 2873 2853 2887 2867
rect 2933 3073 2947 3087
rect 2953 3053 2967 3067
rect 2973 3053 2987 3067
rect 2973 3033 2987 3047
rect 2973 2913 2987 2927
rect 2953 2833 2967 2847
rect 2913 2793 2927 2807
rect 2913 2733 2927 2747
rect 2873 2713 2887 2727
rect 2913 2713 2927 2727
rect 2833 2553 2847 2567
rect 2813 2533 2827 2547
rect 2853 2533 2867 2547
rect 2873 2533 2887 2547
rect 2933 2673 2947 2687
rect 2933 2533 2947 2547
rect 2793 2293 2807 2307
rect 2633 2253 2647 2267
rect 2773 2273 2787 2287
rect 2773 2253 2787 2267
rect 2593 2213 2607 2227
rect 2513 2173 2527 2187
rect 2553 2173 2567 2187
rect 2473 2053 2487 2067
rect 2613 2113 2627 2127
rect 2613 2053 2627 2067
rect 2413 1893 2427 1907
rect 2253 1633 2267 1647
rect 2253 1573 2267 1587
rect 2233 1373 2247 1387
rect 2193 1333 2207 1347
rect 2233 1333 2247 1347
rect 2253 1313 2267 1327
rect 2173 1113 2187 1127
rect 2153 1073 2167 1087
rect 2213 1293 2227 1307
rect 2453 1753 2467 1767
rect 2613 1953 2627 1967
rect 2593 1933 2607 1947
rect 2553 1893 2567 1907
rect 2573 1793 2587 1807
rect 2553 1753 2567 1767
rect 2573 1733 2587 1747
rect 2393 1693 2407 1707
rect 2473 1693 2487 1707
rect 2333 1613 2347 1627
rect 2293 1593 2307 1607
rect 2313 1573 2327 1587
rect 2353 1573 2367 1587
rect 2513 1673 2527 1687
rect 2493 1633 2507 1647
rect 2413 1593 2427 1607
rect 2453 1573 2467 1587
rect 2293 1433 2307 1447
rect 2293 1333 2307 1347
rect 2373 1333 2387 1347
rect 2353 1293 2367 1307
rect 2313 1273 2327 1287
rect 2333 1273 2347 1287
rect 2273 1253 2287 1267
rect 2313 1193 2327 1207
rect 2213 1133 2227 1147
rect 2253 1133 2267 1147
rect 2313 1113 2327 1127
rect 2353 1253 2367 1267
rect 2393 1313 2407 1327
rect 2373 1233 2387 1247
rect 2373 1113 2387 1127
rect 2273 1093 2287 1107
rect 2193 1073 2207 1087
rect 2233 913 2247 927
rect 2133 893 2147 907
rect 2213 893 2227 907
rect 2133 853 2147 867
rect 2153 813 2167 827
rect 2113 793 2127 807
rect 2093 753 2107 767
rect 2173 673 2187 687
rect 2093 653 2107 667
rect 2113 653 2127 667
rect 2073 633 2087 647
rect 2053 593 2067 607
rect 2173 573 2187 587
rect 2073 493 2087 507
rect 1913 393 1927 407
rect 1853 373 1867 387
rect 1993 373 2007 387
rect 1913 333 1927 347
rect 2033 353 2047 367
rect 1893 173 1907 187
rect 1913 153 1927 167
rect 1953 133 1967 147
rect 1933 113 1947 127
rect 2333 1093 2347 1107
rect 2353 1093 2367 1107
rect 2293 913 2307 927
rect 2293 893 2307 907
rect 2273 873 2287 887
rect 2253 653 2267 667
rect 2233 633 2247 647
rect 2313 793 2327 807
rect 2393 1093 2407 1107
rect 2433 1533 2447 1547
rect 2533 1613 2547 1627
rect 2613 1833 2627 1847
rect 2713 2233 2727 2247
rect 2713 2213 2727 2227
rect 2773 2193 2787 2207
rect 2753 2093 2767 2107
rect 2713 1933 2727 1947
rect 2773 1953 2787 1967
rect 2693 1893 2707 1907
rect 2833 2393 2847 2407
rect 2833 2273 2847 2287
rect 2893 2253 2907 2267
rect 2913 2233 2927 2247
rect 2853 2213 2867 2227
rect 2893 2113 2907 2127
rect 2853 2093 2867 2107
rect 2933 2213 2947 2227
rect 2913 2093 2927 2107
rect 2873 2053 2887 2067
rect 2913 2053 2927 2067
rect 2833 2013 2847 2027
rect 2793 1873 2807 1887
rect 2813 1873 2827 1887
rect 2753 1833 2767 1847
rect 2653 1793 2667 1807
rect 2633 1773 2647 1787
rect 2593 1713 2607 1727
rect 2593 1593 2607 1607
rect 2453 1273 2467 1287
rect 2533 1453 2547 1467
rect 2593 1413 2607 1427
rect 2553 1393 2567 1407
rect 2653 1513 2667 1527
rect 2613 1393 2627 1407
rect 2633 1353 2647 1367
rect 2693 1753 2707 1767
rect 2553 1293 2567 1307
rect 2613 1293 2627 1307
rect 2673 1313 2687 1327
rect 2533 1273 2547 1287
rect 2513 1213 2527 1227
rect 2493 1173 2507 1187
rect 2433 1133 2447 1147
rect 2453 1113 2467 1127
rect 2473 1093 2487 1107
rect 2413 1033 2427 1047
rect 2553 1133 2567 1147
rect 2533 1093 2547 1107
rect 2593 1113 2607 1127
rect 2633 1093 2647 1107
rect 2513 1033 2527 1047
rect 2613 1073 2627 1087
rect 2553 893 2567 907
rect 2513 853 2527 867
rect 2633 853 2647 867
rect 2573 833 2587 847
rect 2433 813 2447 827
rect 2373 693 2387 707
rect 2273 633 2287 647
rect 2433 753 2447 767
rect 2353 593 2367 607
rect 2473 613 2487 627
rect 2333 533 2347 547
rect 2293 493 2307 507
rect 2253 413 2267 427
rect 2133 353 2147 367
rect 2213 353 2227 367
rect 2173 193 2187 207
rect 2173 173 2187 187
rect 2113 153 2127 167
rect 2153 153 2167 167
rect 1973 113 1987 127
rect 2073 113 2087 127
rect 2353 393 2367 407
rect 2273 333 2287 347
rect 2293 353 2307 367
rect 2413 353 2427 367
rect 2493 553 2507 567
rect 2773 1813 2787 1827
rect 2753 1753 2767 1767
rect 2713 1733 2727 1747
rect 2713 1613 2727 1627
rect 2813 1853 2827 1867
rect 2793 1793 2807 1807
rect 2833 1813 2847 1827
rect 2873 1813 2887 1827
rect 2853 1793 2867 1807
rect 2893 1773 2907 1787
rect 2813 1753 2827 1767
rect 2913 1733 2927 1747
rect 2813 1713 2827 1727
rect 2913 1713 2927 1727
rect 2793 1613 2807 1627
rect 2713 1553 2727 1567
rect 2733 1573 2747 1587
rect 2753 1533 2767 1547
rect 2793 1533 2807 1547
rect 2733 1413 2747 1427
rect 2713 1313 2727 1327
rect 2733 1313 2747 1327
rect 2773 1293 2787 1307
rect 2713 1273 2727 1287
rect 2773 1273 2787 1287
rect 2693 1193 2707 1207
rect 2733 1213 2747 1227
rect 2753 1193 2767 1207
rect 2713 1173 2727 1187
rect 2753 1113 2767 1127
rect 2673 1093 2687 1107
rect 2733 1093 2747 1107
rect 2893 1653 2907 1667
rect 2853 1633 2867 1647
rect 2853 1513 2867 1527
rect 2833 1393 2847 1407
rect 2913 1533 2927 1547
rect 2993 2773 3007 2787
rect 2993 2713 3007 2727
rect 2973 2593 2987 2607
rect 2993 2593 3007 2607
rect 2973 2533 2987 2547
rect 3093 3393 3107 3407
rect 3073 3273 3087 3287
rect 3053 3213 3067 3227
rect 3033 3193 3047 3207
rect 3033 3113 3047 3127
rect 3253 4633 3267 4647
rect 3413 4713 3427 4727
rect 3413 4673 3427 4687
rect 3353 4613 3367 4627
rect 3293 4593 3307 4607
rect 3213 4553 3227 4567
rect 3213 4533 3227 4547
rect 3253 4533 3267 4547
rect 3213 4493 3227 4507
rect 3233 4193 3247 4207
rect 3273 4173 3287 4187
rect 3233 4153 3247 4167
rect 3213 4113 3227 4127
rect 3233 4113 3247 4127
rect 3193 4093 3207 4107
rect 3173 4013 3187 4027
rect 3213 4053 3227 4067
rect 3273 4093 3287 4107
rect 3253 3993 3267 4007
rect 3313 4493 3327 4507
rect 3353 4473 3367 4487
rect 3373 4473 3387 4487
rect 3333 4433 3347 4447
rect 3333 4393 3347 4407
rect 3313 4273 3327 4287
rect 3353 4173 3367 4187
rect 3373 4193 3387 4207
rect 3413 4193 3427 4207
rect 3333 4153 3347 4167
rect 3373 4153 3387 4167
rect 3313 4073 3327 4087
rect 3333 4073 3347 4087
rect 3293 4033 3307 4047
rect 3333 4053 3347 4067
rect 3353 4033 3367 4047
rect 3313 4013 3327 4027
rect 3273 3973 3287 3987
rect 3253 3953 3267 3967
rect 3233 3873 3247 3887
rect 3233 3833 3247 3847
rect 3253 3833 3267 3847
rect 3213 3713 3227 3727
rect 3233 3733 3247 3747
rect 3313 3973 3327 3987
rect 3293 3813 3307 3827
rect 3333 3813 3347 3827
rect 3293 3753 3307 3767
rect 3313 3733 3327 3747
rect 3453 4753 3467 4767
rect 3473 4753 3487 4767
rect 3473 4693 3487 4707
rect 3513 4913 3527 4927
rect 3573 4913 3587 4927
rect 3853 5633 3867 5647
rect 3953 5633 3967 5647
rect 3933 5593 3947 5607
rect 3773 5573 3787 5587
rect 3713 5533 3727 5547
rect 3733 5533 3747 5547
rect 3793 5513 3807 5527
rect 3753 5493 3767 5507
rect 3773 5493 3787 5507
rect 3733 5433 3747 5447
rect 3673 5393 3687 5407
rect 3693 5413 3707 5427
rect 3713 5413 3727 5427
rect 3733 5413 3747 5427
rect 3713 5393 3727 5407
rect 3633 5193 3647 5207
rect 3693 5173 3707 5187
rect 3653 5133 3667 5147
rect 3713 5093 3727 5107
rect 3573 4893 3587 4907
rect 3613 4893 3627 4907
rect 3553 4853 3567 4867
rect 3493 4673 3507 4687
rect 3533 4653 3547 4667
rect 3453 4633 3467 4647
rect 3493 4633 3507 4647
rect 3453 4513 3467 4527
rect 3473 4513 3487 4527
rect 3513 4493 3527 4507
rect 3533 4473 3547 4487
rect 3553 4453 3567 4467
rect 3513 4393 3527 4407
rect 3453 4193 3467 4207
rect 3493 4193 3507 4207
rect 3533 4193 3547 4207
rect 3473 4153 3487 4167
rect 3393 4093 3407 4107
rect 3433 4093 3447 4107
rect 3393 4073 3407 4087
rect 3373 3833 3387 3847
rect 3353 3793 3367 3807
rect 3713 4873 3727 4887
rect 3673 4853 3687 4867
rect 3653 4733 3667 4747
rect 3593 4713 3607 4727
rect 3633 4673 3647 4687
rect 3653 4673 3667 4687
rect 3613 4653 3627 4667
rect 3633 4633 3647 4647
rect 3653 4593 3667 4607
rect 3653 4513 3667 4527
rect 3593 4473 3607 4487
rect 3633 4473 3647 4487
rect 3593 4433 3607 4447
rect 3653 4433 3667 4447
rect 3633 4413 3647 4427
rect 3613 4393 3627 4407
rect 3633 4373 3647 4387
rect 3593 4253 3607 4267
rect 3573 4233 3587 4247
rect 3513 4153 3527 4167
rect 3553 4153 3567 4167
rect 3493 4113 3507 4127
rect 3493 4093 3507 4107
rect 3433 3993 3447 4007
rect 3413 3973 3427 3987
rect 3553 4053 3567 4067
rect 3693 4813 3707 4827
rect 3993 5593 4007 5607
rect 4073 5593 4087 5607
rect 3973 5553 3987 5567
rect 3973 5533 3987 5547
rect 3953 5513 3967 5527
rect 3853 5493 3867 5507
rect 3953 5493 3967 5507
rect 3973 5493 3987 5507
rect 3913 5473 3927 5487
rect 3833 5453 3847 5467
rect 3813 5433 3827 5447
rect 3793 5413 3807 5427
rect 3893 5433 3907 5447
rect 3833 5413 3847 5427
rect 3853 5413 3867 5427
rect 3773 5373 3787 5387
rect 3773 5173 3787 5187
rect 3793 5153 3807 5167
rect 3833 5033 3847 5047
rect 3773 4993 3787 5007
rect 3833 4993 3847 5007
rect 3873 5393 3887 5407
rect 3893 5393 3907 5407
rect 4133 5573 4147 5587
rect 4273 5613 4287 5627
rect 4233 5593 4247 5607
rect 5073 5773 5087 5787
rect 4833 5673 4847 5687
rect 4973 5673 4987 5687
rect 4713 5653 4727 5667
rect 4733 5653 4747 5667
rect 4873 5653 4887 5667
rect 4893 5653 4907 5667
rect 4453 5633 4467 5647
rect 4473 5613 4487 5627
rect 4493 5633 4507 5647
rect 4553 5633 4567 5647
rect 4513 5553 4527 5567
rect 4533 5513 4547 5527
rect 4433 5473 4447 5487
rect 4313 5453 4327 5467
rect 4373 5453 4387 5467
rect 4093 5433 4107 5447
rect 3993 5373 4007 5387
rect 4113 5413 4127 5427
rect 4153 5433 4167 5447
rect 4153 5393 4167 5407
rect 4233 5413 4247 5427
rect 4253 5393 4267 5407
rect 4353 5413 4367 5427
rect 4373 5393 4387 5407
rect 4413 5393 4427 5407
rect 4133 5373 4147 5387
rect 4053 5353 4067 5367
rect 4073 5353 4087 5367
rect 3973 5253 3987 5267
rect 3973 5193 3987 5207
rect 3913 5173 3927 5187
rect 3893 5153 3907 5167
rect 3913 5093 3927 5107
rect 3853 4973 3867 4987
rect 3813 4933 3827 4947
rect 3833 4913 3847 4927
rect 3933 5053 3947 5067
rect 3953 4973 3967 4987
rect 3873 4813 3887 4827
rect 3793 4793 3807 4807
rect 3913 4773 3927 4787
rect 3813 4713 3827 4727
rect 3753 4693 3767 4707
rect 3753 4673 3767 4687
rect 3833 4693 3847 4707
rect 3733 4633 3747 4647
rect 3813 4633 3827 4647
rect 3713 4593 3727 4607
rect 3693 4473 3707 4487
rect 3693 4433 3707 4447
rect 3673 4213 3687 4227
rect 3593 4173 3607 4187
rect 3633 4173 3647 4187
rect 3573 4033 3587 4047
rect 3453 3933 3467 3947
rect 3373 3753 3387 3767
rect 3353 3733 3367 3747
rect 3333 3713 3347 3727
rect 3293 3673 3307 3687
rect 3333 3673 3347 3687
rect 3253 3633 3267 3647
rect 3273 3633 3287 3647
rect 3173 3573 3187 3587
rect 3193 3513 3207 3527
rect 3173 3493 3187 3507
rect 3213 3493 3227 3507
rect 3193 3473 3207 3487
rect 3253 3493 3267 3507
rect 3233 3473 3247 3487
rect 3253 3453 3267 3467
rect 3153 3393 3167 3407
rect 3113 3333 3127 3347
rect 3133 3333 3147 3347
rect 3193 3333 3207 3347
rect 3233 3333 3247 3347
rect 3153 3313 3167 3327
rect 3153 3253 3167 3267
rect 3093 3173 3107 3187
rect 3093 3153 3107 3167
rect 3133 3153 3147 3167
rect 3073 3033 3087 3047
rect 3153 3073 3167 3087
rect 3133 3033 3147 3047
rect 3073 2993 3087 3007
rect 3113 2973 3127 2987
rect 3133 2913 3147 2927
rect 3133 2873 3147 2887
rect 3033 2813 3047 2827
rect 3113 2813 3127 2827
rect 3033 2773 3047 2787
rect 3073 2773 3087 2787
rect 3113 2773 3127 2787
rect 3033 2733 3047 2747
rect 3313 3573 3327 3587
rect 3333 3473 3347 3487
rect 3353 3493 3367 3507
rect 3413 3733 3427 3747
rect 3433 3713 3447 3727
rect 3453 3733 3467 3747
rect 3393 3573 3407 3587
rect 3393 3533 3407 3547
rect 3413 3533 3427 3547
rect 3373 3473 3387 3487
rect 3333 3453 3347 3467
rect 3353 3453 3367 3467
rect 3533 3953 3547 3967
rect 3573 3953 3587 3967
rect 3493 3913 3507 3927
rect 3513 3813 3527 3827
rect 3553 3753 3567 3767
rect 3573 3733 3587 3747
rect 3553 3673 3567 3687
rect 3533 3573 3547 3587
rect 3493 3533 3507 3547
rect 3513 3533 3527 3547
rect 3553 3553 3567 3567
rect 3413 3453 3427 3467
rect 3313 3393 3327 3407
rect 3293 3333 3307 3347
rect 3313 3313 3327 3327
rect 3293 3273 3307 3287
rect 3233 3253 3247 3267
rect 3193 3153 3207 3167
rect 3273 3133 3287 3147
rect 3213 3113 3227 3127
rect 3273 3073 3287 3087
rect 3253 3053 3267 3067
rect 3233 2993 3247 3007
rect 3293 2933 3307 2947
rect 3273 2833 3287 2847
rect 3293 2833 3307 2847
rect 3173 2793 3187 2807
rect 3253 2793 3267 2807
rect 3153 2773 3167 2787
rect 3213 2773 3227 2787
rect 3093 2733 3107 2747
rect 3133 2733 3147 2747
rect 3053 2673 3067 2687
rect 3173 2653 3187 2667
rect 3193 2593 3207 2607
rect 2973 2313 2987 2327
rect 2953 2113 2967 2127
rect 3033 2533 3047 2547
rect 3093 2553 3107 2567
rect 3153 2553 3167 2567
rect 3073 2453 3087 2467
rect 3013 2413 3027 2427
rect 3093 2373 3107 2387
rect 3053 2313 3067 2327
rect 3013 2293 3027 2307
rect 3033 2273 3047 2287
rect 3033 2253 3047 2267
rect 3033 2133 3047 2147
rect 3033 2053 3047 2067
rect 2953 1993 2967 2007
rect 3053 2013 3067 2027
rect 3033 1993 3047 2007
rect 3053 1993 3067 2007
rect 3013 1933 3027 1947
rect 2993 1853 3007 1867
rect 3033 1813 3047 1827
rect 2973 1793 2987 1807
rect 2953 1773 2967 1787
rect 2933 1413 2947 1427
rect 2873 1393 2887 1407
rect 2913 1373 2927 1387
rect 2853 1353 2867 1367
rect 2913 1353 2927 1367
rect 2813 1293 2827 1307
rect 2833 1293 2847 1307
rect 2873 1313 2887 1327
rect 2893 1293 2907 1307
rect 2853 1273 2867 1287
rect 2793 1213 2807 1227
rect 2813 1173 2827 1187
rect 2993 1753 3007 1767
rect 3033 1753 3047 1767
rect 2993 1633 3007 1647
rect 3073 1953 3087 1967
rect 3153 2513 3167 2527
rect 3233 2733 3247 2747
rect 3413 3433 3427 3447
rect 3353 3353 3367 3367
rect 3413 3353 3427 3367
rect 3393 3253 3407 3267
rect 3373 3233 3387 3247
rect 3333 3213 3347 3227
rect 3353 3193 3367 3207
rect 3353 3153 3367 3167
rect 3333 3113 3347 3127
rect 3393 3073 3407 3087
rect 3373 3033 3387 3047
rect 3393 3013 3407 3027
rect 3393 2993 3407 3007
rect 3373 2933 3387 2947
rect 3313 2773 3327 2787
rect 3373 2773 3387 2787
rect 3313 2733 3327 2747
rect 3333 2753 3347 2767
rect 3253 2713 3267 2727
rect 3353 2713 3367 2727
rect 3293 2673 3307 2687
rect 3313 2673 3327 2687
rect 3233 2593 3247 2607
rect 3193 2553 3207 2567
rect 3273 2553 3287 2567
rect 3173 2493 3187 2507
rect 3213 2513 3227 2527
rect 3253 2513 3267 2527
rect 3273 2513 3287 2527
rect 3213 2493 3227 2507
rect 3193 2473 3207 2487
rect 3193 2413 3207 2427
rect 3193 2353 3207 2367
rect 3173 2333 3187 2347
rect 3193 2333 3207 2347
rect 3293 2453 3307 2467
rect 3253 2393 3267 2407
rect 3233 2353 3247 2367
rect 3193 2253 3207 2267
rect 3213 2253 3227 2267
rect 3113 2233 3127 2247
rect 3153 2233 3167 2247
rect 3193 2233 3207 2247
rect 3133 2173 3147 2187
rect 3173 2093 3187 2107
rect 3213 2073 3227 2087
rect 3193 2033 3207 2047
rect 3173 1933 3187 1947
rect 3153 1873 3167 1887
rect 3093 1813 3107 1827
rect 3113 1813 3127 1827
rect 3093 1773 3107 1787
rect 3073 1733 3087 1747
rect 3033 1613 3047 1627
rect 3053 1613 3067 1627
rect 2973 1573 2987 1587
rect 2973 1533 2987 1547
rect 3013 1513 3027 1527
rect 3033 1373 3047 1387
rect 2993 1353 3007 1367
rect 2973 1293 2987 1307
rect 3113 1753 3127 1767
rect 3173 1713 3187 1727
rect 3473 3493 3487 3507
rect 3513 3493 3527 3507
rect 3453 3473 3467 3487
rect 3493 3473 3507 3487
rect 3493 3433 3507 3447
rect 3453 3413 3467 3427
rect 3553 3373 3567 3387
rect 3613 4153 3627 4167
rect 3653 4153 3667 4167
rect 3773 4613 3787 4627
rect 3813 4553 3827 4567
rect 3753 4453 3767 4467
rect 3793 4473 3807 4487
rect 3813 4453 3827 4467
rect 3773 4213 3787 4227
rect 3733 4173 3747 4187
rect 3633 4073 3647 4087
rect 3713 4073 3727 4087
rect 3733 4073 3747 4087
rect 3713 4053 3727 4067
rect 3793 4193 3807 4207
rect 3853 4673 3867 4687
rect 3893 4633 3907 4647
rect 3893 4613 3907 4627
rect 4033 5173 4047 5187
rect 3993 5153 4007 5167
rect 4013 5113 4027 5127
rect 3993 5073 4007 5087
rect 4013 4973 4027 4987
rect 4053 5153 4067 5167
rect 4093 5053 4107 5067
rect 4053 4953 4067 4967
rect 4033 4913 4047 4927
rect 4073 4913 4087 4927
rect 3973 4853 3987 4867
rect 3953 4793 3967 4807
rect 3953 4693 3967 4707
rect 3933 4593 3947 4607
rect 3933 4553 3947 4567
rect 3893 4493 3907 4507
rect 3853 4453 3867 4467
rect 3873 4433 3887 4447
rect 3913 4253 3927 4267
rect 4013 4693 4027 4707
rect 3993 4653 4007 4667
rect 3973 4233 3987 4247
rect 3913 4213 3927 4227
rect 3833 4193 3847 4207
rect 3933 4193 3947 4207
rect 3973 4173 3987 4187
rect 4073 4633 4087 4647
rect 4033 4593 4047 4607
rect 4013 4493 4027 4507
rect 4213 5353 4227 5367
rect 4273 5333 4287 5347
rect 4253 5173 4267 5187
rect 4193 5133 4207 5147
rect 4213 5153 4227 5167
rect 4253 5133 4267 5147
rect 4173 5113 4187 5127
rect 4133 5013 4147 5027
rect 4133 4973 4147 4987
rect 4233 5033 4247 5047
rect 4233 5013 4247 5027
rect 4113 4913 4127 4927
rect 4193 4933 4207 4947
rect 4173 4913 4187 4927
rect 4213 4913 4227 4927
rect 4153 4753 4167 4767
rect 4173 4693 4187 4707
rect 4173 4673 4187 4687
rect 4133 4633 4147 4647
rect 4173 4633 4187 4647
rect 4413 5213 4427 5227
rect 4293 5153 4307 5167
rect 4333 5153 4347 5167
rect 4353 5133 4367 5147
rect 4373 5133 4387 5147
rect 4313 5113 4327 5127
rect 4393 5073 4407 5087
rect 4373 4973 4387 4987
rect 4273 4953 4287 4967
rect 4293 4953 4307 4967
rect 4273 4893 4287 4907
rect 4273 4873 4287 4887
rect 4273 4713 4287 4727
rect 4353 4913 4367 4927
rect 4373 4913 4387 4927
rect 4333 4813 4347 4827
rect 4293 4673 4307 4687
rect 4333 4673 4347 4687
rect 4253 4613 4267 4627
rect 4233 4593 4247 4607
rect 4233 4573 4247 4587
rect 4113 4533 4127 4547
rect 4053 4513 4067 4527
rect 4093 4513 4107 4527
rect 4113 4493 4127 4507
rect 4033 4433 4047 4447
rect 4153 4413 4167 4427
rect 4033 4233 4047 4247
rect 3993 4153 4007 4167
rect 3873 4073 3887 4087
rect 3793 4053 3807 4067
rect 3773 4033 3787 4047
rect 3753 3993 3767 4007
rect 3673 3953 3687 3967
rect 3713 3933 3727 3947
rect 3633 3793 3647 3807
rect 3713 3733 3727 3747
rect 3633 3693 3647 3707
rect 3613 3673 3627 3687
rect 3633 3613 3647 3627
rect 3613 3573 3627 3587
rect 3693 3693 3707 3707
rect 3673 3633 3687 3647
rect 3673 3613 3687 3627
rect 3653 3553 3667 3567
rect 3693 3533 3707 3547
rect 3653 3493 3667 3507
rect 3593 3393 3607 3407
rect 3573 3313 3587 3327
rect 3453 3273 3467 3287
rect 3433 3173 3447 3187
rect 3433 3113 3447 3127
rect 3473 3253 3487 3267
rect 3473 3133 3487 3147
rect 3453 2993 3467 3007
rect 3433 2953 3447 2967
rect 3533 3233 3547 3247
rect 3533 3213 3547 3227
rect 3513 3153 3527 3167
rect 3553 3193 3567 3207
rect 3673 3453 3687 3467
rect 3613 3273 3627 3287
rect 3693 3413 3707 3427
rect 3693 3393 3707 3407
rect 3673 3253 3687 3267
rect 3593 3233 3607 3247
rect 3633 3233 3647 3247
rect 3653 3213 3667 3227
rect 3693 3213 3707 3227
rect 3693 3193 3707 3207
rect 3613 3153 3627 3167
rect 3573 3133 3587 3147
rect 3613 3133 3627 3147
rect 3493 3033 3507 3047
rect 3553 3033 3567 3047
rect 3513 2993 3527 3007
rect 3533 2993 3547 3007
rect 3473 2793 3487 2807
rect 3513 2793 3527 2807
rect 3413 2773 3427 2787
rect 3433 2773 3447 2787
rect 3433 2733 3447 2747
rect 3413 2713 3427 2727
rect 3393 2673 3407 2687
rect 3333 2653 3347 2667
rect 3373 2653 3387 2667
rect 3373 2553 3387 2567
rect 3453 2693 3467 2707
rect 3353 2513 3367 2527
rect 3393 2513 3407 2527
rect 3433 2513 3447 2527
rect 3353 2493 3367 2507
rect 3333 2473 3347 2487
rect 3333 2353 3347 2367
rect 3273 2293 3287 2307
rect 3313 2293 3327 2307
rect 3253 2273 3267 2287
rect 3273 2253 3287 2267
rect 3293 2273 3307 2287
rect 3313 2213 3327 2227
rect 3433 2453 3447 2467
rect 3393 2433 3407 2447
rect 3413 2433 3427 2447
rect 3373 2353 3387 2367
rect 3373 2293 3387 2307
rect 3393 2293 3407 2307
rect 3253 2173 3267 2187
rect 3333 2173 3347 2187
rect 3353 2173 3367 2187
rect 3293 2113 3307 2127
rect 3313 2113 3327 2127
rect 3273 2093 3287 2107
rect 3253 2073 3267 2087
rect 3233 2053 3247 2067
rect 3273 2053 3287 2067
rect 3253 1973 3267 1987
rect 3213 1793 3227 1807
rect 3193 1673 3207 1687
rect 3353 2093 3367 2107
rect 3313 2033 3327 2047
rect 3333 2033 3347 2047
rect 3313 1813 3327 1827
rect 3293 1773 3307 1787
rect 3293 1733 3307 1747
rect 3253 1713 3267 1727
rect 3513 2733 3527 2747
rect 3493 2713 3507 2727
rect 3473 2673 3487 2687
rect 3473 2653 3487 2667
rect 3473 2553 3487 2567
rect 3473 2473 3487 2487
rect 3453 2353 3467 2367
rect 3413 2273 3427 2287
rect 3473 2313 3487 2327
rect 3393 2213 3407 2227
rect 3393 2173 3407 2187
rect 3413 2173 3427 2187
rect 3433 2153 3447 2167
rect 3373 1833 3387 1847
rect 3373 1813 3387 1827
rect 3413 1813 3427 1827
rect 3353 1773 3367 1787
rect 3313 1673 3327 1687
rect 3113 1593 3127 1607
rect 3113 1573 3127 1587
rect 3113 1533 3127 1547
rect 3213 1653 3227 1667
rect 3233 1653 3247 1667
rect 3133 1513 3147 1527
rect 3233 1633 3247 1647
rect 3233 1573 3247 1587
rect 3393 1793 3407 1807
rect 3393 1753 3407 1767
rect 3413 1693 3427 1707
rect 3693 3113 3707 3127
rect 3653 3053 3667 3067
rect 3633 3033 3647 3047
rect 3673 2993 3687 3007
rect 3733 3713 3747 3727
rect 3733 3653 3747 3667
rect 3833 3973 3847 3987
rect 3893 4033 3907 4047
rect 3853 3933 3867 3947
rect 3773 3913 3787 3927
rect 3813 3833 3827 3847
rect 3833 3753 3847 3767
rect 3773 3733 3787 3747
rect 3793 3653 3807 3667
rect 3833 3653 3847 3667
rect 3773 3573 3787 3587
rect 3713 2833 3727 2847
rect 3753 3513 3767 3527
rect 3773 3473 3787 3487
rect 3833 3493 3847 3507
rect 3793 3453 3807 3467
rect 3833 3393 3847 3407
rect 3833 3233 3847 3247
rect 3833 3213 3847 3227
rect 3773 3153 3787 3167
rect 3793 3153 3807 3167
rect 3753 3053 3767 3067
rect 3773 3013 3787 3027
rect 3653 2793 3667 2807
rect 3593 2733 3607 2747
rect 3613 2733 3627 2747
rect 3573 2713 3587 2727
rect 3593 2693 3607 2707
rect 3553 2673 3567 2687
rect 3533 2653 3547 2667
rect 3573 2653 3587 2667
rect 3513 2493 3527 2507
rect 3493 2253 3507 2267
rect 3493 2233 3507 2247
rect 3473 2113 3487 2127
rect 3453 2073 3467 2087
rect 3453 1973 3467 1987
rect 3433 1553 3447 1567
rect 3253 1473 3267 1487
rect 3273 1473 3287 1487
rect 3113 1393 3127 1407
rect 3053 1353 3067 1367
rect 3193 1353 3207 1367
rect 3013 1313 3027 1327
rect 3033 1293 3047 1307
rect 3153 1313 3167 1327
rect 3133 1293 3147 1307
rect 3033 1273 3047 1287
rect 2953 1173 2967 1187
rect 2773 1093 2787 1107
rect 2893 1113 2907 1127
rect 2873 1033 2887 1047
rect 2953 1133 2967 1147
rect 2933 1113 2947 1127
rect 2993 1173 3007 1187
rect 2973 1073 2987 1087
rect 2913 973 2927 987
rect 2973 933 2987 947
rect 2933 873 2947 887
rect 2773 833 2787 847
rect 2673 813 2687 827
rect 2733 813 2747 827
rect 2853 853 2867 867
rect 2893 853 2907 867
rect 2693 773 2707 787
rect 2813 773 2827 787
rect 2653 753 2667 767
rect 2733 653 2747 667
rect 2873 653 2887 667
rect 2613 613 2627 627
rect 2593 533 2607 547
rect 2733 613 2747 627
rect 2693 533 2707 547
rect 2633 513 2647 527
rect 2593 433 2607 447
rect 2533 413 2547 427
rect 2453 333 2467 347
rect 2313 313 2327 327
rect 2353 313 2367 327
rect 2433 313 2447 327
rect 2373 293 2387 307
rect 2253 173 2267 187
rect 2133 113 2147 127
rect 193 93 207 107
rect 793 93 807 107
rect 1853 93 1867 107
rect 2093 93 2107 107
rect 2333 153 2347 167
rect 2453 153 2467 167
rect 2553 373 2567 387
rect 2533 353 2547 367
rect 2653 453 2667 467
rect 2633 393 2647 407
rect 2713 393 2727 407
rect 2673 333 2687 347
rect 2693 333 2707 347
rect 2573 313 2587 327
rect 2633 293 2647 307
rect 2833 613 2847 627
rect 2793 573 2807 587
rect 2773 513 2787 527
rect 2793 513 2807 527
rect 3053 1133 3067 1147
rect 3073 1113 3087 1127
rect 3113 1113 3127 1127
rect 3093 1073 3107 1087
rect 3193 1233 3207 1247
rect 3173 1213 3187 1227
rect 3153 1153 3167 1167
rect 3153 1073 3167 1087
rect 3133 1053 3147 1067
rect 3113 873 3127 887
rect 3013 833 3027 847
rect 3053 833 3067 847
rect 2953 793 2967 807
rect 2993 793 3007 807
rect 2913 453 2927 467
rect 2833 413 2847 427
rect 2733 353 2747 367
rect 2753 333 2767 347
rect 2513 193 2527 207
rect 2713 193 2727 207
rect 2653 173 2667 187
rect 2613 153 2627 167
rect 2633 133 2647 147
rect 2873 373 2887 387
rect 2873 333 2887 347
rect 2933 333 2947 347
rect 2833 313 2847 327
rect 2893 313 2907 327
rect 2913 313 2927 327
rect 2673 133 2687 147
rect 2713 133 2727 147
rect 2393 113 2407 127
rect 2473 113 2487 127
rect 2913 153 2927 167
rect 2833 133 2847 147
rect 2933 113 2947 127
rect 2773 93 2787 107
rect 2893 93 2907 107
rect 2273 33 2287 47
rect 2673 33 2687 47
rect 2633 13 2647 27
rect 3033 633 3047 647
rect 2973 593 2987 607
rect 2993 613 3007 627
rect 3013 593 3027 607
rect 2973 533 2987 547
rect 3013 353 3027 367
rect 2993 313 3007 327
rect 3133 833 3147 847
rect 3173 833 3187 847
rect 3113 793 3127 807
rect 3153 793 3167 807
rect 3093 653 3107 667
rect 3073 613 3087 627
rect 3113 613 3127 627
rect 3133 633 3147 647
rect 3153 633 3167 647
rect 3093 573 3107 587
rect 3053 393 3067 407
rect 3213 1173 3227 1187
rect 3293 1393 3307 1407
rect 3273 1273 3287 1287
rect 3313 1273 3327 1287
rect 3433 1493 3447 1507
rect 3413 1293 3427 1307
rect 3373 1233 3387 1247
rect 3413 1213 3427 1227
rect 3373 1153 3387 1167
rect 3253 1133 3267 1147
rect 3393 1133 3407 1147
rect 3233 1093 3247 1107
rect 3193 653 3207 667
rect 3313 1113 3327 1127
rect 3273 1053 3287 1067
rect 3253 913 3267 927
rect 3293 853 3307 867
rect 3273 773 3287 787
rect 3333 1033 3347 1047
rect 3633 2673 3647 2687
rect 3733 2793 3747 2807
rect 3693 2773 3707 2787
rect 3713 2753 3727 2767
rect 3753 2753 3767 2767
rect 3673 2733 3687 2747
rect 3733 2733 3747 2747
rect 3673 2713 3687 2727
rect 3653 2553 3667 2567
rect 3613 2513 3627 2527
rect 3573 2473 3587 2487
rect 3573 2293 3587 2307
rect 3533 2253 3547 2267
rect 3573 2253 3587 2267
rect 3513 2193 3527 2207
rect 3593 2173 3607 2187
rect 3533 2093 3547 2107
rect 3573 2093 3587 2107
rect 3513 2053 3527 2067
rect 3553 2053 3567 2067
rect 3693 2673 3707 2687
rect 3673 2493 3687 2507
rect 3653 2473 3667 2487
rect 3673 2393 3687 2407
rect 3633 2373 3647 2387
rect 3653 2373 3667 2387
rect 3633 2253 3647 2267
rect 3773 2733 3787 2747
rect 3713 2573 3727 2587
rect 3753 2573 3767 2587
rect 3833 3053 3847 3067
rect 3813 3033 3827 3047
rect 3833 3013 3847 3027
rect 3813 2933 3827 2947
rect 3833 2893 3847 2907
rect 3933 3993 3947 4007
rect 3973 3993 3987 4007
rect 3893 3813 3907 3827
rect 3913 3773 3927 3787
rect 3893 3633 3907 3647
rect 3893 3613 3907 3627
rect 3873 3593 3887 3607
rect 3873 3513 3887 3527
rect 3913 3513 3927 3527
rect 3913 3373 3927 3387
rect 3893 3233 3907 3247
rect 3873 3193 3887 3207
rect 3913 3193 3927 3207
rect 3913 3173 3927 3187
rect 3873 3073 3887 3087
rect 3873 3033 3887 3047
rect 3893 3033 3907 3047
rect 3893 2993 3907 3007
rect 3873 2973 3887 2987
rect 3853 2813 3867 2827
rect 3873 2813 3887 2827
rect 3813 2773 3827 2787
rect 3793 2693 3807 2707
rect 3833 2633 3847 2647
rect 3833 2613 3847 2627
rect 3813 2573 3827 2587
rect 3793 2533 3807 2547
rect 3733 2513 3747 2527
rect 3753 2513 3767 2527
rect 3793 2513 3807 2527
rect 3713 2433 3727 2447
rect 3693 2373 3707 2387
rect 3773 2473 3787 2487
rect 3753 2353 3767 2367
rect 3733 2273 3747 2287
rect 3673 2253 3687 2267
rect 3693 2253 3707 2267
rect 3653 2233 3667 2247
rect 3653 2213 3667 2227
rect 3633 2073 3647 2087
rect 3553 2033 3567 2047
rect 3613 2033 3627 2047
rect 3593 2013 3607 2027
rect 3493 1913 3507 1927
rect 3533 1913 3547 1927
rect 3493 1853 3507 1867
rect 3573 1813 3587 1827
rect 3493 1793 3507 1807
rect 3473 1733 3487 1747
rect 3473 1693 3487 1707
rect 3473 1553 3487 1567
rect 3473 1533 3487 1547
rect 3453 1453 3467 1467
rect 3453 1373 3467 1387
rect 3453 1293 3467 1307
rect 3453 1273 3467 1287
rect 3433 1193 3447 1207
rect 3433 1133 3447 1147
rect 3433 1013 3447 1027
rect 3413 833 3427 847
rect 3393 813 3407 827
rect 3333 793 3347 807
rect 3413 793 3427 807
rect 3433 773 3447 787
rect 3373 653 3387 667
rect 3413 653 3427 667
rect 3173 613 3187 627
rect 3153 533 3167 547
rect 3173 453 3187 467
rect 3133 413 3147 427
rect 3233 593 3247 607
rect 3253 613 3267 627
rect 3293 613 3307 627
rect 3253 553 3267 567
rect 3213 393 3227 407
rect 3333 613 3347 627
rect 3313 413 3327 427
rect 3153 353 3167 367
rect 3173 353 3187 367
rect 3253 353 3267 367
rect 3153 313 3167 327
rect 3273 313 3287 327
rect 3353 593 3367 607
rect 3353 553 3367 567
rect 3413 393 3427 407
rect 3553 1673 3567 1687
rect 3553 1613 3567 1627
rect 3533 1593 3547 1607
rect 3513 1533 3527 1547
rect 3533 1533 3547 1547
rect 3513 1513 3527 1527
rect 3493 1373 3507 1387
rect 3493 1213 3507 1227
rect 3473 1193 3487 1207
rect 3493 1173 3507 1187
rect 3533 1473 3547 1487
rect 3533 1433 3547 1447
rect 3533 1293 3547 1307
rect 3673 2093 3687 2107
rect 3653 2013 3667 2027
rect 3713 2053 3727 2067
rect 3673 1993 3687 2007
rect 3713 1973 3727 1987
rect 3633 1933 3647 1947
rect 3613 1893 3627 1907
rect 3613 1833 3627 1847
rect 3613 1773 3627 1787
rect 3693 1893 3707 1907
rect 3713 1773 3727 1787
rect 3633 1753 3647 1767
rect 3653 1753 3667 1767
rect 3653 1733 3667 1747
rect 3633 1713 3647 1727
rect 3693 1713 3707 1727
rect 3673 1673 3687 1687
rect 3593 1613 3607 1627
rect 3673 1613 3687 1627
rect 3593 1593 3607 1607
rect 3653 1573 3667 1587
rect 3613 1553 3627 1567
rect 3593 1533 3607 1547
rect 3573 1253 3587 1267
rect 3733 1653 3747 1667
rect 3813 2493 3827 2507
rect 3813 2413 3827 2427
rect 3793 2293 3807 2307
rect 3773 2233 3787 2247
rect 3793 2193 3807 2207
rect 3853 2573 3867 2587
rect 3853 2533 3867 2547
rect 3853 2513 3867 2527
rect 3853 2333 3867 2347
rect 3833 2293 3847 2307
rect 3833 2233 3847 2247
rect 3773 2173 3787 2187
rect 3813 2173 3827 2187
rect 3953 3973 3967 3987
rect 3993 3973 4007 3987
rect 4013 3993 4027 4007
rect 4093 4233 4107 4247
rect 4053 4213 4067 4227
rect 4133 4213 4147 4227
rect 4053 4173 4067 4187
rect 3993 3953 4007 3967
rect 4033 3953 4047 3967
rect 4013 3713 4027 3727
rect 4313 4533 4327 4547
rect 4253 4473 4267 4487
rect 4233 4293 4247 4307
rect 4173 4253 4187 4267
rect 4193 4253 4207 4267
rect 4193 4193 4207 4207
rect 4193 4173 4207 4187
rect 4233 4173 4247 4187
rect 4153 4093 4167 4107
rect 4093 4053 4107 4067
rect 4133 4053 4147 4067
rect 4173 4053 4187 4067
rect 4133 4033 4147 4047
rect 4073 3993 4087 4007
rect 4113 3973 4127 3987
rect 4273 4433 4287 4447
rect 4293 4453 4307 4467
rect 4353 4453 4367 4467
rect 4273 4393 4287 4407
rect 4313 4393 4327 4407
rect 4333 4393 4347 4407
rect 4273 4373 4287 4387
rect 4253 4033 4267 4047
rect 4233 3973 4247 3987
rect 4193 3933 4207 3947
rect 4213 3933 4227 3947
rect 4253 3833 4267 3847
rect 3993 3633 4007 3647
rect 3973 3613 3987 3627
rect 3993 3513 4007 3527
rect 3973 3473 3987 3487
rect 3993 3373 4007 3387
rect 3953 3253 3967 3267
rect 3953 3233 3967 3247
rect 4073 3693 4087 3707
rect 4133 3713 4147 3727
rect 4213 3693 4227 3707
rect 4133 3653 4147 3667
rect 4033 3613 4047 3627
rect 4153 3593 4167 3607
rect 4193 3573 4207 3587
rect 4193 3553 4207 3567
rect 4053 3533 4067 3547
rect 4153 3533 4167 3547
rect 4033 3493 4047 3507
rect 4113 3493 4127 3507
rect 4173 3493 4187 3507
rect 4013 3353 4027 3367
rect 4013 3253 4027 3267
rect 3993 3153 4007 3167
rect 3933 3133 3947 3147
rect 3973 3133 3987 3147
rect 3933 3033 3947 3047
rect 3953 2973 3967 2987
rect 3993 3053 4007 3067
rect 3993 3033 4007 3047
rect 4033 3153 4047 3167
rect 4173 3473 4187 3487
rect 4073 3453 4087 3467
rect 4153 3333 4167 3347
rect 4133 3313 4147 3327
rect 4093 3233 4107 3247
rect 4073 3173 4087 3187
rect 4073 3113 4087 3127
rect 4053 3053 4067 3067
rect 4093 3053 4107 3067
rect 4033 3033 4047 3047
rect 4013 2893 4027 2907
rect 4013 2873 4027 2887
rect 3933 2793 3947 2807
rect 3973 2793 3987 2807
rect 3993 2793 4007 2807
rect 3913 2693 3927 2707
rect 3913 2573 3927 2587
rect 3893 2553 3907 2567
rect 3993 2773 4007 2787
rect 4013 2773 4027 2787
rect 3973 2753 3987 2767
rect 3993 2673 4007 2687
rect 3973 2653 3987 2667
rect 3953 2633 3967 2647
rect 3913 2533 3927 2547
rect 3893 2273 3907 2287
rect 3793 2073 3807 2087
rect 3833 2073 3847 2087
rect 3833 2053 3847 2067
rect 3813 2033 3827 2047
rect 3773 2013 3787 2027
rect 3793 1873 3807 1887
rect 3773 1773 3787 1787
rect 3773 1733 3787 1747
rect 3753 1633 3767 1647
rect 3753 1613 3767 1627
rect 3713 1593 3727 1607
rect 3693 1573 3707 1587
rect 3733 1573 3747 1587
rect 3773 1573 3787 1587
rect 3673 1553 3687 1567
rect 3733 1533 3747 1547
rect 3853 1833 3867 1847
rect 3833 1773 3847 1787
rect 3813 1753 3827 1767
rect 3833 1593 3847 1607
rect 3933 2493 3947 2507
rect 3953 2333 3967 2347
rect 4113 2973 4127 2987
rect 4093 2753 4107 2767
rect 4073 2713 4087 2727
rect 4113 2713 4127 2727
rect 4413 4933 4427 4947
rect 4493 5453 4507 5467
rect 4573 5593 4587 5607
rect 4813 5593 4827 5607
rect 4853 5593 4867 5607
rect 4573 5513 4587 5527
rect 4553 5493 4567 5507
rect 4713 5493 4727 5507
rect 4473 5413 4487 5427
rect 4513 5413 4527 5427
rect 4593 5433 4607 5447
rect 4753 5453 4767 5467
rect 4633 5413 4647 5427
rect 4513 5393 4527 5407
rect 4553 5393 4567 5407
rect 4733 5393 4747 5407
rect 4473 5353 4487 5367
rect 4473 5153 4487 5167
rect 4533 5133 4547 5147
rect 4453 5113 4467 5127
rect 4453 4973 4467 4987
rect 4493 4953 4507 4967
rect 4433 4873 4447 4887
rect 4673 5253 4687 5267
rect 4573 5193 4587 5207
rect 4593 5133 4607 5147
rect 4633 5153 4647 5167
rect 4653 5133 4667 5147
rect 4613 5113 4627 5127
rect 4613 5033 4627 5047
rect 4653 5033 4667 5047
rect 4593 4973 4607 4987
rect 4633 4953 4647 4967
rect 4693 5153 4707 5167
rect 4733 5153 4747 5167
rect 4793 5353 4807 5367
rect 4713 5113 4727 5127
rect 4753 5113 4767 5127
rect 4713 5033 4727 5047
rect 4553 4913 4567 4927
rect 4613 4913 4627 4927
rect 4613 4833 4627 4847
rect 4493 4813 4507 4827
rect 4593 4813 4607 4827
rect 4413 4713 4427 4727
rect 4493 4713 4507 4727
rect 4413 4693 4427 4707
rect 4433 4673 4447 4687
rect 4473 4673 4487 4687
rect 4453 4633 4467 4647
rect 4473 4533 4487 4547
rect 4473 4513 4487 4527
rect 4393 4473 4407 4487
rect 4413 4473 4427 4487
rect 4393 4453 4407 4467
rect 4433 4433 4447 4447
rect 4373 4413 4387 4427
rect 4533 4673 4547 4687
rect 4533 4593 4547 4607
rect 4573 4653 4587 4667
rect 4593 4633 4607 4647
rect 4553 4573 4567 4587
rect 4493 4433 4507 4447
rect 4513 4433 4527 4447
rect 4313 4173 4327 4187
rect 4333 4193 4347 4207
rect 4393 4173 4407 4187
rect 4373 4153 4387 4167
rect 4433 4173 4447 4187
rect 4473 4193 4487 4207
rect 4413 4153 4427 4167
rect 4693 4733 4707 4747
rect 4693 4673 4707 4687
rect 4673 4633 4687 4647
rect 4613 4353 4627 4367
rect 4653 4353 4667 4367
rect 4593 4333 4607 4347
rect 4553 4293 4567 4307
rect 4613 4293 4627 4307
rect 4553 4213 4567 4227
rect 4493 4133 4507 4147
rect 4293 4113 4307 4127
rect 4333 4113 4347 4127
rect 4393 4113 4407 4127
rect 4293 4093 4307 4107
rect 4373 4033 4387 4047
rect 4333 3993 4347 4007
rect 4353 3973 4367 3987
rect 4393 3973 4407 3987
rect 4433 3973 4447 3987
rect 4413 3893 4427 3907
rect 4333 3873 4347 3887
rect 4373 3873 4387 3887
rect 4293 3573 4307 3587
rect 4213 3533 4227 3547
rect 4213 3313 4227 3327
rect 4273 3553 4287 3567
rect 4253 3533 4267 3547
rect 4433 3733 4447 3747
rect 4373 3713 4387 3727
rect 4393 3693 4407 3707
rect 4513 3993 4527 4007
rect 4533 3993 4547 4007
rect 4473 3913 4487 3927
rect 4593 4213 4607 4227
rect 4613 4193 4627 4207
rect 4573 4113 4587 4127
rect 4693 4393 4707 4407
rect 4833 5333 4847 5347
rect 4873 5333 4887 5347
rect 4833 5133 4847 5147
rect 4873 5133 4887 5147
rect 4833 5093 4847 5107
rect 4853 5073 4867 5087
rect 5153 5753 5167 5767
rect 5133 5673 5147 5687
rect 4993 5613 5007 5627
rect 5053 5613 5067 5627
rect 4933 5593 4947 5607
rect 4913 5513 4927 5527
rect 5133 5613 5147 5627
rect 4933 5093 4947 5107
rect 4913 5053 4927 5067
rect 4893 5033 4907 5047
rect 4733 4953 4747 4967
rect 4773 4933 4787 4947
rect 4733 4633 4747 4647
rect 4893 4993 4907 5007
rect 4813 4613 4827 4627
rect 4773 4433 4787 4447
rect 4793 4413 4807 4427
rect 4733 4313 4747 4327
rect 4673 4173 4687 4187
rect 4633 4153 4647 4167
rect 4653 4153 4667 4167
rect 4593 3993 4607 4007
rect 4653 3993 4667 4007
rect 4533 3833 4547 3847
rect 4493 3753 4507 3767
rect 4433 3693 4447 3707
rect 4453 3693 4467 3707
rect 4513 3713 4527 3727
rect 4373 3673 4387 3687
rect 4413 3673 4427 3687
rect 4473 3673 4487 3687
rect 4553 3673 4567 3687
rect 4673 3953 4687 3967
rect 4753 4173 4767 4187
rect 4713 4133 4727 4147
rect 4713 4013 4727 4027
rect 4713 3913 4727 3927
rect 4753 4013 4767 4027
rect 4833 4573 4847 4587
rect 4873 4633 4887 4647
rect 4913 4953 4927 4967
rect 4953 4973 4967 4987
rect 5093 5593 5107 5607
rect 5033 5513 5047 5527
rect 5093 5473 5107 5487
rect 5133 5473 5147 5487
rect 5133 5433 5147 5447
rect 5173 5673 5187 5687
rect 5233 5773 5247 5787
rect 5393 5773 5407 5787
rect 5193 5633 5207 5647
rect 5213 5613 5227 5627
rect 5173 5433 5187 5447
rect 5113 5353 5127 5367
rect 5073 5173 5087 5187
rect 5073 5113 5087 5127
rect 5053 5073 5067 5087
rect 4973 4913 4987 4927
rect 5013 4993 5027 5007
rect 5013 4953 5027 4967
rect 5053 4953 5067 4967
rect 5053 4873 5067 4887
rect 5153 5393 5167 5407
rect 5133 5093 5147 5107
rect 5133 4973 5147 4987
rect 5173 5333 5187 5347
rect 5093 4953 5107 4967
rect 5153 4953 5167 4967
rect 5153 4933 5167 4947
rect 5133 4913 5147 4927
rect 5073 4793 5087 4807
rect 4953 4713 4967 4727
rect 5053 4713 5067 4727
rect 4953 4653 4967 4667
rect 5013 4653 5027 4667
rect 5033 4673 5047 4687
rect 5073 4673 5087 4687
rect 4933 4613 4947 4627
rect 4893 4593 4907 4607
rect 4853 4493 4867 4507
rect 4873 4473 4887 4487
rect 4933 4473 4947 4487
rect 4813 4133 4827 4147
rect 4753 3953 4767 3967
rect 4773 3953 4787 3967
rect 4813 3953 4827 3967
rect 4733 3893 4747 3907
rect 4813 3853 4827 3867
rect 4593 3793 4607 3807
rect 4693 3813 4707 3827
rect 4673 3793 4687 3807
rect 4633 3713 4647 3727
rect 4653 3693 4667 3707
rect 4753 3773 4767 3787
rect 4733 3693 4747 3707
rect 4793 3713 4807 3727
rect 4353 3573 4367 3587
rect 4273 3493 4287 3507
rect 4313 3513 4327 3527
rect 4313 3493 4327 3507
rect 4233 3253 4247 3267
rect 4293 3253 4307 3267
rect 4193 3233 4207 3247
rect 4173 3113 4187 3127
rect 4233 3233 4247 3247
rect 4213 3193 4227 3207
rect 4573 3533 4587 3547
rect 4393 3493 4407 3507
rect 4433 3493 4447 3507
rect 4473 3493 4487 3507
rect 4493 3493 4507 3507
rect 4453 3473 4467 3487
rect 4373 3453 4387 3467
rect 4353 3413 4367 3427
rect 4373 3233 4387 3247
rect 4413 3233 4427 3247
rect 4253 3173 4267 3187
rect 4333 3173 4347 3187
rect 4273 3133 4287 3147
rect 4253 3113 4267 3127
rect 4193 3093 4207 3107
rect 4213 3073 4227 3087
rect 4153 3033 4167 3047
rect 4213 3033 4227 3047
rect 4193 2993 4207 3007
rect 4233 2973 4247 2987
rect 4253 2813 4267 2827
rect 4153 2773 4167 2787
rect 4173 2773 4187 2787
rect 4193 2753 4207 2767
rect 4213 2773 4227 2787
rect 4253 2773 4267 2787
rect 4233 2753 4247 2767
rect 4253 2733 4267 2747
rect 4233 2713 4247 2727
rect 4053 2693 4067 2707
rect 4093 2693 4107 2707
rect 4133 2693 4147 2707
rect 4073 2533 4087 2547
rect 4033 2513 4047 2527
rect 4013 2473 4027 2487
rect 4253 2533 4267 2547
rect 4093 2393 4107 2407
rect 3993 2353 4007 2367
rect 3953 2153 3967 2167
rect 3973 2073 3987 2087
rect 4013 2293 4027 2307
rect 4173 2253 4187 2267
rect 4153 2233 4167 2247
rect 4033 2153 4047 2167
rect 4013 2073 4027 2087
rect 3993 2053 4007 2067
rect 4013 2053 4027 2067
rect 3933 2033 3947 2047
rect 3913 1993 3927 2007
rect 3933 1993 3947 2007
rect 4053 2113 4067 2127
rect 4073 2093 4087 2107
rect 4053 2033 4067 2047
rect 4033 1873 4047 1887
rect 4053 1873 4067 1887
rect 4013 1833 4027 1847
rect 3953 1813 3967 1827
rect 3933 1773 3947 1787
rect 3953 1793 3967 1807
rect 3993 1793 4007 1807
rect 3993 1773 4007 1787
rect 3953 1733 3967 1747
rect 3893 1693 3907 1707
rect 3913 1653 3927 1667
rect 3873 1593 3887 1607
rect 3893 1573 3907 1587
rect 3853 1513 3867 1527
rect 3793 1413 3807 1427
rect 3833 1413 3847 1427
rect 3653 1393 3667 1407
rect 3693 1393 3707 1407
rect 3733 1373 3747 1387
rect 3773 1373 3787 1387
rect 3693 1313 3707 1327
rect 3673 1273 3687 1287
rect 3753 1293 3767 1307
rect 3733 1273 3747 1287
rect 3713 1253 3727 1267
rect 3793 1253 3807 1267
rect 3633 1193 3647 1207
rect 3593 1173 3607 1187
rect 3553 1153 3567 1167
rect 3533 1133 3547 1147
rect 3513 993 3527 1007
rect 3493 973 3507 987
rect 3473 853 3487 867
rect 3473 833 3487 847
rect 3453 353 3467 367
rect 3333 313 3347 327
rect 3433 293 3447 307
rect 3313 193 3327 207
rect 3033 173 3047 187
rect 3193 173 3207 187
rect 2993 113 3007 127
rect 3053 133 3067 147
rect 3073 113 3087 127
rect 3173 133 3187 147
rect 3373 193 3387 207
rect 3213 133 3227 147
rect 3293 133 3307 147
rect 3333 133 3347 147
rect 3393 133 3407 147
rect 3413 153 3427 167
rect 3433 133 3447 147
rect 3153 93 3167 107
rect 2953 13 2967 27
rect 3593 1113 3607 1127
rect 3573 1093 3587 1107
rect 3613 1093 3627 1107
rect 3813 1213 3827 1227
rect 3713 1193 3727 1207
rect 3773 1193 3787 1207
rect 3673 1173 3687 1187
rect 3653 1093 3667 1107
rect 3593 1073 3607 1087
rect 3533 913 3547 927
rect 3513 813 3527 827
rect 3533 793 3547 807
rect 3553 793 3567 807
rect 3553 673 3567 687
rect 3653 1033 3667 1047
rect 3653 913 3667 927
rect 3693 1113 3707 1127
rect 3793 1173 3807 1187
rect 3733 1113 3747 1127
rect 3973 1693 3987 1707
rect 3993 1653 4007 1667
rect 3973 1613 3987 1627
rect 3953 1413 3967 1427
rect 3913 1353 3927 1367
rect 3893 1213 3907 1227
rect 3853 1173 3867 1187
rect 3853 1133 3867 1147
rect 3693 1073 3707 1087
rect 3793 1073 3807 1087
rect 3753 1033 3767 1047
rect 3693 973 3707 987
rect 3793 933 3807 947
rect 3893 1113 3907 1127
rect 3833 1073 3847 1087
rect 3873 1073 3887 1087
rect 3713 853 3727 867
rect 3673 833 3687 847
rect 3673 793 3687 807
rect 3513 633 3527 647
rect 3493 613 3507 627
rect 3533 613 3547 627
rect 3553 633 3567 647
rect 3493 433 3507 447
rect 3633 653 3647 667
rect 3593 633 3607 647
rect 3613 633 3627 647
rect 3673 633 3687 647
rect 3653 593 3667 607
rect 3493 393 3507 407
rect 3573 393 3587 407
rect 3593 393 3607 407
rect 3533 373 3547 387
rect 3693 613 3707 627
rect 3693 453 3707 467
rect 3673 373 3687 387
rect 3813 893 3827 907
rect 3733 833 3747 847
rect 3793 833 3807 847
rect 3753 793 3767 807
rect 3793 793 3807 807
rect 3793 713 3807 727
rect 3853 933 3867 947
rect 3873 893 3887 907
rect 3913 1093 3927 1107
rect 3993 1593 4007 1607
rect 4013 1593 4027 1607
rect 4093 2073 4107 2087
rect 4133 2073 4147 2087
rect 4253 2333 4267 2347
rect 4373 3173 4387 3187
rect 4333 3093 4347 3107
rect 4353 3093 4367 3107
rect 4293 3053 4307 3067
rect 4293 2793 4307 2807
rect 4353 3053 4367 3067
rect 4413 3173 4427 3187
rect 4413 3153 4427 3167
rect 4393 3053 4407 3067
rect 4453 3233 4467 3247
rect 4513 3473 4527 3487
rect 4533 3493 4547 3507
rect 4513 3453 4527 3467
rect 4453 3113 4467 3127
rect 4433 3093 4447 3107
rect 4433 3033 4447 3047
rect 4353 2993 4367 3007
rect 4373 2993 4387 3007
rect 4313 2433 4327 2447
rect 4413 2933 4427 2947
rect 4413 2753 4427 2767
rect 4393 2713 4407 2727
rect 4273 2273 4287 2287
rect 4253 2093 4267 2107
rect 4113 2033 4127 2047
rect 4093 1933 4107 1947
rect 4153 1913 4167 1927
rect 4133 1893 4147 1907
rect 4113 1833 4127 1847
rect 4113 1793 4127 1807
rect 4133 1813 4147 1827
rect 4213 2073 4227 2087
rect 4193 2053 4207 2067
rect 4173 1873 4187 1887
rect 4173 1833 4187 1847
rect 4153 1773 4167 1787
rect 4093 1693 4107 1707
rect 4073 1673 4087 1687
rect 4073 1633 4087 1647
rect 4013 1473 4027 1487
rect 4073 1353 4087 1367
rect 4133 1593 4147 1607
rect 4153 1553 4167 1567
rect 4113 1513 4127 1527
rect 4253 2053 4267 2067
rect 4273 2013 4287 2027
rect 4413 2433 4427 2447
rect 4413 2393 4427 2407
rect 4373 2313 4387 2327
rect 4353 2273 4367 2287
rect 4393 2253 4407 2267
rect 4373 2213 4387 2227
rect 4293 1973 4307 1987
rect 4293 1953 4307 1967
rect 4473 3033 4487 3047
rect 4453 2833 4467 2847
rect 4633 3673 4647 3687
rect 4753 3653 4767 3667
rect 4673 3593 4687 3607
rect 4733 3593 4747 3607
rect 4613 3513 4627 3527
rect 4653 3553 4667 3567
rect 4613 3453 4627 3467
rect 4593 3373 4607 3387
rect 4553 3273 4567 3287
rect 4573 3273 4587 3287
rect 4593 3213 4607 3227
rect 4573 3193 4587 3207
rect 4553 3173 4567 3187
rect 4673 3533 4687 3547
rect 4693 3533 4707 3547
rect 4653 3193 4667 3207
rect 4713 3273 4727 3287
rect 4773 3593 4787 3607
rect 4893 4433 4907 4447
rect 4933 4433 4947 4447
rect 4933 4393 4947 4407
rect 4913 4293 4927 4307
rect 4853 4153 4867 4167
rect 4873 4153 4887 4167
rect 4933 4093 4947 4107
rect 4913 4013 4927 4027
rect 4873 3973 4887 3987
rect 4893 3973 4907 3987
rect 4933 3953 4947 3967
rect 4913 3893 4927 3907
rect 4853 3873 4867 3887
rect 4853 3813 4867 3827
rect 4833 3453 4847 3467
rect 4813 3433 4827 3447
rect 4833 3413 4847 3427
rect 4813 3273 4827 3287
rect 4773 3213 4787 3227
rect 4793 3213 4807 3227
rect 4793 3193 4807 3207
rect 4673 3173 4687 3187
rect 4713 3093 4727 3107
rect 4713 3053 4727 3067
rect 4533 3013 4547 3027
rect 4613 3033 4627 3047
rect 4693 3033 4707 3047
rect 4633 3013 4647 3027
rect 4533 2713 4547 2727
rect 4553 2673 4567 2687
rect 4513 2653 4527 2667
rect 4613 2993 4627 3007
rect 4613 2813 4627 2827
rect 4593 2773 4607 2787
rect 4593 2733 4607 2747
rect 4573 2613 4587 2627
rect 4453 2493 4467 2507
rect 4453 2473 4467 2487
rect 4473 2433 4487 2447
rect 4513 2453 4527 2467
rect 4433 2313 4447 2327
rect 4473 2293 4487 2307
rect 4753 3033 4767 3047
rect 4773 3033 4787 3047
rect 4813 2993 4827 3007
rect 4793 2953 4807 2967
rect 4733 2933 4747 2947
rect 4693 2733 4707 2747
rect 4773 2733 4787 2747
rect 4633 2593 4647 2607
rect 4813 2673 4827 2687
rect 4833 2453 4847 2467
rect 4693 2393 4707 2407
rect 4613 2373 4627 2387
rect 4673 2353 4687 2367
rect 4553 2313 4567 2327
rect 4633 2313 4647 2327
rect 4593 2273 4607 2287
rect 4613 2253 4627 2267
rect 4593 2233 4607 2247
rect 4533 2193 4547 2207
rect 4373 2073 4387 2087
rect 4313 1913 4327 1927
rect 4213 1893 4227 1907
rect 4213 1853 4227 1867
rect 4273 1833 4287 1847
rect 4233 1793 4247 1807
rect 4253 1773 4267 1787
rect 4393 2053 4407 2067
rect 4513 2133 4527 2147
rect 4453 2093 4467 2107
rect 4513 2093 4527 2107
rect 4433 2053 4447 2067
rect 4413 1913 4427 1927
rect 4353 1833 4367 1847
rect 4333 1753 4347 1767
rect 4333 1733 4347 1747
rect 4233 1673 4247 1687
rect 4333 1693 4347 1707
rect 4573 2193 4587 2207
rect 4473 2073 4487 2087
rect 4493 2053 4507 2067
rect 4553 2073 4567 2087
rect 4533 2053 4547 2067
rect 4453 1833 4467 1847
rect 4493 1833 4507 1847
rect 4553 1833 4567 1847
rect 4173 1373 4187 1387
rect 4133 1353 4147 1367
rect 4053 1313 4067 1327
rect 4093 1313 4107 1327
rect 4013 1273 4027 1287
rect 4013 1133 4027 1147
rect 3973 1113 3987 1127
rect 3973 1093 3987 1107
rect 3913 1013 3927 1027
rect 3833 833 3847 847
rect 3813 653 3827 667
rect 3773 633 3787 647
rect 3793 613 3807 627
rect 3733 593 3747 607
rect 3813 513 3827 527
rect 3733 393 3747 407
rect 3793 393 3807 407
rect 3633 353 3647 367
rect 3713 333 3727 347
rect 3553 193 3567 207
rect 3553 173 3567 187
rect 3673 293 3687 307
rect 3733 173 3747 187
rect 3893 853 3907 867
rect 3853 753 3867 767
rect 3893 813 3907 827
rect 3913 833 3927 847
rect 3993 893 4007 907
rect 4093 1133 4107 1147
rect 4113 1113 4127 1127
rect 4053 1053 4067 1067
rect 4153 1313 4167 1327
rect 4193 1313 4207 1327
rect 4173 1273 4187 1287
rect 4213 1233 4227 1247
rect 4213 1193 4227 1207
rect 4153 1113 4167 1127
rect 4173 1113 4187 1127
rect 4013 833 4027 847
rect 4033 853 4047 867
rect 3893 713 3907 727
rect 3873 693 3887 707
rect 3933 653 3947 667
rect 3893 613 3907 627
rect 3913 633 3927 647
rect 4093 873 4107 887
rect 4133 873 4147 887
rect 3993 793 4007 807
rect 4053 793 4067 807
rect 4073 773 4087 787
rect 4033 693 4047 707
rect 3993 613 4007 627
rect 4053 613 4067 627
rect 4073 633 4087 647
rect 3913 533 3927 547
rect 3953 533 3967 547
rect 3853 413 3867 427
rect 3893 413 3907 427
rect 3833 393 3847 407
rect 3853 373 3867 387
rect 3833 333 3847 347
rect 3873 333 3887 347
rect 4013 513 4027 527
rect 4113 853 4127 867
rect 4153 853 4167 867
rect 4213 913 4227 927
rect 4173 833 4187 847
rect 4193 813 4207 827
rect 4133 793 4147 807
rect 4113 433 4127 447
rect 4293 1653 4307 1667
rect 4353 1653 4367 1667
rect 4253 1593 4267 1607
rect 4273 1573 4287 1587
rect 4333 1593 4347 1607
rect 4273 1473 4287 1487
rect 4313 1473 4327 1487
rect 4353 1393 4367 1407
rect 4293 1293 4307 1307
rect 4313 1313 4327 1327
rect 4273 1273 4287 1287
rect 4333 1273 4347 1287
rect 4453 1793 4467 1807
rect 4433 1773 4447 1787
rect 4473 1773 4487 1787
rect 4453 1693 4467 1707
rect 4453 1613 4467 1627
rect 4473 1613 4487 1627
rect 4433 1573 4447 1587
rect 4493 1593 4507 1607
rect 4473 1473 4487 1487
rect 4493 1333 4507 1347
rect 4453 1293 4467 1307
rect 4553 1773 4567 1787
rect 4533 1733 4547 1747
rect 4553 1713 4567 1727
rect 4553 1693 4567 1707
rect 4533 1613 4547 1627
rect 4633 2153 4647 2167
rect 4613 2033 4627 2047
rect 4633 2053 4647 2067
rect 4613 2013 4627 2027
rect 4593 1793 4607 1807
rect 4653 1993 4667 2007
rect 4733 2293 4747 2307
rect 4713 2253 4727 2267
rect 4713 2173 4727 2187
rect 4693 2093 4707 2107
rect 4673 1833 4687 1847
rect 4793 2393 4807 2407
rect 4773 2093 4787 2107
rect 4733 2033 4747 2047
rect 4753 2053 4767 2067
rect 4873 3673 4887 3687
rect 4893 3573 4907 3587
rect 4893 3473 4907 3487
rect 4913 3493 4927 3507
rect 4933 3353 4947 3367
rect 5053 4633 5067 4647
rect 5013 4613 5027 4627
rect 5073 4593 5087 4607
rect 4973 4473 4987 4487
rect 5113 4693 5127 4707
rect 5113 4653 5127 4667
rect 5313 5653 5327 5667
rect 5293 5613 5307 5627
rect 5313 5593 5327 5607
rect 5233 5553 5247 5567
rect 5253 5513 5267 5527
rect 5233 5473 5247 5487
rect 5293 5433 5307 5447
rect 5273 5413 5287 5427
rect 5233 5393 5247 5407
rect 5233 5373 5247 5387
rect 5213 5313 5227 5327
rect 5213 5153 5227 5167
rect 5293 5193 5307 5207
rect 5193 5113 5207 5127
rect 5193 5093 5207 5107
rect 5233 5073 5247 5087
rect 5213 4853 5227 4867
rect 5173 4833 5187 4847
rect 5233 4833 5247 4847
rect 5213 4733 5227 4747
rect 5193 4713 5207 4727
rect 5153 4693 5167 4707
rect 5173 4673 5187 4687
rect 5193 4633 5207 4647
rect 5133 4533 5147 4547
rect 5093 4513 5107 4527
rect 5013 4433 5027 4447
rect 4993 4413 5007 4427
rect 4993 4193 5007 4207
rect 4993 4133 5007 4147
rect 4973 3993 4987 4007
rect 4973 3493 4987 3507
rect 5053 4413 5067 4427
rect 5053 4153 5067 4167
rect 5013 3973 5027 3987
rect 5013 3753 5027 3767
rect 5033 3713 5047 3727
rect 5053 3733 5067 3747
rect 5153 4513 5167 4527
rect 5133 4453 5147 4467
rect 5133 4393 5147 4407
rect 5173 4493 5187 4507
rect 5213 4513 5227 4527
rect 5213 4473 5227 4487
rect 5293 4993 5307 5007
rect 5273 4733 5287 4747
rect 5373 5613 5387 5627
rect 5353 5593 5367 5607
rect 5353 5193 5367 5207
rect 5353 5153 5367 5167
rect 5333 5093 5347 5107
rect 5333 5053 5347 5067
rect 5253 4713 5267 4727
rect 5273 4713 5287 4727
rect 5313 4693 5327 4707
rect 5333 4693 5347 4707
rect 5313 4653 5327 4667
rect 5373 4773 5387 4787
rect 5373 4653 5387 4667
rect 5333 4633 5347 4647
rect 5353 4633 5367 4647
rect 5453 5693 5467 5707
rect 5593 5773 5607 5787
rect 5553 5753 5567 5767
rect 5633 5673 5647 5687
rect 5573 5653 5587 5667
rect 5633 5653 5647 5667
rect 5513 5613 5527 5627
rect 5433 5593 5447 5607
rect 5513 5593 5527 5607
rect 5413 5573 5427 5587
rect 5433 5473 5447 5487
rect 5473 5433 5487 5447
rect 5493 5433 5507 5447
rect 5453 5353 5467 5367
rect 5453 5153 5467 5167
rect 5473 5133 5487 5147
rect 5453 5113 5467 5127
rect 5473 5113 5487 5127
rect 5453 5053 5467 5067
rect 5453 4973 5467 4987
rect 5433 4913 5447 4927
rect 5433 4893 5447 4907
rect 5453 4773 5467 4787
rect 5413 4693 5427 4707
rect 5433 4673 5447 4687
rect 5453 4693 5467 4707
rect 5433 4653 5447 4667
rect 5313 4593 5327 4607
rect 5393 4593 5407 4607
rect 5153 4213 5167 4227
rect 5093 4193 5107 4207
rect 5193 4413 5207 4427
rect 5193 4393 5207 4407
rect 5193 4193 5207 4207
rect 5173 4153 5187 4167
rect 5113 4113 5127 4127
rect 5113 4093 5127 4107
rect 5153 4013 5167 4027
rect 5293 4553 5307 4567
rect 5293 4533 5307 4547
rect 5293 4513 5307 4527
rect 5293 4233 5307 4247
rect 5273 4213 5287 4227
rect 5253 4193 5267 4207
rect 5293 4193 5307 4207
rect 5353 4513 5367 4527
rect 5333 4493 5347 4507
rect 5213 4133 5227 4147
rect 5233 4093 5247 4107
rect 5273 4073 5287 4087
rect 5233 4053 5247 4067
rect 5293 4053 5307 4067
rect 5313 4053 5327 4067
rect 5193 4033 5207 4047
rect 5113 3973 5127 3987
rect 5133 3953 5147 3967
rect 5093 3933 5107 3947
rect 5073 3673 5087 3687
rect 5033 3553 5047 3567
rect 5013 3493 5027 3507
rect 5073 3513 5087 3527
rect 4993 3473 5007 3487
rect 5053 3453 5067 3467
rect 4973 3353 4987 3367
rect 4893 3273 4907 3287
rect 4953 3273 4967 3287
rect 4913 3233 4927 3247
rect 4933 3253 4947 3267
rect 4873 3213 4887 3227
rect 4933 3213 4947 3227
rect 4953 3213 4967 3227
rect 4973 3213 4987 3227
rect 5053 3233 5067 3247
rect 5073 3213 5087 3227
rect 4873 2993 4887 3007
rect 4893 3013 4907 3027
rect 4913 2973 4927 2987
rect 4913 2713 4927 2727
rect 4853 2353 4867 2367
rect 4853 2333 4867 2347
rect 4813 2273 4827 2287
rect 4833 2233 4847 2247
rect 4813 2093 4827 2107
rect 4713 2013 4727 2027
rect 4713 1873 4727 1887
rect 4713 1853 4727 1867
rect 4633 1773 4647 1787
rect 4613 1693 4627 1707
rect 4613 1613 4627 1627
rect 4573 1593 4587 1607
rect 4553 1573 4567 1587
rect 4633 1573 4647 1587
rect 4653 1593 4667 1607
rect 4533 1373 4547 1387
rect 4593 1533 4607 1547
rect 4753 2013 4767 2027
rect 4813 2013 4827 2027
rect 4733 1813 4747 1827
rect 4693 1753 4707 1767
rect 4653 1333 4667 1347
rect 4673 1333 4687 1347
rect 4553 1313 4567 1327
rect 4513 1293 4527 1307
rect 4573 1293 4587 1307
rect 4593 1313 4607 1327
rect 4633 1313 4647 1327
rect 4433 1253 4447 1267
rect 4473 1253 4487 1267
rect 4433 1213 4447 1227
rect 4413 1193 4427 1207
rect 4253 1173 4267 1187
rect 4373 1173 4387 1187
rect 4233 893 4247 907
rect 4353 1153 4367 1167
rect 4393 1153 4407 1167
rect 4353 1133 4367 1147
rect 4313 1113 4327 1127
rect 4333 1093 4347 1107
rect 4453 1133 4467 1147
rect 4573 1273 4587 1287
rect 4493 1153 4507 1167
rect 4533 1153 4547 1167
rect 4493 1113 4507 1127
rect 4453 1093 4467 1107
rect 4513 1093 4527 1107
rect 4413 1073 4427 1087
rect 4793 1873 4807 1887
rect 4793 1793 4807 1807
rect 4753 1753 4767 1767
rect 4813 1773 4827 1787
rect 4773 1733 4787 1747
rect 4773 1673 4787 1687
rect 4813 1693 4827 1707
rect 4793 1633 4807 1647
rect 4793 1613 4807 1627
rect 4753 1593 4767 1607
rect 4773 1593 4787 1607
rect 4733 1553 4747 1567
rect 4773 1513 4787 1527
rect 4733 1493 4747 1507
rect 4753 1413 4767 1427
rect 4713 1333 4727 1347
rect 4733 1313 4747 1327
rect 4893 2313 4907 2327
rect 4893 2293 4907 2307
rect 4873 2253 4887 2267
rect 5133 3913 5147 3927
rect 5133 3793 5147 3807
rect 5153 3753 5167 3767
rect 5153 3693 5167 3707
rect 5113 3673 5127 3687
rect 5213 3873 5227 3887
rect 5173 3573 5187 3587
rect 5133 3513 5147 3527
rect 5153 3513 5167 3527
rect 5153 3473 5167 3487
rect 5173 3493 5187 3507
rect 5113 3453 5127 3467
rect 5133 3453 5147 3467
rect 4993 3033 5007 3047
rect 5033 3033 5047 3047
rect 5013 2993 5027 3007
rect 4973 2973 4987 2987
rect 4953 2773 4967 2787
rect 4973 2753 4987 2767
rect 4953 2733 4967 2747
rect 4993 2733 5007 2747
rect 5013 2753 5027 2767
rect 5053 2753 5067 2767
rect 4933 2293 4947 2307
rect 4993 2713 5007 2727
rect 5053 2673 5067 2687
rect 4973 2433 4987 2447
rect 4913 2273 4927 2287
rect 5193 3453 5207 3467
rect 5153 3253 5167 3267
rect 5153 3233 5167 3247
rect 5113 3053 5127 3067
rect 5173 3053 5187 3067
rect 5133 3033 5147 3047
rect 5193 3013 5207 3027
rect 5113 2993 5127 3007
rect 5173 2973 5187 2987
rect 5133 2773 5147 2787
rect 5153 2753 5167 2767
rect 5173 2773 5187 2787
rect 5173 2733 5187 2747
rect 5133 2433 5147 2447
rect 5073 2333 5087 2347
rect 4973 2253 4987 2267
rect 5053 2273 5067 2287
rect 5093 2273 5107 2287
rect 5133 2273 5147 2287
rect 5113 2253 5127 2267
rect 4933 2233 4947 2247
rect 4893 2173 4907 2187
rect 4953 2133 4967 2147
rect 4873 2073 4887 2087
rect 4913 2073 4927 2087
rect 4853 2033 4867 2047
rect 4853 1833 4867 1847
rect 4833 1653 4847 1667
rect 4893 2053 4907 2067
rect 4933 2053 4947 2067
rect 5033 2193 5047 2207
rect 5033 2173 5047 2187
rect 4993 2153 5007 2167
rect 4893 1853 4907 1867
rect 4913 1793 4927 1807
rect 4933 1813 4947 1827
rect 4913 1733 4927 1747
rect 4853 1613 4867 1627
rect 4873 1613 4887 1627
rect 4893 1593 4907 1607
rect 4933 1613 4947 1627
rect 4833 1553 4847 1567
rect 4853 1553 4867 1567
rect 4813 1533 4827 1547
rect 4873 1513 4887 1527
rect 4813 1393 4827 1407
rect 4853 1393 4867 1407
rect 4853 1373 4867 1387
rect 4893 1313 4907 1327
rect 4693 1273 4707 1287
rect 4793 1273 4807 1287
rect 4793 1253 4807 1267
rect 4653 1173 4667 1187
rect 4693 1173 4707 1187
rect 4613 1133 4627 1147
rect 4653 1093 4667 1107
rect 4673 1093 4687 1107
rect 4593 873 4607 887
rect 4713 1153 4727 1167
rect 4713 1133 4727 1147
rect 4733 1133 4747 1147
rect 4713 1093 4727 1107
rect 4773 1113 4787 1127
rect 4893 1273 4907 1287
rect 4873 1193 4887 1207
rect 4813 1113 4827 1127
rect 4693 1073 4707 1087
rect 4753 1073 4767 1087
rect 4773 1073 4787 1087
rect 4813 1073 4827 1087
rect 4853 1073 4867 1087
rect 4613 853 4627 867
rect 4253 813 4267 827
rect 4313 833 4327 847
rect 4393 833 4407 847
rect 4433 833 4447 847
rect 4513 833 4527 847
rect 4293 793 4307 807
rect 4333 753 4347 767
rect 4353 673 4367 687
rect 4173 653 4187 667
rect 4213 653 4227 667
rect 4373 653 4387 667
rect 4193 613 4207 627
rect 4213 633 4227 647
rect 4233 613 4247 627
rect 4333 613 4347 627
rect 4213 593 4227 607
rect 4213 553 4227 567
rect 4193 433 4207 447
rect 3933 373 3947 387
rect 3913 353 3927 367
rect 3953 353 3967 367
rect 4013 353 4027 367
rect 3993 333 4007 347
rect 4013 253 4027 267
rect 3533 133 3547 147
rect 3673 113 3687 127
rect 3633 93 3647 107
rect 3853 153 3867 167
rect 4053 193 4067 207
rect 3993 113 4007 127
rect 4013 133 4027 147
rect 4153 393 4167 407
rect 4173 393 4187 407
rect 4093 373 4107 387
rect 4133 373 4147 387
rect 4113 353 4127 367
rect 4193 353 4207 367
rect 4213 333 4227 347
rect 4173 313 4187 327
rect 4253 333 4267 347
rect 4273 353 4287 367
rect 4233 293 4247 307
rect 4413 793 4427 807
rect 4533 813 4547 827
rect 4573 833 4587 847
rect 4553 793 4567 807
rect 4513 733 4527 747
rect 4433 693 4447 707
rect 4593 673 4607 687
rect 4473 653 4487 667
rect 4393 613 4407 627
rect 4793 873 4807 887
rect 4873 873 4887 887
rect 4653 853 4667 867
rect 4773 853 4787 867
rect 4693 833 4707 847
rect 4733 833 4747 847
rect 4673 733 4687 747
rect 4733 793 4747 807
rect 4773 793 4787 807
rect 4773 753 4787 767
rect 4713 673 4727 687
rect 4653 653 4667 667
rect 4453 613 4467 627
rect 4573 613 4587 627
rect 4613 613 4627 627
rect 4633 633 4647 647
rect 4813 793 4827 807
rect 4853 773 4867 787
rect 4853 693 4867 707
rect 4833 673 4847 687
rect 4793 653 4807 667
rect 4713 633 4727 647
rect 4733 633 4747 647
rect 4653 613 4667 627
rect 4753 613 4767 627
rect 4773 633 4787 647
rect 4913 1133 4927 1147
rect 4913 1073 4927 1087
rect 4893 853 4907 867
rect 4893 833 4907 847
rect 4973 1833 4987 1847
rect 5053 2133 5067 2147
rect 5013 2113 5027 2127
rect 5133 2233 5147 2247
rect 5073 2113 5087 2127
rect 5093 2113 5107 2127
rect 5113 2113 5127 2127
rect 5013 2073 5027 2087
rect 5073 2033 5087 2047
rect 5013 2013 5027 2027
rect 5073 1913 5087 1927
rect 5033 1833 5047 1847
rect 4993 1813 5007 1827
rect 4973 1793 4987 1807
rect 5013 1773 5027 1787
rect 5053 1773 5067 1787
rect 4993 1753 5007 1767
rect 5053 1753 5067 1767
rect 5093 1753 5107 1767
rect 5013 1673 5027 1687
rect 5013 1613 5027 1627
rect 5033 1533 5047 1547
rect 4993 1513 5007 1527
rect 5033 1453 5047 1467
rect 5013 1293 5027 1307
rect 5013 1273 5027 1287
rect 4993 1233 5007 1247
rect 4973 1133 4987 1147
rect 4993 1133 5007 1147
rect 4953 1073 4967 1087
rect 5013 1053 5027 1067
rect 5013 953 5027 967
rect 4933 873 4947 887
rect 4933 833 4947 847
rect 4953 813 4967 827
rect 4973 833 4987 847
rect 5073 1653 5087 1667
rect 5153 2113 5167 2127
rect 5253 4033 5267 4047
rect 5393 4473 5407 4487
rect 5353 4433 5367 4447
rect 5373 4413 5387 4427
rect 5413 4413 5427 4427
rect 5393 4193 5407 4207
rect 5373 4153 5387 4167
rect 5393 4153 5407 4167
rect 5373 4133 5387 4147
rect 5353 4113 5367 4127
rect 5293 3993 5307 4007
rect 5333 3993 5347 4007
rect 5253 3793 5267 3807
rect 5233 3733 5247 3747
rect 5453 4633 5467 4647
rect 5433 4153 5447 4167
rect 5513 5113 5527 5127
rect 5493 5093 5507 5107
rect 5573 5613 5587 5627
rect 5673 5633 5687 5647
rect 5653 5573 5667 5587
rect 5673 5533 5687 5547
rect 5613 5413 5627 5427
rect 5633 5393 5647 5407
rect 5573 5353 5587 5367
rect 5593 5353 5607 5367
rect 5633 5353 5647 5367
rect 5593 5313 5607 5327
rect 5573 5193 5587 5207
rect 5633 5173 5647 5187
rect 5513 4933 5527 4947
rect 5573 4953 5587 4967
rect 5573 4933 5587 4947
rect 5493 4873 5507 4887
rect 5613 4933 5627 4947
rect 5633 4913 5647 4927
rect 5573 4733 5587 4747
rect 5613 4793 5627 4807
rect 5613 4733 5627 4747
rect 5673 5393 5687 5407
rect 5713 5633 5727 5647
rect 5793 5693 5807 5707
rect 5733 5533 5747 5547
rect 5733 5433 5747 5447
rect 5673 5193 5687 5207
rect 5753 5373 5767 5387
rect 5713 5193 5727 5207
rect 5733 5193 5747 5207
rect 5713 5153 5727 5167
rect 5693 5133 5707 5147
rect 5713 5133 5727 5147
rect 5753 5133 5767 5147
rect 5673 4913 5687 4927
rect 5553 4673 5567 4687
rect 5573 4653 5587 4667
rect 5593 4653 5607 4667
rect 5513 4613 5527 4627
rect 5493 4513 5507 4527
rect 5493 4493 5507 4507
rect 5473 4433 5487 4447
rect 5593 4513 5607 4527
rect 5573 4413 5587 4427
rect 5533 4393 5547 4407
rect 5553 4293 5567 4307
rect 5473 4173 5487 4187
rect 5493 4193 5507 4207
rect 5573 4173 5587 4187
rect 5473 4113 5487 4127
rect 5453 4073 5467 4087
rect 5413 4033 5427 4047
rect 5413 4013 5427 4027
rect 5413 3973 5427 3987
rect 5393 3873 5407 3887
rect 5433 3813 5447 3827
rect 5233 3713 5247 3727
rect 5293 3713 5307 3727
rect 5353 3613 5367 3627
rect 5233 3573 5247 3587
rect 5313 3553 5327 3567
rect 5333 3533 5347 3547
rect 5373 3533 5387 3547
rect 5293 3513 5307 3527
rect 5253 3273 5267 3287
rect 5293 3253 5307 3267
rect 5273 3193 5287 3207
rect 5233 3133 5247 3147
rect 5253 3033 5267 3047
rect 5373 3473 5387 3487
rect 5373 3233 5387 3247
rect 5353 3053 5367 3067
rect 5213 2693 5227 2707
rect 5193 2673 5207 2687
rect 5233 2533 5247 2547
rect 5193 2473 5207 2487
rect 5313 2753 5327 2767
rect 5313 2733 5327 2747
rect 5353 2733 5367 2747
rect 5273 2353 5287 2367
rect 5353 2693 5367 2707
rect 5313 2333 5327 2347
rect 5233 2293 5247 2307
rect 5273 2293 5287 2307
rect 5213 2253 5227 2267
rect 5213 2193 5227 2207
rect 5153 2093 5167 2107
rect 5173 2093 5187 2107
rect 5193 2093 5207 2107
rect 5153 2053 5167 2067
rect 5173 2053 5187 2067
rect 5133 1793 5147 1807
rect 5133 1773 5147 1787
rect 5073 1553 5087 1567
rect 5073 1453 5087 1467
rect 5113 1633 5127 1647
rect 5113 1513 5127 1527
rect 5093 1413 5107 1427
rect 5193 2033 5207 2047
rect 5173 1793 5187 1807
rect 5173 1713 5187 1727
rect 5193 1673 5207 1687
rect 5193 1653 5207 1667
rect 5233 2113 5247 2127
rect 5273 2093 5287 2107
rect 5253 2073 5267 2087
rect 5313 2053 5327 2067
rect 5233 2013 5247 2027
rect 5253 1913 5267 1927
rect 5293 1893 5307 1907
rect 5253 1853 5267 1867
rect 5233 1733 5247 1747
rect 5233 1713 5247 1727
rect 5173 1553 5187 1567
rect 5193 1533 5207 1547
rect 5133 1373 5147 1387
rect 5133 1353 5147 1367
rect 5093 1333 5107 1347
rect 5113 1313 5127 1327
rect 5133 1173 5147 1187
rect 5053 953 5067 967
rect 5033 893 5047 907
rect 5133 893 5147 907
rect 5073 833 5087 847
rect 5033 813 5047 827
rect 5073 793 5087 807
rect 5113 793 5127 807
rect 4913 773 4927 787
rect 5113 773 5127 787
rect 4993 673 5007 687
rect 4873 653 4887 667
rect 4913 653 4927 667
rect 4953 653 4967 667
rect 5093 653 5107 667
rect 4853 633 4867 647
rect 4793 613 4807 627
rect 4833 613 4847 627
rect 4873 613 4887 627
rect 4893 633 4907 647
rect 4813 593 4827 607
rect 4793 493 4807 507
rect 4493 453 4507 467
rect 4533 453 4547 467
rect 4513 393 4527 407
rect 4413 373 4427 387
rect 4373 353 4387 367
rect 4313 313 4327 327
rect 4173 273 4187 287
rect 4133 193 4147 207
rect 4073 153 4087 167
rect 4093 153 4107 167
rect 4113 153 4127 167
rect 4093 113 4107 127
rect 4413 293 4427 307
rect 4333 193 4347 207
rect 4293 153 4307 167
rect 4493 353 4507 367
rect 4513 373 4527 387
rect 4533 353 4547 367
rect 4573 353 4587 367
rect 4593 333 4607 347
rect 4633 353 4647 367
rect 4673 353 4687 367
rect 4733 353 4747 367
rect 4613 313 4627 327
rect 4753 313 4767 327
rect 4573 273 4587 287
rect 4453 253 4467 267
rect 4633 233 4647 247
rect 4593 213 4607 227
rect 4393 113 4407 127
rect 4453 133 4467 147
rect 4513 113 4527 127
rect 4553 133 4567 147
rect 4613 133 4627 147
rect 4573 113 4587 127
rect 4533 93 4547 107
rect 4693 213 4707 227
rect 4753 173 4767 187
rect 4713 153 4727 167
rect 4813 373 4827 387
rect 5173 1433 5187 1447
rect 5153 673 5167 687
rect 5133 653 5147 667
rect 5153 653 5167 667
rect 5133 633 5147 647
rect 5093 473 5107 487
rect 5153 433 5167 447
rect 5133 413 5147 427
rect 5073 393 5087 407
rect 5013 373 5027 387
rect 4893 333 4907 347
rect 4953 353 4967 367
rect 4813 313 4827 327
rect 4973 313 4987 327
rect 4853 233 4867 247
rect 4953 213 4967 227
rect 4873 153 4887 167
rect 4833 133 4847 147
rect 5033 333 5047 347
rect 4993 193 5007 207
rect 5213 1513 5227 1527
rect 5373 2533 5387 2547
rect 5373 2313 5387 2327
rect 5353 2193 5367 2207
rect 5433 3713 5447 3727
rect 5453 3613 5467 3627
rect 5433 3433 5447 3447
rect 5433 3373 5447 3387
rect 5493 4073 5507 4087
rect 5533 4153 5547 4167
rect 5513 4053 5527 4067
rect 5513 4033 5527 4047
rect 5513 3993 5527 4007
rect 5493 3973 5507 3987
rect 5493 3733 5507 3747
rect 5513 3693 5527 3707
rect 5553 3993 5567 4007
rect 5553 3653 5567 3667
rect 5613 4293 5627 4307
rect 5613 3773 5627 3787
rect 5613 3733 5627 3747
rect 5533 3513 5547 3527
rect 5573 3513 5587 3527
rect 5593 3513 5607 3527
rect 5513 3493 5527 3507
rect 5493 3473 5507 3487
rect 5473 3373 5487 3387
rect 5533 3473 5547 3487
rect 5553 3493 5567 3507
rect 5593 3453 5607 3467
rect 5573 3433 5587 3447
rect 5513 3273 5527 3287
rect 5553 3273 5567 3287
rect 5473 3213 5487 3227
rect 5493 3233 5507 3247
rect 5533 3053 5547 3067
rect 5513 3033 5527 3047
rect 5453 2913 5467 2927
rect 5493 2913 5507 2927
rect 5433 2833 5447 2847
rect 5433 2673 5447 2687
rect 5493 2833 5507 2847
rect 5473 2733 5487 2747
rect 5453 2533 5467 2547
rect 5413 2413 5427 2427
rect 5413 2373 5427 2387
rect 5453 2293 5467 2307
rect 5393 2253 5407 2267
rect 5393 2233 5407 2247
rect 5373 2093 5387 2107
rect 5353 2073 5367 2087
rect 5453 2253 5467 2267
rect 5433 2113 5447 2127
rect 5433 2093 5447 2107
rect 5333 1853 5347 1867
rect 5353 1853 5367 1867
rect 5333 1833 5347 1847
rect 5293 1793 5307 1807
rect 5273 1773 5287 1787
rect 5313 1753 5327 1767
rect 5413 2013 5427 2027
rect 5393 1853 5407 1867
rect 5433 1833 5447 1847
rect 5373 1773 5387 1787
rect 5413 1773 5427 1787
rect 5353 1753 5367 1767
rect 5413 1753 5427 1767
rect 5373 1713 5387 1727
rect 5393 1713 5407 1727
rect 5273 1673 5287 1687
rect 5333 1673 5347 1687
rect 5253 1653 5267 1667
rect 5293 1653 5307 1667
rect 5373 1633 5387 1647
rect 5273 1593 5287 1607
rect 5253 1533 5267 1547
rect 5233 1433 5247 1447
rect 5233 1413 5247 1427
rect 5213 1373 5227 1387
rect 5253 1353 5267 1367
rect 5313 1573 5327 1587
rect 5333 1593 5347 1607
rect 5353 1573 5367 1587
rect 5333 1553 5347 1567
rect 5313 1513 5327 1527
rect 5253 1313 5267 1327
rect 5273 1333 5287 1347
rect 5213 1273 5227 1287
rect 5393 1533 5407 1547
rect 5433 1733 5447 1747
rect 5533 2733 5547 2747
rect 5533 2693 5547 2707
rect 5493 2533 5507 2547
rect 5493 2373 5507 2387
rect 5573 2913 5587 2927
rect 5753 5093 5767 5107
rect 5753 4973 5767 4987
rect 5733 4913 5747 4927
rect 5713 4893 5727 4907
rect 5773 4893 5787 4907
rect 5773 4793 5787 4807
rect 5673 4713 5687 4727
rect 5693 4713 5707 4727
rect 5753 4713 5767 4727
rect 5693 4653 5707 4667
rect 5733 4653 5747 4667
rect 5773 4653 5787 4667
rect 5713 4613 5727 4627
rect 5673 4473 5687 4487
rect 5673 4433 5687 4447
rect 5673 4213 5687 4227
rect 5673 4193 5687 4207
rect 5653 4173 5667 4187
rect 5653 4153 5667 4167
rect 5733 4413 5747 4427
rect 5713 4133 5727 4147
rect 5773 4173 5787 4187
rect 5773 4133 5787 4147
rect 5693 4033 5707 4047
rect 5653 3933 5667 3947
rect 5733 3993 5747 4007
rect 5753 3973 5767 3987
rect 5713 3953 5727 3967
rect 5733 3953 5747 3967
rect 5673 3913 5687 3927
rect 5713 3913 5727 3927
rect 5693 3773 5707 3787
rect 5673 3653 5687 3667
rect 5633 3533 5647 3547
rect 5633 3513 5647 3527
rect 5653 3493 5667 3507
rect 5753 3933 5767 3947
rect 5713 3753 5727 3767
rect 5733 3753 5747 3767
rect 5733 3713 5747 3727
rect 5753 3733 5767 3747
rect 5713 3693 5727 3707
rect 5733 3493 5747 3507
rect 5713 3453 5727 3467
rect 5653 3433 5667 3447
rect 5613 3253 5627 3267
rect 5693 3253 5707 3267
rect 5633 3213 5647 3227
rect 5613 3013 5627 3027
rect 5673 3033 5687 3047
rect 5633 2753 5647 2767
rect 5733 2913 5747 2927
rect 5673 2733 5687 2747
rect 5613 2713 5627 2727
rect 5653 2693 5667 2707
rect 5613 2673 5627 2687
rect 5593 2533 5607 2547
rect 5553 2313 5567 2327
rect 5513 2293 5527 2307
rect 5553 2273 5567 2287
rect 5573 2273 5587 2287
rect 5513 2233 5527 2247
rect 5533 2153 5547 2167
rect 5533 2133 5547 2147
rect 5473 2033 5487 2047
rect 5473 2013 5487 2027
rect 5453 1713 5467 1727
rect 5433 1693 5447 1707
rect 5513 2053 5527 2067
rect 5513 2033 5527 2047
rect 5493 1873 5507 1887
rect 5493 1793 5507 1807
rect 5473 1653 5487 1667
rect 5473 1593 5487 1607
rect 5433 1553 5447 1567
rect 5453 1553 5467 1567
rect 5493 1553 5507 1567
rect 5453 1533 5467 1547
rect 5413 1493 5427 1507
rect 5433 1473 5447 1487
rect 5333 1453 5347 1467
rect 5313 1333 5327 1347
rect 5293 1253 5307 1267
rect 5393 1333 5407 1347
rect 5353 1313 5367 1327
rect 5413 1253 5427 1267
rect 5333 1153 5347 1167
rect 5373 1153 5387 1167
rect 5233 1133 5247 1147
rect 5293 1133 5307 1147
rect 5313 1133 5327 1147
rect 5273 1113 5287 1127
rect 5233 873 5247 887
rect 5213 673 5227 687
rect 5213 513 5227 527
rect 5153 373 5167 387
rect 5173 373 5187 387
rect 5133 353 5147 367
rect 5153 333 5167 347
rect 5173 353 5187 367
rect 5193 333 5207 347
rect 5133 313 5147 327
rect 5193 233 5207 247
rect 5093 193 5107 207
rect 5033 173 5047 187
rect 5073 173 5087 187
rect 4973 153 4987 167
rect 4993 133 5007 147
rect 5013 153 5027 167
rect 5033 133 5047 147
rect 5113 153 5127 167
rect 5253 813 5267 827
rect 5253 793 5267 807
rect 5273 793 5287 807
rect 5253 733 5267 747
rect 5413 1133 5427 1147
rect 5373 1113 5387 1127
rect 5313 873 5327 887
rect 5313 833 5327 847
rect 5313 813 5327 827
rect 5293 773 5307 787
rect 5273 673 5287 687
rect 5393 1093 5407 1107
rect 5413 893 5427 907
rect 5373 833 5387 847
rect 5413 813 5427 827
rect 5333 793 5347 807
rect 5393 793 5407 807
rect 5433 733 5447 747
rect 5333 713 5347 727
rect 5273 633 5287 647
rect 5253 613 5267 627
rect 5353 693 5367 707
rect 5373 693 5387 707
rect 5433 693 5447 707
rect 5293 593 5307 607
rect 5333 593 5347 607
rect 5393 613 5407 627
rect 5413 633 5427 647
rect 5633 2333 5647 2347
rect 5653 2253 5667 2267
rect 5633 2233 5647 2247
rect 5713 2533 5727 2547
rect 5713 2293 5727 2307
rect 5693 2273 5707 2287
rect 5733 2273 5747 2287
rect 5633 2053 5647 2067
rect 5533 1793 5547 1807
rect 5533 1773 5547 1787
rect 5533 1593 5547 1607
rect 5513 1473 5527 1487
rect 5593 1753 5607 1767
rect 5573 1733 5587 1747
rect 5573 1633 5587 1647
rect 5713 2233 5727 2247
rect 5673 2193 5687 2207
rect 5733 2193 5747 2207
rect 5733 2173 5747 2187
rect 5753 2133 5767 2147
rect 5673 2093 5687 2107
rect 5733 2093 5747 2107
rect 5713 2053 5727 2067
rect 5733 2073 5747 2087
rect 5673 2033 5687 2047
rect 5693 2033 5707 2047
rect 5653 1793 5667 1807
rect 5633 1613 5647 1627
rect 5653 1593 5667 1607
rect 5573 1573 5587 1587
rect 5553 1553 5567 1567
rect 5613 1573 5627 1587
rect 5593 1553 5607 1567
rect 5613 1533 5627 1547
rect 5573 1393 5587 1407
rect 5533 1373 5547 1387
rect 5553 1353 5567 1367
rect 5493 1333 5507 1347
rect 5493 1313 5507 1327
rect 5473 1173 5487 1187
rect 5473 1133 5487 1147
rect 5493 1133 5507 1147
rect 5533 1133 5547 1147
rect 5513 1113 5527 1127
rect 5593 1333 5607 1347
rect 5593 1193 5607 1207
rect 5593 1173 5607 1187
rect 5573 1073 5587 1087
rect 5493 913 5507 927
rect 5533 913 5547 927
rect 5533 873 5547 887
rect 5473 813 5487 827
rect 5493 833 5507 847
rect 5573 833 5587 847
rect 5733 2033 5747 2047
rect 5773 2033 5787 2047
rect 5713 2013 5727 2027
rect 5693 1973 5707 1987
rect 5673 1533 5687 1547
rect 5653 1393 5667 1407
rect 5653 1373 5667 1387
rect 5633 1333 5647 1347
rect 5713 1613 5727 1627
rect 5693 1353 5707 1367
rect 5633 1273 5647 1287
rect 5633 1193 5647 1207
rect 5613 1113 5627 1127
rect 5673 1173 5687 1187
rect 5673 1153 5687 1167
rect 5713 1133 5727 1147
rect 5673 1093 5687 1107
rect 5693 1093 5707 1107
rect 5713 1093 5727 1107
rect 5653 1073 5667 1087
rect 5613 893 5627 907
rect 5693 873 5707 887
rect 5613 853 5627 867
rect 5653 853 5667 867
rect 5553 813 5567 827
rect 5593 813 5607 827
rect 5493 773 5507 787
rect 5473 733 5487 747
rect 5453 653 5467 667
rect 5473 613 5487 627
rect 5493 533 5507 547
rect 5393 513 5407 527
rect 5253 453 5267 467
rect 5353 453 5367 467
rect 5233 353 5247 367
rect 5213 193 5227 207
rect 5353 413 5367 427
rect 5293 393 5307 407
rect 5333 353 5347 367
rect 5373 393 5387 407
rect 5373 333 5387 347
rect 5353 233 5367 247
rect 5313 213 5327 227
rect 5333 193 5347 207
rect 5593 693 5607 707
rect 5553 673 5567 687
rect 5533 633 5547 647
rect 5573 613 5587 627
rect 5593 633 5607 647
rect 5513 493 5527 507
rect 5413 473 5427 487
rect 5593 473 5607 487
rect 5513 393 5527 407
rect 5553 393 5567 407
rect 5433 373 5447 387
rect 5413 313 5427 327
rect 5233 153 5247 167
rect 5293 153 5307 167
rect 5233 133 5247 147
rect 5353 133 5367 147
rect 5473 353 5487 367
rect 5693 833 5707 847
rect 5673 813 5687 827
rect 5653 733 5667 747
rect 5633 653 5647 667
rect 5613 433 5627 447
rect 5673 713 5687 727
rect 5693 633 5707 647
rect 5653 593 5667 607
rect 5753 1633 5767 1647
rect 5813 5673 5827 5687
rect 5813 3933 5827 3947
rect 5813 3813 5827 3827
rect 5813 2133 5827 2147
rect 5793 1593 5807 1607
rect 5793 1573 5807 1587
rect 5773 1513 5787 1527
rect 5773 1493 5787 1507
rect 5753 1353 5767 1367
rect 5753 1153 5767 1167
rect 5753 1093 5767 1107
rect 5773 1093 5787 1107
rect 5753 873 5767 887
rect 5633 393 5647 407
rect 5613 373 5627 387
rect 5633 353 5647 367
rect 5613 333 5627 347
rect 5493 313 5507 327
rect 5453 173 5467 187
rect 5613 173 5627 187
rect 5493 133 5507 147
rect 5673 533 5687 547
rect 5673 173 5687 187
rect 5733 593 5747 607
rect 5713 393 5727 407
rect 5753 393 5767 407
rect 5733 353 5747 367
rect 5793 353 5807 367
rect 5733 173 5747 187
rect 5593 133 5607 147
rect 5653 133 5667 147
rect 5253 113 5267 127
rect 5373 113 5387 127
rect 5433 113 5447 127
rect 5673 113 5687 127
rect 4633 93 4647 107
<< metal3 >>
rect 5087 5776 5233 5784
rect 5407 5776 5593 5784
rect 5167 5756 5553 5764
rect 5467 5696 5793 5704
rect 4847 5676 4973 5684
rect 5147 5676 5173 5684
rect 5187 5676 5633 5684
rect 5827 5676 5864 5684
rect 467 5656 513 5664
rect 847 5656 1333 5664
rect 1507 5656 1633 5664
rect 1947 5656 2073 5664
rect 2087 5656 2113 5664
rect 2387 5656 2453 5664
rect 2627 5656 2713 5664
rect 2767 5656 2793 5664
rect 2807 5656 2873 5664
rect 2887 5656 3253 5664
rect 3267 5656 3433 5664
rect 3447 5656 3493 5664
rect 3547 5656 4093 5664
rect 4456 5656 4584 5664
rect 4456 5647 4464 5656
rect 127 5636 213 5644
rect 227 5636 244 5644
rect 147 5616 193 5624
rect 236 5624 244 5636
rect 407 5636 533 5644
rect 707 5636 733 5644
rect 907 5636 933 5644
rect 1527 5636 1673 5644
rect 1687 5636 1753 5644
rect 2047 5636 2133 5644
rect 2147 5636 2173 5644
rect 2347 5636 2413 5644
rect 2487 5636 2593 5644
rect 2647 5636 2693 5644
rect 2987 5636 3073 5644
rect 3527 5636 3653 5644
rect 3867 5636 3953 5644
rect 4507 5636 4553 5644
rect 4576 5644 4584 5656
rect 4727 5656 4733 5664
rect 4747 5656 4873 5664
rect 4907 5656 5313 5664
rect 5587 5656 5633 5664
rect 5647 5656 5864 5664
rect 4576 5636 5193 5644
rect 5687 5636 5713 5644
rect 5856 5636 5864 5656
rect 236 5616 373 5624
rect 1216 5624 1224 5633
rect 787 5616 1224 5624
rect 1267 5616 1373 5624
rect 1387 5616 1393 5624
rect 1567 5616 1733 5624
rect 1887 5616 2213 5624
rect 3116 5624 3124 5633
rect 3116 5616 3233 5624
rect 3307 5616 3373 5624
rect 3387 5616 3493 5624
rect 4287 5616 4473 5624
rect 5007 5616 5053 5624
rect 5147 5616 5213 5624
rect 5307 5616 5373 5624
rect 5527 5616 5573 5624
rect 427 5596 493 5604
rect 547 5596 913 5604
rect 1007 5596 1073 5604
rect 1287 5596 1413 5604
rect 1547 5596 1693 5604
rect 1707 5596 1773 5604
rect 1787 5596 1833 5604
rect 1867 5596 1913 5604
rect 2127 5596 2153 5604
rect 2207 5596 2733 5604
rect 3147 5596 3393 5604
rect 3687 5596 3933 5604
rect 4007 5596 4073 5604
rect 4247 5596 4573 5604
rect 4827 5596 4853 5604
rect 4947 5596 5093 5604
rect 5327 5596 5353 5604
rect 5447 5596 5513 5604
rect 727 5576 893 5584
rect 907 5576 1093 5584
rect 1127 5576 1353 5584
rect 1927 5576 2313 5584
rect 3627 5576 3773 5584
rect 3787 5576 4133 5584
rect 5427 5576 5653 5584
rect 667 5556 793 5564
rect 807 5556 813 5564
rect 1827 5556 2273 5564
rect 2287 5556 2313 5564
rect 2787 5556 2813 5564
rect 2827 5556 3973 5564
rect 4527 5556 5233 5564
rect 267 5536 653 5544
rect 667 5536 1053 5544
rect 1067 5536 1393 5544
rect 2387 5536 2773 5544
rect 2787 5536 2873 5544
rect 3007 5536 3713 5544
rect 3747 5536 3973 5544
rect 5687 5536 5733 5544
rect 3407 5516 3793 5524
rect 3967 5516 4533 5524
rect 4587 5516 4913 5524
rect 4927 5516 5033 5524
rect 5047 5516 5253 5524
rect 1387 5496 3753 5504
rect 3787 5496 3853 5504
rect 3867 5496 3953 5504
rect 3987 5496 4553 5504
rect 4567 5496 4713 5504
rect 107 5476 393 5484
rect 547 5476 573 5484
rect 587 5476 693 5484
rect 1627 5476 1633 5484
rect 1647 5476 1693 5484
rect 1987 5476 2553 5484
rect 2567 5476 2933 5484
rect 3547 5476 3913 5484
rect 4447 5476 5093 5484
rect 5107 5476 5133 5484
rect 5247 5476 5433 5484
rect 87 5456 133 5464
rect 147 5456 573 5464
rect 587 5456 773 5464
rect 1147 5456 1173 5464
rect 1747 5456 1853 5464
rect 1867 5456 2053 5464
rect 2107 5456 2233 5464
rect 2247 5456 2413 5464
rect 2507 5456 2513 5464
rect 2527 5456 2853 5464
rect 2927 5456 3013 5464
rect 3027 5456 3253 5464
rect 3567 5456 3833 5464
rect 3847 5456 4313 5464
rect 4387 5456 4493 5464
rect 4507 5456 4753 5464
rect 287 5436 524 5444
rect 96 5407 104 5433
rect 127 5416 193 5424
rect 447 5416 493 5424
rect 516 5407 524 5436
rect 627 5436 833 5444
rect 967 5436 1293 5444
rect 1367 5436 1413 5444
rect 1516 5436 1553 5444
rect 607 5416 673 5424
rect 747 5416 813 5424
rect 867 5416 913 5424
rect 927 5416 933 5424
rect 987 5416 1073 5424
rect 1167 5416 1253 5424
rect 367 5396 413 5404
rect 536 5396 553 5404
rect 67 5376 73 5384
rect 536 5384 544 5396
rect 567 5396 673 5404
rect 1187 5396 1233 5404
rect 87 5376 544 5384
rect 1167 5376 1253 5384
rect 1516 5384 1524 5436
rect 1607 5436 1633 5444
rect 1656 5427 1664 5453
rect 1687 5436 1953 5444
rect 2487 5436 2553 5444
rect 2607 5436 2673 5444
rect 3107 5436 3273 5444
rect 3287 5436 3373 5444
rect 3447 5436 3533 5444
rect 3607 5436 3733 5444
rect 3827 5436 3864 5444
rect 3856 5427 3864 5436
rect 3907 5436 4093 5444
rect 4167 5436 4593 5444
rect 5147 5436 5173 5444
rect 5307 5436 5473 5444
rect 5507 5436 5733 5444
rect 1787 5416 1813 5424
rect 2047 5416 2073 5424
rect 2647 5416 2684 5424
rect 1536 5404 1544 5413
rect 1536 5396 1793 5404
rect 1987 5396 2053 5404
rect 2107 5396 2613 5404
rect 2676 5404 2684 5416
rect 2867 5416 2893 5424
rect 3147 5416 3173 5424
rect 3347 5416 3413 5424
rect 3587 5416 3693 5424
rect 3727 5416 3733 5424
rect 3807 5416 3833 5424
rect 4127 5416 4233 5424
rect 4367 5416 4473 5424
rect 4527 5416 4633 5424
rect 5287 5416 5613 5424
rect 2676 5396 2753 5404
rect 3047 5396 3113 5404
rect 3296 5404 3304 5413
rect 3296 5396 3433 5404
rect 3447 5396 3673 5404
rect 3736 5404 3744 5413
rect 3736 5396 3873 5404
rect 3907 5396 4153 5404
rect 4267 5396 4373 5404
rect 4427 5396 4513 5404
rect 4567 5396 4733 5404
rect 5167 5396 5233 5404
rect 5647 5396 5673 5404
rect 1516 5376 1533 5384
rect 2027 5376 2093 5384
rect 2656 5384 2664 5393
rect 2567 5376 2664 5384
rect 3167 5376 3333 5384
rect 3716 5384 3724 5393
rect 3716 5376 3773 5384
rect 4007 5376 4133 5384
rect 5247 5376 5753 5384
rect 427 5356 453 5364
rect 507 5356 713 5364
rect 4067 5356 4073 5364
rect 4087 5356 4213 5364
rect 4227 5356 4473 5364
rect 4807 5356 5113 5364
rect 5127 5356 5453 5364
rect 5587 5356 5593 5364
rect 5607 5356 5633 5364
rect 407 5336 473 5344
rect 4287 5336 4833 5344
rect 4887 5336 5173 5344
rect 67 5316 93 5324
rect 5227 5316 5593 5324
rect 2187 5296 2333 5304
rect 1567 5276 1593 5284
rect 3507 5256 3973 5264
rect 3987 5256 4673 5264
rect 187 5236 233 5244
rect 167 5216 233 5224
rect 247 5216 613 5224
rect 2027 5216 2193 5224
rect 3567 5216 4413 5224
rect 547 5196 993 5204
rect 2007 5196 2033 5204
rect 2107 5196 2213 5204
rect 2227 5196 2393 5204
rect 2407 5196 2553 5204
rect 3647 5196 3973 5204
rect 3996 5196 4573 5204
rect 96 5176 153 5184
rect 96 5167 104 5176
rect 207 5176 273 5184
rect 327 5176 453 5184
rect 507 5176 613 5184
rect 807 5176 1013 5184
rect 896 5167 904 5176
rect 1067 5176 1293 5184
rect 1707 5176 1893 5184
rect 1927 5176 2053 5184
rect 2067 5176 2313 5184
rect 2367 5176 2473 5184
rect 2827 5176 3553 5184
rect 3707 5176 3773 5184
rect 3996 5184 4004 5196
rect 5307 5196 5353 5204
rect 5587 5196 5673 5204
rect 5696 5196 5713 5204
rect 3927 5176 4004 5184
rect 4056 5176 4253 5184
rect 127 5156 193 5164
rect 367 5156 433 5164
rect 487 5156 573 5164
rect 767 5156 873 5164
rect 1087 5156 1153 5164
rect 1367 5156 1413 5164
rect 1467 5156 1513 5164
rect 1667 5156 1753 5164
rect 1807 5156 1833 5164
rect 2147 5156 2193 5164
rect 2287 5156 2333 5164
rect 2347 5156 2513 5164
rect 2747 5156 2893 5164
rect 3807 5156 3893 5164
rect 4036 5164 4044 5173
rect 4056 5167 4064 5176
rect 5087 5176 5633 5184
rect 4007 5156 4044 5164
rect 4227 5156 4293 5164
rect 4307 5156 4333 5164
rect 4487 5156 4633 5164
rect 4647 5156 4693 5164
rect 4856 5156 5213 5164
rect 427 5136 513 5144
rect 747 5136 813 5144
rect 867 5136 913 5144
rect 1347 5136 1433 5144
rect 1547 5136 1673 5144
rect 1727 5136 1753 5144
rect 1767 5136 1933 5144
rect 1947 5136 2073 5144
rect 2427 5136 2453 5144
rect 2567 5136 2873 5144
rect 2896 5144 2904 5153
rect 2896 5136 2993 5144
rect 3047 5136 3113 5144
rect 3127 5136 3653 5144
rect 3296 5127 3304 5136
rect 4016 5136 4193 5144
rect 4016 5127 4024 5136
rect 4267 5136 4353 5144
rect 4387 5136 4533 5144
rect 4547 5136 4593 5144
rect 4736 5144 4744 5153
rect 4667 5136 4744 5144
rect 4856 5144 4864 5156
rect 5236 5156 5353 5164
rect 4847 5136 4864 5144
rect 5236 5144 5244 5156
rect 5367 5156 5453 5164
rect 5696 5147 5704 5196
rect 5747 5196 5764 5204
rect 5756 5164 5764 5196
rect 5727 5156 5764 5164
rect 4887 5136 5244 5144
rect 5456 5136 5473 5144
rect 5456 5127 5464 5136
rect 5727 5136 5753 5144
rect 147 5116 213 5124
rect 547 5116 593 5124
rect 787 5116 853 5124
rect 907 5116 1133 5124
rect 1147 5116 1313 5124
rect 1327 5116 1353 5124
rect 1707 5116 1773 5124
rect 1787 5116 1873 5124
rect 2387 5116 2493 5124
rect 2507 5116 2553 5124
rect 2627 5116 2673 5124
rect 2687 5116 2713 5124
rect 2927 5116 3133 5124
rect 3387 5116 3513 5124
rect 3527 5116 3553 5124
rect 4187 5116 4313 5124
rect 4327 5116 4453 5124
rect 4627 5116 4713 5124
rect 4727 5116 4753 5124
rect 5087 5116 5193 5124
rect 5487 5116 5513 5124
rect 507 5096 733 5104
rect 767 5096 1033 5104
rect 1047 5096 1133 5104
rect 1147 5096 1273 5104
rect 2127 5096 2153 5104
rect 2167 5096 3033 5104
rect 3727 5096 3913 5104
rect 3927 5096 4833 5104
rect 4947 5096 5133 5104
rect 5207 5096 5333 5104
rect 5507 5096 5753 5104
rect 1127 5076 1153 5084
rect 4007 5076 4393 5084
rect 4407 5076 4853 5084
rect 5067 5076 5233 5084
rect 2367 5056 2653 5064
rect 2667 5056 3933 5064
rect 4107 5056 4913 5064
rect 5347 5056 5453 5064
rect 1787 5036 1913 5044
rect 1927 5036 2093 5044
rect 2107 5036 2433 5044
rect 2847 5036 3833 5044
rect 4247 5036 4613 5044
rect 4627 5036 4653 5044
rect 4727 5036 4893 5044
rect 47 5016 373 5024
rect 1427 5016 2433 5024
rect 2707 5016 2993 5024
rect 3007 5016 3273 5024
rect 4147 5016 4233 5024
rect 3067 4996 3113 5004
rect 3127 4996 3153 5004
rect 3167 4996 3393 5004
rect 3427 4996 3513 5004
rect 3527 4996 3773 5004
rect 3847 4996 4893 5004
rect 5027 4996 5293 5004
rect 87 4976 373 4984
rect 387 4976 413 4984
rect 967 4976 993 4984
rect 1007 4976 1233 4984
rect 1307 4976 1333 4984
rect 1587 4976 1713 4984
rect 1727 4976 1833 4984
rect 2147 4976 2373 4984
rect 2767 4976 2773 4984
rect 2787 4976 2853 4984
rect 3247 4976 3313 4984
rect 3447 4976 3493 4984
rect 3507 4976 3533 4984
rect 3867 4976 3953 4984
rect 3967 4976 4013 4984
rect 4027 4976 4133 4984
rect 4387 4976 4453 4984
rect 4467 4976 4593 4984
rect 4967 4976 5133 4984
rect 5467 4976 5753 4984
rect 176 4956 213 4964
rect 176 4924 184 4956
rect 587 4956 633 4964
rect 707 4956 773 4964
rect 827 4956 893 4964
rect 936 4956 1084 4964
rect 207 4936 233 4944
rect 307 4936 333 4944
rect 396 4927 404 4953
rect 936 4947 944 4956
rect 567 4936 653 4944
rect 807 4936 933 4944
rect 1007 4936 1053 4944
rect 1076 4944 1084 4956
rect 1127 4956 1173 4964
rect 1887 4956 1913 4964
rect 2427 4956 2453 4964
rect 2987 4956 3133 4964
rect 1076 4936 1213 4944
rect 1227 4936 1313 4944
rect 1407 4936 1433 4944
rect 1747 4936 1773 4944
rect 1807 4936 1853 4944
rect 1907 4936 1973 4944
rect 2127 4936 2193 4944
rect 2267 4936 2393 4944
rect 2527 4936 2633 4944
rect 2887 4936 2953 4944
rect 3176 4927 3184 4973
rect 3327 4956 3373 4964
rect 4067 4956 4273 4964
rect 4287 4956 4293 4964
rect 4507 4956 4633 4964
rect 4647 4956 4733 4964
rect 4927 4956 5013 4964
rect 5067 4956 5093 4964
rect 5107 4956 5153 4964
rect 5587 4956 5744 4964
rect 3387 4936 3413 4944
rect 3447 4936 3813 4944
rect 3827 4936 4193 4944
rect 4207 4936 4384 4944
rect 4376 4927 4384 4936
rect 4427 4936 4773 4944
rect 5167 4936 5513 4944
rect 5587 4936 5613 4944
rect 5736 4927 5744 4956
rect 176 4916 213 4924
rect 267 4916 313 4924
rect 327 4916 353 4924
rect 687 4916 773 4924
rect 1467 4916 1493 4924
rect 1507 4916 1533 4924
rect 1647 4916 1813 4924
rect 1927 4916 1953 4924
rect 2167 4916 2493 4924
rect 2547 4916 2593 4924
rect 2767 4916 2873 4924
rect 3527 4916 3573 4924
rect 3756 4916 3833 4924
rect 227 4896 293 4904
rect 607 4896 633 4904
rect 1427 4896 1553 4904
rect 1687 4896 1853 4904
rect 2536 4896 3433 4904
rect 2536 4887 2544 4896
rect 3587 4896 3613 4904
rect 3756 4904 3764 4916
rect 3847 4916 4033 4924
rect 4087 4916 4113 4924
rect 4187 4916 4204 4924
rect 3627 4896 3764 4904
rect 4196 4904 4204 4916
rect 4227 4916 4353 4924
rect 4567 4916 4613 4924
rect 4987 4916 5133 4924
rect 5147 4916 5433 4924
rect 5647 4916 5673 4924
rect 4196 4896 4273 4904
rect 5447 4896 5713 4904
rect 5727 4896 5773 4904
rect 127 4876 293 4884
rect 307 4876 493 4884
rect 1107 4876 1473 4884
rect 3187 4876 3293 4884
rect 3307 4876 3713 4884
rect 4287 4876 4433 4884
rect 5067 4876 5493 4884
rect 2607 4856 3313 4864
rect 3567 4856 3673 4864
rect 3987 4856 5213 4864
rect 147 4836 193 4844
rect 207 4836 553 4844
rect 3147 4836 4613 4844
rect 5187 4836 5233 4844
rect 3707 4816 3873 4824
rect 4347 4816 4493 4824
rect 4507 4816 4593 4824
rect 1827 4796 3433 4804
rect 3807 4796 3953 4804
rect 5087 4796 5613 4804
rect 5627 4796 5773 4804
rect 47 4776 113 4784
rect 187 4776 313 4784
rect 1307 4776 2113 4784
rect 3407 4776 3913 4784
rect 5387 4776 5453 4784
rect 107 4756 153 4764
rect 167 4756 413 4764
rect 427 4756 453 4764
rect 3467 4756 3473 4764
rect 3487 4756 4153 4764
rect 1367 4736 2133 4744
rect 2427 4736 2653 4744
rect 3207 4736 3653 4744
rect 3667 4736 4693 4744
rect 5227 4736 5273 4744
rect 5587 4736 5613 4744
rect 167 4716 193 4724
rect 387 4716 1013 4724
rect 1447 4716 1873 4724
rect 2247 4716 2533 4724
rect 3147 4716 3233 4724
rect 3427 4716 3593 4724
rect 3827 4716 4273 4724
rect 4427 4716 4493 4724
rect 4967 4716 5053 4724
rect 5067 4716 5193 4724
rect 5267 4716 5273 4724
rect 5287 4716 5673 4724
rect 5707 4716 5753 4724
rect 127 4696 264 4704
rect 47 4676 233 4684
rect 256 4664 264 4696
rect 407 4696 504 4704
rect 496 4687 504 4696
rect 527 4696 613 4704
rect 1567 4696 1593 4704
rect 1647 4696 1713 4704
rect 2507 4696 2573 4704
rect 2707 4696 2753 4704
rect 2807 4696 2953 4704
rect 2967 4696 3033 4704
rect 3167 4696 3193 4704
rect 3487 4696 3664 4704
rect 3656 4687 3664 4696
rect 3767 4696 3833 4704
rect 3967 4696 4013 4704
rect 4187 4696 4413 4704
rect 5127 4696 5153 4704
rect 5347 4696 5413 4704
rect 287 4676 373 4684
rect 667 4676 793 4684
rect 807 4676 1013 4684
rect 1167 4676 1213 4684
rect 1267 4676 1353 4684
rect 1367 4676 1493 4684
rect 1547 4676 1573 4684
rect 1787 4676 1993 4684
rect 2087 4676 2353 4684
rect 2407 4676 2433 4684
rect 2527 4676 2813 4684
rect 3087 4676 3253 4684
rect 3347 4676 3413 4684
rect 3507 4676 3633 4684
rect 3767 4676 3853 4684
rect 3867 4676 4173 4684
rect 4307 4676 4333 4684
rect 4347 4676 4433 4684
rect 4487 4676 4533 4684
rect 4707 4676 5033 4684
rect 5087 4676 5173 4684
rect 5316 4684 5324 4693
rect 5316 4676 5433 4684
rect 5456 4684 5464 4693
rect 5456 4676 5553 4684
rect 256 4656 273 4664
rect 467 4656 533 4664
rect 887 4656 1233 4664
rect 1627 4656 1713 4664
rect 1807 4656 1953 4664
rect 2107 4656 2193 4664
rect 2207 4656 2253 4664
rect 2267 4656 2273 4664
rect 2407 4656 2573 4664
rect 2587 4656 2633 4664
rect 2647 4656 2733 4664
rect 2787 4656 2964 4664
rect 127 4636 193 4644
rect 247 4636 313 4644
rect 367 4636 453 4644
rect 1067 4636 1133 4644
rect 1147 4636 1213 4644
rect 1267 4636 1373 4644
rect 1527 4636 1593 4644
rect 1727 4636 2033 4644
rect 2187 4636 2773 4644
rect 2956 4644 2964 4656
rect 3107 4656 3173 4664
rect 3547 4656 3613 4664
rect 4007 4656 4573 4664
rect 4967 4656 5013 4664
rect 5127 4656 5313 4664
rect 5387 4656 5433 4664
rect 5587 4656 5593 4664
rect 5607 4656 5693 4664
rect 5747 4656 5773 4664
rect 2956 4636 3173 4644
rect 3267 4636 3453 4644
rect 3507 4636 3633 4644
rect 3747 4636 3813 4644
rect 3907 4636 4073 4644
rect 4147 4636 4173 4644
rect 4467 4636 4593 4644
rect 4607 4636 4673 4644
rect 4687 4636 4733 4644
rect 4887 4636 5053 4644
rect 5207 4636 5333 4644
rect 5367 4636 5453 4644
rect 267 4616 353 4624
rect 1327 4616 1473 4624
rect 1607 4616 2244 4624
rect 527 4596 833 4604
rect 847 4596 893 4604
rect 907 4596 1673 4604
rect 2236 4604 2244 4616
rect 2327 4616 2673 4624
rect 2927 4616 3353 4624
rect 3787 4616 3893 4624
rect 4096 4616 4253 4624
rect 2236 4596 2513 4604
rect 2687 4596 3293 4604
rect 3307 4596 3653 4604
rect 3727 4596 3933 4604
rect 4096 4604 4104 4616
rect 4827 4616 4933 4624
rect 5027 4616 5513 4624
rect 5527 4616 5713 4624
rect 4047 4596 4104 4604
rect 4247 4596 4533 4604
rect 4907 4596 5073 4604
rect 5327 4596 5393 4604
rect 147 4576 493 4584
rect 1387 4576 1433 4584
rect 1847 4576 2093 4584
rect 2467 4576 2673 4584
rect 2687 4576 2893 4584
rect 2907 4576 3013 4584
rect 4247 4576 4553 4584
rect 4567 4576 4833 4584
rect 247 4556 413 4564
rect 427 4556 693 4564
rect 1007 4556 1933 4564
rect 2287 4556 2593 4564
rect 2767 4556 2833 4564
rect 2847 4556 3213 4564
rect 3827 4556 3933 4564
rect 3947 4556 5293 4564
rect 507 4536 573 4544
rect 647 4536 653 4544
rect 667 4536 853 4544
rect 867 4536 933 4544
rect 1287 4536 1393 4544
rect 1407 4536 1433 4544
rect 1447 4536 1753 4544
rect 1827 4536 2173 4544
rect 3227 4536 3253 4544
rect 4127 4536 4313 4544
rect 4327 4536 4473 4544
rect 5147 4536 5293 4544
rect 587 4516 713 4524
rect 907 4516 1533 4524
rect 1667 4516 1973 4524
rect 2027 4516 2493 4524
rect 2507 4516 2573 4524
rect 2887 4516 2913 4524
rect 3127 4516 3453 4524
rect 3467 4516 3473 4524
rect 3667 4516 4053 4524
rect 4067 4516 4093 4524
rect 4487 4516 5093 4524
rect 5167 4516 5213 4524
rect 5307 4516 5353 4524
rect 5507 4516 5593 4524
rect 107 4496 153 4504
rect 267 4496 353 4504
rect 687 4496 773 4504
rect 787 4496 813 4504
rect 827 4496 893 4504
rect 1187 4496 1273 4504
rect 1296 4496 1313 4504
rect 56 4424 64 4493
rect 116 4476 293 4484
rect 116 4467 124 4476
rect 307 4476 393 4484
rect 607 4476 673 4484
rect 727 4476 824 4484
rect 287 4456 333 4464
rect 387 4456 413 4464
rect 567 4456 693 4464
rect 707 4456 793 4464
rect 816 4464 824 4476
rect 947 4476 1013 4484
rect 1296 4484 1304 4496
rect 1807 4496 2213 4504
rect 2487 4496 2613 4504
rect 2727 4496 2853 4504
rect 3027 4496 3133 4504
rect 3147 4496 3213 4504
rect 3227 4496 3313 4504
rect 3527 4496 3893 4504
rect 4027 4496 4113 4504
rect 4867 4496 5173 4504
rect 5187 4496 5333 4504
rect 1187 4476 1304 4484
rect 1467 4476 1493 4484
rect 1567 4476 1913 4484
rect 1927 4476 2013 4484
rect 2047 4476 2173 4484
rect 2227 4476 2764 4484
rect 2756 4467 2764 4476
rect 2887 4476 2993 4484
rect 3387 4476 3533 4484
rect 3547 4476 3584 4484
rect 816 4456 913 4464
rect 927 4456 993 4464
rect 1047 4456 1153 4464
rect 1207 4456 1333 4464
rect 1347 4456 1413 4464
rect 1447 4456 1713 4464
rect 1847 4456 1933 4464
rect 2067 4456 2153 4464
rect 2367 4456 2413 4464
rect 2447 4456 2473 4464
rect 2527 4456 2733 4464
rect 2947 4456 2973 4464
rect 3356 4464 3364 4473
rect 3356 4456 3553 4464
rect 3576 4464 3584 4476
rect 3607 4476 3633 4484
rect 3707 4476 3793 4484
rect 4267 4476 4393 4484
rect 4427 4476 4524 4484
rect 3576 4456 3753 4464
rect 76 4444 84 4453
rect 3656 4447 3664 4456
rect 3827 4456 3853 4464
rect 4307 4456 4353 4464
rect 4367 4456 4393 4464
rect 4516 4447 4524 4476
rect 4887 4476 4933 4484
rect 4947 4476 4973 4484
rect 5227 4476 5393 4484
rect 5496 4464 5504 4493
rect 5147 4456 5504 4464
rect 5676 4447 5684 4473
rect 76 4436 173 4444
rect 187 4436 213 4444
rect 347 4436 393 4444
rect 467 4436 533 4444
rect 1087 4436 1293 4444
rect 1307 4436 1353 4444
rect 1796 4436 1813 4444
rect 56 4416 73 4424
rect 256 4424 264 4433
rect 1796 4427 1804 4436
rect 2607 4436 2713 4444
rect 3007 4436 3333 4444
rect 3347 4436 3593 4444
rect 3707 4436 3873 4444
rect 4047 4436 4273 4444
rect 4447 4436 4493 4444
rect 4787 4436 4893 4444
rect 4947 4436 5013 4444
rect 5367 4436 5473 4444
rect 256 4416 333 4424
rect 1107 4416 1153 4424
rect 1527 4416 1553 4424
rect 1567 4416 1593 4424
rect 2076 4424 2084 4433
rect 2067 4416 2084 4424
rect 2347 4416 3633 4424
rect 4167 4416 4373 4424
rect 4807 4416 4993 4424
rect 5067 4416 5193 4424
rect 5387 4416 5413 4424
rect 5587 4416 5733 4424
rect 1707 4396 2333 4404
rect 2667 4396 3333 4404
rect 3527 4396 3613 4404
rect 4287 4396 4313 4404
rect 4327 4396 4333 4404
rect 4707 4396 4933 4404
rect 4947 4396 5133 4404
rect 5207 4396 5533 4404
rect 1827 4376 1853 4384
rect 2647 4376 3153 4384
rect 3647 4376 4273 4384
rect 1367 4356 2333 4364
rect 2747 4356 3033 4364
rect 4627 4356 4653 4364
rect 1487 4336 2373 4344
rect 2467 4336 2933 4344
rect 2947 4336 2993 4344
rect 3047 4336 4593 4344
rect 2227 4316 2413 4324
rect 2427 4316 4733 4324
rect 907 4296 2433 4304
rect 2707 4296 4233 4304
rect 4567 4296 4613 4304
rect 4627 4296 4913 4304
rect 5567 4296 5613 4304
rect 1687 4276 1853 4284
rect 2167 4276 2193 4284
rect 2967 4276 3313 4284
rect 387 4256 433 4264
rect 1267 4256 1293 4264
rect 1327 4256 1733 4264
rect 1847 4256 1893 4264
rect 1947 4256 2093 4264
rect 2127 4256 2353 4264
rect 2467 4256 2513 4264
rect 2727 4256 3593 4264
rect 3927 4256 4173 4264
rect 4187 4256 4193 4264
rect 1187 4236 1373 4244
rect 1527 4236 2053 4244
rect 2187 4236 2233 4244
rect 2276 4236 2493 4244
rect 816 4216 1033 4224
rect 816 4207 824 4216
rect 1047 4216 1213 4224
rect 1267 4216 1293 4224
rect 1487 4216 1653 4224
rect 1767 4216 1793 4224
rect 2047 4216 2073 4224
rect 2276 4224 2284 4236
rect 2836 4236 2893 4244
rect 2836 4227 2844 4236
rect 3027 4236 3573 4244
rect 3987 4236 4033 4244
rect 4047 4236 4093 4244
rect 5307 4236 5524 4244
rect 2147 4216 2284 4224
rect 2407 4216 2713 4224
rect 147 4196 213 4204
rect 227 4196 273 4204
rect 467 4196 593 4204
rect 767 4196 813 4204
rect 867 4196 913 4204
rect 1147 4196 1233 4204
rect 47 4176 113 4184
rect 156 4176 173 4184
rect 156 4164 164 4176
rect 267 4176 333 4184
rect 736 4184 744 4193
rect 736 4176 833 4184
rect 1076 4184 1084 4193
rect 1356 4187 1364 4213
rect 2636 4207 2644 4216
rect 2727 4216 2773 4224
rect 2887 4216 2953 4224
rect 3687 4216 3773 4224
rect 3816 4216 3913 4224
rect 1387 4196 1433 4204
rect 1547 4196 1613 4204
rect 1787 4196 1933 4204
rect 1947 4196 1973 4204
rect 2027 4196 2124 4204
rect 2116 4187 2124 4196
rect 2167 4196 2193 4204
rect 2216 4196 2593 4204
rect 1076 4176 1273 4184
rect 1607 4176 1673 4184
rect 1747 4176 1873 4184
rect 2067 4176 2093 4184
rect 2216 4184 2224 4196
rect 2727 4196 2913 4204
rect 3247 4196 3264 4204
rect 2127 4176 2224 4184
rect 2247 4176 2273 4184
rect 2367 4176 2433 4184
rect 2607 4176 3033 4184
rect 147 4156 164 4164
rect 187 4156 233 4164
rect 247 4156 573 4164
rect 827 4156 913 4164
rect 927 4156 933 4164
rect 947 4156 1053 4164
rect 1207 4156 1613 4164
rect 1727 4156 1813 4164
rect 1907 4156 1993 4164
rect 2007 4156 2133 4164
rect 2307 4156 2333 4164
rect 2487 4156 2873 4164
rect 2907 4156 3113 4164
rect 3127 4156 3233 4164
rect 3256 4164 3264 4196
rect 3296 4196 3373 4204
rect 3296 4184 3304 4196
rect 3427 4196 3453 4204
rect 3507 4196 3533 4204
rect 3816 4204 3824 4216
rect 4067 4216 4133 4224
rect 4567 4216 4593 4224
rect 5167 4216 5184 4224
rect 3807 4196 3824 4204
rect 3847 4196 3933 4204
rect 4207 4196 4333 4204
rect 4347 4196 4444 4204
rect 4436 4187 4444 4196
rect 4487 4196 4613 4204
rect 5007 4196 5093 4204
rect 3287 4176 3304 4184
rect 3316 4176 3353 4184
rect 3316 4164 3324 4176
rect 3607 4176 3633 4184
rect 3647 4176 3733 4184
rect 3987 4176 4053 4184
rect 4207 4176 4233 4184
rect 4327 4176 4393 4184
rect 4687 4176 4753 4184
rect 5176 4184 5184 4216
rect 5287 4216 5304 4224
rect 5296 4207 5304 4216
rect 5207 4196 5253 4204
rect 5407 4196 5493 4204
rect 5516 4204 5524 4236
rect 5687 4216 5704 4224
rect 5516 4196 5673 4204
rect 5176 4176 5464 4184
rect 3256 4156 3324 4164
rect 3347 4156 3373 4164
rect 3487 4156 3513 4164
rect 3527 4156 3553 4164
rect 3627 4156 3653 4164
rect 3667 4156 3993 4164
rect 4387 4156 4413 4164
rect 4647 4156 4653 4164
rect 4667 4156 4853 4164
rect 4887 4156 5053 4164
rect 5187 4156 5373 4164
rect 5407 4156 5433 4164
rect 5456 4164 5464 4176
rect 5487 4176 5573 4184
rect 5696 4184 5704 4216
rect 5667 4176 5704 4184
rect 5456 4156 5533 4164
rect 5776 4164 5784 4173
rect 5667 4156 5784 4164
rect 227 4136 253 4144
rect 587 4136 1693 4144
rect 1716 4136 2413 4144
rect 67 4116 113 4124
rect 247 4116 413 4124
rect 427 4116 553 4124
rect 567 4116 653 4124
rect 1107 4116 1253 4124
rect 1567 4116 1613 4124
rect 1716 4124 1724 4136
rect 2427 4136 2553 4144
rect 2687 4136 2713 4144
rect 2867 4136 4493 4144
rect 4507 4136 4713 4144
rect 4827 4136 4993 4144
rect 5227 4136 5373 4144
rect 5727 4136 5773 4144
rect 1647 4116 1724 4124
rect 2407 4116 2513 4124
rect 2527 4116 2693 4124
rect 2767 4116 2953 4124
rect 3087 4116 3133 4124
rect 3167 4116 3213 4124
rect 3247 4116 3493 4124
rect 4307 4116 4333 4124
rect 4407 4116 4573 4124
rect 4587 4116 5113 4124
rect 5367 4116 5473 4124
rect 67 4096 93 4104
rect 107 4096 433 4104
rect 447 4096 453 4104
rect 647 4096 733 4104
rect 747 4096 1973 4104
rect 2067 4096 2253 4104
rect 2327 4096 2413 4104
rect 2847 4096 3053 4104
rect 3067 4096 3193 4104
rect 3287 4096 3393 4104
rect 3447 4096 3493 4104
rect 4167 4096 4293 4104
rect 4947 4096 5113 4104
rect 5127 4096 5233 4104
rect 167 4076 293 4084
rect 1247 4076 2833 4084
rect 2856 4076 3313 4084
rect 367 4056 413 4064
rect 427 4056 593 4064
rect 607 4056 1993 4064
rect 2856 4064 2864 4076
rect 3347 4076 3393 4084
rect 3647 4076 3713 4084
rect 3747 4076 3873 4084
rect 3887 4076 5273 4084
rect 5467 4076 5493 4084
rect 2047 4056 2864 4064
rect 2987 4056 3153 4064
rect 3227 4056 3333 4064
rect 3347 4056 3553 4064
rect 3727 4056 3793 4064
rect 3807 4056 4093 4064
rect 4147 4056 4173 4064
rect 5247 4056 5293 4064
rect 5327 4056 5513 4064
rect 167 4036 193 4044
rect 307 4036 553 4044
rect 567 4036 613 4044
rect 887 4036 953 4044
rect 967 4036 1493 4044
rect 1547 4036 1553 4044
rect 1567 4036 1813 4044
rect 2167 4036 2813 4044
rect 2887 4036 3133 4044
rect 3307 4036 3353 4044
rect 3587 4036 3773 4044
rect 3907 4036 4133 4044
rect 4147 4036 4253 4044
rect 4387 4036 5193 4044
rect 5267 4036 5413 4044
rect 5527 4036 5693 4044
rect 107 4016 173 4024
rect 987 4016 1093 4024
rect 1287 4016 1333 4024
rect 1347 4016 1633 4024
rect 1667 4016 1753 4024
rect 1767 4016 1833 4024
rect 2187 4016 2273 4024
rect 2287 4016 2493 4024
rect 2887 4016 2993 4024
rect 3047 4016 3093 4024
rect 3187 4016 3284 4024
rect 76 3984 84 4013
rect 167 3996 213 4004
rect 607 3996 713 4004
rect 867 3996 913 4004
rect 1407 3996 1453 4004
rect 1467 3996 1613 4004
rect 1887 3996 2293 4004
rect 2307 3996 2333 4004
rect 2387 3996 2433 4004
rect 2647 3996 2673 4004
rect 2827 3996 3253 4004
rect 76 3976 93 3984
rect 207 3976 253 3984
rect 267 3976 333 3984
rect 487 3976 553 3984
rect 747 3976 833 3984
rect 856 3976 1344 3984
rect 147 3956 173 3964
rect 856 3964 864 3976
rect 727 3956 864 3964
rect 987 3956 1073 3964
rect 1227 3956 1313 3964
rect 1336 3964 1344 3976
rect 1647 3976 1693 3984
rect 1867 3976 1893 3984
rect 1987 3976 2073 3984
rect 2207 3976 2233 3984
rect 1336 3956 2133 3964
rect 1167 3936 1313 3944
rect 1387 3936 1553 3944
rect 1987 3936 2013 3944
rect 2156 3944 2164 3973
rect 2416 3964 2424 3973
rect 2327 3956 2424 3964
rect 2476 3964 2484 3993
rect 3276 3987 3284 4016
rect 3327 4016 4713 4024
rect 4767 4016 4913 4024
rect 5167 4016 5413 4024
rect 3447 3996 3753 4004
rect 3947 3996 3973 4004
rect 4027 3996 4073 4004
rect 4087 3996 4333 4004
rect 4547 3996 4593 4004
rect 4667 3996 4973 4004
rect 5307 3996 5333 4004
rect 5347 3996 5513 4004
rect 5567 3996 5733 4004
rect 2507 3976 2613 3984
rect 2627 3976 2753 3984
rect 2787 3976 2913 3984
rect 2967 3976 2993 3984
rect 3327 3976 3413 3984
rect 3536 3976 3833 3984
rect 3536 3967 3544 3976
rect 3847 3976 3953 3984
rect 4007 3976 4113 3984
rect 4127 3976 4233 3984
rect 4247 3976 4353 3984
rect 4407 3976 4433 3984
rect 4516 3984 4524 3993
rect 4516 3976 4873 3984
rect 4816 3967 4824 3976
rect 4907 3976 5013 3984
rect 5036 3976 5113 3984
rect 2476 3956 2493 3964
rect 2527 3956 2553 3964
rect 2607 3956 2633 3964
rect 2767 3956 2793 3964
rect 2987 3956 3033 3964
rect 3267 3956 3484 3964
rect 2696 3944 2704 3953
rect 2156 3936 2873 3944
rect 2936 3944 2944 3953
rect 2936 3936 2953 3944
rect 3067 3936 3453 3944
rect 3476 3944 3484 3956
rect 3587 3956 3673 3964
rect 4007 3956 4033 3964
rect 4687 3956 4753 3964
rect 4767 3956 4773 3964
rect 5036 3964 5044 3976
rect 5427 3976 5493 3984
rect 4947 3956 5044 3964
rect 5147 3956 5713 3964
rect 5756 3964 5764 3973
rect 5747 3956 5764 3964
rect 3476 3936 3713 3944
rect 3867 3936 4193 3944
rect 4207 3936 4213 3944
rect 5107 3936 5653 3944
rect 5767 3936 5813 3944
rect 2467 3916 2613 3924
rect 2627 3916 2673 3924
rect 3007 3916 3493 3924
rect 3787 3916 4473 3924
rect 4727 3916 5133 3924
rect 5687 3916 5713 3924
rect 1307 3896 2993 3904
rect 3027 3896 4413 3904
rect 4747 3896 4913 3904
rect 2407 3876 2453 3884
rect 2487 3876 2513 3884
rect 2547 3876 2613 3884
rect 2667 3876 2953 3884
rect 2967 3876 3224 3884
rect 1107 3856 1253 3864
rect 1687 3856 2753 3864
rect 3216 3864 3224 3876
rect 3247 3876 4333 3884
rect 4387 3876 4853 3884
rect 5227 3876 5393 3884
rect 3216 3856 4813 3864
rect 1307 3836 3113 3844
rect 3147 3836 3233 3844
rect 3267 3836 3373 3844
rect 3827 3836 4253 3844
rect 4267 3836 4533 3844
rect 1087 3816 1173 3824
rect 2387 3816 2733 3824
rect 3307 3816 3333 3824
rect 3527 3816 3893 3824
rect 4707 3816 4853 3824
rect 5447 3816 5813 3824
rect 1047 3796 1213 3804
rect 2067 3796 2073 3804
rect 2087 3796 2393 3804
rect 2487 3796 2653 3804
rect 2827 3796 2953 3804
rect 3127 3796 3353 3804
rect 3647 3796 4593 3804
rect 4687 3796 5133 3804
rect 5147 3796 5253 3804
rect 67 3776 113 3784
rect 2707 3776 3913 3784
rect 3927 3776 4753 3784
rect 5627 3776 5693 3784
rect 127 3756 244 3764
rect 236 3747 244 3756
rect 967 3756 1013 3764
rect 1127 3756 1173 3764
rect 1256 3756 1333 3764
rect 1256 3747 1264 3756
rect 1407 3756 1533 3764
rect 1827 3756 1873 3764
rect 1907 3756 1993 3764
rect 2007 3756 2133 3764
rect 2347 3756 2573 3764
rect 2847 3756 3293 3764
rect 3387 3756 3553 3764
rect 3847 3756 4493 3764
rect 5027 3756 5153 3764
rect 5167 3756 5713 3764
rect 5747 3756 5784 3764
rect 87 3736 184 3744
rect 176 3724 184 3736
rect 207 3736 224 3744
rect 216 3724 224 3736
rect 247 3736 313 3744
rect 667 3736 733 3744
rect 747 3736 993 3744
rect 1167 3736 1193 3744
rect 1347 3736 1433 3744
rect 1687 3736 1873 3744
rect 1887 3736 2033 3744
rect 2067 3736 2173 3744
rect 2327 3736 2424 3744
rect 176 3716 204 3724
rect 216 3716 293 3724
rect 87 3696 133 3704
rect 196 3704 204 3716
rect 427 3716 493 3724
rect 607 3716 813 3724
rect 1116 3724 1124 3733
rect 867 3716 924 3724
rect 1116 3716 1233 3724
rect 196 3696 213 3704
rect 267 3696 333 3704
rect 447 3696 453 3704
rect 467 3696 533 3704
rect 567 3696 713 3704
rect 816 3704 824 3713
rect 747 3696 824 3704
rect 847 3696 893 3704
rect 916 3704 924 3716
rect 1427 3716 1453 3724
rect 1467 3716 1493 3724
rect 916 3696 1013 3704
rect 1376 3704 1384 3713
rect 1147 3696 1384 3704
rect 1396 3704 1404 3713
rect 1516 3707 1524 3733
rect 2416 3727 2424 3736
rect 2576 3736 2693 3744
rect 1587 3716 1733 3724
rect 1907 3716 1993 3724
rect 2107 3716 2273 3724
rect 2467 3716 2553 3724
rect 1396 3696 1433 3704
rect 1567 3696 1753 3704
rect 1967 3696 2093 3704
rect 2127 3696 2293 3704
rect 2576 3704 2584 3736
rect 2807 3736 3033 3744
rect 3247 3736 3313 3744
rect 3367 3736 3413 3744
rect 3467 3736 3573 3744
rect 3727 3736 3773 3744
rect 5067 3736 5233 3744
rect 5247 3736 5493 3744
rect 5627 3736 5753 3744
rect 2687 3716 2704 3724
rect 2487 3696 2584 3704
rect 2696 3704 2704 3716
rect 2727 3716 2833 3724
rect 3076 3724 3084 3733
rect 2927 3716 3213 3724
rect 3347 3716 3433 3724
rect 3747 3716 4013 3724
rect 4027 3716 4133 3724
rect 4436 3724 4444 3733
rect 4416 3716 4444 3724
rect 2696 3696 2713 3704
rect 2947 3696 2993 3704
rect 3047 3696 3113 3704
rect 3647 3696 3693 3704
rect 4087 3696 4213 3704
rect 4376 3687 4384 3713
rect 4416 3704 4424 3716
rect 4527 3716 4633 3724
rect 4807 3716 5033 3724
rect 5247 3716 5293 3724
rect 5307 3716 5364 3724
rect 4407 3696 4424 3704
rect 4447 3696 4453 3704
rect 4467 3696 4653 3704
rect 4747 3696 5153 3704
rect 5356 3704 5364 3716
rect 5447 3716 5544 3724
rect 5356 3696 5513 3704
rect 5536 3704 5544 3716
rect 5776 3724 5784 3756
rect 5747 3716 5784 3724
rect 5536 3696 5713 3704
rect 627 3676 773 3684
rect 1027 3676 1093 3684
rect 1276 3676 1484 3684
rect 1276 3664 1284 3676
rect 587 3656 1284 3664
rect 1296 3656 1393 3664
rect 1296 3644 1304 3656
rect 1476 3664 1484 3676
rect 1507 3676 1653 3684
rect 1987 3676 2033 3684
rect 2047 3676 2593 3684
rect 2707 3676 2793 3684
rect 2807 3676 2833 3684
rect 2987 3676 3133 3684
rect 3307 3676 3333 3684
rect 3567 3676 3613 3684
rect 4427 3676 4473 3684
rect 4567 3676 4633 3684
rect 4887 3676 5073 3684
rect 5087 3676 5113 3684
rect 1476 3656 1933 3664
rect 1947 3656 1993 3664
rect 2267 3656 2513 3664
rect 2527 3656 2633 3664
rect 2647 3656 2933 3664
rect 3087 3656 3733 3664
rect 3807 3656 3833 3664
rect 4147 3656 4753 3664
rect 5567 3656 5673 3664
rect 727 3636 1304 3644
rect 1327 3636 1373 3644
rect 1567 3636 1593 3644
rect 1907 3636 2433 3644
rect 2527 3636 2733 3644
rect 3267 3636 3273 3644
rect 3287 3636 3673 3644
rect 3907 3636 3993 3644
rect 1207 3616 1213 3624
rect 1227 3616 1273 3624
rect 1607 3616 2213 3624
rect 2607 3616 2733 3624
rect 2747 3616 3633 3624
rect 3687 3616 3893 3624
rect 3987 3616 4033 3624
rect 5367 3616 5453 3624
rect 107 3596 213 3604
rect 1387 3596 3073 3604
rect 3107 3596 3873 3604
rect 4167 3596 4673 3604
rect 4747 3596 4773 3604
rect 107 3576 273 3584
rect 307 3576 413 3584
rect 687 3576 893 3584
rect 907 3576 973 3584
rect 1767 3576 2253 3584
rect 2407 3576 2433 3584
rect 2907 3576 3173 3584
rect 3327 3576 3393 3584
rect 3547 3576 3613 3584
rect 3627 3576 3773 3584
rect 4207 3576 4293 3584
rect 4367 3576 4893 3584
rect 5187 3576 5233 3584
rect 147 3556 373 3564
rect 507 3556 1113 3564
rect 1727 3556 1993 3564
rect 2287 3556 3553 3564
rect 3667 3556 4193 3564
rect 4287 3556 4653 3564
rect 5047 3556 5313 3564
rect 116 3536 213 3544
rect 116 3507 124 3536
rect 387 3536 613 3544
rect 967 3536 1053 3544
rect 1667 3536 1713 3544
rect 1927 3536 1953 3544
rect 2187 3536 2333 3544
rect 2347 3536 2393 3544
rect 3007 3536 3033 3544
rect 3067 3536 3393 3544
rect 3427 3536 3493 3544
rect 3707 3536 4053 3544
rect 4167 3536 4213 3544
rect 4267 3536 4573 3544
rect 4687 3536 4693 3544
rect 4707 3536 5333 3544
rect 5387 3536 5633 3544
rect 147 3516 204 3524
rect 196 3507 204 3516
rect 267 3516 293 3524
rect 487 3516 593 3524
rect 927 3516 1093 3524
rect 1107 3516 1153 3524
rect 1347 3516 1413 3524
rect 1536 3516 1673 3524
rect 1536 3507 1544 3516
rect 1847 3516 2013 3524
rect 2067 3516 2153 3524
rect 2167 3516 2293 3524
rect 247 3496 273 3504
rect 407 3496 453 3504
rect 947 3496 993 3504
rect 1287 3496 1333 3504
rect 1587 3496 1613 3504
rect 1787 3496 1853 3504
rect 1887 3496 1913 3504
rect 2027 3496 2093 3504
rect 2147 3496 2173 3504
rect 76 3484 84 3493
rect -24 3476 553 3484
rect 1036 3484 1044 3493
rect 927 3476 1044 3484
rect 1187 3476 1253 3484
rect 1367 3476 1393 3484
rect 1456 3484 1464 3493
rect 1456 3476 1613 3484
rect 1667 3476 1693 3484
rect 1707 3476 1813 3484
rect 1987 3476 2213 3484
rect 2236 3484 2244 3516
rect 2367 3516 2533 3524
rect 2587 3516 2813 3524
rect 2887 3516 3053 3524
rect 3516 3524 3524 3533
rect 3207 3516 3524 3524
rect 3656 3516 3753 3524
rect 3656 3507 3664 3516
rect 3776 3516 3873 3524
rect 2267 3496 2333 3504
rect 2387 3496 2453 3504
rect 2476 3496 2673 3504
rect 2476 3484 2484 3496
rect 2696 3496 2733 3504
rect 2696 3487 2704 3496
rect 2807 3496 2873 3504
rect 3067 3496 3173 3504
rect 3227 3496 3253 3504
rect 3316 3496 3353 3504
rect 2236 3476 2484 3484
rect 2567 3476 2653 3484
rect 2727 3476 2833 3484
rect 2867 3476 3193 3484
rect 3316 3484 3324 3496
rect 3367 3496 3473 3504
rect 3527 3496 3653 3504
rect 3776 3487 3784 3516
rect 4007 3516 4313 3524
rect 4327 3516 4613 3524
rect 5087 3516 5133 3524
rect 5147 3516 5153 3524
rect 5307 3516 5533 3524
rect 5587 3516 5593 3524
rect 5607 3516 5633 3524
rect 3916 3504 3924 3513
rect 3847 3496 4033 3504
rect 4127 3496 4173 3504
rect 4187 3496 4273 3504
rect 4327 3496 4393 3504
rect 4447 3496 4473 3504
rect 4507 3496 4533 3504
rect 4927 3496 4973 3504
rect 5027 3496 5173 3504
rect 5527 3496 5553 3504
rect 5667 3496 5733 3504
rect 3247 3476 3324 3484
rect 3347 3476 3364 3484
rect 147 3456 173 3464
rect 807 3456 893 3464
rect 1107 3456 1293 3464
rect 1436 3464 1444 3473
rect 3356 3467 3364 3476
rect 3387 3476 3453 3484
rect 3507 3476 3764 3484
rect 1427 3456 1444 3464
rect 1647 3456 1753 3464
rect 1947 3456 2353 3464
rect 3027 3456 3053 3464
rect 3127 3456 3204 3464
rect 107 3436 113 3444
rect 567 3436 593 3444
rect 827 3436 873 3444
rect 887 3436 953 3444
rect 1307 3436 1373 3444
rect 2047 3436 2273 3444
rect 3196 3444 3204 3456
rect 3267 3456 3333 3464
rect 3427 3456 3673 3464
rect 3756 3464 3764 3476
rect 3987 3476 4173 3484
rect 4467 3476 4513 3484
rect 4527 3476 4893 3484
rect 4907 3476 4993 3484
rect 5167 3476 5373 3484
rect 5507 3476 5533 3484
rect 3756 3456 3793 3464
rect 4087 3456 4373 3464
rect 4527 3456 4613 3464
rect 4847 3456 5053 3464
rect 5127 3456 5133 3464
rect 5147 3456 5193 3464
rect 5607 3456 5713 3464
rect 2287 3436 3184 3444
rect 3196 3436 3413 3444
rect 2567 3416 2913 3424
rect 3176 3424 3184 3436
rect 3436 3436 3493 3444
rect 3436 3424 3444 3436
rect 4827 3436 5433 3444
rect 5587 3436 5653 3444
rect 3176 3416 3444 3424
rect 3467 3416 3693 3424
rect 4367 3416 4833 3424
rect 1487 3396 2113 3404
rect 3107 3396 3153 3404
rect 3236 3396 3313 3404
rect 2007 3376 2853 3384
rect 3236 3384 3244 3396
rect 3327 3396 3593 3404
rect 3707 3396 3833 3404
rect 2927 3376 3244 3384
rect 3567 3376 3913 3384
rect 4007 3376 4593 3384
rect 5447 3376 5473 3384
rect 1047 3356 2553 3364
rect 2667 3356 3353 3364
rect 3427 3356 4013 3364
rect 4947 3356 4973 3364
rect 2767 3336 2793 3344
rect 2807 3336 3113 3344
rect 3147 3336 3193 3344
rect 3247 3336 3293 3344
rect 3307 3336 4153 3344
rect 1087 3316 1233 3324
rect 2627 3316 2753 3324
rect 3047 3316 3153 3324
rect 3327 3316 3573 3324
rect 4147 3316 4213 3324
rect 367 3296 413 3304
rect 667 3296 673 3304
rect 687 3296 833 3304
rect 847 3296 1353 3304
rect 1787 3296 1933 3304
rect 2087 3296 2313 3304
rect 2327 3296 2413 3304
rect 2687 3296 2873 3304
rect 2927 3296 3324 3304
rect 267 3276 313 3284
rect 327 3276 393 3284
rect 1187 3276 1253 3284
rect 1267 3276 1493 3284
rect 1567 3276 1733 3284
rect 1656 3267 1664 3276
rect 1827 3276 2013 3284
rect 2207 3276 2253 3284
rect 2587 3276 2653 3284
rect 2787 3276 3073 3284
rect 3087 3276 3293 3284
rect 3316 3284 3324 3296
rect 3316 3276 3453 3284
rect 3467 3276 3613 3284
rect 4567 3276 4573 3284
rect 4587 3276 4713 3284
rect 4727 3276 4813 3284
rect 4827 3276 4893 3284
rect 4907 3276 4953 3284
rect 4967 3276 5253 3284
rect 5527 3276 5553 3284
rect 87 3256 273 3264
rect 327 3256 553 3264
rect 707 3256 873 3264
rect 887 3256 913 3264
rect 927 3256 953 3264
rect 1007 3256 1093 3264
rect 1227 3256 1473 3264
rect 1587 3256 1613 3264
rect 1927 3256 2133 3264
rect 2207 3256 2233 3264
rect 2487 3256 2713 3264
rect 2816 3256 2933 3264
rect 2816 3247 2824 3256
rect 2976 3256 3153 3264
rect 107 3236 173 3244
rect 227 3236 313 3244
rect 427 3236 513 3244
rect 1127 3236 1213 3244
rect 1267 3236 1373 3244
rect 1447 3236 1593 3244
rect 1647 3236 1713 3244
rect 1807 3236 2084 3244
rect 147 3216 173 3224
rect 247 3216 273 3224
rect 407 3216 453 3224
rect 727 3216 753 3224
rect 767 3216 913 3224
rect 1236 3224 1244 3233
rect 1187 3216 1244 3224
rect 1527 3216 1673 3224
rect 2076 3224 2084 3236
rect 2107 3236 2173 3244
rect 2767 3236 2793 3244
rect 2847 3236 2913 3244
rect 2076 3216 2193 3224
rect 2247 3216 2293 3224
rect 2407 3216 2573 3224
rect 2596 3224 2604 3233
rect 2596 3216 2693 3224
rect 107 3196 253 3204
rect 887 3196 973 3204
rect 1507 3196 1553 3204
rect 1807 3196 1893 3204
rect 1907 3196 1933 3204
rect 2227 3196 2373 3204
rect 2667 3196 2733 3204
rect 2976 3204 2984 3256
rect 3167 3256 3233 3264
rect 3407 3256 3473 3264
rect 3687 3256 3953 3264
rect 4027 3256 4233 3264
rect 4307 3256 4484 3264
rect 3387 3236 3533 3244
rect 3547 3236 3593 3244
rect 3847 3236 3893 3244
rect 3967 3236 4093 3244
rect 4207 3236 4233 3244
rect 4427 3236 4453 3244
rect 4476 3244 4484 3256
rect 4947 3256 5153 3264
rect 5307 3256 5613 3264
rect 5627 3256 5693 3264
rect 4476 3236 4913 3244
rect 5067 3236 5153 3244
rect 5387 3236 5493 3244
rect 3027 3216 3053 3224
rect 3347 3216 3533 3224
rect 2867 3196 2984 3204
rect 3047 3196 3353 3204
rect 3367 3196 3553 3204
rect 3636 3204 3644 3233
rect 3667 3216 3693 3224
rect 4376 3224 4384 3233
rect 3847 3216 4384 3224
rect 4607 3216 4773 3224
rect 4807 3216 4824 3224
rect 3636 3196 3693 3204
rect 3887 3196 3913 3204
rect 4227 3196 4573 3204
rect 4667 3196 4793 3204
rect 4816 3204 4824 3216
rect 4887 3216 4933 3224
rect 4967 3216 4973 3224
rect 4987 3216 5073 3224
rect 5087 3216 5473 3224
rect 5487 3216 5633 3224
rect 4816 3196 5273 3204
rect 87 3176 113 3184
rect 647 3176 973 3184
rect 1147 3176 1233 3184
rect 1247 3176 1793 3184
rect 2567 3176 2653 3184
rect 2927 3176 3093 3184
rect 3447 3176 3913 3184
rect 4087 3176 4253 3184
rect 4347 3176 4373 3184
rect 4427 3176 4553 3184
rect 4567 3176 4673 3184
rect 867 3156 933 3164
rect 947 3156 993 3164
rect 1007 3156 1213 3164
rect 1767 3156 1893 3164
rect 2327 3156 2613 3164
rect 2627 3156 3093 3164
rect 3147 3156 3193 3164
rect 3207 3156 3353 3164
rect 3527 3156 3613 3164
rect 3627 3156 3773 3164
rect 3807 3156 3993 3164
rect 4047 3156 4413 3164
rect 27 3136 1033 3144
rect 1187 3136 1233 3144
rect 1347 3136 1613 3144
rect 1847 3136 2033 3144
rect 2347 3136 2593 3144
rect 2607 3136 2853 3144
rect 3287 3136 3473 3144
rect 3587 3136 3613 3144
rect 3947 3136 3973 3144
rect 4287 3136 5233 3144
rect 587 3116 1124 3124
rect 867 3096 1073 3104
rect 1116 3104 1124 3116
rect 1147 3116 1293 3124
rect 1407 3116 1533 3124
rect 2187 3116 2253 3124
rect 2367 3116 2433 3124
rect 2527 3116 2573 3124
rect 2707 3116 2753 3124
rect 3047 3116 3213 3124
rect 3347 3116 3433 3124
rect 3707 3116 4073 3124
rect 4187 3116 4253 3124
rect 4267 3116 4453 3124
rect 1116 3096 1593 3104
rect 2147 3096 2513 3104
rect 2647 3096 4193 3104
rect 4207 3096 4333 3104
rect 4367 3096 4433 3104
rect 4447 3096 4713 3104
rect 407 3076 664 3084
rect 367 3056 573 3064
rect 587 3056 633 3064
rect 167 3036 253 3044
rect 307 3036 473 3044
rect 547 3036 613 3044
rect 656 3027 664 3076
rect 1027 3076 1153 3084
rect 1507 3076 1733 3084
rect 1747 3076 1933 3084
rect 2047 3076 2113 3084
rect 2127 3076 2633 3084
rect 2687 3076 2773 3084
rect 2787 3076 2873 3084
rect 2887 3076 2933 3084
rect 3167 3076 3273 3084
rect 3287 3076 3393 3084
rect 3887 3076 4213 3084
rect 687 3056 1173 3064
rect 1287 3056 1313 3064
rect 1527 3056 1573 3064
rect 1587 3056 1673 3064
rect 1987 3056 2073 3064
rect 2087 3056 2353 3064
rect 2487 3056 2553 3064
rect 2587 3056 2953 3064
rect 716 3036 773 3044
rect -24 3016 13 3024
rect 327 3016 513 3024
rect 567 3016 653 3024
rect 127 2996 213 3004
rect 267 2996 413 3004
rect 716 3004 724 3036
rect 827 3036 944 3044
rect 936 3027 944 3036
rect 967 3036 1293 3044
rect 1336 3036 1633 3044
rect 1336 3027 1344 3036
rect 1847 3036 1924 3044
rect 1916 3027 1924 3036
rect 2027 3036 2233 3044
rect 2416 3044 2424 3053
rect 2416 3036 2653 3044
rect 747 3016 753 3024
rect 767 3016 793 3024
rect 987 3016 1033 3024
rect 1547 3016 1653 3024
rect 1727 3016 1773 3024
rect 1827 3016 1873 3024
rect 2127 3016 2253 3024
rect 667 2996 724 3004
rect 836 3004 844 3013
rect 807 2996 844 3004
rect 1096 2987 1104 3013
rect 1167 2996 1413 3004
rect 1427 2996 1473 3004
rect 1707 2996 1733 3004
rect 2276 3004 2284 3033
rect 2416 3027 2424 3036
rect 2367 3016 2393 3024
rect 2456 3016 2533 3024
rect 2456 3004 2464 3016
rect 2696 3007 2704 3056
rect 2987 3056 3164 3064
rect 2787 3036 2844 3044
rect 2736 3024 2744 3033
rect 2836 3024 2844 3036
rect 2867 3036 2973 3044
rect 3087 3036 3133 3044
rect 3156 3044 3164 3056
rect 3267 3056 3653 3064
rect 3767 3056 3833 3064
rect 3847 3056 3993 3064
rect 4107 3056 4293 3064
rect 4367 3056 4393 3064
rect 4727 3056 5113 3064
rect 5187 3056 5264 3064
rect 3156 3036 3373 3044
rect 3507 3036 3544 3044
rect 2736 3016 2784 3024
rect 2836 3016 2873 3024
rect 2167 2996 2464 3004
rect 2487 2996 2673 3004
rect 2776 3004 2784 3016
rect 3536 3024 3544 3036
rect 3567 3036 3633 3044
rect 3827 3036 3873 3044
rect 3907 3036 3933 3044
rect 4007 3036 4033 3044
rect 3407 3016 3524 3024
rect 3536 3016 3773 3024
rect 3516 3007 3524 3016
rect 4056 3024 4064 3053
rect 5256 3047 5264 3056
rect 5367 3056 5533 3064
rect 4227 3036 4433 3044
rect 4447 3036 4473 3044
rect 4707 3036 4753 3044
rect 4787 3036 4993 3044
rect 5047 3036 5133 3044
rect 5527 3036 5673 3044
rect 3847 3016 4064 3024
rect 4156 3024 4164 3033
rect 4156 3016 4533 3024
rect 4616 3007 4624 3033
rect 4647 3016 4893 3024
rect 5207 3016 5613 3024
rect 2776 2996 3073 3004
rect 3087 2996 3233 3004
rect 3407 2996 3453 3004
rect 3547 2996 3673 3004
rect 3687 2996 3893 3004
rect 4207 2996 4353 3004
rect 4367 2996 4373 3004
rect 4827 2996 4873 3004
rect 5027 2996 5113 3004
rect 87 2976 113 2984
rect 227 2976 373 2984
rect 767 2976 1073 2984
rect 1567 2976 1693 2984
rect 1707 2976 1973 2984
rect 2727 2976 3113 2984
rect 3887 2976 3953 2984
rect 3967 2976 4113 2984
rect 4127 2976 4233 2984
rect 4927 2976 4973 2984
rect 4987 2976 5173 2984
rect 667 2956 1113 2964
rect 1127 2956 1273 2964
rect 1507 2956 1653 2964
rect 2207 2956 2713 2964
rect 2907 2956 3433 2964
rect 3676 2956 4793 2964
rect 607 2936 713 2944
rect 727 2936 1153 2944
rect 1987 2936 3293 2944
rect 3676 2944 3684 2956
rect 3387 2936 3684 2944
rect 3716 2936 3813 2944
rect 1047 2916 1393 2924
rect 2247 2916 2433 2924
rect 2447 2916 2593 2924
rect 2987 2916 3133 2924
rect 3716 2924 3724 2936
rect 4427 2936 4733 2944
rect 3176 2916 3724 2924
rect 487 2896 2133 2904
rect 3176 2904 3184 2916
rect 5467 2916 5493 2924
rect 5587 2916 5733 2924
rect 2207 2896 3184 2904
rect 3847 2896 4013 2904
rect 1627 2876 2853 2884
rect 2867 2876 2893 2884
rect 3147 2876 4013 2884
rect 1927 2856 2033 2864
rect 2787 2856 2873 2864
rect 1167 2836 2953 2844
rect 2967 2836 3273 2844
rect 3307 2836 3713 2844
rect 3727 2836 4453 2844
rect 5447 2836 5493 2844
rect 507 2816 853 2824
rect 1307 2816 2053 2824
rect 2127 2816 2173 2824
rect 2587 2816 3033 2824
rect 3127 2816 3853 2824
rect 3867 2816 3873 2824
rect 4267 2816 4613 2824
rect 87 2796 253 2804
rect 787 2796 813 2804
rect 827 2796 893 2804
rect 1947 2796 1993 2804
rect 2187 2796 2313 2804
rect 2447 2796 2753 2804
rect 2847 2796 2913 2804
rect 3187 2796 3253 2804
rect 3487 2796 3513 2804
rect 3667 2796 3733 2804
rect 3947 2796 3973 2804
rect 4007 2796 4293 2804
rect 76 2776 113 2784
rect 76 2744 84 2776
rect 316 2776 373 2784
rect 316 2764 324 2776
rect 627 2776 713 2784
rect 727 2776 793 2784
rect 807 2776 893 2784
rect 947 2776 1073 2784
rect 1327 2776 2013 2784
rect 2227 2776 2373 2784
rect 2387 2776 2453 2784
rect 2647 2776 2673 2784
rect 2767 2776 2993 2784
rect 3007 2776 3033 2784
rect 3087 2776 3113 2784
rect 3167 2776 3213 2784
rect 3236 2776 3313 2784
rect 107 2756 324 2764
rect 347 2756 413 2764
rect 467 2756 533 2764
rect 607 2756 653 2764
rect 847 2756 933 2764
rect 1287 2756 1333 2764
rect 1347 2756 1373 2764
rect 1427 2756 1473 2764
rect 1487 2756 1513 2764
rect 1636 2756 1813 2764
rect 1636 2747 1644 2756
rect 1827 2756 1953 2764
rect 2196 2764 2204 2773
rect 2196 2756 2224 2764
rect 2216 2747 2224 2756
rect 2367 2756 2413 2764
rect 2427 2756 2653 2764
rect 2816 2756 2833 2764
rect 76 2736 93 2744
rect 127 2736 153 2744
rect 227 2736 493 2744
rect 567 2736 573 2744
rect 587 2736 673 2744
rect 747 2736 773 2744
rect 1007 2736 1313 2744
rect 1407 2736 1493 2744
rect 1567 2736 1633 2744
rect 1656 2736 1773 2744
rect 207 2716 393 2724
rect 487 2716 753 2724
rect 907 2716 953 2724
rect 1656 2724 1664 2736
rect 1967 2736 1993 2744
rect 2167 2736 2193 2744
rect 2467 2736 2693 2744
rect 1347 2716 1664 2724
rect 1687 2716 1833 2724
rect 2307 2716 2653 2724
rect 2816 2707 2824 2756
rect 3236 2764 3244 2776
rect 3387 2776 3413 2784
rect 3447 2776 3693 2784
rect 3827 2776 3993 2784
rect 4027 2776 4153 2784
rect 4167 2776 4173 2784
rect 4227 2776 4253 2784
rect 4967 2776 5133 2784
rect 5187 2776 5864 2784
rect 3036 2756 3244 2764
rect 3036 2747 3044 2756
rect 3727 2756 3753 2764
rect 3987 2756 4093 2764
rect 4107 2756 4193 2764
rect 4247 2756 4413 2764
rect 2847 2736 2913 2744
rect 3107 2736 3133 2744
rect 3247 2736 3313 2744
rect 3336 2744 3344 2753
rect 4596 2747 4604 2773
rect 4987 2756 5013 2764
rect 5067 2756 5153 2764
rect 5176 2756 5313 2764
rect 5176 2747 5184 2756
rect 3336 2736 3433 2744
rect 3527 2736 3593 2744
rect 3627 2736 3673 2744
rect 3687 2736 3733 2744
rect 3787 2736 4253 2744
rect 4707 2736 4773 2744
rect 4967 2736 4993 2744
rect 5327 2736 5353 2744
rect 5487 2736 5533 2744
rect 5636 2744 5644 2753
rect 5636 2736 5673 2744
rect 2887 2716 2913 2724
rect 2927 2716 2993 2724
rect 3267 2716 3344 2724
rect 447 2696 633 2704
rect 647 2696 733 2704
rect 747 2696 933 2704
rect 1307 2696 1653 2704
rect 1767 2696 1793 2704
rect 2267 2696 2313 2704
rect 2327 2696 2473 2704
rect 2507 2696 2733 2704
rect 3336 2704 3344 2716
rect 3367 2716 3413 2724
rect 3427 2716 3493 2724
rect 3507 2716 3573 2724
rect 3687 2716 4073 2724
rect 4127 2716 4233 2724
rect 4407 2716 4533 2724
rect 4547 2716 4913 2724
rect 5007 2716 5613 2724
rect 3336 2696 3453 2704
rect 3607 2696 3793 2704
rect 3927 2696 4053 2704
rect 4107 2696 4133 2704
rect 5227 2696 5353 2704
rect 5547 2696 5653 2704
rect 547 2676 673 2684
rect 727 2676 873 2684
rect 1207 2676 2933 2684
rect 3067 2676 3293 2684
rect 3327 2676 3393 2684
rect 3487 2676 3553 2684
rect 3567 2676 3633 2684
rect 3707 2676 3993 2684
rect 4567 2676 4813 2684
rect 4827 2676 5053 2684
rect 5067 2676 5193 2684
rect 5207 2676 5433 2684
rect 5447 2676 5613 2684
rect 187 2656 273 2664
rect 287 2656 353 2664
rect 367 2656 633 2664
rect 1247 2656 1353 2664
rect 1367 2656 1593 2664
rect 1607 2656 1684 2664
rect 1587 2636 1653 2644
rect 1676 2644 1684 2656
rect 1787 2656 1913 2664
rect 2107 2656 3173 2664
rect 3347 2656 3373 2664
rect 3487 2656 3533 2664
rect 3587 2656 3884 2664
rect 1676 2636 3833 2644
rect 3876 2644 3884 2656
rect 3987 2656 4513 2664
rect 3876 2636 3953 2644
rect 1587 2616 1913 2624
rect 1927 2616 2513 2624
rect 2527 2616 3833 2624
rect 3847 2616 4573 2624
rect 167 2596 373 2604
rect 807 2596 993 2604
rect 1187 2596 1644 2604
rect 247 2576 473 2584
rect 487 2576 533 2584
rect 667 2576 753 2584
rect 767 2576 873 2584
rect 1107 2576 1173 2584
rect 1636 2584 1644 2596
rect 1667 2596 1693 2604
rect 1867 2596 1933 2604
rect 2207 2596 2313 2604
rect 2327 2596 2413 2604
rect 2587 2596 2613 2604
rect 2647 2596 2973 2604
rect 3007 2596 3193 2604
rect 3247 2596 4633 2604
rect 1636 2576 1973 2584
rect 2067 2576 2273 2584
rect 2367 2576 2553 2584
rect 2727 2576 2744 2584
rect 316 2556 393 2564
rect 187 2536 293 2544
rect 316 2544 324 2556
rect 656 2556 673 2564
rect 307 2536 324 2544
rect 347 2536 373 2544
rect 387 2536 433 2544
rect 656 2544 664 2556
rect 827 2556 973 2564
rect 996 2556 1093 2564
rect 567 2536 664 2544
rect 747 2536 773 2544
rect 887 2536 913 2544
rect 996 2544 1004 2556
rect 1427 2556 1693 2564
rect 1827 2556 1873 2564
rect 2147 2556 2233 2564
rect 2387 2556 2433 2564
rect 2627 2556 2673 2564
rect 2696 2556 2713 2564
rect 947 2536 1004 2544
rect 1127 2536 1193 2544
rect 1247 2536 1413 2544
rect 1547 2536 1613 2544
rect 1767 2536 1793 2544
rect 127 2516 173 2524
rect 287 2516 353 2524
rect 367 2516 413 2524
rect 987 2516 1033 2524
rect 1287 2516 1353 2524
rect 1527 2516 1553 2524
rect 1647 2516 1993 2524
rect 2016 2524 2024 2553
rect 2047 2536 2093 2544
rect 2127 2536 2144 2544
rect 2016 2516 2113 2524
rect 2136 2524 2144 2536
rect 2167 2536 2333 2544
rect 2507 2536 2593 2544
rect 2696 2544 2704 2556
rect 2736 2544 2744 2576
rect 2787 2576 3713 2584
rect 3767 2576 3813 2584
rect 3867 2576 3913 2584
rect 2847 2556 2884 2564
rect 2876 2547 2884 2556
rect 3107 2556 3153 2564
rect 3207 2556 3273 2564
rect 3387 2556 3473 2564
rect 3667 2556 3744 2564
rect 2616 2536 2704 2544
rect 2716 2536 2744 2544
rect 2136 2516 2164 2524
rect 2156 2507 2164 2516
rect 2187 2516 2293 2524
rect 2367 2516 2393 2524
rect 2447 2516 2473 2524
rect 2616 2524 2624 2536
rect 2716 2527 2724 2536
rect 2827 2536 2853 2544
rect 2947 2536 2973 2544
rect 3047 2536 3264 2544
rect 3256 2527 3264 2536
rect 3736 2527 3744 2556
rect 3807 2536 3853 2544
rect 3896 2544 3904 2553
rect 3896 2536 3913 2544
rect 4087 2536 4253 2544
rect 4267 2536 5233 2544
rect 5387 2536 5453 2544
rect 5467 2536 5493 2544
rect 5607 2536 5713 2544
rect 2507 2516 2624 2524
rect 3167 2516 3213 2524
rect 3287 2516 3353 2524
rect 3447 2516 3613 2524
rect 3627 2516 3704 2524
rect 1227 2496 1333 2504
rect 1347 2496 1473 2504
rect 1547 2496 1573 2504
rect 1727 2496 1793 2504
rect 2447 2496 2453 2504
rect 2467 2496 2753 2504
rect 3187 2496 3213 2504
rect 3236 2496 3353 2504
rect 1567 2476 1733 2484
rect 1747 2476 1764 2484
rect 1807 2476 1833 2484
rect 1856 2476 1893 2484
rect 1507 2456 1693 2464
rect 1856 2464 1864 2476
rect 1907 2476 2253 2484
rect 2347 2476 2493 2484
rect 2607 2476 2693 2484
rect 3236 2484 3244 2496
rect 3396 2504 3404 2513
rect 3396 2496 3513 2504
rect 3527 2496 3673 2504
rect 3696 2504 3704 2516
rect 3767 2516 3793 2524
rect 3867 2516 4033 2524
rect 3696 2496 3813 2504
rect 3947 2496 4453 2504
rect 3207 2476 3244 2484
rect 3347 2476 3473 2484
rect 3587 2476 3653 2484
rect 3787 2476 4013 2484
rect 4467 2476 5193 2484
rect 1747 2456 1864 2464
rect 1887 2456 2213 2464
rect 2247 2456 3073 2464
rect 3307 2456 3433 2464
rect 4527 2456 4833 2464
rect 167 2436 253 2444
rect 767 2436 893 2444
rect 1207 2436 1873 2444
rect 2076 2436 2773 2444
rect 2076 2424 2084 2436
rect 3176 2436 3393 2444
rect 1007 2416 2084 2424
rect 2107 2416 2553 2424
rect 3176 2424 3184 2436
rect 3427 2436 3713 2444
rect 4327 2436 4413 2444
rect 4427 2436 4473 2444
rect 4987 2436 5133 2444
rect 3027 2416 3184 2424
rect 3207 2416 3744 2424
rect 1107 2396 2833 2404
rect 3267 2396 3673 2404
rect 3736 2404 3744 2416
rect 3827 2416 5413 2424
rect 3736 2396 4093 2404
rect 4107 2396 4413 2404
rect 4427 2396 4693 2404
rect 4707 2396 4793 2404
rect 1467 2376 1973 2384
rect 2187 2376 2373 2384
rect 3107 2376 3633 2384
rect 3667 2376 3693 2384
rect 4627 2376 5413 2384
rect 5427 2376 5493 2384
rect 1647 2356 1684 2364
rect 1407 2336 1653 2344
rect 1676 2344 1684 2356
rect 1767 2356 2133 2364
rect 2527 2356 3193 2364
rect 3247 2356 3333 2364
rect 3387 2356 3453 2364
rect 3767 2356 3993 2364
rect 4687 2356 4853 2364
rect 4867 2356 5273 2364
rect 1676 2336 1713 2344
rect 1727 2336 1833 2344
rect 2127 2336 3173 2344
rect 3207 2336 3853 2344
rect 3967 2336 4253 2344
rect 4867 2336 5073 2344
rect 5327 2336 5633 2344
rect 307 2316 353 2324
rect 1607 2316 2053 2324
rect 2167 2316 2193 2324
rect 2987 2316 3044 2324
rect -24 2284 -16 2304
rect 87 2296 224 2304
rect 216 2287 224 2296
rect 247 2296 313 2304
rect 687 2296 893 2304
rect 907 2296 1013 2304
rect 1127 2296 1253 2304
rect 1347 2296 1413 2304
rect 1447 2296 1473 2304
rect 1727 2296 1864 2304
rect 1856 2287 1864 2296
rect 1887 2296 1913 2304
rect 1927 2296 2013 2304
rect 2147 2296 2653 2304
rect 2807 2296 3013 2304
rect 3036 2304 3044 2316
rect 3067 2316 3473 2324
rect 4387 2316 4433 2324
rect 4447 2316 4553 2324
rect 4647 2316 4893 2324
rect 5387 2316 5553 2324
rect 3036 2296 3273 2304
rect 3327 2296 3373 2304
rect 3407 2296 3573 2304
rect 3716 2296 3793 2304
rect -24 2276 93 2284
rect 236 2276 333 2284
rect -24 2256 73 2264
rect 236 2264 244 2276
rect 427 2276 453 2284
rect 827 2276 853 2284
rect 1287 2276 1453 2284
rect 1527 2276 1553 2284
rect 1567 2276 1713 2284
rect 1887 2276 2073 2284
rect 2467 2276 2533 2284
rect 2787 2276 2804 2284
rect 167 2256 244 2264
rect 267 2256 293 2264
rect 307 2256 313 2264
rect 636 2264 644 2273
rect 447 2256 644 2264
rect 967 2256 1153 2264
rect 1507 2256 1693 2264
rect 1736 2247 1744 2273
rect 1807 2256 1893 2264
rect 1927 2256 2033 2264
rect 2047 2256 2113 2264
rect 2647 2256 2773 2264
rect 2796 2264 2804 2276
rect 2847 2276 3033 2284
rect 3267 2276 3293 2284
rect 3307 2276 3413 2284
rect 3716 2284 3724 2296
rect 3847 2296 4013 2304
rect 4487 2296 4733 2304
rect 4907 2296 4933 2304
rect 5247 2296 5273 2304
rect 5467 2296 5513 2304
rect 5527 2296 5713 2304
rect 3676 2276 3724 2284
rect 3676 2267 3684 2276
rect 3747 2276 3893 2284
rect 4287 2276 4353 2284
rect 4827 2276 4913 2284
rect 4927 2276 5053 2284
rect 5107 2276 5133 2284
rect 5567 2276 5573 2284
rect 5587 2276 5664 2284
rect 2796 2256 2893 2264
rect 3047 2256 3193 2264
rect 3227 2256 3273 2264
rect 3507 2256 3533 2264
rect 3587 2256 3633 2264
rect 3707 2256 4164 2264
rect 4156 2247 4164 2256
rect 4187 2256 4393 2264
rect 4596 2247 4604 2273
rect 5656 2267 5664 2276
rect 5707 2276 5733 2284
rect 4627 2256 4713 2264
rect 4887 2256 4973 2264
rect 5127 2256 5213 2264
rect 5407 2256 5453 2264
rect 387 2236 473 2244
rect 507 2236 533 2244
rect 547 2236 653 2244
rect 1047 2236 1073 2244
rect 1307 2236 1433 2244
rect 1447 2236 1573 2244
rect 1767 2236 2173 2244
rect 2276 2236 2333 2244
rect 467 2216 513 2224
rect 587 2216 633 2224
rect 1067 2216 1093 2224
rect 1187 2216 1293 2224
rect 1427 2216 1513 2224
rect 1627 2216 1753 2224
rect 1796 2216 1813 2224
rect 347 2196 593 2204
rect 627 2196 773 2204
rect 1796 2204 1804 2216
rect 2276 2224 2284 2236
rect 2727 2236 2913 2244
rect 2927 2236 3113 2244
rect 3167 2236 3193 2244
rect 3507 2236 3653 2244
rect 3787 2236 3833 2244
rect 4847 2236 4933 2244
rect 5147 2236 5393 2244
rect 5527 2236 5633 2244
rect 5647 2236 5713 2244
rect 2107 2216 2284 2224
rect 2347 2216 2593 2224
rect 2727 2216 2853 2224
rect 2947 2216 3313 2224
rect 3327 2216 3393 2224
rect 3667 2216 4373 2224
rect 1727 2196 1804 2204
rect 1827 2196 1993 2204
rect 2787 2196 3513 2204
rect 3527 2196 3793 2204
rect 4547 2196 4573 2204
rect 4587 2196 5033 2204
rect 5227 2196 5353 2204
rect 5687 2196 5733 2204
rect 427 2176 473 2184
rect 1847 2176 1893 2184
rect 2287 2176 2513 2184
rect 2567 2176 3133 2184
rect 3267 2176 3333 2184
rect 3367 2176 3393 2184
rect 3427 2176 3593 2184
rect 3787 2176 3813 2184
rect 4727 2176 4893 2184
rect 5047 2176 5733 2184
rect 127 2156 1873 2164
rect 2167 2156 2233 2164
rect 2247 2156 2433 2164
rect 2447 2156 3433 2164
rect 3447 2156 3953 2164
rect 4047 2156 4633 2164
rect 5007 2156 5533 2164
rect 587 2136 913 2144
rect 1487 2136 1593 2144
rect 2436 2136 3033 2144
rect 87 2116 793 2124
rect 927 2116 1353 2124
rect 1587 2116 1773 2124
rect 1867 2116 1933 2124
rect 2436 2124 2444 2136
rect 3456 2136 4513 2144
rect 1987 2116 2444 2124
rect 2627 2116 2893 2124
rect 2967 2116 3293 2124
rect 3456 2124 3464 2136
rect 4967 2136 5053 2144
rect 5547 2136 5753 2144
rect 5767 2136 5813 2144
rect 3327 2116 3464 2124
rect 3487 2116 4053 2124
rect 5027 2116 5073 2124
rect 5107 2116 5113 2124
rect 5127 2116 5153 2124
rect 5247 2116 5433 2124
rect 5696 2116 5764 2124
rect 207 2096 273 2104
rect 307 2096 373 2104
rect 807 2096 893 2104
rect 1287 2096 1393 2104
rect 1527 2096 1693 2104
rect 1707 2096 1773 2104
rect 1787 2096 1893 2104
rect 2427 2096 2753 2104
rect 2867 2096 2913 2104
rect 3187 2096 3273 2104
rect 3287 2096 3344 2104
rect 427 2076 613 2084
rect 687 2076 753 2084
rect 847 2076 1113 2084
rect 1147 2076 1213 2084
rect 1267 2076 1393 2084
rect 1407 2076 1473 2084
rect 1496 2076 1653 2084
rect 1496 2067 1504 2076
rect 1687 2076 1933 2084
rect 2007 2076 2093 2084
rect 2207 2076 2884 2084
rect 2876 2067 2884 2076
rect 3227 2076 3253 2084
rect 3336 2084 3344 2096
rect 3367 2096 3533 2104
rect 3587 2096 3673 2104
rect 4087 2096 4253 2104
rect 4467 2096 4513 2104
rect 4707 2096 4773 2104
rect 4827 2096 5153 2104
rect 5207 2096 5273 2104
rect 5387 2096 5433 2104
rect 5636 2096 5673 2104
rect 3336 2076 3453 2084
rect 3467 2076 3524 2084
rect 3516 2067 3524 2076
rect 3647 2076 3793 2084
rect 3807 2076 3833 2084
rect 3987 2076 4013 2084
rect 4107 2076 4133 2084
rect 4147 2076 4213 2084
rect 4387 2076 4473 2084
rect 4496 2076 4553 2084
rect 4496 2067 4504 2076
rect 4887 2076 4913 2084
rect 4936 2076 5013 2084
rect 4936 2067 4944 2076
rect 5176 2084 5184 2093
rect 5156 2076 5184 2084
rect 5156 2067 5164 2076
rect 5267 2076 5353 2084
rect 5636 2067 5644 2096
rect 407 2056 473 2064
rect 827 2056 913 2064
rect 1007 2056 1073 2064
rect 1087 2056 1193 2064
rect 1247 2056 1273 2064
rect 1287 2056 1373 2064
rect 1547 2056 1633 2064
rect 1687 2056 1873 2064
rect 1927 2056 2053 2064
rect 2087 2056 2113 2064
rect 2487 2056 2613 2064
rect 2927 2056 3033 2064
rect 3247 2056 3273 2064
rect 3567 2056 3713 2064
rect 3847 2056 3993 2064
rect 4007 2056 4013 2064
rect 4207 2056 4253 2064
rect 4407 2056 4433 2064
rect 4547 2056 4633 2064
rect 4767 2056 4893 2064
rect 5187 2056 5313 2064
rect 5527 2056 5544 2064
rect 207 2036 233 2044
rect 256 2024 264 2053
rect 296 2044 304 2053
rect 296 2036 513 2044
rect 787 2036 853 2044
rect 907 2036 1053 2044
rect 1667 2036 1693 2044
rect 1767 2036 2073 2044
rect 2307 2036 3184 2044
rect 256 2016 293 2024
rect 307 2016 353 2024
rect 427 2016 713 2024
rect 827 2016 933 2024
rect 1096 2024 1104 2033
rect 967 2016 1613 2024
rect 1687 2016 1833 2024
rect 1856 2016 2353 2024
rect 1856 2004 1864 2016
rect 2847 2016 3053 2024
rect 3176 2024 3184 2036
rect 3207 2036 3313 2044
rect 3347 2036 3553 2044
rect 3627 2036 3813 2044
rect 3827 2036 3933 2044
rect 4067 2036 4113 2044
rect 4627 2036 4733 2044
rect 4747 2036 4853 2044
rect 5087 2036 5193 2044
rect 5487 2036 5513 2044
rect 5536 2044 5544 2056
rect 5696 2047 5704 2116
rect 5716 2096 5733 2104
rect 5716 2067 5724 2096
rect 5756 2084 5764 2116
rect 5747 2076 5764 2084
rect 5536 2036 5673 2044
rect 5747 2036 5773 2044
rect 3176 2016 3593 2024
rect 3607 2016 3653 2024
rect 3787 2016 4273 2024
rect 4627 2016 4713 2024
rect 4767 2016 4813 2024
rect 5027 2016 5233 2024
rect 5427 2016 5473 2024
rect 5487 2016 5713 2024
rect 127 1996 1864 2004
rect 2307 1996 2373 2004
rect 2967 1996 3033 2004
rect 3067 1996 3673 2004
rect 3687 1996 3913 2004
rect 3947 1996 4653 2004
rect 1487 1976 1713 1984
rect 2027 1976 3253 1984
rect 3467 1976 3713 1984
rect 4307 1976 5693 1984
rect 287 1956 333 1964
rect 1847 1956 2253 1964
rect 2627 1956 2773 1964
rect 2787 1956 3073 1964
rect 3087 1956 4293 1964
rect 387 1936 653 1944
rect 1407 1936 1573 1944
rect 1767 1936 1973 1944
rect 2067 1936 2333 1944
rect 2607 1936 2713 1944
rect 3027 1936 3173 1944
rect 3647 1936 4093 1944
rect 4107 1936 4244 1944
rect 1927 1916 3493 1924
rect 3547 1916 4153 1924
rect 4236 1924 4244 1936
rect 4236 1916 4313 1924
rect 4327 1916 4413 1924
rect 5087 1916 5253 1924
rect 2427 1896 2553 1904
rect 2707 1896 3613 1904
rect 3707 1896 4133 1904
rect 4227 1896 5293 1904
rect 407 1876 513 1884
rect 1027 1876 1933 1884
rect 1987 1876 2793 1884
rect 2827 1876 3153 1884
rect 3807 1876 4033 1884
rect 4067 1876 4173 1884
rect 4187 1876 4713 1884
rect 4807 1876 5493 1884
rect 227 1856 713 1864
rect 1707 1856 1853 1864
rect 2827 1856 2993 1864
rect 3507 1856 4213 1864
rect 4727 1856 4893 1864
rect 4907 1856 5253 1864
rect 5267 1856 5333 1864
rect 5367 1856 5393 1864
rect 207 1836 333 1844
rect 347 1836 493 1844
rect 727 1836 1133 1844
rect 1247 1836 2113 1844
rect 2227 1836 2613 1844
rect 2767 1836 3373 1844
rect 3387 1836 3613 1844
rect 3867 1836 4013 1844
rect 4127 1836 4173 1844
rect 4187 1836 4273 1844
rect 4367 1836 4453 1844
rect 4507 1836 4553 1844
rect 4687 1836 4853 1844
rect 4987 1836 5033 1844
rect 5347 1836 5433 1844
rect 127 1816 213 1824
rect 247 1816 264 1824
rect 107 1796 193 1804
rect 236 1784 244 1793
rect 147 1776 244 1784
rect 127 1756 213 1764
rect 256 1744 264 1816
rect 376 1804 384 1813
rect 356 1796 384 1804
rect 356 1787 364 1796
rect 416 1784 424 1813
rect 387 1776 424 1784
rect 516 1784 524 1833
rect 547 1816 953 1824
rect 1867 1816 1953 1824
rect 1967 1816 2153 1824
rect 2207 1816 2253 1824
rect 2787 1816 2833 1824
rect 2887 1816 3033 1824
rect 3056 1816 3093 1824
rect 567 1796 593 1804
rect 607 1796 833 1804
rect 947 1796 1033 1804
rect 1107 1796 1173 1804
rect 1187 1796 1233 1804
rect 1287 1796 1333 1804
rect 1647 1796 1753 1804
rect 2247 1796 2273 1804
rect 2587 1796 2653 1804
rect 2807 1796 2853 1804
rect 3056 1804 3064 1816
rect 3127 1816 3313 1824
rect 3387 1816 3413 1824
rect 3587 1816 3953 1824
rect 4147 1816 4733 1824
rect 4947 1816 4993 1824
rect 2987 1796 3064 1804
rect 3407 1796 3493 1804
rect 4007 1796 4113 1804
rect 4247 1796 4453 1804
rect 4467 1796 4593 1804
rect 4807 1796 4824 1804
rect 516 1776 553 1784
rect 707 1776 804 1784
rect 427 1756 684 1764
rect 227 1736 264 1744
rect 427 1736 473 1744
rect 676 1744 684 1756
rect 727 1756 773 1764
rect 796 1764 804 1776
rect 827 1776 973 1784
rect 1127 1776 1253 1784
rect 1267 1776 1393 1784
rect 1507 1776 1533 1784
rect 1547 1776 1553 1784
rect 1627 1776 1733 1784
rect 2187 1776 2633 1784
rect 2647 1776 2893 1784
rect 2967 1776 3093 1784
rect 3216 1784 3224 1793
rect 3107 1776 3224 1784
rect 3307 1776 3353 1784
rect 3627 1776 3713 1784
rect 3727 1776 3773 1784
rect 3847 1776 3933 1784
rect 3956 1784 3964 1793
rect 4816 1787 4824 1796
rect 4927 1796 4973 1804
rect 5016 1796 5133 1804
rect 5016 1787 5024 1796
rect 5187 1796 5284 1804
rect 5276 1787 5284 1796
rect 5307 1796 5384 1804
rect 5376 1787 5384 1796
rect 5507 1796 5533 1804
rect 5667 1796 5864 1804
rect 3956 1776 3993 1784
rect 4167 1776 4253 1784
rect 4447 1776 4473 1784
rect 4567 1776 4633 1784
rect 5067 1776 5133 1784
rect 5427 1776 5533 1784
rect 796 1756 993 1764
rect 1047 1756 1133 1764
rect 1147 1756 1193 1764
rect 1447 1756 1513 1764
rect 1527 1756 1773 1764
rect 1787 1756 1833 1764
rect 2467 1756 2553 1764
rect 2707 1756 2753 1764
rect 2827 1756 2993 1764
rect 3047 1756 3113 1764
rect 3407 1756 3633 1764
rect 3667 1756 3813 1764
rect 3827 1756 4333 1764
rect 4707 1756 4753 1764
rect 5007 1756 5053 1764
rect 5067 1756 5093 1764
rect 5327 1756 5353 1764
rect 5367 1756 5413 1764
rect 5427 1756 5593 1764
rect 527 1736 664 1744
rect 676 1736 853 1744
rect 267 1716 353 1724
rect 527 1716 553 1724
rect 656 1724 664 1736
rect 967 1736 1053 1744
rect 1367 1736 1413 1744
rect 1507 1736 1813 1744
rect 1947 1736 2573 1744
rect 2727 1736 2913 1744
rect 3087 1736 3293 1744
rect 3487 1736 3653 1744
rect 3787 1736 3953 1744
rect 4347 1736 4533 1744
rect 4547 1736 4773 1744
rect 4787 1736 4913 1744
rect 4927 1736 5233 1744
rect 5247 1736 5433 1744
rect 5447 1736 5573 1744
rect 656 1716 1313 1724
rect 1387 1716 1873 1724
rect 2607 1716 2813 1724
rect 2927 1716 3173 1724
rect 3267 1716 3633 1724
rect 3647 1716 3693 1724
rect 4336 1716 4553 1724
rect 4336 1707 4344 1716
rect 5187 1716 5233 1724
rect 5247 1716 5373 1724
rect 5407 1716 5453 1724
rect 147 1696 733 1704
rect 1867 1696 2233 1704
rect 2407 1696 2473 1704
rect 3427 1696 3473 1704
rect 3487 1696 3893 1704
rect 3987 1696 4093 1704
rect 4467 1696 4553 1704
rect 4627 1696 4813 1704
rect 5256 1696 5433 1704
rect 207 1676 293 1684
rect 1147 1676 1313 1684
rect 1447 1676 1593 1684
rect 1807 1676 1913 1684
rect 1936 1676 1993 1684
rect 947 1656 1093 1664
rect 1936 1664 1944 1676
rect 2527 1676 3193 1684
rect 3276 1676 3313 1684
rect 1107 1656 1944 1664
rect 2907 1656 3213 1664
rect 3247 1656 3264 1664
rect 87 1636 573 1644
rect 587 1636 613 1644
rect 1307 1636 2253 1644
rect 2507 1636 2853 1644
rect 3007 1636 3233 1644
rect 327 1616 373 1624
rect 567 1616 693 1624
rect 747 1616 753 1624
rect 767 1616 893 1624
rect 987 1616 1293 1624
rect 1347 1616 1453 1624
rect 1587 1616 1633 1624
rect 1747 1616 1833 1624
rect 2047 1616 2333 1624
rect 2547 1616 2713 1624
rect 2807 1616 3033 1624
rect 3047 1616 3053 1624
rect 287 1596 384 1604
rect 376 1587 384 1596
rect 887 1596 1033 1604
rect 1167 1596 1373 1604
rect 1607 1596 1633 1604
rect 2307 1596 2413 1604
rect 2607 1596 2724 1604
rect 47 1576 113 1584
rect 287 1576 353 1584
rect 507 1576 533 1584
rect 787 1576 853 1584
rect 927 1576 973 1584
rect 1047 1576 1173 1584
rect 1567 1576 1653 1584
rect 2136 1584 2144 1593
rect 2047 1576 2144 1584
rect 2267 1576 2313 1584
rect 2367 1576 2453 1584
rect -24 1556 13 1564
rect 147 1556 213 1564
rect 256 1564 264 1573
rect 2716 1567 2724 1596
rect 3096 1596 3113 1604
rect 2747 1576 2973 1584
rect 256 1556 393 1564
rect 607 1556 633 1564
rect 1207 1556 1253 1564
rect 1267 1556 1313 1564
rect 1487 1556 1773 1564
rect 3096 1564 3104 1596
rect 3127 1576 3233 1584
rect 3096 1556 3124 1564
rect 96 1544 104 1553
rect 3116 1547 3124 1556
rect 96 1536 113 1544
rect 207 1536 233 1544
rect 367 1536 753 1544
rect 2447 1536 2753 1544
rect 2767 1536 2793 1544
rect 2927 1536 2973 1544
rect 87 1516 373 1524
rect 967 1516 1253 1524
rect 2667 1516 2853 1524
rect 3027 1516 3133 1524
rect 27 1496 1393 1504
rect 3256 1487 3264 1656
rect 3276 1487 3284 1676
rect 3567 1676 3673 1684
rect 4087 1676 4233 1684
rect 4787 1676 5013 1684
rect 5256 1684 5264 1696
rect 5207 1676 5264 1684
rect 5287 1676 5333 1684
rect 3747 1656 3913 1664
rect 4007 1656 4293 1664
rect 4367 1656 4833 1664
rect 5087 1656 5193 1664
rect 5207 1656 5253 1664
rect 5307 1656 5473 1664
rect 3767 1636 4073 1644
rect 4096 1636 4793 1644
rect 3567 1616 3593 1624
rect 3687 1616 3753 1624
rect 4096 1624 4104 1636
rect 5127 1636 5373 1644
rect 5587 1636 5753 1644
rect 3987 1616 4104 1624
rect 4467 1616 4473 1624
rect 4547 1616 4613 1624
rect 4807 1616 4853 1624
rect 4887 1616 4933 1624
rect 5027 1616 5364 1624
rect 3547 1596 3593 1604
rect 3676 1596 3713 1604
rect 3676 1584 3684 1596
rect 3847 1596 3873 1604
rect 4007 1596 4013 1604
rect 4027 1596 4124 1604
rect 3667 1576 3684 1584
rect 3707 1576 3733 1584
rect 3787 1576 3893 1584
rect 3447 1556 3473 1564
rect 3627 1556 3673 1564
rect 4116 1564 4124 1596
rect 4147 1596 4253 1604
rect 4347 1596 4493 1604
rect 4507 1596 4573 1604
rect 4667 1596 4753 1604
rect 4856 1596 4893 1604
rect 4287 1576 4433 1584
rect 4447 1576 4553 1584
rect 4567 1576 4633 1584
rect 4776 1584 4784 1593
rect 4647 1576 4784 1584
rect 4856 1567 4864 1596
rect 5287 1596 5333 1604
rect 5356 1587 5364 1616
rect 5647 1616 5713 1624
rect 5487 1596 5533 1604
rect 5667 1596 5793 1604
rect 5327 1576 5344 1584
rect 5336 1567 5344 1576
rect 5456 1576 5573 1584
rect 5456 1567 5464 1576
rect 5627 1576 5793 1584
rect 4116 1556 4153 1564
rect 4747 1556 4833 1564
rect 5087 1556 5173 1564
rect 5347 1556 5433 1564
rect 5507 1556 5553 1564
rect 5567 1556 5593 1564
rect 3487 1536 3513 1544
rect 3547 1536 3593 1544
rect 3747 1536 4593 1544
rect 4607 1536 4813 1544
rect 4827 1536 5033 1544
rect 5207 1536 5253 1544
rect 5407 1536 5453 1544
rect 5627 1536 5673 1544
rect 3527 1516 3853 1524
rect 3867 1516 4113 1524
rect 4787 1516 4873 1524
rect 4887 1516 4993 1524
rect 5127 1516 5213 1524
rect 5327 1516 5773 1524
rect 3447 1496 4733 1504
rect 5427 1496 5773 1504
rect 307 1476 393 1484
rect 2047 1476 2113 1484
rect 3547 1476 4013 1484
rect 4027 1476 4273 1484
rect 4287 1476 4313 1484
rect 4327 1476 4473 1484
rect 5447 1476 5513 1484
rect 327 1456 353 1464
rect 2547 1456 3453 1464
rect 3467 1456 5033 1464
rect 5047 1456 5073 1464
rect 5087 1456 5333 1464
rect 2307 1436 3533 1444
rect 5187 1436 5233 1444
rect 127 1416 313 1424
rect 1387 1416 2593 1424
rect 2607 1416 2733 1424
rect 2747 1416 2933 1424
rect 3807 1416 3833 1424
rect 3967 1416 4753 1424
rect 5107 1416 5233 1424
rect 2567 1396 2613 1404
rect 2847 1396 2873 1404
rect 3127 1396 3293 1404
rect 3667 1396 3693 1404
rect 3707 1396 4353 1404
rect 4827 1396 4853 1404
rect 5587 1396 5653 1404
rect 1707 1376 1753 1384
rect 1767 1376 1793 1384
rect 1807 1376 2073 1384
rect 2147 1376 2233 1384
rect 2927 1376 3033 1384
rect 3467 1376 3493 1384
rect 3747 1376 3773 1384
rect 3787 1376 4173 1384
rect 4547 1376 4853 1384
rect 5147 1376 5213 1384
rect 5547 1376 5653 1384
rect 827 1356 913 1364
rect 927 1356 1013 1364
rect 1716 1356 1733 1364
rect 1716 1347 1724 1356
rect 1747 1356 1984 1364
rect 1976 1347 1984 1356
rect 2647 1356 2853 1364
rect 2867 1356 2913 1364
rect 3007 1356 3053 1364
rect 3207 1356 3913 1364
rect 4087 1356 4133 1364
rect 5147 1356 5253 1364
rect 5267 1356 5553 1364
rect 5707 1356 5753 1364
rect 207 1336 473 1344
rect 516 1336 533 1344
rect 107 1316 193 1324
rect 247 1316 273 1324
rect 407 1316 493 1324
rect 516 1307 524 1336
rect 887 1336 953 1344
rect 967 1336 1193 1344
rect 1467 1336 1673 1344
rect 1887 1336 1933 1344
rect 2027 1336 2193 1344
rect 2247 1336 2293 1344
rect 2387 1336 4493 1344
rect 4507 1336 4653 1344
rect 4667 1336 4673 1344
rect 4727 1336 5093 1344
rect 5107 1336 5273 1344
rect 5287 1336 5313 1344
rect 5407 1336 5493 1344
rect 5607 1336 5633 1344
rect 547 1316 573 1324
rect 587 1316 673 1324
rect 1067 1316 1133 1324
rect 1187 1316 1213 1324
rect 1567 1316 1693 1324
rect 1707 1316 1953 1324
rect 2067 1316 2253 1324
rect 2407 1316 2673 1324
rect 2747 1316 2873 1324
rect 2887 1316 3013 1324
rect 3027 1316 3153 1324
rect 3707 1316 3764 1324
rect 267 1296 433 1304
rect 567 1296 633 1304
rect 647 1296 793 1304
rect 1167 1296 1293 1304
rect 2227 1296 2353 1304
rect 2567 1296 2613 1304
rect 2716 1287 2724 1313
rect 3756 1307 3764 1316
rect 4107 1316 4153 1324
rect 4567 1316 4593 1324
rect 4647 1316 4733 1324
rect 4907 1316 5113 1324
rect 5267 1316 5353 1324
rect 5376 1316 5493 1324
rect 2787 1296 2813 1304
rect 2847 1296 2893 1304
rect 2987 1296 3033 1304
rect 3147 1296 3413 1304
rect 3467 1296 3533 1304
rect 4056 1304 4064 1313
rect 4196 1304 4204 1313
rect 4056 1296 4293 1304
rect 4316 1304 4324 1313
rect 4316 1296 4453 1304
rect 4527 1296 4573 1304
rect 5376 1304 5384 1316
rect 5027 1296 5384 1304
rect 387 1276 553 1284
rect 1267 1276 1313 1284
rect 2007 1276 2093 1284
rect 2107 1276 2313 1284
rect 2347 1276 2453 1284
rect 2467 1276 2533 1284
rect 2787 1276 2853 1284
rect 3047 1276 3273 1284
rect 3327 1276 3453 1284
rect 3687 1276 3733 1284
rect 4027 1276 4173 1284
rect 4287 1276 4333 1284
rect 4587 1276 4693 1284
rect 4807 1276 4893 1284
rect 4907 1276 5013 1284
rect 5227 1276 5633 1284
rect 187 1256 233 1264
rect 327 1256 373 1264
rect 467 1256 513 1264
rect 547 1256 653 1264
rect 2107 1256 2273 1264
rect 2367 1256 3573 1264
rect 3727 1256 3793 1264
rect 4447 1256 4473 1264
rect 4487 1256 4793 1264
rect 5307 1256 5413 1264
rect 127 1236 273 1244
rect 287 1236 473 1244
rect 1807 1236 2373 1244
rect 3207 1236 3373 1244
rect 4227 1236 4993 1244
rect 147 1216 213 1224
rect 227 1216 533 1224
rect 2527 1216 2733 1224
rect 2807 1216 3173 1224
rect 3427 1216 3493 1224
rect 3827 1216 3893 1224
rect 3907 1216 4433 1224
rect 2327 1196 2693 1204
rect 2767 1196 3433 1204
rect 3487 1196 3633 1204
rect 3647 1196 3713 1204
rect 3787 1196 4213 1204
rect 4427 1196 4873 1204
rect 5607 1196 5633 1204
rect 107 1176 433 1184
rect 1567 1176 1613 1184
rect 1627 1176 2013 1184
rect 2087 1176 2493 1184
rect 2727 1176 2813 1184
rect 2827 1176 2953 1184
rect 2967 1176 2993 1184
rect 3007 1176 3213 1184
rect 3507 1176 3593 1184
rect 3607 1176 3673 1184
rect 3807 1176 3853 1184
rect 4267 1176 4373 1184
rect 4667 1176 4693 1184
rect 5147 1176 5473 1184
rect 5607 1176 5673 1184
rect 227 1156 293 1164
rect 667 1156 773 1164
rect 787 1156 933 1164
rect 1147 1156 1433 1164
rect 1527 1156 1633 1164
rect 3167 1156 3373 1164
rect 3567 1156 4353 1164
rect 4407 1156 4493 1164
rect 4507 1156 4533 1164
rect 4547 1156 4713 1164
rect 5347 1156 5373 1164
rect 5687 1156 5753 1164
rect 47 1136 173 1144
rect 447 1136 613 1144
rect 687 1136 893 1144
rect 947 1136 993 1144
rect 1207 1136 1273 1144
rect 1287 1136 1333 1144
rect 1387 1136 1533 1144
rect 1847 1136 2213 1144
rect 2227 1136 2253 1144
rect 2447 1136 2553 1144
rect 2967 1136 3053 1144
rect 3236 1136 3253 1144
rect 176 1116 353 1124
rect 87 1096 153 1104
rect 176 1104 184 1116
rect 407 1116 613 1124
rect 847 1116 1053 1124
rect 1227 1116 2033 1124
rect 2187 1116 2313 1124
rect 2387 1116 2453 1124
rect 2607 1116 2753 1124
rect 2907 1116 2933 1124
rect 3087 1116 3113 1124
rect 3236 1107 3244 1136
rect 3407 1136 3433 1144
rect 3547 1136 3853 1144
rect 4027 1136 4093 1144
rect 4367 1136 4453 1144
rect 4627 1136 4664 1144
rect 3327 1116 3593 1124
rect 3707 1116 3733 1124
rect 3907 1116 3973 1124
rect 4127 1116 4153 1124
rect 4187 1116 4313 1124
rect 4336 1116 4493 1124
rect 4336 1107 4344 1116
rect 4656 1107 4664 1136
rect 4727 1136 4733 1144
rect 4747 1136 4913 1144
rect 4927 1136 4973 1144
rect 5007 1136 5233 1144
rect 5307 1136 5313 1144
rect 5327 1136 5413 1144
rect 5427 1136 5473 1144
rect 5507 1136 5533 1144
rect 5727 1136 5784 1144
rect 4787 1116 4813 1124
rect 5287 1116 5373 1124
rect 5396 1116 5513 1124
rect 5396 1107 5404 1116
rect 5627 1116 5744 1124
rect 167 1096 184 1104
rect 207 1096 273 1104
rect 296 1096 373 1104
rect 296 1084 304 1096
rect 387 1096 493 1104
rect 787 1096 873 1104
rect 1127 1096 1293 1104
rect 1307 1096 1373 1104
rect 1547 1096 1913 1104
rect 2067 1096 2113 1104
rect 2287 1096 2333 1104
rect 2367 1096 2393 1104
rect 2487 1096 2533 1104
rect 2647 1096 2673 1104
rect 2747 1096 2773 1104
rect 3627 1096 3653 1104
rect 3927 1096 3973 1104
rect 4467 1096 4513 1104
rect 4687 1096 4713 1104
rect 5687 1096 5693 1104
rect 5707 1096 5713 1104
rect 5736 1104 5744 1116
rect 5776 1107 5784 1136
rect 5736 1096 5753 1104
rect 87 1076 304 1084
rect 327 1076 453 1084
rect 547 1076 593 1084
rect 647 1076 673 1084
rect 707 1076 893 1084
rect 1036 1084 1044 1093
rect 1036 1076 1253 1084
rect 1267 1076 1413 1084
rect 1467 1076 1753 1084
rect 1887 1076 1933 1084
rect 2016 1084 2024 1093
rect 1967 1076 2153 1084
rect 2207 1076 2613 1084
rect 2627 1076 2973 1084
rect 3107 1076 3153 1084
rect 3576 1084 3584 1093
rect 3576 1076 3593 1084
rect 3607 1076 3693 1084
rect 3807 1076 3833 1084
rect 3887 1076 4413 1084
rect 4707 1076 4753 1084
rect 4787 1076 4813 1084
rect 4867 1076 4913 1084
rect 4927 1076 4953 1084
rect 5587 1076 5653 1084
rect 1267 1056 1493 1064
rect 1867 1056 1893 1064
rect 2087 1056 3133 1064
rect 3287 1056 4053 1064
rect 4067 1056 5013 1064
rect 1307 1036 1353 1044
rect 2427 1036 2513 1044
rect 2887 1036 3333 1044
rect 3667 1036 3753 1044
rect 367 1016 393 1024
rect 427 1016 633 1024
rect 647 1016 673 1024
rect 3447 1016 3913 1024
rect 1827 996 3513 1004
rect 2927 976 3493 984
rect 3507 976 3693 984
rect 487 956 513 964
rect 3516 956 5013 964
rect 3516 944 3524 956
rect 5027 956 5053 964
rect 2987 936 3524 944
rect 3807 936 3853 944
rect 2247 916 2293 924
rect 3267 916 3533 924
rect 3667 916 4213 924
rect 5507 916 5533 924
rect 587 896 613 904
rect 627 896 733 904
rect 2147 896 2213 904
rect 2307 896 2553 904
rect 3827 896 3873 904
rect 3896 896 3993 904
rect 147 876 173 884
rect 887 876 1213 884
rect 1347 876 1364 884
rect 96 856 233 864
rect 96 847 104 856
rect 447 856 553 864
rect 687 856 713 864
rect 727 856 793 864
rect 916 856 1133 864
rect 916 847 924 856
rect 1356 864 1364 876
rect 1447 876 1853 884
rect 2016 876 2273 884
rect 1356 856 1373 864
rect 1427 856 1453 864
rect 1487 856 1553 864
rect 1647 856 1713 864
rect 2016 864 2024 876
rect 2947 876 3113 884
rect 3896 884 3904 896
rect 4007 896 4233 904
rect 5047 896 5133 904
rect 5427 896 5613 904
rect 3127 876 3904 884
rect 4107 876 4133 884
rect 4607 876 4793 884
rect 4887 876 4933 884
rect 5247 876 5313 884
rect 5547 876 5684 884
rect 1907 856 2024 864
rect 2047 856 2053 864
rect 2067 856 2133 864
rect 2527 856 2633 864
rect 2867 856 2893 864
rect 3307 856 3473 864
rect 3727 856 3893 864
rect 4047 856 4113 864
rect 4127 856 4153 864
rect 4627 856 4653 864
rect 4667 856 4773 864
rect 4907 856 5613 864
rect 5627 856 5653 864
rect 5676 864 5684 876
rect 5707 876 5753 884
rect 5676 856 5724 864
rect 147 836 193 844
rect 387 836 513 844
rect 567 836 853 844
rect 967 836 1013 844
rect 1087 836 1133 844
rect 1367 836 1573 844
rect 1787 836 1833 844
rect 1847 836 1913 844
rect 1927 836 1973 844
rect 2587 836 2773 844
rect 3027 836 3053 844
rect 3147 836 3173 844
rect 3427 836 3473 844
rect 3687 836 3733 844
rect 3807 836 3833 844
rect 3927 836 4013 844
rect 4187 836 4313 844
rect 4407 836 4433 844
rect 4527 836 4573 844
rect 4707 836 4733 844
rect 4756 836 4893 844
rect 267 816 313 824
rect 507 816 613 824
rect 827 816 893 824
rect 1196 824 1204 833
rect 1027 816 1204 824
rect 1227 816 1293 824
rect 1747 816 1813 824
rect 1887 816 2013 824
rect 2027 816 2073 824
rect 2167 816 2433 824
rect 2687 816 2733 824
rect 3407 816 3444 824
rect 127 796 213 804
rect 247 796 273 804
rect 347 796 373 804
rect 407 796 533 804
rect 547 796 933 804
rect 1107 796 1233 804
rect 1467 796 1613 804
rect 1787 796 2113 804
rect 2127 796 2313 804
rect 2967 796 2993 804
rect 3127 796 3153 804
rect 3347 796 3413 804
rect 3436 804 3444 816
rect 3527 816 3893 824
rect 4207 816 4253 824
rect 4756 824 4764 836
rect 4907 836 4933 844
rect 4987 836 5073 844
rect 4547 816 4764 824
rect 4967 816 5033 824
rect 3436 796 3533 804
rect 3567 796 3673 804
rect 3687 796 3753 804
rect 3807 796 3993 804
rect 4007 796 4053 804
rect 4147 796 4293 804
rect 4307 796 4413 804
rect 4567 796 4733 804
rect 4787 796 4813 804
rect 5056 804 5064 836
rect 5327 836 5373 844
rect 5396 836 5493 844
rect 5267 816 5313 824
rect 5396 807 5404 836
rect 5587 836 5693 844
rect 5427 816 5473 824
rect 5567 816 5593 824
rect 5716 824 5724 856
rect 5687 816 5724 824
rect 4827 796 5073 804
rect 5127 796 5253 804
rect 5287 796 5333 804
rect 667 776 733 784
rect 747 776 953 784
rect 1767 776 1993 784
rect 2707 776 2813 784
rect 2827 776 3273 784
rect 3447 776 4073 784
rect 4867 776 4913 784
rect 4927 776 5113 784
rect 5307 776 5493 784
rect 687 756 773 764
rect 787 756 1033 764
rect 1987 756 2093 764
rect 2447 756 2653 764
rect 3867 756 4333 764
rect 4347 756 4773 764
rect 1347 736 1953 744
rect 2007 736 4513 744
rect 4527 736 4673 744
rect 5267 736 5433 744
rect 5447 736 5473 744
rect 5487 736 5653 744
rect 147 716 353 724
rect 3807 716 3893 724
rect 5347 716 5673 724
rect 1467 696 1813 704
rect 1867 696 2373 704
rect 3887 696 4033 704
rect 4047 696 4433 704
rect 4867 696 5353 704
rect 5367 696 5373 704
rect 5447 696 5593 704
rect 947 676 1113 684
rect 1127 676 1213 684
rect 1227 676 1533 684
rect 1827 676 2173 684
rect 3567 676 4353 684
rect 4367 676 4593 684
rect 4727 676 4833 684
rect 4847 676 4993 684
rect 5167 676 5213 684
rect 5287 676 5553 684
rect 167 656 273 664
rect 467 656 653 664
rect 987 656 993 664
rect 1007 656 1184 664
rect 127 636 533 644
rect 296 627 304 636
rect 1107 636 1153 644
rect 1176 644 1184 656
rect 1407 656 1513 664
rect 1667 656 1933 664
rect 2007 656 2093 664
rect 2127 656 2253 664
rect 2747 656 2844 664
rect 1176 636 1353 644
rect 1236 627 1244 636
rect 1527 636 1673 644
rect 1727 636 1733 644
rect 1747 636 1993 644
rect 2087 636 2233 644
rect 2247 636 2273 644
rect 2836 627 2844 656
rect 2887 656 3093 664
rect 3107 656 3193 664
rect 3207 656 3373 664
rect 3427 656 3633 664
rect 3827 656 3933 664
rect 4187 656 4213 664
rect 4387 656 4473 664
rect 4667 656 4793 664
rect 4887 656 4913 664
rect 4927 656 4953 664
rect 5107 656 5133 664
rect 5167 656 5453 664
rect 5467 656 5633 664
rect 3047 636 3133 644
rect 3167 636 3513 644
rect 3567 636 3593 644
rect 3687 636 3773 644
rect 4087 636 4204 644
rect 67 616 93 624
rect 107 616 253 624
rect 327 616 393 624
rect 607 616 673 624
rect 696 616 793 624
rect 47 596 73 604
rect 516 604 524 613
rect 427 596 633 604
rect 696 604 704 616
rect 987 616 1013 624
rect 1147 616 1193 624
rect 1427 616 1533 624
rect 1607 616 1653 624
rect 1707 616 1773 624
rect 1867 616 1913 624
rect 1967 616 1993 624
rect 2356 616 2473 624
rect 2356 607 2364 616
rect 2627 616 2733 624
rect 2747 616 2824 624
rect 647 596 704 604
rect 867 596 1073 604
rect 1207 596 1553 604
rect 1727 596 1833 604
rect 1847 596 2053 604
rect 2816 604 2824 616
rect 3007 616 3073 624
rect 3127 616 3173 624
rect 3307 616 3333 624
rect 3347 616 3493 624
rect 3616 624 3624 633
rect 3547 616 3664 624
rect 2816 596 2973 604
rect 3027 596 3233 604
rect 3256 604 3264 613
rect 3256 596 3353 604
rect 87 576 153 584
rect 687 576 773 584
rect 787 576 1313 584
rect 1427 576 1793 584
rect 2187 576 2793 584
rect 2807 576 3093 584
rect 3496 584 3504 613
rect 3656 607 3664 616
rect 3707 616 3793 624
rect 3807 616 3893 624
rect 3916 604 3924 633
rect 4196 627 4204 636
rect 4647 636 4713 644
rect 4787 636 4853 644
rect 5147 636 5273 644
rect 5296 636 5413 644
rect 4007 616 4053 624
rect 4216 607 4224 633
rect 4247 616 4333 624
rect 4407 616 4453 624
rect 4627 616 4653 624
rect 4736 624 4744 633
rect 4676 616 4744 624
rect 3747 596 3924 604
rect 4576 604 4584 613
rect 4676 604 4684 616
rect 4767 616 4793 624
rect 4847 616 4873 624
rect 4236 596 4684 604
rect 4236 584 4244 596
rect 4896 604 4904 633
rect 5296 624 5304 636
rect 5427 636 5533 644
rect 5607 636 5693 644
rect 5267 616 5304 624
rect 5407 616 5473 624
rect 5487 616 5573 624
rect 4827 596 4904 604
rect 5307 596 5333 604
rect 5667 596 5733 604
rect 3496 576 4244 584
rect 1247 556 1373 564
rect 1387 556 1473 564
rect 1847 556 2493 564
rect 3267 556 3353 564
rect 3367 556 4213 564
rect 167 536 453 544
rect 467 536 513 544
rect 1127 536 1153 544
rect 2347 536 2593 544
rect 2607 536 2693 544
rect 2707 536 2973 544
rect 2987 536 3153 544
rect 3927 536 3953 544
rect 5507 536 5673 544
rect 2647 516 2773 524
rect 2787 516 2793 524
rect 3827 516 4013 524
rect 5227 516 5393 524
rect 2087 496 2293 504
rect 4807 496 5513 504
rect 5107 476 5413 484
rect 5427 476 5593 484
rect 2667 456 2913 464
rect 3187 456 3693 464
rect 4507 456 4533 464
rect 5267 456 5353 464
rect 2607 436 3493 444
rect 4127 436 4193 444
rect 5167 436 5613 444
rect 307 416 553 424
rect 1027 416 1633 424
rect 2267 416 2533 424
rect 2847 416 3133 424
rect 3147 416 3313 424
rect 3867 416 3893 424
rect 5147 416 5353 424
rect 747 396 813 404
rect 1487 396 1913 404
rect 2367 396 2633 404
rect 2727 396 3053 404
rect 3227 396 3413 404
rect 3507 396 3573 404
rect 3607 396 3733 404
rect 3807 396 3833 404
rect 4136 396 4153 404
rect 4136 387 4144 396
rect 4187 396 4513 404
rect 5087 396 5293 404
rect 5387 396 5513 404
rect 5527 396 5553 404
rect 5567 396 5633 404
rect 5727 396 5753 404
rect 216 376 413 384
rect 216 367 224 376
rect 556 376 793 384
rect 107 356 213 364
rect 267 356 293 364
rect 467 356 533 364
rect 556 364 564 376
rect 967 376 1033 384
rect 1047 376 1073 384
rect 1116 376 1353 384
rect 547 356 564 364
rect 1007 356 1093 364
rect 1116 364 1124 376
rect 1407 376 1513 384
rect 1527 376 1593 384
rect 1667 376 1693 384
rect 1787 376 1853 384
rect 1867 376 1993 384
rect 2007 376 2553 384
rect 2567 376 2873 384
rect 2887 376 3533 384
rect 3547 376 3673 384
rect 3867 376 3933 384
rect 3947 376 4093 384
rect 4147 376 4413 384
rect 4527 376 4813 384
rect 5027 376 5144 384
rect 5136 367 5144 376
rect 5187 376 5433 384
rect 5627 376 5644 384
rect 1107 356 1124 364
rect 1387 356 1453 364
rect 1627 356 1713 364
rect 2047 356 2133 364
rect 2227 356 2293 364
rect 2307 356 2413 364
rect 2547 356 2733 364
rect 3027 356 3153 364
rect 3187 356 3253 364
rect 3467 356 3633 364
rect 3927 356 3953 364
rect 4027 356 4113 364
rect 4207 356 4244 364
rect 127 336 313 344
rect 327 336 373 344
rect 416 344 424 353
rect 416 336 653 344
rect 976 344 984 353
rect 947 336 984 344
rect 1267 336 1333 344
rect 1687 336 1733 344
rect 1827 336 1913 344
rect 1927 336 2273 344
rect 2467 336 2673 344
rect 2707 336 2753 344
rect 2887 336 2933 344
rect 3727 336 3833 344
rect 3887 336 3993 344
rect 4007 336 4213 344
rect 4236 344 4244 356
rect 4387 356 4484 364
rect 4236 336 4253 344
rect 267 316 293 324
rect 307 316 433 324
rect 1547 316 1613 324
rect 2327 316 2353 324
rect 2447 316 2573 324
rect 2847 316 2893 324
rect 2927 316 2993 324
rect 3167 316 3273 324
rect 3287 316 3333 324
rect 4276 324 4284 353
rect 4476 344 4484 356
rect 4507 356 4533 364
rect 4587 356 4633 364
rect 4687 356 4733 364
rect 4896 356 4953 364
rect 4896 347 4904 356
rect 5156 364 5164 373
rect 5636 367 5644 376
rect 5156 356 5173 364
rect 5247 356 5333 364
rect 5747 356 5793 364
rect 4476 336 4593 344
rect 5047 336 5153 344
rect 5207 336 5373 344
rect 5476 344 5484 353
rect 5476 336 5613 344
rect 4187 316 4284 324
rect 4327 316 4613 324
rect 4767 316 4813 324
rect 4987 316 5133 324
rect 5427 316 5493 324
rect 347 296 393 304
rect 987 296 1053 304
rect 1067 296 1633 304
rect 2387 296 2633 304
rect 3447 296 3673 304
rect 3687 296 4233 304
rect 4247 296 4413 304
rect 827 276 1073 284
rect 1087 276 1193 284
rect 4187 276 4573 284
rect 287 256 373 264
rect 387 256 593 264
rect 4027 256 4453 264
rect 487 236 573 244
rect 4647 236 4853 244
rect 5207 236 5353 244
rect 527 216 833 224
rect 847 216 913 224
rect 927 216 1013 224
rect 4607 216 4693 224
rect 4707 216 4953 224
rect 4967 216 5313 224
rect 427 196 553 204
rect 567 196 673 204
rect 867 196 1133 204
rect 1607 196 2173 204
rect 2527 196 2713 204
rect 3327 196 3373 204
rect 3387 196 3553 204
rect 4067 196 4133 204
rect 4147 196 4333 204
rect 4347 196 4993 204
rect 5016 196 5093 204
rect 167 176 213 184
rect 227 176 533 184
rect 587 176 633 184
rect 647 176 873 184
rect 907 176 1173 184
rect 1247 176 1313 184
rect 1347 176 1433 184
rect 1747 176 1893 184
rect 2187 176 2253 184
rect 2667 176 3033 184
rect 3207 176 3553 184
rect 3567 176 3733 184
rect 5016 184 5024 196
rect 5227 196 5333 204
rect 4767 176 5024 184
rect 5047 176 5073 184
rect 5087 176 5453 184
rect 5627 176 5673 184
rect 5687 176 5733 184
rect 107 156 173 164
rect 656 156 953 164
rect 656 147 664 156
rect 1287 156 1293 164
rect 1307 156 1413 164
rect 1707 156 1793 164
rect 1807 156 1913 164
rect 2127 156 2153 164
rect 2167 156 2333 164
rect 2347 156 2453 164
rect 2476 156 2613 164
rect 96 136 113 144
rect 96 124 104 136
rect 147 136 193 144
rect 407 136 473 144
rect 567 136 653 144
rect 707 136 833 144
rect 887 136 1193 144
rect 1207 136 1233 144
rect 1587 136 1673 144
rect 1727 136 1753 144
rect 2476 144 2484 156
rect 2636 156 2913 164
rect 2636 147 2644 156
rect 2936 156 3413 164
rect 1967 136 2484 144
rect 2687 136 2713 144
rect 2936 144 2944 156
rect 3867 156 4073 164
rect 4107 156 4113 164
rect 4127 156 4293 164
rect 4307 156 4713 164
rect 4887 156 4973 164
rect 5027 156 5113 164
rect 5127 156 5233 164
rect 5247 156 5293 164
rect 2847 136 2944 144
rect 2936 127 2944 136
rect 3067 136 3173 144
rect 3227 136 3293 144
rect 3347 136 3393 144
rect 3447 136 3533 144
rect 3676 136 4013 144
rect 3676 127 3684 136
rect 4467 136 4553 144
rect 4567 136 4604 144
rect 87 116 104 124
rect 127 116 153 124
rect 187 116 233 124
rect 847 116 893 124
rect 907 116 933 124
rect 967 116 1033 124
rect 1047 116 1493 124
rect 1987 116 2073 124
rect 2147 116 2393 124
rect 2407 116 2473 124
rect 3007 116 3073 124
rect 4007 116 4093 124
rect 4407 116 4513 124
rect 4596 124 4604 136
rect 4627 136 4833 144
rect 5007 136 5033 144
rect 5056 136 5233 144
rect 5056 124 5064 136
rect 5367 136 5493 144
rect 5607 136 5653 144
rect 4596 116 5064 124
rect 5267 116 5373 124
rect 5447 116 5673 124
rect 207 96 793 104
rect 1936 104 1944 113
rect 1867 96 2093 104
rect 2787 96 2893 104
rect 2907 96 3153 104
rect 3647 96 4533 104
rect 4576 104 4584 113
rect 4576 96 4633 104
rect 2287 36 2673 44
rect 2647 16 2953 24
<< m1p >>
rect 4 5762 5816 5778
rect 44 5522 156 5538
rect 184 5522 316 5538
rect 344 5522 456 5538
rect 484 5522 596 5538
rect 624 5522 756 5538
rect 764 5522 1036 5538
rect 1044 5522 1176 5538
rect 1184 5522 1316 5538
rect 1324 5522 1456 5538
rect 1464 5522 1596 5538
rect 1624 5522 1736 5538
rect 1764 5522 1876 5538
rect 1904 5522 2136 5538
rect 2144 5522 2256 5538
rect 2284 5522 2396 5538
rect 2424 5522 2536 5538
rect 2544 5522 3196 5538
rect 3204 5522 3616 5538
rect 3624 5522 3896 5538
rect 3924 5522 4036 5538
rect 4044 5522 4416 5538
rect 4424 5522 5396 5538
rect 5424 5522 5796 5538
rect 4 5282 5816 5298
rect 44 5042 156 5058
rect 184 5042 296 5058
rect 324 5042 696 5058
rect 704 5042 836 5058
rect 844 5042 976 5058
rect 984 5042 1116 5058
rect 1124 5042 1356 5058
rect 1384 5042 1496 5058
rect 1524 5042 1776 5058
rect 1784 5042 2816 5058
rect 2824 5042 2936 5058
rect 2944 5042 3076 5058
rect 3084 5042 3196 5058
rect 3224 5042 3336 5058
rect 3344 5042 3476 5058
rect 3484 5042 3616 5058
rect 3624 5042 3736 5058
rect 3744 5042 3876 5058
rect 3884 5042 3976 5058
rect 4004 5042 4116 5058
rect 4144 5042 4256 5058
rect 4284 5042 4416 5058
rect 4444 5042 4676 5058
rect 4684 5042 5556 5058
rect 5564 5042 5676 5058
rect 5684 5042 5816 5058
rect 4 4802 5816 4818
rect 44 4562 156 4578
rect 184 4562 296 4578
rect 324 4562 436 4578
rect 464 4562 736 4578
rect 744 4562 856 4578
rect 864 4562 976 4578
rect 984 4562 1076 4578
rect 1084 4562 1456 4578
rect 1464 4562 2696 4578
rect 2704 4562 3276 4578
rect 3284 4562 3416 4578
rect 3424 4562 3556 4578
rect 3564 4562 3696 4578
rect 3704 4562 3836 4578
rect 3844 4562 3956 4578
rect 3984 4562 4096 4578
rect 4104 4562 4216 4578
rect 4224 4562 4336 4578
rect 4364 4562 4496 4578
rect 4504 4562 5616 4578
rect 5624 4562 5756 4578
rect 4 4322 5816 4338
rect 44 4082 776 4098
rect 784 4082 916 4098
rect 924 4082 1016 4098
rect 1024 4082 1156 4098
rect 1184 4082 1316 4098
rect 1324 4082 1556 4098
rect 1564 4082 1676 4098
rect 1684 4082 1796 4098
rect 1804 4082 1936 4098
rect 1944 4082 2076 4098
rect 2104 4082 2216 4098
rect 2244 4082 2356 4098
rect 2384 4082 2496 4098
rect 2524 4082 2756 4098
rect 2764 4082 3036 4098
rect 3044 4082 3496 4098
rect 3504 4082 4836 4098
rect 4844 4082 5076 4098
rect 5084 4082 5816 4098
rect 4 3842 5816 3858
rect 44 3602 156 3618
rect 164 3602 296 3618
rect 304 3602 936 3618
rect 944 3602 1076 3618
rect 1104 3602 1216 3618
rect 1224 3602 1336 3618
rect 1364 3602 1476 3618
rect 1504 3602 1616 3618
rect 1644 3602 2216 3618
rect 2224 3602 2356 3618
rect 2364 3602 2496 3618
rect 2504 3602 2616 3618
rect 2644 3602 2756 3618
rect 2764 3602 2876 3618
rect 2884 3602 3016 3618
rect 3024 3602 3136 3618
rect 3164 3602 3276 3618
rect 3284 3602 3716 3618
rect 3724 3602 3856 3618
rect 3864 3602 3956 3618
rect 3984 3602 4476 3618
rect 4484 3602 4836 3618
rect 4864 3602 4956 3618
rect 4984 3602 5096 3618
rect 5104 3602 5776 3618
rect 4 3362 5816 3378
rect 44 3122 356 3138
rect 364 3122 476 3138
rect 484 3122 616 3138
rect 624 3122 756 3138
rect 764 3122 896 3138
rect 904 3122 1036 3138
rect 1044 3122 1176 3138
rect 1184 3122 1416 3138
rect 1444 3122 1556 3138
rect 1584 3122 1716 3138
rect 1724 3122 1856 3138
rect 1884 3122 1996 3138
rect 2004 3122 2776 3138
rect 2784 3122 2916 3138
rect 2924 3122 3056 3138
rect 3064 3122 3176 3138
rect 3184 3122 3316 3138
rect 3324 3122 3436 3138
rect 3444 3122 3576 3138
rect 3584 3122 3716 3138
rect 3724 3122 3856 3138
rect 3864 3122 4696 3138
rect 4704 3122 4836 3138
rect 4844 3122 4956 3138
rect 4964 3122 5316 3138
rect 5324 3122 5776 3138
rect 4 2882 5816 2898
rect 44 2642 136 2658
rect 144 2642 376 2658
rect 384 2642 516 2658
rect 524 2642 896 2658
rect 904 2642 1036 2658
rect 1044 2642 1156 2658
rect 1184 2642 5776 2658
rect 4 2402 5816 2418
rect 44 2162 156 2178
rect 164 2162 556 2178
rect 564 2162 696 2178
rect 724 2162 836 2178
rect 864 2162 976 2178
rect 984 2162 2816 2178
rect 2844 2162 2956 2178
rect 2984 2162 3076 2178
rect 3104 2162 3216 2178
rect 3244 2162 3356 2178
rect 3364 2162 3476 2178
rect 3504 2162 3636 2178
rect 3664 2162 3756 2178
rect 3784 2162 4996 2178
rect 5004 2162 5796 2178
rect 4 1922 5816 1938
rect 44 1682 176 1698
rect 184 1682 316 1698
rect 324 1682 456 1698
rect 464 1682 596 1698
rect 624 1682 716 1698
rect 744 1682 976 1698
rect 984 1682 1376 1698
rect 1384 1682 1516 1698
rect 1524 1682 2656 1698
rect 2684 1682 2776 1698
rect 2804 1682 2916 1698
rect 2944 1682 4716 1698
rect 4724 1682 4836 1698
rect 4844 1682 4956 1698
rect 4984 1682 5116 1698
rect 5144 1682 5796 1698
rect 4 1442 5816 1458
rect 44 1202 996 1218
rect 1004 1202 1116 1218
rect 1124 1202 1236 1218
rect 1244 1202 1356 1218
rect 1384 1202 1476 1218
rect 1484 1202 1596 1218
rect 1624 1202 2116 1218
rect 2124 1202 2516 1218
rect 2544 1202 2676 1218
rect 2704 1202 3436 1218
rect 3444 1202 4256 1218
rect 4264 1202 4396 1218
rect 4404 1202 4556 1218
rect 4564 1202 4696 1218
rect 4704 1202 4956 1218
rect 4964 1202 5056 1218
rect 5084 1202 5176 1218
rect 5184 1202 5296 1218
rect 5324 1202 5436 1218
rect 5464 1202 5576 1218
rect 5584 1202 5796 1218
rect 4 962 5816 978
rect 44 722 156 738
rect 184 722 316 738
rect 324 722 456 738
rect 464 722 596 738
rect 604 722 736 738
rect 744 722 856 738
rect 884 722 1016 738
rect 1024 722 1156 738
rect 1164 722 1296 738
rect 1304 722 1436 738
rect 1444 722 3176 738
rect 3204 722 3316 738
rect 3344 722 3456 738
rect 3464 722 3576 738
rect 3604 722 3716 738
rect 3724 722 3836 738
rect 3844 722 3976 738
rect 3984 722 4376 738
rect 4404 722 5336 738
rect 5344 722 5616 738
rect 5624 722 5736 738
rect 4 482 5816 498
rect 44 242 156 258
rect 184 242 296 258
rect 344 242 456 258
rect 484 242 596 258
rect 624 242 736 258
rect 764 242 876 258
rect 904 242 2836 258
rect 2864 242 2976 258
rect 2984 242 3236 258
rect 3244 242 3356 258
rect 3364 242 3476 258
rect 3504 242 4056 258
rect 4064 242 4776 258
rect 4804 242 4916 258
rect 4924 242 5536 258
rect 5564 242 5796 258
rect 4 2 5816 18
<< m2p >>
rect 513 5653 527 5667
rect 553 5653 567 5667
rect 793 5653 807 5667
rect 833 5653 847 5667
rect 1373 5653 1387 5667
rect 1493 5653 1507 5667
rect 1533 5653 1547 5667
rect 1793 5653 1807 5667
rect 1833 5653 1847 5667
rect 2453 5653 2467 5667
rect 2493 5653 2507 5667
rect 2573 5653 2587 5667
rect 2613 5653 2627 5667
rect 2713 5653 2727 5667
rect 2753 5653 2767 5667
rect 2833 5653 2847 5667
rect 2873 5653 2887 5667
rect 3253 5653 3267 5667
rect 3493 5653 3507 5667
rect 3533 5653 3547 5667
rect 5073 5653 5087 5667
rect 5113 5653 5127 5667
rect 5173 5653 5187 5667
rect 5213 5653 5227 5667
rect 5533 5653 5547 5667
rect 5573 5653 5587 5667
rect 73 5633 87 5647
rect 113 5633 127 5647
rect 213 5633 227 5647
rect 253 5633 267 5647
rect 393 5633 407 5647
rect 433 5633 447 5647
rect 493 5633 507 5647
rect 533 5633 547 5647
rect 653 5633 667 5647
rect 693 5633 707 5647
rect 813 5633 827 5647
rect 933 5633 947 5647
rect 973 5633 987 5647
rect 1213 5633 1227 5647
rect 1513 5633 1527 5647
rect 1553 5633 1567 5647
rect 1673 5633 1687 5647
rect 1713 5633 1727 5647
rect 1813 5633 1827 5647
rect 1853 5633 1867 5647
rect 1933 5633 1947 5647
rect 2033 5633 2047 5647
rect 2073 5633 2087 5647
rect 2173 5633 2187 5647
rect 2213 5633 2227 5647
rect 2293 5633 2307 5647
rect 2333 5633 2347 5647
rect 2473 5633 2487 5647
rect 2593 5633 2607 5647
rect 2633 5633 2647 5647
rect 2733 5633 2747 5647
rect 2773 5633 2787 5647
rect 2853 5633 2867 5647
rect 2973 5633 2987 5647
rect 3073 5633 3087 5647
rect 3113 5633 3127 5647
rect 3513 5633 3527 5647
rect 3553 5633 3567 5647
rect 3653 5633 3667 5647
rect 3753 5633 3767 5647
rect 3853 5633 3867 5647
rect 3953 5633 3967 5647
rect 3993 5633 4007 5647
rect 4093 5633 4107 5647
rect 4453 5633 4467 5647
rect 4493 5633 4507 5647
rect 4593 5633 4607 5647
rect 4733 5633 4747 5647
rect 4833 5633 4847 5647
rect 4933 5633 4947 5647
rect 4973 5633 4987 5647
rect 5093 5633 5107 5647
rect 5193 5633 5207 5647
rect 5313 5633 5327 5647
rect 5353 5633 5367 5647
rect 5453 5633 5467 5647
rect 5553 5633 5567 5647
rect 5673 5633 5687 5647
rect 93 5613 107 5627
rect 133 5613 147 5627
rect 193 5613 207 5627
rect 233 5613 247 5627
rect 373 5613 387 5627
rect 673 5613 687 5627
rect 713 5613 727 5627
rect 913 5613 927 5627
rect 1053 5613 1067 5627
rect 1093 5613 1107 5627
rect 1253 5613 1267 5627
rect 1353 5613 1367 5627
rect 1413 5613 1427 5627
rect 1653 5613 1667 5627
rect 2053 5613 2067 5627
rect 2093 5613 2107 5627
rect 2153 5613 2167 5627
rect 2193 5613 2207 5627
rect 2353 5613 2367 5627
rect 3093 5613 3107 5627
rect 3133 5613 3147 5627
rect 3233 5613 3247 5627
rect 3293 5613 3307 5627
rect 3373 5613 3387 5627
rect 3413 5613 3427 5627
rect 3933 5613 3947 5627
rect 3973 5613 3987 5627
rect 4153 5613 4167 5627
rect 4233 5613 4247 5627
rect 4273 5613 4287 5627
rect 4473 5613 4487 5627
rect 4513 5613 4527 5627
rect 4953 5613 4967 5627
rect 4993 5613 5007 5627
rect 5293 5613 5307 5627
rect 5333 5613 5347 5627
rect 413 5593 427 5607
rect 953 5593 967 5607
rect 1073 5593 1087 5607
rect 1273 5593 1287 5607
rect 1693 5593 1707 5607
rect 1913 5593 1927 5607
rect 2313 5593 2327 5607
rect 2993 5593 3007 5607
rect 3393 5593 3407 5607
rect 3673 5593 3687 5607
rect 3773 5593 3787 5607
rect 3833 5593 3847 5607
rect 4073 5593 4087 5607
rect 4853 5593 4867 5607
rect 5433 5593 5447 5607
rect 5653 5593 5667 5607
rect 1133 5453 1147 5467
rect 1393 5453 1407 5467
rect 2233 5453 2247 5467
rect 3013 5453 3027 5467
rect 3513 5453 3527 5467
rect 3853 5453 3867 5467
rect 4493 5453 4507 5467
rect 4613 5453 4627 5467
rect 5093 5453 5107 5467
rect 93 5433 107 5447
rect 133 5433 147 5447
rect 793 5433 807 5447
rect 833 5433 847 5447
rect 1093 5433 1107 5447
rect 1373 5433 1387 5447
rect 1413 5433 1427 5447
rect 1633 5433 1647 5447
rect 1673 5433 1687 5447
rect 2313 5433 2327 5447
rect 2373 5433 2387 5447
rect 2433 5433 2447 5447
rect 2473 5433 2487 5447
rect 2873 5433 2887 5447
rect 2913 5433 2927 5447
rect 3533 5433 3547 5447
rect 3813 5433 3827 5447
rect 4093 5433 4107 5447
rect 4133 5433 4147 5447
rect 4533 5433 4547 5447
rect 4713 5433 4727 5447
rect 4753 5433 4767 5447
rect 4833 5433 4847 5447
rect 4913 5433 4927 5447
rect 4953 5433 4967 5447
rect 5173 5433 5187 5447
rect 5253 5433 5267 5447
rect 5293 5433 5307 5447
rect 5433 5433 5447 5447
rect 5473 5433 5487 5447
rect 73 5413 87 5427
rect 113 5413 127 5427
rect 253 5413 267 5427
rect 293 5413 307 5427
rect 393 5413 407 5427
rect 433 5413 447 5427
rect 533 5413 547 5427
rect 573 5413 587 5427
rect 653 5413 667 5427
rect 693 5413 707 5427
rect 813 5413 827 5427
rect 853 5413 867 5427
rect 933 5413 947 5427
rect 973 5413 987 5427
rect 1113 5413 1127 5427
rect 1153 5413 1167 5427
rect 1213 5413 1227 5427
rect 1253 5413 1267 5427
rect 1533 5413 1547 5427
rect 1573 5413 1587 5427
rect 1653 5413 1667 5427
rect 1693 5413 1707 5427
rect 1813 5413 1827 5427
rect 1853 5413 1867 5427
rect 1953 5413 1967 5427
rect 1993 5413 2007 5427
rect 2073 5413 2087 5427
rect 2213 5413 2227 5427
rect 2453 5413 2467 5427
rect 2493 5413 2507 5427
rect 2633 5413 2647 5427
rect 2673 5413 2687 5427
rect 2773 5413 2787 5427
rect 2813 5413 2827 5427
rect 2893 5413 2907 5427
rect 2933 5413 2947 5427
rect 3033 5413 3047 5427
rect 3133 5413 3147 5427
rect 3253 5413 3267 5427
rect 3293 5413 3307 5427
rect 3413 5413 3427 5427
rect 3573 5413 3587 5427
rect 3693 5413 3707 5427
rect 3733 5413 3747 5427
rect 3833 5413 3847 5427
rect 3873 5413 3887 5427
rect 3953 5413 3967 5427
rect 4073 5413 4087 5427
rect 4113 5413 4127 5427
rect 4233 5413 4247 5427
rect 4353 5413 4367 5427
rect 4393 5413 4407 5427
rect 4473 5413 4487 5427
rect 4513 5413 4527 5427
rect 4633 5413 4647 5427
rect 4733 5413 4747 5427
rect 4773 5413 4787 5427
rect 5113 5413 5127 5427
rect 5453 5413 5467 5427
rect 5493 5413 5507 5427
rect 5613 5413 5627 5427
rect 5733 5413 5747 5427
rect 233 5393 247 5407
rect 273 5393 287 5407
rect 373 5393 387 5407
rect 413 5393 427 5407
rect 513 5393 527 5407
rect 553 5393 567 5407
rect 673 5393 687 5407
rect 713 5393 727 5407
rect 953 5393 967 5407
rect 993 5393 1007 5407
rect 1233 5393 1247 5407
rect 1273 5393 1287 5407
rect 1513 5393 1527 5407
rect 1553 5393 1567 5407
rect 1793 5393 1807 5407
rect 1833 5393 1847 5407
rect 1933 5393 1947 5407
rect 1973 5393 1987 5407
rect 2053 5393 2067 5407
rect 2093 5393 2107 5407
rect 2333 5393 2347 5407
rect 2613 5393 2627 5407
rect 2653 5393 2667 5407
rect 2753 5393 2767 5407
rect 2793 5393 2807 5407
rect 3113 5393 3127 5407
rect 3153 5393 3167 5407
rect 3273 5393 3287 5407
rect 3313 5393 3327 5407
rect 3393 5393 3407 5407
rect 3433 5393 3447 5407
rect 3673 5393 3687 5407
rect 3713 5393 3727 5407
rect 3933 5393 3947 5407
rect 3973 5393 3987 5407
rect 4213 5393 4227 5407
rect 4253 5393 4267 5407
rect 4333 5393 4347 5407
rect 4373 5393 4387 5407
rect 5593 5393 5607 5407
rect 5633 5393 5647 5407
rect 5713 5393 5727 5407
rect 5753 5393 5767 5407
rect 73 5173 87 5187
rect 113 5173 127 5187
rect 453 5173 467 5187
rect 493 5173 507 5187
rect 873 5173 887 5187
rect 913 5173 927 5187
rect 1013 5173 1027 5187
rect 1053 5173 1067 5187
rect 1253 5173 1267 5187
rect 1293 5173 1307 5187
rect 2173 5173 2187 5187
rect 2213 5173 2227 5187
rect 2313 5173 2327 5187
rect 2353 5173 2367 5187
rect 3013 5173 3027 5187
rect 3633 5173 3647 5187
rect 3673 5173 3687 5187
rect 3773 5173 3787 5187
rect 3813 5173 3827 5187
rect 3913 5173 3927 5187
rect 3953 5173 3967 5187
rect 4033 5173 4047 5187
rect 4073 5173 4087 5187
rect 4573 5173 4587 5187
rect 4613 5173 4627 5187
rect 5593 5173 5607 5187
rect 5633 5173 5647 5187
rect 5693 5173 5707 5187
rect 5733 5173 5747 5187
rect 93 5153 107 5167
rect 133 5153 147 5167
rect 193 5153 207 5167
rect 233 5153 247 5167
rect 353 5153 367 5167
rect 473 5153 487 5167
rect 513 5153 527 5167
rect 573 5153 587 5167
rect 613 5153 627 5167
rect 753 5153 767 5167
rect 793 5153 807 5167
rect 853 5153 867 5167
rect 893 5153 907 5167
rect 1033 5153 1047 5167
rect 1073 5153 1087 5167
rect 1153 5153 1167 5167
rect 1273 5153 1287 5167
rect 1313 5153 1327 5167
rect 1413 5153 1427 5167
rect 1453 5153 1467 5167
rect 1553 5153 1567 5167
rect 1653 5153 1667 5167
rect 1693 5153 1707 5167
rect 1833 5153 1847 5167
rect 1893 5153 1907 5167
rect 2053 5153 2067 5167
rect 2093 5153 2107 5167
rect 2193 5153 2207 5167
rect 2333 5153 2347 5167
rect 2373 5153 2387 5167
rect 2473 5153 2487 5167
rect 2513 5153 2527 5167
rect 2593 5153 2607 5167
rect 2693 5153 2707 5167
rect 2733 5153 2747 5167
rect 2853 5153 2867 5167
rect 2893 5153 2907 5167
rect 3273 5153 3287 5167
rect 3513 5153 3527 5167
rect 3553 5153 3567 5167
rect 3653 5153 3667 5167
rect 3793 5153 3807 5167
rect 3933 5153 3947 5167
rect 4013 5153 4027 5167
rect 4053 5153 4067 5167
rect 4173 5153 4187 5167
rect 4213 5153 4227 5167
rect 4333 5153 4347 5167
rect 4373 5153 4387 5167
rect 4473 5153 4487 5167
rect 4593 5153 4607 5167
rect 4633 5153 4647 5167
rect 4693 5153 4707 5167
rect 4733 5153 4747 5167
rect 5213 5153 5227 5167
rect 5253 5153 5267 5167
rect 5353 5153 5367 5167
rect 5453 5153 5467 5167
rect 5493 5153 5507 5167
rect 5613 5153 5627 5167
rect 5713 5153 5727 5167
rect 253 5133 267 5147
rect 633 5133 647 5147
rect 733 5133 747 5147
rect 1433 5133 1447 5147
rect 1473 5133 1487 5147
rect 1673 5133 1687 5147
rect 1713 5133 1727 5147
rect 1873 5133 1887 5147
rect 1933 5133 1947 5147
rect 2033 5133 2047 5147
rect 2073 5133 2087 5147
rect 2113 5133 2127 5147
rect 2453 5133 2467 5147
rect 2713 5133 2727 5147
rect 2753 5133 2767 5147
rect 2873 5133 2887 5147
rect 2913 5133 2927 5147
rect 2993 5133 3007 5147
rect 3053 5133 3067 5147
rect 3113 5133 3127 5147
rect 3153 5133 3167 5147
rect 3373 5133 3387 5147
rect 3413 5133 3427 5147
rect 3533 5133 3547 5147
rect 3573 5133 3587 5147
rect 4193 5133 4207 5147
rect 4233 5133 4247 5147
rect 4313 5133 4327 5147
rect 4353 5133 4367 5147
rect 4753 5133 4767 5147
rect 4833 5133 4847 5147
rect 4873 5133 4887 5147
rect 4933 5133 4947 5147
rect 5013 5133 5027 5147
rect 5053 5133 5067 5147
rect 5193 5133 5207 5147
rect 5233 5133 5247 5147
rect 5433 5133 5447 5147
rect 5473 5133 5487 5147
rect 213 5113 227 5127
rect 333 5113 347 5127
rect 593 5113 607 5127
rect 773 5113 787 5127
rect 1133 5113 1147 5127
rect 1573 5113 1587 5127
rect 2493 5113 2507 5127
rect 2613 5113 2627 5127
rect 3133 5113 3147 5127
rect 3293 5113 3307 5127
rect 3393 5113 3407 5127
rect 4453 5113 4467 5127
rect 4713 5113 4727 5127
rect 4853 5113 4867 5127
rect 5333 5113 5347 5127
rect 1073 4973 1087 4987
rect 1333 4973 1347 4987
rect 1833 4973 1847 4987
rect 2133 4973 2147 4987
rect 2273 4973 2287 4987
rect 2653 4973 2667 4987
rect 2853 4973 2867 4987
rect 3433 4973 3447 4987
rect 3513 4973 3527 4987
rect 3693 4973 3707 4987
rect 3953 4973 3967 4987
rect 4453 4973 4467 4987
rect 4613 4973 4627 4987
rect 93 4953 107 4967
rect 133 4953 147 4967
rect 473 4953 487 4967
rect 513 4953 527 4967
rect 773 4953 787 4967
rect 813 4953 827 4967
rect 913 4953 927 4967
rect 953 4953 967 4967
rect 1033 4953 1047 4967
rect 1193 4953 1207 4967
rect 1233 4953 1247 4967
rect 1713 4953 1727 4967
rect 1753 4953 1767 4967
rect 1873 4953 1887 4967
rect 2093 4953 2107 4967
rect 2373 4953 2387 4967
rect 2413 4953 2427 4967
rect 3133 4953 3147 4967
rect 3173 4953 3187 4967
rect 3273 4953 3287 4967
rect 3313 4953 3327 4967
rect 3393 4953 3407 4967
rect 3533 4953 3547 4967
rect 3673 4953 3687 4967
rect 3713 4953 3727 4967
rect 4313 4953 4327 4967
rect 4373 4953 4387 4967
rect 4473 4953 4487 4967
rect 4593 4953 4607 4967
rect 4633 4953 4647 4967
rect 4753 4953 4767 4967
rect 4793 4953 4807 4967
rect 4833 4953 4847 4967
rect 4913 4953 4927 4967
rect 4953 4953 4967 4967
rect 5093 4953 5107 4967
rect 5133 4953 5147 4967
rect 5213 4953 5227 4967
rect 5293 4953 5307 4967
rect 5333 4953 5347 4967
rect 73 4933 87 4947
rect 113 4933 127 4947
rect 233 4933 247 4947
rect 273 4933 287 4947
rect 333 4933 347 4947
rect 373 4933 387 4947
rect 493 4933 507 4947
rect 533 4933 547 4947
rect 653 4933 667 4947
rect 753 4933 767 4947
rect 793 4933 807 4947
rect 893 4933 907 4947
rect 933 4933 947 4947
rect 1053 4933 1067 4947
rect 1093 4933 1107 4947
rect 1173 4933 1187 4947
rect 1213 4933 1227 4947
rect 1313 4933 1327 4947
rect 1433 4933 1447 4947
rect 1573 4933 1587 4947
rect 1613 4933 1627 4947
rect 1693 4933 1707 4947
rect 1733 4933 1747 4947
rect 1813 4933 1827 4947
rect 1853 4933 1867 4947
rect 1973 4933 1987 4947
rect 2113 4933 2127 4947
rect 2153 4933 2167 4947
rect 2253 4933 2267 4947
rect 2353 4933 2367 4947
rect 2393 4933 2407 4947
rect 2513 4933 2527 4947
rect 2553 4933 2567 4947
rect 2633 4933 2647 4947
rect 2773 4933 2787 4947
rect 2873 4933 2887 4947
rect 2953 4933 2967 4947
rect 2993 4933 3007 4947
rect 3113 4933 3127 4947
rect 3153 4933 3167 4947
rect 3253 4933 3267 4947
rect 3293 4933 3307 4947
rect 3413 4933 3427 4947
rect 3453 4933 3467 4947
rect 3573 4933 3587 4947
rect 3813 4933 3827 4947
rect 3853 4933 3867 4947
rect 3933 4933 3947 4947
rect 4013 4933 4027 4947
rect 4053 4933 4067 4947
rect 4153 4933 4167 4947
rect 4193 4933 4207 4947
rect 4513 4933 4527 4947
rect 4733 4933 4747 4947
rect 4773 4933 4787 4947
rect 5113 4933 5127 4947
rect 5153 4933 5167 4947
rect 5513 4933 5527 4947
rect 5613 4933 5627 4947
rect 5753 4933 5767 4947
rect 213 4913 227 4927
rect 253 4913 267 4927
rect 353 4913 367 4927
rect 393 4913 407 4927
rect 633 4913 647 4927
rect 673 4913 687 4927
rect 1413 4913 1427 4927
rect 1453 4913 1467 4927
rect 1553 4913 1567 4927
rect 1593 4913 1607 4927
rect 1953 4913 1967 4927
rect 1993 4913 2007 4927
rect 2493 4913 2507 4927
rect 2533 4913 2547 4927
rect 2753 4913 2767 4927
rect 2793 4913 2807 4927
rect 2973 4913 2987 4927
rect 3013 4913 3027 4927
rect 3793 4913 3807 4927
rect 3833 4913 3847 4927
rect 4033 4913 4047 4927
rect 4073 4913 4087 4927
rect 4173 4913 4187 4927
rect 4213 4913 4227 4927
rect 4333 4913 4347 4927
rect 5493 4913 5507 4927
rect 5533 4913 5547 4927
rect 5593 4913 5607 4927
rect 5633 4913 5647 4927
rect 5733 4913 5747 4927
rect 5773 4913 5787 4927
rect 213 4693 227 4707
rect 253 4693 267 4707
rect 473 4693 487 4707
rect 513 4693 527 4707
rect 613 4693 627 4707
rect 653 4693 667 4707
rect 773 4693 787 4707
rect 813 4693 827 4707
rect 1593 4693 1607 4707
rect 1633 4693 1647 4707
rect 1873 4693 1887 4707
rect 1913 4693 1927 4707
rect 2133 4693 2147 4707
rect 2173 4693 2187 4707
rect 2373 4693 2387 4707
rect 2413 4693 2427 4707
rect 2493 4693 2507 4707
rect 2533 4693 2547 4707
rect 2753 4693 2767 4707
rect 2793 4693 2807 4707
rect 3193 4693 3207 4707
rect 3233 4693 3247 4707
rect 3313 4693 3327 4707
rect 3353 4693 3367 4707
rect 3593 4693 3607 4707
rect 3633 4693 3647 4707
rect 3873 4693 3887 4707
rect 3913 4693 3927 4707
rect 4013 4693 4027 4707
rect 4053 4693 4067 4707
rect 4273 4693 4287 4707
rect 4413 4693 4427 4707
rect 4453 4693 4467 4707
rect 4553 4693 4567 4707
rect 4593 4693 4607 4707
rect 5153 4693 5167 4707
rect 5193 4693 5207 4707
rect 5273 4693 5287 4707
rect 5313 4693 5327 4707
rect 5413 4693 5427 4707
rect 5453 4693 5467 4707
rect 5533 4693 5547 4707
rect 5573 4693 5587 4707
rect 5673 4693 5687 4707
rect 5713 4693 5727 4707
rect 93 4673 107 4687
rect 133 4673 147 4687
rect 233 4673 247 4687
rect 273 4673 287 4687
rect 333 4673 347 4687
rect 373 4673 387 4687
rect 493 4673 507 4687
rect 633 4673 647 4687
rect 673 4673 687 4687
rect 793 4673 807 4687
rect 833 4673 847 4687
rect 913 4673 927 4687
rect 1013 4673 1027 4687
rect 1113 4673 1127 4687
rect 1213 4673 1227 4687
rect 1253 4673 1267 4687
rect 1353 4673 1367 4687
rect 1393 4673 1407 4687
rect 1493 4673 1507 4687
rect 1573 4673 1587 4687
rect 1613 4673 1627 4687
rect 1733 4673 1747 4687
rect 1773 4673 1787 4687
rect 1893 4673 1907 4687
rect 1993 4673 2007 4687
rect 2033 4673 2047 4687
rect 2153 4673 2167 4687
rect 2193 4673 2207 4687
rect 2393 4673 2407 4687
rect 2513 4673 2527 4687
rect 2733 4673 2747 4687
rect 2773 4673 2787 4687
rect 3033 4673 3047 4687
rect 3073 4673 3087 4687
rect 3213 4673 3227 4687
rect 3333 4673 3347 4687
rect 3373 4673 3387 4687
rect 3473 4673 3487 4687
rect 3513 4673 3527 4687
rect 3613 4673 3627 4687
rect 3653 4673 3667 4687
rect 3753 4673 3767 4687
rect 3793 4673 3807 4687
rect 3853 4673 3867 4687
rect 3893 4673 3907 4687
rect 3993 4673 4007 4687
rect 4033 4673 4047 4687
rect 4153 4673 4167 4687
rect 4433 4673 4447 4687
rect 4473 4673 4487 4687
rect 4533 4673 4547 4687
rect 4573 4673 4587 4687
rect 4693 4673 4707 4687
rect 5033 4673 5047 4687
rect 5073 4673 5087 4687
rect 5173 4673 5187 4687
rect 5293 4673 5307 4687
rect 5433 4673 5447 4687
rect 5553 4673 5567 4687
rect 5693 4673 5707 4687
rect 5733 4673 5747 4687
rect 73 4653 87 4667
rect 393 4653 407 4667
rect 1233 4653 1247 4667
rect 1273 4653 1287 4667
rect 1333 4653 1347 4667
rect 1373 4653 1387 4667
rect 1753 4653 1767 4667
rect 1793 4653 1807 4667
rect 1973 4653 1987 4667
rect 2013 4653 2027 4667
rect 2273 4653 2287 4667
rect 2313 4653 2327 4667
rect 2633 4653 2647 4667
rect 2673 4653 2687 4667
rect 2893 4653 2907 4667
rect 2933 4653 2947 4667
rect 3013 4653 3027 4667
rect 3053 4653 3067 4667
rect 3093 4653 3107 4667
rect 3453 4653 3467 4667
rect 3733 4653 3747 4667
rect 4253 4653 4267 4667
rect 4313 4653 4327 4667
rect 4753 4653 4767 4667
rect 4833 4653 4847 4667
rect 4873 4653 4887 4667
rect 5013 4653 5027 4667
rect 5053 4653 5067 4667
rect 113 4633 127 4647
rect 353 4633 367 4647
rect 893 4633 907 4647
rect 993 4633 1007 4647
rect 1133 4633 1147 4647
rect 1473 4633 1487 4647
rect 2913 4633 2927 4647
rect 3493 4633 3507 4647
rect 3773 4633 3787 4647
rect 4133 4633 4147 4647
rect 4673 4633 4687 4647
rect 353 4493 367 4507
rect 773 4493 787 4507
rect 893 4493 907 4507
rect 1053 4493 1067 4507
rect 1313 4493 1327 4507
rect 1433 4493 1447 4507
rect 1933 4493 1947 4507
rect 2753 4493 2767 4507
rect 2853 4493 2867 4507
rect 3213 4493 3227 4507
rect 3813 4493 3827 4507
rect 4753 4493 4767 4507
rect 5493 4493 5507 4507
rect 93 4473 107 4487
rect 133 4473 147 4487
rect 393 4473 407 4487
rect 533 4473 547 4487
rect 573 4473 587 4487
rect 673 4473 687 4487
rect 713 4473 727 4487
rect 933 4473 947 4487
rect 1273 4473 1287 4487
rect 1493 4473 1507 4487
rect 1533 4473 1547 4487
rect 1913 4473 1927 4487
rect 1953 4473 1967 4487
rect 2833 4473 2847 4487
rect 2873 4473 2887 4487
rect 3313 4473 3327 4487
rect 3353 4473 3367 4487
rect 3473 4473 3487 4487
rect 3533 4473 3547 4487
rect 3793 4473 3807 4487
rect 4013 4473 4027 4487
rect 4053 4473 4067 4487
rect 4113 4473 4127 4487
rect 4173 4473 4187 4487
rect 4413 4473 4427 4487
rect 4453 4473 4467 4487
rect 4973 4473 4987 4487
rect 5013 4473 5027 4487
rect 5093 4473 5107 4487
rect 5173 4473 5187 4487
rect 5213 4473 5227 4487
rect 5353 4473 5367 4487
rect 5393 4473 5407 4487
rect 5513 4473 5527 4487
rect 5673 4473 5687 4487
rect 5713 4473 5727 4487
rect 73 4453 87 4467
rect 113 4453 127 4467
rect 233 4453 247 4467
rect 273 4453 287 4467
rect 333 4453 347 4467
rect 373 4453 387 4467
rect 513 4453 527 4467
rect 553 4453 567 4467
rect 653 4453 667 4467
rect 693 4453 707 4467
rect 793 4453 807 4467
rect 873 4453 887 4467
rect 913 4453 927 4467
rect 1033 4453 1047 4467
rect 1153 4453 1167 4467
rect 1193 4453 1207 4467
rect 1293 4453 1307 4467
rect 1333 4453 1347 4467
rect 1413 4453 1427 4467
rect 1513 4453 1527 4467
rect 1553 4453 1567 4467
rect 1673 4453 1687 4467
rect 1793 4453 1807 4467
rect 1833 4453 1847 4467
rect 2053 4453 2067 4467
rect 2093 4453 2107 4467
rect 2213 4453 2227 4467
rect 2253 4453 2267 4467
rect 2353 4453 2367 4467
rect 2473 4453 2487 4467
rect 2513 4453 2527 4467
rect 2573 4453 2587 4467
rect 2613 4453 2627 4467
rect 2733 4453 2747 4467
rect 2973 4453 2987 4467
rect 3013 4453 3027 4467
rect 3113 4453 3127 4467
rect 3153 4453 3167 4467
rect 3233 4453 3247 4467
rect 3333 4453 3347 4467
rect 3373 4453 3387 4467
rect 3633 4453 3647 4467
rect 3753 4453 3767 4467
rect 3893 4453 3907 4467
rect 4293 4453 4307 4467
rect 4393 4453 4407 4467
rect 4433 4453 4447 4467
rect 4533 4453 4547 4467
rect 4673 4453 4687 4467
rect 4773 4453 4787 4467
rect 4873 4453 4887 4467
rect 4993 4453 5007 4467
rect 5033 4453 5047 4467
rect 5373 4453 5387 4467
rect 5413 4453 5427 4467
rect 5553 4453 5567 4467
rect 5653 4453 5667 4467
rect 5693 4453 5707 4467
rect 213 4433 227 4447
rect 253 4433 267 4447
rect 1133 4433 1147 4447
rect 1173 4433 1187 4447
rect 1653 4433 1667 4447
rect 1693 4433 1707 4447
rect 1773 4433 1787 4447
rect 1813 4433 1827 4447
rect 2033 4433 2047 4447
rect 2073 4433 2087 4447
rect 2193 4433 2207 4447
rect 2233 4433 2247 4447
rect 2333 4433 2347 4447
rect 2373 4433 2387 4447
rect 2453 4433 2467 4447
rect 2493 4433 2507 4447
rect 2593 4433 2607 4447
rect 2633 4433 2647 4447
rect 2953 4433 2967 4447
rect 2993 4433 3007 4447
rect 3093 4433 3107 4447
rect 3133 4433 3147 4447
rect 3493 4433 3507 4447
rect 3613 4433 3627 4447
rect 3653 4433 3667 4447
rect 3873 4433 3887 4447
rect 3913 4433 3927 4447
rect 4153 4433 4167 4447
rect 4273 4433 4287 4447
rect 4313 4433 4327 4447
rect 4513 4433 4527 4447
rect 4553 4433 4567 4447
rect 4653 4433 4667 4447
rect 4693 4433 4707 4447
rect 4853 4433 4867 4447
rect 4893 4433 4907 4447
rect 393 4213 407 4227
rect 433 4213 447 4227
rect 533 4213 547 4227
rect 573 4213 587 4227
rect 1213 4213 1227 4227
rect 1253 4213 1267 4227
rect 1353 4213 1367 4227
rect 1393 4213 1407 4227
rect 1473 4213 1487 4227
rect 1513 4213 1527 4227
rect 1713 4213 1727 4227
rect 1753 4213 1767 4227
rect 1853 4213 1867 4227
rect 1893 4213 1907 4227
rect 1993 4213 2007 4227
rect 2033 4213 2047 4227
rect 2133 4213 2147 4227
rect 2173 4213 2187 4227
rect 2573 4213 2587 4227
rect 2613 4213 2627 4227
rect 2833 4213 2847 4227
rect 2873 4213 2887 4227
rect 2953 4213 2967 4227
rect 2993 4213 3007 4227
rect 3633 4213 3647 4227
rect 3673 4213 3687 4227
rect 3773 4213 3787 4227
rect 3813 4213 3827 4227
rect 3913 4213 3927 4227
rect 3953 4213 3967 4227
rect 4053 4213 4067 4227
rect 4093 4213 4107 4227
rect 4173 4213 4187 4227
rect 4213 4213 4227 4227
rect 93 4193 107 4207
rect 133 4193 147 4207
rect 233 4193 247 4207
rect 273 4193 287 4207
rect 413 4193 427 4207
rect 453 4193 467 4207
rect 553 4193 567 4207
rect 593 4193 607 4207
rect 673 4193 687 4207
rect 813 4193 827 4207
rect 853 4193 867 4207
rect 953 4193 967 4207
rect 1073 4193 1087 4207
rect 1113 4193 1127 4207
rect 1233 4193 1247 4207
rect 1273 4193 1287 4207
rect 1373 4193 1387 4207
rect 1493 4193 1507 4207
rect 1733 4193 1747 4207
rect 1773 4193 1787 4207
rect 1873 4193 1887 4207
rect 1913 4193 1927 4207
rect 1973 4193 1987 4207
rect 2013 4193 2027 4207
rect 2113 4193 2127 4207
rect 2153 4193 2167 4207
rect 2413 4193 2427 4207
rect 2453 4193 2467 4207
rect 2593 4193 2607 4207
rect 2633 4193 2647 4207
rect 2713 4193 2727 4207
rect 2813 4193 2827 4207
rect 2853 4193 2867 4207
rect 2973 4193 2987 4207
rect 3073 4193 3087 4207
rect 3113 4193 3127 4207
rect 3213 4193 3227 4207
rect 3253 4193 3267 4207
rect 3373 4193 3387 4207
rect 3413 4193 3427 4207
rect 3533 4193 3547 4207
rect 3613 4193 3627 4207
rect 3653 4193 3667 4207
rect 3753 4193 3767 4207
rect 3793 4193 3807 4207
rect 3933 4193 3947 4207
rect 4073 4193 4087 4207
rect 4193 4193 4207 4207
rect 4293 4193 4307 4207
rect 4333 4193 4347 4207
rect 4473 4193 4487 4207
rect 4573 4193 4587 4207
rect 4613 4193 4627 4207
rect 4733 4193 4747 4207
rect 4773 4193 4787 4207
rect 4993 4193 5007 4207
rect 5093 4193 5107 4207
rect 5133 4193 5147 4207
rect 5253 4193 5267 4207
rect 5293 4193 5307 4207
rect 5393 4193 5407 4207
rect 5493 4193 5507 4207
rect 5533 4193 5547 4207
rect 113 4173 127 4187
rect 153 4173 167 4187
rect 253 4173 267 4187
rect 293 4173 307 4187
rect 713 4173 727 4187
rect 833 4173 847 4187
rect 873 4173 887 4187
rect 1053 4173 1067 4187
rect 1593 4173 1607 4187
rect 1633 4173 1647 4187
rect 2273 4173 2287 4187
rect 2313 4173 2327 4187
rect 2433 4173 2447 4187
rect 2473 4173 2487 4187
rect 3133 4173 3147 4187
rect 3273 4173 3287 4187
rect 3353 4173 3367 4187
rect 3393 4173 3407 4187
rect 4313 4173 4327 4187
rect 4353 4173 4367 4187
rect 4433 4173 4447 4187
rect 4593 4173 4607 4187
rect 4633 4173 4647 4187
rect 4713 4173 4727 4187
rect 4753 4173 4767 4187
rect 4853 4173 4867 4187
rect 4893 4173 4907 4187
rect 5153 4173 5167 4187
rect 5233 4173 5247 4187
rect 5273 4173 5287 4187
rect 5473 4173 5487 4187
rect 5513 4173 5527 4187
rect 5653 4173 5667 4187
rect 5693 4173 5707 4187
rect 5773 4173 5787 4187
rect 733 4153 747 4167
rect 933 4153 947 4167
rect 1093 4153 1107 4167
rect 1613 4153 1627 4167
rect 2293 4153 2307 4167
rect 2693 4153 2707 4167
rect 3093 4153 3107 4167
rect 3233 4153 3247 4167
rect 3513 4153 3527 4167
rect 4413 4153 4427 4167
rect 4873 4153 4887 4167
rect 4973 4153 4987 4167
rect 5113 4153 5127 4167
rect 5373 4153 5387 4167
rect 93 4013 107 4027
rect 353 4013 367 4027
rect 453 4013 467 4027
rect 613 4013 627 4027
rect 753 4013 767 4027
rect 953 4013 967 4027
rect 1533 4013 1547 4027
rect 1633 4013 1647 4027
rect 1753 4013 1767 4027
rect 3093 4013 3107 4027
rect 3333 4013 3347 4027
rect 3733 4013 3747 4027
rect 4133 4013 4147 4027
rect 4613 4013 4627 4027
rect 5013 4013 5027 4027
rect 5153 4013 5167 4027
rect 173 3993 187 4007
rect 213 3993 227 4007
rect 493 3993 507 4007
rect 593 3993 607 4007
rect 633 3993 647 4007
rect 813 3993 827 4007
rect 853 3993 867 4007
rect 1193 3993 1207 4007
rect 1233 3993 1247 4007
rect 1273 3993 1287 4007
rect 1613 3993 1627 4007
rect 1653 3993 1667 4007
rect 1993 3993 2007 4007
rect 2033 3993 2047 4007
rect 2433 3993 2447 4007
rect 2473 3993 2487 4007
rect 3433 3993 3447 4007
rect 3473 3993 3487 4007
rect 3713 3993 3727 4007
rect 3973 3993 3987 4007
rect 4013 3993 4027 4007
rect 4093 3993 4107 4007
rect 4333 3993 4347 4007
rect 4373 3993 4387 4007
rect 4473 3993 4487 4007
rect 4513 3993 4527 4007
rect 4633 3993 4647 4007
rect 5193 3993 5207 4007
rect 5273 3993 5287 4007
rect 5313 3993 5327 4007
rect 5433 3993 5447 4007
rect 5513 3993 5527 4007
rect 5553 3993 5567 4007
rect 5693 3993 5707 4007
rect 5733 3993 5747 4007
rect 73 3973 87 3987
rect 193 3973 207 3987
rect 233 3973 247 3987
rect 333 3973 347 3987
rect 433 3973 447 3987
rect 473 3973 487 3987
rect 733 3973 747 3987
rect 833 3973 847 3987
rect 873 3973 887 3987
rect 973 3973 987 3987
rect 1053 3973 1067 3987
rect 1093 3973 1107 3987
rect 1213 3973 1227 3987
rect 1253 3973 1267 3987
rect 1393 3973 1407 3987
rect 1513 3973 1527 3987
rect 1733 3973 1747 3987
rect 1813 3973 1827 3987
rect 1853 3973 1867 3987
rect 1973 3973 1987 3987
rect 2013 3973 2027 3987
rect 2153 3973 2167 3987
rect 2193 3973 2207 3987
rect 2253 3973 2267 3987
rect 2293 3973 2307 3987
rect 2413 3973 2427 3987
rect 2453 3973 2467 3987
rect 2573 3973 2587 3987
rect 2673 3973 2687 3987
rect 2773 3973 2787 3987
rect 2813 3973 2827 3987
rect 2913 3973 2927 3987
rect 2953 3973 2967 3987
rect 3073 3973 3087 3987
rect 3193 3973 3207 3987
rect 3233 3973 3247 3987
rect 3313 3973 3327 3987
rect 3413 3973 3427 3987
rect 3453 3973 3467 3987
rect 3553 3973 3567 3987
rect 3673 3973 3687 3987
rect 3833 3973 3847 3987
rect 3953 3973 3967 3987
rect 3993 3973 4007 3987
rect 4113 3973 4127 3987
rect 4153 3973 4167 3987
rect 4233 3973 4247 3987
rect 4353 3973 4367 3987
rect 4393 3973 4407 3987
rect 4493 3973 4507 3987
rect 4533 3973 4547 3987
rect 4673 3973 4687 3987
rect 4793 3973 4807 3987
rect 4873 3973 4887 3987
rect 4913 3973 4927 3987
rect 5033 3973 5047 3987
rect 5133 3973 5147 3987
rect 5713 3973 5727 3987
rect 5753 3973 5767 3987
rect 1073 3953 1087 3967
rect 1113 3953 1127 3967
rect 1373 3953 1387 3967
rect 1413 3953 1427 3967
rect 1833 3953 1847 3967
rect 1873 3953 1887 3967
rect 2133 3953 2147 3967
rect 2173 3953 2187 3967
rect 2273 3953 2287 3967
rect 2313 3953 2327 3967
rect 2553 3953 2567 3967
rect 2593 3953 2607 3967
rect 2653 3953 2667 3967
rect 2693 3953 2707 3967
rect 2793 3953 2807 3967
rect 2833 3953 2847 3967
rect 2933 3953 2947 3967
rect 2973 3953 2987 3967
rect 3173 3953 3187 3967
rect 3213 3953 3227 3967
rect 3533 3953 3547 3967
rect 3573 3953 3587 3967
rect 3813 3953 3827 3967
rect 3853 3953 3867 3967
rect 4213 3953 4227 3967
rect 4253 3953 4267 3967
rect 4773 3953 4787 3967
rect 4813 3953 4827 3967
rect 4893 3953 4907 3967
rect 4933 3953 4947 3967
rect 73 3733 87 3747
rect 113 3733 127 3747
rect 193 3733 207 3747
rect 233 3733 247 3747
rect 693 3733 707 3747
rect 733 3733 747 3747
rect 1113 3733 1127 3747
rect 1153 3733 1167 3747
rect 1253 3733 1267 3747
rect 1293 3733 1307 3747
rect 1773 3733 1787 3747
rect 1813 3733 1827 3747
rect 1873 3733 1887 3747
rect 1913 3733 1927 3747
rect 2133 3733 2147 3747
rect 2173 3733 2187 3747
rect 2273 3733 2287 3747
rect 2313 3733 2327 3747
rect 2533 3733 2547 3747
rect 2573 3733 2587 3747
rect 3033 3733 3047 3747
rect 3073 3733 3087 3747
rect 3193 3733 3207 3747
rect 3233 3733 3247 3747
rect 3413 3733 3427 3747
rect 3453 3733 3467 3747
rect 3773 3733 3787 3747
rect 3813 3733 3827 3747
rect 4493 3733 4507 3747
rect 4533 3733 4547 3747
rect 5013 3733 5027 3747
rect 5053 3733 5067 3747
rect 5713 3733 5727 3747
rect 5753 3733 5767 3747
rect 93 3713 107 3727
rect 213 3713 227 3727
rect 253 3713 267 3727
rect 353 3713 367 3727
rect 413 3713 427 3727
rect 553 3713 567 3727
rect 593 3713 607 3727
rect 713 3713 727 3727
rect 813 3713 827 3727
rect 853 3713 867 3727
rect 993 3713 1007 3727
rect 1033 3713 1047 3727
rect 1133 3713 1147 3727
rect 1233 3713 1247 3727
rect 1273 3713 1287 3727
rect 1373 3713 1387 3727
rect 1413 3713 1427 3727
rect 1533 3713 1547 3727
rect 1573 3713 1587 3727
rect 1673 3713 1687 3727
rect 1793 3713 1807 3727
rect 1893 3713 1907 3727
rect 2053 3713 2067 3727
rect 2153 3713 2167 3727
rect 2253 3713 2267 3727
rect 2293 3713 2307 3727
rect 2413 3713 2427 3727
rect 2453 3713 2467 3727
rect 2553 3713 2567 3727
rect 2673 3713 2687 3727
rect 2713 3713 2727 3727
rect 2813 3713 2827 3727
rect 2913 3713 2927 3727
rect 2953 3713 2967 3727
rect 3053 3713 3067 3727
rect 3213 3713 3227 3727
rect 3313 3713 3327 3727
rect 3393 3713 3407 3727
rect 3433 3713 3447 3727
rect 3553 3713 3567 3727
rect 3793 3713 3807 3727
rect 3913 3713 3927 3727
rect 4013 3713 4027 3727
rect 4373 3713 4387 3727
rect 4413 3713 4427 3727
rect 4513 3713 4527 3727
rect 4753 3713 4767 3727
rect 4793 3713 4807 3727
rect 4873 3713 4887 3727
rect 5033 3713 5047 3727
rect 5133 3713 5147 3727
rect 5233 3713 5247 3727
rect 5373 3713 5387 3727
rect 5733 3713 5747 3727
rect 393 3693 407 3707
rect 453 3693 467 3707
rect 573 3693 587 3707
rect 613 3693 627 3707
rect 793 3693 807 3707
rect 833 3693 847 3707
rect 973 3693 987 3707
rect 1013 3693 1027 3707
rect 1053 3693 1067 3707
rect 1433 3693 1447 3707
rect 1513 3693 1527 3707
rect 1553 3693 1567 3707
rect 2013 3693 2027 3707
rect 2433 3693 2447 3707
rect 2473 3693 2487 3707
rect 2653 3693 2667 3707
rect 2693 3693 2707 3707
rect 2933 3693 2947 3707
rect 2973 3693 2987 3707
rect 3653 3693 3667 3707
rect 3693 3693 3707 3707
rect 4073 3693 4087 3707
rect 4153 3693 4167 3707
rect 4193 3693 4207 3707
rect 4353 3693 4367 3707
rect 4393 3693 4407 3707
rect 4433 3693 4447 3707
rect 4613 3693 4627 3707
rect 4653 3693 4667 3707
rect 4733 3693 4747 3707
rect 4773 3693 4787 3707
rect 4893 3693 4907 3707
rect 5433 3693 5447 3707
rect 5513 3693 5527 3707
rect 5553 3693 5567 3707
rect 1393 3673 1407 3687
rect 1653 3673 1667 3687
rect 1993 3673 2007 3687
rect 2833 3673 2847 3687
rect 3333 3673 3347 3687
rect 3533 3673 3547 3687
rect 3673 3673 3687 3687
rect 3893 3673 3907 3687
rect 4033 3673 4047 3687
rect 4633 3673 4647 3687
rect 5113 3673 5127 3687
rect 213 3533 227 3547
rect 333 3533 347 3547
rect 1713 3533 1727 3547
rect 1953 3533 1967 3547
rect 2433 3533 2447 3547
rect 3893 3533 3907 3547
rect 4153 3533 4167 3547
rect 93 3513 107 3527
rect 133 3513 147 3527
rect 253 3513 267 3527
rect 433 3513 447 3527
rect 473 3513 487 3527
rect 973 3513 987 3527
rect 1013 3513 1027 3527
rect 1513 3513 1527 3527
rect 1553 3513 1567 3527
rect 1673 3513 1687 3527
rect 1993 3513 2007 3527
rect 2113 3513 2127 3527
rect 2153 3513 2167 3527
rect 2233 3513 2247 3527
rect 2273 3513 2287 3527
rect 2393 3513 2407 3527
rect 2533 3513 2547 3527
rect 2593 3513 2607 3527
rect 2813 3513 2827 3527
rect 2853 3513 2867 3527
rect 2953 3513 2967 3527
rect 2993 3513 3007 3527
rect 3493 3513 3507 3527
rect 3533 3513 3547 3527
rect 3633 3513 3647 3527
rect 3673 3513 3687 3527
rect 3753 3513 3767 3527
rect 3813 3513 3827 3527
rect 3873 3513 3887 3527
rect 3913 3513 3927 3527
rect 4053 3513 4067 3527
rect 4093 3513 4107 3527
rect 4253 3513 4267 3527
rect 4293 3513 4307 3527
rect 4613 3513 4627 3527
rect 4693 3513 4707 3527
rect 4733 3513 4747 3527
rect 5033 3513 5047 3527
rect 5073 3513 5087 3527
rect 5313 3513 5327 3527
rect 5353 3513 5367 3527
rect 5433 3513 5447 3527
rect 5633 3513 5647 3527
rect 5673 3513 5687 3527
rect 73 3493 87 3507
rect 113 3493 127 3507
rect 193 3493 207 3507
rect 233 3493 247 3507
rect 353 3493 367 3507
rect 453 3493 467 3507
rect 493 3493 507 3507
rect 573 3493 587 3507
rect 613 3493 627 3507
rect 773 3493 787 3507
rect 893 3493 907 3507
rect 993 3493 1007 3507
rect 1033 3493 1047 3507
rect 1153 3493 1167 3507
rect 1193 3493 1207 3507
rect 1273 3493 1287 3507
rect 1413 3493 1427 3507
rect 1453 3493 1467 3507
rect 1533 3493 1547 3507
rect 1573 3493 1587 3507
rect 1693 3493 1707 3507
rect 1733 3493 1747 3507
rect 1833 3493 1847 3507
rect 1873 3493 1887 3507
rect 1933 3493 1947 3507
rect 1973 3493 1987 3507
rect 2093 3493 2107 3507
rect 2133 3493 2147 3507
rect 2253 3493 2267 3507
rect 2293 3493 2307 3507
rect 2413 3493 2427 3507
rect 2453 3493 2467 3507
rect 2673 3493 2687 3507
rect 2793 3493 2807 3507
rect 2833 3493 2847 3507
rect 3093 3493 3107 3507
rect 3173 3493 3187 3507
rect 3213 3493 3227 3507
rect 3353 3493 3367 3507
rect 3393 3493 3407 3507
rect 3473 3493 3487 3507
rect 3513 3493 3527 3507
rect 3613 3493 3627 3507
rect 3653 3493 3667 3507
rect 4033 3493 4047 3507
rect 4073 3493 4087 3507
rect 4173 3493 4187 3507
rect 4273 3493 4287 3507
rect 4313 3493 4327 3507
rect 4433 3493 4447 3507
rect 4533 3493 4547 3507
rect 4913 3493 4927 3507
rect 5013 3493 5027 3507
rect 5053 3493 5067 3507
rect 5173 3493 5187 3507
rect 5553 3493 5567 3507
rect 5653 3493 5667 3507
rect 5693 3493 5707 3507
rect 593 3473 607 3487
rect 633 3473 647 3487
rect 753 3473 767 3487
rect 793 3473 807 3487
rect 873 3473 887 3487
rect 913 3473 927 3487
rect 1133 3473 1147 3487
rect 1173 3473 1187 3487
rect 1253 3473 1267 3487
rect 1293 3473 1307 3487
rect 1393 3473 1407 3487
rect 1433 3473 1447 3487
rect 1813 3473 1827 3487
rect 1853 3473 1867 3487
rect 2553 3473 2567 3487
rect 2653 3473 2667 3487
rect 2693 3473 2707 3487
rect 3073 3473 3087 3487
rect 3113 3473 3127 3487
rect 3193 3473 3207 3487
rect 3233 3473 3247 3487
rect 3333 3473 3347 3487
rect 3373 3473 3387 3487
rect 3773 3473 3787 3487
rect 4413 3473 4427 3487
rect 4453 3473 4467 3487
rect 4513 3473 4527 3487
rect 4553 3473 4567 3487
rect 4893 3473 4907 3487
rect 4933 3473 4947 3487
rect 5153 3473 5167 3487
rect 5193 3473 5207 3487
rect 5533 3473 5547 3487
rect 5573 3473 5587 3487
rect 393 3253 407 3267
rect 433 3253 447 3267
rect 693 3253 707 3267
rect 833 3253 847 3267
rect 873 3253 887 3267
rect 953 3253 967 3267
rect 993 3253 1007 3267
rect 1093 3253 1107 3267
rect 1133 3253 1147 3267
rect 1473 3253 1487 3267
rect 1513 3253 1527 3267
rect 1613 3253 1627 3267
rect 1653 3253 1667 3267
rect 1913 3253 1927 3267
rect 1953 3253 1967 3267
rect 2153 3253 2167 3267
rect 2193 3253 2207 3267
rect 2313 3253 2327 3267
rect 2413 3253 2427 3267
rect 2453 3253 2467 3267
rect 2833 3253 2847 3267
rect 2873 3253 2887 3267
rect 2973 3253 2987 3267
rect 3013 3253 3027 3267
rect 3113 3253 3127 3267
rect 3153 3253 3167 3267
rect 3253 3253 3267 3267
rect 3293 3253 3307 3267
rect 3473 3253 3487 3267
rect 3513 3253 3527 3267
rect 4893 3253 4907 3267
rect 4933 3253 4947 3267
rect 5253 3253 5267 3267
rect 5293 3253 5307 3267
rect 5653 3253 5667 3267
rect 5693 3253 5707 3267
rect 73 3233 87 3247
rect 173 3233 187 3247
rect 213 3233 227 3247
rect 313 3233 327 3247
rect 413 3233 427 3247
rect 513 3233 527 3247
rect 553 3233 567 3247
rect 853 3233 867 3247
rect 973 3233 987 3247
rect 1013 3233 1027 3247
rect 1113 3233 1127 3247
rect 1153 3233 1167 3247
rect 1213 3233 1227 3247
rect 1253 3233 1267 3247
rect 1373 3233 1387 3247
rect 1493 3233 1507 3247
rect 1533 3233 1547 3247
rect 1633 3233 1647 3247
rect 1673 3233 1687 3247
rect 1773 3233 1787 3247
rect 1813 3233 1827 3247
rect 1933 3233 1947 3247
rect 2053 3233 2067 3247
rect 2093 3233 2107 3247
rect 2173 3233 2187 3247
rect 2433 3233 2447 3247
rect 2553 3233 2567 3247
rect 2593 3233 2607 3247
rect 2713 3233 2727 3247
rect 2753 3233 2767 3247
rect 2813 3233 2827 3247
rect 2853 3233 2867 3247
rect 2953 3233 2967 3247
rect 2993 3233 3007 3247
rect 3133 3233 3147 3247
rect 3273 3233 3287 3247
rect 3373 3233 3387 3247
rect 3493 3233 3507 3247
rect 3533 3233 3547 3247
rect 3593 3233 3607 3247
rect 3633 3233 3647 3247
rect 3753 3233 3767 3247
rect 3793 3233 3807 3247
rect 3893 3233 3907 3247
rect 4233 3233 4247 3247
rect 4273 3233 4287 3247
rect 4373 3233 4387 3247
rect 4413 3233 4427 3247
rect 4753 3233 4767 3247
rect 4793 3233 4807 3247
rect 4913 3233 4927 3247
rect 5013 3233 5027 3247
rect 5053 3233 5067 3247
rect 5153 3233 5167 3247
rect 5273 3233 5287 3247
rect 5373 3233 5387 3247
rect 5493 3233 5507 3247
rect 5533 3233 5547 3247
rect 5673 3233 5687 3247
rect 193 3213 207 3227
rect 233 3213 247 3227
rect 573 3213 587 3227
rect 653 3213 667 3227
rect 713 3213 727 3227
rect 1273 3213 1287 3227
rect 1753 3213 1767 3227
rect 2033 3213 2047 3227
rect 2293 3213 2307 3227
rect 2353 3213 2367 3227
rect 2573 3213 2587 3227
rect 2613 3213 2627 3227
rect 2693 3213 2707 3227
rect 3653 3213 3667 3227
rect 3773 3213 3787 3227
rect 3813 3213 3827 3227
rect 3953 3213 3967 3227
rect 4033 3213 4047 3227
rect 4073 3213 4087 3227
rect 4213 3213 4227 3227
rect 4253 3213 4267 3227
rect 4353 3213 4367 3227
rect 4393 3213 4407 3227
rect 4473 3213 4487 3227
rect 4553 3213 4567 3227
rect 4593 3213 4607 3227
rect 4733 3213 4747 3227
rect 4773 3213 4787 3227
rect 5033 3213 5047 3227
rect 5073 3213 5087 3227
rect 5473 3213 5487 3227
rect 5513 3213 5527 3227
rect 93 3193 107 3207
rect 333 3193 347 3207
rect 533 3193 547 3207
rect 1233 3193 1247 3207
rect 1393 3193 1407 3207
rect 1793 3193 1807 3207
rect 2073 3193 2087 3207
rect 2733 3193 2747 3207
rect 3353 3193 3367 3207
rect 3613 3193 3627 3207
rect 3873 3193 3887 3207
rect 5173 3193 5187 3207
rect 5353 3193 5367 3207
rect 1233 3053 1247 3067
rect 1673 3053 1687 3067
rect 2413 3053 2427 3067
rect 2553 3053 2567 3067
rect 2873 3053 2887 3067
rect 2953 3053 2967 3067
rect 3333 3053 3347 3067
rect 3833 3053 3847 3067
rect 4073 3053 4087 3067
rect 93 3033 107 3047
rect 153 3033 167 3047
rect 533 3033 547 3047
rect 573 3033 587 3047
rect 633 3033 647 3047
rect 673 3033 687 3047
rect 773 3033 787 3047
rect 813 3033 827 3047
rect 913 3033 927 3047
rect 953 3033 967 3047
rect 1213 3033 1227 3047
rect 1253 3033 1267 3047
rect 1313 3033 1327 3047
rect 1353 3033 1367 3047
rect 1633 3033 1647 3047
rect 1793 3033 1807 3047
rect 1833 3033 1847 3047
rect 1893 3033 1907 3047
rect 1933 3033 1947 3047
rect 2093 3033 2107 3047
rect 2133 3033 2147 3047
rect 2233 3033 2247 3047
rect 2273 3033 2287 3047
rect 2373 3033 2387 3047
rect 2513 3033 2527 3047
rect 2653 3033 2667 3047
rect 2693 3033 2707 3047
rect 2733 3033 2747 3047
rect 2853 3033 2867 3047
rect 2933 3033 2947 3047
rect 2973 3033 2987 3047
rect 3213 3033 3227 3047
rect 3273 3033 3287 3047
rect 3353 3033 3367 3047
rect 3513 3033 3527 3047
rect 3553 3033 3567 3047
rect 3653 3033 3667 3047
rect 3693 3033 3707 3047
rect 3813 3033 3827 3047
rect 3933 3033 3947 3047
rect 3993 3033 4007 3047
rect 4053 3033 4067 3047
rect 4093 3033 4107 3047
rect 4353 3033 4367 3047
rect 4393 3033 4407 3047
rect 4473 3033 4487 3047
rect 4573 3033 4587 3047
rect 4613 3033 4627 3047
rect 4713 3033 4727 3047
rect 4753 3033 4767 3047
rect 5133 3033 5147 3047
rect 5173 3033 5187 3047
rect 5253 3033 5267 3047
rect 5553 3033 5567 3047
rect 5633 3033 5647 3047
rect 5673 3033 5687 3047
rect 233 3013 247 3027
rect 273 3013 287 3027
rect 393 3013 407 3027
rect 513 3013 527 3027
rect 553 3013 567 3027
rect 653 3013 667 3027
rect 693 3013 707 3027
rect 793 3013 807 3027
rect 833 3013 847 3027
rect 933 3013 947 3027
rect 973 3013 987 3027
rect 1093 3013 1107 3027
rect 1333 3013 1347 3027
rect 1373 3013 1387 3027
rect 1493 3013 1507 3027
rect 1533 3013 1547 3027
rect 1653 3013 1667 3027
rect 1693 3013 1707 3027
rect 1773 3013 1787 3027
rect 1813 3013 1827 3027
rect 1913 3013 1927 3027
rect 1953 3013 1967 3027
rect 2073 3013 2087 3027
rect 2113 3013 2127 3027
rect 2213 3013 2227 3027
rect 2253 3013 2267 3027
rect 2393 3013 2407 3027
rect 2433 3013 2447 3027
rect 2533 3013 2547 3027
rect 2573 3013 2587 3027
rect 2673 3013 2687 3027
rect 2713 3013 2727 3027
rect 2813 3013 2827 3027
rect 3093 3013 3107 3027
rect 3393 3013 3407 3027
rect 3493 3013 3507 3027
rect 3533 3013 3547 3027
rect 3633 3013 3647 3027
rect 3673 3013 3687 3027
rect 3773 3013 3787 3027
rect 4173 3013 4187 3027
rect 4213 3013 4227 3027
rect 4593 3013 4607 3027
rect 4633 3013 4647 3027
rect 4733 3013 4747 3027
rect 4773 3013 4787 3027
rect 4893 3013 4907 3027
rect 4993 3013 5007 3027
rect 5353 3013 5367 3027
rect 5493 3013 5507 3027
rect 113 2993 127 3007
rect 253 2993 267 3007
rect 293 2993 307 3007
rect 373 2993 387 3007
rect 413 2993 427 3007
rect 1073 2993 1087 3007
rect 1113 2993 1127 3007
rect 1473 2993 1487 3007
rect 1513 2993 1527 3007
rect 3073 2993 3087 3007
rect 3113 2993 3127 3007
rect 3233 2993 3247 3007
rect 3953 2993 3967 3007
rect 4193 2993 4207 3007
rect 4233 2993 4247 3007
rect 4873 2993 4887 3007
rect 4913 2993 4927 3007
rect 4973 2993 4987 3007
rect 5013 2993 5027 3007
rect 73 2773 87 2787
rect 113 2773 127 2787
rect 573 2773 587 2787
rect 613 2773 627 2787
rect 713 2773 727 2787
rect 813 2773 827 2787
rect 853 2773 867 2787
rect 1073 2773 1087 2787
rect 1113 2773 1127 2787
rect 1793 2773 1807 2787
rect 1933 2773 1947 2787
rect 1973 2773 1987 2787
rect 2213 2773 2227 2787
rect 2333 2773 2347 2787
rect 2373 2773 2387 2787
rect 2593 2773 2607 2787
rect 2633 2773 2647 2787
rect 2753 2773 2767 2787
rect 3033 2773 3047 2787
rect 3073 2773 3087 2787
rect 3153 2773 3167 2787
rect 3193 2773 3207 2787
rect 3453 2773 3467 2787
rect 3693 2773 3707 2787
rect 3733 2773 3747 2787
rect 3813 2773 3827 2787
rect 3853 2773 3867 2787
rect 4173 2773 4187 2787
rect 4213 2773 4227 2787
rect 5133 2773 5147 2787
rect 5173 2773 5187 2787
rect 93 2753 107 2767
rect 193 2753 207 2767
rect 233 2753 247 2767
rect 333 2753 347 2767
rect 413 2753 427 2767
rect 453 2753 467 2767
rect 593 2753 607 2767
rect 833 2753 847 2767
rect 933 2753 947 2767
rect 973 2753 987 2767
rect 1093 2753 1107 2767
rect 1233 2753 1247 2767
rect 1273 2753 1287 2767
rect 1373 2753 1387 2767
rect 1413 2753 1427 2767
rect 1513 2753 1527 2767
rect 1953 2753 1967 2767
rect 2053 2753 2067 2767
rect 2093 2753 2107 2767
rect 2353 2753 2367 2767
rect 2613 2753 2627 2767
rect 2653 2753 2667 2767
rect 2893 2753 2907 2767
rect 2933 2753 2947 2767
rect 3053 2753 3067 2767
rect 3093 2753 3107 2767
rect 3173 2753 3187 2767
rect 3293 2753 3307 2767
rect 3333 2753 3347 2767
rect 3673 2753 3687 2767
rect 3713 2753 3727 2767
rect 3833 2753 3847 2767
rect 3973 2753 3987 2767
rect 4053 2753 4067 2767
rect 4093 2753 4107 2767
rect 4193 2753 4207 2767
rect 4293 2753 4307 2767
rect 4413 2753 4427 2767
rect 5013 2753 5027 2767
rect 5053 2753 5067 2767
rect 5153 2753 5167 2767
rect 5253 2753 5267 2767
rect 5293 2753 5307 2767
rect 5633 2753 5647 2767
rect 5673 2753 5687 2767
rect 173 2733 187 2747
rect 213 2733 227 2747
rect 473 2733 487 2747
rect 673 2733 687 2747
rect 733 2733 747 2747
rect 993 2733 1007 2747
rect 1253 2733 1267 2747
rect 1293 2733 1307 2747
rect 1353 2733 1367 2747
rect 1393 2733 1407 2747
rect 1553 2733 1567 2747
rect 1633 2733 1647 2747
rect 1673 2733 1687 2747
rect 1773 2733 1787 2747
rect 1833 2733 1847 2747
rect 2033 2733 2047 2747
rect 2073 2733 2087 2747
rect 2193 2733 2207 2747
rect 2253 2733 2267 2747
rect 2453 2733 2467 2747
rect 2493 2733 2507 2747
rect 2733 2733 2747 2747
rect 2793 2733 2807 2747
rect 2873 2733 2887 2747
rect 2913 2733 2927 2747
rect 3313 2733 3327 2747
rect 3353 2733 3367 2747
rect 3433 2733 3447 2747
rect 3493 2733 3507 2747
rect 3553 2733 3567 2747
rect 3593 2733 3607 2747
rect 3953 2733 3967 2747
rect 4073 2733 4087 2747
rect 4113 2733 4127 2747
rect 4313 2733 4327 2747
rect 4473 2733 4487 2747
rect 4553 2733 4567 2747
rect 4593 2733 4607 2747
rect 4773 2733 4787 2747
rect 4813 2733 4827 2747
rect 4893 2733 4907 2747
rect 4993 2733 5007 2747
rect 5033 2733 5047 2747
rect 5353 2733 5367 2747
rect 5433 2733 5447 2747
rect 5473 2733 5487 2747
rect 5613 2733 5627 2747
rect 5653 2733 5667 2747
rect 353 2713 367 2727
rect 433 2713 447 2727
rect 953 2713 967 2727
rect 1573 2713 1587 2727
rect 1653 2713 1667 2727
rect 2473 2713 2487 2727
rect 3573 2713 3587 2727
rect 4393 2713 4407 2727
rect 93 2573 107 2587
rect 153 2573 167 2587
rect 313 2573 327 2587
rect 533 2573 547 2587
rect 653 2573 667 2587
rect 933 2573 947 2587
rect 1593 2573 1607 2587
rect 2313 2573 2327 2587
rect 2873 2573 2887 2587
rect 2993 2573 3007 2587
rect 3913 2573 3927 2587
rect 4253 2573 4267 2587
rect 4633 2573 4647 2587
rect 273 2553 287 2567
rect 633 2553 647 2567
rect 673 2553 687 2567
rect 753 2553 767 2567
rect 793 2553 807 2567
rect 973 2553 987 2567
rect 1093 2553 1107 2567
rect 1133 2553 1147 2567
rect 1313 2553 1327 2567
rect 1373 2553 1387 2567
rect 1693 2553 1707 2567
rect 1733 2553 1747 2567
rect 1873 2553 1887 2567
rect 1913 2553 1927 2567
rect 1973 2553 1987 2567
rect 2013 2553 2027 2567
rect 2273 2553 2287 2567
rect 2573 2553 2587 2567
rect 2613 2553 2627 2567
rect 2673 2553 2687 2567
rect 2713 2553 2727 2567
rect 2833 2553 2847 2567
rect 3053 2553 3067 2567
rect 3093 2553 3107 2567
rect 3473 2553 3487 2567
rect 3533 2553 3547 2567
rect 3733 2553 3747 2567
rect 3773 2553 3787 2567
rect 3813 2553 3827 2567
rect 3893 2553 3907 2567
rect 3933 2553 3947 2567
rect 5013 2553 5027 2567
rect 5053 2553 5067 2567
rect 5133 2553 5147 2567
rect 5733 2553 5747 2567
rect 73 2533 87 2547
rect 173 2533 187 2547
rect 293 2533 307 2547
rect 333 2533 347 2547
rect 393 2533 407 2547
rect 433 2533 447 2547
rect 553 2533 567 2547
rect 773 2533 787 2547
rect 813 2533 827 2547
rect 913 2533 927 2547
rect 953 2533 967 2547
rect 1073 2533 1087 2547
rect 1113 2533 1127 2547
rect 1233 2533 1247 2547
rect 1493 2533 1507 2547
rect 1533 2533 1547 2547
rect 1613 2533 1627 2547
rect 1713 2533 1727 2547
rect 1753 2533 1767 2547
rect 1853 2533 1867 2547
rect 1893 2533 1907 2547
rect 1993 2533 2007 2547
rect 2033 2533 2047 2547
rect 2153 2533 2167 2547
rect 2193 2533 2207 2547
rect 2293 2533 2307 2547
rect 2333 2533 2347 2547
rect 2413 2533 2427 2547
rect 2553 2533 2567 2547
rect 2593 2533 2607 2547
rect 2693 2533 2707 2547
rect 2733 2533 2747 2547
rect 2853 2533 2867 2547
rect 2893 2533 2907 2547
rect 2973 2533 2987 2547
rect 3073 2533 3087 2547
rect 3113 2533 3127 2547
rect 3233 2533 3247 2547
rect 3373 2533 3387 2547
rect 3413 2533 3427 2547
rect 3633 2533 3647 2547
rect 3753 2533 3767 2547
rect 3793 2533 3807 2547
rect 3993 2533 4007 2547
rect 4073 2533 4087 2547
rect 4373 2533 4387 2547
rect 4513 2533 4527 2547
rect 4813 2533 4827 2547
rect 4893 2533 4907 2547
rect 5233 2533 5247 2547
rect 5373 2533 5387 2547
rect 5493 2533 5507 2547
rect 5633 2533 5647 2547
rect 5713 2533 5727 2547
rect 413 2513 427 2527
rect 453 2513 467 2527
rect 1213 2513 1227 2527
rect 1253 2513 1267 2527
rect 1353 2513 1367 2527
rect 1473 2513 1487 2527
rect 1513 2513 1527 2527
rect 2133 2513 2147 2527
rect 2173 2513 2187 2527
rect 2393 2513 2407 2527
rect 2433 2513 2447 2527
rect 3213 2513 3227 2527
rect 3253 2513 3267 2527
rect 3353 2513 3367 2527
rect 3393 2513 3407 2527
rect 3513 2513 3527 2527
rect 3613 2513 3627 2527
rect 3653 2513 3667 2527
rect 4413 2513 4427 2527
rect 4473 2513 4487 2527
rect 193 2293 207 2307
rect 233 2293 247 2307
rect 313 2293 327 2307
rect 353 2293 367 2307
rect 753 2293 767 2307
rect 793 2293 807 2307
rect 893 2293 907 2307
rect 933 2293 947 2307
rect 1253 2293 1267 2307
rect 1293 2293 1307 2307
rect 1833 2293 1847 2307
rect 1873 2293 1887 2307
rect 1973 2293 1987 2307
rect 2013 2293 2027 2307
rect 2493 2293 2507 2307
rect 3013 2293 3027 2307
rect 3053 2293 3067 2307
rect 3133 2293 3147 2307
rect 3173 2293 3187 2307
rect 3673 2293 3687 2307
rect 3713 2293 3727 2307
rect 4313 2293 4327 2307
rect 4433 2293 4447 2307
rect 4693 2293 4707 2307
rect 4733 2293 4747 2307
rect 5193 2293 5207 2307
rect 5233 2293 5247 2307
rect 5413 2293 5427 2307
rect 5453 2293 5467 2307
rect 213 2273 227 2287
rect 253 2273 267 2287
rect 333 2273 347 2287
rect 453 2273 467 2287
rect 493 2273 507 2287
rect 593 2273 607 2287
rect 633 2273 647 2287
rect 773 2273 787 2287
rect 813 2273 827 2287
rect 913 2273 927 2287
rect 1013 2273 1027 2287
rect 1133 2273 1147 2287
rect 1273 2273 1287 2287
rect 1313 2273 1327 2287
rect 1413 2273 1427 2287
rect 1453 2273 1467 2287
rect 1553 2273 1567 2287
rect 1593 2273 1607 2287
rect 1713 2273 1727 2287
rect 1753 2273 1767 2287
rect 1853 2273 1867 2287
rect 1893 2273 1907 2287
rect 1993 2273 2007 2287
rect 2033 2273 2047 2287
rect 2073 2273 2087 2287
rect 2153 2273 2167 2287
rect 2453 2273 2467 2287
rect 2733 2273 2747 2287
rect 2773 2273 2787 2287
rect 2873 2273 2887 2287
rect 2913 2273 2927 2287
rect 3033 2273 3047 2287
rect 3153 2273 3167 2287
rect 3293 2273 3307 2287
rect 3333 2273 3347 2287
rect 3553 2273 3567 2287
rect 3593 2273 3607 2287
rect 3693 2273 3707 2287
rect 3893 2273 3907 2287
rect 3973 2273 3987 2287
rect 4273 2273 4287 2287
rect 4553 2273 4567 2287
rect 4593 2273 4607 2287
rect 4713 2273 4727 2287
rect 4953 2273 4967 2287
rect 5053 2273 5067 2287
rect 5093 2273 5107 2287
rect 5213 2273 5227 2287
rect 5313 2273 5327 2287
rect 5433 2273 5447 2287
rect 5553 2273 5567 2287
rect 5633 2273 5647 2287
rect 5693 2273 5707 2287
rect 73 2253 87 2267
rect 113 2253 127 2267
rect 433 2253 447 2267
rect 473 2253 487 2267
rect 613 2253 627 2267
rect 653 2253 667 2267
rect 1053 2253 1067 2267
rect 1153 2253 1167 2267
rect 1393 2253 1407 2267
rect 1573 2253 1587 2267
rect 1613 2253 1627 2267
rect 1693 2253 1707 2267
rect 2593 2253 2607 2267
rect 2633 2253 2647 2267
rect 2713 2253 2727 2267
rect 2753 2253 2767 2267
rect 2853 2253 2867 2267
rect 2893 2253 2907 2267
rect 3273 2253 3287 2267
rect 3393 2253 3407 2267
rect 3433 2253 3447 2267
rect 3533 2253 3547 2267
rect 3573 2253 3587 2267
rect 3793 2253 3807 2267
rect 3833 2253 3847 2267
rect 4393 2253 4407 2267
rect 4453 2253 4467 2267
rect 4533 2253 4547 2267
rect 4573 2253 4587 2267
rect 4613 2253 4627 2267
rect 4833 2253 4847 2267
rect 4873 2253 4887 2267
rect 5033 2253 5047 2267
rect 5073 2253 5087 2267
rect 5113 2253 5127 2267
rect 5333 2253 5347 2267
rect 5653 2253 5667 2267
rect 5713 2253 5727 2267
rect 1073 2233 1087 2247
rect 1433 2233 1447 2247
rect 1733 2233 1747 2247
rect 2333 2233 2347 2247
rect 3313 2233 3327 2247
rect 3413 2233 3427 2247
rect 4153 2233 4167 2247
rect 4933 2233 4947 2247
rect 5533 2233 5547 2247
rect 373 2093 387 2107
rect 533 2093 547 2107
rect 793 2093 807 2107
rect 1513 2093 1527 2107
rect 1893 2093 1907 2107
rect 2613 2093 2627 2107
rect 3273 2093 3287 2107
rect 3533 2093 3547 2107
rect 5153 2093 5167 2107
rect 5273 2093 5287 2107
rect 5493 2093 5507 2107
rect 5633 2093 5647 2107
rect 93 2073 107 2087
rect 133 2073 147 2087
rect 413 2073 427 2087
rect 633 2073 647 2087
rect 673 2073 687 2087
rect 753 2073 767 2087
rect 1213 2073 1227 2087
rect 1253 2073 1267 2087
rect 1353 2073 1367 2087
rect 1393 2073 1407 2087
rect 1473 2073 1487 2087
rect 1733 2073 1747 2087
rect 1773 2073 1787 2087
rect 1933 2073 1947 2087
rect 2093 2073 2107 2087
rect 2153 2073 2167 2087
rect 2853 2073 2867 2087
rect 2893 2073 2907 2087
rect 3253 2073 3267 2087
rect 3293 2073 3307 2087
rect 3393 2073 3407 2087
rect 3453 2073 3467 2087
rect 3573 2073 3587 2087
rect 3693 2073 3707 2087
rect 3973 2073 3987 2087
rect 4093 2073 4107 2087
rect 4153 2073 4167 2087
rect 4373 2073 4387 2087
rect 4413 2073 4427 2087
rect 4473 2073 4487 2087
rect 4513 2073 4527 2087
rect 4913 2073 4927 2087
rect 4953 2073 4967 2087
rect 5053 2073 5067 2087
rect 5093 2073 5107 2087
rect 5253 2073 5267 2087
rect 5293 2073 5307 2087
rect 5693 2073 5707 2087
rect 5733 2073 5747 2087
rect 253 2053 267 2067
rect 293 2053 307 2067
rect 353 2053 367 2067
rect 393 2053 407 2067
rect 513 2053 527 2067
rect 613 2053 627 2067
rect 653 2053 667 2067
rect 773 2053 787 2067
rect 813 2053 827 2067
rect 873 2053 887 2067
rect 913 2053 927 2067
rect 1073 2053 1087 2067
rect 1113 2053 1127 2067
rect 1193 2053 1207 2067
rect 1233 2053 1247 2067
rect 1333 2053 1347 2067
rect 1373 2053 1387 2067
rect 1493 2053 1507 2067
rect 1533 2053 1547 2067
rect 1633 2053 1647 2067
rect 1673 2053 1687 2067
rect 1753 2053 1767 2067
rect 1793 2053 1807 2067
rect 1873 2053 1887 2067
rect 1913 2053 1927 2067
rect 2053 2053 2067 2067
rect 2113 2053 2127 2067
rect 2273 2053 2287 2067
rect 2313 2053 2327 2067
rect 2353 2053 2367 2067
rect 2433 2053 2447 2067
rect 2733 2053 2747 2067
rect 2873 2053 2887 2067
rect 2913 2053 2927 2067
rect 3033 2053 3047 2067
rect 3133 2053 3147 2067
rect 3513 2053 3527 2067
rect 3553 2053 3567 2067
rect 3713 2053 3727 2067
rect 3793 2053 3807 2067
rect 3833 2053 3847 2067
rect 3953 2053 3967 2067
rect 4253 2053 4267 2067
rect 4353 2053 4367 2067
rect 4393 2053 4407 2067
rect 4493 2053 4507 2067
rect 4533 2053 4547 2067
rect 4633 2053 4647 2067
rect 4753 2053 4767 2067
rect 4893 2053 4907 2067
rect 4933 2053 4947 2067
rect 5033 2053 5047 2067
rect 5073 2053 5087 2067
rect 5173 2053 5187 2067
rect 5393 2053 5407 2067
rect 5513 2053 5527 2067
rect 5613 2053 5627 2067
rect 5713 2053 5727 2067
rect 5753 2053 5767 2067
rect 233 2033 247 2047
rect 273 2033 287 2047
rect 893 2033 907 2047
rect 933 2033 947 2047
rect 1053 2033 1067 2047
rect 1093 2033 1107 2047
rect 1613 2033 1627 2047
rect 1653 2033 1667 2047
rect 2253 2033 2267 2047
rect 2293 2033 2307 2047
rect 2773 2033 2787 2047
rect 3013 2033 3027 2047
rect 3053 2033 3067 2047
rect 3113 2033 3127 2047
rect 3153 2033 3167 2047
rect 3413 2033 3427 2047
rect 3813 2033 3827 2047
rect 3853 2033 3867 2047
rect 4113 2033 4127 2047
rect 4233 2033 4247 2047
rect 4273 2033 4287 2047
rect 4613 2033 4627 2047
rect 4653 2033 4667 2047
rect 4733 2033 4747 2047
rect 4773 2033 4787 2047
rect 5373 2033 5387 2047
rect 5413 2033 5427 2047
rect 73 1813 87 1827
rect 113 1813 127 1827
rect 493 1813 507 1827
rect 533 1813 547 1827
rect 1853 1813 1867 1827
rect 1893 1813 1907 1827
rect 1973 1813 1987 1827
rect 2013 1813 2027 1827
rect 2613 1813 2627 1827
rect 2693 1813 2707 1827
rect 2733 1813 2747 1827
rect 2833 1813 2847 1827
rect 2873 1813 2887 1827
rect 4093 1813 4107 1827
rect 4133 1813 4147 1827
rect 4373 1813 4387 1827
rect 4413 1813 4427 1827
rect 4653 1813 4667 1827
rect 4893 1813 4907 1827
rect 4933 1813 4947 1827
rect 93 1793 107 1807
rect 133 1793 147 1807
rect 193 1793 207 1807
rect 233 1793 247 1807
rect 353 1793 367 1807
rect 393 1793 407 1807
rect 513 1793 527 1807
rect 553 1793 567 1807
rect 753 1793 767 1807
rect 793 1793 807 1807
rect 933 1793 947 1807
rect 1053 1793 1067 1807
rect 1093 1793 1107 1807
rect 1193 1793 1207 1807
rect 1233 1793 1247 1807
rect 1333 1793 1347 1807
rect 1433 1793 1447 1807
rect 1473 1793 1487 1807
rect 1573 1793 1587 1807
rect 1613 1793 1627 1807
rect 1713 1793 1727 1807
rect 1753 1793 1767 1807
rect 1873 1793 1887 1807
rect 1993 1793 2007 1807
rect 2113 1793 2127 1807
rect 2153 1793 2167 1807
rect 2193 1793 2207 1807
rect 2273 1793 2287 1807
rect 2573 1793 2587 1807
rect 2713 1793 2727 1807
rect 2853 1793 2867 1807
rect 2893 1793 2907 1807
rect 2973 1793 2987 1807
rect 3013 1793 3027 1807
rect 3213 1793 3227 1807
rect 3273 1793 3287 1807
rect 3393 1793 3407 1807
rect 3493 1793 3507 1807
rect 3533 1793 3547 1807
rect 3653 1793 3667 1807
rect 3693 1793 3707 1807
rect 3813 1793 3827 1807
rect 3853 1793 3867 1807
rect 3953 1793 3967 1807
rect 3993 1793 4007 1807
rect 4113 1793 4127 1807
rect 4233 1793 4247 1807
rect 4273 1793 4287 1807
rect 4393 1793 4407 1807
rect 4493 1793 4507 1807
rect 4533 1793 4547 1807
rect 4913 1793 4927 1807
rect 5033 1793 5047 1807
rect 5073 1793 5087 1807
rect 5173 1793 5187 1807
rect 5393 1793 5407 1807
rect 5433 1793 5447 1807
rect 5533 1793 5547 1807
rect 5573 1793 5587 1807
rect 5653 1793 5667 1807
rect 5693 1793 5707 1807
rect 253 1773 267 1787
rect 373 1773 387 1787
rect 413 1773 427 1787
rect 653 1773 667 1787
rect 693 1773 707 1787
rect 813 1773 827 1787
rect 1073 1773 1087 1787
rect 1113 1773 1127 1787
rect 1213 1773 1227 1787
rect 1253 1773 1267 1787
rect 1453 1773 1467 1787
rect 1493 1773 1507 1787
rect 1553 1773 1567 1787
rect 1593 1773 1607 1787
rect 1733 1773 1747 1787
rect 1773 1773 1787 1787
rect 2993 1773 3007 1787
rect 3033 1773 3047 1787
rect 3093 1773 3107 1787
rect 3133 1773 3147 1787
rect 3233 1773 3247 1787
rect 3293 1773 3307 1787
rect 3473 1773 3487 1787
rect 3513 1773 3527 1787
rect 3553 1773 3567 1787
rect 3673 1773 3687 1787
rect 3713 1773 3727 1787
rect 3833 1773 3847 1787
rect 3873 1773 3887 1787
rect 3933 1773 3947 1787
rect 3973 1773 3987 1787
rect 4213 1773 4227 1787
rect 4253 1773 4267 1787
rect 4293 1773 4307 1787
rect 4473 1773 4487 1787
rect 4513 1773 4527 1787
rect 4633 1773 4647 1787
rect 4693 1773 4707 1787
rect 4773 1773 4787 1787
rect 4813 1773 4827 1787
rect 5013 1773 5027 1787
rect 5053 1773 5067 1787
rect 5093 1773 5107 1787
rect 5273 1773 5287 1787
rect 5313 1773 5327 1787
rect 5373 1773 5387 1787
rect 5413 1773 5427 1787
rect 5553 1773 5567 1787
rect 5593 1773 5607 1787
rect 213 1753 227 1767
rect 673 1753 687 1767
rect 773 1753 787 1767
rect 953 1753 967 1767
rect 1353 1753 1367 1767
rect 2453 1753 2467 1767
rect 3113 1753 3127 1767
rect 3413 1753 3427 1767
rect 4793 1753 4807 1767
rect 5193 1753 5207 1767
rect 5293 1753 5307 1767
rect 373 1613 387 1627
rect 553 1613 567 1627
rect 753 1613 767 1627
rect 1293 1613 1307 1627
rect 1573 1613 1587 1627
rect 2033 1613 2047 1627
rect 3233 1613 3247 1627
rect 3633 1613 3647 1627
rect 413 1593 427 1607
rect 513 1593 527 1607
rect 893 1593 907 1607
rect 933 1593 947 1607
rect 1273 1593 1287 1607
rect 1313 1593 1327 1607
rect 1413 1593 1427 1607
rect 1453 1593 1467 1607
rect 1633 1593 1647 1607
rect 1673 1593 1687 1607
rect 1713 1593 1727 1607
rect 2293 1593 2307 1607
rect 2333 1593 2347 1607
rect 2593 1593 2607 1607
rect 2633 1593 2647 1607
rect 2853 1593 2867 1607
rect 2893 1593 2907 1607
rect 2993 1593 3007 1607
rect 3033 1593 3047 1607
rect 3593 1593 3607 1607
rect 3713 1593 3727 1607
rect 3753 1593 3767 1607
rect 3873 1593 3887 1607
rect 3913 1593 3927 1607
rect 3993 1593 4007 1607
rect 4053 1593 4067 1607
rect 4253 1593 4267 1607
rect 4293 1593 4307 1607
rect 4333 1593 4347 1607
rect 4413 1593 4427 1607
rect 4453 1593 4467 1607
rect 4493 1593 4507 1607
rect 4573 1593 4587 1607
rect 4613 1593 4627 1607
rect 4653 1593 4667 1607
rect 4853 1593 4867 1607
rect 4893 1593 4907 1607
rect 5013 1593 5027 1607
rect 5073 1593 5087 1607
rect 5293 1593 5307 1607
rect 5333 1593 5347 1607
rect 5373 1593 5387 1607
rect 5753 1593 5767 1607
rect 73 1573 87 1587
rect 113 1573 127 1587
rect 253 1573 267 1587
rect 293 1573 307 1587
rect 353 1573 367 1587
rect 393 1573 407 1587
rect 533 1573 547 1587
rect 573 1573 587 1587
rect 653 1573 667 1587
rect 773 1573 787 1587
rect 873 1573 887 1587
rect 913 1573 927 1587
rect 1033 1573 1047 1587
rect 1073 1573 1087 1587
rect 1173 1573 1187 1587
rect 1553 1573 1567 1587
rect 1653 1573 1667 1587
rect 1693 1573 1707 1587
rect 1773 1573 1787 1587
rect 1853 1573 1867 1587
rect 2153 1573 2167 1587
rect 2313 1573 2327 1587
rect 2353 1573 2367 1587
rect 2453 1573 2467 1587
rect 2573 1573 2587 1587
rect 2613 1573 2627 1587
rect 2733 1573 2747 1587
rect 2833 1573 2847 1587
rect 2873 1573 2887 1587
rect 2973 1573 2987 1587
rect 3013 1573 3027 1587
rect 3113 1573 3127 1587
rect 3413 1573 3427 1587
rect 3493 1573 3507 1587
rect 3613 1573 3627 1587
rect 3653 1573 3667 1587
rect 3733 1573 3747 1587
rect 3773 1573 3787 1587
rect 4133 1573 4147 1587
rect 4273 1573 4287 1587
rect 4313 1573 4327 1587
rect 4433 1573 4447 1587
rect 4473 1573 4487 1587
rect 4593 1573 4607 1587
rect 4633 1573 4647 1587
rect 4753 1573 4767 1587
rect 4873 1573 4887 1587
rect 4913 1573 4927 1587
rect 5153 1573 5167 1587
rect 5193 1573 5207 1587
rect 5313 1573 5327 1587
rect 5353 1573 5367 1587
rect 5473 1573 5487 1587
rect 5573 1573 5587 1587
rect 5613 1573 5627 1587
rect 5773 1573 5787 1587
rect 93 1553 107 1567
rect 133 1553 147 1567
rect 233 1553 247 1567
rect 273 1553 287 1567
rect 633 1553 647 1567
rect 673 1553 687 1567
rect 1013 1553 1027 1567
rect 1053 1553 1067 1567
rect 1153 1553 1167 1567
rect 1193 1553 1207 1567
rect 2193 1553 2207 1567
rect 2433 1553 2447 1567
rect 2473 1553 2487 1567
rect 2713 1553 2727 1567
rect 2753 1553 2767 1567
rect 3073 1553 3087 1567
rect 4013 1553 4027 1567
rect 4113 1553 4127 1567
rect 4153 1553 4167 1567
rect 4733 1553 4747 1567
rect 4773 1553 4787 1567
rect 5033 1553 5047 1567
rect 5173 1553 5187 1567
rect 5213 1553 5227 1567
rect 5453 1553 5467 1567
rect 5493 1553 5507 1567
rect 5593 1553 5607 1567
rect 5633 1553 5647 1567
rect 73 1333 87 1347
rect 113 1333 127 1347
rect 353 1333 367 1347
rect 393 1333 407 1347
rect 813 1333 827 1347
rect 913 1333 927 1347
rect 953 1333 967 1347
rect 1153 1333 1167 1347
rect 1193 1333 1207 1347
rect 1273 1333 1287 1347
rect 1313 1333 1327 1347
rect 1413 1333 1427 1347
rect 1453 1333 1467 1347
rect 1533 1333 1547 1347
rect 1573 1333 1587 1347
rect 1673 1333 1687 1347
rect 1713 1333 1727 1347
rect 1793 1333 1807 1347
rect 1833 1333 1847 1347
rect 1933 1333 1947 1347
rect 1973 1333 1987 1347
rect 2193 1333 2207 1347
rect 2233 1333 2247 1347
rect 2333 1333 2347 1347
rect 2373 1333 2387 1347
rect 4713 1333 4727 1347
rect 4753 1333 4767 1347
rect 5093 1333 5107 1347
rect 5133 1333 5147 1347
rect 5233 1333 5247 1347
rect 5273 1333 5287 1347
rect 93 1313 107 1327
rect 133 1313 147 1327
rect 193 1313 207 1327
rect 233 1313 247 1327
rect 373 1313 387 1327
rect 413 1313 427 1327
rect 493 1313 507 1327
rect 533 1313 547 1327
rect 633 1313 647 1327
rect 673 1313 687 1327
rect 933 1313 947 1327
rect 1053 1313 1067 1327
rect 1133 1313 1147 1327
rect 1173 1313 1187 1327
rect 1293 1313 1307 1327
rect 1433 1313 1447 1327
rect 1553 1313 1567 1327
rect 1693 1313 1707 1327
rect 1733 1313 1747 1327
rect 1813 1313 1827 1327
rect 1953 1313 1967 1327
rect 1993 1313 2007 1327
rect 2073 1313 2087 1327
rect 2213 1313 2227 1327
rect 2253 1313 2267 1327
rect 2353 1313 2367 1327
rect 2393 1313 2407 1327
rect 2473 1313 2487 1327
rect 2593 1313 2607 1327
rect 2633 1313 2647 1327
rect 2713 1313 2727 1327
rect 2753 1313 2767 1327
rect 2873 1313 2887 1327
rect 2913 1313 2927 1327
rect 3013 1313 3027 1327
rect 3053 1313 3067 1327
rect 3153 1313 3167 1327
rect 3193 1313 3207 1327
rect 3293 1313 3307 1327
rect 3393 1313 3407 1327
rect 3653 1313 3667 1327
rect 3693 1313 3707 1327
rect 3773 1313 3787 1327
rect 3813 1313 3827 1327
rect 3913 1313 3927 1327
rect 4013 1313 4027 1327
rect 4053 1313 4067 1327
rect 4153 1313 4167 1327
rect 4193 1313 4207 1327
rect 4313 1313 4327 1327
rect 4353 1313 4367 1327
rect 4433 1313 4447 1327
rect 4473 1313 4487 1327
rect 4593 1313 4607 1327
rect 4633 1313 4647 1327
rect 4733 1313 4747 1327
rect 4853 1313 4867 1327
rect 4893 1313 4907 1327
rect 5113 1313 5127 1327
rect 5253 1313 5267 1327
rect 5353 1313 5367 1327
rect 5393 1313 5407 1327
rect 5493 1313 5507 1327
rect 5533 1313 5547 1327
rect 5653 1313 5667 1327
rect 5693 1313 5707 1327
rect 253 1293 267 1307
rect 513 1293 527 1307
rect 553 1293 567 1307
rect 653 1293 667 1307
rect 693 1293 707 1307
rect 793 1293 807 1307
rect 853 1293 867 1307
rect 2613 1293 2627 1307
rect 2653 1293 2667 1307
rect 2773 1293 2787 1307
rect 2893 1293 2907 1307
rect 2933 1293 2947 1307
rect 3033 1293 3047 1307
rect 3073 1293 3087 1307
rect 3173 1293 3187 1307
rect 3213 1293 3227 1307
rect 3493 1293 3507 1307
rect 3533 1293 3547 1307
rect 3633 1293 3647 1307
rect 3753 1293 3767 1307
rect 3793 1293 3807 1307
rect 4033 1293 4047 1307
rect 4073 1293 4087 1307
rect 4173 1293 4187 1307
rect 4213 1293 4227 1307
rect 4293 1293 4307 1307
rect 4453 1293 4467 1307
rect 4493 1293 4507 1307
rect 4573 1293 4587 1307
rect 4613 1293 4627 1307
rect 4833 1293 4847 1307
rect 4873 1293 4887 1307
rect 4973 1293 4987 1307
rect 5013 1293 5027 1307
rect 5373 1293 5387 1307
rect 5413 1293 5427 1307
rect 5473 1293 5487 1307
rect 5513 1293 5527 1307
rect 5633 1293 5647 1307
rect 5673 1293 5687 1307
rect 213 1273 227 1287
rect 1073 1273 1087 1287
rect 2093 1273 2107 1287
rect 2453 1273 2467 1287
rect 2733 1273 2747 1287
rect 3313 1273 3327 1287
rect 3373 1273 3387 1287
rect 3673 1273 3687 1287
rect 3933 1273 3947 1287
rect 4333 1273 4347 1287
rect 4993 1273 5007 1287
rect 93 1133 107 1147
rect 173 1133 187 1147
rect 893 1133 907 1147
rect 1193 1133 1207 1147
rect 1273 1133 1287 1147
rect 1433 1133 1447 1147
rect 1533 1133 1547 1147
rect 1633 1133 1647 1147
rect 2713 1133 2727 1147
rect 2833 1133 2847 1147
rect 2953 1133 2967 1147
rect 3233 1133 3247 1147
rect 3373 1133 3387 1147
rect 3493 1133 3507 1147
rect 4093 1133 4107 1147
rect 4193 1133 4207 1147
rect 4353 1133 4367 1147
rect 4653 1133 4667 1147
rect 4993 1133 5007 1147
rect 5093 1133 5107 1147
rect 5493 1133 5507 1147
rect 5773 1133 5787 1147
rect 213 1113 227 1127
rect 293 1113 307 1127
rect 333 1113 347 1127
rect 433 1113 447 1127
rect 473 1113 487 1127
rect 713 1113 727 1127
rect 753 1113 767 1127
rect 933 1113 947 1127
rect 1053 1113 1067 1127
rect 1093 1113 1107 1127
rect 1313 1113 1327 1127
rect 1513 1113 1527 1127
rect 1553 1113 1567 1127
rect 2033 1113 2047 1127
rect 2073 1113 2087 1127
rect 2453 1113 2467 1127
rect 2493 1113 2507 1127
rect 2813 1113 2827 1127
rect 2853 1113 2867 1127
rect 2933 1113 2947 1127
rect 2973 1113 2987 1127
rect 3053 1113 3067 1127
rect 3113 1113 3127 1127
rect 3213 1113 3227 1127
rect 3253 1113 3267 1127
rect 3353 1113 3367 1127
rect 3393 1113 3407 1127
rect 3593 1113 3607 1127
rect 3633 1113 3647 1127
rect 3733 1113 3747 1127
rect 3773 1113 3787 1127
rect 4073 1113 4087 1127
rect 4113 1113 4127 1127
rect 4313 1113 4327 1127
rect 4493 1113 4507 1127
rect 4533 1113 4547 1127
rect 4613 1113 4627 1127
rect 4733 1113 4747 1127
rect 4773 1113 4787 1127
rect 4873 1113 4887 1127
rect 4913 1113 4927 1127
rect 5373 1113 5387 1127
rect 5413 1113 5427 1127
rect 5473 1113 5487 1127
rect 5513 1113 5527 1127
rect 73 1093 87 1107
rect 153 1093 167 1107
rect 193 1093 207 1107
rect 313 1093 327 1107
rect 353 1093 367 1107
rect 453 1093 467 1107
rect 493 1093 507 1107
rect 613 1093 627 1107
rect 653 1093 667 1107
rect 733 1093 747 1107
rect 773 1093 787 1107
rect 873 1093 887 1107
rect 913 1093 927 1107
rect 1033 1093 1047 1107
rect 1073 1093 1087 1107
rect 1173 1093 1187 1107
rect 1253 1093 1267 1107
rect 1293 1093 1307 1107
rect 1413 1093 1427 1107
rect 1653 1093 1667 1107
rect 1773 1093 1787 1107
rect 1813 1093 1827 1107
rect 1913 1093 1927 1107
rect 2013 1093 2027 1107
rect 2053 1093 2067 1107
rect 2173 1093 2187 1107
rect 2213 1093 2227 1107
rect 2313 1093 2327 1107
rect 2353 1093 2367 1107
rect 2433 1093 2447 1107
rect 2473 1093 2487 1107
rect 2593 1093 2607 1107
rect 2633 1093 2647 1107
rect 2733 1093 2747 1107
rect 3473 1093 3487 1107
rect 3573 1093 3587 1107
rect 3613 1093 3627 1107
rect 3713 1093 3727 1107
rect 3753 1093 3767 1107
rect 3853 1093 3867 1107
rect 3973 1093 3987 1107
rect 4213 1093 4227 1107
rect 4333 1093 4347 1107
rect 4373 1093 4387 1107
rect 4473 1093 4487 1107
rect 4513 1093 4527 1107
rect 4633 1093 4647 1107
rect 4673 1093 4687 1107
rect 4753 1093 4767 1107
rect 4793 1093 4807 1107
rect 5013 1093 5027 1107
rect 5113 1093 5127 1107
rect 5233 1093 5247 1107
rect 5353 1093 5367 1107
rect 5393 1093 5407 1107
rect 5633 1093 5647 1107
rect 5673 1093 5687 1107
rect 5753 1093 5767 1107
rect 593 1073 607 1087
rect 633 1073 647 1087
rect 1753 1073 1767 1087
rect 1793 1073 1807 1087
rect 1893 1073 1907 1087
rect 1933 1073 1947 1087
rect 2153 1073 2167 1087
rect 2193 1073 2207 1087
rect 2293 1073 2307 1087
rect 2333 1073 2347 1087
rect 2573 1073 2587 1087
rect 2613 1073 2627 1087
rect 3093 1073 3107 1087
rect 3833 1073 3847 1087
rect 3873 1073 3887 1087
rect 3953 1073 3967 1087
rect 3993 1073 4007 1087
rect 5213 1073 5227 1087
rect 5253 1073 5267 1087
rect 5613 1073 5627 1087
rect 5653 1073 5667 1087
rect 73 853 87 867
rect 113 853 127 867
rect 353 853 367 867
rect 393 853 407 867
rect 633 853 647 867
rect 673 853 687 867
rect 1053 853 1067 867
rect 1093 853 1107 867
rect 1333 853 1347 867
rect 1373 853 1387 867
rect 1553 853 1567 867
rect 1593 853 1607 867
rect 1713 853 1727 867
rect 1753 853 1767 867
rect 1853 853 1867 867
rect 1893 853 1907 867
rect 1993 853 2007 867
rect 2033 853 2047 867
rect 2293 853 2307 867
rect 2513 853 2527 867
rect 2553 853 2567 867
rect 2753 853 2767 867
rect 2793 853 2807 867
rect 2893 853 2907 867
rect 2933 853 2947 867
rect 3253 853 3267 867
rect 3293 853 3307 867
rect 3993 853 4007 867
rect 4033 853 4047 867
rect 93 833 107 847
rect 133 833 147 847
rect 193 833 207 847
rect 233 833 247 847
rect 373 833 387 847
rect 413 833 427 847
rect 513 833 527 847
rect 553 833 567 847
rect 653 833 667 847
rect 693 833 707 847
rect 753 833 767 847
rect 793 833 807 847
rect 913 833 927 847
rect 953 833 967 847
rect 1073 833 1087 847
rect 1113 833 1127 847
rect 1193 833 1207 847
rect 1233 833 1247 847
rect 1353 833 1367 847
rect 1393 833 1407 847
rect 1473 833 1487 847
rect 1573 833 1587 847
rect 1733 833 1747 847
rect 1773 833 1787 847
rect 1873 833 1887 847
rect 1913 833 1927 847
rect 1973 833 1987 847
rect 2013 833 2027 847
rect 2133 833 2147 847
rect 2173 833 2187 847
rect 2413 833 2427 847
rect 2533 833 2547 847
rect 2633 833 2647 847
rect 2773 833 2787 847
rect 2913 833 2927 847
rect 3033 833 3047 847
rect 3133 833 3147 847
rect 3273 833 3287 847
rect 3653 833 3667 847
rect 3693 833 3707 847
rect 3773 833 3787 847
rect 3873 833 3887 847
rect 3913 833 3927 847
rect 4013 833 4027 847
rect 4133 833 4147 847
rect 4173 833 4187 847
rect 4273 833 4287 847
rect 4313 833 4327 847
rect 4433 833 4447 847
rect 4533 833 4547 847
rect 4573 833 4587 847
rect 4653 833 4667 847
rect 4693 833 4707 847
rect 4933 833 4947 847
rect 4973 833 4987 847
rect 5053 833 5067 847
rect 5093 833 5107 847
rect 5213 833 5227 847
rect 5373 833 5387 847
rect 5493 833 5507 847
rect 5533 833 5547 847
rect 5653 833 5667 847
rect 5693 833 5707 847
rect 253 813 267 827
rect 493 813 507 827
rect 813 813 827 827
rect 933 813 947 827
rect 973 813 987 827
rect 1173 813 1187 827
rect 1213 813 1227 827
rect 2113 813 2127 827
rect 2153 813 2167 827
rect 2253 813 2267 827
rect 2313 813 2327 827
rect 2673 813 2687 827
rect 3393 813 3407 827
rect 3433 813 3447 827
rect 3513 813 3527 827
rect 3553 813 3567 827
rect 3633 813 3647 827
rect 3893 813 3907 827
rect 3933 813 3947 827
rect 4153 813 4167 827
rect 4193 813 4207 827
rect 4293 813 4307 827
rect 4333 813 4347 827
rect 4553 813 4567 827
rect 4593 813 4607 827
rect 4713 813 4727 827
rect 4813 813 4827 827
rect 4853 813 4867 827
rect 4953 813 4967 827
rect 4993 813 5007 827
rect 5113 813 5127 827
rect 5253 813 5267 827
rect 5473 813 5487 827
rect 5513 813 5527 827
rect 5553 813 5567 827
rect 5633 813 5647 827
rect 5673 813 5687 827
rect 213 793 227 807
rect 533 793 547 807
rect 773 793 787 807
rect 1453 793 1467 807
rect 2393 793 2407 807
rect 2693 793 2707 807
rect 3013 793 3027 807
rect 3153 793 3167 807
rect 3413 793 3427 807
rect 3533 793 3547 807
rect 3673 793 3687 807
rect 3793 793 3807 807
rect 4413 793 4427 807
rect 4673 793 4687 807
rect 5073 793 5087 807
rect 5273 793 5287 807
rect 5393 793 5407 807
rect 273 653 287 667
rect 653 653 667 667
rect 1213 653 1227 667
rect 1393 653 1407 667
rect 1933 653 1947 667
rect 2093 653 2107 667
rect 2253 653 2267 667
rect 2733 653 2747 667
rect 3093 653 3107 667
rect 4033 653 4047 667
rect 4353 653 4367 667
rect 4473 653 4487 667
rect 4993 653 5007 667
rect 5673 653 5687 667
rect 233 633 247 647
rect 533 633 547 647
rect 573 633 587 647
rect 693 633 707 647
rect 953 633 967 647
rect 993 633 1007 647
rect 1253 633 1267 647
rect 1353 633 1367 647
rect 1673 633 1687 647
rect 1713 633 1727 647
rect 1973 633 1987 647
rect 2073 633 2087 647
rect 2113 633 2127 647
rect 2233 633 2247 647
rect 2313 633 2327 647
rect 2373 633 2387 647
rect 2713 633 2727 647
rect 2753 633 2767 647
rect 2813 633 2827 647
rect 2853 633 2867 647
rect 3133 633 3147 647
rect 3513 633 3527 647
rect 3553 633 3567 647
rect 3773 633 3787 647
rect 3813 633 3827 647
rect 3873 633 3887 647
rect 3913 633 3927 647
rect 4073 633 4087 647
rect 4173 633 4187 647
rect 4213 633 4227 647
rect 4433 633 4447 647
rect 4593 633 4607 647
rect 4633 633 4647 647
rect 4733 633 4747 647
rect 4773 633 4787 647
rect 4853 633 4867 647
rect 4893 633 4907 647
rect 5113 633 5127 647
rect 5153 633 5167 647
rect 5273 633 5287 647
rect 5313 633 5327 647
rect 5373 633 5387 647
rect 5413 633 5427 647
rect 5553 633 5567 647
rect 5593 633 5607 647
rect 5653 633 5667 647
rect 5693 633 5707 647
rect 93 613 107 627
rect 133 613 147 627
rect 253 613 267 627
rect 293 613 307 627
rect 393 613 407 627
rect 433 613 447 627
rect 513 613 527 627
rect 553 613 567 627
rect 633 613 647 627
rect 673 613 687 627
rect 793 613 807 627
rect 933 613 947 627
rect 973 613 987 627
rect 1093 613 1107 627
rect 1133 613 1147 627
rect 1193 613 1207 627
rect 1233 613 1247 627
rect 1373 613 1387 627
rect 1413 613 1427 627
rect 1493 613 1507 627
rect 1533 613 1547 627
rect 1653 613 1667 627
rect 1693 613 1707 627
rect 1813 613 1827 627
rect 1853 613 1867 627
rect 1913 613 1927 627
rect 1953 613 1967 627
rect 2193 613 2207 627
rect 2473 613 2487 627
rect 2613 613 2627 627
rect 2833 613 2847 627
rect 2873 613 2887 627
rect 2993 613 3007 627
rect 3073 613 3087 627
rect 3113 613 3127 627
rect 3253 613 3267 627
rect 3293 613 3307 627
rect 3373 613 3387 627
rect 3493 613 3507 627
rect 3533 613 3547 627
rect 3633 613 3647 627
rect 3753 613 3767 627
rect 3793 613 3807 627
rect 3893 613 3907 627
rect 3933 613 3947 627
rect 4013 613 4027 627
rect 4053 613 4067 627
rect 4193 613 4207 627
rect 4233 613 4247 627
rect 4333 613 4347 627
rect 4453 613 4467 627
rect 4493 613 4507 627
rect 4573 613 4587 627
rect 4613 613 4627 627
rect 4713 613 4727 627
rect 4753 613 4767 627
rect 4873 613 4887 627
rect 4913 613 4927 627
rect 5013 613 5027 627
rect 5253 613 5267 627
rect 5293 613 5307 627
rect 5393 613 5407 627
rect 5433 613 5447 627
rect 5533 613 5547 627
rect 5573 613 5587 627
rect 73 593 87 607
rect 113 593 127 607
rect 373 593 387 607
rect 413 593 427 607
rect 773 593 787 607
rect 813 593 827 607
rect 1073 593 1087 607
rect 1113 593 1127 607
rect 1513 593 1527 607
rect 1553 593 1567 607
rect 1793 593 1807 607
rect 1833 593 1847 607
rect 2353 593 2367 607
rect 2453 593 2467 607
rect 2493 593 2507 607
rect 2593 593 2607 607
rect 2633 593 2647 607
rect 2973 593 2987 607
rect 3013 593 3027 607
rect 3233 593 3247 607
rect 3273 593 3287 607
rect 3353 593 3367 607
rect 3393 593 3407 607
rect 3613 593 3627 607
rect 3653 593 3667 607
rect 73 373 87 387
rect 113 373 127 387
rect 513 373 527 387
rect 553 373 567 387
rect 673 373 687 387
rect 793 373 807 387
rect 833 373 847 387
rect 1073 373 1087 387
rect 1113 373 1127 387
rect 1353 373 1367 387
rect 1393 373 1407 387
rect 1773 373 1787 387
rect 2513 373 2527 387
rect 2553 373 2567 387
rect 3813 373 3827 387
rect 3853 373 3867 387
rect 3933 373 3947 387
rect 3973 373 3987 387
rect 4093 373 4107 387
rect 4133 373 4147 387
rect 4473 373 4487 387
rect 4513 373 4527 387
rect 5713 373 5727 387
rect 5753 373 5767 387
rect 93 353 107 367
rect 133 353 147 367
rect 213 353 227 367
rect 253 353 267 367
rect 373 353 387 367
rect 413 353 427 367
rect 533 353 547 367
rect 573 353 587 367
rect 813 353 827 367
rect 853 353 867 367
rect 953 353 967 367
rect 993 353 1007 367
rect 1053 353 1067 367
rect 1093 353 1107 367
rect 1213 353 1227 367
rect 1373 353 1387 367
rect 1413 353 1427 367
rect 1513 353 1527 367
rect 1613 353 1627 367
rect 1653 353 1667 367
rect 2033 353 2047 367
rect 2133 353 2147 367
rect 2173 353 2187 367
rect 2293 353 2307 367
rect 2333 353 2347 367
rect 2413 353 2427 367
rect 2533 353 2547 367
rect 2573 353 2587 367
rect 2653 353 2667 367
rect 2693 353 2707 367
rect 2793 353 2807 367
rect 3013 353 3027 367
rect 3133 353 3147 367
rect 3173 353 3187 367
rect 3253 353 3267 367
rect 3293 353 3307 367
rect 3413 353 3427 367
rect 3533 353 3547 367
rect 3573 353 3587 367
rect 3653 353 3667 367
rect 3693 353 3707 367
rect 3833 353 3847 367
rect 3873 353 3887 367
rect 3953 353 3967 367
rect 4113 353 4127 367
rect 4153 353 4167 367
rect 4233 353 4247 367
rect 4273 353 4287 367
rect 4373 353 4387 367
rect 4493 353 4507 367
rect 4593 353 4607 367
rect 4633 353 4647 367
rect 4733 353 4747 367
rect 4833 353 4847 367
rect 4873 353 4887 367
rect 4953 353 4967 367
rect 5013 353 5027 367
rect 5133 353 5147 367
rect 5173 353 5187 367
rect 5293 353 5307 367
rect 5333 353 5347 367
rect 5473 353 5487 367
rect 5513 353 5527 367
rect 5593 353 5607 367
rect 5633 353 5647 367
rect 5733 353 5747 367
rect 233 333 247 347
rect 273 333 287 347
rect 393 333 407 347
rect 433 333 447 347
rect 653 333 667 347
rect 713 333 727 347
rect 933 333 947 347
rect 1253 333 1267 347
rect 1633 333 1647 347
rect 1673 333 1687 347
rect 1753 333 1767 347
rect 1813 333 1827 347
rect 1873 333 1887 347
rect 1913 333 1927 347
rect 2153 333 2167 347
rect 2193 333 2207 347
rect 2273 333 2287 347
rect 2633 333 2647 347
rect 2673 333 2687 347
rect 2893 333 2907 347
rect 2933 333 2947 347
rect 3113 333 3127 347
rect 3313 333 3327 347
rect 3513 333 3527 347
rect 3553 333 3567 347
rect 3713 333 3727 347
rect 4253 333 4267 347
rect 4293 333 4307 347
rect 4613 333 4627 347
rect 4653 333 4667 347
rect 4853 333 4867 347
rect 4893 333 4907 347
rect 4973 333 4987 347
rect 5033 333 5047 347
rect 5153 333 5167 347
rect 5193 333 5207 347
rect 5273 333 5287 347
rect 5313 333 5327 347
rect 5453 333 5467 347
rect 5573 333 5587 347
rect 5613 333 5627 347
rect 973 313 987 327
rect 1273 313 1287 327
rect 1533 313 1547 327
rect 1893 313 1907 327
rect 2013 313 2027 327
rect 2313 313 2327 327
rect 2433 313 2447 327
rect 2813 313 2827 327
rect 2913 313 2927 327
rect 2993 313 3007 327
rect 3153 313 3167 327
rect 3273 313 3287 327
rect 3433 313 3447 327
rect 3673 313 3687 327
rect 4393 313 4407 327
rect 4753 313 4767 327
rect 5493 313 5507 327
rect 213 173 227 187
rect 413 173 427 187
rect 913 173 927 187
rect 1173 173 1187 187
rect 1313 173 1327 187
rect 1593 173 1607 187
rect 2653 173 2667 187
rect 3313 173 3327 187
rect 3553 173 3567 187
rect 4313 173 4327 187
rect 5093 173 5107 187
rect 5473 173 5487 187
rect 5613 173 5627 187
rect 253 153 267 167
rect 373 153 387 167
rect 533 153 547 167
rect 573 153 587 167
rect 633 153 647 167
rect 673 153 687 167
rect 1013 153 1027 167
rect 1053 153 1067 167
rect 1213 153 1227 167
rect 1293 153 1307 167
rect 1333 153 1347 167
rect 1413 153 1427 167
rect 1473 153 1487 167
rect 1693 153 1707 167
rect 1733 153 1747 167
rect 2213 153 2227 167
rect 2253 153 2267 167
rect 2453 153 2467 167
rect 2513 153 2527 167
rect 2613 153 2627 167
rect 2753 153 2767 167
rect 2813 153 2827 167
rect 3373 153 3387 167
rect 3413 153 3427 167
rect 3753 153 3767 167
rect 3793 153 3807 167
rect 3853 153 3867 167
rect 3893 153 3907 167
rect 4113 153 4127 167
rect 4173 153 4187 167
rect 4293 153 4307 167
rect 4333 153 4347 167
rect 4713 153 4727 167
rect 4753 153 4767 167
rect 4973 153 4987 167
rect 5013 153 5027 167
rect 5073 153 5087 167
rect 5113 153 5127 167
rect 5333 153 5347 167
rect 5393 153 5407 167
rect 93 133 107 147
rect 133 133 147 147
rect 193 133 207 147
rect 233 133 247 147
rect 393 133 407 147
rect 433 133 447 147
rect 513 133 527 147
rect 553 133 567 147
rect 653 133 667 147
rect 693 133 707 147
rect 813 133 827 147
rect 853 133 867 147
rect 933 133 947 147
rect 1033 133 1047 147
rect 1073 133 1087 147
rect 1153 133 1167 147
rect 1193 133 1207 147
rect 1573 133 1587 147
rect 1673 133 1687 147
rect 1713 133 1727 147
rect 1833 133 1847 147
rect 1913 133 1927 147
rect 1953 133 1967 147
rect 2113 133 2127 147
rect 2153 133 2167 147
rect 2373 133 2387 147
rect 2633 133 2647 147
rect 2673 133 2687 147
rect 2913 133 2927 147
rect 3053 133 3067 147
rect 3173 133 3187 147
rect 3213 133 3227 147
rect 3293 133 3307 147
rect 3393 133 3407 147
rect 3433 133 3447 147
rect 3533 133 3547 147
rect 3653 133 3667 147
rect 4013 133 4027 147
rect 4413 133 4427 147
rect 4553 133 4567 147
rect 4593 133 4607 147
rect 4693 133 4707 147
rect 4733 133 4747 147
rect 4833 133 4847 147
rect 4953 133 4967 147
rect 4993 133 5007 147
rect 5233 133 5247 147
rect 5313 133 5327 147
rect 5373 133 5387 147
rect 5493 133 5507 147
rect 5593 133 5607 147
rect 5693 133 5707 147
rect 73 113 87 127
rect 113 113 127 127
rect 793 113 807 127
rect 833 113 847 127
rect 1453 113 1467 127
rect 1813 113 1827 127
rect 1853 113 1867 127
rect 1933 113 1947 127
rect 1973 113 1987 127
rect 2093 113 2107 127
rect 2133 113 2147 127
rect 2353 113 2367 127
rect 2393 113 2407 127
rect 2493 113 2507 127
rect 2773 113 2787 127
rect 2893 113 2907 127
rect 2933 113 2947 127
rect 3033 113 3047 127
rect 3073 113 3087 127
rect 3153 113 3167 127
rect 3193 113 3207 127
rect 3633 113 3647 127
rect 3673 113 3687 127
rect 3993 113 4007 127
rect 4033 113 4047 127
rect 4153 113 4167 127
rect 4393 113 4407 127
rect 4433 113 4447 127
rect 4533 113 4547 127
rect 4573 113 4587 127
rect 4813 113 4827 127
rect 4853 113 4867 127
rect 5213 113 5227 127
rect 5253 113 5267 127
rect 5673 113 5687 127
rect 5713 113 5727 127
<< labels >>
flabel metal1 s 5822 2 5882 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 5737 5817 5743 5823 3 FreeSans 16 90 0 0 ABCmd_i[7]
port 2 nsew
flabel metal2 s 5697 5817 5703 5823 3 FreeSans 16 90 0 0 ABCmd_i[6]
port 3 nsew
flabel metal2 s 5637 5817 5643 5823 3 FreeSans 16 90 0 0 ABCmd_i[5]
port 4 nsew
flabel metal2 s 5597 5817 5603 5823 3 FreeSans 16 90 0 0 ABCmd_i[4]
port 5 nsew
flabel metal2 s 5557 5817 5563 5823 3 FreeSans 16 90 0 0 ABCmd_i[3]
port 6 nsew
flabel metal3 s 5856 2776 5864 2784 3 FreeSans 16 0 0 0 ABCmd_i[2]
port 7 nsew
flabel metal3 s 5856 5636 5864 5644 3 FreeSans 16 0 0 0 ABCmd_i[1]
port 8 nsew
flabel metal3 s 5856 5676 5864 5684 3 FreeSans 16 0 0 0 ABCmd_i[0]
port 9 nsew
flabel metal2 s 3897 -23 3903 -17 7 FreeSans 16 270 0 0 ACC_o[7]
port 10 nsew
flabel metal2 s 3857 -23 3863 -17 7 FreeSans 16 270 0 0 ACC_o[6]
port 11 nsew
flabel metal2 s 3757 -23 3763 -17 7 FreeSans 16 270 0 0 ACC_o[5]
port 12 nsew
flabel metal2 s 3497 -23 3503 -17 7 FreeSans 16 270 0 0 ACC_o[4]
port 13 nsew
flabel metal2 s 2677 -23 2683 -17 7 FreeSans 16 270 0 0 ACC_o[3]
port 14 nsew
flabel metal3 s -24 2296 -16 2304 7 FreeSans 16 0 0 0 ACC_o[2]
port 15 nsew
flabel metal3 s -24 2256 -16 2264 7 FreeSans 16 0 0 0 ACC_o[1]
port 16 nsew
flabel metal3 s -24 1556 -16 1564 7 FreeSans 16 0 0 0 ACC_o[0]
port 17 nsew
flabel metal2 s 2637 -23 2643 -17 7 FreeSans 16 270 0 0 Flag_i
port 18 nsew
flabel metal2 s 5197 5817 5203 5823 3 FreeSans 16 90 0 0 LoadA_i
port 19 nsew
flabel metal2 s 5237 5817 5243 5823 3 FreeSans 16 90 0 0 LoadB_i
port 20 nsew
flabel metal2 s 5517 5817 5523 5823 3 FreeSans 16 90 0 0 LoadCmd_i
port 21 nsew
flabel metal3 s -24 3016 -16 3024 7 FreeSans 16 0 0 0 MulH_i
port 22 nsew
flabel metal3 s -24 3476 -16 3484 7 FreeSans 16 0 0 0 MulL_i
port 23 nsew
flabel metal2 s 4717 5817 4723 5823 3 FreeSans 16 90 0 0 clk
port 24 nsew
flabel metal3 s 5856 1796 5864 1804 3 FreeSans 16 0 0 0 reset
port 25 nsew
rlabel nsubstratencontact 44 488 44 488 0 FILL_1__1036_.vdd
rlabel metal1 24 242 56 258 0 FILL_1__1036_.gnd
rlabel nsubstratencontact 44 12 44 12 0 FILL_1__1014_.vdd
rlabel metal1 24 242 56 258 0 FILL_1__1014_.gnd
rlabel nsubstratencontact 24 488 24 488 0 FILL_0__1036_.vdd
rlabel metal1 4 242 36 258 0 FILL_0__1036_.gnd
rlabel nsubstratencontact 24 12 24 12 0 FILL_0__1014_.vdd
rlabel metal1 4 242 36 258 0 FILL_0__1014_.gnd
rlabel metal1 44 242 156 258 0 _1036_.gnd
rlabel metal1 44 482 156 498 0 _1036_.vdd
rlabel metal2 133 353 147 367 0 _1036_.A
rlabel metal2 113 373 127 387 0 _1036_.B
rlabel metal2 93 353 107 367 0 _1036_.C
rlabel metal2 73 373 87 387 0 _1036_.Y
rlabel metal1 44 242 156 258 0 _1014_.gnd
rlabel metal1 44 2 156 18 0 _1014_.vdd
rlabel metal2 133 133 147 147 0 _1014_.A
rlabel metal2 113 113 127 127 0 _1014_.B
rlabel metal2 93 133 107 147 0 _1014_.C
rlabel metal2 73 113 87 127 0 _1014_.Y
rlabel nsubstratencontact 184 488 184 488 0 FILL_1__1032_.vdd
rlabel metal1 164 242 196 258 0 FILL_1__1032_.gnd
rlabel nsubstratencontact 176 12 176 12 0 FILL_1__1029_.vdd
rlabel metal1 164 242 196 258 0 FILL_1__1029_.gnd
rlabel nsubstratencontact 164 488 164 488 0 FILL_0__1032_.vdd
rlabel metal1 144 242 176 258 0 FILL_0__1032_.gnd
rlabel nsubstratencontact 156 12 156 12 0 FILL_0__1029_.vdd
rlabel metal1 144 242 176 258 0 FILL_0__1029_.gnd
rlabel metal1 184 242 296 258 0 _1032_.gnd
rlabel metal1 184 482 296 498 0 _1032_.vdd
rlabel metal2 273 333 287 347 0 _1032_.A
rlabel metal2 253 353 267 367 0 _1032_.B
rlabel metal2 213 353 227 367 0 _1032_.C
rlabel metal2 233 333 247 347 0 _1032_.Y
rlabel metal1 184 242 296 258 0 _1029_.gnd
rlabel metal1 184 2 296 18 0 _1029_.vdd
rlabel metal2 193 133 207 147 0 _1029_.A
rlabel metal2 213 173 227 187 0 _1029_.B
rlabel metal2 233 133 247 147 0 _1029_.C
rlabel metal2 253 153 267 167 0 _1029_.Y
rlabel nsubstratencontact 344 488 344 488 0 FILL_2__1056_.vdd
rlabel metal1 324 242 356 258 0 FILL_2__1056_.gnd
rlabel nsubstratencontact 344 12 344 12 0 FILL_2__1030_.vdd
rlabel metal1 324 242 356 258 0 FILL_2__1030_.gnd
rlabel nsubstratencontact 324 488 324 488 0 FILL_1__1056_.vdd
rlabel metal1 304 242 336 258 0 FILL_1__1056_.gnd
rlabel nsubstratencontact 324 12 324 12 0 FILL_1__1030_.vdd
rlabel metal1 304 242 336 258 0 FILL_1__1030_.gnd
rlabel nsubstratencontact 304 488 304 488 0 FILL_0__1056_.vdd
rlabel metal1 284 242 316 258 0 FILL_0__1056_.gnd
rlabel nsubstratencontact 304 12 304 12 0 FILL_0__1030_.vdd
rlabel metal1 284 242 316 258 0 FILL_0__1030_.gnd
rlabel metal1 344 242 456 258 0 _1056_.gnd
rlabel metal1 344 482 456 498 0 _1056_.vdd
rlabel metal2 433 333 447 347 0 _1056_.A
rlabel metal2 413 353 427 367 0 _1056_.B
rlabel metal2 373 353 387 367 0 _1056_.C
rlabel metal2 393 333 407 347 0 _1056_.Y
rlabel metal1 344 242 456 258 0 _1030_.gnd
rlabel metal1 344 2 456 18 0 _1030_.vdd
rlabel metal2 433 133 447 147 0 _1030_.A
rlabel metal2 413 173 427 187 0 _1030_.B
rlabel metal2 393 133 407 147 0 _1030_.C
rlabel metal2 373 153 387 167 0 _1030_.Y
rlabel nsubstratencontact 484 12 484 12 0 FILL_1__1013_.vdd
rlabel metal1 464 242 496 258 0 FILL_1__1013_.gnd
rlabel nsubstratencontact 484 488 484 488 0 FILL_1__1010_.vdd
rlabel metal1 464 242 496 258 0 FILL_1__1010_.gnd
rlabel nsubstratencontact 464 12 464 12 0 FILL_0__1013_.vdd
rlabel metal1 444 242 476 258 0 FILL_0__1013_.gnd
rlabel nsubstratencontact 464 488 464 488 0 FILL_0__1010_.vdd
rlabel metal1 444 242 476 258 0 FILL_0__1010_.gnd
rlabel metal1 484 242 596 258 0 _1013_.gnd
rlabel metal1 484 2 596 18 0 _1013_.vdd
rlabel metal2 573 153 587 167 0 _1013_.A
rlabel metal2 553 133 567 147 0 _1013_.B
rlabel metal2 513 133 527 147 0 _1013_.C
rlabel metal2 533 153 547 167 0 _1013_.Y
rlabel metal1 484 242 596 258 0 _1010_.gnd
rlabel metal1 484 482 596 498 0 _1010_.vdd
rlabel metal2 573 353 587 367 0 _1010_.A
rlabel metal2 553 373 567 387 0 _1010_.B
rlabel metal2 533 353 547 367 0 _1010_.C
rlabel metal2 513 373 527 387 0 _1010_.Y
rlabel nsubstratencontact 624 488 624 488 0 FILL_1__1031_.vdd
rlabel metal1 604 242 636 258 0 FILL_1__1031_.gnd
rlabel nsubstratencontact 616 12 616 12 0 FILL_1__1006_.vdd
rlabel metal1 604 242 636 258 0 FILL_1__1006_.gnd
rlabel nsubstratencontact 604 488 604 488 0 FILL_0__1031_.vdd
rlabel metal1 584 242 616 258 0 FILL_0__1031_.gnd
rlabel nsubstratencontact 596 12 596 12 0 FILL_0__1006_.vdd
rlabel metal1 584 242 616 258 0 FILL_0__1006_.gnd
rlabel metal1 624 242 736 258 0 _1031_.gnd
rlabel metal1 624 482 736 498 0 _1031_.vdd
rlabel metal2 713 333 727 347 0 _1031_.A
rlabel metal2 653 333 667 347 0 _1031_.Y
rlabel metal2 673 373 687 387 0 _1031_.B
rlabel metal1 624 242 736 258 0 _1006_.gnd
rlabel metal1 624 2 736 18 0 _1006_.vdd
rlabel metal2 633 153 647 167 0 _1006_.A
rlabel metal2 653 133 667 147 0 _1006_.B
rlabel metal2 693 133 707 147 0 _1006_.C
rlabel metal2 673 153 687 167 0 _1006_.Y
rlabel nsubstratencontact 764 12 764 12 0 FILL_1__1012_.vdd
rlabel metal1 744 242 776 258 0 FILL_1__1012_.gnd
rlabel nsubstratencontact 764 488 764 488 0 FILL_1__1009_.vdd
rlabel metal1 744 242 776 258 0 FILL_1__1009_.gnd
rlabel nsubstratencontact 744 12 744 12 0 FILL_0__1012_.vdd
rlabel metal1 724 242 756 258 0 FILL_0__1012_.gnd
rlabel nsubstratencontact 744 488 744 488 0 FILL_0__1009_.vdd
rlabel metal1 724 242 756 258 0 FILL_0__1009_.gnd
rlabel nsubstratencontact 884 488 884 488 0 FILL_0__1087_.vdd
rlabel metal1 864 242 896 258 0 FILL_0__1087_.gnd
rlabel nsubstratencontact 876 12 876 12 0 FILL_0__1005_.vdd
rlabel metal1 864 242 896 258 0 FILL_0__1005_.gnd
rlabel metal1 764 242 876 258 0 _1012_.gnd
rlabel metal1 764 2 876 18 0 _1012_.vdd
rlabel metal2 853 133 867 147 0 _1012_.A
rlabel metal2 833 113 847 127 0 _1012_.B
rlabel metal2 813 133 827 147 0 _1012_.C
rlabel metal2 793 113 807 127 0 _1012_.Y
rlabel metal1 764 242 876 258 0 _1009_.gnd
rlabel metal1 764 482 876 498 0 _1009_.vdd
rlabel metal2 853 353 867 367 0 _1009_.A
rlabel metal2 833 373 847 387 0 _1009_.B
rlabel metal2 813 353 827 367 0 _1009_.C
rlabel metal2 793 373 807 387 0 _1009_.Y
rlabel nsubstratencontact 904 488 904 488 0 FILL_1__1087_.vdd
rlabel metal1 884 242 916 258 0 FILL_1__1087_.gnd
rlabel nsubstratencontact 996 12 996 12 0 FILL_1__1070_.vdd
rlabel metal1 984 242 1016 258 0 FILL_1__1070_.gnd
rlabel nsubstratencontact 896 12 896 12 0 FILL_1__1005_.vdd
rlabel metal1 884 242 916 258 0 FILL_1__1005_.gnd
rlabel nsubstratencontact 1016 488 1016 488 0 FILL_0__1073_.vdd
rlabel metal1 1004 242 1036 258 0 FILL_0__1073_.gnd
rlabel nsubstratencontact 976 12 976 12 0 FILL_0__1070_.vdd
rlabel metal1 964 242 996 258 0 FILL_0__1070_.gnd
rlabel metal1 904 242 1016 258 0 _1087_.gnd
rlabel metal1 904 482 1016 498 0 _1087_.vdd
rlabel metal2 993 353 1007 367 0 _1087_.A
rlabel metal2 973 313 987 327 0 _1087_.B
rlabel metal2 953 353 967 367 0 _1087_.C
rlabel metal2 933 333 947 347 0 _1087_.Y
rlabel metal1 1004 242 1116 258 0 _1070_.gnd
rlabel metal1 1004 2 1116 18 0 _1070_.vdd
rlabel metal2 1013 153 1027 167 0 _1070_.A
rlabel metal2 1033 133 1047 147 0 _1070_.B
rlabel metal2 1073 133 1087 147 0 _1070_.C
rlabel metal2 1053 153 1067 167 0 _1070_.Y
rlabel metal1 904 242 976 258 0 _1005_.gnd
rlabel metal1 904 2 976 18 0 _1005_.vdd
rlabel metal2 913 173 927 187 0 _1005_.A
rlabel metal2 933 133 947 147 0 _1005_.Y
rlabel nsubstratencontact 1036 488 1036 488 0 FILL_1__1073_.vdd
rlabel metal1 1024 242 1056 258 0 FILL_1__1073_.gnd
rlabel nsubstratencontact 1136 12 1136 12 0 FILL_1__1057_.vdd
rlabel metal1 1124 242 1156 258 0 FILL_1__1057_.gnd
rlabel nsubstratencontact 1116 12 1116 12 0 FILL_0__1057_.vdd
rlabel metal1 1104 242 1136 258 0 FILL_0__1057_.gnd
rlabel metal1 1044 242 1156 258 0 _1073_.gnd
rlabel metal1 1044 482 1156 498 0 _1073_.vdd
rlabel metal2 1053 353 1067 367 0 _1073_.A
rlabel metal2 1073 373 1087 387 0 _1073_.B
rlabel metal2 1093 353 1107 367 0 _1073_.C
rlabel metal2 1113 373 1127 387 0 _1073_.Y
rlabel nsubstratencontact 1184 488 1184 488 0 FILL_1__1007_.vdd
rlabel metal1 1164 242 1196 258 0 FILL_1__1007_.gnd
rlabel nsubstratencontact 1164 488 1164 488 0 FILL_0__1007_.vdd
rlabel metal1 1144 242 1176 258 0 FILL_0__1007_.gnd
rlabel nsubstratencontact 1256 12 1256 12 0 FILL_0__1002_.vdd
rlabel metal1 1244 242 1276 258 0 FILL_0__1002_.gnd
rlabel metal1 1144 242 1256 258 0 _1057_.gnd
rlabel metal1 1144 2 1256 18 0 _1057_.vdd
rlabel metal2 1153 133 1167 147 0 _1057_.A
rlabel metal2 1173 173 1187 187 0 _1057_.B
rlabel metal2 1193 133 1207 147 0 _1057_.C
rlabel metal2 1213 153 1227 167 0 _1057_.Y
rlabel metal1 1184 242 1296 258 0 _1007_.gnd
rlabel metal1 1184 482 1296 498 0 _1007_.vdd
rlabel metal2 1273 313 1287 327 0 _1007_.A
rlabel metal2 1253 333 1267 347 0 _1007_.B
rlabel metal2 1213 353 1227 367 0 _1007_.Y
rlabel nsubstratencontact 1324 488 1324 488 0 FILL_1__1071_.vdd
rlabel metal1 1304 242 1336 258 0 FILL_1__1071_.gnd
rlabel nsubstratencontact 1396 12 1396 12 0 FILL_1__1003_.vdd
rlabel metal1 1384 242 1416 258 0 FILL_1__1003_.gnd
rlabel nsubstratencontact 1276 12 1276 12 0 FILL_1__1002_.vdd
rlabel metal1 1264 242 1296 258 0 FILL_1__1002_.gnd
rlabel nsubstratencontact 1304 488 1304 488 0 FILL_0__1071_.vdd
rlabel metal1 1284 242 1316 258 0 FILL_0__1071_.gnd
rlabel nsubstratencontact 1376 12 1376 12 0 FILL_0__1003_.vdd
rlabel metal1 1364 242 1396 258 0 FILL_0__1003_.gnd
rlabel metal1 1324 242 1436 258 0 _1071_.gnd
rlabel metal1 1324 482 1436 498 0 _1071_.vdd
rlabel metal2 1413 353 1427 367 0 _1071_.A
rlabel metal2 1393 373 1407 387 0 _1071_.B
rlabel metal2 1373 353 1387 367 0 _1071_.C
rlabel metal2 1353 373 1367 387 0 _1071_.Y
rlabel metal1 1284 242 1376 258 0 _1002_.gnd
rlabel metal1 1284 2 1376 18 0 _1002_.vdd
rlabel metal2 1333 153 1347 167 0 _1002_.B
rlabel metal2 1293 153 1307 167 0 _1002_.A
rlabel metal2 1313 173 1327 187 0 _1002_.Y
rlabel nsubstratencontact 1484 488 1484 488 0 FILL_2__1063_.vdd
rlabel metal1 1464 242 1496 258 0 FILL_2__1063_.gnd
rlabel nsubstratencontact 1464 488 1464 488 0 FILL_1__1063_.vdd
rlabel metal1 1444 242 1476 258 0 FILL_1__1063_.gnd
rlabel nsubstratencontact 1524 12 1524 12 0 FILL_0__1883_.vdd
rlabel metal1 1504 242 1536 258 0 FILL_0__1883_.gnd
rlabel nsubstratencontact 1444 488 1444 488 0 FILL_0__1063_.vdd
rlabel metal1 1424 242 1456 258 0 FILL_0__1063_.gnd
rlabel metal1 1484 242 1556 258 0 _1063_.gnd
rlabel metal1 1484 482 1556 498 0 _1063_.vdd
rlabel metal2 1533 313 1547 327 0 _1063_.A
rlabel metal2 1513 353 1527 367 0 _1063_.Y
rlabel metal1 1404 242 1516 258 0 _1003_.gnd
rlabel metal1 1404 2 1516 18 0 _1003_.vdd
rlabel metal2 1413 153 1427 167 0 _1003_.A
rlabel metal2 1473 153 1487 167 0 _1003_.Y
rlabel metal2 1453 113 1467 127 0 _1003_.B
rlabel nsubstratencontact 1644 12 1644 12 0 FILL_1__1884_.vdd
rlabel metal1 1624 242 1656 258 0 FILL_1__1884_.gnd
rlabel nsubstratencontact 1544 12 1544 12 0 FILL_1__1883_.vdd
rlabel metal1 1524 242 1556 258 0 FILL_1__1883_.gnd
rlabel nsubstratencontact 1584 488 1584 488 0 FILL_1__1072_.vdd
rlabel metal1 1564 242 1596 258 0 FILL_1__1072_.gnd
rlabel nsubstratencontact 1624 12 1624 12 0 FILL_0__1884_.vdd
rlabel metal1 1604 242 1636 258 0 FILL_0__1884_.gnd
rlabel nsubstratencontact 1564 488 1564 488 0 FILL_0__1072_.vdd
rlabel metal1 1544 242 1576 258 0 FILL_0__1072_.gnd
rlabel metal1 1544 242 1616 258 0 _1883_.gnd
rlabel metal1 1544 2 1616 18 0 _1883_.vdd
rlabel metal2 1593 173 1607 187 0 _1883_.A
rlabel metal2 1573 133 1587 147 0 _1883_.Y
rlabel metal1 1584 242 1696 258 0 _1072_.gnd
rlabel metal1 1584 482 1696 498 0 _1072_.vdd
rlabel metal2 1673 333 1687 347 0 _1072_.A
rlabel metal2 1653 353 1667 367 0 _1072_.B
rlabel metal2 1613 353 1627 367 0 _1072_.C
rlabel metal2 1633 333 1647 347 0 _1072_.Y
rlabel nsubstratencontact 1784 12 1784 12 0 FILL_1__1887_.vdd
rlabel metal1 1764 242 1796 258 0 FILL_1__1887_.gnd
rlabel nsubstratencontact 1724 488 1724 488 0 FILL_1__1876_.vdd
rlabel metal1 1704 242 1736 258 0 FILL_1__1876_.gnd
rlabel nsubstratencontact 1764 12 1764 12 0 FILL_0__1887_.vdd
rlabel metal1 1744 242 1776 258 0 FILL_0__1887_.gnd
rlabel nsubstratencontact 1704 488 1704 488 0 FILL_0__1876_.vdd
rlabel metal1 1684 242 1716 258 0 FILL_0__1876_.gnd
rlabel metal1 1644 242 1756 258 0 _1884_.gnd
rlabel metal1 1644 2 1756 18 0 _1884_.vdd
rlabel metal2 1733 153 1747 167 0 _1884_.A
rlabel metal2 1713 133 1727 147 0 _1884_.B
rlabel metal2 1673 133 1687 147 0 _1884_.C
rlabel metal2 1693 153 1707 167 0 _1884_.Y
rlabel metal1 1724 242 1836 258 0 _1876_.gnd
rlabel metal1 1724 482 1836 498 0 _1876_.vdd
rlabel metal2 1813 333 1827 347 0 _1876_.A
rlabel metal2 1753 333 1767 347 0 _1876_.Y
rlabel metal2 1773 373 1787 387 0 _1876_.B
rlabel nsubstratencontact 1896 12 1896 12 0 FILL_1__1886_.vdd
rlabel metal1 1884 242 1916 258 0 FILL_1__1886_.gnd
rlabel nsubstratencontact 1856 488 1856 488 0 FILL_1__1875_.vdd
rlabel metal1 1844 242 1876 258 0 FILL_1__1875_.gnd
rlabel nsubstratencontact 1876 12 1876 12 0 FILL_0__1886_.vdd
rlabel metal1 1864 242 1896 258 0 FILL_0__1886_.gnd
rlabel nsubstratencontact 1836 488 1836 488 0 FILL_0__1875_.vdd
rlabel metal1 1824 242 1856 258 0 FILL_0__1875_.gnd
rlabel metal1 1784 242 1876 258 0 _1887_.gnd
rlabel metal1 1784 2 1876 18 0 _1887_.vdd
rlabel metal2 1853 113 1867 127 0 _1887_.A
rlabel metal2 1813 113 1827 127 0 _1887_.B
rlabel metal2 1833 133 1847 147 0 _1887_.Y
rlabel metal1 1864 242 1956 258 0 _1875_.gnd
rlabel metal1 1864 482 1956 498 0 _1875_.vdd
rlabel metal2 1913 333 1927 347 0 _1875_.B
rlabel metal2 1873 333 1887 347 0 _1875_.A
rlabel metal2 1893 313 1907 327 0 _1875_.Y
rlabel nsubstratencontact 1996 488 1996 488 0 FILL_2__1846_.vdd
rlabel metal1 1984 242 2016 258 0 FILL_2__1846_.gnd
rlabel nsubstratencontact 1976 488 1976 488 0 FILL_1__1846_.vdd
rlabel metal1 1964 242 1996 258 0 FILL_1__1846_.gnd
rlabel nsubstratencontact 2024 12 2024 12 0 FILL_0__1885_.vdd
rlabel metal1 2004 242 2036 258 0 FILL_0__1885_.gnd
rlabel nsubstratencontact 1956 488 1956 488 0 FILL_0__1846_.vdd
rlabel metal1 1944 242 1976 258 0 FILL_0__1846_.gnd
rlabel metal1 1904 242 2016 258 0 _1886_.gnd
rlabel metal1 1904 2 2016 18 0 _1886_.vdd
rlabel metal2 1913 133 1927 147 0 _1886_.A
rlabel metal2 1933 113 1947 127 0 _1886_.B
rlabel metal2 1953 133 1967 147 0 _1886_.C
rlabel metal2 1973 113 1987 127 0 _1886_.Y
rlabel metal1 2004 242 2076 258 0 _1846_.gnd
rlabel metal1 2004 482 2076 498 0 _1846_.vdd
rlabel metal2 2013 313 2027 327 0 _1846_.A
rlabel metal2 2033 353 2047 367 0 _1846_.Y
rlabel nsubstratencontact 2064 12 2064 12 0 FILL_2__1885_.vdd
rlabel metal1 2044 242 2076 258 0 FILL_2__1885_.gnd
rlabel nsubstratencontact 2044 12 2044 12 0 FILL_1__1885_.vdd
rlabel metal1 2024 242 2056 258 0 FILL_1__1885_.gnd
rlabel nsubstratencontact 2104 488 2104 488 0 FILL_1__1847_.vdd
rlabel metal1 2084 242 2116 258 0 FILL_1__1847_.gnd
rlabel nsubstratencontact 2084 488 2084 488 0 FILL_0__1847_.vdd
rlabel metal1 2064 242 2096 258 0 FILL_0__1847_.gnd
rlabel metal1 2064 242 2176 258 0 _1885_.gnd
rlabel metal1 2064 2 2176 18 0 _1885_.vdd
rlabel metal2 2153 133 2167 147 0 _1885_.A
rlabel metal2 2133 113 2147 127 0 _1885_.B
rlabel metal2 2113 133 2127 147 0 _1885_.C
rlabel metal2 2093 113 2107 127 0 _1885_.Y
rlabel metal1 2104 242 2216 258 0 _1847_.gnd
rlabel metal1 2104 482 2216 498 0 _1847_.vdd
rlabel metal2 2193 333 2207 347 0 _1847_.A
rlabel metal2 2173 353 2187 367 0 _1847_.B
rlabel metal2 2133 353 2147 367 0 _1847_.C
rlabel metal2 2153 333 2167 347 0 _1847_.Y
rlabel nsubstratencontact 2196 12 2196 12 0 FILL_1__1893_.vdd
rlabel metal1 2184 242 2216 258 0 FILL_1__1893_.gnd
rlabel nsubstratencontact 2244 488 2244 488 0 FILL_1__1874_.vdd
rlabel metal1 2224 242 2256 258 0 FILL_1__1874_.gnd
rlabel nsubstratencontact 2176 12 2176 12 0 FILL_0__1893_.vdd
rlabel metal1 2164 242 2196 258 0 FILL_0__1893_.gnd
rlabel nsubstratencontact 2224 488 2224 488 0 FILL_0__1874_.vdd
rlabel metal1 2204 242 2236 258 0 FILL_0__1874_.gnd
rlabel metal1 2204 242 2296 258 0 _1893_.gnd
rlabel metal1 2204 2 2296 18 0 _1893_.vdd
rlabel metal2 2213 153 2227 167 0 _1893_.A
rlabel metal2 2253 153 2267 167 0 _1893_.Y
rlabel metal1 2244 242 2356 258 0 _1874_.gnd
rlabel metal1 2244 482 2356 498 0 _1874_.vdd
rlabel metal2 2333 353 2347 367 0 _1874_.A
rlabel metal2 2313 313 2327 327 0 _1874_.B
rlabel metal2 2293 353 2307 367 0 _1874_.C
rlabel metal2 2273 333 2287 347 0 _1874_.Y
rlabel nsubstratencontact 2324 12 2324 12 0 FILL_1__1857_.vdd
rlabel metal1 2304 242 2336 258 0 FILL_1__1857_.gnd
rlabel nsubstratencontact 2384 488 2384 488 0 FILL_1__1834_.vdd
rlabel metal1 2364 242 2396 258 0 FILL_1__1834_.gnd
rlabel nsubstratencontact 2304 12 2304 12 0 FILL_0__1857_.vdd
rlabel metal1 2284 242 2316 258 0 FILL_0__1857_.gnd
rlabel nsubstratencontact 2364 488 2364 488 0 FILL_0__1834_.vdd
rlabel metal1 2344 242 2376 258 0 FILL_0__1834_.gnd
rlabel metal1 2324 242 2416 258 0 _1857_.gnd
rlabel metal1 2324 2 2416 18 0 _1857_.vdd
rlabel metal2 2393 113 2407 127 0 _1857_.A
rlabel metal2 2353 113 2367 127 0 _1857_.B
rlabel metal2 2373 133 2387 147 0 _1857_.Y
rlabel metal1 2384 242 2456 258 0 _1834_.gnd
rlabel metal1 2384 482 2456 498 0 _1834_.vdd
rlabel metal2 2433 313 2447 327 0 _1834_.A
rlabel metal2 2413 353 2427 367 0 _1834_.Y
rlabel nsubstratencontact 2436 12 2436 12 0 FILL_1__1849_.vdd
rlabel metal1 2424 242 2456 258 0 FILL_1__1849_.gnd
rlabel nsubstratencontact 2484 488 2484 488 0 FILL_1__1848_.vdd
rlabel metal1 2464 242 2496 258 0 FILL_1__1848_.gnd
rlabel nsubstratencontact 2416 12 2416 12 0 FILL_0__1849_.vdd
rlabel metal1 2404 242 2436 258 0 FILL_0__1849_.gnd
rlabel nsubstratencontact 2464 488 2464 488 0 FILL_0__1848_.vdd
rlabel metal1 2444 242 2476 258 0 FILL_0__1848_.gnd
rlabel metal1 2444 242 2556 258 0 _1849_.gnd
rlabel metal1 2444 2 2556 18 0 _1849_.vdd
rlabel metal2 2453 153 2467 167 0 _1849_.A
rlabel metal2 2513 153 2527 167 0 _1849_.Y
rlabel metal2 2493 113 2507 127 0 _1849_.B
rlabel metal1 2484 242 2596 258 0 _1848_.gnd
rlabel metal1 2484 482 2596 498 0 _1848_.vdd
rlabel metal2 2573 353 2587 367 0 _1848_.A
rlabel metal2 2553 373 2567 387 0 _1848_.B
rlabel metal2 2533 353 2547 367 0 _1848_.C
rlabel metal2 2513 373 2527 387 0 _1848_.Y
rlabel nsubstratencontact 2584 12 2584 12 0 FILL_1__1873_.vdd
rlabel metal1 2564 242 2596 258 0 FILL_1__1873_.gnd
rlabel nsubstratencontact 2616 488 2616 488 0 FILL_1__1870_.vdd
rlabel metal1 2604 242 2636 258 0 FILL_1__1870_.gnd
rlabel nsubstratencontact 2564 12 2564 12 0 FILL_0__1873_.vdd
rlabel metal1 2544 242 2576 258 0 FILL_0__1873_.gnd
rlabel nsubstratencontact 2596 488 2596 488 0 FILL_0__1870_.vdd
rlabel metal1 2584 242 2616 258 0 FILL_0__1870_.gnd
rlabel metal1 2584 242 2696 258 0 _1873_.gnd
rlabel metal1 2584 2 2696 18 0 _1873_.vdd
rlabel metal2 2673 133 2687 147 0 _1873_.A
rlabel metal2 2653 173 2667 187 0 _1873_.B
rlabel metal2 2633 133 2647 147 0 _1873_.C
rlabel metal2 2613 153 2627 167 0 _1873_.Y
rlabel metal1 2624 242 2736 258 0 _1870_.gnd
rlabel metal1 2624 482 2736 498 0 _1870_.vdd
rlabel metal2 2633 333 2647 347 0 _1870_.A
rlabel metal2 2653 353 2667 367 0 _1870_.B
rlabel metal2 2693 353 2707 367 0 _1870_.C
rlabel metal2 2673 333 2687 347 0 _1870_.Y
rlabel nsubstratencontact 2724 12 2724 12 0 FILL_1__1869_.vdd
rlabel metal1 2704 242 2736 258 0 FILL_1__1869_.gnd
rlabel nsubstratencontact 2764 488 2764 488 0 FILL_1__1829_.vdd
rlabel metal1 2744 242 2776 258 0 FILL_1__1829_.gnd
rlabel nsubstratencontact 2704 12 2704 12 0 FILL_0__1869_.vdd
rlabel metal1 2684 242 2716 258 0 FILL_0__1869_.gnd
rlabel nsubstratencontact 2744 488 2744 488 0 FILL_0__1829_.vdd
rlabel metal1 2724 242 2756 258 0 FILL_0__1829_.gnd
rlabel metal1 2724 242 2836 258 0 _1869_.gnd
rlabel metal1 2724 2 2836 18 0 _1869_.vdd
rlabel metal2 2813 153 2827 167 0 _1869_.A
rlabel metal2 2753 153 2767 167 0 _1869_.Y
rlabel metal2 2773 113 2787 127 0 _1869_.B
rlabel metal1 2764 242 2836 258 0 _1829_.gnd
rlabel metal1 2764 482 2836 498 0 _1829_.vdd
rlabel metal2 2813 313 2827 327 0 _1829_.A
rlabel metal2 2793 353 2807 367 0 _1829_.Y
rlabel nsubstratencontact 2876 12 2876 12 0 FILL_2__1872_.vdd
rlabel metal1 2864 242 2896 258 0 FILL_2__1872_.gnd
rlabel nsubstratencontact 2856 12 2856 12 0 FILL_1__1872_.vdd
rlabel metal1 2844 242 2876 258 0 FILL_1__1872_.gnd
rlabel nsubstratencontact 2864 488 2864 488 0 FILL_1__1861_.vdd
rlabel metal1 2844 242 2876 258 0 FILL_1__1861_.gnd
rlabel nsubstratencontact 2836 12 2836 12 0 FILL_0__1872_.vdd
rlabel metal1 2824 242 2856 258 0 FILL_0__1872_.gnd
rlabel nsubstratencontact 2844 488 2844 488 0 FILL_0__1861_.vdd
rlabel metal1 2824 242 2856 258 0 FILL_0__1861_.gnd
rlabel metal1 2884 242 2976 258 0 _1872_.gnd
rlabel metal1 2884 2 2976 18 0 _1872_.vdd
rlabel metal2 2893 113 2907 127 0 _1872_.A
rlabel metal2 2933 113 2947 127 0 _1872_.B
rlabel metal2 2913 133 2927 147 0 _1872_.Y
rlabel metal1 2864 242 2956 258 0 _1861_.gnd
rlabel metal1 2864 482 2956 498 0 _1861_.vdd
rlabel metal2 2893 333 2907 347 0 _1861_.B
rlabel metal2 2933 333 2947 347 0 _1861_.A
rlabel metal2 2913 313 2927 327 0 _1861_.Y
rlabel nsubstratencontact 2976 488 2976 488 0 FILL_1__1865_.vdd
rlabel metal1 2964 242 2996 258 0 FILL_1__1865_.gnd
rlabel nsubstratencontact 3004 12 3004 12 0 FILL_1__1862_.vdd
rlabel metal1 2984 242 3016 258 0 FILL_1__1862_.gnd
rlabel nsubstratencontact 2956 488 2956 488 0 FILL_0__1865_.vdd
rlabel metal1 2944 242 2976 258 0 FILL_0__1865_.gnd
rlabel nsubstratencontact 2984 12 2984 12 0 FILL_0__1862_.vdd
rlabel metal1 2964 242 2996 258 0 FILL_0__1862_.gnd
rlabel metal1 2984 242 3056 258 0 _1865_.gnd
rlabel metal1 2984 482 3056 498 0 _1865_.vdd
rlabel metal2 2993 313 3007 327 0 _1865_.A
rlabel metal2 3013 353 3027 367 0 _1865_.Y
rlabel metal1 3004 242 3096 258 0 _1862_.gnd
rlabel metal1 3004 2 3096 18 0 _1862_.vdd
rlabel metal2 3073 113 3087 127 0 _1862_.A
rlabel metal2 3033 113 3047 127 0 _1862_.B
rlabel metal2 3053 133 3067 147 0 _1862_.Y
rlabel nsubstratencontact 3124 12 3124 12 0 FILL_1__1864_.vdd
rlabel metal1 3104 242 3136 258 0 FILL_1__1864_.gnd
rlabel nsubstratencontact 3084 488 3084 488 0 FILL_1__1835_.vdd
rlabel metal1 3064 242 3096 258 0 FILL_1__1835_.gnd
rlabel nsubstratencontact 3104 12 3104 12 0 FILL_0__1864_.vdd
rlabel metal1 3084 242 3116 258 0 FILL_0__1864_.gnd
rlabel nsubstratencontact 3064 488 3064 488 0 FILL_0__1835_.vdd
rlabel metal1 3044 242 3076 258 0 FILL_0__1835_.gnd
rlabel metal1 3124 242 3236 258 0 _1864_.gnd
rlabel metal1 3124 2 3236 18 0 _1864_.vdd
rlabel metal2 3213 133 3227 147 0 _1864_.A
rlabel metal2 3193 113 3207 127 0 _1864_.B
rlabel metal2 3173 133 3187 147 0 _1864_.C
rlabel metal2 3153 113 3167 127 0 _1864_.Y
rlabel metal1 3084 242 3196 258 0 _1835_.gnd
rlabel metal1 3084 482 3196 498 0 _1835_.vdd
rlabel metal2 3173 353 3187 367 0 _1835_.A
rlabel metal2 3153 313 3167 327 0 _1835_.B
rlabel metal2 3133 353 3147 367 0 _1835_.C
rlabel metal2 3113 333 3127 347 0 _1835_.Y
rlabel nsubstratencontact 3236 488 3236 488 0 FILL_2__1866_.vdd
rlabel metal1 3224 242 3256 258 0 FILL_2__1866_.gnd
rlabel nsubstratencontact 3216 488 3216 488 0 FILL_1__1866_.vdd
rlabel metal1 3204 242 3236 258 0 FILL_1__1866_.gnd
rlabel nsubstratencontact 3264 12 3264 12 0 FILL_1__1860_.vdd
rlabel metal1 3244 242 3276 258 0 FILL_1__1860_.gnd
rlabel nsubstratencontact 3196 488 3196 488 0 FILL_0__1866_.vdd
rlabel metal1 3184 242 3216 258 0 FILL_0__1866_.gnd
rlabel nsubstratencontact 3244 12 3244 12 0 FILL_0__1860_.vdd
rlabel metal1 3224 242 3256 258 0 FILL_0__1860_.gnd
rlabel metal1 3244 242 3356 258 0 _1866_.gnd
rlabel metal1 3244 482 3356 498 0 _1866_.vdd
rlabel metal2 3253 353 3267 367 0 _1866_.A
rlabel metal2 3273 313 3287 327 0 _1866_.B
rlabel metal2 3293 353 3307 367 0 _1866_.C
rlabel metal2 3313 333 3327 347 0 _1866_.Y
rlabel metal1 3264 242 3336 258 0 _1860_.gnd
rlabel metal1 3264 2 3336 18 0 _1860_.vdd
rlabel metal2 3313 173 3327 187 0 _1860_.A
rlabel metal2 3293 133 3307 147 0 _1860_.Y
rlabel nsubstratencontact 3356 12 3356 12 0 FILL_1__1868_.vdd
rlabel metal1 3344 242 3376 258 0 FILL_1__1868_.gnd
rlabel nsubstratencontact 3384 488 3384 488 0 FILL_1__1739_.vdd
rlabel metal1 3364 242 3396 258 0 FILL_1__1739_.gnd
rlabel nsubstratencontact 3336 12 3336 12 0 FILL_0__1868_.vdd
rlabel metal1 3324 242 3356 258 0 FILL_0__1868_.gnd
rlabel nsubstratencontact 3364 488 3364 488 0 FILL_0__1739_.vdd
rlabel metal1 3344 242 3376 258 0 FILL_0__1739_.gnd
rlabel metal1 3364 242 3476 258 0 _1868_.gnd
rlabel metal1 3364 2 3476 18 0 _1868_.vdd
rlabel metal2 3373 153 3387 167 0 _1868_.A
rlabel metal2 3393 133 3407 147 0 _1868_.B
rlabel metal2 3433 133 3447 147 0 _1868_.C
rlabel metal2 3413 153 3427 167 0 _1868_.Y
rlabel metal1 3384 242 3456 258 0 _1739_.gnd
rlabel metal1 3384 482 3456 498 0 _1739_.vdd
rlabel metal2 3433 313 3447 327 0 _1739_.A
rlabel metal2 3413 353 3427 367 0 _1739_.Y
rlabel nsubstratencontact 3496 488 3496 488 0 FILL_2__1859_.vdd
rlabel metal1 3484 242 3516 258 0 FILL_2__1859_.gnd
rlabel nsubstratencontact 3504 12 3504 12 0 FILL_1__1867_.vdd
rlabel metal1 3484 242 3516 258 0 FILL_1__1867_.gnd
rlabel nsubstratencontact 3476 488 3476 488 0 FILL_1__1859_.vdd
rlabel metal1 3464 242 3496 258 0 FILL_1__1859_.gnd
rlabel nsubstratencontact 3484 12 3484 12 0 FILL_0__1867_.vdd
rlabel metal1 3464 242 3496 258 0 FILL_0__1867_.gnd
rlabel nsubstratencontact 3456 488 3456 488 0 FILL_0__1859_.vdd
rlabel metal1 3444 242 3476 258 0 FILL_0__1859_.gnd
rlabel metal1 3504 242 3576 258 0 _1867_.gnd
rlabel metal1 3504 2 3576 18 0 _1867_.vdd
rlabel metal2 3553 173 3567 187 0 _1867_.A
rlabel metal2 3533 133 3547 147 0 _1867_.Y
rlabel metal1 3504 242 3616 258 0 _1859_.gnd
rlabel metal1 3504 482 3616 498 0 _1859_.vdd
rlabel metal2 3513 333 3527 347 0 _1859_.A
rlabel metal2 3533 353 3547 367 0 _1859_.B
rlabel metal2 3573 353 3587 367 0 _1859_.C
rlabel metal2 3553 333 3567 347 0 _1859_.Y
rlabel nsubstratencontact 3636 488 3636 488 0 FILL_1__1778_.vdd
rlabel metal1 3624 242 3656 258 0 FILL_1__1778_.gnd
rlabel nsubstratencontact 3604 12 3604 12 0 FILL_1__1758_.vdd
rlabel metal1 3584 242 3616 258 0 FILL_1__1758_.gnd
rlabel nsubstratencontact 3616 488 3616 488 0 FILL_0__1778_.vdd
rlabel metal1 3604 242 3636 258 0 FILL_0__1778_.gnd
rlabel nsubstratencontact 3584 12 3584 12 0 FILL_0__1758_.vdd
rlabel metal1 3564 242 3596 258 0 FILL_0__1758_.gnd
rlabel metal1 3644 242 3756 258 0 _1778_.gnd
rlabel metal1 3644 482 3756 498 0 _1778_.vdd
rlabel metal2 3653 353 3667 367 0 _1778_.A
rlabel metal2 3673 313 3687 327 0 _1778_.B
rlabel metal2 3693 353 3707 367 0 _1778_.C
rlabel metal2 3713 333 3727 347 0 _1778_.Y
rlabel metal1 3604 242 3696 258 0 _1758_.gnd
rlabel metal1 3604 2 3696 18 0 _1758_.vdd
rlabel metal2 3673 113 3687 127 0 _1758_.A
rlabel metal2 3633 113 3647 127 0 _1758_.B
rlabel metal2 3653 133 3667 147 0 _1758_.Y
rlabel nsubstratencontact 3724 12 3724 12 0 FILL_1__1895_.vdd
rlabel metal1 3704 242 3736 258 0 FILL_1__1895_.gnd
rlabel nsubstratencontact 3784 488 3784 488 0 FILL_1__1779_.vdd
rlabel metal1 3764 242 3796 258 0 FILL_1__1779_.gnd
rlabel nsubstratencontact 3704 12 3704 12 0 FILL_0__1895_.vdd
rlabel metal1 3684 242 3716 258 0 FILL_0__1895_.gnd
rlabel nsubstratencontact 3764 488 3764 488 0 FILL_0__1779_.vdd
rlabel metal1 3744 242 3776 258 0 FILL_0__1779_.gnd
rlabel metal1 3724 242 3816 258 0 _1895_.gnd
rlabel metal1 3724 2 3816 18 0 _1895_.vdd
rlabel metal2 3793 153 3807 167 0 _1895_.A
rlabel metal2 3753 153 3767 167 0 _1895_.Y
rlabel metal1 3784 242 3896 258 0 _1779_.gnd
rlabel metal1 3784 482 3896 498 0 _1779_.vdd
rlabel metal2 3873 353 3887 367 0 _1779_.A
rlabel metal2 3853 373 3867 387 0 _1779_.B
rlabel metal2 3833 353 3847 367 0 _1779_.C
rlabel metal2 3813 373 3827 387 0 _1779_.Y
rlabel nsubstratencontact 3836 12 3836 12 0 FILL_1__1897_.vdd
rlabel metal1 3824 242 3856 258 0 FILL_1__1897_.gnd
rlabel nsubstratencontact 3916 488 3916 488 0 FILL_1__1775_.vdd
rlabel metal1 3904 242 3936 258 0 FILL_1__1775_.gnd
rlabel nsubstratencontact 3816 12 3816 12 0 FILL_0__1897_.vdd
rlabel metal1 3804 242 3836 258 0 FILL_0__1897_.gnd
rlabel nsubstratencontact 3896 488 3896 488 0 FILL_0__1775_.vdd
rlabel metal1 3884 242 3916 258 0 FILL_0__1775_.gnd
rlabel metal1 3844 242 3936 258 0 _1897_.gnd
rlabel metal1 3844 2 3936 18 0 _1897_.vdd
rlabel metal2 3853 153 3867 167 0 _1897_.A
rlabel metal2 3893 153 3907 167 0 _1897_.Y
rlabel nsubstratencontact 4044 488 4044 488 0 FILL_1__1774_.vdd
rlabel metal1 4024 242 4056 258 0 FILL_1__1774_.gnd
rlabel nsubstratencontact 3964 12 3964 12 0 FILL_1__1754_.vdd
rlabel metal1 3944 242 3976 258 0 FILL_1__1754_.gnd
rlabel nsubstratencontact 4024 488 4024 488 0 FILL_0__1774_.vdd
rlabel metal1 4004 242 4036 258 0 FILL_0__1774_.gnd
rlabel nsubstratencontact 3944 12 3944 12 0 FILL_0__1754_.vdd
rlabel metal1 3924 242 3956 258 0 FILL_0__1754_.gnd
rlabel metal1 3924 242 4016 258 0 _1775_.gnd
rlabel metal1 3924 482 4016 498 0 _1775_.vdd
rlabel metal2 3933 373 3947 387 0 _1775_.A
rlabel metal2 3973 373 3987 387 0 _1775_.B
rlabel metal2 3953 353 3967 367 0 _1775_.Y
rlabel metal1 3964 242 4056 258 0 _1754_.gnd
rlabel metal1 3964 2 4056 18 0 _1754_.vdd
rlabel metal2 4033 113 4047 127 0 _1754_.A
rlabel metal2 3993 113 4007 127 0 _1754_.B
rlabel metal2 4013 133 4027 147 0 _1754_.Y
rlabel nsubstratencontact 4064 488 4064 488 0 FILL_2__1774_.vdd
rlabel metal1 4044 242 4076 258 0 FILL_2__1774_.gnd
rlabel nsubstratencontact 4096 12 4096 12 0 FILL_2__1761_.vdd
rlabel metal1 4084 242 4116 258 0 FILL_2__1761_.gnd
rlabel nsubstratencontact 4076 12 4076 12 0 FILL_1__1761_.vdd
rlabel metal1 4064 242 4096 258 0 FILL_1__1761_.gnd
rlabel nsubstratencontact 4184 488 4184 488 0 FILL_0__1795_.vdd
rlabel metal1 4164 242 4196 258 0 FILL_0__1795_.gnd
rlabel nsubstratencontact 4056 12 4056 12 0 FILL_0__1761_.vdd
rlabel metal1 4044 242 4076 258 0 FILL_0__1761_.gnd
rlabel metal1 4064 242 4176 258 0 _1774_.gnd
rlabel metal1 4064 482 4176 498 0 _1774_.vdd
rlabel metal2 4153 353 4167 367 0 _1774_.A
rlabel metal2 4133 373 4147 387 0 _1774_.B
rlabel metal2 4113 353 4127 367 0 _1774_.C
rlabel metal2 4093 373 4107 387 0 _1774_.Y
rlabel metal1 4104 242 4216 258 0 _1761_.gnd
rlabel metal1 4104 2 4216 18 0 _1761_.vdd
rlabel metal2 4113 153 4127 167 0 _1761_.A
rlabel metal2 4173 153 4187 167 0 _1761_.Y
rlabel metal2 4153 113 4167 127 0 _1761_.B
rlabel nsubstratencontact 4264 12 4264 12 0 FILL_2__1794_.vdd
rlabel metal1 4244 242 4276 258 0 FILL_2__1794_.gnd
rlabel nsubstratencontact 4204 488 4204 488 0 FILL_1__1795_.vdd
rlabel metal1 4184 242 4216 258 0 FILL_1__1795_.gnd
rlabel nsubstratencontact 4244 12 4244 12 0 FILL_1__1794_.vdd
rlabel metal1 4224 242 4256 258 0 FILL_1__1794_.gnd
rlabel nsubstratencontact 4224 12 4224 12 0 FILL_0__1794_.vdd
rlabel metal1 4204 242 4236 258 0 FILL_0__1794_.gnd
rlabel metal1 4204 242 4316 258 0 _1795_.gnd
rlabel metal1 4204 482 4316 498 0 _1795_.vdd
rlabel metal2 4293 333 4307 347 0 _1795_.A
rlabel metal2 4273 353 4287 367 0 _1795_.B
rlabel metal2 4233 353 4247 367 0 _1795_.C
rlabel metal2 4253 333 4267 347 0 _1795_.Y
rlabel metal1 4264 242 4356 258 0 _1794_.gnd
rlabel metal1 4264 2 4356 18 0 _1794_.vdd
rlabel metal2 4293 153 4307 167 0 _1794_.B
rlabel metal2 4333 153 4347 167 0 _1794_.A
rlabel metal2 4313 173 4327 187 0 _1794_.Y
rlabel nsubstratencontact 4344 488 4344 488 0 FILL_1__1772_.vdd
rlabel metal1 4324 242 4356 258 0 FILL_1__1772_.gnd
rlabel nsubstratencontact 4376 12 4376 12 0 FILL_1__1738_.vdd
rlabel metal1 4364 242 4396 258 0 FILL_1__1738_.gnd
rlabel nsubstratencontact 4424 488 4424 488 0 FILL_0__1780_.vdd
rlabel metal1 4404 242 4436 258 0 FILL_0__1780_.gnd
rlabel nsubstratencontact 4324 488 4324 488 0 FILL_0__1772_.vdd
rlabel metal1 4304 242 4336 258 0 FILL_0__1772_.gnd
rlabel nsubstratencontact 4356 12 4356 12 0 FILL_0__1738_.vdd
rlabel metal1 4344 242 4376 258 0 FILL_0__1738_.gnd
rlabel metal1 4344 242 4416 258 0 _1772_.gnd
rlabel metal1 4344 482 4416 498 0 _1772_.vdd
rlabel metal2 4393 313 4407 327 0 _1772_.A
rlabel metal2 4373 353 4387 367 0 _1772_.Y
rlabel metal1 4384 242 4476 258 0 _1738_.gnd
rlabel metal1 4384 2 4476 18 0 _1738_.vdd
rlabel metal2 4393 113 4407 127 0 _1738_.A
rlabel metal2 4433 113 4447 127 0 _1738_.B
rlabel metal2 4413 133 4427 147 0 _1738_.Y
rlabel nsubstratencontact 4444 488 4444 488 0 FILL_1__1780_.vdd
rlabel metal1 4424 242 4456 258 0 FILL_1__1780_.gnd
rlabel nsubstratencontact 4504 12 4504 12 0 FILL_1__1757_.vdd
rlabel metal1 4484 242 4516 258 0 FILL_1__1757_.gnd
rlabel nsubstratencontact 4544 488 4544 488 0 FILL_0__1773_.vdd
rlabel metal1 4524 242 4556 258 0 FILL_0__1773_.gnd
rlabel nsubstratencontact 4484 12 4484 12 0 FILL_0__1757_.vdd
rlabel metal1 4464 242 4496 258 0 FILL_0__1757_.gnd
rlabel metal1 4444 242 4536 258 0 _1780_.gnd
rlabel metal1 4444 482 4536 498 0 _1780_.vdd
rlabel metal2 4513 373 4527 387 0 _1780_.A
rlabel metal2 4473 373 4487 387 0 _1780_.B
rlabel metal2 4493 353 4507 367 0 _1780_.Y
rlabel metal1 4504 242 4616 258 0 _1757_.gnd
rlabel metal1 4504 2 4616 18 0 _1757_.vdd
rlabel metal2 4593 133 4607 147 0 _1757_.A
rlabel metal2 4573 113 4587 127 0 _1757_.B
rlabel metal2 4553 133 4567 147 0 _1757_.C
rlabel metal2 4533 113 4547 127 0 _1757_.Y
rlabel nsubstratencontact 4564 488 4564 488 0 FILL_1__1773_.vdd
rlabel metal1 4544 242 4576 258 0 FILL_1__1773_.gnd
rlabel nsubstratencontact 4664 12 4664 12 0 FILL_2__1741_.vdd
rlabel metal1 4644 242 4676 258 0 FILL_2__1741_.gnd
rlabel nsubstratencontact 4704 488 4704 488 0 FILL_1__1760_.vdd
rlabel metal1 4684 242 4716 258 0 FILL_1__1760_.gnd
rlabel nsubstratencontact 4644 12 4644 12 0 FILL_1__1741_.vdd
rlabel metal1 4624 242 4656 258 0 FILL_1__1741_.gnd
rlabel nsubstratencontact 4684 488 4684 488 0 FILL_0__1760_.vdd
rlabel metal1 4664 242 4696 258 0 FILL_0__1760_.gnd
rlabel nsubstratencontact 4624 12 4624 12 0 FILL_0__1741_.vdd
rlabel metal1 4604 242 4636 258 0 FILL_0__1741_.gnd
rlabel metal1 4564 242 4676 258 0 _1773_.gnd
rlabel metal1 4564 482 4676 498 0 _1773_.vdd
rlabel metal2 4653 333 4667 347 0 _1773_.A
rlabel metal2 4633 353 4647 367 0 _1773_.B
rlabel metal2 4593 353 4607 367 0 _1773_.C
rlabel metal2 4613 333 4627 347 0 _1773_.Y
rlabel metal1 4664 242 4776 258 0 _1741_.gnd
rlabel metal1 4664 2 4776 18 0 _1741_.vdd
rlabel metal2 4753 153 4767 167 0 _1741_.A
rlabel metal2 4733 133 4747 147 0 _1741_.B
rlabel metal2 4693 133 4707 147 0 _1741_.C
rlabel metal2 4713 153 4727 167 0 _1741_.Y
rlabel nsubstratencontact 4804 488 4804 488 0 FILL_1__1756_.vdd
rlabel metal1 4784 242 4816 258 0 FILL_1__1756_.gnd
rlabel nsubstratencontact 4796 12 4796 12 0 FILL_1__1737_.vdd
rlabel metal1 4784 242 4816 258 0 FILL_1__1737_.gnd
rlabel nsubstratencontact 4784 488 4784 488 0 FILL_0__1756_.vdd
rlabel metal1 4764 242 4796 258 0 FILL_0__1756_.gnd
rlabel nsubstratencontact 4776 12 4776 12 0 FILL_0__1737_.vdd
rlabel metal1 4764 242 4796 258 0 FILL_0__1737_.gnd
rlabel metal1 4704 242 4776 258 0 _1760_.gnd
rlabel metal1 4704 482 4776 498 0 _1760_.vdd
rlabel metal2 4753 313 4767 327 0 _1760_.A
rlabel metal2 4733 353 4747 367 0 _1760_.Y
rlabel metal1 4804 242 4916 258 0 _1756_.gnd
rlabel metal1 4804 482 4916 498 0 _1756_.vdd
rlabel metal2 4893 333 4907 347 0 _1756_.A
rlabel metal2 4873 353 4887 367 0 _1756_.B
rlabel metal2 4833 353 4847 367 0 _1756_.C
rlabel metal2 4853 333 4867 347 0 _1756_.Y
rlabel metal1 4804 242 4896 258 0 _1737_.gnd
rlabel metal1 4804 2 4896 18 0 _1737_.vdd
rlabel metal2 4813 113 4827 127 0 _1737_.A
rlabel metal2 4853 113 4867 127 0 _1737_.B
rlabel metal2 4833 133 4847 147 0 _1737_.Y
rlabel nsubstratencontact 4936 488 4936 488 0 FILL_1__1753_.vdd
rlabel metal1 4924 242 4956 258 0 FILL_1__1753_.gnd
rlabel nsubstratencontact 4924 12 4924 12 0 FILL_1__1736_.vdd
rlabel metal1 4904 242 4936 258 0 FILL_1__1736_.gnd
rlabel nsubstratencontact 4916 488 4916 488 0 FILL_0__1753_.vdd
rlabel metal1 4904 242 4936 258 0 FILL_0__1753_.gnd
rlabel nsubstratencontact 4904 12 4904 12 0 FILL_0__1736_.vdd
rlabel metal1 4884 242 4916 258 0 FILL_0__1736_.gnd
rlabel metal1 4944 242 5076 258 0 _1753_.gnd
rlabel metal1 4944 482 5075 498 0 _1753_.vdd
rlabel metal2 4953 353 4967 367 0 _1753_.S
rlabel metal2 4973 333 4987 347 0 _1753_.B
rlabel metal2 5013 353 5027 367 0 _1753_.Y
rlabel metal2 5033 333 5047 347 0 _1753_.A
rlabel metal1 4924 242 5036 258 0 _1736_.gnd
rlabel metal1 4924 2 5036 18 0 _1736_.vdd
rlabel metal2 5013 153 5027 167 0 _1736_.A
rlabel metal2 4993 133 5007 147 0 _1736_.B
rlabel metal2 4953 133 4967 147 0 _1736_.C
rlabel metal2 4973 153 4987 167 0 _1736_.Y
rlabel nsubstratencontact 5056 12 5056 12 0 FILL_1__1740_.vdd
rlabel metal1 5044 242 5076 258 0 FILL_1__1740_.gnd
rlabel nsubstratencontact 5036 12 5036 12 0 FILL_0__1740_.vdd
rlabel metal1 5024 242 5056 258 0 FILL_0__1740_.gnd
rlabel nsubstratencontact 5104 488 5104 488 0 FILL_1__1752_.vdd
rlabel metal1 5084 242 5116 258 0 FILL_1__1752_.gnd
rlabel nsubstratencontact 5184 12 5184 12 0 FILL_1__1726_.vdd
rlabel metal1 5164 242 5196 258 0 FILL_1__1726_.gnd
rlabel nsubstratencontact 5084 488 5084 488 0 FILL_0__1752_.vdd
rlabel metal1 5064 242 5096 258 0 FILL_0__1752_.gnd
rlabel nsubstratencontact 5164 12 5164 12 0 FILL_0__1726_.vdd
rlabel metal1 5144 242 5176 258 0 FILL_0__1726_.gnd
rlabel metal1 5104 242 5216 258 0 _1752_.gnd
rlabel metal1 5104 482 5216 498 0 _1752_.vdd
rlabel metal2 5193 333 5207 347 0 _1752_.A
rlabel metal2 5173 353 5187 367 0 _1752_.B
rlabel metal2 5133 353 5147 367 0 _1752_.C
rlabel metal2 5153 333 5167 347 0 _1752_.Y
rlabel metal1 5064 242 5156 258 0 _1740_.gnd
rlabel metal1 5064 2 5156 18 0 _1740_.vdd
rlabel metal2 5113 153 5127 167 0 _1740_.B
rlabel metal2 5073 153 5087 167 0 _1740_.A
rlabel metal2 5093 173 5107 187 0 _1740_.Y
rlabel metal1 5184 242 5276 258 0 _1726_.gnd
rlabel metal1 5184 2 5276 18 0 _1726_.vdd
rlabel metal2 5253 113 5267 127 0 _1726_.A
rlabel metal2 5213 113 5227 127 0 _1726_.B
rlabel metal2 5233 133 5247 147 0 _1726_.Y
rlabel nsubstratencontact 5256 488 5256 488 0 FILL_2__1735_.vdd
rlabel metal1 5244 242 5276 258 0 FILL_2__1735_.gnd
rlabel nsubstratencontact 5236 488 5236 488 0 FILL_1__1735_.vdd
rlabel metal1 5224 242 5256 258 0 FILL_1__1735_.gnd
rlabel nsubstratencontact 5296 12 5296 12 0 FILL_1__1725_.vdd
rlabel metal1 5284 242 5316 258 0 FILL_1__1725_.gnd
rlabel nsubstratencontact 5216 488 5216 488 0 FILL_0__1735_.vdd
rlabel metal1 5204 242 5236 258 0 FILL_0__1735_.gnd
rlabel nsubstratencontact 5276 12 5276 12 0 FILL_0__1725_.vdd
rlabel metal1 5264 242 5296 258 0 FILL_0__1725_.gnd
rlabel metal1 5264 242 5376 258 0 _1735_.gnd
rlabel metal1 5264 482 5376 498 0 _1735_.vdd
rlabel metal2 5273 333 5287 347 0 _1735_.A
rlabel metal2 5293 353 5307 367 0 _1735_.B
rlabel metal2 5333 353 5347 367 0 _1735_.C
rlabel metal2 5313 333 5327 347 0 _1735_.Y
rlabel metal1 5304 242 5436 258 0 _1725_.gnd
rlabel metal1 5304 2 5435 18 0 _1725_.vdd
rlabel metal2 5313 133 5327 147 0 _1725_.S
rlabel metal2 5333 153 5347 167 0 _1725_.B
rlabel metal2 5373 133 5387 147 0 _1725_.Y
rlabel metal2 5393 153 5407 167 0 _1725_.A
rlabel nsubstratencontact 5424 488 5424 488 0 FILL_2__1722_.vdd
rlabel metal1 5404 242 5436 258 0 FILL_2__1722_.gnd
rlabel nsubstratencontact 5456 12 5456 12 0 FILL_1__1723_.vdd
rlabel metal1 5444 242 5476 258 0 FILL_1__1723_.gnd
rlabel nsubstratencontact 5404 488 5404 488 0 FILL_1__1722_.vdd
rlabel metal1 5384 242 5416 258 0 FILL_1__1722_.gnd
rlabel nsubstratencontact 5436 12 5436 12 0 FILL_0__1723_.vdd
rlabel metal1 5424 242 5456 258 0 FILL_0__1723_.gnd
rlabel nsubstratencontact 5384 488 5384 488 0 FILL_0__1722_.vdd
rlabel metal1 5364 242 5396 258 0 FILL_0__1722_.gnd
rlabel metal1 5464 242 5536 258 0 _1723_.gnd
rlabel metal1 5464 2 5536 18 0 _1723_.vdd
rlabel metal2 5473 173 5487 187 0 _1723_.A
rlabel metal2 5493 133 5507 147 0 _1723_.Y
rlabel metal1 5424 242 5536 258 0 _1722_.gnd
rlabel metal1 5424 482 5536 498 0 _1722_.vdd
rlabel metal2 5513 353 5527 367 0 _1722_.A
rlabel metal2 5493 313 5507 327 0 _1722_.B
rlabel metal2 5473 353 5487 367 0 _1722_.C
rlabel metal2 5453 333 5467 347 0 _1722_.Y
rlabel nsubstratencontact 5556 488 5556 488 0 FILL_1__1721_.vdd
rlabel metal1 5544 242 5576 258 0 FILL_1__1721_.gnd
rlabel nsubstratencontact 5564 12 5564 12 0 FILL_1__1612_.vdd
rlabel metal1 5544 242 5576 258 0 FILL_1__1612_.gnd
rlabel nsubstratencontact 5536 488 5536 488 0 FILL_0__1721_.vdd
rlabel metal1 5524 242 5556 258 0 FILL_0__1721_.gnd
rlabel nsubstratencontact 5544 12 5544 12 0 FILL_0__1612_.vdd
rlabel metal1 5524 242 5556 258 0 FILL_0__1612_.gnd
rlabel nsubstratencontact 5656 12 5656 12 0 FILL_1__1701_.vdd
rlabel metal1 5644 242 5676 258 0 FILL_1__1701_.gnd
rlabel nsubstratencontact 5676 488 5676 488 0 FILL_0__1731_.vdd
rlabel metal1 5664 242 5696 258 0 FILL_0__1731_.gnd
rlabel nsubstratencontact 5636 12 5636 12 0 FILL_0__1701_.vdd
rlabel metal1 5624 242 5656 258 0 FILL_0__1701_.gnd
rlabel metal1 5564 242 5676 258 0 _1721_.gnd
rlabel metal1 5564 482 5676 498 0 _1721_.vdd
rlabel metal2 5573 333 5587 347 0 _1721_.A
rlabel metal2 5593 353 5607 367 0 _1721_.B
rlabel metal2 5633 353 5647 367 0 _1721_.C
rlabel metal2 5613 333 5627 347 0 _1721_.Y
rlabel metal1 5664 242 5756 258 0 _1701_.gnd
rlabel metal1 5664 2 5756 18 0 _1701_.vdd
rlabel metal2 5673 113 5687 127 0 _1701_.A
rlabel metal2 5713 113 5727 127 0 _1701_.B
rlabel metal2 5693 133 5707 147 0 _1701_.Y
rlabel metal1 5564 242 5636 258 0 _1612_.gnd
rlabel metal1 5564 2 5636 18 0 _1612_.vdd
rlabel metal2 5613 173 5627 187 0 _1612_.A
rlabel metal2 5593 133 5607 147 0 _1612_.Y
rlabel nsubstratencontact 5696 488 5696 488 0 FILL_1__1731_.vdd
rlabel metal1 5684 242 5716 258 0 FILL_1__1731_.gnd
rlabel nsubstratencontact 5796 488 5796 488 0 FILL86850x3750.vdd
rlabel metal1 5784 242 5816 258 0 FILL86850x3750.gnd
rlabel nsubstratencontact 5804 12 5804 12 0 FILL86850x150.vdd
rlabel metal1 5784 242 5816 258 0 FILL86850x150.gnd
rlabel nsubstratencontact 5784 12 5784 12 0 FILL86550x150.vdd
rlabel metal1 5764 242 5796 258 0 FILL86550x150.gnd
rlabel nsubstratencontact 5764 12 5764 12 0 FILL86250x150.vdd
rlabel metal1 5744 242 5776 258 0 FILL86250x150.gnd
rlabel metal1 5704 242 5796 258 0 _1731_.gnd
rlabel metal1 5704 482 5796 498 0 _1731_.vdd
rlabel metal2 5713 373 5727 387 0 _1731_.A
rlabel metal2 5753 373 5767 387 0 _1731_.B
rlabel metal2 5733 353 5747 367 0 _1731_.Y
rlabel nsubstratencontact 44 492 44 492 0 FILL_1__1048_.vdd
rlabel metal1 24 722 56 738 0 FILL_1__1048_.gnd
rlabel nsubstratencontact 24 492 24 492 0 FILL_0__1048_.vdd
rlabel metal1 4 722 36 738 0 FILL_0__1048_.gnd
rlabel metal1 44 722 156 738 0 _1048_.gnd
rlabel metal1 44 482 156 498 0 _1048_.vdd
rlabel metal2 133 613 147 627 0 _1048_.A
rlabel metal2 113 593 127 607 0 _1048_.B
rlabel metal2 93 613 107 627 0 _1048_.C
rlabel metal2 73 593 87 607 0 _1048_.Y
rlabel nsubstratencontact 204 492 204 492 0 FILL_2__1037_.vdd
rlabel metal1 184 722 216 738 0 FILL_2__1037_.gnd
rlabel nsubstratencontact 184 492 184 492 0 FILL_1__1037_.vdd
rlabel metal1 164 722 196 738 0 FILL_1__1037_.gnd
rlabel nsubstratencontact 164 492 164 492 0 FILL_0__1037_.vdd
rlabel metal1 144 722 176 738 0 FILL_0__1037_.gnd
rlabel metal1 204 722 316 738 0 _1037_.gnd
rlabel metal1 204 482 316 498 0 _1037_.vdd
rlabel metal2 293 613 307 627 0 _1037_.A
rlabel metal2 273 653 287 667 0 _1037_.B
rlabel metal2 253 613 267 627 0 _1037_.C
rlabel metal2 233 633 247 647 0 _1037_.Y
rlabel nsubstratencontact 344 492 344 492 0 FILL_1__1028_.vdd
rlabel metal1 324 722 356 738 0 FILL_1__1028_.gnd
rlabel nsubstratencontact 324 492 324 492 0 FILL_0__1028_.vdd
rlabel metal1 304 722 336 738 0 FILL_0__1028_.gnd
rlabel metal1 344 722 456 738 0 _1028_.gnd
rlabel metal1 344 482 456 498 0 _1028_.vdd
rlabel metal2 433 613 447 627 0 _1028_.A
rlabel metal2 413 593 427 607 0 _1028_.B
rlabel metal2 393 613 407 627 0 _1028_.C
rlabel metal2 373 593 387 607 0 _1028_.Y
rlabel nsubstratencontact 484 492 484 492 0 FILL_1__1035_.vdd
rlabel metal1 464 722 496 738 0 FILL_1__1035_.gnd
rlabel nsubstratencontact 464 492 464 492 0 FILL_0__1035_.vdd
rlabel metal1 444 722 476 738 0 FILL_0__1035_.gnd
rlabel metal1 484 722 596 738 0 _1035_.gnd
rlabel metal1 484 482 596 498 0 _1035_.vdd
rlabel metal2 573 633 587 647 0 _1035_.A
rlabel metal2 553 613 567 627 0 _1035_.B
rlabel metal2 513 613 527 627 0 _1035_.C
rlabel metal2 533 633 547 647 0 _1035_.Y
rlabel nsubstratencontact 616 492 616 492 0 FILL_1__1095_.vdd
rlabel metal1 604 722 636 738 0 FILL_1__1095_.gnd
rlabel nsubstratencontact 596 492 596 492 0 FILL_0__1095_.vdd
rlabel metal1 584 722 616 738 0 FILL_0__1095_.gnd
rlabel metal1 624 722 736 738 0 _1095_.gnd
rlabel metal1 624 482 736 498 0 _1095_.vdd
rlabel metal2 633 613 647 627 0 _1095_.A
rlabel metal2 653 653 667 667 0 _1095_.B
rlabel metal2 673 613 687 627 0 _1095_.C
rlabel metal2 693 633 707 647 0 _1095_.Y
rlabel nsubstratencontact 756 492 756 492 0 FILL_1__1027_.vdd
rlabel metal1 744 722 776 738 0 FILL_1__1027_.gnd
rlabel nsubstratencontact 736 492 736 492 0 FILL_0__1027_.vdd
rlabel metal1 724 722 756 738 0 FILL_0__1027_.gnd
rlabel nsubstratencontact 884 492 884 492 0 FILL_1__1096_.vdd
rlabel metal1 864 722 896 738 0 FILL_1__1096_.gnd
rlabel nsubstratencontact 864 492 864 492 0 FILL_0__1096_.vdd
rlabel metal1 844 722 876 738 0 FILL_0__1096_.gnd
rlabel metal1 764 722 856 738 0 _1027_.gnd
rlabel metal1 764 482 856 498 0 _1027_.vdd
rlabel metal2 773 593 787 607 0 _1027_.A
rlabel metal2 813 593 827 607 0 _1027_.B
rlabel metal2 793 613 807 627 0 _1027_.Y
rlabel nsubstratencontact 904 492 904 492 0 FILL_2__1096_.vdd
rlabel metal1 884 722 916 738 0 FILL_2__1096_.gnd
rlabel nsubstratencontact 1024 492 1024 492 0 FILL_0__1086_.vdd
rlabel metal1 1004 722 1036 738 0 FILL_0__1086_.gnd
rlabel metal1 904 722 1016 738 0 _1096_.gnd
rlabel metal1 904 482 1016 498 0 _1096_.vdd
rlabel metal2 993 633 1007 647 0 _1096_.A
rlabel metal2 973 613 987 627 0 _1096_.B
rlabel metal2 933 613 947 627 0 _1096_.C
rlabel metal2 953 633 967 647 0 _1096_.Y
rlabel nsubstratencontact 1044 492 1044 492 0 FILL_1__1086_.vdd
rlabel metal1 1024 722 1056 738 0 FILL_1__1086_.gnd
rlabel metal1 1044 722 1156 738 0 _1086_.gnd
rlabel metal1 1044 482 1156 498 0 _1086_.vdd
rlabel metal2 1133 613 1147 627 0 _1086_.A
rlabel metal2 1113 593 1127 607 0 _1086_.B
rlabel metal2 1093 613 1107 627 0 _1086_.C
rlabel metal2 1073 593 1087 607 0 _1086_.Y
rlabel nsubstratencontact 1176 492 1176 492 0 FILL_1__1209_.vdd
rlabel metal1 1164 722 1196 738 0 FILL_1__1209_.gnd
rlabel nsubstratencontact 1156 492 1156 492 0 FILL_0__1209_.vdd
rlabel metal1 1144 722 1176 738 0 FILL_0__1209_.gnd
rlabel metal1 1184 722 1296 738 0 _1209_.gnd
rlabel metal1 1184 482 1296 498 0 _1209_.vdd
rlabel metal2 1193 613 1207 627 0 _1209_.A
rlabel metal2 1213 653 1227 667 0 _1209_.B
rlabel metal2 1233 613 1247 627 0 _1209_.C
rlabel metal2 1253 633 1267 647 0 _1209_.Y
rlabel nsubstratencontact 1324 492 1324 492 0 FILL_1__1088_.vdd
rlabel metal1 1304 722 1336 738 0 FILL_1__1088_.gnd
rlabel nsubstratencontact 1304 492 1304 492 0 FILL_0__1088_.vdd
rlabel metal1 1284 722 1316 738 0 FILL_0__1088_.gnd
rlabel metal1 1324 722 1436 738 0 _1088_.gnd
rlabel metal1 1324 482 1436 498 0 _1088_.vdd
rlabel metal2 1413 613 1427 627 0 _1088_.A
rlabel metal2 1393 653 1407 667 0 _1088_.B
rlabel metal2 1373 613 1387 627 0 _1088_.C
rlabel metal2 1353 633 1367 647 0 _1088_.Y
rlabel nsubstratencontact 1476 492 1476 492 0 FILL_2__1069_.vdd
rlabel metal1 1464 722 1496 738 0 FILL_2__1069_.gnd
rlabel nsubstratencontact 1456 492 1456 492 0 FILL_1__1069_.vdd
rlabel metal1 1444 722 1476 738 0 FILL_1__1069_.gnd
rlabel nsubstratencontact 1436 492 1436 492 0 FILL_0__1069_.vdd
rlabel metal1 1424 722 1456 738 0 FILL_0__1069_.gnd
rlabel metal1 1484 722 1596 738 0 _1069_.gnd
rlabel metal1 1484 482 1596 498 0 _1069_.vdd
rlabel metal2 1493 613 1507 627 0 _1069_.A
rlabel metal2 1513 593 1527 607 0 _1069_.B
rlabel metal2 1533 613 1547 627 0 _1069_.C
rlabel metal2 1553 593 1567 607 0 _1069_.Y
rlabel nsubstratencontact 1624 492 1624 492 0 FILL_1__1064_.vdd
rlabel metal1 1604 722 1636 738 0 FILL_1__1064_.gnd
rlabel nsubstratencontact 1604 492 1604 492 0 FILL_0__1064_.vdd
rlabel metal1 1584 722 1616 738 0 FILL_0__1064_.gnd
rlabel metal1 1624 722 1736 738 0 _1064_.gnd
rlabel metal1 1624 482 1736 498 0 _1064_.vdd
rlabel metal2 1713 633 1727 647 0 _1064_.A
rlabel metal2 1693 613 1707 627 0 _1064_.B
rlabel metal2 1653 613 1667 627 0 _1064_.C
rlabel metal2 1673 633 1687 647 0 _1064_.Y
rlabel nsubstratencontact 1764 492 1764 492 0 FILL_1__1068_.vdd
rlabel metal1 1744 722 1776 738 0 FILL_1__1068_.gnd
rlabel nsubstratencontact 1744 492 1744 492 0 FILL_0__1068_.vdd
rlabel metal1 1724 722 1756 738 0 FILL_0__1068_.gnd
rlabel metal1 1764 722 1876 738 0 _1068_.gnd
rlabel metal1 1764 482 1876 498 0 _1068_.vdd
rlabel metal2 1853 613 1867 627 0 _1068_.A
rlabel metal2 1833 593 1847 607 0 _1068_.B
rlabel metal2 1813 613 1827 627 0 _1068_.C
rlabel metal2 1793 593 1807 607 0 _1068_.Y
rlabel nsubstratencontact 1896 492 1896 492 0 FILL_1__1221_.vdd
rlabel metal1 1884 722 1916 738 0 FILL_1__1221_.gnd
rlabel nsubstratencontact 1876 492 1876 492 0 FILL_0__1221_.vdd
rlabel metal1 1864 722 1896 738 0 FILL_0__1221_.gnd
rlabel nsubstratencontact 2024 492 2024 492 0 FILL_0__1060_.vdd
rlabel metal1 2004 722 2036 738 0 FILL_0__1060_.gnd
rlabel metal1 1904 722 2016 738 0 _1221_.gnd
rlabel metal1 1904 482 2016 498 0 _1221_.vdd
rlabel metal2 1913 613 1927 627 0 _1221_.A
rlabel metal2 1933 653 1947 667 0 _1221_.B
rlabel metal2 1953 613 1967 627 0 _1221_.C
rlabel metal2 1973 633 1987 647 0 _1221_.Y
rlabel nsubstratencontact 2164 492 2164 492 0 FILL_1__1065_.vdd
rlabel metal1 2144 722 2176 738 0 FILL_1__1065_.gnd
rlabel nsubstratencontact 2044 492 2044 492 0 FILL_1__1060_.vdd
rlabel metal1 2024 722 2056 738 0 FILL_1__1060_.gnd
rlabel nsubstratencontact 2144 492 2144 492 0 FILL_0__1065_.vdd
rlabel metal1 2124 722 2156 738 0 FILL_0__1065_.gnd
rlabel metal1 2044 722 2136 738 0 _1060_.gnd
rlabel metal1 2044 482 2136 498 0 _1060_.vdd
rlabel metal2 2073 633 2087 647 0 _1060_.B
rlabel metal2 2113 633 2127 647 0 _1060_.A
rlabel metal2 2093 653 2107 667 0 _1060_.Y
rlabel nsubstratencontact 2276 492 2276 492 0 FILL_0__1889_.vdd
rlabel metal1 2264 722 2296 738 0 FILL_0__1889_.gnd
rlabel metal1 2164 722 2276 738 0 _1065_.gnd
rlabel metal1 2164 482 2276 498 0 _1065_.vdd
rlabel metal2 2253 653 2267 667 0 _1065_.A
rlabel metal2 2233 633 2247 647 0 _1065_.B
rlabel metal2 2193 613 2207 627 0 _1065_.Y
rlabel nsubstratencontact 2296 492 2296 492 0 FILL_1__1889_.vdd
rlabel metal1 2284 722 2316 738 0 FILL_1__1889_.gnd
rlabel metal1 2304 722 2416 738 0 _1889_.gnd
rlabel metal1 2304 482 2416 498 0 _1889_.vdd
rlabel metal2 2313 633 2327 647 0 _1889_.A
rlabel metal2 2373 633 2387 647 0 _1889_.Y
rlabel metal2 2353 593 2367 607 0 _1889_.B
rlabel nsubstratencontact 2436 492 2436 492 0 FILL_1__1888_.vdd
rlabel metal1 2424 722 2456 738 0 FILL_1__1888_.gnd
rlabel nsubstratencontact 2416 492 2416 492 0 FILL_0__1888_.vdd
rlabel metal1 2404 722 2436 738 0 FILL_0__1888_.gnd
rlabel metal1 2444 722 2536 738 0 _1888_.gnd
rlabel metal1 2444 482 2536 498 0 _1888_.vdd
rlabel metal2 2453 593 2467 607 0 _1888_.A
rlabel metal2 2493 593 2507 607 0 _1888_.B
rlabel metal2 2473 613 2487 627 0 _1888_.Y
rlabel nsubstratencontact 2544 492 2544 492 0 FILL_0__1830_.vdd
rlabel metal1 2524 722 2556 738 0 FILL_0__1830_.gnd
rlabel nsubstratencontact 2564 492 2564 492 0 FILL_1__1830_.vdd
rlabel metal1 2544 722 2576 738 0 FILL_1__1830_.gnd
rlabel nsubstratencontact 2664 492 2664 492 0 FILL_0__1853_.vdd
rlabel metal1 2644 722 2676 738 0 FILL_0__1853_.gnd
rlabel metal1 2564 722 2656 738 0 _1830_.gnd
rlabel metal1 2564 482 2656 498 0 _1830_.vdd
rlabel metal2 2633 593 2647 607 0 _1830_.A
rlabel metal2 2593 593 2607 607 0 _1830_.B
rlabel metal2 2613 613 2627 627 0 _1830_.Y
rlabel nsubstratencontact 2684 492 2684 492 0 FILL_1__1853_.vdd
rlabel metal1 2664 722 2696 738 0 FILL_1__1853_.gnd
rlabel nsubstratencontact 2776 492 2776 492 0 FILL_0__1854_.vdd
rlabel metal1 2764 722 2796 738 0 FILL_0__1854_.gnd
rlabel metal1 2684 722 2776 738 0 _1853_.gnd
rlabel metal1 2684 482 2776 498 0 _1853_.vdd
rlabel metal2 2713 633 2727 647 0 _1853_.B
rlabel metal2 2753 633 2767 647 0 _1853_.A
rlabel metal2 2733 653 2747 667 0 _1853_.Y
rlabel nsubstratencontact 2796 492 2796 492 0 FILL_1__1854_.vdd
rlabel metal1 2784 722 2816 738 0 FILL_1__1854_.gnd
rlabel metal1 2804 722 2916 738 0 _1854_.gnd
rlabel metal1 2804 482 2916 498 0 _1854_.vdd
rlabel metal2 2813 633 2827 647 0 _1854_.A
rlabel metal2 2833 613 2847 627 0 _1854_.B
rlabel metal2 2873 613 2887 627 0 _1854_.C
rlabel metal2 2853 633 2867 647 0 _1854_.Y
rlabel nsubstratencontact 2944 492 2944 492 0 FILL_1__1832_.vdd
rlabel metal1 2924 722 2956 738 0 FILL_1__1832_.gnd
rlabel nsubstratencontact 3036 492 3036 492 0 FILL_0__1871_.vdd
rlabel metal1 3024 722 3056 738 0 FILL_0__1871_.gnd
rlabel nsubstratencontact 2924 492 2924 492 0 FILL_0__1832_.vdd
rlabel metal1 2904 722 2936 738 0 FILL_0__1832_.gnd
rlabel metal1 2944 722 3036 738 0 _1832_.gnd
rlabel metal1 2944 482 3036 498 0 _1832_.vdd
rlabel metal2 3013 593 3027 607 0 _1832_.A
rlabel metal2 2973 593 2987 607 0 _1832_.B
rlabel metal2 2993 613 3007 627 0 _1832_.Y
rlabel nsubstratencontact 3056 492 3056 492 0 FILL_1__1871_.vdd
rlabel metal1 3044 722 3076 738 0 FILL_1__1871_.gnd
rlabel metal1 3064 722 3176 738 0 _1871_.gnd
rlabel metal1 3064 482 3176 498 0 _1871_.vdd
rlabel metal2 3073 613 3087 627 0 _1871_.A
rlabel metal2 3093 653 3107 667 0 _1871_.B
rlabel metal2 3113 613 3127 627 0 _1871_.C
rlabel metal2 3133 633 3147 647 0 _1871_.Y
rlabel nsubstratencontact 3204 492 3204 492 0 FILL_1__1831_.vdd
rlabel metal1 3184 722 3216 738 0 FILL_1__1831_.gnd
rlabel nsubstratencontact 3184 492 3184 492 0 FILL_0__1831_.vdd
rlabel metal1 3164 722 3196 738 0 FILL_0__1831_.gnd
rlabel metal1 3204 722 3316 738 0 _1831_.gnd
rlabel metal1 3204 482 3316 498 0 _1831_.vdd
rlabel metal2 3293 613 3307 627 0 _1831_.A
rlabel metal2 3273 593 3287 607 0 _1831_.B
rlabel metal2 3253 613 3267 627 0 _1831_.C
rlabel metal2 3233 593 3247 607 0 _1831_.Y
rlabel nsubstratencontact 3336 492 3336 492 0 FILL_1__1816_.vdd
rlabel metal1 3324 722 3356 738 0 FILL_1__1816_.gnd
rlabel nsubstratencontact 3316 492 3316 492 0 FILL_0__1816_.vdd
rlabel metal1 3304 722 3336 738 0 FILL_0__1816_.gnd
rlabel metal1 3344 722 3436 738 0 _1816_.gnd
rlabel metal1 3344 482 3436 498 0 _1816_.vdd
rlabel metal2 3353 593 3367 607 0 _1816_.A
rlabel metal2 3393 593 3407 607 0 _1816_.B
rlabel metal2 3373 613 3387 627 0 _1816_.Y
rlabel nsubstratencontact 3464 492 3464 492 0 FILL_1__1818_.vdd
rlabel metal1 3444 722 3476 738 0 FILL_1__1818_.gnd
rlabel nsubstratencontact 3444 492 3444 492 0 FILL_0__1818_.vdd
rlabel metal1 3424 722 3456 738 0 FILL_0__1818_.gnd
rlabel metal1 3464 722 3576 738 0 _1818_.gnd
rlabel metal1 3464 482 3576 498 0 _1818_.vdd
rlabel metal2 3553 633 3567 647 0 _1818_.A
rlabel metal2 3533 613 3547 627 0 _1818_.B
rlabel metal2 3493 613 3507 627 0 _1818_.C
rlabel metal2 3513 633 3527 647 0 _1818_.Y
rlabel nsubstratencontact 3596 492 3596 492 0 FILL_1__1815_.vdd
rlabel metal1 3584 722 3616 738 0 FILL_1__1815_.gnd
rlabel nsubstratencontact 3576 492 3576 492 0 FILL_0__1815_.vdd
rlabel metal1 3564 722 3596 738 0 FILL_0__1815_.gnd
rlabel metal1 3604 722 3696 738 0 _1815_.gnd
rlabel metal1 3604 482 3696 498 0 _1815_.vdd
rlabel metal2 3613 593 3627 607 0 _1815_.A
rlabel metal2 3653 593 3667 607 0 _1815_.B
rlabel metal2 3633 613 3647 627 0 _1815_.Y
rlabel nsubstratencontact 3724 492 3724 492 0 FILL_1__1845_.vdd
rlabel metal1 3704 722 3736 738 0 FILL_1__1845_.gnd
rlabel nsubstratencontact 3704 492 3704 492 0 FILL_0__1845_.vdd
rlabel metal1 3684 722 3716 738 0 FILL_0__1845_.gnd
rlabel metal1 3724 722 3836 738 0 _1845_.gnd
rlabel metal1 3724 482 3836 498 0 _1845_.vdd
rlabel metal2 3813 633 3827 647 0 _1845_.A
rlabel metal2 3793 613 3807 627 0 _1845_.B
rlabel metal2 3753 613 3767 627 0 _1845_.C
rlabel metal2 3773 633 3787 647 0 _1845_.Y
rlabel nsubstratencontact 3856 492 3856 492 0 FILL_1__1844_.vdd
rlabel metal1 3844 722 3876 738 0 FILL_1__1844_.gnd
rlabel nsubstratencontact 3836 492 3836 492 0 FILL_0__1844_.vdd
rlabel metal1 3824 722 3856 738 0 FILL_0__1844_.gnd
rlabel metal1 3864 722 3976 738 0 _1844_.gnd
rlabel metal1 3864 482 3976 498 0 _1844_.vdd
rlabel metal2 3873 633 3887 647 0 _1844_.A
rlabel metal2 3893 613 3907 627 0 _1844_.B
rlabel metal2 3933 613 3947 627 0 _1844_.C
rlabel metal2 3913 633 3927 647 0 _1844_.Y
rlabel nsubstratencontact 3996 492 3996 492 0 FILL_1__1793_.vdd
rlabel metal1 3984 722 4016 738 0 FILL_1__1793_.gnd
rlabel nsubstratencontact 3976 492 3976 492 0 FILL_0__1793_.vdd
rlabel metal1 3964 722 3996 738 0 FILL_0__1793_.gnd
rlabel metal1 4004 722 4116 738 0 _1793_.gnd
rlabel metal1 4004 482 4116 498 0 _1793_.vdd
rlabel metal2 4013 613 4027 627 0 _1793_.A
rlabel metal2 4033 653 4047 667 0 _1793_.B
rlabel metal2 4053 613 4067 627 0 _1793_.C
rlabel metal2 4073 633 4087 647 0 _1793_.Y
rlabel nsubstratencontact 4156 492 4156 492 0 FILL_2__1813_.vdd
rlabel metal1 4144 722 4176 738 0 FILL_2__1813_.gnd
rlabel nsubstratencontact 4136 492 4136 492 0 FILL_1__1813_.vdd
rlabel metal1 4124 722 4156 738 0 FILL_1__1813_.gnd
rlabel nsubstratencontact 4116 492 4116 492 0 FILL_0__1813_.vdd
rlabel metal1 4104 722 4136 738 0 FILL_0__1813_.gnd
rlabel metal1 4164 722 4276 738 0 _1813_.gnd
rlabel metal1 4164 482 4276 498 0 _1813_.vdd
rlabel metal2 4173 633 4187 647 0 _1813_.A
rlabel metal2 4193 613 4207 627 0 _1813_.B
rlabel metal2 4233 613 4247 627 0 _1813_.C
rlabel metal2 4213 633 4227 647 0 _1813_.Y
rlabel nsubstratencontact 4304 492 4304 492 0 FILL_1__1812_.vdd
rlabel metal1 4284 722 4316 738 0 FILL_1__1812_.gnd
rlabel nsubstratencontact 4284 492 4284 492 0 FILL_0__1812_.vdd
rlabel metal1 4264 722 4296 738 0 FILL_0__1812_.gnd
rlabel nsubstratencontact 4404 492 4404 492 0 FILL_1__1782_.vdd
rlabel metal1 4384 722 4416 738 0 FILL_1__1782_.gnd
rlabel nsubstratencontact 4384 492 4384 492 0 FILL_0__1782_.vdd
rlabel metal1 4364 722 4396 738 0 FILL_0__1782_.gnd
rlabel metal1 4304 722 4376 738 0 _1812_.gnd
rlabel metal1 4304 482 4376 498 0 _1812_.vdd
rlabel metal2 4353 653 4367 667 0 _1812_.A
rlabel metal2 4333 613 4347 627 0 _1812_.Y
rlabel metal1 4404 722 4516 738 0 _1782_.gnd
rlabel metal1 4404 482 4516 498 0 _1782_.vdd
rlabel metal2 4493 613 4507 627 0 _1782_.A
rlabel metal2 4473 653 4487 667 0 _1782_.B
rlabel metal2 4453 613 4467 627 0 _1782_.C
rlabel metal2 4433 633 4447 647 0 _1782_.Y
rlabel nsubstratencontact 4544 492 4544 492 0 FILL_1__1811_.vdd
rlabel metal1 4524 722 4556 738 0 FILL_1__1811_.gnd
rlabel nsubstratencontact 4524 492 4524 492 0 FILL_0__1811_.vdd
rlabel metal1 4504 722 4536 738 0 FILL_0__1811_.gnd
rlabel metal1 4544 722 4656 738 0 _1811_.gnd
rlabel metal1 4544 482 4656 498 0 _1811_.vdd
rlabel metal2 4633 633 4647 647 0 _1811_.A
rlabel metal2 4613 613 4627 627 0 _1811_.B
rlabel metal2 4573 613 4587 627 0 _1811_.C
rlabel metal2 4593 633 4607 647 0 _1811_.Y
rlabel nsubstratencontact 4684 492 4684 492 0 FILL_1__1810_.vdd
rlabel metal1 4664 722 4696 738 0 FILL_1__1810_.gnd
rlabel nsubstratencontact 4664 492 4664 492 0 FILL_0__1810_.vdd
rlabel metal1 4644 722 4676 738 0 FILL_0__1810_.gnd
rlabel nsubstratencontact 4796 492 4796 492 0 FILL_0__1755_.vdd
rlabel metal1 4784 722 4816 738 0 FILL_0__1755_.gnd
rlabel metal1 4684 722 4796 738 0 _1810_.gnd
rlabel metal1 4684 482 4796 498 0 _1810_.vdd
rlabel metal2 4773 633 4787 647 0 _1810_.A
rlabel metal2 4753 613 4767 627 0 _1810_.B
rlabel metal2 4713 613 4727 627 0 _1810_.C
rlabel metal2 4733 633 4747 647 0 _1810_.Y
rlabel nsubstratencontact 4836 492 4836 492 0 FILL_2__1755_.vdd
rlabel metal1 4824 722 4856 738 0 FILL_2__1755_.gnd
rlabel nsubstratencontact 4816 492 4816 492 0 FILL_1__1755_.vdd
rlabel metal1 4804 722 4836 738 0 FILL_1__1755_.gnd
rlabel metal1 4844 722 4956 738 0 _1755_.gnd
rlabel metal1 4844 482 4956 498 0 _1755_.vdd
rlabel metal2 4853 633 4867 647 0 _1755_.A
rlabel metal2 4873 613 4887 627 0 _1755_.B
rlabel metal2 4913 613 4927 627 0 _1755_.C
rlabel metal2 4893 633 4907 647 0 _1755_.Y
rlabel nsubstratencontact 4976 492 4976 492 0 FILL_1__1751_.vdd
rlabel metal1 4964 722 4996 738 0 FILL_1__1751_.gnd
rlabel nsubstratencontact 5056 492 5056 492 0 FILL_0_BUFX2_insert14.vdd
rlabel metal1 5044 722 5076 738 0 FILL_0_BUFX2_insert14.gnd
rlabel nsubstratencontact 4956 492 4956 492 0 FILL_0__1751_.vdd
rlabel metal1 4944 722 4976 738 0 FILL_0__1751_.gnd
rlabel metal1 4984 722 5056 738 0 _1751_.gnd
rlabel metal1 4984 482 5056 498 0 _1751_.vdd
rlabel metal2 4993 653 5007 667 0 _1751_.A
rlabel metal2 5013 613 5027 627 0 _1751_.Y
rlabel nsubstratencontact 5096 492 5096 492 0 FILL_2_BUFX2_insert14.vdd
rlabel metal1 5084 722 5116 738 0 FILL_2_BUFX2_insert14.gnd
rlabel nsubstratencontact 5076 492 5076 492 0 FILL_1_BUFX2_insert14.vdd
rlabel metal1 5064 722 5096 738 0 FILL_1_BUFX2_insert14.gnd
rlabel metal1 5104 722 5196 738 0 BUFX2_insert14.gnd
rlabel metal1 5104 482 5196 498 0 BUFX2_insert14.vdd
rlabel metal2 5113 633 5127 647 0 BUFX2_insert14.A
rlabel metal2 5153 633 5167 647 0 BUFX2_insert14.Y
rlabel nsubstratencontact 5224 492 5224 492 0 FILL_1__1713_.vdd
rlabel metal1 5204 722 5236 738 0 FILL_1__1713_.gnd
rlabel nsubstratencontact 5204 492 5204 492 0 FILL_0__1713_.vdd
rlabel metal1 5184 722 5216 738 0 FILL_0__1713_.gnd
rlabel metal1 5224 722 5336 738 0 _1713_.gnd
rlabel metal1 5224 482 5336 498 0 _1713_.vdd
rlabel metal2 5313 633 5327 647 0 _1713_.A
rlabel metal2 5293 613 5307 627 0 _1713_.B
rlabel metal2 5253 613 5267 627 0 _1713_.C
rlabel metal2 5273 633 5287 647 0 _1713_.Y
rlabel nsubstratencontact 5356 492 5356 492 0 FILL_1__1706_.vdd
rlabel metal1 5344 722 5376 738 0 FILL_1__1706_.gnd
rlabel nsubstratencontact 5336 492 5336 492 0 FILL_0__1706_.vdd
rlabel metal1 5324 722 5356 738 0 FILL_0__1706_.gnd
rlabel metal1 5364 722 5476 738 0 _1706_.gnd
rlabel metal1 5364 482 5476 498 0 _1706_.vdd
rlabel metal2 5373 633 5387 647 0 _1706_.A
rlabel metal2 5393 613 5407 627 0 _1706_.B
rlabel metal2 5433 613 5447 627 0 _1706_.C
rlabel metal2 5413 633 5427 647 0 _1706_.Y
rlabel nsubstratencontact 5504 492 5504 492 0 FILL_1__1707_.vdd
rlabel metal1 5484 722 5516 738 0 FILL_1__1707_.gnd
rlabel nsubstratencontact 5484 492 5484 492 0 FILL_0__1707_.vdd
rlabel metal1 5464 722 5496 738 0 FILL_0__1707_.gnd
rlabel metal1 5504 722 5616 738 0 _1707_.gnd
rlabel metal1 5504 482 5616 498 0 _1707_.vdd
rlabel metal2 5593 633 5607 647 0 _1707_.A
rlabel metal2 5573 613 5587 627 0 _1707_.B
rlabel metal2 5533 613 5547 627 0 _1707_.C
rlabel metal2 5553 633 5567 647 0 _1707_.Y
rlabel metal1 5644 722 5736 738 0 _1712_.gnd
rlabel metal1 5644 482 5736 498 0 _1712_.vdd
rlabel metal2 5693 633 5707 647 0 _1712_.B
rlabel metal2 5653 633 5667 647 0 _1712_.A
rlabel metal2 5673 653 5687 667 0 _1712_.Y
rlabel nsubstratencontact 5744 492 5744 492 0 FILL85950x7350.vdd
rlabel metal1 5724 722 5756 738 0 FILL85950x7350.gnd
rlabel nsubstratencontact 5764 492 5764 492 0 FILL86250x7350.vdd
rlabel metal1 5744 722 5776 738 0 FILL86250x7350.gnd
rlabel nsubstratencontact 5784 492 5784 492 0 FILL86550x7350.vdd
rlabel metal1 5764 722 5796 738 0 FILL86550x7350.gnd
rlabel nsubstratencontact 5804 492 5804 492 0 FILL86850x7350.vdd
rlabel metal1 5784 722 5816 738 0 FILL86850x7350.gnd
rlabel nsubstratencontact 5616 492 5616 492 0 FILL_0__1712_.vdd
rlabel metal1 5604 722 5636 738 0 FILL_0__1712_.gnd
rlabel nsubstratencontact 5636 492 5636 492 0 FILL_1__1712_.vdd
rlabel metal1 5624 722 5656 738 0 FILL_1__1712_.gnd
rlabel nsubstratencontact 44 968 44 968 0 FILL_1__1049_.vdd
rlabel metal1 24 722 56 738 0 FILL_1__1049_.gnd
rlabel nsubstratencontact 24 968 24 968 0 FILL_0__1049_.vdd
rlabel metal1 4 722 36 738 0 FILL_0__1049_.gnd
rlabel metal1 44 722 156 738 0 _1049_.gnd
rlabel metal1 44 962 156 978 0 _1049_.vdd
rlabel metal2 133 833 147 847 0 _1049_.A
rlabel metal2 113 853 127 867 0 _1049_.B
rlabel metal2 93 833 107 847 0 _1049_.C
rlabel metal2 73 853 87 867 0 _1049_.Y
rlabel nsubstratencontact 176 968 176 968 0 FILL_1__1033_.vdd
rlabel metal1 164 722 196 738 0 FILL_1__1033_.gnd
rlabel nsubstratencontact 156 968 156 968 0 FILL_0__1033_.vdd
rlabel metal1 144 722 176 738 0 FILL_0__1033_.gnd
rlabel metal1 184 722 296 738 0 _1033_.gnd
rlabel metal1 184 962 296 978 0 _1033_.vdd
rlabel metal2 193 833 207 847 0 _1033_.A
rlabel metal2 213 793 227 807 0 _1033_.B
rlabel metal2 233 833 247 847 0 _1033_.C
rlabel metal2 253 813 267 827 0 _1033_.Y
rlabel nsubstratencontact 324 968 324 968 0 FILL_1__1114_.vdd
rlabel metal1 304 722 336 738 0 FILL_1__1114_.gnd
rlabel nsubstratencontact 304 968 304 968 0 FILL_0__1114_.vdd
rlabel metal1 284 722 316 738 0 FILL_0__1114_.gnd
rlabel metal1 324 722 436 738 0 _1114_.gnd
rlabel metal1 324 962 436 978 0 _1114_.vdd
rlabel metal2 413 833 427 847 0 _1114_.A
rlabel metal2 393 853 407 867 0 _1114_.B
rlabel metal2 373 833 387 847 0 _1114_.C
rlabel metal2 353 853 367 867 0 _1114_.Y
rlabel nsubstratencontact 464 968 464 968 0 FILL_1__1094_.vdd
rlabel metal1 444 722 476 738 0 FILL_1__1094_.gnd
rlabel nsubstratencontact 444 968 444 968 0 FILL_0__1094_.vdd
rlabel metal1 424 722 456 738 0 FILL_0__1094_.gnd
rlabel metal1 464 722 576 738 0 _1094_.gnd
rlabel metal1 464 962 576 978 0 _1094_.vdd
rlabel metal2 553 833 567 847 0 _1094_.A
rlabel metal2 533 793 547 807 0 _1094_.B
rlabel metal2 513 833 527 847 0 _1094_.C
rlabel metal2 493 813 507 827 0 _1094_.Y
rlabel nsubstratencontact 604 968 604 968 0 FILL_1__1113_.vdd
rlabel metal1 584 722 616 738 0 FILL_1__1113_.gnd
rlabel nsubstratencontact 584 968 584 968 0 FILL_0__1113_.vdd
rlabel metal1 564 722 596 738 0 FILL_0__1113_.gnd
rlabel metal1 604 722 716 738 0 _1113_.gnd
rlabel metal1 604 962 716 978 0 _1113_.vdd
rlabel metal2 693 833 707 847 0 _1113_.A
rlabel metal2 673 853 687 867 0 _1113_.B
rlabel metal2 653 833 667 847 0 _1113_.C
rlabel metal2 633 853 647 867 0 _1113_.Y
rlabel nsubstratencontact 736 968 736 968 0 FILL_1__1098_.vdd
rlabel metal1 724 722 756 738 0 FILL_1__1098_.gnd
rlabel nsubstratencontact 716 968 716 968 0 FILL_0__1098_.vdd
rlabel metal1 704 722 736 738 0 FILL_0__1098_.gnd
rlabel metal1 744 722 856 738 0 _1098_.gnd
rlabel metal1 744 962 856 978 0 _1098_.vdd
rlabel metal2 753 833 767 847 0 _1098_.A
rlabel metal2 773 793 787 807 0 _1098_.B
rlabel metal2 793 833 807 847 0 _1098_.C
rlabel metal2 813 813 827 827 0 _1098_.Y
rlabel nsubstratencontact 884 968 884 968 0 FILL_1__1093_.vdd
rlabel metal1 864 722 896 738 0 FILL_1__1093_.gnd
rlabel nsubstratencontact 864 968 864 968 0 FILL_0__1093_.vdd
rlabel metal1 844 722 876 738 0 FILL_0__1093_.gnd
rlabel nsubstratencontact 1024 968 1024 968 0 FILL_1__1097_.vdd
rlabel metal1 1004 722 1036 738 0 FILL_1__1097_.gnd
rlabel nsubstratencontact 1004 968 1004 968 0 FILL_0__1097_.vdd
rlabel metal1 984 722 1016 738 0 FILL_0__1097_.gnd
rlabel metal1 884 722 996 738 0 _1093_.gnd
rlabel metal1 884 962 996 978 0 _1093_.vdd
rlabel metal2 973 813 987 827 0 _1093_.A
rlabel metal2 953 833 967 847 0 _1093_.B
rlabel metal2 913 833 927 847 0 _1093_.C
rlabel metal2 933 813 947 827 0 _1093_.Y
rlabel nsubstratencontact 1136 968 1136 968 0 FILL_0__1236_.vdd
rlabel metal1 1124 722 1156 738 0 FILL_0__1236_.gnd
rlabel metal1 1024 722 1136 738 0 _1097_.gnd
rlabel metal1 1024 962 1136 978 0 _1097_.vdd
rlabel metal2 1113 833 1127 847 0 _1097_.A
rlabel metal2 1093 853 1107 867 0 _1097_.B
rlabel metal2 1073 833 1087 847 0 _1097_.C
rlabel metal2 1053 853 1067 867 0 _1097_.Y
rlabel nsubstratencontact 1156 968 1156 968 0 FILL_1__1236_.vdd
rlabel metal1 1144 722 1176 738 0 FILL_1__1236_.gnd
rlabel metal1 1164 722 1276 738 0 _1236_.gnd
rlabel metal1 1164 962 1276 978 0 _1236_.vdd
rlabel metal2 1173 813 1187 827 0 _1236_.A
rlabel metal2 1193 833 1207 847 0 _1236_.B
rlabel metal2 1233 833 1247 847 0 _1236_.C
rlabel metal2 1213 813 1227 827 0 _1236_.Y
rlabel nsubstratencontact 1304 968 1304 968 0 FILL_1__1026_.vdd
rlabel metal1 1284 722 1316 738 0 FILL_1__1026_.gnd
rlabel nsubstratencontact 1284 968 1284 968 0 FILL_0__1026_.vdd
rlabel metal1 1264 722 1296 738 0 FILL_0__1026_.gnd
rlabel metal1 1304 722 1416 738 0 _1026_.gnd
rlabel metal1 1304 962 1416 978 0 _1026_.vdd
rlabel metal2 1393 833 1407 847 0 _1026_.A
rlabel metal2 1373 853 1387 867 0 _1026_.B
rlabel metal2 1353 833 1367 847 0 _1026_.C
rlabel metal2 1333 853 1347 867 0 _1026_.Y
rlabel nsubstratencontact 1436 968 1436 968 0 FILL_1__1023_.vdd
rlabel metal1 1424 722 1456 738 0 FILL_1__1023_.gnd
rlabel nsubstratencontact 1516 968 1516 968 0 FILL_0__1025_.vdd
rlabel metal1 1504 722 1536 738 0 FILL_0__1025_.gnd
rlabel nsubstratencontact 1416 968 1416 968 0 FILL_0__1023_.vdd
rlabel metal1 1404 722 1436 738 0 FILL_0__1023_.gnd
rlabel metal1 1444 722 1516 738 0 _1023_.gnd
rlabel metal1 1444 962 1516 978 0 _1023_.vdd
rlabel metal2 1453 793 1467 807 0 _1023_.A
rlabel metal2 1473 833 1487 847 0 _1023_.Y
rlabel nsubstratencontact 1536 968 1536 968 0 FILL_1__1025_.vdd
rlabel metal1 1524 722 1556 738 0 FILL_1__1025_.gnd
rlabel nsubstratencontact 1644 968 1644 968 0 FILL_0__1004_.vdd
rlabel metal1 1624 722 1656 738 0 FILL_0__1004_.gnd
rlabel metal1 1544 722 1636 738 0 _1025_.gnd
rlabel metal1 1544 962 1636 978 0 _1025_.vdd
rlabel metal2 1553 853 1567 867 0 _1025_.A
rlabel metal2 1593 853 1607 867 0 _1025_.B
rlabel metal2 1573 833 1587 847 0 _1025_.Y
rlabel nsubstratencontact 1684 968 1684 968 0 FILL_2__1004_.vdd
rlabel metal1 1664 722 1696 738 0 FILL_2__1004_.gnd
rlabel nsubstratencontact 1664 968 1664 968 0 FILL_1__1004_.vdd
rlabel metal1 1644 722 1676 738 0 FILL_1__1004_.gnd
rlabel metal1 1684 722 1796 738 0 _1004_.gnd
rlabel metal1 1684 962 1796 978 0 _1004_.vdd
rlabel metal2 1773 833 1787 847 0 _1004_.A
rlabel metal2 1753 853 1767 867 0 _1004_.B
rlabel metal2 1733 833 1747 847 0 _1004_.C
rlabel metal2 1713 853 1727 867 0 _1004_.Y
rlabel nsubstratencontact 1824 968 1824 968 0 FILL_1__1000_.vdd
rlabel metal1 1804 722 1836 738 0 FILL_1__1000_.gnd
rlabel nsubstratencontact 1804 968 1804 968 0 FILL_0__1000_.vdd
rlabel metal1 1784 722 1816 738 0 FILL_0__1000_.gnd
rlabel metal1 1824 722 1936 738 0 _1000_.gnd
rlabel metal1 1824 962 1936 978 0 _1000_.vdd
rlabel metal2 1913 833 1927 847 0 _1000_.A
rlabel metal2 1893 853 1907 867 0 _1000_.B
rlabel metal2 1873 833 1887 847 0 _1000_.C
rlabel metal2 1853 853 1867 867 0 _1000_.Y
rlabel nsubstratencontact 1956 968 1956 968 0 FILL_1__1062_.vdd
rlabel metal1 1944 722 1976 738 0 FILL_1__1062_.gnd
rlabel nsubstratencontact 1936 968 1936 968 0 FILL_0__1062_.vdd
rlabel metal1 1924 722 1956 738 0 FILL_0__1062_.gnd
rlabel metal1 1964 722 2076 738 0 _1062_.gnd
rlabel metal1 1964 962 2076 978 0 _1062_.vdd
rlabel metal2 1973 833 1987 847 0 _1062_.A
rlabel metal2 1993 853 2007 867 0 _1062_.B
rlabel metal2 2013 833 2027 847 0 _1062_.C
rlabel metal2 2033 853 2047 867 0 _1062_.Y
rlabel nsubstratencontact 2096 968 2096 968 0 FILL_1__1228_.vdd
rlabel metal1 2084 722 2116 738 0 FILL_1__1228_.gnd
rlabel nsubstratencontact 2076 968 2076 968 0 FILL_0__1228_.vdd
rlabel metal1 2064 722 2096 738 0 FILL_0__1228_.gnd
rlabel metal1 2104 722 2216 738 0 _1228_.gnd
rlabel metal1 2104 962 2216 978 0 _1228_.vdd
rlabel metal2 2113 813 2127 827 0 _1228_.A
rlabel metal2 2133 833 2147 847 0 _1228_.B
rlabel metal2 2173 833 2187 847 0 _1228_.C
rlabel metal2 2153 813 2167 827 0 _1228_.Y
rlabel nsubstratencontact 2236 968 2236 968 0 FILL_1__1061_.vdd
rlabel metal1 2224 722 2256 738 0 FILL_1__1061_.gnd
rlabel nsubstratencontact 2216 968 2216 968 0 FILL_0__1061_.vdd
rlabel metal1 2204 722 2236 738 0 FILL_0__1061_.gnd
rlabel metal1 2244 722 2356 738 0 _1061_.gnd
rlabel metal1 2244 962 2356 978 0 _1061_.vdd
rlabel metal2 2253 813 2267 827 0 _1061_.A
rlabel metal2 2313 813 2327 827 0 _1061_.Y
rlabel metal2 2293 853 2307 867 0 _1061_.B
rlabel nsubstratencontact 2376 968 2376 968 0 FILL_1__1483_.vdd
rlabel metal1 2364 722 2396 738 0 FILL_1__1483_.gnd
rlabel nsubstratencontact 2356 968 2356 968 0 FILL_0__1483_.vdd
rlabel metal1 2344 722 2376 738 0 FILL_0__1483_.gnd
rlabel metal1 2384 722 2456 738 0 _1483_.gnd
rlabel metal1 2384 962 2456 978 0 _1483_.vdd
rlabel metal2 2393 793 2407 807 0 _1483_.A
rlabel metal2 2413 833 2427 847 0 _1483_.Y
rlabel nsubstratencontact 2484 968 2484 968 0 FILL_1__1882_.vdd
rlabel metal1 2464 722 2496 738 0 FILL_1__1882_.gnd
rlabel nsubstratencontact 2464 968 2464 968 0 FILL_0__1882_.vdd
rlabel metal1 2444 722 2476 738 0 FILL_0__1882_.gnd
rlabel metal1 2484 722 2576 738 0 _1882_.gnd
rlabel metal1 2484 962 2576 978 0 _1882_.vdd
rlabel metal2 2553 853 2567 867 0 _1882_.A
rlabel metal2 2513 853 2527 867 0 _1882_.B
rlabel metal2 2533 833 2547 847 0 _1882_.Y
rlabel nsubstratencontact 2604 968 2604 968 0 FILL_1__1881_.vdd
rlabel metal1 2584 722 2616 738 0 FILL_1__1881_.gnd
rlabel nsubstratencontact 2584 968 2584 968 0 FILL_0__1881_.vdd
rlabel metal1 2564 722 2596 738 0 FILL_0__1881_.gnd
rlabel metal1 2604 722 2716 738 0 _1881_.gnd
rlabel metal1 2604 962 2716 978 0 _1881_.vdd
rlabel metal2 2693 793 2707 807 0 _1881_.A
rlabel metal2 2673 813 2687 827 0 _1881_.B
rlabel metal2 2633 833 2647 847 0 _1881_.Y
rlabel nsubstratencontact 2736 968 2736 968 0 FILL_1__1880_.vdd
rlabel metal1 2724 722 2756 738 0 FILL_1__1880_.gnd
rlabel nsubstratencontact 2716 968 2716 968 0 FILL_0__1880_.vdd
rlabel metal1 2704 722 2736 738 0 FILL_0__1880_.gnd
rlabel metal1 2744 722 2836 738 0 _1880_.gnd
rlabel metal1 2744 962 2836 978 0 _1880_.vdd
rlabel metal2 2753 853 2767 867 0 _1880_.A
rlabel metal2 2793 853 2807 867 0 _1880_.B
rlabel metal2 2773 833 2787 847 0 _1880_.Y
rlabel nsubstratencontact 2864 968 2864 968 0 FILL_1__1858_.vdd
rlabel metal1 2844 722 2876 738 0 FILL_1__1858_.gnd
rlabel nsubstratencontact 2844 968 2844 968 0 FILL_0__1858_.vdd
rlabel metal1 2824 722 2856 738 0 FILL_0__1858_.gnd
rlabel metal1 2864 722 2956 738 0 _1858_.gnd
rlabel metal1 2864 962 2956 978 0 _1858_.vdd
rlabel metal2 2933 853 2947 867 0 _1858_.A
rlabel metal2 2893 853 2907 867 0 _1858_.B
rlabel metal2 2913 833 2927 847 0 _1858_.Y
rlabel nsubstratencontact 2996 968 2996 968 0 FILL_2__1833_.vdd
rlabel metal1 2984 722 3016 738 0 FILL_2__1833_.gnd
rlabel nsubstratencontact 2976 968 2976 968 0 FILL_1__1833_.vdd
rlabel metal1 2964 722 2996 738 0 FILL_1__1833_.gnd
rlabel nsubstratencontact 2956 968 2956 968 0 FILL_0__1833_.vdd
rlabel metal1 2944 722 2976 738 0 FILL_0__1833_.gnd
rlabel metal1 3004 722 3076 738 0 _1833_.gnd
rlabel metal1 3004 962 3076 978 0 _1833_.vdd
rlabel metal2 3013 793 3027 807 0 _1833_.A
rlabel metal2 3033 833 3047 847 0 _1833_.Y
rlabel nsubstratencontact 3104 968 3104 968 0 FILL_1__1777_.vdd
rlabel metal1 3084 722 3116 738 0 FILL_1__1777_.gnd
rlabel nsubstratencontact 3084 968 3084 968 0 FILL_0__1777_.vdd
rlabel metal1 3064 722 3096 738 0 FILL_0__1777_.gnd
rlabel metal1 3104 722 3176 738 0 _1777_.gnd
rlabel metal1 3104 962 3176 978 0 _1777_.vdd
rlabel metal2 3153 793 3167 807 0 _1777_.A
rlabel metal2 3133 833 3147 847 0 _1777_.Y
rlabel nsubstratencontact 3224 968 3224 968 0 FILL_2__1879_.vdd
rlabel metal1 3204 722 3236 738 0 FILL_2__1879_.gnd
rlabel nsubstratencontact 3204 968 3204 968 0 FILL_1__1879_.vdd
rlabel metal1 3184 722 3216 738 0 FILL_1__1879_.gnd
rlabel nsubstratencontact 3184 968 3184 968 0 FILL_0__1879_.vdd
rlabel metal1 3164 722 3196 738 0 FILL_0__1879_.gnd
rlabel metal1 3224 722 3316 738 0 _1879_.gnd
rlabel metal1 3224 962 3316 978 0 _1879_.vdd
rlabel metal2 3293 853 3307 867 0 _1879_.A
rlabel metal2 3253 853 3267 867 0 _1879_.B
rlabel metal2 3273 833 3287 847 0 _1879_.Y
rlabel nsubstratencontact 3364 968 3364 968 0 FILL_2__1800_.vdd
rlabel metal1 3344 722 3376 738 0 FILL_2__1800_.gnd
rlabel nsubstratencontact 3344 968 3344 968 0 FILL_1__1800_.vdd
rlabel metal1 3324 722 3356 738 0 FILL_1__1800_.gnd
rlabel nsubstratencontact 3324 968 3324 968 0 FILL_0__1800_.vdd
rlabel metal1 3304 722 3336 738 0 FILL_0__1800_.gnd
rlabel nsubstratencontact 3464 968 3464 968 0 FILL_0__1799_.vdd
rlabel metal1 3444 722 3476 738 0 FILL_0__1799_.gnd
rlabel metal1 3364 722 3456 738 0 _1800_.gnd
rlabel metal1 3364 962 3456 978 0 _1800_.vdd
rlabel metal2 3393 813 3407 827 0 _1800_.B
rlabel metal2 3433 813 3447 827 0 _1800_.A
rlabel metal2 3413 793 3427 807 0 _1800_.Y
rlabel nsubstratencontact 3484 968 3484 968 0 FILL_1__1799_.vdd
rlabel metal1 3464 722 3496 738 0 FILL_1__1799_.gnd
rlabel metal1 3484 722 3576 738 0 _1799_.gnd
rlabel metal1 3484 962 3576 978 0 _1799_.vdd
rlabel metal2 3513 813 3527 827 0 _1799_.B
rlabel metal2 3553 813 3567 827 0 _1799_.A
rlabel metal2 3533 793 3547 807 0 _1799_.Y
rlabel nsubstratencontact 3604 968 3604 968 0 FILL_1__1814_.vdd
rlabel metal1 3584 722 3616 738 0 FILL_1__1814_.gnd
rlabel nsubstratencontact 3584 968 3584 968 0 FILL_0__1814_.vdd
rlabel metal1 3564 722 3596 738 0 FILL_0__1814_.gnd
rlabel metal1 3604 722 3716 738 0 _1814_.gnd
rlabel metal1 3604 962 3716 978 0 _1814_.vdd
rlabel metal2 3693 833 3707 847 0 _1814_.A
rlabel metal2 3673 793 3687 807 0 _1814_.B
rlabel metal2 3653 833 3667 847 0 _1814_.C
rlabel metal2 3633 813 3647 827 0 _1814_.Y
rlabel nsubstratencontact 3744 968 3744 968 0 FILL_1__1798_.vdd
rlabel metal1 3724 722 3756 738 0 FILL_1__1798_.gnd
rlabel nsubstratencontact 3724 968 3724 968 0 FILL_0__1798_.vdd
rlabel metal1 3704 722 3736 738 0 FILL_0__1798_.gnd
rlabel metal1 3744 722 3816 738 0 _1798_.gnd
rlabel metal1 3744 962 3816 978 0 _1798_.vdd
rlabel metal2 3793 793 3807 807 0 _1798_.A
rlabel metal2 3773 833 3787 847 0 _1798_.Y
rlabel nsubstratencontact 3844 968 3844 968 0 FILL_1__1797_.vdd
rlabel metal1 3824 722 3856 738 0 FILL_1__1797_.gnd
rlabel nsubstratencontact 3824 968 3824 968 0 FILL_0__1797_.vdd
rlabel metal1 3804 722 3836 738 0 FILL_0__1797_.gnd
rlabel metal1 3844 722 3956 738 0 _1797_.gnd
rlabel metal1 3844 962 3956 978 0 _1797_.vdd
rlabel metal2 3933 813 3947 827 0 _1797_.A
rlabel metal2 3913 833 3927 847 0 _1797_.B
rlabel metal2 3873 833 3887 847 0 _1797_.C
rlabel metal2 3893 813 3907 827 0 _1797_.Y
rlabel nsubstratencontact 3976 968 3976 968 0 FILL_1__1796_.vdd
rlabel metal1 3964 722 3996 738 0 FILL_1__1796_.gnd
rlabel nsubstratencontact 3956 968 3956 968 0 FILL_0__1796_.vdd
rlabel metal1 3944 722 3976 738 0 FILL_0__1796_.gnd
rlabel metal1 3984 722 4076 738 0 _1796_.gnd
rlabel metal1 3984 962 4076 978 0 _1796_.vdd
rlabel metal2 3993 853 4007 867 0 _1796_.A
rlabel metal2 4033 853 4047 867 0 _1796_.B
rlabel metal2 4013 833 4027 847 0 _1796_.Y
rlabel nsubstratencontact 4104 968 4104 968 0 FILL_1__1771_.vdd
rlabel metal1 4084 722 4116 738 0 FILL_1__1771_.gnd
rlabel nsubstratencontact 4084 968 4084 968 0 FILL_0__1771_.vdd
rlabel metal1 4064 722 4096 738 0 FILL_0__1771_.gnd
rlabel metal1 4104 722 4216 738 0 _1771_.gnd
rlabel metal1 4104 962 4216 978 0 _1771_.vdd
rlabel metal2 4193 813 4207 827 0 _1771_.A
rlabel metal2 4173 833 4187 847 0 _1771_.B
rlabel metal2 4133 833 4147 847 0 _1771_.C
rlabel metal2 4153 813 4167 827 0 _1771_.Y
rlabel nsubstratencontact 4244 968 4244 968 0 FILL_1__1770_.vdd
rlabel metal1 4224 722 4256 738 0 FILL_1__1770_.gnd
rlabel nsubstratencontact 4224 968 4224 968 0 FILL_0__1770_.vdd
rlabel metal1 4204 722 4236 738 0 FILL_0__1770_.gnd
rlabel metal1 4244 722 4356 738 0 _1770_.gnd
rlabel metal1 4244 962 4356 978 0 _1770_.vdd
rlabel metal2 4333 813 4347 827 0 _1770_.A
rlabel metal2 4313 833 4327 847 0 _1770_.B
rlabel metal2 4273 833 4287 847 0 _1770_.C
rlabel metal2 4293 813 4307 827 0 _1770_.Y
rlabel nsubstratencontact 4396 968 4396 968 0 FILL_2__1781_.vdd
rlabel metal1 4384 722 4416 738 0 FILL_2__1781_.gnd
rlabel nsubstratencontact 4376 968 4376 968 0 FILL_1__1781_.vdd
rlabel metal1 4364 722 4396 738 0 FILL_1__1781_.gnd
rlabel nsubstratencontact 4356 968 4356 968 0 FILL_0__1781_.vdd
rlabel metal1 4344 722 4376 738 0 FILL_0__1781_.gnd
rlabel metal1 4404 722 4476 738 0 _1781_.gnd
rlabel metal1 4404 962 4476 978 0 _1781_.vdd
rlabel metal2 4413 793 4427 807 0 _1781_.A
rlabel metal2 4433 833 4447 847 0 _1781_.Y
rlabel nsubstratencontact 4504 968 4504 968 0 FILL_1__1749_.vdd
rlabel metal1 4484 722 4516 738 0 FILL_1__1749_.gnd
rlabel nsubstratencontact 4484 968 4484 968 0 FILL_0__1749_.vdd
rlabel metal1 4464 722 4496 738 0 FILL_0__1749_.gnd
rlabel metal1 4504 722 4616 738 0 _1749_.gnd
rlabel metal1 4504 962 4616 978 0 _1749_.vdd
rlabel metal2 4593 813 4607 827 0 _1749_.A
rlabel metal2 4573 833 4587 847 0 _1749_.B
rlabel metal2 4533 833 4547 847 0 _1749_.C
rlabel metal2 4553 813 4567 827 0 _1749_.Y
rlabel nsubstratencontact 4636 968 4636 968 0 FILL_1__1750_.vdd
rlabel metal1 4624 722 4656 738 0 FILL_1__1750_.gnd
rlabel nsubstratencontact 4616 968 4616 968 0 FILL_0__1750_.vdd
rlabel metal1 4604 722 4636 738 0 FILL_0__1750_.gnd
rlabel metal1 4644 722 4756 738 0 _1750_.gnd
rlabel metal1 4644 962 4756 978 0 _1750_.vdd
rlabel metal2 4653 833 4667 847 0 _1750_.A
rlabel metal2 4673 793 4687 807 0 _1750_.B
rlabel metal2 4693 833 4707 847 0 _1750_.C
rlabel metal2 4713 813 4727 827 0 _1750_.Y
rlabel nsubstratencontact 4784 968 4784 968 0 FILL_1_BUFX2_insert13.vdd
rlabel metal1 4764 722 4796 738 0 FILL_1_BUFX2_insert13.gnd
rlabel nsubstratencontact 4764 968 4764 968 0 FILL_0_BUFX2_insert13.vdd
rlabel metal1 4744 722 4776 738 0 FILL_0_BUFX2_insert13.gnd
rlabel metal1 4784 722 4876 738 0 BUFX2_insert13.gnd
rlabel metal1 4784 962 4876 978 0 BUFX2_insert13.vdd
rlabel metal2 4853 813 4867 827 0 BUFX2_insert13.A
rlabel metal2 4813 813 4827 827 0 BUFX2_insert13.Y
rlabel nsubstratencontact 4904 968 4904 968 0 FILL_1__1703_.vdd
rlabel metal1 4884 722 4916 738 0 FILL_1__1703_.gnd
rlabel nsubstratencontact 4884 968 4884 968 0 FILL_0__1703_.vdd
rlabel metal1 4864 722 4896 738 0 FILL_0__1703_.gnd
rlabel metal1 4904 722 5016 738 0 _1703_.gnd
rlabel metal1 4904 962 5016 978 0 _1703_.vdd
rlabel metal2 4993 813 5007 827 0 _1703_.A
rlabel metal2 4973 833 4987 847 0 _1703_.B
rlabel metal2 4933 833 4947 847 0 _1703_.C
rlabel metal2 4953 813 4967 827 0 _1703_.Y
rlabel nsubstratencontact 5036 968 5036 968 0 FILL_1__1704_.vdd
rlabel metal1 5024 722 5056 738 0 FILL_1__1704_.gnd
rlabel nsubstratencontact 5016 968 5016 968 0 FILL_0__1704_.vdd
rlabel metal1 5004 722 5036 738 0 FILL_0__1704_.gnd
rlabel metal1 5044 722 5156 738 0 _1704_.gnd
rlabel metal1 5044 962 5156 978 0 _1704_.vdd
rlabel metal2 5053 833 5067 847 0 _1704_.A
rlabel metal2 5073 793 5087 807 0 _1704_.B
rlabel metal2 5093 833 5107 847 0 _1704_.C
rlabel metal2 5113 813 5127 827 0 _1704_.Y
rlabel nsubstratencontact 5184 968 5184 968 0 FILL_1__1708_.vdd
rlabel metal1 5164 722 5196 738 0 FILL_1__1708_.gnd
rlabel nsubstratencontact 5164 968 5164 968 0 FILL_0__1708_.vdd
rlabel metal1 5144 722 5176 738 0 FILL_0__1708_.gnd
rlabel metal1 5184 722 5296 738 0 _1708_.gnd
rlabel metal1 5184 962 5296 978 0 _1708_.vdd
rlabel metal2 5273 793 5287 807 0 _1708_.A
rlabel metal2 5253 813 5267 827 0 _1708_.B
rlabel metal2 5213 833 5227 847 0 _1708_.Y
rlabel nsubstratencontact 5344 968 5344 968 0 FILL_2__1689_.vdd
rlabel metal1 5324 722 5356 738 0 FILL_2__1689_.gnd
rlabel nsubstratencontact 5324 968 5324 968 0 FILL_1__1689_.vdd
rlabel metal1 5304 722 5336 738 0 FILL_1__1689_.gnd
rlabel nsubstratencontact 5304 968 5304 968 0 FILL_0__1689_.vdd
rlabel metal1 5284 722 5316 738 0 FILL_0__1689_.gnd
rlabel metal1 5344 722 5416 738 0 _1689_.gnd
rlabel metal1 5344 962 5416 978 0 _1689_.vdd
rlabel metal2 5393 793 5407 807 0 _1689_.A
rlabel metal2 5373 833 5387 847 0 _1689_.Y
rlabel nsubstratencontact 5444 968 5444 968 0 FILL_1__1734_.vdd
rlabel metal1 5424 722 5456 738 0 FILL_1__1734_.gnd
rlabel nsubstratencontact 5424 968 5424 968 0 FILL_0__1734_.vdd
rlabel metal1 5404 722 5436 738 0 FILL_0__1734_.gnd
rlabel metal1 5444 722 5576 738 0 _1734_.gnd
rlabel metal1 5444 962 5576 978 0 _1734_.vdd
rlabel metal2 5553 813 5567 827 0 _1734_.A
rlabel metal2 5533 833 5547 847 0 _1734_.B
rlabel metal2 5473 813 5487 827 0 _1734_.C
rlabel metal2 5493 833 5507 847 0 _1734_.D
rlabel metal2 5513 813 5527 827 0 _1734_.Y
rlabel metal1 5624 722 5736 738 0 _1728_.gnd
rlabel metal1 5624 962 5736 978 0 _1728_.vdd
rlabel metal2 5633 813 5647 827 0 _1728_.A
rlabel metal2 5653 833 5667 847 0 _1728_.B
rlabel metal2 5693 833 5707 847 0 _1728_.C
rlabel metal2 5673 813 5687 827 0 _1728_.Y
rlabel nsubstratencontact 5736 968 5736 968 0 FILL85950x10950.vdd
rlabel metal1 5724 722 5756 738 0 FILL85950x10950.gnd
rlabel nsubstratencontact 5756 968 5756 968 0 FILL86250x10950.vdd
rlabel metal1 5744 722 5776 738 0 FILL86250x10950.gnd
rlabel nsubstratencontact 5776 968 5776 968 0 FILL86550x10950.vdd
rlabel metal1 5764 722 5796 738 0 FILL86550x10950.gnd
rlabel nsubstratencontact 5796 968 5796 968 0 FILL86850x10950.vdd
rlabel metal1 5784 722 5816 738 0 FILL86850x10950.gnd
rlabel nsubstratencontact 5576 968 5576 968 0 FILL_0__1728_.vdd
rlabel metal1 5564 722 5596 738 0 FILL_0__1728_.gnd
rlabel nsubstratencontact 5596 968 5596 968 0 FILL_1__1728_.vdd
rlabel metal1 5584 722 5616 738 0 FILL_1__1728_.gnd
rlabel nsubstratencontact 5616 968 5616 968 0 FILL_2__1728_.vdd
rlabel metal1 5604 722 5636 738 0 FILL_2__1728_.gnd
rlabel nsubstratencontact 136 972 136 972 0 FILL_1__1055_.vdd
rlabel metal1 124 1202 156 1218 0 FILL_1__1055_.gnd
rlabel nsubstratencontact 44 972 44 972 0 FILL_1__1046_.vdd
rlabel metal1 24 1202 56 1218 0 FILL_1__1046_.gnd
rlabel nsubstratencontact 116 972 116 972 0 FILL_0__1055_.vdd
rlabel metal1 104 1202 136 1218 0 FILL_0__1055_.gnd
rlabel nsubstratencontact 24 972 24 972 0 FILL_0__1046_.vdd
rlabel metal1 4 1202 36 1218 0 FILL_0__1046_.gnd
rlabel metal1 44 1202 116 1218 0 _1046_.gnd
rlabel metal1 44 962 116 978 0 _1046_.vdd
rlabel metal2 93 1133 107 1147 0 _1046_.A
rlabel metal2 73 1093 87 1107 0 _1046_.Y
rlabel nsubstratencontact 256 972 256 972 0 FILL_0__1047_.vdd
rlabel metal1 244 1202 276 1218 0 FILL_0__1047_.gnd
rlabel metal1 144 1202 256 1218 0 _1055_.gnd
rlabel metal1 144 962 256 978 0 _1055_.vdd
rlabel metal2 153 1093 167 1107 0 _1055_.A
rlabel metal2 173 1133 187 1147 0 _1055_.B
rlabel metal2 193 1093 207 1107 0 _1055_.C
rlabel metal2 213 1113 227 1127 0 _1055_.Y
rlabel nsubstratencontact 276 972 276 972 0 FILL_1__1047_.vdd
rlabel metal1 264 1202 296 1218 0 FILL_1__1047_.gnd
rlabel metal1 284 1202 396 1218 0 _1047_.gnd
rlabel metal1 284 962 396 978 0 _1047_.vdd
rlabel metal2 293 1113 307 1127 0 _1047_.A
rlabel metal2 313 1093 327 1107 0 _1047_.B
rlabel metal2 353 1093 367 1107 0 _1047_.C
rlabel metal2 333 1113 347 1127 0 _1047_.Y
rlabel nsubstratencontact 416 972 416 972 0 FILL_1__1118_.vdd
rlabel metal1 404 1202 436 1218 0 FILL_1__1118_.gnd
rlabel nsubstratencontact 396 972 396 972 0 FILL_0__1118_.vdd
rlabel metal1 384 1202 416 1218 0 FILL_0__1118_.gnd
rlabel metal1 424 1202 536 1218 0 _1118_.gnd
rlabel metal1 424 962 536 978 0 _1118_.vdd
rlabel metal2 433 1113 447 1127 0 _1118_.A
rlabel metal2 453 1093 467 1107 0 _1118_.B
rlabel metal2 493 1093 507 1107 0 _1118_.C
rlabel metal2 473 1113 487 1127 0 _1118_.Y
rlabel nsubstratencontact 564 972 564 972 0 FILL_1__1119_.vdd
rlabel metal1 544 1202 576 1218 0 FILL_1__1119_.gnd
rlabel nsubstratencontact 544 972 544 972 0 FILL_0__1119_.vdd
rlabel metal1 524 1202 556 1218 0 FILL_0__1119_.gnd
rlabel metal1 564 1202 676 1218 0 _1119_.gnd
rlabel metal1 564 962 676 978 0 _1119_.vdd
rlabel metal2 653 1093 667 1107 0 _1119_.A
rlabel metal2 633 1073 647 1087 0 _1119_.B
rlabel metal2 613 1093 627 1107 0 _1119_.C
rlabel metal2 593 1073 607 1087 0 _1119_.Y
rlabel nsubstratencontact 696 972 696 972 0 FILL_1__1112_.vdd
rlabel metal1 684 1202 716 1218 0 FILL_1__1112_.gnd
rlabel nsubstratencontact 676 972 676 972 0 FILL_0__1112_.vdd
rlabel metal1 664 1202 696 1218 0 FILL_0__1112_.gnd
rlabel metal1 704 1202 816 1218 0 _1112_.gnd
rlabel metal1 704 962 816 978 0 _1112_.vdd
rlabel metal2 713 1113 727 1127 0 _1112_.A
rlabel metal2 733 1093 747 1107 0 _1112_.B
rlabel metal2 773 1093 787 1107 0 _1112_.C
rlabel metal2 753 1113 767 1127 0 _1112_.Y
rlabel nsubstratencontact 856 972 856 972 0 FILL_2__1246_.vdd
rlabel metal1 844 1202 876 1218 0 FILL_2__1246_.gnd
rlabel nsubstratencontact 836 972 836 972 0 FILL_1__1246_.vdd
rlabel metal1 824 1202 856 1218 0 FILL_1__1246_.gnd
rlabel nsubstratencontact 816 972 816 972 0 FILL_0__1246_.vdd
rlabel metal1 804 1202 836 1218 0 FILL_0__1246_.gnd
rlabel metal1 864 1202 976 1218 0 _1246_.gnd
rlabel metal1 864 962 976 978 0 _1246_.vdd
rlabel metal2 873 1093 887 1107 0 _1246_.A
rlabel metal2 893 1133 907 1147 0 _1246_.B
rlabel metal2 913 1093 927 1107 0 _1246_.C
rlabel metal2 933 1113 947 1127 0 _1246_.Y
rlabel nsubstratencontact 1004 972 1004 972 0 FILL_1__1022_.vdd
rlabel metal1 984 1202 1016 1218 0 FILL_1__1022_.gnd
rlabel nsubstratencontact 984 972 984 972 0 FILL_0__1022_.vdd
rlabel metal1 964 1202 996 1218 0 FILL_0__1022_.gnd
rlabel metal1 1004 1202 1116 1218 0 _1022_.gnd
rlabel metal1 1004 962 1116 978 0 _1022_.vdd
rlabel metal2 1093 1113 1107 1127 0 _1022_.A
rlabel metal2 1073 1093 1087 1107 0 _1022_.B
rlabel metal2 1033 1093 1047 1107 0 _1022_.C
rlabel metal2 1053 1113 1067 1127 0 _1022_.Y
rlabel nsubstratencontact 1144 972 1144 972 0 FILL_1__1021_.vdd
rlabel metal1 1124 1202 1156 1218 0 FILL_1__1021_.gnd
rlabel nsubstratencontact 1124 972 1124 972 0 FILL_0__1021_.vdd
rlabel metal1 1104 1202 1136 1218 0 FILL_0__1021_.gnd
rlabel nsubstratencontact 1236 972 1236 972 0 FILL_1__1101_.vdd
rlabel metal1 1224 1202 1256 1218 0 FILL_1__1101_.gnd
rlabel nsubstratencontact 1216 972 1216 972 0 FILL_0__1101_.vdd
rlabel metal1 1204 1202 1236 1218 0 FILL_0__1101_.gnd
rlabel metal1 1244 1202 1356 1218 0 _1101_.gnd
rlabel metal1 1244 962 1356 978 0 _1101_.vdd
rlabel metal2 1253 1093 1267 1107 0 _1101_.A
rlabel metal2 1273 1133 1287 1147 0 _1101_.B
rlabel metal2 1293 1093 1307 1107 0 _1101_.C
rlabel metal2 1313 1113 1327 1127 0 _1101_.Y
rlabel metal1 1144 1202 1216 1218 0 _1021_.gnd
rlabel metal1 1144 962 1216 978 0 _1021_.vdd
rlabel metal2 1193 1133 1207 1147 0 _1021_.A
rlabel metal2 1173 1093 1187 1107 0 _1021_.Y
rlabel nsubstratencontact 1384 972 1384 972 0 FILL_1__1016_.vdd
rlabel metal1 1364 1202 1396 1218 0 FILL_1__1016_.gnd
rlabel nsubstratencontact 1364 972 1364 972 0 FILL_0__1016_.vdd
rlabel metal1 1344 1202 1376 1218 0 FILL_0__1016_.gnd
rlabel metal1 1384 1202 1456 1218 0 _1016_.gnd
rlabel metal1 1384 962 1456 978 0 _1016_.vdd
rlabel metal2 1433 1133 1447 1147 0 _1016_.A
rlabel metal2 1413 1093 1427 1107 0 _1016_.Y
rlabel nsubstratencontact 1484 972 1484 972 0 FILL_1__1019_.vdd
rlabel metal1 1464 1202 1496 1218 0 FILL_1__1019_.gnd
rlabel nsubstratencontact 1464 972 1464 972 0 FILL_0__1019_.vdd
rlabel metal1 1444 1202 1476 1218 0 FILL_0__1019_.gnd
rlabel metal1 1484 1202 1576 1218 0 _1019_.gnd
rlabel metal1 1484 962 1576 978 0 _1019_.vdd
rlabel metal2 1513 1113 1527 1127 0 _1019_.B
rlabel metal2 1553 1113 1567 1127 0 _1019_.A
rlabel metal2 1533 1133 1547 1147 0 _1019_.Y
rlabel nsubstratencontact 1616 972 1616 972 0 FILL_2__1024_.vdd
rlabel metal1 1604 1202 1636 1218 0 FILL_2__1024_.gnd
rlabel nsubstratencontact 1596 972 1596 972 0 FILL_1__1024_.vdd
rlabel metal1 1584 1202 1616 1218 0 FILL_1__1024_.gnd
rlabel nsubstratencontact 1576 972 1576 972 0 FILL_0__1024_.vdd
rlabel metal1 1564 1202 1596 1218 0 FILL_0__1024_.gnd
rlabel metal1 1624 1202 1696 1218 0 _1024_.gnd
rlabel metal1 1624 962 1696 978 0 _1024_.vdd
rlabel metal2 1633 1133 1647 1147 0 _1024_.A
rlabel metal2 1653 1093 1667 1107 0 _1024_.Y
rlabel nsubstratencontact 1724 972 1724 972 0 FILL_1__1015_.vdd
rlabel metal1 1704 1202 1736 1218 0 FILL_1__1015_.gnd
rlabel nsubstratencontact 1704 972 1704 972 0 FILL_0__1015_.vdd
rlabel metal1 1684 1202 1716 1218 0 FILL_0__1015_.gnd
rlabel metal1 1724 1202 1836 1218 0 _1015_.gnd
rlabel metal1 1724 962 1836 978 0 _1015_.vdd
rlabel metal2 1813 1093 1827 1107 0 _1015_.A
rlabel metal2 1793 1073 1807 1087 0 _1015_.B
rlabel metal2 1773 1093 1787 1107 0 _1015_.C
rlabel metal2 1753 1073 1767 1087 0 _1015_.Y
rlabel nsubstratencontact 1864 972 1864 972 0 FILL_1__1085_.vdd
rlabel metal1 1844 1202 1876 1218 0 FILL_1__1085_.gnd
rlabel nsubstratencontact 1844 972 1844 972 0 FILL_0__1085_.vdd
rlabel metal1 1824 1202 1856 1218 0 FILL_0__1085_.gnd
rlabel metal1 1864 1202 1956 1218 0 _1085_.gnd
rlabel metal1 1864 962 1956 978 0 _1085_.vdd
rlabel metal2 1933 1073 1947 1087 0 _1085_.A
rlabel metal2 1893 1073 1907 1087 0 _1085_.B
rlabel metal2 1913 1093 1927 1107 0 _1085_.Y
rlabel nsubstratencontact 1984 972 1984 972 0 FILL_1__1008_.vdd
rlabel metal1 1964 1202 1996 1218 0 FILL_1__1008_.gnd
rlabel nsubstratencontact 1964 972 1964 972 0 FILL_0__1008_.vdd
rlabel metal1 1944 1202 1976 1218 0 FILL_0__1008_.gnd
rlabel metal1 1984 1202 2096 1218 0 _1008_.gnd
rlabel metal1 1984 962 2096 978 0 _1008_.vdd
rlabel metal2 2073 1113 2087 1127 0 _1008_.A
rlabel metal2 2053 1093 2067 1107 0 _1008_.B
rlabel metal2 2013 1093 2027 1107 0 _1008_.C
rlabel metal2 2033 1113 2047 1127 0 _1008_.Y
rlabel nsubstratencontact 2124 972 2124 972 0 FILL_1__1001_.vdd
rlabel metal1 2104 1202 2136 1218 0 FILL_1__1001_.gnd
rlabel nsubstratencontact 2104 972 2104 972 0 FILL_0__1001_.vdd
rlabel metal1 2084 1202 2116 1218 0 FILL_0__1001_.gnd
rlabel metal1 2124 1202 2236 1218 0 _1001_.gnd
rlabel metal1 2124 962 2236 978 0 _1001_.vdd
rlabel metal2 2213 1093 2227 1107 0 _1001_.A
rlabel metal2 2193 1073 2207 1087 0 _1001_.B
rlabel metal2 2173 1093 2187 1107 0 _1001_.C
rlabel metal2 2153 1073 2167 1087 0 _1001_.Y
rlabel nsubstratencontact 2264 972 2264 972 0 FILL_1__1058_.vdd
rlabel metal1 2244 1202 2276 1218 0 FILL_1__1058_.gnd
rlabel nsubstratencontact 2244 972 2244 972 0 FILL_0__1058_.vdd
rlabel metal1 2224 1202 2256 1218 0 FILL_0__1058_.gnd
rlabel metal1 2264 1202 2376 1218 0 _1058_.gnd
rlabel metal1 2264 962 2376 978 0 _1058_.vdd
rlabel metal2 2353 1093 2367 1107 0 _1058_.A
rlabel metal2 2333 1073 2347 1087 0 _1058_.B
rlabel metal2 2313 1093 2327 1107 0 _1058_.C
rlabel metal2 2293 1073 2307 1087 0 _1058_.Y
rlabel nsubstratencontact 2404 972 2404 972 0 FILL_1__1067_.vdd
rlabel metal1 2384 1202 2416 1218 0 FILL_1__1067_.gnd
rlabel nsubstratencontact 2384 972 2384 972 0 FILL_0__1067_.vdd
rlabel metal1 2364 1202 2396 1218 0 FILL_0__1067_.gnd
rlabel nsubstratencontact 2524 972 2524 972 0 FILL_0__1059_.vdd
rlabel metal1 2504 1202 2536 1218 0 FILL_0__1059_.gnd
rlabel metal1 2404 1202 2516 1218 0 _1067_.gnd
rlabel metal1 2404 962 2516 978 0 _1067_.vdd
rlabel metal2 2493 1113 2507 1127 0 _1067_.A
rlabel metal2 2473 1093 2487 1107 0 _1067_.B
rlabel metal2 2433 1093 2447 1107 0 _1067_.C
rlabel metal2 2453 1113 2467 1127 0 _1067_.Y
rlabel nsubstratencontact 2544 972 2544 972 0 FILL_1__1059_.vdd
rlabel metal1 2524 1202 2556 1218 0 FILL_1__1059_.gnd
rlabel nsubstratencontact 2656 972 2656 972 0 FILL_0__1272_.vdd
rlabel metal1 2644 1202 2676 1218 0 FILL_0__1272_.gnd
rlabel metal1 2544 1202 2656 1218 0 _1059_.gnd
rlabel metal1 2544 962 2656 978 0 _1059_.vdd
rlabel metal2 2633 1093 2647 1107 0 _1059_.A
rlabel metal2 2613 1073 2627 1087 0 _1059_.B
rlabel metal2 2593 1093 2607 1107 0 _1059_.C
rlabel metal2 2573 1073 2587 1087 0 _1059_.Y
rlabel nsubstratencontact 2696 972 2696 972 0 FILL_2__1272_.vdd
rlabel metal1 2684 1202 2716 1218 0 FILL_2__1272_.gnd
rlabel nsubstratencontact 2676 972 2676 972 0 FILL_1__1272_.vdd
rlabel metal1 2664 1202 2696 1218 0 FILL_1__1272_.gnd
rlabel nsubstratencontact 2776 972 2776 972 0 FILL_0__1532_.vdd
rlabel metal1 2764 1202 2796 1218 0 FILL_0__1532_.gnd
rlabel metal1 2704 1202 2776 1218 0 _1272_.gnd
rlabel metal1 2704 962 2776 978 0 _1272_.vdd
rlabel metal2 2713 1133 2727 1147 0 _1272_.A
rlabel metal2 2733 1093 2747 1107 0 _1272_.Y
rlabel nsubstratencontact 2796 972 2796 972 0 FILL_1__1532_.vdd
rlabel metal1 2784 1202 2816 1218 0 FILL_1__1532_.gnd
rlabel nsubstratencontact 2896 972 2896 972 0 FILL_0__1855_.vdd
rlabel metal1 2884 1202 2916 1218 0 FILL_0__1855_.gnd
rlabel metal1 2804 1202 2896 1218 0 _1532_.gnd
rlabel metal1 2804 962 2896 978 0 _1532_.vdd
rlabel metal2 2853 1113 2867 1127 0 _1532_.B
rlabel metal2 2813 1113 2827 1127 0 _1532_.A
rlabel metal2 2833 1133 2847 1147 0 _1532_.Y
rlabel nsubstratencontact 3036 972 3036 972 0 FILL_1__1856_.vdd
rlabel metal1 3024 1202 3056 1218 0 FILL_1__1856_.gnd
rlabel nsubstratencontact 2916 972 2916 972 0 FILL_1__1855_.vdd
rlabel metal1 2904 1202 2936 1218 0 FILL_1__1855_.gnd
rlabel nsubstratencontact 3016 972 3016 972 0 FILL_0__1856_.vdd
rlabel metal1 3004 1202 3036 1218 0 FILL_0__1856_.gnd
rlabel metal1 2924 1202 3016 1218 0 _1855_.gnd
rlabel metal1 2924 962 3016 978 0 _1855_.vdd
rlabel metal2 2973 1113 2987 1127 0 _1855_.B
rlabel metal2 2933 1113 2947 1127 0 _1855_.A
rlabel metal2 2953 1133 2967 1147 0 _1855_.Y
rlabel nsubstratencontact 3164 972 3164 972 0 FILL_0__1271_.vdd
rlabel metal1 3144 1202 3176 1218 0 FILL_0__1271_.gnd
rlabel metal1 3044 1202 3156 1218 0 _1856_.gnd
rlabel metal1 3044 962 3156 978 0 _1856_.vdd
rlabel metal2 3053 1113 3067 1127 0 _1856_.A
rlabel metal2 3113 1113 3127 1127 0 _1856_.Y
rlabel metal2 3093 1073 3107 1087 0 _1856_.B
rlabel nsubstratencontact 3184 972 3184 972 0 FILL_1__1271_.vdd
rlabel metal1 3164 1202 3196 1218 0 FILL_1__1271_.gnd
rlabel nsubstratencontact 3284 972 3284 972 0 FILL_0__1852_.vdd
rlabel metal1 3264 1202 3296 1218 0 FILL_0__1852_.gnd
rlabel metal1 3184 1202 3276 1218 0 _1271_.gnd
rlabel metal1 3184 962 3276 978 0 _1271_.vdd
rlabel metal2 3213 1113 3227 1127 0 _1271_.B
rlabel metal2 3253 1113 3267 1127 0 _1271_.A
rlabel metal2 3233 1133 3247 1147 0 _1271_.Y
rlabel nsubstratencontact 3324 972 3324 972 0 FILL_2__1852_.vdd
rlabel metal1 3304 1202 3336 1218 0 FILL_2__1852_.gnd
rlabel nsubstratencontact 3304 972 3304 972 0 FILL_1__1852_.vdd
rlabel metal1 3284 1202 3316 1218 0 FILL_1__1852_.gnd
rlabel nsubstratencontact 3424 972 3424 972 0 FILL_0__1877_.vdd
rlabel metal1 3404 1202 3436 1218 0 FILL_0__1877_.gnd
rlabel metal1 3324 1202 3416 1218 0 _1852_.gnd
rlabel metal1 3324 962 3416 978 0 _1852_.vdd
rlabel metal2 3353 1113 3367 1127 0 _1852_.B
rlabel metal2 3393 1113 3407 1127 0 _1852_.A
rlabel metal2 3373 1133 3387 1147 0 _1852_.Y
rlabel nsubstratencontact 3444 972 3444 972 0 FILL_1__1877_.vdd
rlabel metal1 3424 1202 3456 1218 0 FILL_1__1877_.gnd
rlabel nsubstratencontact 3544 972 3544 972 0 FILL_1__1828_.vdd
rlabel metal1 3524 1202 3556 1218 0 FILL_1__1828_.gnd
rlabel nsubstratencontact 3524 972 3524 972 0 FILL_0__1828_.vdd
rlabel metal1 3504 1202 3536 1218 0 FILL_0__1828_.gnd
rlabel metal1 3444 1202 3516 1218 0 _1877_.gnd
rlabel metal1 3444 962 3516 978 0 _1877_.vdd
rlabel metal2 3493 1133 3507 1147 0 _1877_.A
rlabel metal2 3473 1093 3487 1107 0 _1877_.Y
rlabel nsubstratencontact 3664 972 3664 972 0 FILL_0__1827_.vdd
rlabel metal1 3644 1202 3676 1218 0 FILL_0__1827_.gnd
rlabel metal1 3544 1202 3656 1218 0 _1828_.gnd
rlabel metal1 3544 962 3656 978 0 _1828_.vdd
rlabel metal2 3633 1113 3647 1127 0 _1828_.A
rlabel metal2 3613 1093 3627 1107 0 _1828_.B
rlabel metal2 3573 1093 3587 1107 0 _1828_.C
rlabel metal2 3593 1113 3607 1127 0 _1828_.Y
rlabel nsubstratencontact 3684 972 3684 972 0 FILL_1__1827_.vdd
rlabel metal1 3664 1202 3696 1218 0 FILL_1__1827_.gnd
rlabel nsubstratencontact 3796 972 3796 972 0 FILL_0__1878_.vdd
rlabel metal1 3784 1202 3816 1218 0 FILL_0__1878_.gnd
rlabel metal1 3684 1202 3796 1218 0 _1827_.gnd
rlabel metal1 3684 962 3796 978 0 _1827_.vdd
rlabel metal2 3773 1113 3787 1127 0 _1827_.A
rlabel metal2 3753 1093 3767 1107 0 _1827_.B
rlabel metal2 3713 1093 3727 1107 0 _1827_.C
rlabel metal2 3733 1113 3747 1127 0 _1827_.Y
rlabel nsubstratencontact 3816 972 3816 972 0 FILL_1__1878_.vdd
rlabel metal1 3804 1202 3836 1218 0 FILL_1__1878_.gnd
rlabel nsubstratencontact 3916 972 3916 972 0 FILL_0__1851_.vdd
rlabel metal1 3904 1202 3936 1218 0 FILL_0__1851_.gnd
rlabel metal1 3824 1202 3916 1218 0 _1878_.gnd
rlabel metal1 3824 962 3916 978 0 _1878_.vdd
rlabel metal2 3833 1073 3847 1087 0 _1878_.A
rlabel metal2 3873 1073 3887 1087 0 _1878_.B
rlabel metal2 3853 1093 3867 1107 0 _1878_.Y
rlabel nsubstratencontact 3936 972 3936 972 0 FILL_1__1851_.vdd
rlabel metal1 3924 1202 3956 1218 0 FILL_1__1851_.gnd
rlabel nsubstratencontact 4036 972 4036 972 0 FILL_0__1850_.vdd
rlabel metal1 4024 1202 4056 1218 0 FILL_0__1850_.gnd
rlabel metal1 3944 1202 4036 1218 0 _1851_.gnd
rlabel metal1 3944 962 4036 978 0 _1851_.vdd
rlabel metal2 3953 1073 3967 1087 0 _1851_.A
rlabel metal2 3993 1073 4007 1087 0 _1851_.B
rlabel metal2 3973 1093 3987 1107 0 _1851_.Y
rlabel nsubstratencontact 4056 972 4056 972 0 FILL_1__1850_.vdd
rlabel metal1 4044 1202 4076 1218 0 FILL_1__1850_.gnd
rlabel nsubstratencontact 4176 972 4176 972 0 FILL_1__1801_.vdd
rlabel metal1 4164 1202 4196 1218 0 FILL_1__1801_.gnd
rlabel nsubstratencontact 4156 972 4156 972 0 FILL_0__1801_.vdd
rlabel metal1 4144 1202 4176 1218 0 FILL_0__1801_.gnd
rlabel metal1 4064 1202 4156 1218 0 _1850_.gnd
rlabel metal1 4064 962 4156 978 0 _1850_.vdd
rlabel metal2 4113 1113 4127 1127 0 _1850_.B
rlabel metal2 4073 1113 4087 1127 0 _1850_.A
rlabel metal2 4093 1133 4107 1147 0 _1850_.Y
rlabel nsubstratencontact 4284 972 4284 972 0 FILL_1__1769_.vdd
rlabel metal1 4264 1202 4296 1218 0 FILL_1__1769_.gnd
rlabel nsubstratencontact 4264 972 4264 972 0 FILL_0__1769_.vdd
rlabel metal1 4244 1202 4276 1218 0 FILL_0__1769_.gnd
rlabel metal1 4184 1202 4256 1218 0 _1801_.gnd
rlabel metal1 4184 962 4256 978 0 _1801_.vdd
rlabel metal2 4193 1133 4207 1147 0 _1801_.A
rlabel metal2 4213 1093 4227 1107 0 _1801_.Y
rlabel metal1 4284 1202 4396 1218 0 _1769_.gnd
rlabel metal1 4284 962 4396 978 0 _1769_.vdd
rlabel metal2 4373 1093 4387 1107 0 _1769_.A
rlabel metal2 4353 1133 4367 1147 0 _1769_.B
rlabel metal2 4333 1093 4347 1107 0 _1769_.C
rlabel metal2 4313 1113 4327 1127 0 _1769_.Y
rlabel nsubstratencontact 4424 972 4424 972 0 FILL_1__1768_.vdd
rlabel metal1 4404 1202 4436 1218 0 FILL_1__1768_.gnd
rlabel nsubstratencontact 4404 972 4404 972 0 FILL_0__1768_.vdd
rlabel metal1 4384 1202 4416 1218 0 FILL_0__1768_.gnd
rlabel nsubstratencontact 4444 972 4444 972 0 FILL_2__1768_.vdd
rlabel metal1 4424 1202 4456 1218 0 FILL_2__1768_.gnd
rlabel metal1 4444 1202 4556 1218 0 _1768_.gnd
rlabel metal1 4444 962 4556 978 0 _1768_.vdd
rlabel metal2 4533 1113 4547 1127 0 _1768_.A
rlabel metal2 4513 1093 4527 1107 0 _1768_.B
rlabel metal2 4473 1093 4487 1107 0 _1768_.C
rlabel metal2 4493 1113 4507 1127 0 _1768_.Y
rlabel nsubstratencontact 4564 972 4564 972 0 FILL_0__1809_.vdd
rlabel metal1 4544 1202 4576 1218 0 FILL_0__1809_.gnd
rlabel nsubstratencontact 4584 972 4584 972 0 FILL_1__1809_.vdd
rlabel metal1 4564 1202 4596 1218 0 FILL_1__1809_.gnd
rlabel metal1 4584 1202 4696 1218 0 _1809_.gnd
rlabel metal1 4584 962 4696 978 0 _1809_.vdd
rlabel metal2 4673 1093 4687 1107 0 _1809_.A
rlabel metal2 4653 1133 4667 1147 0 _1809_.B
rlabel metal2 4633 1093 4647 1107 0 _1809_.C
rlabel metal2 4613 1113 4627 1127 0 _1809_.Y
rlabel nsubstratencontact 4716 972 4716 972 0 FILL_1__1808_.vdd
rlabel metal1 4704 1202 4736 1218 0 FILL_1__1808_.gnd
rlabel nsubstratencontact 4696 972 4696 972 0 FILL_0__1808_.vdd
rlabel metal1 4684 1202 4716 1218 0 FILL_0__1808_.gnd
rlabel metal1 4724 1202 4836 1218 0 _1808_.gnd
rlabel metal1 4724 962 4836 978 0 _1808_.vdd
rlabel metal2 4733 1113 4747 1127 0 _1808_.A
rlabel metal2 4753 1093 4767 1107 0 _1808_.B
rlabel metal2 4793 1093 4807 1107 0 _1808_.C
rlabel metal2 4773 1113 4787 1127 0 _1808_.Y
rlabel nsubstratencontact 4856 972 4856 972 0 FILL_1_BUFX2_insert11.vdd
rlabel metal1 4844 1202 4876 1218 0 FILL_1_BUFX2_insert11.gnd
rlabel nsubstratencontact 4836 972 4836 972 0 FILL_0_BUFX2_insert11.vdd
rlabel metal1 4824 1202 4856 1218 0 FILL_0_BUFX2_insert11.gnd
rlabel metal1 4864 1202 4956 1218 0 BUFX2_insert11.gnd
rlabel metal1 4864 962 4956 978 0 BUFX2_insert11.vdd
rlabel metal2 4873 1113 4887 1127 0 BUFX2_insert11.A
rlabel metal2 4913 1113 4927 1127 0 BUFX2_insert11.Y
rlabel nsubstratencontact 4976 972 4976 972 0 FILL_1__1711_.vdd
rlabel metal1 4964 1202 4996 1218 0 FILL_1__1711_.gnd
rlabel nsubstratencontact 4956 972 4956 972 0 FILL_0__1711_.vdd
rlabel metal1 4944 1202 4976 1218 0 FILL_0__1711_.gnd
rlabel nsubstratencontact 5056 972 5056 972 0 FILL_0__1685_.vdd
rlabel metal1 5044 1202 5076 1218 0 FILL_0__1685_.gnd
rlabel metal1 4984 1202 5056 1218 0 _1711_.gnd
rlabel metal1 4984 962 5056 978 0 _1711_.vdd
rlabel metal2 4993 1133 5007 1147 0 _1711_.A
rlabel metal2 5013 1093 5027 1107 0 _1711_.Y
rlabel nsubstratencontact 5184 972 5184 972 0 FILL_1__1710_.vdd
rlabel metal1 5164 1202 5196 1218 0 FILL_1__1710_.gnd
rlabel nsubstratencontact 5076 972 5076 972 0 FILL_1__1685_.vdd
rlabel metal1 5064 1202 5096 1218 0 FILL_1__1685_.gnd
rlabel nsubstratencontact 5164 972 5164 972 0 FILL_0__1710_.vdd
rlabel metal1 5144 1202 5176 1218 0 FILL_0__1710_.gnd
rlabel metal1 5084 1202 5156 1218 0 _1685_.gnd
rlabel metal1 5084 962 5156 978 0 _1685_.vdd
rlabel metal2 5093 1133 5107 1147 0 _1685_.A
rlabel metal2 5113 1093 5127 1107 0 _1685_.Y
rlabel nsubstratencontact 5304 972 5304 972 0 FILL_1__1709_.vdd
rlabel metal1 5284 1202 5316 1218 0 FILL_1__1709_.gnd
rlabel nsubstratencontact 5284 972 5284 972 0 FILL_0__1709_.vdd
rlabel metal1 5264 1202 5296 1218 0 FILL_0__1709_.gnd
rlabel metal1 5184 1202 5276 1218 0 _1710_.gnd
rlabel metal1 5184 962 5276 978 0 _1710_.vdd
rlabel metal2 5253 1073 5267 1087 0 _1710_.A
rlabel metal2 5213 1073 5227 1087 0 _1710_.B
rlabel metal2 5233 1093 5247 1107 0 _1710_.Y
rlabel nsubstratencontact 5324 972 5324 972 0 FILL_2__1709_.vdd
rlabel metal1 5304 1202 5336 1218 0 FILL_2__1709_.gnd
rlabel nsubstratencontact 5436 972 5436 972 0 FILL_0__1688_.vdd
rlabel metal1 5424 1202 5456 1218 0 FILL_0__1688_.gnd
rlabel metal1 5324 1202 5436 1218 0 _1709_.gnd
rlabel metal1 5324 962 5436 978 0 _1709_.vdd
rlabel metal2 5413 1113 5427 1127 0 _1709_.A
rlabel metal2 5393 1093 5407 1107 0 _1709_.B
rlabel metal2 5353 1093 5367 1107 0 _1709_.C
rlabel metal2 5373 1113 5387 1127 0 _1709_.Y
rlabel nsubstratencontact 5456 972 5456 972 0 FILL_1__1688_.vdd
rlabel metal1 5444 1202 5476 1218 0 FILL_1__1688_.gnd
rlabel nsubstratencontact 5564 972 5564 972 0 FILL_0__1733_.vdd
rlabel metal1 5544 1202 5576 1218 0 FILL_0__1733_.gnd
rlabel metal1 5464 1202 5556 1218 0 _1688_.gnd
rlabel metal1 5464 962 5556 978 0 _1688_.vdd
rlabel metal2 5513 1113 5527 1127 0 _1688_.B
rlabel metal2 5473 1113 5487 1127 0 _1688_.A
rlabel metal2 5493 1133 5507 1147 0 _1688_.Y
rlabel metal1 5724 1202 5796 1218 0 _1597_.gnd
rlabel metal1 5724 962 5796 978 0 _1597_.vdd
rlabel metal2 5773 1133 5787 1147 0 _1597_.A
rlabel metal2 5753 1093 5767 1107 0 _1597_.Y
rlabel metal1 5584 1202 5696 1218 0 _1733_.gnd
rlabel metal1 5584 962 5696 978 0 _1733_.vdd
rlabel metal2 5673 1093 5687 1107 0 _1733_.A
rlabel metal2 5653 1073 5667 1087 0 _1733_.B
rlabel metal2 5633 1093 5647 1107 0 _1733_.C
rlabel metal2 5613 1073 5627 1087 0 _1733_.Y
rlabel nsubstratencontact 5804 972 5804 972 0 FILL86850x14550.vdd
rlabel metal1 5784 1202 5816 1218 0 FILL86850x14550.gnd
rlabel nsubstratencontact 5704 972 5704 972 0 FILL_0__1597_.vdd
rlabel metal1 5684 1202 5716 1218 0 FILL_0__1597_.gnd
rlabel nsubstratencontact 5724 972 5724 972 0 FILL_1__1597_.vdd
rlabel metal1 5704 1202 5736 1218 0 FILL_1__1597_.gnd
rlabel nsubstratencontact 5584 972 5584 972 0 FILL_1__1733_.vdd
rlabel metal1 5564 1202 5596 1218 0 FILL_1__1733_.gnd
rlabel nsubstratencontact 44 1448 44 1448 0 FILL_1__1121_.vdd
rlabel metal1 24 1202 56 1218 0 FILL_1__1121_.gnd
rlabel nsubstratencontact 24 1448 24 1448 0 FILL_0__1121_.vdd
rlabel metal1 4 1202 36 1218 0 FILL_0__1121_.gnd
rlabel metal1 44 1202 156 1218 0 _1121_.gnd
rlabel metal1 44 1442 156 1458 0 _1121_.vdd
rlabel metal2 133 1313 147 1327 0 _1121_.A
rlabel metal2 113 1333 127 1347 0 _1121_.B
rlabel metal2 93 1313 107 1327 0 _1121_.C
rlabel metal2 73 1333 87 1347 0 _1121_.Y
rlabel nsubstratencontact 176 1448 176 1448 0 FILL_1__1123_.vdd
rlabel metal1 164 1202 196 1218 0 FILL_1__1123_.gnd
rlabel nsubstratencontact 156 1448 156 1448 0 FILL_0__1123_.vdd
rlabel metal1 144 1202 176 1218 0 FILL_0__1123_.gnd
rlabel metal1 184 1202 296 1218 0 _1123_.gnd
rlabel metal1 184 1442 296 1458 0 _1123_.vdd
rlabel metal2 193 1313 207 1327 0 _1123_.A
rlabel metal2 213 1273 227 1287 0 _1123_.B
rlabel metal2 233 1313 247 1327 0 _1123_.C
rlabel metal2 253 1293 267 1307 0 _1123_.Y
rlabel nsubstratencontact 324 1448 324 1448 0 FILL_1__1116_.vdd
rlabel metal1 304 1202 336 1218 0 FILL_1__1116_.gnd
rlabel nsubstratencontact 304 1448 304 1448 0 FILL_0__1116_.vdd
rlabel metal1 284 1202 316 1218 0 FILL_0__1116_.gnd
rlabel metal1 324 1202 436 1218 0 _1116_.gnd
rlabel metal1 324 1442 436 1458 0 _1116_.vdd
rlabel metal2 413 1313 427 1327 0 _1116_.A
rlabel metal2 393 1333 407 1347 0 _1116_.B
rlabel metal2 373 1313 387 1327 0 _1116_.C
rlabel metal2 353 1333 367 1347 0 _1116_.Y
rlabel nsubstratencontact 464 1448 464 1448 0 FILL_1__1195_.vdd
rlabel metal1 444 1202 476 1218 0 FILL_1__1195_.gnd
rlabel nsubstratencontact 444 1448 444 1448 0 FILL_0__1195_.vdd
rlabel metal1 424 1202 456 1218 0 FILL_0__1195_.gnd
rlabel metal1 464 1202 576 1218 0 _1195_.gnd
rlabel metal1 464 1442 576 1458 0 _1195_.vdd
rlabel metal2 553 1293 567 1307 0 _1195_.A
rlabel metal2 533 1313 547 1327 0 _1195_.B
rlabel metal2 493 1313 507 1327 0 _1195_.C
rlabel metal2 513 1293 527 1307 0 _1195_.Y
rlabel nsubstratencontact 604 1448 604 1448 0 FILL_1__1120_.vdd
rlabel metal1 584 1202 616 1218 0 FILL_1__1120_.gnd
rlabel nsubstratencontact 584 1448 584 1448 0 FILL_0__1120_.vdd
rlabel metal1 564 1202 596 1218 0 FILL_0__1120_.gnd
rlabel metal1 604 1202 716 1218 0 _1120_.gnd
rlabel metal1 604 1442 716 1458 0 _1120_.vdd
rlabel metal2 693 1293 707 1307 0 _1120_.A
rlabel metal2 673 1313 687 1327 0 _1120_.B
rlabel metal2 633 1313 647 1327 0 _1120_.C
rlabel metal2 653 1293 667 1307 0 _1120_.Y
rlabel nsubstratencontact 764 1448 764 1448 0 FILL_2__1115_.vdd
rlabel metal1 744 1202 776 1218 0 FILL_2__1115_.gnd
rlabel nsubstratencontact 744 1448 744 1448 0 FILL_1__1115_.vdd
rlabel metal1 724 1202 756 1218 0 FILL_1__1115_.gnd
rlabel nsubstratencontact 724 1448 724 1448 0 FILL_0__1115_.vdd
rlabel metal1 704 1202 736 1218 0 FILL_0__1115_.gnd
rlabel nsubstratencontact 876 1448 876 1448 0 FILL_0__1111_.vdd
rlabel metal1 864 1202 896 1218 0 FILL_0__1111_.gnd
rlabel metal1 764 1202 876 1218 0 _1115_.gnd
rlabel metal1 764 1442 876 1458 0 _1115_.vdd
rlabel metal2 853 1293 867 1307 0 _1115_.A
rlabel metal2 793 1293 807 1307 0 _1115_.Y
rlabel metal2 813 1333 827 1347 0 _1115_.B
rlabel nsubstratencontact 896 1448 896 1448 0 FILL_1__1111_.vdd
rlabel metal1 884 1202 916 1218 0 FILL_1__1111_.gnd
rlabel nsubstratencontact 1024 1448 1024 1448 0 FILL_1__1100_.vdd
rlabel metal1 1004 1202 1036 1218 0 FILL_1__1100_.gnd
rlabel nsubstratencontact 1004 1448 1004 1448 0 FILL_0__1100_.vdd
rlabel metal1 984 1202 1016 1218 0 FILL_0__1100_.gnd
rlabel metal1 904 1202 996 1218 0 _1111_.gnd
rlabel metal1 904 1442 996 1458 0 _1111_.vdd
rlabel metal2 913 1333 927 1347 0 _1111_.A
rlabel metal2 953 1333 967 1347 0 _1111_.B
rlabel metal2 933 1313 947 1327 0 _1111_.Y
rlabel nsubstratencontact 1116 1448 1116 1448 0 FILL_1__1107_.vdd
rlabel metal1 1104 1202 1136 1218 0 FILL_1__1107_.gnd
rlabel nsubstratencontact 1096 1448 1096 1448 0 FILL_0__1107_.vdd
rlabel metal1 1084 1202 1116 1218 0 FILL_0__1107_.gnd
rlabel metal1 1124 1202 1236 1218 0 _1107_.gnd
rlabel metal1 1124 1442 1236 1458 0 _1107_.vdd
rlabel metal2 1133 1313 1147 1327 0 _1107_.A
rlabel metal2 1153 1333 1167 1347 0 _1107_.B
rlabel metal2 1173 1313 1187 1327 0 _1107_.C
rlabel metal2 1193 1333 1207 1347 0 _1107_.Y
rlabel metal1 1024 1202 1096 1218 0 _1100_.gnd
rlabel metal1 1024 1442 1096 1458 0 _1100_.vdd
rlabel metal2 1073 1273 1087 1287 0 _1100_.A
rlabel metal2 1053 1313 1067 1327 0 _1100_.Y
rlabel nsubstratencontact 1256 1448 1256 1448 0 FILL_1__1106_.vdd
rlabel metal1 1244 1202 1276 1218 0 FILL_1__1106_.gnd
rlabel nsubstratencontact 1236 1448 1236 1448 0 FILL_0__1106_.vdd
rlabel metal1 1224 1202 1256 1218 0 FILL_0__1106_.gnd
rlabel nsubstratencontact 1384 1448 1384 1448 0 FILL_1__1092_.vdd
rlabel metal1 1364 1202 1396 1218 0 FILL_1__1092_.gnd
rlabel nsubstratencontact 1364 1448 1364 1448 0 FILL_0__1092_.vdd
rlabel metal1 1344 1202 1376 1218 0 FILL_0__1092_.gnd
rlabel metal1 1264 1202 1356 1218 0 _1106_.gnd
rlabel metal1 1264 1442 1356 1458 0 _1106_.vdd
rlabel metal2 1273 1333 1287 1347 0 _1106_.A
rlabel metal2 1313 1333 1327 1347 0 _1106_.B
rlabel metal2 1293 1313 1307 1327 0 _1106_.Y
rlabel metal1 1384 1202 1476 1218 0 _1092_.gnd
rlabel metal1 1384 1442 1476 1458 0 _1092_.vdd
rlabel metal2 1453 1333 1467 1347 0 _1092_.A
rlabel metal2 1413 1333 1427 1347 0 _1092_.B
rlabel metal2 1433 1313 1447 1327 0 _1092_.Y
rlabel nsubstratencontact 1504 1448 1504 1448 0 FILL_1__1083_.vdd
rlabel metal1 1484 1202 1516 1218 0 FILL_1__1083_.gnd
rlabel nsubstratencontact 1484 1448 1484 1448 0 FILL_0__1083_.vdd
rlabel metal1 1464 1202 1496 1218 0 FILL_0__1083_.gnd
rlabel metal1 1504 1202 1596 1218 0 _1083_.gnd
rlabel metal1 1504 1442 1596 1458 0 _1083_.vdd
rlabel metal2 1573 1333 1587 1347 0 _1083_.A
rlabel metal2 1533 1333 1547 1347 0 _1083_.B
rlabel metal2 1553 1313 1567 1327 0 _1083_.Y
rlabel nsubstratencontact 1644 1448 1644 1448 0 FILL_2__1089_.vdd
rlabel metal1 1624 1202 1656 1218 0 FILL_2__1089_.gnd
rlabel nsubstratencontact 1624 1448 1624 1448 0 FILL_1__1089_.vdd
rlabel metal1 1604 1202 1636 1218 0 FILL_1__1089_.gnd
rlabel nsubstratencontact 1604 1448 1604 1448 0 FILL_0__1089_.vdd
rlabel metal1 1584 1202 1616 1218 0 FILL_0__1089_.gnd
rlabel nsubstratencontact 1776 1448 1776 1448 0 FILL_1__1081_.vdd
rlabel metal1 1764 1202 1796 1218 0 FILL_1__1081_.gnd
rlabel nsubstratencontact 1756 1448 1756 1448 0 FILL_0__1081_.vdd
rlabel metal1 1744 1202 1776 1218 0 FILL_0__1081_.gnd
rlabel metal1 1644 1202 1756 1218 0 _1089_.gnd
rlabel metal1 1644 1442 1756 1458 0 _1089_.vdd
rlabel metal2 1733 1313 1747 1327 0 _1089_.A
rlabel metal2 1713 1333 1727 1347 0 _1089_.B
rlabel metal2 1693 1313 1707 1327 0 _1089_.C
rlabel metal2 1673 1333 1687 1347 0 _1089_.Y
rlabel nsubstratencontact 1904 1448 1904 1448 0 FILL_1__1084_.vdd
rlabel metal1 1884 1202 1916 1218 0 FILL_1__1084_.gnd
rlabel nsubstratencontact 1884 1448 1884 1448 0 FILL_0__1084_.vdd
rlabel metal1 1864 1202 1896 1218 0 FILL_0__1084_.gnd
rlabel metal1 1784 1202 1876 1218 0 _1081_.gnd
rlabel metal1 1784 1442 1876 1458 0 _1081_.vdd
rlabel metal2 1793 1333 1807 1347 0 _1081_.A
rlabel metal2 1833 1333 1847 1347 0 _1081_.B
rlabel metal2 1813 1313 1827 1327 0 _1081_.Y
rlabel nsubstratencontact 2024 1448 2024 1448 0 FILL_0__1075_.vdd
rlabel metal1 2004 1202 2036 1218 0 FILL_0__1075_.gnd
rlabel metal1 1904 1202 2016 1218 0 _1084_.gnd
rlabel metal1 1904 1442 2016 1458 0 _1084_.vdd
rlabel metal2 1993 1313 2007 1327 0 _1084_.A
rlabel metal2 1973 1333 1987 1347 0 _1084_.B
rlabel metal2 1953 1313 1967 1327 0 _1084_.C
rlabel metal2 1933 1333 1947 1347 0 _1084_.Y
rlabel nsubstratencontact 2164 1448 2164 1448 0 FILL_2__1017_.vdd
rlabel metal1 2144 1202 2176 1218 0 FILL_2__1017_.gnd
rlabel nsubstratencontact 2044 1448 2044 1448 0 FILL_1__1075_.vdd
rlabel metal1 2024 1202 2056 1218 0 FILL_1__1075_.gnd
rlabel nsubstratencontact 2144 1448 2144 1448 0 FILL_1__1017_.vdd
rlabel metal1 2124 1202 2156 1218 0 FILL_1__1017_.gnd
rlabel nsubstratencontact 2124 1448 2124 1448 0 FILL_0__1017_.vdd
rlabel metal1 2104 1202 2136 1218 0 FILL_0__1017_.gnd
rlabel metal1 2044 1202 2116 1218 0 _1075_.gnd
rlabel metal1 2044 1442 2116 1458 0 _1075_.vdd
rlabel metal2 2093 1273 2107 1287 0 _1075_.A
rlabel metal2 2073 1313 2087 1327 0 _1075_.Y
rlabel nsubstratencontact 2284 1448 2284 1448 0 FILL_0__1074_.vdd
rlabel metal1 2264 1202 2296 1218 0 FILL_0__1074_.gnd
rlabel metal1 2164 1202 2276 1218 0 _1017_.gnd
rlabel metal1 2164 1442 2276 1458 0 _1017_.vdd
rlabel metal2 2253 1313 2267 1327 0 _1017_.A
rlabel metal2 2233 1333 2247 1347 0 _1017_.B
rlabel metal2 2213 1313 2227 1327 0 _1017_.C
rlabel metal2 2193 1333 2207 1347 0 _1017_.Y
rlabel nsubstratencontact 2304 1448 2304 1448 0 FILL_1__1074_.vdd
rlabel metal1 2284 1202 2316 1218 0 FILL_1__1074_.gnd
rlabel metal1 2304 1202 2416 1218 0 _1074_.gnd
rlabel metal1 2304 1442 2416 1458 0 _1074_.vdd
rlabel metal2 2393 1313 2407 1327 0 _1074_.A
rlabel metal2 2373 1333 2387 1347 0 _1074_.B
rlabel metal2 2353 1313 2367 1327 0 _1074_.C
rlabel metal2 2333 1333 2347 1347 0 _1074_.Y
rlabel nsubstratencontact 2436 1448 2436 1448 0 FILL_1__944_.vdd
rlabel metal1 2424 1202 2456 1218 0 FILL_1__944_.gnd
rlabel nsubstratencontact 2524 1448 2524 1448 0 FILL_0__1533_.vdd
rlabel metal1 2504 1202 2536 1218 0 FILL_0__1533_.gnd
rlabel nsubstratencontact 2416 1448 2416 1448 0 FILL_0__944_.vdd
rlabel metal1 2404 1202 2436 1218 0 FILL_0__944_.gnd
rlabel metal1 2444 1202 2516 1218 0 _944_.gnd
rlabel metal1 2444 1442 2516 1458 0 _944_.vdd
rlabel metal2 2453 1273 2467 1287 0 _944_.A
rlabel metal2 2473 1313 2487 1327 0 _944_.Y
rlabel nsubstratencontact 2544 1448 2544 1448 0 FILL_1__1533_.vdd
rlabel metal1 2524 1202 2556 1218 0 FILL_1__1533_.gnd
rlabel nsubstratencontact 2564 1448 2564 1448 0 FILL_2__1533_.vdd
rlabel metal1 2544 1202 2576 1218 0 FILL_2__1533_.gnd
rlabel metal1 2564 1202 2676 1218 0 _1533_.gnd
rlabel metal1 2564 1442 2676 1458 0 _1533_.vdd
rlabel metal2 2653 1293 2667 1307 0 _1533_.A
rlabel metal2 2633 1313 2647 1327 0 _1533_.B
rlabel metal2 2593 1313 2607 1327 0 _1533_.C
rlabel metal2 2613 1293 2627 1307 0 _1533_.Y
rlabel nsubstratencontact 2696 1448 2696 1448 0 FILL_1__1485_.vdd
rlabel metal1 2684 1202 2716 1218 0 FILL_1__1485_.gnd
rlabel nsubstratencontact 2676 1448 2676 1448 0 FILL_0__1485_.vdd
rlabel metal1 2664 1202 2696 1218 0 FILL_0__1485_.gnd
rlabel metal1 2704 1202 2816 1218 0 _1485_.gnd
rlabel metal1 2704 1442 2816 1458 0 _1485_.vdd
rlabel metal2 2713 1313 2727 1327 0 _1485_.A
rlabel metal2 2733 1273 2747 1287 0 _1485_.B
rlabel metal2 2753 1313 2767 1327 0 _1485_.C
rlabel metal2 2773 1293 2787 1307 0 _1485_.Y
rlabel nsubstratencontact 2844 1448 2844 1448 0 FILL_1__1274_.vdd
rlabel metal1 2824 1202 2856 1218 0 FILL_1__1274_.gnd
rlabel nsubstratencontact 2824 1448 2824 1448 0 FILL_0__1274_.vdd
rlabel metal1 2804 1202 2836 1218 0 FILL_0__1274_.gnd
rlabel metal1 2844 1202 2956 1218 0 _1274_.gnd
rlabel metal1 2844 1442 2956 1458 0 _1274_.vdd
rlabel metal2 2933 1293 2947 1307 0 _1274_.A
rlabel metal2 2913 1313 2927 1327 0 _1274_.B
rlabel metal2 2873 1313 2887 1327 0 _1274_.C
rlabel metal2 2893 1293 2907 1307 0 _1274_.Y
rlabel nsubstratencontact 2984 1448 2984 1448 0 FILL_1__1431_.vdd
rlabel metal1 2964 1202 2996 1218 0 FILL_1__1431_.gnd
rlabel nsubstratencontact 2964 1448 2964 1448 0 FILL_0__1431_.vdd
rlabel metal1 2944 1202 2976 1218 0 FILL_0__1431_.gnd
rlabel metal1 2984 1202 3096 1218 0 _1431_.gnd
rlabel metal1 2984 1442 3096 1458 0 _1431_.vdd
rlabel metal2 3073 1293 3087 1307 0 _1431_.A
rlabel metal2 3053 1313 3067 1327 0 _1431_.B
rlabel metal2 3013 1313 3027 1327 0 _1431_.C
rlabel metal2 3033 1293 3047 1307 0 _1431_.Y
rlabel nsubstratencontact 3124 1448 3124 1448 0 FILL_1__1484_.vdd
rlabel metal1 3104 1202 3136 1218 0 FILL_1__1484_.gnd
rlabel nsubstratencontact 3104 1448 3104 1448 0 FILL_0__1484_.vdd
rlabel metal1 3084 1202 3116 1218 0 FILL_0__1484_.gnd
rlabel metal1 3124 1202 3236 1218 0 _1484_.gnd
rlabel metal1 3124 1442 3236 1458 0 _1484_.vdd
rlabel metal2 3213 1293 3227 1307 0 _1484_.A
rlabel metal2 3193 1313 3207 1327 0 _1484_.B
rlabel metal2 3153 1313 3167 1327 0 _1484_.C
rlabel metal2 3173 1293 3187 1307 0 _1484_.Y
rlabel nsubstratencontact 3264 1448 3264 1448 0 FILL_1__1759_.vdd
rlabel metal1 3244 1202 3276 1218 0 FILL_1__1759_.gnd
rlabel nsubstratencontact 3244 1448 3244 1448 0 FILL_0__1759_.vdd
rlabel metal1 3224 1202 3256 1218 0 FILL_0__1759_.gnd
rlabel metal1 3264 1202 3336 1218 0 _1759_.gnd
rlabel metal1 3264 1442 3336 1458 0 _1759_.vdd
rlabel metal2 3313 1273 3327 1287 0 _1759_.A
rlabel metal2 3293 1313 3307 1327 0 _1759_.Y
rlabel nsubstratencontact 3356 1448 3356 1448 0 FILL_1__1817_.vdd
rlabel metal1 3344 1202 3376 1218 0 FILL_1__1817_.gnd
rlabel nsubstratencontact 3336 1448 3336 1448 0 FILL_0__1817_.vdd
rlabel metal1 3324 1202 3356 1218 0 FILL_0__1817_.gnd
rlabel metal1 3364 1202 3436 1218 0 _1817_.gnd
rlabel metal1 3364 1442 3436 1458 0 _1817_.vdd
rlabel metal2 3373 1273 3387 1287 0 _1817_.A
rlabel metal2 3393 1313 3407 1327 0 _1817_.Y
rlabel nsubstratencontact 3464 1448 3464 1448 0 FILL_1__1894_.vdd
rlabel metal1 3444 1202 3476 1218 0 FILL_1__1894_.gnd
rlabel nsubstratencontact 3444 1448 3444 1448 0 FILL_0__1894_.vdd
rlabel metal1 3424 1202 3456 1218 0 FILL_0__1894_.gnd
rlabel metal1 3464 1202 3556 1218 0 _1894_.gnd
rlabel metal1 3464 1442 3556 1458 0 _1894_.vdd
rlabel metal2 3533 1293 3547 1307 0 _1894_.A
rlabel metal2 3493 1293 3507 1307 0 _1894_.Y
rlabel nsubstratencontact 3604 1448 3604 1448 0 FILL_2__1826_.vdd
rlabel metal1 3584 1202 3616 1218 0 FILL_2__1826_.gnd
rlabel nsubstratencontact 3584 1448 3584 1448 0 FILL_1__1826_.vdd
rlabel metal1 3564 1202 3596 1218 0 FILL_1__1826_.gnd
rlabel nsubstratencontact 3564 1448 3564 1448 0 FILL_0__1826_.vdd
rlabel metal1 3544 1202 3576 1218 0 FILL_0__1826_.gnd
rlabel metal1 3604 1202 3716 1218 0 _1826_.gnd
rlabel metal1 3604 1442 3716 1458 0 _1826_.vdd
rlabel metal2 3693 1313 3707 1327 0 _1826_.A
rlabel metal2 3673 1273 3687 1287 0 _1826_.B
rlabel metal2 3653 1313 3667 1327 0 _1826_.C
rlabel metal2 3633 1293 3647 1307 0 _1826_.Y
rlabel nsubstratencontact 3736 1448 3736 1448 0 FILL_1__1825_.vdd
rlabel metal1 3724 1202 3756 1218 0 FILL_1__1825_.gnd
rlabel nsubstratencontact 3716 1448 3716 1448 0 FILL_0__1825_.vdd
rlabel metal1 3704 1202 3736 1218 0 FILL_0__1825_.gnd
rlabel metal1 3744 1202 3856 1218 0 _1825_.gnd
rlabel metal1 3744 1442 3856 1458 0 _1825_.vdd
rlabel metal2 3753 1293 3767 1307 0 _1825_.A
rlabel metal2 3773 1313 3787 1327 0 _1825_.B
rlabel metal2 3813 1313 3827 1327 0 _1825_.C
rlabel metal2 3793 1293 3807 1307 0 _1825_.Y
rlabel nsubstratencontact 3884 1448 3884 1448 0 FILL_1__1776_.vdd
rlabel metal1 3864 1202 3896 1218 0 FILL_1__1776_.gnd
rlabel nsubstratencontact 3864 1448 3864 1448 0 FILL_0__1776_.vdd
rlabel metal1 3844 1202 3876 1218 0 FILL_0__1776_.gnd
rlabel metal1 3884 1202 3956 1218 0 _1776_.gnd
rlabel metal1 3884 1442 3956 1458 0 _1776_.vdd
rlabel metal2 3933 1273 3947 1287 0 _1776_.A
rlabel metal2 3913 1313 3927 1327 0 _1776_.Y
rlabel nsubstratencontact 3984 1448 3984 1448 0 FILL_1__1792_.vdd
rlabel metal1 3964 1202 3996 1218 0 FILL_1__1792_.gnd
rlabel nsubstratencontact 3964 1448 3964 1448 0 FILL_0__1792_.vdd
rlabel metal1 3944 1202 3976 1218 0 FILL_0__1792_.gnd
rlabel metal1 3984 1202 4096 1218 0 _1792_.gnd
rlabel metal1 3984 1442 4096 1458 0 _1792_.vdd
rlabel metal2 4073 1293 4087 1307 0 _1792_.A
rlabel metal2 4053 1313 4067 1327 0 _1792_.B
rlabel metal2 4013 1313 4027 1327 0 _1792_.C
rlabel metal2 4033 1293 4047 1307 0 _1792_.Y
rlabel nsubstratencontact 4124 1448 4124 1448 0 FILL_1__1791_.vdd
rlabel metal1 4104 1202 4136 1218 0 FILL_1__1791_.gnd
rlabel nsubstratencontact 4104 1448 4104 1448 0 FILL_0__1791_.vdd
rlabel metal1 4084 1202 4116 1218 0 FILL_0__1791_.gnd
rlabel metal1 4124 1202 4236 1218 0 _1791_.gnd
rlabel metal1 4124 1442 4236 1458 0 _1791_.vdd
rlabel metal2 4213 1293 4227 1307 0 _1791_.A
rlabel metal2 4193 1313 4207 1327 0 _1791_.B
rlabel metal2 4153 1313 4167 1327 0 _1791_.C
rlabel metal2 4173 1293 4187 1307 0 _1791_.Y
rlabel nsubstratencontact 4264 1448 4264 1448 0 FILL_1__1790_.vdd
rlabel metal1 4244 1202 4276 1218 0 FILL_1__1790_.gnd
rlabel nsubstratencontact 4244 1448 4244 1448 0 FILL_0__1790_.vdd
rlabel metal1 4224 1202 4256 1218 0 FILL_0__1790_.gnd
rlabel metal1 4264 1202 4376 1218 0 _1790_.gnd
rlabel metal1 4264 1442 4376 1458 0 _1790_.vdd
rlabel metal2 4353 1313 4367 1327 0 _1790_.A
rlabel metal2 4333 1273 4347 1287 0 _1790_.B
rlabel metal2 4313 1313 4327 1327 0 _1790_.C
rlabel metal2 4293 1293 4307 1307 0 _1790_.Y
rlabel nsubstratencontact 4404 1448 4404 1448 0 FILL_1__1789_.vdd
rlabel metal1 4384 1202 4416 1218 0 FILL_1__1789_.gnd
rlabel nsubstratencontact 4384 1448 4384 1448 0 FILL_0__1789_.vdd
rlabel metal1 4364 1202 4396 1218 0 FILL_0__1789_.gnd
rlabel metal1 4404 1202 4516 1218 0 _1789_.gnd
rlabel metal1 4404 1442 4516 1458 0 _1789_.vdd
rlabel metal2 4493 1293 4507 1307 0 _1789_.A
rlabel metal2 4473 1313 4487 1327 0 _1789_.B
rlabel metal2 4433 1313 4447 1327 0 _1789_.C
rlabel metal2 4453 1293 4467 1307 0 _1789_.Y
rlabel nsubstratencontact 4536 1448 4536 1448 0 FILL_1__1807_.vdd
rlabel metal1 4524 1202 4556 1218 0 FILL_1__1807_.gnd
rlabel nsubstratencontact 4516 1448 4516 1448 0 FILL_0__1807_.vdd
rlabel metal1 4504 1202 4536 1218 0 FILL_0__1807_.gnd
rlabel nsubstratencontact 4556 1448 4556 1448 0 FILL_2__1807_.vdd
rlabel metal1 4544 1202 4576 1218 0 FILL_2__1807_.gnd
rlabel nsubstratencontact 4676 1448 4676 1448 0 FILL_0__1802_.vdd
rlabel metal1 4664 1202 4696 1218 0 FILL_0__1802_.gnd
rlabel metal1 4564 1202 4676 1218 0 _1807_.gnd
rlabel metal1 4564 1442 4676 1458 0 _1807_.vdd
rlabel metal2 4573 1293 4587 1307 0 _1807_.A
rlabel metal2 4593 1313 4607 1327 0 _1807_.B
rlabel metal2 4633 1313 4647 1327 0 _1807_.C
rlabel metal2 4613 1293 4627 1307 0 _1807_.Y
rlabel nsubstratencontact 4696 1448 4696 1448 0 FILL_1__1802_.vdd
rlabel metal1 4684 1202 4716 1218 0 FILL_1__1802_.gnd
rlabel nsubstratencontact 4796 1448 4796 1448 0 FILL_0__1841_.vdd
rlabel metal1 4784 1202 4816 1218 0 FILL_0__1841_.gnd
rlabel metal1 4704 1202 4796 1218 0 _1802_.gnd
rlabel metal1 4704 1442 4796 1458 0 _1802_.vdd
rlabel metal2 4713 1333 4727 1347 0 _1802_.A
rlabel metal2 4753 1333 4767 1347 0 _1802_.B
rlabel metal2 4733 1313 4747 1327 0 _1802_.Y
rlabel nsubstratencontact 4816 1448 4816 1448 0 FILL_1__1841_.vdd
rlabel metal1 4804 1202 4836 1218 0 FILL_1__1841_.gnd
rlabel metal1 4824 1202 4936 1218 0 _1841_.gnd
rlabel metal1 4824 1442 4936 1458 0 _1841_.vdd
rlabel metal2 4833 1293 4847 1307 0 _1841_.A
rlabel metal2 4853 1313 4867 1327 0 _1841_.B
rlabel metal2 4893 1313 4907 1327 0 _1841_.C
rlabel metal2 4873 1293 4887 1307 0 _1841_.Y
rlabel nsubstratencontact 4956 1448 4956 1448 0 FILL_1__1705_.vdd
rlabel metal1 4944 1202 4976 1218 0 FILL_1__1705_.gnd
rlabel nsubstratencontact 5056 1448 5056 1448 0 FILL_0__1836_.vdd
rlabel metal1 5044 1202 5076 1218 0 FILL_0__1836_.gnd
rlabel nsubstratencontact 4936 1448 4936 1448 0 FILL_0__1705_.vdd
rlabel metal1 4924 1202 4956 1218 0 FILL_0__1705_.gnd
rlabel metal1 4964 1202 5056 1218 0 _1705_.gnd
rlabel metal1 4964 1442 5056 1458 0 _1705_.vdd
rlabel metal2 5013 1293 5027 1307 0 _1705_.B
rlabel metal2 4973 1293 4987 1307 0 _1705_.A
rlabel metal2 4993 1273 5007 1287 0 _1705_.Y
rlabel nsubstratencontact 5076 1448 5076 1448 0 FILL_1__1836_.vdd
rlabel metal1 5064 1202 5096 1218 0 FILL_1__1836_.gnd
rlabel nsubstratencontact 5184 1448 5184 1448 0 FILL_0__1714_.vdd
rlabel metal1 5164 1202 5196 1218 0 FILL_0__1714_.gnd
rlabel metal1 5084 1202 5176 1218 0 _1836_.gnd
rlabel metal1 5084 1442 5176 1458 0 _1836_.vdd
rlabel metal2 5093 1333 5107 1347 0 _1836_.A
rlabel metal2 5133 1333 5147 1347 0 _1836_.B
rlabel metal2 5113 1313 5127 1327 0 _1836_.Y
rlabel nsubstratencontact 5204 1448 5204 1448 0 FILL_1__1714_.vdd
rlabel metal1 5184 1202 5216 1218 0 FILL_1__1714_.gnd
rlabel nsubstratencontact 5304 1448 5304 1448 0 FILL_0__1720_.vdd
rlabel metal1 5284 1202 5316 1218 0 FILL_0__1720_.gnd
rlabel metal1 5204 1202 5296 1218 0 _1714_.gnd
rlabel metal1 5204 1442 5296 1458 0 _1714_.vdd
rlabel metal2 5273 1333 5287 1347 0 _1714_.A
rlabel metal2 5233 1333 5247 1347 0 _1714_.B
rlabel metal2 5253 1313 5267 1327 0 _1714_.Y
rlabel nsubstratencontact 5324 1448 5324 1448 0 FILL_1__1720_.vdd
rlabel metal1 5304 1202 5336 1218 0 FILL_1__1720_.gnd
rlabel nsubstratencontact 5436 1448 5436 1448 0 FILL_0__1687_.vdd
rlabel metal1 5424 1202 5456 1218 0 FILL_0__1687_.gnd
rlabel metal1 5324 1202 5436 1218 0 _1720_.gnd
rlabel metal1 5324 1442 5436 1458 0 _1720_.vdd
rlabel metal2 5413 1293 5427 1307 0 _1720_.A
rlabel metal2 5393 1313 5407 1327 0 _1720_.B
rlabel metal2 5353 1313 5367 1327 0 _1720_.C
rlabel metal2 5373 1293 5387 1307 0 _1720_.Y
rlabel nsubstratencontact 5456 1448 5456 1448 0 FILL_1__1687_.vdd
rlabel metal1 5444 1202 5476 1218 0 FILL_1__1687_.gnd
rlabel metal1 5464 1202 5576 1218 0 _1687_.gnd
rlabel metal1 5464 1442 5576 1458 0 _1687_.vdd
rlabel metal2 5473 1293 5487 1307 0 _1687_.A
rlabel metal2 5493 1313 5507 1327 0 _1687_.B
rlabel metal2 5533 1313 5547 1327 0 _1687_.C
rlabel metal2 5513 1293 5527 1307 0 _1687_.Y
rlabel metal1 5624 1202 5736 1218 0 _1702_.gnd
rlabel metal1 5624 1442 5736 1458 0 _1702_.vdd
rlabel metal2 5633 1293 5647 1307 0 _1702_.A
rlabel metal2 5653 1313 5667 1327 0 _1702_.B
rlabel metal2 5693 1313 5707 1327 0 _1702_.C
rlabel metal2 5673 1293 5687 1307 0 _1702_.Y
rlabel nsubstratencontact 5736 1448 5736 1448 0 FILL85950x18150.vdd
rlabel metal1 5724 1202 5756 1218 0 FILL85950x18150.gnd
rlabel nsubstratencontact 5756 1448 5756 1448 0 FILL86250x18150.vdd
rlabel metal1 5744 1202 5776 1218 0 FILL86250x18150.gnd
rlabel nsubstratencontact 5776 1448 5776 1448 0 FILL86550x18150.vdd
rlabel metal1 5764 1202 5796 1218 0 FILL86550x18150.gnd
rlabel nsubstratencontact 5796 1448 5796 1448 0 FILL86850x18150.vdd
rlabel metal1 5784 1202 5816 1218 0 FILL86850x18150.gnd
rlabel nsubstratencontact 5576 1448 5576 1448 0 FILL_0__1702_.vdd
rlabel metal1 5564 1202 5596 1218 0 FILL_0__1702_.gnd
rlabel nsubstratencontact 5596 1448 5596 1448 0 FILL_1__1702_.vdd
rlabel metal1 5584 1202 5616 1218 0 FILL_1__1702_.gnd
rlabel nsubstratencontact 5616 1448 5616 1448 0 FILL_2__1702_.vdd
rlabel metal1 5604 1202 5636 1218 0 FILL_2__1702_.gnd
rlabel nsubstratencontact 56 1452 56 1452 0 FILL_2__1050_.vdd
rlabel metal1 44 1682 76 1698 0 FILL_2__1050_.gnd
rlabel nsubstratencontact 36 1452 36 1452 0 FILL_1__1050_.vdd
rlabel metal1 24 1682 56 1698 0 FILL_1__1050_.gnd
rlabel nsubstratencontact 16 1452 16 1452 0 FILL_0__1050_.vdd
rlabel metal1 4 1682 36 1698 0 FILL_0__1050_.gnd
rlabel metal1 64 1682 176 1698 0 _1050_.gnd
rlabel metal1 64 1442 176 1458 0 _1050_.vdd
rlabel metal2 73 1573 87 1587 0 _1050_.A
rlabel metal2 93 1553 107 1567 0 _1050_.B
rlabel metal2 113 1573 127 1587 0 _1050_.C
rlabel metal2 133 1553 147 1567 0 _1050_.Y
rlabel nsubstratencontact 204 1452 204 1452 0 FILL_1__1117_.vdd
rlabel metal1 184 1682 216 1698 0 FILL_1__1117_.gnd
rlabel nsubstratencontact 184 1452 184 1452 0 FILL_0__1117_.vdd
rlabel metal1 164 1682 196 1698 0 FILL_0__1117_.gnd
rlabel metal1 204 1682 316 1698 0 _1117_.gnd
rlabel metal1 204 1442 316 1458 0 _1117_.vdd
rlabel metal2 293 1573 307 1587 0 _1117_.A
rlabel metal2 273 1553 287 1567 0 _1117_.B
rlabel metal2 253 1573 267 1587 0 _1117_.C
rlabel metal2 233 1553 247 1567 0 _1117_.Y
rlabel nsubstratencontact 336 1452 336 1452 0 FILL_1__1124_.vdd
rlabel metal1 324 1682 356 1698 0 FILL_1__1124_.gnd
rlabel nsubstratencontact 316 1452 316 1452 0 FILL_0__1124_.vdd
rlabel metal1 304 1682 336 1698 0 FILL_0__1124_.gnd
rlabel metal1 344 1682 456 1698 0 _1124_.gnd
rlabel metal1 344 1442 456 1458 0 _1124_.vdd
rlabel metal2 353 1573 367 1587 0 _1124_.A
rlabel metal2 373 1613 387 1627 0 _1124_.B
rlabel metal2 393 1573 407 1587 0 _1124_.C
rlabel metal2 413 1593 427 1607 0 _1124_.Y
rlabel nsubstratencontact 484 1452 484 1452 0 FILL_1__1352_.vdd
rlabel metal1 464 1682 496 1698 0 FILL_1__1352_.gnd
rlabel nsubstratencontact 464 1452 464 1452 0 FILL_0__1352_.vdd
rlabel metal1 444 1682 476 1698 0 FILL_0__1352_.gnd
rlabel metal1 484 1682 596 1698 0 _1352_.gnd
rlabel metal1 484 1442 596 1458 0 _1352_.vdd
rlabel metal2 573 1573 587 1587 0 _1352_.A
rlabel metal2 553 1613 567 1627 0 _1352_.B
rlabel metal2 533 1573 547 1587 0 _1352_.C
rlabel metal2 513 1593 527 1607 0 _1352_.Y
rlabel nsubstratencontact 616 1452 616 1452 0 FILL_1__1284_.vdd
rlabel metal1 604 1682 636 1698 0 FILL_1__1284_.gnd
rlabel nsubstratencontact 596 1452 596 1452 0 FILL_0__1284_.vdd
rlabel metal1 584 1682 616 1698 0 FILL_0__1284_.gnd
rlabel metal1 624 1682 716 1698 0 _1284_.gnd
rlabel metal1 624 1442 716 1458 0 _1284_.vdd
rlabel metal2 633 1553 647 1567 0 _1284_.A
rlabel metal2 673 1553 687 1567 0 _1284_.B
rlabel metal2 653 1573 667 1587 0 _1284_.Y
rlabel nsubstratencontact 736 1452 736 1452 0 FILL_1__1251_.vdd
rlabel metal1 724 1682 756 1698 0 FILL_1__1251_.gnd
rlabel nsubstratencontact 716 1452 716 1452 0 FILL_0__1251_.vdd
rlabel metal1 704 1682 736 1698 0 FILL_0__1251_.gnd
rlabel metal1 744 1682 816 1698 0 _1251_.gnd
rlabel metal1 744 1442 816 1458 0 _1251_.vdd
rlabel metal2 753 1613 767 1627 0 _1251_.A
rlabel metal2 773 1573 787 1587 0 _1251_.Y
rlabel nsubstratencontact 844 1452 844 1452 0 FILL_1__1194_.vdd
rlabel metal1 824 1682 856 1698 0 FILL_1__1194_.gnd
rlabel nsubstratencontact 824 1452 824 1452 0 FILL_0__1194_.vdd
rlabel metal1 804 1682 836 1698 0 FILL_0__1194_.gnd
rlabel metal1 844 1682 956 1698 0 _1194_.gnd
rlabel metal1 844 1442 956 1458 0 _1194_.vdd
rlabel metal2 933 1593 947 1607 0 _1194_.A
rlabel metal2 913 1573 927 1587 0 _1194_.B
rlabel metal2 873 1573 887 1587 0 _1194_.C
rlabel metal2 893 1593 907 1607 0 _1194_.Y
rlabel nsubstratencontact 984 1452 984 1452 0 FILL_1__1110_.vdd
rlabel metal1 964 1682 996 1698 0 FILL_1__1110_.gnd
rlabel nsubstratencontact 964 1452 964 1452 0 FILL_0__1110_.vdd
rlabel metal1 944 1682 976 1698 0 FILL_0__1110_.gnd
rlabel metal1 984 1682 1096 1698 0 _1110_.gnd
rlabel metal1 984 1442 1096 1458 0 _1110_.vdd
rlabel metal2 1073 1573 1087 1587 0 _1110_.A
rlabel metal2 1053 1553 1067 1567 0 _1110_.B
rlabel metal2 1033 1573 1047 1587 0 _1110_.C
rlabel metal2 1013 1553 1027 1567 0 _1110_.Y
rlabel nsubstratencontact 1124 1452 1124 1452 0 FILL_1__1108_.vdd
rlabel metal1 1104 1682 1136 1698 0 FILL_1__1108_.gnd
rlabel nsubstratencontact 1104 1452 1104 1452 0 FILL_0__1108_.vdd
rlabel metal1 1084 1682 1116 1698 0 FILL_0__1108_.gnd
rlabel nsubstratencontact 1216 1452 1216 1452 0 FILL_0__1193_.vdd
rlabel metal1 1204 1682 1236 1698 0 FILL_0__1193_.gnd
rlabel metal1 1124 1682 1216 1698 0 _1108_.gnd
rlabel metal1 1124 1442 1216 1458 0 _1108_.vdd
rlabel metal2 1193 1553 1207 1567 0 _1108_.A
rlabel metal2 1153 1553 1167 1567 0 _1108_.B
rlabel metal2 1173 1573 1187 1587 0 _1108_.Y
rlabel nsubstratencontact 1256 1452 1256 1452 0 FILL_2__1193_.vdd
rlabel metal1 1244 1682 1276 1698 0 FILL_2__1193_.gnd
rlabel nsubstratencontact 1236 1452 1236 1452 0 FILL_1__1193_.vdd
rlabel metal1 1224 1682 1256 1698 0 FILL_1__1193_.gnd
rlabel metal1 1264 1682 1356 1698 0 _1193_.gnd
rlabel metal1 1264 1442 1356 1458 0 _1193_.vdd
rlabel metal2 1313 1593 1327 1607 0 _1193_.B
rlabel metal2 1273 1593 1287 1607 0 _1193_.A
rlabel metal2 1293 1613 1307 1627 0 _1193_.Y
rlabel nsubstratencontact 1384 1452 1384 1452 0 FILL_1__1890_.vdd
rlabel metal1 1364 1682 1396 1698 0 FILL_1__1890_.gnd
rlabel nsubstratencontact 1364 1452 1364 1452 0 FILL_0__1890_.vdd
rlabel metal1 1344 1682 1376 1698 0 FILL_0__1890_.gnd
rlabel metal1 1384 1682 1476 1698 0 _1890_.gnd
rlabel metal1 1384 1442 1476 1458 0 _1890_.vdd
rlabel metal2 1453 1593 1467 1607 0 _1890_.A
rlabel metal2 1413 1593 1427 1607 0 _1890_.Y
rlabel nsubstratencontact 1524 1452 1524 1452 0 FILL_2__1082_.vdd
rlabel metal1 1504 1682 1536 1698 0 FILL_2__1082_.gnd
rlabel nsubstratencontact 1504 1452 1504 1452 0 FILL_1__1082_.vdd
rlabel metal1 1484 1682 1516 1698 0 FILL_1__1082_.gnd
rlabel nsubstratencontact 1484 1452 1484 1452 0 FILL_0__1082_.vdd
rlabel metal1 1464 1682 1496 1698 0 FILL_0__1082_.gnd
rlabel metal1 1524 1682 1596 1698 0 _1082_.gnd
rlabel metal1 1524 1442 1596 1458 0 _1082_.vdd
rlabel metal2 1573 1613 1587 1627 0 _1082_.A
rlabel metal2 1553 1573 1567 1587 0 _1082_.Y
rlabel metal1 1624 1682 1756 1698 0 _1201_.gnd
rlabel metal1 1624 1442 1756 1458 0 _1201_.vdd
rlabel metal2 1633 1593 1647 1607 0 _1201_.A
rlabel metal2 1653 1573 1667 1587 0 _1201_.B
rlabel metal2 1713 1593 1727 1607 0 _1201_.C
rlabel metal2 1693 1573 1707 1587 0 _1201_.D
rlabel metal2 1673 1593 1687 1607 0 _1201_.Y
rlabel metal1 1744 1682 2236 1698 0 _1661_.gnd
rlabel metal1 1744 1442 2236 1458 0 _1661_.vdd
rlabel metal2 2153 1573 2167 1587 0 _1661_.S
rlabel metal2 2033 1613 2047 1627 0 _1661_.D
rlabel metal2 1853 1573 1867 1587 0 _1661_.CLK
rlabel metal2 2193 1553 2207 1567 0 _1661_.R
rlabel metal2 1773 1573 1787 1587 0 _1661_.Q
rlabel nsubstratencontact 1596 1452 1596 1452 0 FILL_0__1201_.vdd
rlabel metal1 1584 1682 1616 1698 0 FILL_0__1201_.gnd
rlabel nsubstratencontact 1616 1452 1616 1452 0 FILL_1__1201_.vdd
rlabel metal1 1604 1682 1636 1698 0 FILL_1__1201_.gnd
rlabel metal1 2424 1682 2516 1698 0 _1277_.gnd
rlabel metal1 2424 1442 2516 1458 0 _1277_.vdd
rlabel metal2 2433 1553 2447 1567 0 _1277_.A
rlabel metal2 2473 1553 2487 1567 0 _1277_.B
rlabel metal2 2453 1573 2467 1587 0 _1277_.Y
rlabel metal1 2284 1682 2396 1698 0 _1278_.gnd
rlabel metal1 2284 1442 2396 1458 0 _1278_.vdd
rlabel metal2 2293 1593 2307 1607 0 _1278_.A
rlabel metal2 2313 1573 2327 1587 0 _1278_.B
rlabel metal2 2353 1573 2367 1587 0 _1278_.C
rlabel metal2 2333 1593 2347 1607 0 _1278_.Y
rlabel nsubstratencontact 2396 1452 2396 1452 0 FILL_0__1277_.vdd
rlabel metal1 2384 1682 2416 1698 0 FILL_0__1277_.gnd
rlabel nsubstratencontact 2236 1452 2236 1452 0 FILL_0__1278_.vdd
rlabel metal1 2224 1682 2256 1698 0 FILL_0__1278_.gnd
rlabel nsubstratencontact 2524 1452 2524 1452 0 FILL_0__1534_.vdd
rlabel metal1 2504 1682 2536 1698 0 FILL_0__1534_.gnd
rlabel nsubstratencontact 2416 1452 2416 1452 0 FILL_1__1277_.vdd
rlabel metal1 2404 1682 2436 1698 0 FILL_1__1277_.gnd
rlabel nsubstratencontact 2256 1452 2256 1452 0 FILL_1__1278_.vdd
rlabel metal1 2244 1682 2276 1698 0 FILL_1__1278_.gnd
rlabel nsubstratencontact 2544 1452 2544 1452 0 FILL_1__1534_.vdd
rlabel metal1 2524 1682 2556 1698 0 FILL_1__1534_.gnd
rlabel nsubstratencontact 2276 1452 2276 1452 0 FILL_2__1278_.vdd
rlabel metal1 2264 1682 2296 1698 0 FILL_2__1278_.gnd
rlabel nsubstratencontact 2664 1452 2664 1452 0 FILL_0__1535_.vdd
rlabel metal1 2644 1682 2676 1698 0 FILL_0__1535_.gnd
rlabel metal1 2544 1682 2656 1698 0 _1534_.gnd
rlabel metal1 2544 1442 2656 1458 0 _1534_.vdd
rlabel metal2 2633 1593 2647 1607 0 _1534_.A
rlabel metal2 2613 1573 2627 1587 0 _1534_.B
rlabel metal2 2573 1573 2587 1587 0 _1534_.C
rlabel metal2 2593 1593 2607 1607 0 _1534_.Y
rlabel nsubstratencontact 2684 1452 2684 1452 0 FILL_1__1535_.vdd
rlabel metal1 2664 1682 2696 1698 0 FILL_1__1535_.gnd
rlabel nsubstratencontact 2784 1452 2784 1452 0 FILL_0__1276_.vdd
rlabel metal1 2764 1682 2796 1698 0 FILL_0__1276_.gnd
rlabel metal1 2684 1682 2776 1698 0 _1535_.gnd
rlabel metal1 2684 1442 2776 1458 0 _1535_.vdd
rlabel metal2 2753 1553 2767 1567 0 _1535_.A
rlabel metal2 2713 1553 2727 1567 0 _1535_.B
rlabel metal2 2733 1573 2747 1587 0 _1535_.Y
rlabel nsubstratencontact 2804 1452 2804 1452 0 FILL_1__1276_.vdd
rlabel metal1 2784 1682 2816 1698 0 FILL_1__1276_.gnd
rlabel metal1 2804 1682 2916 1698 0 _1276_.gnd
rlabel metal1 2804 1442 2916 1458 0 _1276_.vdd
rlabel metal2 2893 1593 2907 1607 0 _1276_.A
rlabel metal2 2873 1573 2887 1587 0 _1276_.B
rlabel metal2 2833 1573 2847 1587 0 _1276_.C
rlabel metal2 2853 1593 2867 1607 0 _1276_.Y
rlabel nsubstratencontact 2944 1452 2944 1452 0 FILL_1__1536_.vdd
rlabel metal1 2924 1682 2956 1698 0 FILL_1__1536_.gnd
rlabel nsubstratencontact 2924 1452 2924 1452 0 FILL_0__1536_.vdd
rlabel metal1 2904 1682 2936 1698 0 FILL_0__1536_.gnd
rlabel metal1 2944 1682 3056 1698 0 _1536_.gnd
rlabel metal1 2944 1442 3056 1458 0 _1536_.vdd
rlabel metal2 3033 1593 3047 1607 0 _1536_.A
rlabel metal2 3013 1573 3027 1587 0 _1536_.B
rlabel metal2 2973 1573 2987 1587 0 _1536_.C
rlabel metal2 2993 1593 3007 1607 0 _1536_.Y
rlabel metal1 3044 1682 3536 1698 0 _1665_.gnd
rlabel metal1 3044 1442 3536 1458 0 _1665_.vdd
rlabel metal2 3113 1573 3127 1587 0 _1665_.S
rlabel metal2 3233 1613 3247 1627 0 _1665_.D
rlabel metal2 3413 1573 3427 1587 0 _1665_.CLK
rlabel metal2 3073 1553 3087 1567 0 _1665_.R
rlabel metal2 3493 1573 3507 1587 0 _1665_.Q
rlabel nsubstratencontact 3544 1452 3544 1452 0 FILL_0__1843_.vdd
rlabel metal1 3524 1682 3556 1698 0 FILL_0__1843_.gnd
rlabel nsubstratencontact 3564 1452 3564 1452 0 FILL_1__1843_.vdd
rlabel metal1 3544 1682 3576 1698 0 FILL_1__1843_.gnd
rlabel metal1 3564 1682 3676 1698 0 _1843_.gnd
rlabel metal1 3564 1442 3676 1458 0 _1843_.vdd
rlabel metal2 3653 1573 3667 1587 0 _1843_.A
rlabel metal2 3633 1613 3647 1627 0 _1843_.B
rlabel metal2 3613 1573 3627 1587 0 _1843_.C
rlabel metal2 3593 1593 3607 1607 0 _1843_.Y
rlabel nsubstratencontact 3696 1452 3696 1452 0 FILL_1__1842_.vdd
rlabel metal1 3684 1682 3716 1698 0 FILL_1__1842_.gnd
rlabel nsubstratencontact 3676 1452 3676 1452 0 FILL_0__1842_.vdd
rlabel metal1 3664 1682 3696 1698 0 FILL_0__1842_.gnd
rlabel metal1 3704 1682 3816 1698 0 _1842_.gnd
rlabel metal1 3704 1442 3816 1458 0 _1842_.vdd
rlabel metal2 3713 1593 3727 1607 0 _1842_.A
rlabel metal2 3733 1573 3747 1587 0 _1842_.B
rlabel metal2 3773 1573 3787 1587 0 _1842_.C
rlabel metal2 3753 1593 3767 1607 0 _1842_.Y
rlabel nsubstratencontact 3844 1452 3844 1452 0 FILL_1__1896_.vdd
rlabel metal1 3824 1682 3856 1698 0 FILL_1__1896_.gnd
rlabel nsubstratencontact 3824 1452 3824 1452 0 FILL_0__1896_.vdd
rlabel metal1 3804 1682 3836 1698 0 FILL_0__1896_.gnd
rlabel metal1 3844 1682 3936 1698 0 _1896_.gnd
rlabel metal1 3844 1442 3936 1458 0 _1896_.vdd
rlabel metal2 3913 1593 3927 1607 0 _1896_.A
rlabel metal2 3873 1593 3887 1607 0 _1896_.Y
rlabel nsubstratencontact 3964 1452 3964 1452 0 FILL_1__1784_.vdd
rlabel metal1 3944 1682 3976 1698 0 FILL_1__1784_.gnd
rlabel nsubstratencontact 3944 1452 3944 1452 0 FILL_0__1784_.vdd
rlabel metal1 3924 1682 3956 1698 0 FILL_0__1784_.gnd
rlabel metal1 3964 1682 4076 1698 0 _1784_.gnd
rlabel metal1 3964 1442 4076 1458 0 _1784_.vdd
rlabel metal2 4053 1593 4067 1607 0 _1784_.A
rlabel metal2 3993 1593 4007 1607 0 _1784_.Y
rlabel metal2 4013 1553 4027 1567 0 _1784_.B
rlabel nsubstratencontact 4096 1452 4096 1452 0 FILL_1__1785_.vdd
rlabel metal1 4084 1682 4116 1698 0 FILL_1__1785_.gnd
rlabel nsubstratencontact 4204 1452 4204 1452 0 FILL_0__1786_.vdd
rlabel metal1 4184 1682 4216 1698 0 FILL_0__1786_.gnd
rlabel nsubstratencontact 4076 1452 4076 1452 0 FILL_0__1785_.vdd
rlabel metal1 4064 1682 4096 1698 0 FILL_0__1785_.gnd
rlabel metal1 4104 1682 4196 1698 0 _1785_.gnd
rlabel metal1 4104 1442 4196 1458 0 _1785_.vdd
rlabel metal2 4113 1553 4127 1567 0 _1785_.A
rlabel metal2 4153 1553 4167 1567 0 _1785_.B
rlabel metal2 4133 1573 4147 1587 0 _1785_.Y
rlabel nsubstratencontact 4224 1452 4224 1452 0 FILL_1__1786_.vdd
rlabel metal1 4204 1682 4236 1698 0 FILL_1__1786_.gnd
rlabel metal1 4224 1682 4356 1698 0 _1786_.gnd
rlabel metal1 4224 1442 4356 1458 0 _1786_.vdd
rlabel metal2 4333 1593 4347 1607 0 _1786_.A
rlabel metal2 4313 1573 4327 1587 0 _1786_.B
rlabel metal2 4253 1593 4267 1607 0 _1786_.C
rlabel metal2 4273 1573 4287 1587 0 _1786_.D
rlabel metal2 4293 1593 4307 1607 0 _1786_.Y
rlabel nsubstratencontact 4384 1452 4384 1452 0 FILL_1__1805_.vdd
rlabel metal1 4364 1682 4396 1698 0 FILL_1__1805_.gnd
rlabel nsubstratencontact 4364 1452 4364 1452 0 FILL_0__1805_.vdd
rlabel metal1 4344 1682 4376 1698 0 FILL_0__1805_.gnd
rlabel metal1 4384 1682 4516 1698 0 _1805_.gnd
rlabel metal1 4384 1442 4516 1458 0 _1805_.vdd
rlabel metal2 4493 1593 4507 1607 0 _1805_.A
rlabel metal2 4473 1573 4487 1587 0 _1805_.B
rlabel metal2 4413 1593 4427 1607 0 _1805_.C
rlabel metal2 4433 1573 4447 1587 0 _1805_.D
rlabel metal2 4453 1593 4467 1607 0 _1805_.Y
rlabel nsubstratencontact 4556 1452 4556 1452 0 FILL_2__1839_.vdd
rlabel metal1 4544 1682 4576 1698 0 FILL_2__1839_.gnd
rlabel nsubstratencontact 4536 1452 4536 1452 0 FILL_1__1839_.vdd
rlabel metal1 4524 1682 4556 1698 0 FILL_1__1839_.gnd
rlabel nsubstratencontact 4516 1452 4516 1452 0 FILL_0__1839_.vdd
rlabel metal1 4504 1682 4536 1698 0 FILL_0__1839_.gnd
rlabel nsubstratencontact 4696 1452 4696 1452 0 FILL_0__1838_.vdd
rlabel metal1 4684 1682 4716 1698 0 FILL_0__1838_.gnd
rlabel metal1 4564 1682 4696 1698 0 _1839_.gnd
rlabel metal1 4564 1442 4696 1458 0 _1839_.vdd
rlabel metal2 4573 1593 4587 1607 0 _1839_.A
rlabel metal2 4593 1573 4607 1587 0 _1839_.B
rlabel metal2 4653 1593 4667 1607 0 _1839_.C
rlabel metal2 4633 1573 4647 1587 0 _1839_.D
rlabel metal2 4613 1593 4627 1607 0 _1839_.Y
rlabel nsubstratencontact 4836 1452 4836 1452 0 FILL_1__1840_.vdd
rlabel metal1 4824 1682 4856 1698 0 FILL_1__1840_.gnd
rlabel nsubstratencontact 4716 1452 4716 1452 0 FILL_1__1838_.vdd
rlabel metal1 4704 1682 4736 1698 0 FILL_1__1838_.gnd
rlabel nsubstratencontact 4816 1452 4816 1452 0 FILL_0__1840_.vdd
rlabel metal1 4804 1682 4836 1698 0 FILL_0__1840_.gnd
rlabel metal1 4724 1682 4816 1698 0 _1838_.gnd
rlabel metal1 4724 1442 4816 1458 0 _1838_.vdd
rlabel metal2 4733 1553 4747 1567 0 _1838_.A
rlabel metal2 4773 1553 4787 1567 0 _1838_.B
rlabel metal2 4753 1573 4767 1587 0 _1838_.Y
rlabel nsubstratencontact 4984 1452 4984 1452 0 FILL_1__1837_.vdd
rlabel metal1 4964 1682 4996 1698 0 FILL_1__1837_.gnd
rlabel nsubstratencontact 4964 1452 4964 1452 0 FILL_0__1837_.vdd
rlabel metal1 4944 1682 4976 1698 0 FILL_0__1837_.gnd
rlabel metal1 4844 1682 4956 1698 0 _1840_.gnd
rlabel metal1 4844 1442 4956 1458 0 _1840_.vdd
rlabel metal2 4853 1593 4867 1607 0 _1840_.A
rlabel metal2 4873 1573 4887 1587 0 _1840_.B
rlabel metal2 4913 1573 4927 1587 0 _1840_.C
rlabel metal2 4893 1593 4907 1607 0 _1840_.Y
rlabel metal1 4984 1682 5096 1698 0 _1837_.gnd
rlabel metal1 4984 1442 5096 1458 0 _1837_.vdd
rlabel metal2 5073 1593 5087 1607 0 _1837_.A
rlabel metal2 5013 1593 5027 1607 0 _1837_.Y
rlabel metal2 5033 1553 5047 1567 0 _1837_.B
rlabel nsubstratencontact 5136 1452 5136 1452 0 FILL_2__1715_.vdd
rlabel metal1 5124 1682 5156 1698 0 FILL_2__1715_.gnd
rlabel nsubstratencontact 5116 1452 5116 1452 0 FILL_1__1715_.vdd
rlabel metal1 5104 1682 5136 1698 0 FILL_1__1715_.gnd
rlabel nsubstratencontact 5096 1452 5096 1452 0 FILL_0__1715_.vdd
rlabel metal1 5084 1682 5116 1698 0 FILL_0__1715_.gnd
rlabel metal1 5144 1682 5256 1698 0 _1715_.gnd
rlabel metal1 5144 1442 5256 1458 0 _1715_.vdd
rlabel metal2 5153 1573 5167 1587 0 _1715_.A
rlabel metal2 5173 1553 5187 1567 0 _1715_.B
rlabel metal2 5193 1573 5207 1587 0 _1715_.C
rlabel metal2 5213 1553 5227 1567 0 _1715_.Y
rlabel nsubstratencontact 5276 1452 5276 1452 0 FILL_1__1716_.vdd
rlabel metal1 5264 1682 5296 1698 0 FILL_1__1716_.gnd
rlabel nsubstratencontact 5256 1452 5256 1452 0 FILL_0__1716_.vdd
rlabel metal1 5244 1682 5276 1698 0 FILL_0__1716_.gnd
rlabel metal1 5284 1682 5416 1698 0 _1716_.gnd
rlabel metal1 5284 1442 5416 1458 0 _1716_.vdd
rlabel metal2 5293 1593 5307 1607 0 _1716_.A
rlabel metal2 5313 1573 5327 1587 0 _1716_.B
rlabel metal2 5373 1593 5387 1607 0 _1716_.C
rlabel metal2 5353 1573 5367 1587 0 _1716_.D
rlabel metal2 5333 1593 5347 1607 0 _1716_.Y
rlabel nsubstratencontact 5436 1452 5436 1452 0 FILL_1__1700_.vdd
rlabel metal1 5424 1682 5456 1698 0 FILL_1__1700_.gnd
rlabel nsubstratencontact 5416 1452 5416 1452 0 FILL_0__1700_.vdd
rlabel metal1 5404 1682 5436 1698 0 FILL_0__1700_.gnd
rlabel metal1 5444 1682 5536 1698 0 _1700_.gnd
rlabel metal1 5444 1442 5536 1458 0 _1700_.vdd
rlabel metal2 5453 1553 5467 1567 0 _1700_.A
rlabel metal2 5493 1553 5507 1567 0 _1700_.B
rlabel metal2 5473 1573 5487 1587 0 _1700_.Y
rlabel nsubstratencontact 5556 1452 5556 1452 0 FILL_1__1732_.vdd
rlabel metal1 5544 1682 5576 1698 0 FILL_1__1732_.gnd
rlabel nsubstratencontact 5536 1452 5536 1452 0 FILL_0__1732_.vdd
rlabel metal1 5524 1682 5556 1698 0 FILL_0__1732_.gnd
rlabel metal1 5724 1682 5796 1698 0 _1696_.gnd
rlabel metal1 5724 1442 5796 1458 0 _1696_.vdd
rlabel metal2 5773 1573 5787 1587 0 _1696_.A
rlabel metal2 5753 1593 5767 1607 0 _1696_.Y
rlabel metal1 5564 1682 5676 1698 0 _1732_.gnd
rlabel metal1 5564 1442 5676 1458 0 _1732_.vdd
rlabel metal2 5573 1573 5587 1587 0 _1732_.A
rlabel metal2 5593 1553 5607 1567 0 _1732_.B
rlabel metal2 5613 1573 5627 1587 0 _1732_.C
rlabel metal2 5633 1553 5647 1567 0 _1732_.Y
rlabel nsubstratencontact 5804 1452 5804 1452 0 FILL86850x21750.vdd
rlabel metal1 5784 1682 5816 1698 0 FILL86850x21750.gnd
rlabel nsubstratencontact 5684 1452 5684 1452 0 FILL_0__1696_.vdd
rlabel metal1 5664 1682 5696 1698 0 FILL_0__1696_.gnd
rlabel nsubstratencontact 5704 1452 5704 1452 0 FILL_1__1696_.vdd
rlabel metal1 5684 1682 5716 1698 0 FILL_1__1696_.gnd
rlabel nsubstratencontact 5724 1452 5724 1452 0 FILL_2__1696_.vdd
rlabel metal1 5704 1682 5736 1698 0 FILL_2__1696_.gnd
rlabel nsubstratencontact 44 1928 44 1928 0 FILL_1__1258_.vdd
rlabel metal1 24 1682 56 1698 0 FILL_1__1258_.gnd
rlabel nsubstratencontact 24 1928 24 1928 0 FILL_0__1258_.vdd
rlabel metal1 4 1682 36 1698 0 FILL_0__1258_.gnd
rlabel metal1 44 1682 156 1698 0 _1258_.gnd
rlabel metal1 44 1922 156 1938 0 _1258_.vdd
rlabel metal2 133 1793 147 1807 0 _1258_.A
rlabel metal2 113 1813 127 1827 0 _1258_.B
rlabel metal2 93 1793 107 1807 0 _1258_.C
rlabel metal2 73 1813 87 1827 0 _1258_.Y
rlabel nsubstratencontact 176 1928 176 1928 0 FILL_1__1250_.vdd
rlabel metal1 164 1682 196 1698 0 FILL_1__1250_.gnd
rlabel nsubstratencontact 156 1928 156 1928 0 FILL_0__1250_.vdd
rlabel metal1 144 1682 176 1698 0 FILL_0__1250_.gnd
rlabel metal1 184 1682 296 1698 0 _1250_.gnd
rlabel metal1 184 1922 296 1938 0 _1250_.vdd
rlabel metal2 193 1793 207 1807 0 _1250_.A
rlabel metal2 213 1753 227 1767 0 _1250_.B
rlabel metal2 233 1793 247 1807 0 _1250_.C
rlabel metal2 253 1773 267 1787 0 _1250_.Y
rlabel nsubstratencontact 324 1928 324 1928 0 FILL_1__1353_.vdd
rlabel metal1 304 1682 336 1698 0 FILL_1__1353_.gnd
rlabel nsubstratencontact 304 1928 304 1928 0 FILL_0__1353_.vdd
rlabel metal1 284 1682 316 1698 0 FILL_0__1353_.gnd
rlabel metal1 324 1682 436 1698 0 _1353_.gnd
rlabel metal1 324 1922 436 1938 0 _1353_.vdd
rlabel metal2 413 1773 427 1787 0 _1353_.A
rlabel metal2 393 1793 407 1807 0 _1353_.B
rlabel metal2 353 1793 367 1807 0 _1353_.C
rlabel metal2 373 1773 387 1787 0 _1353_.Y
rlabel nsubstratencontact 464 1928 464 1928 0 FILL_1__1245_.vdd
rlabel metal1 444 1682 476 1698 0 FILL_1__1245_.gnd
rlabel nsubstratencontact 444 1928 444 1928 0 FILL_0__1245_.vdd
rlabel metal1 424 1682 456 1698 0 FILL_0__1245_.gnd
rlabel metal1 464 1682 576 1698 0 _1245_.gnd
rlabel metal1 464 1922 576 1938 0 _1245_.vdd
rlabel metal2 553 1793 567 1807 0 _1245_.A
rlabel metal2 533 1813 547 1827 0 _1245_.B
rlabel metal2 513 1793 527 1807 0 _1245_.C
rlabel metal2 493 1813 507 1827 0 _1245_.Y
rlabel nsubstratencontact 624 1928 624 1928 0 FILL_2__1285_.vdd
rlabel metal1 604 1682 636 1698 0 FILL_2__1285_.gnd
rlabel nsubstratencontact 604 1928 604 1928 0 FILL_1__1285_.vdd
rlabel metal1 584 1682 616 1698 0 FILL_1__1285_.gnd
rlabel nsubstratencontact 584 1928 584 1928 0 FILL_0__1285_.vdd
rlabel metal1 564 1682 596 1698 0 FILL_0__1285_.gnd
rlabel metal1 624 1682 716 1698 0 _1285_.gnd
rlabel metal1 624 1922 716 1938 0 _1285_.vdd
rlabel metal2 653 1773 667 1787 0 _1285_.B
rlabel metal2 693 1773 707 1787 0 _1285_.A
rlabel metal2 673 1753 687 1767 0 _1285_.Y
rlabel nsubstratencontact 736 1928 736 1928 0 FILL_1__1286_.vdd
rlabel metal1 724 1682 756 1698 0 FILL_1__1286_.gnd
rlabel nsubstratencontact 716 1928 716 1928 0 FILL_0__1286_.vdd
rlabel metal1 704 1682 736 1698 0 FILL_0__1286_.gnd
rlabel metal1 744 1682 856 1698 0 _1286_.gnd
rlabel metal1 744 1922 856 1938 0 _1286_.vdd
rlabel metal2 753 1793 767 1807 0 _1286_.A
rlabel metal2 773 1753 787 1767 0 _1286_.B
rlabel metal2 793 1793 807 1807 0 _1286_.C
rlabel metal2 813 1773 827 1787 0 _1286_.Y
rlabel nsubstratencontact 884 1928 884 1928 0 FILL_1__1102_.vdd
rlabel metal1 864 1682 896 1698 0 FILL_1__1102_.gnd
rlabel nsubstratencontact 864 1928 864 1928 0 FILL_0__1102_.vdd
rlabel metal1 844 1682 876 1698 0 FILL_0__1102_.gnd
rlabel nsubstratencontact 1024 1928 1024 1928 0 FILL_2__1109_.vdd
rlabel metal1 1004 1682 1036 1698 0 FILL_2__1109_.gnd
rlabel nsubstratencontact 904 1928 904 1928 0 FILL_2__1102_.vdd
rlabel metal1 884 1682 916 1698 0 FILL_2__1102_.gnd
rlabel nsubstratencontact 1004 1928 1004 1928 0 FILL_1__1109_.vdd
rlabel metal1 984 1682 1016 1698 0 FILL_1__1109_.gnd
rlabel nsubstratencontact 984 1928 984 1928 0 FILL_0__1109_.vdd
rlabel metal1 964 1682 996 1698 0 FILL_0__1109_.gnd
rlabel metal1 904 1682 976 1698 0 _1102_.gnd
rlabel metal1 904 1922 976 1938 0 _1102_.vdd
rlabel metal2 953 1753 967 1767 0 _1102_.A
rlabel metal2 933 1793 947 1807 0 _1102_.Y
rlabel nsubstratencontact 1144 1928 1144 1928 0 FILL_0__1103_.vdd
rlabel metal1 1124 1682 1156 1698 0 FILL_0__1103_.gnd
rlabel metal1 1024 1682 1136 1698 0 _1109_.gnd
rlabel metal1 1024 1922 1136 1938 0 _1109_.vdd
rlabel metal2 1113 1773 1127 1787 0 _1109_.A
rlabel metal2 1093 1793 1107 1807 0 _1109_.B
rlabel metal2 1053 1793 1067 1807 0 _1109_.C
rlabel metal2 1073 1773 1087 1787 0 _1109_.Y
rlabel nsubstratencontact 1164 1928 1164 1928 0 FILL_1__1103_.vdd
rlabel metal1 1144 1682 1176 1698 0 FILL_1__1103_.gnd
rlabel metal1 1164 1682 1276 1698 0 _1103_.gnd
rlabel metal1 1164 1922 1276 1938 0 _1103_.vdd
rlabel metal2 1253 1773 1267 1787 0 _1103_.A
rlabel metal2 1233 1793 1247 1807 0 _1103_.B
rlabel metal2 1193 1793 1207 1807 0 _1103_.C
rlabel metal2 1213 1773 1227 1787 0 _1103_.Y
rlabel nsubstratencontact 1304 1928 1304 1928 0 FILL_1__1105_.vdd
rlabel metal1 1284 1682 1316 1698 0 FILL_1__1105_.gnd
rlabel nsubstratencontact 1404 1928 1404 1928 0 FILL_1__1020_.vdd
rlabel metal1 1384 1682 1416 1698 0 FILL_1__1020_.gnd
rlabel nsubstratencontact 1284 1928 1284 1928 0 FILL_0__1105_.vdd
rlabel metal1 1264 1682 1296 1698 0 FILL_0__1105_.gnd
rlabel nsubstratencontact 1384 1928 1384 1928 0 FILL_0__1020_.vdd
rlabel metal1 1364 1682 1396 1698 0 FILL_0__1020_.gnd
rlabel metal1 1304 1682 1376 1698 0 _1105_.gnd
rlabel metal1 1304 1922 1376 1938 0 _1105_.vdd
rlabel metal2 1353 1753 1367 1767 0 _1105_.A
rlabel metal2 1333 1793 1347 1807 0 _1105_.Y
rlabel nsubstratencontact 1516 1928 1516 1928 0 FILL_0__1091_.vdd
rlabel metal1 1504 1682 1536 1698 0 FILL_0__1091_.gnd
rlabel metal1 1404 1682 1516 1698 0 _1020_.gnd
rlabel metal1 1404 1922 1516 1938 0 _1020_.vdd
rlabel metal2 1493 1773 1507 1787 0 _1020_.A
rlabel metal2 1473 1793 1487 1807 0 _1020_.B
rlabel metal2 1433 1793 1447 1807 0 _1020_.C
rlabel metal2 1453 1773 1467 1787 0 _1020_.Y
rlabel nsubstratencontact 1536 1928 1536 1928 0 FILL_1__1091_.vdd
rlabel metal1 1524 1682 1556 1698 0 FILL_1__1091_.gnd
rlabel metal1 1544 1682 1656 1698 0 _1091_.gnd
rlabel metal1 1544 1922 1656 1938 0 _1091_.vdd
rlabel metal2 1553 1773 1567 1787 0 _1091_.A
rlabel metal2 1573 1793 1587 1807 0 _1091_.B
rlabel metal2 1613 1793 1627 1807 0 _1091_.C
rlabel metal2 1593 1773 1607 1787 0 _1091_.Y
rlabel nsubstratencontact 1684 1928 1684 1928 0 FILL_1__1080_.vdd
rlabel metal1 1664 1682 1696 1698 0 FILL_1__1080_.gnd
rlabel nsubstratencontact 1664 1928 1664 1928 0 FILL_0__1080_.vdd
rlabel metal1 1644 1682 1676 1698 0 FILL_0__1080_.gnd
rlabel metal1 1684 1682 1796 1698 0 _1080_.gnd
rlabel metal1 1684 1922 1796 1938 0 _1080_.vdd
rlabel metal2 1773 1773 1787 1787 0 _1080_.A
rlabel metal2 1753 1793 1767 1807 0 _1080_.B
rlabel metal2 1713 1793 1727 1807 0 _1080_.C
rlabel metal2 1733 1773 1747 1787 0 _1080_.Y
rlabel nsubstratencontact 1824 1928 1824 1928 0 FILL_1__1104_.vdd
rlabel metal1 1804 1682 1836 1698 0 FILL_1__1104_.gnd
rlabel nsubstratencontact 1804 1928 1804 1928 0 FILL_0__1104_.vdd
rlabel metal1 1784 1682 1816 1698 0 FILL_0__1104_.gnd
rlabel metal1 1824 1682 1916 1698 0 _1104_.gnd
rlabel metal1 1824 1922 1916 1938 0 _1104_.vdd
rlabel metal2 1893 1813 1907 1827 0 _1104_.A
rlabel metal2 1853 1813 1867 1827 0 _1104_.B
rlabel metal2 1873 1793 1887 1807 0 _1104_.Y
rlabel nsubstratencontact 1944 1928 1944 1928 0 FILL_1__1099_.vdd
rlabel metal1 1924 1682 1956 1698 0 FILL_1__1099_.gnd
rlabel nsubstratencontact 1924 1928 1924 1928 0 FILL_0__1099_.vdd
rlabel metal1 1904 1682 1936 1698 0 FILL_0__1099_.gnd
rlabel metal1 1944 1682 2036 1698 0 _1099_.gnd
rlabel metal1 1944 1922 2036 1938 0 _1099_.vdd
rlabel metal2 2013 1813 2027 1827 0 _1099_.A
rlabel metal2 1973 1813 1987 1827 0 _1099_.B
rlabel metal2 1993 1793 2007 1807 0 _1099_.Y
rlabel metal1 2084 1682 2176 1698 0 _1043_.gnd
rlabel metal1 2084 1922 2176 1938 0 _1043_.vdd
rlabel metal2 2153 1793 2167 1807 0 _1043_.A
rlabel metal2 2113 1793 2127 1807 0 _1043_.Y
rlabel metal1 2164 1682 2656 1698 0 _1664_.gnd
rlabel metal1 2164 1922 2656 1938 0 _1664_.vdd
rlabel metal2 2573 1793 2587 1807 0 _1664_.S
rlabel metal2 2453 1753 2467 1767 0 _1664_.D
rlabel metal2 2273 1793 2287 1807 0 _1664_.CLK
rlabel metal2 2613 1813 2627 1827 0 _1664_.R
rlabel metal2 2193 1793 2207 1807 0 _1664_.Q
rlabel nsubstratencontact 2044 1928 2044 1928 0 FILL_0__1043_.vdd
rlabel metal1 2024 1682 2056 1698 0 FILL_0__1043_.gnd
rlabel nsubstratencontact 2064 1928 2064 1928 0 FILL_1__1043_.vdd
rlabel metal1 2044 1682 2076 1698 0 FILL_1__1043_.gnd
rlabel nsubstratencontact 2084 1928 2084 1928 0 FILL_2__1043_.vdd
rlabel metal1 2064 1682 2096 1698 0 FILL_2__1043_.gnd
rlabel metal1 2684 1682 2776 1698 0 _1066_.gnd
rlabel metal1 2684 1922 2776 1938 0 _1066_.vdd
rlabel metal2 2693 1813 2707 1827 0 _1066_.A
rlabel metal2 2733 1813 2747 1827 0 _1066_.B
rlabel metal2 2713 1793 2727 1807 0 _1066_.Y
rlabel metal1 2804 1682 2916 1698 0 _1275_.gnd
rlabel metal1 2804 1922 2916 1938 0 _1275_.vdd
rlabel metal2 2893 1793 2907 1807 0 _1275_.A
rlabel metal2 2873 1813 2887 1827 0 _1275_.B
rlabel metal2 2853 1793 2867 1807 0 _1275_.C
rlabel metal2 2833 1813 2847 1827 0 _1275_.Y
rlabel metal1 2944 1682 3056 1698 0 _1432_.gnd
rlabel metal1 2944 1922 3056 1938 0 _1432_.vdd
rlabel metal2 3033 1773 3047 1787 0 _1432_.A
rlabel metal2 3013 1793 3027 1807 0 _1432_.B
rlabel metal2 2973 1793 2987 1807 0 _1432_.C
rlabel metal2 2993 1773 3007 1787 0 _1432_.Y
rlabel nsubstratencontact 2656 1928 2656 1928 0 FILL_0__1066_.vdd
rlabel metal1 2644 1682 2676 1698 0 FILL_0__1066_.gnd
rlabel nsubstratencontact 2784 1928 2784 1928 0 FILL_0__1275_.vdd
rlabel metal1 2764 1682 2796 1698 0 FILL_0__1275_.gnd
rlabel nsubstratencontact 2924 1928 2924 1928 0 FILL_0__1432_.vdd
rlabel metal1 2904 1682 2936 1698 0 FILL_0__1432_.gnd
rlabel nsubstratencontact 2676 1928 2676 1928 0 FILL_1__1066_.vdd
rlabel metal1 2664 1682 2696 1698 0 FILL_1__1066_.gnd
rlabel nsubstratencontact 2804 1928 2804 1928 0 FILL_1__1275_.vdd
rlabel metal1 2784 1682 2816 1698 0 FILL_1__1275_.gnd
rlabel nsubstratencontact 2944 1928 2944 1928 0 FILL_1__1432_.vdd
rlabel metal1 2924 1682 2956 1698 0 FILL_1__1432_.gnd
rlabel nsubstratencontact 3076 1928 3076 1928 0 FILL_1__1430_.vdd
rlabel metal1 3064 1682 3096 1698 0 FILL_1__1430_.gnd
rlabel nsubstratencontact 3056 1928 3056 1928 0 FILL_0__1430_.vdd
rlabel metal1 3044 1682 3076 1698 0 FILL_0__1430_.gnd
rlabel nsubstratencontact 3176 1928 3176 1928 0 FILL_0__1281_.vdd
rlabel metal1 3164 1682 3196 1698 0 FILL_0__1281_.gnd
rlabel metal1 3084 1682 3176 1698 0 _1430_.gnd
rlabel metal1 3084 1922 3176 1938 0 _1430_.vdd
rlabel metal2 3133 1773 3147 1787 0 _1430_.B
rlabel metal2 3093 1773 3107 1787 0 _1430_.A
rlabel metal2 3113 1753 3127 1767 0 _1430_.Y
rlabel nsubstratencontact 3196 1928 3196 1928 0 FILL_1__1281_.vdd
rlabel metal1 3184 1682 3216 1698 0 FILL_1__1281_.gnd
rlabel metal1 3204 1682 3336 1698 0 _1281_.gnd
rlabel metal1 3204 1922 3335 1938 0 _1281_.vdd
rlabel metal2 3213 1793 3227 1807 0 _1281_.S
rlabel metal2 3233 1773 3247 1787 0 _1281_.B
rlabel metal2 3273 1793 3287 1807 0 _1281_.Y
rlabel metal2 3293 1773 3307 1787 0 _1281_.A
rlabel nsubstratencontact 3456 1928 3456 1928 0 FILL_1__1824_.vdd
rlabel metal1 3444 1682 3476 1698 0 FILL_1__1824_.gnd
rlabel nsubstratencontact 3364 1928 3364 1928 0 FILL_1__1819_.vdd
rlabel metal1 3344 1682 3376 1698 0 FILL_1__1819_.gnd
rlabel nsubstratencontact 3436 1928 3436 1928 0 FILL_0__1824_.vdd
rlabel metal1 3424 1682 3456 1698 0 FILL_0__1824_.gnd
rlabel nsubstratencontact 3344 1928 3344 1928 0 FILL_0__1819_.vdd
rlabel metal1 3324 1682 3356 1698 0 FILL_0__1819_.gnd
rlabel metal1 3464 1682 3596 1698 0 _1824_.gnd
rlabel metal1 3464 1922 3596 1938 0 _1824_.vdd
rlabel metal2 3473 1773 3487 1787 0 _1824_.A
rlabel metal2 3493 1793 3507 1807 0 _1824_.B
rlabel metal2 3553 1773 3567 1787 0 _1824_.C
rlabel metal2 3513 1773 3527 1787 0 _1824_.Y
rlabel metal2 3533 1793 3547 1807 0 _1824_.D
rlabel metal1 3364 1682 3436 1698 0 _1819_.gnd
rlabel metal1 3364 1922 3436 1938 0 _1819_.vdd
rlabel metal2 3413 1753 3427 1767 0 _1819_.A
rlabel metal2 3393 1793 3407 1807 0 _1819_.Y
rlabel nsubstratencontact 3624 1928 3624 1928 0 FILL_1__1823_.vdd
rlabel metal1 3604 1682 3636 1698 0 FILL_1__1823_.gnd
rlabel nsubstratencontact 3604 1928 3604 1928 0 FILL_0__1823_.vdd
rlabel metal1 3584 1682 3616 1698 0 FILL_0__1823_.gnd
rlabel metal1 3624 1682 3736 1698 0 _1823_.gnd
rlabel metal1 3624 1922 3736 1938 0 _1823_.vdd
rlabel metal2 3713 1773 3727 1787 0 _1823_.A
rlabel metal2 3693 1793 3707 1807 0 _1823_.B
rlabel metal2 3653 1793 3667 1807 0 _1823_.C
rlabel metal2 3673 1773 3687 1787 0 _1823_.Y
rlabel nsubstratencontact 3784 1928 3784 1928 0 FILL_2__1787_.vdd
rlabel metal1 3764 1682 3796 1698 0 FILL_2__1787_.gnd
rlabel nsubstratencontact 3764 1928 3764 1928 0 FILL_1__1787_.vdd
rlabel metal1 3744 1682 3776 1698 0 FILL_1__1787_.gnd
rlabel nsubstratencontact 3744 1928 3744 1928 0 FILL_0__1787_.vdd
rlabel metal1 3724 1682 3756 1698 0 FILL_0__1787_.gnd
rlabel metal1 3784 1682 3896 1698 0 _1787_.gnd
rlabel metal1 3784 1922 3896 1938 0 _1787_.vdd
rlabel metal2 3873 1773 3887 1787 0 _1787_.A
rlabel metal2 3853 1793 3867 1807 0 _1787_.B
rlabel metal2 3813 1793 3827 1807 0 _1787_.C
rlabel metal2 3833 1773 3847 1787 0 _1787_.Y
rlabel nsubstratencontact 3916 1928 3916 1928 0 FILL_1__1788_.vdd
rlabel metal1 3904 1682 3936 1698 0 FILL_1__1788_.gnd
rlabel nsubstratencontact 3896 1928 3896 1928 0 FILL_0__1788_.vdd
rlabel metal1 3884 1682 3916 1698 0 FILL_0__1788_.gnd
rlabel nsubstratencontact 4044 1928 4044 1928 0 FILL_0__1783_.vdd
rlabel metal1 4024 1682 4056 1698 0 FILL_0__1783_.gnd
rlabel metal1 3924 1682 4036 1698 0 _1788_.gnd
rlabel metal1 3924 1922 4036 1938 0 _1788_.vdd
rlabel metal2 3933 1773 3947 1787 0 _1788_.A
rlabel metal2 3953 1793 3967 1807 0 _1788_.B
rlabel metal2 3993 1793 4007 1807 0 _1788_.C
rlabel metal2 3973 1773 3987 1787 0 _1788_.Y
rlabel nsubstratencontact 4184 1928 4184 1928 0 FILL_1__1822_.vdd
rlabel metal1 4164 1682 4196 1698 0 FILL_1__1822_.gnd
rlabel nsubstratencontact 4064 1928 4064 1928 0 FILL_1__1783_.vdd
rlabel metal1 4044 1682 4076 1698 0 FILL_1__1783_.gnd
rlabel nsubstratencontact 4164 1928 4164 1928 0 FILL_0__1822_.vdd
rlabel metal1 4144 1682 4176 1698 0 FILL_0__1822_.gnd
rlabel metal1 4184 1682 4316 1698 0 _1822_.gnd
rlabel metal1 4184 1922 4316 1938 0 _1822_.vdd
rlabel metal2 4293 1773 4307 1787 0 _1822_.A
rlabel metal2 4273 1793 4287 1807 0 _1822_.B
rlabel metal2 4213 1773 4227 1787 0 _1822_.C
rlabel metal2 4233 1793 4247 1807 0 _1822_.D
rlabel metal2 4253 1773 4267 1787 0 _1822_.Y
rlabel metal1 4064 1682 4156 1698 0 _1783_.gnd
rlabel metal1 4064 1922 4156 1938 0 _1783_.vdd
rlabel metal2 4133 1813 4147 1827 0 _1783_.A
rlabel metal2 4093 1813 4107 1827 0 _1783_.B
rlabel metal2 4113 1793 4127 1807 0 _1783_.Y
rlabel nsubstratencontact 4344 1928 4344 1928 0 FILL_1__1804_.vdd
rlabel metal1 4324 1682 4356 1698 0 FILL_1__1804_.gnd
rlabel nsubstratencontact 4324 1928 4324 1928 0 FILL_0__1804_.vdd
rlabel metal1 4304 1682 4336 1698 0 FILL_0__1804_.gnd
rlabel nsubstratencontact 4456 1928 4456 1928 0 FILL_1__1806_.vdd
rlabel metal1 4444 1682 4476 1698 0 FILL_1__1806_.gnd
rlabel nsubstratencontact 4436 1928 4436 1928 0 FILL_0__1806_.vdd
rlabel metal1 4424 1682 4456 1698 0 FILL_0__1806_.gnd
rlabel metal1 4464 1682 4576 1698 0 _1806_.gnd
rlabel metal1 4464 1922 4576 1938 0 _1806_.vdd
rlabel metal2 4473 1773 4487 1787 0 _1806_.A
rlabel metal2 4493 1793 4507 1807 0 _1806_.B
rlabel metal2 4533 1793 4547 1807 0 _1806_.C
rlabel metal2 4513 1773 4527 1787 0 _1806_.Y
rlabel metal1 4344 1682 4436 1698 0 _1804_.gnd
rlabel metal1 4344 1922 4436 1938 0 _1804_.vdd
rlabel metal2 4413 1813 4427 1827 0 _1804_.A
rlabel metal2 4373 1813 4387 1827 0 _1804_.B
rlabel metal2 4393 1793 4407 1807 0 _1804_.Y
rlabel nsubstratencontact 4604 1928 4604 1928 0 FILL_1__1803_.vdd
rlabel metal1 4584 1682 4616 1698 0 FILL_1__1803_.gnd
rlabel nsubstratencontact 4584 1928 4584 1928 0 FILL_0__1803_.vdd
rlabel metal1 4564 1682 4596 1698 0 FILL_0__1803_.gnd
rlabel metal1 4604 1682 4716 1698 0 _1803_.gnd
rlabel metal1 4604 1922 4716 1938 0 _1803_.vdd
rlabel metal2 4693 1773 4707 1787 0 _1803_.A
rlabel metal2 4633 1773 4647 1787 0 _1803_.Y
rlabel metal2 4653 1813 4667 1827 0 _1803_.B
rlabel nsubstratencontact 4744 1928 4744 1928 0 FILL_1__1863_.vdd
rlabel metal1 4724 1682 4756 1698 0 FILL_1__1863_.gnd
rlabel nsubstratencontact 4724 1928 4724 1928 0 FILL_0__1863_.vdd
rlabel metal1 4704 1682 4736 1698 0 FILL_0__1863_.gnd
rlabel nsubstratencontact 4844 1928 4844 1928 0 FILL_0__1693_.vdd
rlabel metal1 4824 1682 4856 1698 0 FILL_0__1693_.gnd
rlabel metal1 4744 1682 4836 1698 0 _1863_.gnd
rlabel metal1 4744 1922 4836 1938 0 _1863_.vdd
rlabel metal2 4773 1773 4787 1787 0 _1863_.B
rlabel metal2 4813 1773 4827 1787 0 _1863_.A
rlabel metal2 4793 1753 4807 1767 0 _1863_.Y
rlabel nsubstratencontact 4984 1928 4984 1928 0 FILL_1__1695_.vdd
rlabel metal1 4964 1682 4996 1698 0 FILL_1__1695_.gnd
rlabel nsubstratencontact 4864 1928 4864 1928 0 FILL_1__1693_.vdd
rlabel metal1 4844 1682 4876 1698 0 FILL_1__1693_.gnd
rlabel nsubstratencontact 4964 1928 4964 1928 0 FILL_0__1695_.vdd
rlabel metal1 4944 1682 4976 1698 0 FILL_0__1695_.gnd
rlabel metal1 4984 1682 5116 1698 0 _1695_.gnd
rlabel metal1 4984 1922 5116 1938 0 _1695_.vdd
rlabel metal2 5093 1773 5107 1787 0 _1695_.A
rlabel metal2 5073 1793 5087 1807 0 _1695_.B
rlabel metal2 5013 1773 5027 1787 0 _1695_.C
rlabel metal2 5033 1793 5047 1807 0 _1695_.D
rlabel metal2 5053 1773 5067 1787 0 _1695_.Y
rlabel metal1 4864 1682 4956 1698 0 _1693_.gnd
rlabel metal1 4864 1922 4956 1938 0 _1693_.vdd
rlabel metal2 4933 1813 4947 1827 0 _1693_.A
rlabel metal2 4893 1813 4907 1827 0 _1693_.B
rlabel metal2 4913 1793 4927 1807 0 _1693_.Y
rlabel nsubstratencontact 5144 1928 5144 1928 0 FILL_1__1717_.vdd
rlabel metal1 5124 1682 5156 1698 0 FILL_1__1717_.gnd
rlabel nsubstratencontact 5124 1928 5124 1928 0 FILL_0__1717_.vdd
rlabel metal1 5104 1682 5136 1698 0 FILL_0__1717_.gnd
rlabel metal1 5144 1682 5216 1698 0 _1717_.gnd
rlabel metal1 5144 1922 5216 1938 0 _1717_.vdd
rlabel metal2 5193 1753 5207 1767 0 _1717_.A
rlabel metal2 5173 1793 5187 1807 0 _1717_.Y
rlabel nsubstratencontact 5244 1928 5244 1928 0 FILL_1__1718_.vdd
rlabel metal1 5224 1682 5256 1698 0 FILL_1__1718_.gnd
rlabel nsubstratencontact 5224 1928 5224 1928 0 FILL_0__1718_.vdd
rlabel metal1 5204 1682 5236 1698 0 FILL_0__1718_.gnd
rlabel metal1 5244 1682 5336 1698 0 _1718_.gnd
rlabel metal1 5244 1922 5336 1938 0 _1718_.vdd
rlabel metal2 5273 1773 5287 1787 0 _1718_.B
rlabel metal2 5313 1773 5327 1787 0 _1718_.A
rlabel metal2 5293 1753 5307 1767 0 _1718_.Y
rlabel nsubstratencontact 5356 1928 5356 1928 0 FILL_1__1719_.vdd
rlabel metal1 5344 1682 5376 1698 0 FILL_1__1719_.gnd
rlabel nsubstratencontact 5336 1928 5336 1928 0 FILL_0__1719_.vdd
rlabel metal1 5324 1682 5356 1698 0 FILL_0__1719_.gnd
rlabel metal1 5364 1682 5476 1698 0 _1719_.gnd
rlabel metal1 5364 1922 5476 1938 0 _1719_.vdd
rlabel metal2 5373 1773 5387 1787 0 _1719_.A
rlabel metal2 5393 1793 5407 1807 0 _1719_.B
rlabel metal2 5433 1793 5447 1807 0 _1719_.C
rlabel metal2 5413 1773 5427 1787 0 _1719_.Y
rlabel nsubstratencontact 5504 1928 5504 1928 0 FILL_1__1699_.vdd
rlabel metal1 5484 1682 5516 1698 0 FILL_1__1699_.gnd
rlabel nsubstratencontact 5484 1928 5484 1928 0 FILL_0__1699_.vdd
rlabel metal1 5464 1682 5496 1698 0 FILL_0__1699_.gnd
rlabel metal1 5504 1682 5616 1698 0 _1699_.gnd
rlabel metal1 5504 1922 5616 1938 0 _1699_.vdd
rlabel metal2 5593 1773 5607 1787 0 _1699_.A
rlabel metal2 5573 1793 5587 1807 0 _1699_.B
rlabel metal2 5533 1793 5547 1807 0 _1699_.C
rlabel metal2 5553 1773 5567 1787 0 _1699_.Y
rlabel metal1 5644 1682 5736 1698 0 _1596_.gnd
rlabel metal1 5644 1922 5736 1938 0 _1596_.vdd
rlabel metal2 5653 1793 5667 1807 0 _1596_.A
rlabel metal2 5693 1793 5707 1807 0 _1596_.Y
rlabel nsubstratencontact 5736 1928 5736 1928 0 FILL85950x25350.vdd
rlabel metal1 5724 1682 5756 1698 0 FILL85950x25350.gnd
rlabel nsubstratencontact 5756 1928 5756 1928 0 FILL86250x25350.vdd
rlabel metal1 5744 1682 5776 1698 0 FILL86250x25350.gnd
rlabel nsubstratencontact 5776 1928 5776 1928 0 FILL86550x25350.vdd
rlabel metal1 5764 1682 5796 1698 0 FILL86550x25350.gnd
rlabel nsubstratencontact 5796 1928 5796 1928 0 FILL86850x25350.vdd
rlabel metal1 5784 1682 5816 1698 0 FILL86850x25350.gnd
rlabel nsubstratencontact 5616 1928 5616 1928 0 FILL_0__1596_.vdd
rlabel metal1 5604 1682 5636 1698 0 FILL_0__1596_.gnd
rlabel nsubstratencontact 5636 1928 5636 1928 0 FILL_1__1596_.vdd
rlabel metal1 5624 1682 5656 1698 0 FILL_1__1596_.gnd
rlabel nsubstratencontact 64 1932 64 1932 0 FILL_2__1892_.vdd
rlabel metal1 44 2162 76 2178 0 FILL_2__1892_.gnd
rlabel nsubstratencontact 44 1932 44 1932 0 FILL_1__1892_.vdd
rlabel metal1 24 2162 56 2178 0 FILL_1__1892_.gnd
rlabel nsubstratencontact 24 1932 24 1932 0 FILL_0__1892_.vdd
rlabel metal1 4 2162 36 2178 0 FILL_0__1892_.gnd
rlabel metal1 64 2162 156 2178 0 _1892_.gnd
rlabel metal1 64 1922 156 1938 0 _1892_.vdd
rlabel metal2 133 2073 147 2087 0 _1892_.A
rlabel metal2 93 2073 107 2087 0 _1892_.Y
rlabel nsubstratencontact 204 1932 204 1932 0 FILL_2__1122_.vdd
rlabel metal1 184 2162 216 2178 0 FILL_2__1122_.gnd
rlabel nsubstratencontact 184 1932 184 1932 0 FILL_1__1122_.vdd
rlabel metal1 164 2162 196 2178 0 FILL_1__1122_.gnd
rlabel nsubstratencontact 164 1932 164 1932 0 FILL_0__1122_.vdd
rlabel metal1 144 2162 176 2178 0 FILL_0__1122_.gnd
rlabel metal1 204 2162 316 2178 0 _1122_.gnd
rlabel metal1 204 1922 316 1938 0 _1122_.vdd
rlabel metal2 293 2053 307 2067 0 _1122_.A
rlabel metal2 273 2033 287 2047 0 _1122_.B
rlabel metal2 253 2053 267 2067 0 _1122_.C
rlabel metal2 233 2033 247 2047 0 _1122_.Y
rlabel nsubstratencontact 336 1932 336 1932 0 FILL_1__1192_.vdd
rlabel metal1 324 2162 356 2178 0 FILL_1__1192_.gnd
rlabel nsubstratencontact 316 1932 316 1932 0 FILL_0__1192_.vdd
rlabel metal1 304 2162 336 2178 0 FILL_0__1192_.gnd
rlabel metal1 344 2162 456 2178 0 _1192_.gnd
rlabel metal1 344 1922 456 1938 0 _1192_.vdd
rlabel metal2 353 2053 367 2067 0 _1192_.A
rlabel metal2 373 2093 387 2107 0 _1192_.B
rlabel metal2 393 2053 407 2067 0 _1192_.C
rlabel metal2 413 2073 427 2087 0 _1192_.Y
rlabel nsubstratencontact 484 1932 484 1932 0 FILL_1__1054_.vdd
rlabel metal1 464 2162 496 2178 0 FILL_1__1054_.gnd
rlabel nsubstratencontact 464 1932 464 1932 0 FILL_0__1054_.vdd
rlabel metal1 444 2162 476 2178 0 FILL_0__1054_.gnd
rlabel metal1 484 2162 556 2178 0 _1054_.gnd
rlabel metal1 484 1922 556 1938 0 _1054_.vdd
rlabel metal2 533 2093 547 2107 0 _1054_.A
rlabel metal2 513 2053 527 2067 0 _1054_.Y
rlabel nsubstratencontact 584 1932 584 1932 0 FILL_1__1255_.vdd
rlabel metal1 564 2162 596 2178 0 FILL_1__1255_.gnd
rlabel nsubstratencontact 564 1932 564 1932 0 FILL_0__1255_.vdd
rlabel metal1 544 2162 576 2178 0 FILL_0__1255_.gnd
rlabel metal1 584 2162 696 2178 0 _1255_.gnd
rlabel metal1 584 1922 696 1938 0 _1255_.vdd
rlabel metal2 673 2073 687 2087 0 _1255_.A
rlabel metal2 653 2053 667 2067 0 _1255_.B
rlabel metal2 613 2053 627 2067 0 _1255_.C
rlabel metal2 633 2073 647 2087 0 _1255_.Y
rlabel nsubstratencontact 724 1932 724 1932 0 FILL_1__1254_.vdd
rlabel metal1 704 2162 736 2178 0 FILL_1__1254_.gnd
rlabel nsubstratencontact 704 1932 704 1932 0 FILL_0__1254_.vdd
rlabel metal1 684 2162 716 2178 0 FILL_0__1254_.gnd
rlabel metal1 724 2162 836 2178 0 _1254_.gnd
rlabel metal1 724 1922 836 1938 0 _1254_.vdd
rlabel metal2 813 2053 827 2067 0 _1254_.A
rlabel metal2 793 2093 807 2107 0 _1254_.B
rlabel metal2 773 2053 787 2067 0 _1254_.C
rlabel metal2 753 2073 767 2087 0 _1254_.Y
rlabel nsubstratencontact 856 1932 856 1932 0 FILL_1__1257_.vdd
rlabel metal1 844 2162 876 2178 0 FILL_1__1257_.gnd
rlabel nsubstratencontact 836 1932 836 1932 0 FILL_0__1257_.vdd
rlabel metal1 824 2162 856 2178 0 FILL_0__1257_.gnd
rlabel metal1 864 2162 976 2178 0 _1257_.gnd
rlabel metal1 864 1922 976 1938 0 _1257_.vdd
rlabel metal2 873 2053 887 2067 0 _1257_.A
rlabel metal2 893 2033 907 2047 0 _1257_.B
rlabel metal2 913 2053 927 2067 0 _1257_.C
rlabel metal2 933 2033 947 2047 0 _1257_.Y
rlabel nsubstratencontact 1024 1932 1024 1932 0 FILL_2__1252_.vdd
rlabel metal1 1004 2162 1036 2178 0 FILL_2__1252_.gnd
rlabel nsubstratencontact 1004 1932 1004 1932 0 FILL_1__1252_.vdd
rlabel metal1 984 2162 1016 2178 0 FILL_1__1252_.gnd
rlabel nsubstratencontact 984 1932 984 1932 0 FILL_0__1252_.vdd
rlabel metal1 964 2162 996 2178 0 FILL_0__1252_.gnd
rlabel nsubstratencontact 1144 1932 1144 1932 0 FILL_0__1249_.vdd
rlabel metal1 1124 2162 1156 2178 0 FILL_0__1249_.gnd
rlabel metal1 1024 2162 1136 2178 0 _1252_.gnd
rlabel metal1 1024 1922 1136 1938 0 _1252_.vdd
rlabel metal2 1113 2053 1127 2067 0 _1252_.A
rlabel metal2 1093 2033 1107 2047 0 _1252_.B
rlabel metal2 1073 2053 1087 2067 0 _1252_.C
rlabel metal2 1053 2033 1067 2047 0 _1252_.Y
rlabel nsubstratencontact 1164 1932 1164 1932 0 FILL_1__1249_.vdd
rlabel metal1 1144 2162 1176 2178 0 FILL_1__1249_.gnd
rlabel metal1 1164 2162 1276 2178 0 _1249_.gnd
rlabel metal1 1164 1922 1276 1938 0 _1249_.vdd
rlabel metal2 1253 2073 1267 2087 0 _1249_.A
rlabel metal2 1233 2053 1247 2067 0 _1249_.B
rlabel metal2 1193 2053 1207 2067 0 _1249_.C
rlabel metal2 1213 2073 1227 2087 0 _1249_.Y
rlabel nsubstratencontact 1304 1932 1304 1932 0 FILL_1__1253_.vdd
rlabel metal1 1284 2162 1316 2178 0 FILL_1__1253_.gnd
rlabel nsubstratencontact 1284 1932 1284 1932 0 FILL_0__1253_.vdd
rlabel metal1 1264 2162 1296 2178 0 FILL_0__1253_.gnd
rlabel metal1 1304 2162 1416 2178 0 _1253_.gnd
rlabel metal1 1304 1922 1416 1938 0 _1253_.vdd
rlabel metal2 1393 2073 1407 2087 0 _1253_.A
rlabel metal2 1373 2053 1387 2067 0 _1253_.B
rlabel metal2 1333 2053 1347 2067 0 _1253_.C
rlabel metal2 1353 2073 1367 2087 0 _1253_.Y
rlabel nsubstratencontact 1444 1932 1444 1932 0 FILL_1__1247_.vdd
rlabel metal1 1424 2162 1456 2178 0 FILL_1__1247_.gnd
rlabel nsubstratencontact 1424 1932 1424 1932 0 FILL_0__1247_.vdd
rlabel metal1 1404 2162 1436 2178 0 FILL_0__1247_.gnd
rlabel metal1 1444 2162 1556 2178 0 _1247_.gnd
rlabel metal1 1444 1922 1556 1938 0 _1247_.vdd
rlabel metal2 1533 2053 1547 2067 0 _1247_.A
rlabel metal2 1513 2093 1527 2107 0 _1247_.B
rlabel metal2 1493 2053 1507 2067 0 _1247_.C
rlabel metal2 1473 2073 1487 2087 0 _1247_.Y
rlabel nsubstratencontact 1584 1932 1584 1932 0 FILL_1__1244_.vdd
rlabel metal1 1564 2162 1596 2178 0 FILL_1__1244_.gnd
rlabel nsubstratencontact 1716 1932 1716 1932 0 FILL_1__1243_.vdd
rlabel metal1 1704 2162 1736 2178 0 FILL_1__1243_.gnd
rlabel nsubstratencontact 1564 1932 1564 1932 0 FILL_0__1244_.vdd
rlabel metal1 1544 2162 1576 2178 0 FILL_0__1244_.gnd
rlabel nsubstratencontact 1696 1932 1696 1932 0 FILL_0__1243_.vdd
rlabel metal1 1684 2162 1716 2178 0 FILL_0__1243_.gnd
rlabel metal1 1584 2162 1696 2178 0 _1244_.gnd
rlabel metal1 1584 1922 1696 1938 0 _1244_.vdd
rlabel metal2 1673 2053 1687 2067 0 _1244_.A
rlabel metal2 1653 2033 1667 2047 0 _1244_.B
rlabel metal2 1633 2053 1647 2067 0 _1244_.C
rlabel metal2 1613 2033 1627 2047 0 _1244_.Y
rlabel nsubstratencontact 1856 1932 1856 1932 0 FILL_1__1290_.vdd
rlabel metal1 1844 2162 1876 2178 0 FILL_1__1290_.gnd
rlabel nsubstratencontact 1836 1932 1836 1932 0 FILL_0__1290_.vdd
rlabel metal1 1824 2162 1856 2178 0 FILL_0__1290_.gnd
rlabel metal1 1864 2162 1976 2178 0 _1290_.gnd
rlabel metal1 1864 1922 1976 1938 0 _1290_.vdd
rlabel metal2 1873 2053 1887 2067 0 _1290_.A
rlabel metal2 1893 2093 1907 2107 0 _1290_.B
rlabel metal2 1913 2053 1927 2067 0 _1290_.C
rlabel metal2 1933 2073 1947 2087 0 _1290_.Y
rlabel metal1 1724 2162 1836 2178 0 _1243_.gnd
rlabel metal1 1724 1922 1836 1938 0 _1243_.vdd
rlabel metal2 1733 2073 1747 2087 0 _1243_.A
rlabel metal2 1753 2053 1767 2067 0 _1243_.B
rlabel metal2 1793 2053 1807 2067 0 _1243_.C
rlabel metal2 1773 2073 1787 2087 0 _1243_.Y
rlabel nsubstratencontact 2004 1932 2004 1932 0 FILL_1__1289_.vdd
rlabel metal1 1984 2162 2016 2178 0 FILL_1__1289_.gnd
rlabel nsubstratencontact 1984 1932 1984 1932 0 FILL_0__1289_.vdd
rlabel metal1 1964 2162 1996 2178 0 FILL_0__1289_.gnd
rlabel metal1 2004 1922 2196 1938 0 _1289_.vdd
rlabel metal2 2153 2073 2167 2087 0 _1289_.A
rlabel metal2 2113 2053 2127 2067 0 _1289_.B
rlabel metal2 2093 2073 2107 2087 0 _1289_.C
rlabel metal2 2053 2053 2067 2067 0 _1289_.Y
rlabel metal1 2004 2162 2196 2178 0 _1289_.gnd
rlabel metal1 2224 2162 2336 2178 0 _1018_.gnd
rlabel metal1 2224 1922 2336 1938 0 _1018_.vdd
rlabel metal2 2313 2053 2327 2067 0 _1018_.A
rlabel metal2 2293 2033 2307 2047 0 _1018_.B
rlabel metal2 2273 2053 2287 2067 0 _1018_.C
rlabel metal2 2253 2033 2267 2047 0 _1018_.Y
rlabel metal1 2324 2162 2816 2178 0 _1663_.gnd
rlabel metal1 2324 1922 2816 1938 0 _1663_.vdd
rlabel metal2 2733 2053 2747 2067 0 _1663_.S
rlabel metal2 2613 2093 2627 2107 0 _1663_.D
rlabel metal2 2433 2053 2447 2067 0 _1663_.CLK
rlabel metal2 2773 2033 2787 2047 0 _1663_.R
rlabel metal2 2353 2053 2367 2067 0 _1663_.Q
rlabel nsubstratencontact 2204 1932 2204 1932 0 FILL_0__1018_.vdd
rlabel metal1 2184 2162 2216 2178 0 FILL_0__1018_.gnd
rlabel nsubstratencontact 2224 1932 2224 1932 0 FILL_1__1018_.vdd
rlabel metal1 2204 2162 2236 2178 0 FILL_1__1018_.gnd
rlabel metal1 2984 2162 3076 2178 0 _1433_.gnd
rlabel metal1 2984 1922 3076 1938 0 _1433_.vdd
rlabel metal2 3053 2033 3067 2047 0 _1433_.A
rlabel metal2 3013 2033 3027 2047 0 _1433_.B
rlabel metal2 3033 2053 3047 2067 0 _1433_.Y
rlabel metal1 2844 2162 2956 2178 0 _1434_.gnd
rlabel metal1 2844 1922 2956 1938 0 _1434_.vdd
rlabel metal2 2853 2073 2867 2087 0 _1434_.A
rlabel metal2 2873 2053 2887 2067 0 _1434_.B
rlabel metal2 2913 2053 2927 2067 0 _1434_.C
rlabel metal2 2893 2073 2907 2087 0 _1434_.Y
rlabel nsubstratencontact 2964 1932 2964 1932 0 FILL_0__1433_.vdd
rlabel metal1 2944 2162 2976 2178 0 FILL_0__1433_.gnd
rlabel nsubstratencontact 2816 1932 2816 1932 0 FILL_0__1434_.vdd
rlabel metal1 2804 2162 2836 2178 0 FILL_0__1434_.gnd
rlabel nsubstratencontact 2984 1932 2984 1932 0 FILL_1__1433_.vdd
rlabel metal1 2964 2162 2996 2178 0 FILL_1__1433_.gnd
rlabel nsubstratencontact 2836 1932 2836 1932 0 FILL_1__1434_.vdd
rlabel metal1 2824 2162 2856 2178 0 FILL_1__1434_.gnd
rlabel nsubstratencontact 3096 1932 3096 1932 0 FILL_1__1570_.vdd
rlabel metal1 3084 2162 3116 2178 0 FILL_1__1570_.gnd
rlabel nsubstratencontact 3076 1932 3076 1932 0 FILL_0__1570_.vdd
rlabel metal1 3064 2162 3096 2178 0 FILL_0__1570_.gnd
rlabel metal1 3104 2162 3196 2178 0 _1570_.gnd
rlabel metal1 3104 1922 3196 1938 0 _1570_.vdd
rlabel metal2 3113 2033 3127 2047 0 _1570_.A
rlabel metal2 3153 2033 3167 2047 0 _1570_.B
rlabel metal2 3133 2053 3147 2067 0 _1570_.Y
rlabel nsubstratencontact 3236 1932 3236 1932 0 FILL_2__1540_.vdd
rlabel metal1 3224 2162 3256 2178 0 FILL_2__1540_.gnd
rlabel nsubstratencontact 3216 1932 3216 1932 0 FILL_1__1540_.vdd
rlabel metal1 3204 2162 3236 2178 0 FILL_1__1540_.gnd
rlabel nsubstratencontact 3196 1932 3196 1932 0 FILL_0__1540_.vdd
rlabel metal1 3184 2162 3216 2178 0 FILL_0__1540_.gnd
rlabel metal1 3244 2162 3336 2178 0 _1540_.gnd
rlabel metal1 3244 1922 3336 1938 0 _1540_.vdd
rlabel metal2 3293 2073 3307 2087 0 _1540_.B
rlabel metal2 3253 2073 3267 2087 0 _1540_.A
rlabel metal2 3273 2093 3287 2107 0 _1540_.Y
rlabel nsubstratencontact 3364 1932 3364 1932 0 FILL_1__1541_.vdd
rlabel metal1 3344 2162 3376 2178 0 FILL_1__1541_.gnd
rlabel nsubstratencontact 3344 1932 3344 1932 0 FILL_0__1541_.vdd
rlabel metal1 3324 2162 3356 2178 0 FILL_0__1541_.gnd
rlabel metal1 3364 2162 3476 2178 0 _1541_.gnd
rlabel metal1 3364 1922 3476 1938 0 _1541_.vdd
rlabel metal2 3453 2073 3467 2087 0 _1541_.A
rlabel metal2 3393 2073 3407 2087 0 _1541_.Y
rlabel metal2 3413 2033 3427 2047 0 _1541_.B
rlabel nsubstratencontact 3496 1932 3496 1932 0 FILL_1__1594_.vdd
rlabel metal1 3484 2162 3516 2178 0 FILL_1__1594_.gnd
rlabel nsubstratencontact 3476 1932 3476 1932 0 FILL_0__1594_.vdd
rlabel metal1 3464 2162 3496 2178 0 FILL_0__1594_.gnd
rlabel metal1 3504 2162 3616 2178 0 _1594_.gnd
rlabel metal1 3504 1922 3616 1938 0 _1594_.vdd
rlabel metal2 3513 2053 3527 2067 0 _1594_.A
rlabel metal2 3533 2093 3547 2107 0 _1594_.B
rlabel metal2 3553 2053 3567 2067 0 _1594_.C
rlabel metal2 3573 2073 3587 2087 0 _1594_.Y
rlabel nsubstratencontact 3664 1932 3664 1932 0 FILL_2__920_.vdd
rlabel metal1 3644 2162 3676 2178 0 FILL_2__920_.gnd
rlabel nsubstratencontact 3644 1932 3644 1932 0 FILL_1__920_.vdd
rlabel metal1 3624 2162 3656 2178 0 FILL_1__920_.gnd
rlabel nsubstratencontact 3624 1932 3624 1932 0 FILL_0__920_.vdd
rlabel metal1 3604 2162 3636 2178 0 FILL_0__920_.gnd
rlabel nsubstratencontact 3776 1932 3776 1932 0 FILL_2__1076_.vdd
rlabel metal1 3764 2162 3796 2178 0 FILL_2__1076_.gnd
rlabel nsubstratencontact 3756 1932 3756 1932 0 FILL_1__1076_.vdd
rlabel metal1 3744 2162 3776 2178 0 FILL_1__1076_.gnd
rlabel nsubstratencontact 3736 1932 3736 1932 0 FILL_0__1076_.vdd
rlabel metal1 3724 2162 3756 2178 0 FILL_0__1076_.gnd
rlabel metal1 3784 2162 3896 2178 0 _1076_.gnd
rlabel metal1 3784 1922 3896 1938 0 _1076_.vdd
rlabel metal2 3793 2053 3807 2067 0 _1076_.A
rlabel metal2 3813 2033 3827 2047 0 _1076_.B
rlabel metal2 3833 2053 3847 2067 0 _1076_.C
rlabel metal2 3853 2033 3867 2047 0 _1076_.Y
rlabel metal1 3664 2162 3736 2178 0 _920_.gnd
rlabel metal1 3664 1922 3736 1938 0 _920_.vdd
rlabel metal2 3713 2053 3727 2067 0 _920_.A
rlabel metal2 3693 2073 3707 2087 0 _920_.Y
rlabel nsubstratencontact 3916 1932 3916 1932 0 FILL_1__933_.vdd
rlabel metal1 3904 2162 3936 2178 0 FILL_1__933_.gnd
rlabel nsubstratencontact 3896 1932 3896 1932 0 FILL_0__933_.vdd
rlabel metal1 3884 2162 3916 2178 0 FILL_0__933_.gnd
rlabel nsubstratencontact 3936 1932 3936 1932 0 FILL_2__933_.vdd
rlabel metal1 3924 2162 3956 2178 0 FILL_2__933_.gnd
rlabel nsubstratencontact 4044 1932 4044 1932 0 FILL_1__1820_.vdd
rlabel metal1 4024 2162 4056 2178 0 FILL_1__1820_.gnd
rlabel nsubstratencontact 4024 1932 4024 1932 0 FILL_0__1820_.vdd
rlabel metal1 4004 2162 4036 2178 0 FILL_0__1820_.gnd
rlabel metal1 3944 2162 4016 2178 0 _933_.gnd
rlabel metal1 3944 1922 4016 1938 0 _933_.vdd
rlabel metal2 3953 2053 3967 2067 0 _933_.A
rlabel metal2 3973 2073 3987 2087 0 _933_.Y
rlabel nsubstratencontact 4064 1932 4064 1932 0 FILL_2__1820_.vdd
rlabel metal1 4044 2162 4076 2178 0 FILL_2__1820_.gnd
rlabel nsubstratencontact 4184 1932 4184 1932 0 FILL_0__1821_.vdd
rlabel metal1 4164 2162 4196 2178 0 FILL_0__1821_.gnd
rlabel metal1 4064 2162 4176 2178 0 _1820_.gnd
rlabel metal1 4064 1922 4176 1938 0 _1820_.vdd
rlabel metal2 4153 2073 4167 2087 0 _1820_.A
rlabel metal2 4093 2073 4107 2087 0 _1820_.Y
rlabel metal2 4113 2033 4127 2047 0 _1820_.B
rlabel nsubstratencontact 4204 1932 4204 1932 0 FILL_1__1821_.vdd
rlabel metal1 4184 2162 4216 2178 0 FILL_1__1821_.gnd
rlabel nsubstratencontact 4304 1932 4304 1932 0 FILL_0__1766_.vdd
rlabel metal1 4284 2162 4316 2178 0 FILL_0__1766_.gnd
rlabel metal1 4204 2162 4296 2178 0 _1821_.gnd
rlabel metal1 4204 1922 4296 1938 0 _1821_.vdd
rlabel metal2 4273 2033 4287 2047 0 _1821_.A
rlabel metal2 4233 2033 4247 2047 0 _1821_.B
rlabel metal2 4253 2053 4267 2067 0 _1821_.Y
rlabel nsubstratencontact 4324 1932 4324 1932 0 FILL_1__1766_.vdd
rlabel metal1 4304 2162 4336 2178 0 FILL_1__1766_.gnd
rlabel metal1 4324 2162 4436 2178 0 _1766_.gnd
rlabel metal1 4324 1922 4436 1938 0 _1766_.vdd
rlabel metal2 4413 2073 4427 2087 0 _1766_.A
rlabel metal2 4393 2053 4407 2067 0 _1766_.B
rlabel metal2 4353 2053 4367 2067 0 _1766_.C
rlabel metal2 4373 2073 4387 2087 0 _1766_.Y
rlabel nsubstratencontact 4456 1932 4456 1932 0 FILL_1__1767_.vdd
rlabel metal1 4444 2162 4476 2178 0 FILL_1__1767_.gnd
rlabel nsubstratencontact 4436 1932 4436 1932 0 FILL_0__1767_.vdd
rlabel metal1 4424 2162 4456 2178 0 FILL_0__1767_.gnd
rlabel metal1 4464 2162 4576 2178 0 _1767_.gnd
rlabel metal1 4464 1922 4576 1938 0 _1767_.vdd
rlabel metal2 4473 2073 4487 2087 0 _1767_.A
rlabel metal2 4493 2053 4507 2067 0 _1767_.B
rlabel metal2 4533 2053 4547 2067 0 _1767_.C
rlabel metal2 4513 2073 4527 2087 0 _1767_.Y
rlabel nsubstratencontact 4596 1932 4596 1932 0 FILL_1__1762_.vdd
rlabel metal1 4584 2162 4616 2178 0 FILL_1__1762_.gnd
rlabel nsubstratencontact 4576 1932 4576 1932 0 FILL_0__1762_.vdd
rlabel metal1 4564 2162 4596 2178 0 FILL_0__1762_.gnd
rlabel metal1 4604 2162 4696 2178 0 _1762_.gnd
rlabel metal1 4604 1922 4696 1938 0 _1762_.vdd
rlabel metal2 4613 2033 4627 2047 0 _1762_.A
rlabel metal2 4653 2033 4667 2047 0 _1762_.B
rlabel metal2 4633 2053 4647 2067 0 _1762_.Y
rlabel nsubstratencontact 4716 1932 4716 1932 0 FILL_1__1742_.vdd
rlabel metal1 4704 2162 4736 2178 0 FILL_1__1742_.gnd
rlabel nsubstratencontact 4696 1932 4696 1932 0 FILL_0__1742_.vdd
rlabel metal1 4684 2162 4716 2178 0 FILL_0__1742_.gnd
rlabel metal1 4724 2162 4816 2178 0 _1742_.gnd
rlabel metal1 4724 1922 4816 1938 0 _1742_.vdd
rlabel metal2 4733 2033 4747 2047 0 _1742_.A
rlabel metal2 4773 2033 4787 2047 0 _1742_.B
rlabel metal2 4753 2053 4767 2067 0 _1742_.Y
rlabel nsubstratencontact 4864 1932 4864 1932 0 FILL_2__1748_.vdd
rlabel metal1 4844 2162 4876 2178 0 FILL_2__1748_.gnd
rlabel nsubstratencontact 4844 1932 4844 1932 0 FILL_1__1748_.vdd
rlabel metal1 4824 2162 4856 2178 0 FILL_1__1748_.gnd
rlabel nsubstratencontact 4824 1932 4824 1932 0 FILL_0__1748_.vdd
rlabel metal1 4804 2162 4836 2178 0 FILL_0__1748_.gnd
rlabel metal1 4864 2162 4976 2178 0 _1748_.gnd
rlabel metal1 4864 1922 4976 1938 0 _1748_.vdd
rlabel metal2 4953 2073 4967 2087 0 _1748_.A
rlabel metal2 4933 2053 4947 2067 0 _1748_.B
rlabel metal2 4893 2053 4907 2067 0 _1748_.C
rlabel metal2 4913 2073 4927 2087 0 _1748_.Y
rlabel nsubstratencontact 5004 1932 5004 1932 0 FILL_1__1747_.vdd
rlabel metal1 4984 2162 5016 2178 0 FILL_1__1747_.gnd
rlabel nsubstratencontact 4984 1932 4984 1932 0 FILL_0__1747_.vdd
rlabel metal1 4964 2162 4996 2178 0 FILL_0__1747_.gnd
rlabel metal1 5004 2162 5116 2178 0 _1747_.gnd
rlabel metal1 5004 1922 5116 1938 0 _1747_.vdd
rlabel metal2 5093 2073 5107 2087 0 _1747_.A
rlabel metal2 5073 2053 5087 2067 0 _1747_.B
rlabel metal2 5033 2053 5047 2067 0 _1747_.C
rlabel metal2 5053 2073 5067 2087 0 _1747_.Y
rlabel nsubstratencontact 5136 1932 5136 1932 0 FILL_1__1743_.vdd
rlabel metal1 5124 2162 5156 2178 0 FILL_1__1743_.gnd
rlabel nsubstratencontact 5116 1932 5116 1932 0 FILL_0__1743_.vdd
rlabel metal1 5104 2162 5136 2178 0 FILL_0__1743_.gnd
rlabel metal1 5144 2162 5216 2178 0 _1743_.gnd
rlabel metal1 5144 1922 5216 1938 0 _1743_.vdd
rlabel metal2 5153 2093 5167 2107 0 _1743_.A
rlabel metal2 5173 2053 5187 2067 0 _1743_.Y
rlabel nsubstratencontact 5236 1932 5236 1932 0 FILL_1__1744_.vdd
rlabel metal1 5224 2162 5256 2178 0 FILL_1__1744_.gnd
rlabel nsubstratencontact 5216 1932 5216 1932 0 FILL_0__1744_.vdd
rlabel metal1 5204 2162 5236 2178 0 FILL_0__1744_.gnd
rlabel metal1 5244 2162 5336 2178 0 _1744_.gnd
rlabel metal1 5244 1922 5336 1938 0 _1744_.vdd
rlabel metal2 5293 2073 5307 2087 0 _1744_.B
rlabel metal2 5253 2073 5267 2087 0 _1744_.A
rlabel metal2 5273 2093 5287 2107 0 _1744_.Y
rlabel nsubstratencontact 5356 1932 5356 1932 0 FILL_1__1691_.vdd
rlabel metal1 5344 2162 5376 2178 0 FILL_1__1691_.gnd
rlabel nsubstratencontact 5336 1932 5336 1932 0 FILL_0__1691_.vdd
rlabel metal1 5324 2162 5356 2178 0 FILL_0__1691_.gnd
rlabel metal1 5364 2162 5456 2178 0 _1691_.gnd
rlabel metal1 5364 1922 5456 1938 0 _1691_.vdd
rlabel metal2 5373 2033 5387 2047 0 _1691_.A
rlabel metal2 5413 2033 5427 2047 0 _1691_.B
rlabel metal2 5393 2053 5407 2067 0 _1691_.Y
rlabel nsubstratencontact 5476 1932 5476 1932 0 FILL_1__1698_.vdd
rlabel metal1 5464 2162 5496 2178 0 FILL_1__1698_.gnd
rlabel nsubstratencontact 5456 1932 5456 1932 0 FILL_0__1698_.vdd
rlabel metal1 5444 2162 5476 2178 0 FILL_0__1698_.gnd
rlabel nsubstratencontact 5564 1932 5564 1932 0 FILL_0__1600_.vdd
rlabel metal1 5544 2162 5576 2178 0 FILL_0__1600_.gnd
rlabel metal1 5484 2162 5556 2178 0 _1698_.gnd
rlabel metal1 5484 1922 5556 1938 0 _1698_.vdd
rlabel metal2 5493 2093 5507 2107 0 _1698_.A
rlabel metal2 5513 2053 5527 2067 0 _1698_.Y
rlabel metal1 5584 2162 5656 2178 0 _1600_.gnd
rlabel metal1 5584 1922 5656 1938 0 _1600_.vdd
rlabel metal2 5633 2093 5647 2107 0 _1600_.A
rlabel metal2 5613 2053 5627 2067 0 _1600_.Y
rlabel metal1 5684 2162 5796 2178 0 _1730_.gnd
rlabel metal1 5684 1922 5796 1938 0 _1730_.vdd
rlabel metal2 5693 2073 5707 2087 0 _1730_.A
rlabel metal2 5713 2053 5727 2067 0 _1730_.B
rlabel metal2 5753 2053 5767 2067 0 _1730_.C
rlabel metal2 5733 2073 5747 2087 0 _1730_.Y
rlabel nsubstratencontact 5804 1932 5804 1932 0 FILL86850x28950.vdd
rlabel metal1 5784 2162 5816 2178 0 FILL86850x28950.gnd
rlabel nsubstratencontact 5656 1932 5656 1932 0 FILL_0__1730_.vdd
rlabel metal1 5644 2162 5676 2178 0 FILL_0__1730_.gnd
rlabel nsubstratencontact 5584 1932 5584 1932 0 FILL_1__1600_.vdd
rlabel metal1 5564 2162 5596 2178 0 FILL_1__1600_.gnd
rlabel nsubstratencontact 5676 1932 5676 1932 0 FILL_1__1730_.vdd
rlabel metal1 5664 2162 5696 2178 0 FILL_1__1730_.gnd
rlabel nsubstratencontact 44 2408 44 2408 0 FILL_1__1891_.vdd
rlabel metal1 24 2162 56 2178 0 FILL_1__1891_.gnd
rlabel nsubstratencontact 24 2408 24 2408 0 FILL_0__1891_.vdd
rlabel metal1 4 2162 36 2178 0 FILL_0__1891_.gnd
rlabel nsubstratencontact 144 2408 144 2408 0 FILL_0__1166_.vdd
rlabel metal1 124 2162 156 2178 0 FILL_0__1166_.gnd
rlabel metal1 44 2162 136 2178 0 _1891_.gnd
rlabel metal1 44 2402 136 2418 0 _1891_.vdd
rlabel metal2 113 2253 127 2267 0 _1891_.A
rlabel metal2 73 2253 87 2267 0 _1891_.Y
rlabel nsubstratencontact 164 2408 164 2408 0 FILL_1__1166_.vdd
rlabel metal1 144 2162 176 2178 0 FILL_1__1166_.gnd
rlabel metal1 164 2162 276 2178 0 _1166_.gnd
rlabel metal1 164 2402 276 2418 0 _1166_.vdd
rlabel metal2 253 2273 267 2287 0 _1166_.A
rlabel metal2 233 2293 247 2307 0 _1166_.B
rlabel metal2 213 2273 227 2287 0 _1166_.C
rlabel metal2 193 2293 207 2307 0 _1166_.Y
rlabel nsubstratencontact 296 2408 296 2408 0 FILL_1__1051_.vdd
rlabel metal1 284 2162 316 2178 0 FILL_1__1051_.gnd
rlabel nsubstratencontact 276 2408 276 2408 0 FILL_0__1051_.vdd
rlabel metal1 264 2162 296 2178 0 FILL_0__1051_.gnd
rlabel metal1 304 2162 396 2178 0 _1051_.gnd
rlabel metal1 304 2402 396 2418 0 _1051_.vdd
rlabel metal2 313 2293 327 2307 0 _1051_.A
rlabel metal2 353 2293 367 2307 0 _1051_.B
rlabel metal2 333 2273 347 2287 0 _1051_.Y
rlabel nsubstratencontact 416 2408 416 2408 0 FILL_1__1125_.vdd
rlabel metal1 404 2162 436 2178 0 FILL_1__1125_.gnd
rlabel nsubstratencontact 396 2408 396 2408 0 FILL_0__1125_.vdd
rlabel metal1 384 2162 416 2178 0 FILL_0__1125_.gnd
rlabel metal1 424 2162 536 2178 0 _1125_.gnd
rlabel metal1 424 2402 536 2418 0 _1125_.vdd
rlabel metal2 433 2253 447 2267 0 _1125_.A
rlabel metal2 453 2273 467 2287 0 _1125_.B
rlabel metal2 493 2273 507 2287 0 _1125_.C
rlabel metal2 473 2253 487 2267 0 _1125_.Y
rlabel nsubstratencontact 564 2408 564 2408 0 FILL_1__1256_.vdd
rlabel metal1 544 2162 576 2178 0 FILL_1__1256_.gnd
rlabel nsubstratencontact 544 2408 544 2408 0 FILL_0__1256_.vdd
rlabel metal1 524 2162 556 2178 0 FILL_0__1256_.gnd
rlabel metal1 564 2162 676 2178 0 _1256_.gnd
rlabel metal1 564 2402 676 2418 0 _1256_.vdd
rlabel metal2 653 2253 667 2267 0 _1256_.A
rlabel metal2 633 2273 647 2287 0 _1256_.B
rlabel metal2 593 2273 607 2287 0 _1256_.C
rlabel metal2 613 2253 627 2267 0 _1256_.Y
rlabel nsubstratencontact 724 2408 724 2408 0 FILL_2__1259_.vdd
rlabel metal1 704 2162 736 2178 0 FILL_2__1259_.gnd
rlabel nsubstratencontact 704 2408 704 2408 0 FILL_1__1259_.vdd
rlabel metal1 684 2162 716 2178 0 FILL_1__1259_.gnd
rlabel nsubstratencontact 684 2408 684 2408 0 FILL_0__1259_.vdd
rlabel metal1 664 2162 696 2178 0 FILL_0__1259_.gnd
rlabel metal1 724 2162 836 2178 0 _1259_.gnd
rlabel metal1 724 2402 836 2418 0 _1259_.vdd
rlabel metal2 813 2273 827 2287 0 _1259_.A
rlabel metal2 793 2293 807 2307 0 _1259_.B
rlabel metal2 773 2273 787 2287 0 _1259_.C
rlabel metal2 753 2293 767 2307 0 _1259_.Y
rlabel nsubstratencontact 864 2408 864 2408 0 FILL_1__1045_.vdd
rlabel metal1 844 2162 876 2178 0 FILL_1__1045_.gnd
rlabel nsubstratencontact 844 2408 844 2408 0 FILL_0__1045_.vdd
rlabel metal1 824 2162 856 2178 0 FILL_0__1045_.gnd
rlabel metal1 864 2162 956 2178 0 _1045_.gnd
rlabel metal1 864 2402 956 2418 0 _1045_.vdd
rlabel metal2 933 2293 947 2307 0 _1045_.A
rlabel metal2 893 2293 907 2307 0 _1045_.B
rlabel metal2 913 2273 927 2287 0 _1045_.Y
rlabel nsubstratencontact 984 2408 984 2408 0 FILL_1__1040_.vdd
rlabel metal1 964 2162 996 2178 0 FILL_1__1040_.gnd
rlabel nsubstratencontact 964 2408 964 2408 0 FILL_0__1040_.vdd
rlabel metal1 944 2162 976 2178 0 FILL_0__1040_.gnd
rlabel metal1 984 2162 1096 2178 0 _1040_.gnd
rlabel metal1 984 2402 1096 2418 0 _1040_.vdd
rlabel metal2 1073 2233 1087 2247 0 _1040_.A
rlabel metal2 1053 2253 1067 2267 0 _1040_.B
rlabel metal2 1013 2273 1027 2287 0 _1040_.Y
rlabel nsubstratencontact 1116 2408 1116 2408 0 FILL_1__1273_.vdd
rlabel metal1 1104 2162 1136 2178 0 FILL_1__1273_.gnd
rlabel nsubstratencontact 1096 2408 1096 2408 0 FILL_0__1273_.vdd
rlabel metal1 1084 2162 1116 2178 0 FILL_0__1273_.gnd
rlabel metal1 1124 2162 1196 2178 0 _1273_.gnd
rlabel metal1 1124 2402 1196 2418 0 _1273_.vdd
rlabel metal2 1133 2273 1147 2287 0 _1273_.A
rlabel metal2 1153 2253 1167 2267 0 _1273_.Y
rlabel nsubstratencontact 1224 2408 1224 2408 0 FILL_1__1240_.vdd
rlabel metal1 1204 2162 1236 2178 0 FILL_1__1240_.gnd
rlabel nsubstratencontact 1204 2408 1204 2408 0 FILL_0__1240_.vdd
rlabel metal1 1184 2162 1216 2178 0 FILL_0__1240_.gnd
rlabel metal1 1224 2162 1336 2178 0 _1240_.gnd
rlabel metal1 1224 2402 1336 2418 0 _1240_.vdd
rlabel metal2 1313 2273 1327 2287 0 _1240_.A
rlabel metal2 1293 2293 1307 2307 0 _1240_.B
rlabel metal2 1273 2273 1287 2287 0 _1240_.C
rlabel metal2 1253 2293 1267 2307 0 _1240_.Y
rlabel nsubstratencontact 1364 2408 1364 2408 0 FILL_1__1248_.vdd
rlabel metal1 1344 2162 1376 2178 0 FILL_1__1248_.gnd
rlabel nsubstratencontact 1344 2408 1344 2408 0 FILL_0__1248_.vdd
rlabel metal1 1324 2162 1356 2178 0 FILL_0__1248_.gnd
rlabel metal1 1364 2162 1476 2178 0 _1248_.gnd
rlabel metal1 1364 2402 1476 2418 0 _1248_.vdd
rlabel metal2 1453 2273 1467 2287 0 _1248_.A
rlabel metal2 1433 2233 1447 2247 0 _1248_.B
rlabel metal2 1413 2273 1427 2287 0 _1248_.C
rlabel metal2 1393 2253 1407 2267 0 _1248_.Y
rlabel nsubstratencontact 1524 2408 1524 2408 0 FILL_2__1239_.vdd
rlabel metal1 1504 2162 1536 2178 0 FILL_2__1239_.gnd
rlabel nsubstratencontact 1504 2408 1504 2408 0 FILL_1__1239_.vdd
rlabel metal1 1484 2162 1516 2178 0 FILL_1__1239_.gnd
rlabel nsubstratencontact 1484 2408 1484 2408 0 FILL_0__1239_.vdd
rlabel metal1 1464 2162 1496 2178 0 FILL_0__1239_.gnd
rlabel nsubstratencontact 1644 2408 1644 2408 0 FILL_0__1340_.vdd
rlabel metal1 1624 2162 1656 2178 0 FILL_0__1340_.gnd
rlabel metal1 1524 2162 1636 2178 0 _1239_.gnd
rlabel metal1 1524 2402 1636 2418 0 _1239_.vdd
rlabel metal2 1613 2253 1627 2267 0 _1239_.A
rlabel metal2 1593 2273 1607 2287 0 _1239_.B
rlabel metal2 1553 2273 1567 2287 0 _1239_.C
rlabel metal2 1573 2253 1587 2267 0 _1239_.Y
rlabel nsubstratencontact 1664 2408 1664 2408 0 FILL_1__1340_.vdd
rlabel metal1 1644 2162 1676 2178 0 FILL_1__1340_.gnd
rlabel nsubstratencontact 1784 2408 1784 2408 0 FILL_0__1242_.vdd
rlabel metal1 1764 2162 1796 2178 0 FILL_0__1242_.gnd
rlabel metal1 1664 2162 1776 2178 0 _1340_.gnd
rlabel metal1 1664 2402 1776 2418 0 _1340_.vdd
rlabel metal2 1753 2273 1767 2287 0 _1340_.A
rlabel metal2 1733 2233 1747 2247 0 _1340_.B
rlabel metal2 1713 2273 1727 2287 0 _1340_.C
rlabel metal2 1693 2253 1707 2267 0 _1340_.Y
rlabel nsubstratencontact 1804 2408 1804 2408 0 FILL_1__1242_.vdd
rlabel metal1 1784 2162 1816 2178 0 FILL_1__1242_.gnd
rlabel metal1 1804 2162 1916 2178 0 _1242_.gnd
rlabel metal1 1804 2402 1916 2418 0 _1242_.vdd
rlabel metal2 1893 2273 1907 2287 0 _1242_.A
rlabel metal2 1873 2293 1887 2307 0 _1242_.B
rlabel metal2 1853 2273 1867 2287 0 _1242_.C
rlabel metal2 1833 2293 1847 2307 0 _1242_.Y
rlabel nsubstratencontact 1944 2408 1944 2408 0 FILL_1__1235_.vdd
rlabel metal1 1924 2162 1956 2178 0 FILL_1__1235_.gnd
rlabel nsubstratencontact 1924 2408 1924 2408 0 FILL_0__1235_.vdd
rlabel metal1 1904 2162 1936 2178 0 FILL_0__1235_.gnd
rlabel metal1 1944 2162 2056 2178 0 _1235_.gnd
rlabel metal1 1944 2402 2056 2418 0 _1235_.vdd
rlabel metal2 2033 2273 2047 2287 0 _1235_.A
rlabel metal2 2013 2293 2027 2307 0 _1235_.B
rlabel metal2 1993 2273 2007 2287 0 _1235_.C
rlabel metal2 1973 2293 1987 2307 0 _1235_.Y
rlabel metal1 2044 2162 2536 2178 0 _1662_.gnd
rlabel metal1 2044 2402 2536 2418 0 _1662_.vdd
rlabel metal2 2453 2273 2467 2287 0 _1662_.S
rlabel metal2 2333 2233 2347 2247 0 _1662_.D
rlabel metal2 2153 2273 2167 2287 0 _1662_.CLK
rlabel metal2 2493 2293 2507 2307 0 _1662_.R
rlabel metal2 2073 2273 2087 2287 0 _1662_.Q
rlabel nsubstratencontact 2544 2408 2544 2408 0 FILL_0_BUFX2_insert9.vdd
rlabel metal1 2524 2162 2556 2178 0 FILL_0_BUFX2_insert9.gnd
rlabel nsubstratencontact 2564 2408 2564 2408 0 FILL_1_BUFX2_insert9.vdd
rlabel metal1 2544 2162 2576 2178 0 FILL_1_BUFX2_insert9.gnd
rlabel nsubstratencontact 2656 2408 2656 2408 0 FILL_0__1487_.vdd
rlabel metal1 2644 2162 2676 2178 0 FILL_0__1487_.gnd
rlabel metal1 2564 2162 2656 2178 0 BUFX2_insert9.gnd
rlabel metal1 2564 2402 2656 2418 0 BUFX2_insert9.vdd
rlabel metal2 2633 2253 2647 2267 0 BUFX2_insert9.A
rlabel metal2 2593 2253 2607 2267 0 BUFX2_insert9.Y
rlabel nsubstratencontact 2696 2408 2696 2408 0 FILL_2__1487_.vdd
rlabel metal1 2684 2162 2716 2178 0 FILL_2__1487_.gnd
rlabel nsubstratencontact 2676 2408 2676 2408 0 FILL_1__1487_.vdd
rlabel metal1 2664 2162 2696 2178 0 FILL_1__1487_.gnd
rlabel metal1 2704 2162 2816 2178 0 _1487_.gnd
rlabel metal1 2704 2402 2816 2418 0 _1487_.vdd
rlabel metal2 2713 2253 2727 2267 0 _1487_.A
rlabel metal2 2733 2273 2747 2287 0 _1487_.B
rlabel metal2 2773 2273 2787 2287 0 _1487_.C
rlabel metal2 2753 2253 2767 2267 0 _1487_.Y
rlabel nsubstratencontact 2836 2408 2836 2408 0 FILL_1__1486_.vdd
rlabel metal1 2824 2162 2856 2178 0 FILL_1__1486_.gnd
rlabel nsubstratencontact 2816 2408 2816 2408 0 FILL_0__1486_.vdd
rlabel metal1 2804 2162 2836 2178 0 FILL_0__1486_.gnd
rlabel metal1 2844 2162 2956 2178 0 _1486_.gnd
rlabel metal1 2844 2402 2956 2418 0 _1486_.vdd
rlabel metal2 2853 2253 2867 2267 0 _1486_.A
rlabel metal2 2873 2273 2887 2287 0 _1486_.B
rlabel metal2 2913 2273 2927 2287 0 _1486_.C
rlabel metal2 2893 2253 2907 2267 0 _1486_.Y
rlabel nsubstratencontact 2984 2408 2984 2408 0 FILL_1__1038_.vdd
rlabel metal1 2964 2162 2996 2178 0 FILL_1__1038_.gnd
rlabel nsubstratencontact 2964 2408 2964 2408 0 FILL_0__1038_.vdd
rlabel metal1 2944 2162 2976 2178 0 FILL_0__1038_.gnd
rlabel metal1 2984 2162 3076 2178 0 _1038_.gnd
rlabel metal1 2984 2402 3076 2418 0 _1038_.vdd
rlabel metal2 3053 2293 3067 2307 0 _1038_.A
rlabel metal2 3013 2293 3027 2307 0 _1038_.B
rlabel metal2 3033 2273 3047 2287 0 _1038_.Y
rlabel nsubstratencontact 3116 2408 3116 2408 0 FILL_2__1572_.vdd
rlabel metal1 3104 2162 3136 2178 0 FILL_2__1572_.gnd
rlabel nsubstratencontact 3096 2408 3096 2408 0 FILL_1__1572_.vdd
rlabel metal1 3084 2162 3116 2178 0 FILL_1__1572_.gnd
rlabel nsubstratencontact 3076 2408 3076 2408 0 FILL_0__1572_.vdd
rlabel metal1 3064 2162 3096 2178 0 FILL_0__1572_.gnd
rlabel metal1 3124 2162 3216 2178 0 _1572_.gnd
rlabel metal1 3124 2402 3216 2418 0 _1572_.vdd
rlabel metal2 3133 2293 3147 2307 0 _1572_.A
rlabel metal2 3173 2293 3187 2307 0 _1572_.B
rlabel metal2 3153 2273 3167 2287 0 _1572_.Y
rlabel nsubstratencontact 3244 2408 3244 2408 0 FILL_1__1282_.vdd
rlabel metal1 3224 2162 3256 2178 0 FILL_1__1282_.gnd
rlabel nsubstratencontact 3224 2408 3224 2408 0 FILL_0__1282_.vdd
rlabel metal1 3204 2162 3236 2178 0 FILL_0__1282_.gnd
rlabel metal1 3244 2162 3356 2178 0 _1282_.gnd
rlabel metal1 3244 2402 3356 2418 0 _1282_.vdd
rlabel metal2 3333 2273 3347 2287 0 _1282_.A
rlabel metal2 3313 2233 3327 2247 0 _1282_.B
rlabel metal2 3293 2273 3307 2287 0 _1282_.C
rlabel metal2 3273 2253 3287 2267 0 _1282_.Y
rlabel nsubstratencontact 3376 2408 3376 2408 0 FILL_1__1428_.vdd
rlabel metal1 3364 2162 3396 2178 0 FILL_1__1428_.gnd
rlabel nsubstratencontact 3356 2408 3356 2408 0 FILL_0__1428_.vdd
rlabel metal1 3344 2162 3376 2178 0 FILL_0__1428_.gnd
rlabel metal1 3384 2162 3476 2178 0 _1428_.gnd
rlabel metal1 3384 2402 3476 2418 0 _1428_.vdd
rlabel metal2 3433 2253 3447 2267 0 _1428_.B
rlabel metal2 3393 2253 3407 2267 0 _1428_.A
rlabel metal2 3413 2233 3427 2247 0 _1428_.Y
rlabel nsubstratencontact 3516 2408 3516 2408 0 FILL_2__1429_.vdd
rlabel metal1 3504 2162 3536 2178 0 FILL_2__1429_.gnd
rlabel nsubstratencontact 3496 2408 3496 2408 0 FILL_1__1429_.vdd
rlabel metal1 3484 2162 3516 2178 0 FILL_1__1429_.gnd
rlabel nsubstratencontact 3476 2408 3476 2408 0 FILL_0__1429_.vdd
rlabel metal1 3464 2162 3496 2178 0 FILL_0__1429_.gnd
rlabel metal1 3524 2162 3636 2178 0 _1429_.gnd
rlabel metal1 3524 2402 3636 2418 0 _1429_.vdd
rlabel metal2 3533 2253 3547 2267 0 _1429_.A
rlabel metal2 3553 2273 3567 2287 0 _1429_.B
rlabel metal2 3593 2273 3607 2287 0 _1429_.C
rlabel metal2 3573 2253 3587 2267 0 _1429_.Y
rlabel metal1 3664 2162 3756 2178 0 _1588_.gnd
rlabel metal1 3664 2402 3756 2418 0 _1588_.vdd
rlabel metal2 3673 2293 3687 2307 0 _1588_.A
rlabel metal2 3713 2293 3727 2307 0 _1588_.B
rlabel metal2 3693 2273 3707 2287 0 _1588_.Y
rlabel metal1 3864 2162 4356 2178 0 _1667_.gnd
rlabel metal1 3864 2402 4356 2418 0 _1667_.vdd
rlabel metal2 4273 2273 4287 2287 0 _1667_.S
rlabel metal2 4153 2233 4167 2247 0 _1667_.D
rlabel metal2 3973 2273 3987 2287 0 _1667_.CLK
rlabel metal2 4313 2293 4327 2307 0 _1667_.R
rlabel metal2 3893 2273 3907 2287 0 _1667_.Q
rlabel metal1 3784 2162 3876 2178 0 BUFX2_insert5.gnd
rlabel metal1 3784 2402 3876 2418 0 BUFX2_insert5.vdd
rlabel metal2 3793 2253 3807 2267 0 BUFX2_insert5.A
rlabel metal2 3833 2253 3847 2267 0 BUFX2_insert5.Y
rlabel nsubstratencontact 3636 2408 3636 2408 0 FILL_0__1588_.vdd
rlabel metal1 3624 2162 3656 2178 0 FILL_0__1588_.gnd
rlabel nsubstratencontact 3756 2408 3756 2408 0 FILL_0_BUFX2_insert5.vdd
rlabel metal1 3744 2162 3776 2178 0 FILL_0_BUFX2_insert5.gnd
rlabel nsubstratencontact 3656 2408 3656 2408 0 FILL_1__1588_.vdd
rlabel metal1 3644 2162 3676 2178 0 FILL_1__1588_.gnd
rlabel nsubstratencontact 3776 2408 3776 2408 0 FILL_1_BUFX2_insert5.vdd
rlabel metal1 3764 2162 3796 2178 0 FILL_1_BUFX2_insert5.gnd
rlabel metal1 4384 2162 4496 2178 0 _1763_.gnd
rlabel metal1 4384 2402 4496 2418 0 _1763_.vdd
rlabel metal2 4393 2253 4407 2267 0 _1763_.A
rlabel metal2 4453 2253 4467 2267 0 _1763_.Y
rlabel metal2 4433 2293 4447 2307 0 _1763_.B
rlabel metal1 4524 2162 4656 2178 0 _1765_.gnd
rlabel metal1 4524 2402 4656 2418 0 _1765_.vdd
rlabel metal2 4533 2253 4547 2267 0 _1765_.A
rlabel metal2 4553 2273 4567 2287 0 _1765_.B
rlabel metal2 4613 2253 4627 2267 0 _1765_.C
rlabel metal2 4593 2273 4607 2287 0 _1765_.D
rlabel metal2 4573 2253 4587 2267 0 _1765_.Y
rlabel nsubstratencontact 4356 2408 4356 2408 0 FILL_0__1763_.vdd
rlabel metal1 4344 2162 4376 2178 0 FILL_0__1763_.gnd
rlabel nsubstratencontact 4496 2408 4496 2408 0 FILL_0__1765_.vdd
rlabel metal1 4484 2162 4516 2178 0 FILL_0__1765_.gnd
rlabel nsubstratencontact 4376 2408 4376 2408 0 FILL_1__1763_.vdd
rlabel metal1 4364 2162 4396 2178 0 FILL_1__1763_.gnd
rlabel nsubstratencontact 4516 2408 4516 2408 0 FILL_1__1765_.vdd
rlabel metal1 4504 2162 4536 2178 0 FILL_1__1765_.gnd
rlabel nsubstratencontact 4676 2408 4676 2408 0 FILL_1__1764_.vdd
rlabel metal1 4664 2162 4696 2178 0 FILL_1__1764_.gnd
rlabel nsubstratencontact 4656 2408 4656 2408 0 FILL_0__1764_.vdd
rlabel metal1 4644 2162 4676 2178 0 FILL_0__1764_.gnd
rlabel metal1 4684 2162 4776 2178 0 _1764_.gnd
rlabel metal1 4684 2402 4776 2418 0 _1764_.vdd
rlabel metal2 4693 2293 4707 2307 0 _1764_.A
rlabel metal2 4733 2293 4747 2307 0 _1764_.B
rlabel metal2 4713 2273 4727 2287 0 _1764_.Y
rlabel nsubstratencontact 4804 2408 4804 2408 0 FILL_1_BUFX2_insert12.vdd
rlabel metal1 4784 2162 4816 2178 0 FILL_1_BUFX2_insert12.gnd
rlabel nsubstratencontact 4784 2408 4784 2408 0 FILL_0_BUFX2_insert12.vdd
rlabel metal1 4764 2162 4796 2178 0 FILL_0_BUFX2_insert12.gnd
rlabel metal1 4804 2162 4896 2178 0 BUFX2_insert12.gnd
rlabel metal1 4804 2402 4896 2418 0 BUFX2_insert12.vdd
rlabel metal2 4873 2253 4887 2267 0 BUFX2_insert12.A
rlabel metal2 4833 2253 4847 2267 0 BUFX2_insert12.Y
rlabel nsubstratencontact 4916 2408 4916 2408 0 FILL_1__1603_.vdd
rlabel metal1 4904 2162 4936 2178 0 FILL_1__1603_.gnd
rlabel nsubstratencontact 4996 2408 4996 2408 0 FILL_0__1746_.vdd
rlabel metal1 4984 2162 5016 2178 0 FILL_0__1746_.gnd
rlabel nsubstratencontact 4896 2408 4896 2408 0 FILL_0__1603_.vdd
rlabel metal1 4884 2162 4916 2178 0 FILL_0__1603_.gnd
rlabel metal1 4924 2162 4996 2178 0 _1603_.gnd
rlabel metal1 4924 2402 4996 2418 0 _1603_.vdd
rlabel metal2 4933 2233 4947 2247 0 _1603_.A
rlabel metal2 4953 2273 4967 2287 0 _1603_.Y
rlabel nsubstratencontact 5016 2408 5016 2408 0 FILL_1__1746_.vdd
rlabel metal1 5004 2162 5036 2178 0 FILL_1__1746_.gnd
rlabel metal1 5024 2162 5156 2178 0 _1746_.gnd
rlabel metal1 5024 2402 5156 2418 0 _1746_.vdd
rlabel metal2 5033 2253 5047 2267 0 _1746_.A
rlabel metal2 5053 2273 5067 2287 0 _1746_.B
rlabel metal2 5113 2253 5127 2267 0 _1746_.C
rlabel metal2 5093 2273 5107 2287 0 _1746_.D
rlabel metal2 5073 2253 5087 2267 0 _1746_.Y
rlabel nsubstratencontact 5156 2408 5156 2408 0 FILL_0__1745_.vdd
rlabel metal1 5144 2162 5176 2178 0 FILL_0__1745_.gnd
rlabel nsubstratencontact 5176 2408 5176 2408 0 FILL_1__1745_.vdd
rlabel metal1 5164 2162 5196 2178 0 FILL_1__1745_.gnd
rlabel metal1 5184 2162 5276 2178 0 _1745_.gnd
rlabel metal1 5184 2402 5276 2418 0 _1745_.vdd
rlabel metal2 5193 2293 5207 2307 0 _1745_.A
rlabel metal2 5233 2293 5247 2307 0 _1745_.B
rlabel metal2 5213 2273 5227 2287 0 _1745_.Y
rlabel nsubstratencontact 5296 2408 5296 2408 0 FILL_1__1692_.vdd
rlabel metal1 5284 2162 5316 2178 0 FILL_1__1692_.gnd
rlabel nsubstratencontact 5376 2408 5376 2408 0 FILL_0__1694_.vdd
rlabel metal1 5364 2162 5396 2178 0 FILL_0__1694_.gnd
rlabel nsubstratencontact 5276 2408 5276 2408 0 FILL_0__1692_.vdd
rlabel metal1 5264 2162 5296 2178 0 FILL_0__1692_.gnd
rlabel metal1 5304 2162 5376 2178 0 _1692_.gnd
rlabel metal1 5304 2402 5376 2418 0 _1692_.vdd
rlabel metal2 5313 2273 5327 2287 0 _1692_.A
rlabel metal2 5333 2253 5347 2267 0 _1692_.Y
rlabel nsubstratencontact 5396 2408 5396 2408 0 FILL_1__1694_.vdd
rlabel metal1 5384 2162 5416 2178 0 FILL_1__1694_.gnd
rlabel metal1 5404 2162 5496 2178 0 _1694_.gnd
rlabel metal1 5404 2402 5496 2418 0 _1694_.vdd
rlabel metal2 5413 2293 5427 2307 0 _1694_.A
rlabel metal2 5453 2293 5467 2307 0 _1694_.B
rlabel metal2 5433 2273 5447 2287 0 _1694_.Y
rlabel nsubstratencontact 5516 2408 5516 2408 0 FILL_1__1697_.vdd
rlabel metal1 5504 2162 5536 2178 0 FILL_1__1697_.gnd
rlabel nsubstratencontact 5496 2408 5496 2408 0 FILL_0__1697_.vdd
rlabel metal1 5484 2162 5516 2178 0 FILL_0__1697_.gnd
rlabel metal1 5524 2162 5596 2178 0 _1697_.gnd
rlabel metal1 5524 2402 5596 2418 0 _1697_.vdd
rlabel metal2 5533 2233 5547 2247 0 _1697_.A
rlabel metal2 5553 2273 5567 2287 0 _1697_.Y
rlabel metal1 5624 2162 5756 2178 0 _1729_.gnd
rlabel metal1 5624 2402 5755 2418 0 _1729_.vdd
rlabel metal2 5633 2273 5647 2287 0 _1729_.S
rlabel metal2 5653 2253 5667 2267 0 _1729_.B
rlabel metal2 5693 2273 5707 2287 0 _1729_.Y
rlabel metal2 5713 2253 5727 2267 0 _1729_.A
rlabel nsubstratencontact 5756 2408 5756 2408 0 FILL86250x32550.vdd
rlabel metal1 5744 2162 5776 2178 0 FILL86250x32550.gnd
rlabel nsubstratencontact 5776 2408 5776 2408 0 FILL86550x32550.vdd
rlabel metal1 5764 2162 5796 2178 0 FILL86550x32550.gnd
rlabel nsubstratencontact 5796 2408 5796 2408 0 FILL86850x32550.vdd
rlabel metal1 5784 2162 5816 2178 0 FILL86850x32550.gnd
rlabel nsubstratencontact 5596 2408 5596 2408 0 FILL_0__1729_.vdd
rlabel metal1 5584 2162 5616 2178 0 FILL_0__1729_.gnd
rlabel nsubstratencontact 5616 2408 5616 2408 0 FILL_1__1729_.vdd
rlabel metal1 5604 2162 5636 2178 0 FILL_1__1729_.gnd
rlabel nsubstratencontact 44 2412 44 2412 0 FILL_1__1165_.vdd
rlabel metal1 24 2642 56 2658 0 FILL_1__1165_.gnd
rlabel nsubstratencontact 136 2412 136 2412 0 FILL_1__1053_.vdd
rlabel metal1 124 2642 156 2658 0 FILL_1__1053_.gnd
rlabel nsubstratencontact 24 2412 24 2412 0 FILL_0__1165_.vdd
rlabel metal1 4 2642 36 2658 0 FILL_0__1165_.gnd
rlabel nsubstratencontact 116 2412 116 2412 0 FILL_0__1053_.vdd
rlabel metal1 104 2642 136 2658 0 FILL_0__1053_.gnd
rlabel metal1 44 2642 116 2658 0 _1165_.gnd
rlabel metal1 44 2402 116 2418 0 _1165_.vdd
rlabel metal2 93 2573 107 2587 0 _1165_.A
rlabel metal2 73 2533 87 2547 0 _1165_.Y
rlabel nsubstratencontact 244 2412 244 2412 0 FILL_1__1127_.vdd
rlabel metal1 224 2642 256 2658 0 FILL_1__1127_.gnd
rlabel nsubstratencontact 224 2412 224 2412 0 FILL_0__1127_.vdd
rlabel metal1 204 2642 236 2658 0 FILL_0__1127_.gnd
rlabel metal1 244 2642 356 2658 0 _1127_.gnd
rlabel metal1 244 2402 356 2418 0 _1127_.vdd
rlabel metal2 333 2533 347 2547 0 _1127_.A
rlabel metal2 313 2573 327 2587 0 _1127_.B
rlabel metal2 293 2533 307 2547 0 _1127_.C
rlabel metal2 273 2553 287 2567 0 _1127_.Y
rlabel metal1 144 2642 216 2658 0 _1053_.gnd
rlabel metal1 144 2402 216 2418 0 _1053_.vdd
rlabel metal2 153 2573 167 2587 0 _1053_.A
rlabel metal2 173 2533 187 2547 0 _1053_.Y
rlabel nsubstratencontact 376 2412 376 2412 0 FILL_1__1126_.vdd
rlabel metal1 364 2642 396 2658 0 FILL_1__1126_.gnd
rlabel nsubstratencontact 356 2412 356 2412 0 FILL_0__1126_.vdd
rlabel metal1 344 2642 376 2658 0 FILL_0__1126_.gnd
rlabel nsubstratencontact 496 2412 496 2412 0 FILL_0__1262_.vdd
rlabel metal1 484 2642 516 2658 0 FILL_0__1262_.gnd
rlabel metal1 384 2642 496 2658 0 _1126_.gnd
rlabel metal1 384 2402 496 2418 0 _1126_.vdd
rlabel metal2 393 2533 407 2547 0 _1126_.A
rlabel metal2 413 2513 427 2527 0 _1126_.B
rlabel metal2 433 2533 447 2547 0 _1126_.C
rlabel metal2 453 2513 467 2527 0 _1126_.Y
rlabel nsubstratencontact 516 2412 516 2412 0 FILL_1__1262_.vdd
rlabel metal1 504 2642 536 2658 0 FILL_1__1262_.gnd
rlabel nsubstratencontact 616 2412 616 2412 0 FILL_1__1591_.vdd
rlabel metal1 604 2642 636 2658 0 FILL_1__1591_.gnd
rlabel nsubstratencontact 596 2412 596 2412 0 FILL_0__1591_.vdd
rlabel metal1 584 2642 616 2658 0 FILL_0__1591_.gnd
rlabel metal1 624 2642 716 2658 0 _1591_.gnd
rlabel metal1 624 2402 716 2418 0 _1591_.vdd
rlabel metal2 673 2553 687 2567 0 _1591_.B
rlabel metal2 633 2553 647 2567 0 _1591_.A
rlabel metal2 653 2573 667 2587 0 _1591_.Y
rlabel metal1 524 2642 596 2658 0 _1262_.gnd
rlabel metal1 524 2402 596 2418 0 _1262_.vdd
rlabel metal2 533 2573 547 2587 0 _1262_.A
rlabel metal2 553 2533 567 2547 0 _1262_.Y
rlabel nsubstratencontact 736 2412 736 2412 0 FILL_1__1593_.vdd
rlabel metal1 724 2642 756 2658 0 FILL_1__1593_.gnd
rlabel nsubstratencontact 716 2412 716 2412 0 FILL_0__1593_.vdd
rlabel metal1 704 2642 736 2658 0 FILL_0__1593_.gnd
rlabel metal1 744 2642 856 2658 0 _1593_.gnd
rlabel metal1 744 2402 856 2418 0 _1593_.vdd
rlabel metal2 753 2553 767 2567 0 _1593_.A
rlabel metal2 773 2533 787 2547 0 _1593_.B
rlabel metal2 813 2533 827 2547 0 _1593_.C
rlabel metal2 793 2553 807 2567 0 _1593_.Y
rlabel nsubstratencontact 876 2412 876 2412 0 FILL_1__1592_.vdd
rlabel metal1 864 2642 896 2658 0 FILL_1__1592_.gnd
rlabel nsubstratencontact 856 2412 856 2412 0 FILL_0__1592_.vdd
rlabel metal1 844 2642 876 2658 0 FILL_0__1592_.gnd
rlabel nsubstratencontact 896 2412 896 2412 0 FILL_2__1592_.vdd
rlabel metal1 884 2642 916 2658 0 FILL_2__1592_.gnd
rlabel nsubstratencontact 1024 2412 1024 2412 0 FILL_0__1044_.vdd
rlabel metal1 1004 2642 1036 2658 0 FILL_0__1044_.gnd
rlabel metal1 904 2642 1016 2658 0 _1592_.gnd
rlabel metal1 904 2402 1016 2418 0 _1592_.vdd
rlabel metal2 913 2533 927 2547 0 _1592_.A
rlabel metal2 933 2573 947 2587 0 _1592_.B
rlabel metal2 953 2533 967 2547 0 _1592_.C
rlabel metal2 973 2553 987 2567 0 _1592_.Y
rlabel nsubstratencontact 1044 2412 1044 2412 0 FILL_1__1044_.vdd
rlabel metal1 1024 2642 1056 2658 0 FILL_1__1044_.gnd
rlabel metal1 1044 2642 1156 2658 0 _1044_.gnd
rlabel metal1 1044 2402 1156 2418 0 _1044_.vdd
rlabel metal2 1133 2553 1147 2567 0 _1044_.A
rlabel metal2 1113 2533 1127 2547 0 _1044_.B
rlabel metal2 1073 2533 1087 2547 0 _1044_.C
rlabel metal2 1093 2553 1107 2567 0 _1044_.Y
rlabel nsubstratencontact 1184 2412 1184 2412 0 FILL_1__1208_.vdd
rlabel metal1 1164 2642 1196 2658 0 FILL_1__1208_.gnd
rlabel nsubstratencontact 1164 2412 1164 2412 0 FILL_0__1208_.vdd
rlabel metal1 1144 2642 1176 2658 0 FILL_0__1208_.gnd
rlabel metal1 1184 2642 1276 2658 0 _1208_.gnd
rlabel metal1 1184 2402 1276 2418 0 _1208_.vdd
rlabel metal2 1253 2513 1267 2527 0 _1208_.A
rlabel metal2 1213 2513 1227 2527 0 _1208_.B
rlabel metal2 1233 2533 1247 2547 0 _1208_.Y
rlabel nsubstratencontact 1296 2412 1296 2412 0 FILL_1__1241_.vdd
rlabel metal1 1284 2642 1316 2658 0 FILL_1__1241_.gnd
rlabel nsubstratencontact 1276 2412 1276 2412 0 FILL_0__1241_.vdd
rlabel metal1 1264 2642 1296 2658 0 FILL_0__1241_.gnd
rlabel metal1 1304 2642 1416 2658 0 _1241_.gnd
rlabel metal1 1304 2402 1416 2418 0 _1241_.vdd
rlabel metal2 1313 2553 1327 2567 0 _1241_.A
rlabel metal2 1373 2553 1387 2567 0 _1241_.Y
rlabel metal2 1353 2513 1367 2527 0 _1241_.B
rlabel nsubstratencontact 1444 2412 1444 2412 0 FILL_1__1204_.vdd
rlabel metal1 1424 2642 1456 2658 0 FILL_1__1204_.gnd
rlabel nsubstratencontact 1424 2412 1424 2412 0 FILL_0__1204_.vdd
rlabel metal1 1404 2642 1436 2658 0 FILL_0__1204_.gnd
rlabel metal1 1444 2642 1556 2658 0 _1204_.gnd
rlabel metal1 1444 2402 1556 2418 0 _1204_.vdd
rlabel metal2 1533 2533 1547 2547 0 _1204_.A
rlabel metal2 1513 2513 1527 2527 0 _1204_.B
rlabel metal2 1493 2533 1507 2547 0 _1204_.C
rlabel metal2 1473 2513 1487 2527 0 _1204_.Y
rlabel nsubstratencontact 1576 2412 1576 2412 0 FILL_1__1199_.vdd
rlabel metal1 1564 2642 1596 2658 0 FILL_1__1199_.gnd
rlabel nsubstratencontact 1556 2412 1556 2412 0 FILL_0__1199_.vdd
rlabel metal1 1544 2642 1576 2658 0 FILL_0__1199_.gnd
rlabel metal1 1584 2642 1656 2658 0 _1199_.gnd
rlabel metal1 1584 2402 1656 2418 0 _1199_.vdd
rlabel metal2 1593 2573 1607 2587 0 _1199_.A
rlabel metal2 1613 2533 1627 2547 0 _1199_.Y
rlabel nsubstratencontact 1676 2412 1676 2412 0 FILL_1__1341_.vdd
rlabel metal1 1664 2642 1696 2658 0 FILL_1__1341_.gnd
rlabel nsubstratencontact 1656 2412 1656 2412 0 FILL_0__1341_.vdd
rlabel metal1 1644 2642 1676 2658 0 FILL_0__1341_.gnd
rlabel metal1 1684 2642 1796 2658 0 _1341_.gnd
rlabel metal1 1684 2402 1796 2418 0 _1341_.vdd
rlabel metal2 1693 2553 1707 2567 0 _1341_.A
rlabel metal2 1713 2533 1727 2547 0 _1341_.B
rlabel metal2 1753 2533 1767 2547 0 _1341_.C
rlabel metal2 1733 2553 1747 2567 0 _1341_.Y
rlabel nsubstratencontact 1824 2412 1824 2412 0 FILL_1__1203_.vdd
rlabel metal1 1804 2642 1836 2658 0 FILL_1__1203_.gnd
rlabel nsubstratencontact 1804 2412 1804 2412 0 FILL_0__1203_.vdd
rlabel metal1 1784 2642 1816 2658 0 FILL_0__1203_.gnd
rlabel metal1 1824 2642 1936 2658 0 _1203_.gnd
rlabel metal1 1824 2402 1936 2418 0 _1203_.vdd
rlabel metal2 1913 2553 1927 2567 0 _1203_.A
rlabel metal2 1893 2533 1907 2547 0 _1203_.B
rlabel metal2 1853 2533 1867 2547 0 _1203_.C
rlabel metal2 1873 2553 1887 2567 0 _1203_.Y
rlabel nsubstratencontact 1956 2412 1956 2412 0 FILL_1__1571_.vdd
rlabel metal1 1944 2642 1976 2658 0 FILL_1__1571_.gnd
rlabel nsubstratencontact 1936 2412 1936 2412 0 FILL_0__1571_.vdd
rlabel metal1 1924 2642 1956 2658 0 FILL_0__1571_.gnd
rlabel metal1 1964 2642 2076 2658 0 _1571_.gnd
rlabel metal1 1964 2402 2076 2418 0 _1571_.vdd
rlabel metal2 1973 2553 1987 2567 0 _1571_.A
rlabel metal2 1993 2533 2007 2547 0 _1571_.B
rlabel metal2 2033 2533 2047 2547 0 _1571_.C
rlabel metal2 2013 2553 2027 2567 0 _1571_.Y
rlabel nsubstratencontact 2104 2412 2104 2412 0 FILL_1__1230_.vdd
rlabel metal1 2084 2642 2116 2658 0 FILL_1__1230_.gnd
rlabel nsubstratencontact 2084 2412 2084 2412 0 FILL_0__1230_.vdd
rlabel metal1 2064 2642 2096 2658 0 FILL_0__1230_.gnd
rlabel metal1 2104 2642 2216 2658 0 _1230_.gnd
rlabel metal1 2104 2402 2216 2418 0 _1230_.vdd
rlabel metal2 2193 2533 2207 2547 0 _1230_.A
rlabel metal2 2173 2513 2187 2527 0 _1230_.B
rlabel metal2 2153 2533 2167 2547 0 _1230_.C
rlabel metal2 2133 2513 2147 2527 0 _1230_.Y
rlabel nsubstratencontact 2244 2412 2244 2412 0 FILL_1__1238_.vdd
rlabel metal1 2224 2642 2256 2658 0 FILL_1__1238_.gnd
rlabel nsubstratencontact 2224 2412 2224 2412 0 FILL_0__1238_.vdd
rlabel metal1 2204 2642 2236 2658 0 FILL_0__1238_.gnd
rlabel metal1 2244 2642 2356 2658 0 _1238_.gnd
rlabel metal1 2244 2402 2356 2418 0 _1238_.vdd
rlabel metal2 2333 2533 2347 2547 0 _1238_.A
rlabel metal2 2313 2573 2327 2587 0 _1238_.B
rlabel metal2 2293 2533 2307 2547 0 _1238_.C
rlabel metal2 2273 2553 2287 2567 0 _1238_.Y
rlabel nsubstratencontact 2376 2412 2376 2412 0 FILL_1__1227_.vdd
rlabel metal1 2364 2642 2396 2658 0 FILL_1__1227_.gnd
rlabel nsubstratencontact 2356 2412 2356 2412 0 FILL_0__1227_.vdd
rlabel metal1 2344 2642 2376 2658 0 FILL_0__1227_.gnd
rlabel metal1 2384 2642 2476 2658 0 _1227_.gnd
rlabel metal1 2384 2402 2476 2418 0 _1227_.vdd
rlabel metal2 2393 2513 2407 2527 0 _1227_.A
rlabel metal2 2433 2513 2447 2527 0 _1227_.B
rlabel metal2 2413 2533 2427 2547 0 _1227_.Y
rlabel nsubstratencontact 2524 2412 2524 2412 0 FILL_2__1233_.vdd
rlabel metal1 2504 2642 2536 2658 0 FILL_2__1233_.gnd
rlabel nsubstratencontact 2504 2412 2504 2412 0 FILL_1__1233_.vdd
rlabel metal1 2484 2642 2516 2658 0 FILL_1__1233_.gnd
rlabel nsubstratencontact 2484 2412 2484 2412 0 FILL_0__1233_.vdd
rlabel metal1 2464 2642 2496 2658 0 FILL_0__1233_.gnd
rlabel metal1 2524 2642 2636 2658 0 _1233_.gnd
rlabel metal1 2524 2402 2636 2418 0 _1233_.vdd
rlabel metal2 2613 2553 2627 2567 0 _1233_.A
rlabel metal2 2593 2533 2607 2547 0 _1233_.B
rlabel metal2 2553 2533 2567 2547 0 _1233_.C
rlabel metal2 2573 2553 2587 2567 0 _1233_.Y
rlabel nsubstratencontact 2656 2412 2656 2412 0 FILL_1__1229_.vdd
rlabel metal1 2644 2642 2676 2658 0 FILL_1__1229_.gnd
rlabel nsubstratencontact 2636 2412 2636 2412 0 FILL_0__1229_.vdd
rlabel metal1 2624 2642 2656 2658 0 FILL_0__1229_.gnd
rlabel nsubstratencontact 2784 2412 2784 2412 0 FILL_0__1482_.vdd
rlabel metal1 2764 2642 2796 2658 0 FILL_0__1482_.gnd
rlabel metal1 2664 2642 2776 2658 0 _1229_.gnd
rlabel metal1 2664 2402 2776 2418 0 _1229_.vdd
rlabel metal2 2673 2553 2687 2567 0 _1229_.A
rlabel metal2 2693 2533 2707 2547 0 _1229_.B
rlabel metal2 2733 2533 2747 2547 0 _1229_.C
rlabel metal2 2713 2553 2727 2567 0 _1229_.Y
rlabel nsubstratencontact 2804 2412 2804 2412 0 FILL_1__1482_.vdd
rlabel metal1 2784 2642 2816 2658 0 FILL_1__1482_.gnd
rlabel metal1 2804 2642 2916 2658 0 _1482_.gnd
rlabel metal1 2804 2402 2916 2418 0 _1482_.vdd
rlabel metal2 2893 2533 2907 2547 0 _1482_.A
rlabel metal2 2873 2573 2887 2587 0 _1482_.B
rlabel metal2 2853 2533 2867 2547 0 _1482_.C
rlabel metal2 2833 2553 2847 2567 0 _1482_.Y
rlabel nsubstratencontact 3036 2412 3036 2412 0 FILL_1__1542_.vdd
rlabel metal1 3024 2642 3056 2658 0 FILL_1__1542_.gnd
rlabel nsubstratencontact 2944 2412 2944 2412 0 FILL_1__1179_.vdd
rlabel metal1 2924 2642 2956 2658 0 FILL_1__1179_.gnd
rlabel nsubstratencontact 3016 2412 3016 2412 0 FILL_0__1542_.vdd
rlabel metal1 3004 2642 3036 2658 0 FILL_0__1542_.gnd
rlabel nsubstratencontact 2924 2412 2924 2412 0 FILL_0__1179_.vdd
rlabel metal1 2904 2642 2936 2658 0 FILL_0__1179_.gnd
rlabel metal1 2944 2642 3016 2658 0 _1179_.gnd
rlabel metal1 2944 2402 3016 2418 0 _1179_.vdd
rlabel metal2 2993 2573 3007 2587 0 _1179_.A
rlabel metal2 2973 2533 2987 2547 0 _1179_.Y
rlabel nsubstratencontact 3156 2412 3156 2412 0 FILL_0__1566_.vdd
rlabel metal1 3144 2642 3176 2658 0 FILL_0__1566_.gnd
rlabel metal1 3044 2642 3156 2658 0 _1542_.gnd
rlabel metal1 3044 2402 3156 2418 0 _1542_.vdd
rlabel metal2 3053 2553 3067 2567 0 _1542_.A
rlabel metal2 3073 2533 3087 2547 0 _1542_.B
rlabel metal2 3113 2533 3127 2547 0 _1542_.C
rlabel metal2 3093 2553 3107 2567 0 _1542_.Y
rlabel nsubstratencontact 3196 2412 3196 2412 0 FILL_2__1566_.vdd
rlabel metal1 3184 2642 3216 2658 0 FILL_2__1566_.gnd
rlabel nsubstratencontact 3176 2412 3176 2412 0 FILL_1__1566_.vdd
rlabel metal1 3164 2642 3196 2658 0 FILL_1__1566_.gnd
rlabel metal1 3204 2642 3296 2658 0 _1566_.gnd
rlabel metal1 3204 2402 3296 2418 0 _1566_.vdd
rlabel metal2 3213 2513 3227 2527 0 _1566_.A
rlabel metal2 3253 2513 3267 2527 0 _1566_.B
rlabel metal2 3233 2533 3247 2547 0 _1566_.Y
rlabel nsubstratencontact 3324 2412 3324 2412 0 FILL_1__1178_.vdd
rlabel metal1 3304 2642 3336 2658 0 FILL_1__1178_.gnd
rlabel nsubstratencontact 3304 2412 3304 2412 0 FILL_0__1178_.vdd
rlabel metal1 3284 2642 3316 2658 0 FILL_0__1178_.gnd
rlabel metal1 3324 2642 3436 2658 0 _1178_.gnd
rlabel metal1 3324 2402 3436 2418 0 _1178_.vdd
rlabel metal2 3413 2533 3427 2547 0 _1178_.A
rlabel metal2 3393 2513 3407 2527 0 _1178_.B
rlabel metal2 3373 2533 3387 2547 0 _1178_.C
rlabel metal2 3353 2513 3367 2527 0 _1178_.Y
rlabel nsubstratencontact 3456 2412 3456 2412 0 FILL_1__1427_.vdd
rlabel metal1 3444 2642 3476 2658 0 FILL_1__1427_.gnd
rlabel nsubstratencontact 3436 2412 3436 2412 0 FILL_0__1427_.vdd
rlabel metal1 3424 2642 3456 2658 0 FILL_0__1427_.gnd
rlabel metal1 3464 2642 3576 2658 0 _1427_.gnd
rlabel metal1 3464 2402 3576 2418 0 _1427_.vdd
rlabel metal2 3473 2553 3487 2567 0 _1427_.A
rlabel metal2 3533 2553 3547 2567 0 _1427_.Y
rlabel metal2 3513 2513 3527 2527 0 _1427_.B
rlabel nsubstratencontact 3716 2412 3716 2412 0 FILL_1__1595_.vdd
rlabel metal1 3704 2642 3736 2658 0 FILL_1__1595_.gnd
rlabel nsubstratencontact 3596 2412 3596 2412 0 FILL_1__1173_.vdd
rlabel metal1 3584 2642 3616 2658 0 FILL_1__1173_.gnd
rlabel nsubstratencontact 3696 2412 3696 2412 0 FILL_0__1595_.vdd
rlabel metal1 3684 2642 3716 2658 0 FILL_0__1595_.gnd
rlabel nsubstratencontact 3576 2412 3576 2412 0 FILL_0__1173_.vdd
rlabel metal1 3564 2642 3596 2658 0 FILL_0__1173_.gnd
rlabel metal1 3724 2642 3856 2658 0 _1595_.gnd
rlabel metal1 3724 2402 3856 2418 0 _1595_.vdd
rlabel metal2 3733 2553 3747 2567 0 _1595_.A
rlabel metal2 3753 2533 3767 2547 0 _1595_.B
rlabel metal2 3813 2553 3827 2567 0 _1595_.C
rlabel metal2 3793 2533 3807 2547 0 _1595_.D
rlabel metal2 3773 2553 3787 2567 0 _1595_.Y
rlabel metal1 3604 2642 3696 2658 0 _1173_.gnd
rlabel metal1 3604 2402 3696 2418 0 _1173_.vdd
rlabel metal2 3613 2513 3627 2527 0 _1173_.A
rlabel metal2 3653 2513 3667 2527 0 _1173_.B
rlabel metal2 3633 2533 3647 2547 0 _1173_.Y
rlabel nsubstratencontact 3876 2412 3876 2412 0 FILL_1__1590_.vdd
rlabel metal1 3864 2642 3896 2658 0 FILL_1__1590_.gnd
rlabel nsubstratencontact 3856 2412 3856 2412 0 FILL_0__1590_.vdd
rlabel metal1 3844 2642 3876 2658 0 FILL_0__1590_.gnd
rlabel metal1 3884 2642 3976 2658 0 _1590_.gnd
rlabel metal1 3884 2402 3976 2418 0 _1590_.vdd
rlabel metal2 3933 2553 3947 2567 0 _1590_.B
rlabel metal2 3893 2553 3907 2567 0 _1590_.A
rlabel metal2 3913 2573 3927 2587 0 _1590_.Y
rlabel metal1 3964 2642 4456 2658 0 _1668_.gnd
rlabel metal1 3964 2402 4456 2418 0 _1668_.vdd
rlabel metal2 4373 2533 4387 2547 0 _1668_.S
rlabel metal2 4253 2573 4267 2587 0 _1668_.D
rlabel metal2 4073 2533 4087 2547 0 _1668_.CLK
rlabel metal2 4413 2513 4427 2527 0 _1668_.R
rlabel metal2 3993 2533 4007 2547 0 _1668_.Q
rlabel metal1 4444 2642 4936 2658 0 _1666_.gnd
rlabel metal1 4444 2402 4936 2418 0 _1666_.vdd
rlabel metal2 4513 2533 4527 2547 0 _1666_.S
rlabel metal2 4633 2573 4647 2587 0 _1666_.D
rlabel metal2 4813 2533 4827 2547 0 _1666_.CLK
rlabel metal2 4473 2513 4487 2527 0 _1666_.R
rlabel metal2 4893 2533 4907 2547 0 _1666_.Q
rlabel metal1 4924 2642 5176 2658 0 _1655_.gnd
rlabel metal1 4924 2402 5176 2418 0 _1655_.vdd
rlabel metal2 5013 2553 5027 2567 0 _1655_.D
rlabel metal2 5053 2553 5067 2567 0 _1655_.CLK
rlabel metal2 5133 2553 5147 2567 0 _1655_.Q
rlabel metal1 5204 2642 5416 2658 0 CLKBUF1_insert0.gnd
rlabel metal1 5204 2402 5416 2418 0 CLKBUF1_insert0.vdd
rlabel metal2 5373 2533 5387 2547 0 CLKBUF1_insert0.A
rlabel metal2 5233 2533 5247 2547 0 CLKBUF1_insert0.Y
rlabel metal1 5464 2642 5676 2658 0 CLKBUF1_insert1.gnd
rlabel metal1 5464 2402 5676 2418 0 CLKBUF1_insert1.vdd
rlabel metal2 5493 2533 5507 2547 0 CLKBUF1_insert1.A
rlabel metal2 5633 2533 5647 2547 0 CLKBUF1_insert1.Y
rlabel nsubstratencontact 5184 2412 5184 2412 0 FILL_0_CLKBUF1_insert0.vdd
rlabel metal1 5164 2642 5196 2658 0 FILL_0_CLKBUF1_insert0.gnd
rlabel nsubstratencontact 5416 2412 5416 2412 0 FILL_0_CLKBUF1_insert1.vdd
rlabel metal1 5404 2642 5436 2658 0 FILL_0_CLKBUF1_insert1.gnd
rlabel nsubstratencontact 5204 2412 5204 2412 0 FILL_1_CLKBUF1_insert0.vdd
rlabel metal1 5184 2642 5216 2658 0 FILL_1_CLKBUF1_insert0.gnd
rlabel nsubstratencontact 5436 2412 5436 2412 0 FILL_1_CLKBUF1_insert1.vdd
rlabel metal1 5424 2642 5456 2658 0 FILL_1_CLKBUF1_insert1.gnd
rlabel nsubstratencontact 5456 2412 5456 2412 0 FILL_2_CLKBUF1_insert1.vdd
rlabel metal1 5444 2642 5476 2658 0 FILL_2_CLKBUF1_insert1.gnd
rlabel metal1 5704 2642 5776 2658 0 _1690_.gnd
rlabel metal1 5704 2402 5776 2418 0 _1690_.vdd
rlabel metal2 5713 2533 5727 2547 0 _1690_.A
rlabel metal2 5733 2553 5747 2567 0 _1690_.Y
rlabel nsubstratencontact 5784 2412 5784 2412 0 FILL86550x36150.vdd
rlabel metal1 5764 2642 5796 2658 0 FILL86550x36150.gnd
rlabel nsubstratencontact 5804 2412 5804 2412 0 FILL86850x36150.vdd
rlabel metal1 5784 2642 5816 2658 0 FILL86850x36150.gnd
rlabel nsubstratencontact 5676 2412 5676 2412 0 FILL_0__1690_.vdd
rlabel metal1 5664 2642 5696 2658 0 FILL_0__1690_.gnd
rlabel nsubstratencontact 5696 2412 5696 2412 0 FILL_1__1690_.vdd
rlabel metal1 5684 2642 5716 2658 0 FILL_1__1690_.gnd
rlabel nsubstratencontact 44 2888 44 2888 0 FILL_1__1052_.vdd
rlabel metal1 24 2642 56 2658 0 FILL_1__1052_.gnd
rlabel nsubstratencontact 136 2888 136 2888 0 FILL_0__1191_.vdd
rlabel metal1 124 2642 156 2658 0 FILL_0__1191_.gnd
rlabel nsubstratencontact 24 2888 24 2888 0 FILL_0__1052_.vdd
rlabel metal1 4 2642 36 2658 0 FILL_0__1052_.gnd
rlabel metal1 44 2642 136 2658 0 _1052_.gnd
rlabel metal1 44 2882 136 2898 0 _1052_.vdd
rlabel metal2 113 2773 127 2787 0 _1052_.A
rlabel metal2 73 2773 87 2787 0 _1052_.B
rlabel metal2 93 2753 107 2767 0 _1052_.Y
rlabel nsubstratencontact 156 2888 156 2888 0 FILL_1__1191_.vdd
rlabel metal1 144 2642 176 2658 0 FILL_1__1191_.gnd
rlabel metal1 164 2642 276 2658 0 _1191_.gnd
rlabel metal1 164 2882 276 2898 0 _1191_.vdd
rlabel metal2 173 2733 187 2747 0 _1191_.A
rlabel metal2 193 2753 207 2767 0 _1191_.B
rlabel metal2 233 2753 247 2767 0 _1191_.C
rlabel metal2 213 2733 227 2747 0 _1191_.Y
rlabel nsubstratencontact 304 2888 304 2888 0 FILL_1__1263_.vdd
rlabel metal1 284 2642 316 2658 0 FILL_1__1263_.gnd
rlabel nsubstratencontact 376 2888 376 2888 0 FILL_0__1267_.vdd
rlabel metal1 364 2642 396 2658 0 FILL_0__1267_.gnd
rlabel nsubstratencontact 284 2888 284 2888 0 FILL_0__1263_.vdd
rlabel metal1 264 2642 296 2658 0 FILL_0__1263_.gnd
rlabel metal1 304 2642 376 2658 0 _1263_.gnd
rlabel metal1 304 2882 376 2898 0 _1263_.vdd
rlabel metal2 353 2713 367 2727 0 _1263_.A
rlabel metal2 333 2753 347 2767 0 _1263_.Y
rlabel nsubstratencontact 396 2888 396 2888 0 FILL_1__1267_.vdd
rlabel metal1 384 2642 416 2658 0 FILL_1__1267_.gnd
rlabel metal1 404 2642 516 2658 0 _1267_.gnd
rlabel metal1 404 2882 516 2898 0 _1267_.vdd
rlabel metal2 413 2753 427 2767 0 _1267_.A
rlabel metal2 433 2713 447 2727 0 _1267_.B
rlabel metal2 453 2753 467 2767 0 _1267_.C
rlabel metal2 473 2733 487 2747 0 _1267_.Y
rlabel nsubstratencontact 524 2888 524 2888 0 FILL_0__1268_.vdd
rlabel metal1 504 2642 536 2658 0 FILL_0__1268_.gnd
rlabel nsubstratencontact 544 2888 544 2888 0 FILL_1__1268_.vdd
rlabel metal1 524 2642 556 2658 0 FILL_1__1268_.gnd
rlabel nsubstratencontact 636 2888 636 2888 0 FILL_0__1260_.vdd
rlabel metal1 624 2642 656 2658 0 FILL_0__1260_.gnd
rlabel metal1 544 2642 636 2658 0 _1268_.gnd
rlabel metal1 544 2882 636 2898 0 _1268_.vdd
rlabel metal2 613 2773 627 2787 0 _1268_.A
rlabel metal2 573 2773 587 2787 0 _1268_.B
rlabel metal2 593 2753 607 2767 0 _1268_.Y
rlabel nsubstratencontact 656 2888 656 2888 0 FILL_1__1260_.vdd
rlabel metal1 644 2642 676 2658 0 FILL_1__1260_.gnd
rlabel metal1 664 2642 776 2658 0 _1260_.gnd
rlabel metal1 664 2882 776 2898 0 _1260_.vdd
rlabel metal2 673 2733 687 2747 0 _1260_.A
rlabel metal2 733 2733 747 2747 0 _1260_.Y
rlabel metal2 713 2773 727 2787 0 _1260_.B
rlabel nsubstratencontact 796 2888 796 2888 0 FILL_1__1261_.vdd
rlabel metal1 784 2642 816 2658 0 FILL_1__1261_.gnd
rlabel nsubstratencontact 776 2888 776 2888 0 FILL_0__1261_.vdd
rlabel metal1 764 2642 796 2658 0 FILL_0__1261_.gnd
rlabel metal1 804 2642 896 2658 0 _1261_.gnd
rlabel metal1 804 2882 896 2898 0 _1261_.vdd
rlabel metal2 813 2773 827 2787 0 _1261_.A
rlabel metal2 853 2773 867 2787 0 _1261_.B
rlabel metal2 833 2753 847 2767 0 _1261_.Y
rlabel nsubstratencontact 916 2888 916 2888 0 FILL_1__1358_.vdd
rlabel metal1 904 2642 936 2658 0 FILL_1__1358_.gnd
rlabel nsubstratencontact 896 2888 896 2888 0 FILL_0__1358_.vdd
rlabel metal1 884 2642 916 2658 0 FILL_0__1358_.gnd
rlabel metal1 924 2642 1036 2658 0 _1358_.gnd
rlabel metal1 924 2882 1036 2898 0 _1358_.vdd
rlabel metal2 933 2753 947 2767 0 _1358_.A
rlabel metal2 953 2713 967 2727 0 _1358_.B
rlabel metal2 973 2753 987 2767 0 _1358_.C
rlabel metal2 993 2733 1007 2747 0 _1358_.Y
rlabel nsubstratencontact 1056 2888 1056 2888 0 FILL_1__1270_.vdd
rlabel metal1 1044 2642 1076 2658 0 FILL_1__1270_.gnd
rlabel nsubstratencontact 1036 2888 1036 2888 0 FILL_0__1270_.vdd
rlabel metal1 1024 2642 1056 2658 0 FILL_0__1270_.gnd
rlabel metal1 1064 2642 1156 2658 0 _1270_.gnd
rlabel metal1 1064 2882 1156 2898 0 _1270_.vdd
rlabel metal2 1073 2773 1087 2787 0 _1270_.A
rlabel metal2 1113 2773 1127 2787 0 _1270_.B
rlabel metal2 1093 2753 1107 2767 0 _1270_.Y
rlabel nsubstratencontact 1204 2888 1204 2888 0 FILL_2__1207_.vdd
rlabel metal1 1184 2642 1216 2658 0 FILL_2__1207_.gnd
rlabel nsubstratencontact 1184 2888 1184 2888 0 FILL_1__1207_.vdd
rlabel metal1 1164 2642 1196 2658 0 FILL_1__1207_.gnd
rlabel nsubstratencontact 1164 2888 1164 2888 0 FILL_0__1207_.vdd
rlabel metal1 1144 2642 1176 2658 0 FILL_0__1207_.gnd
rlabel metal1 1204 2642 1316 2658 0 _1207_.gnd
rlabel metal1 1204 2882 1316 2898 0 _1207_.vdd
rlabel metal2 1293 2733 1307 2747 0 _1207_.A
rlabel metal2 1273 2753 1287 2767 0 _1207_.B
rlabel metal2 1233 2753 1247 2767 0 _1207_.C
rlabel metal2 1253 2733 1267 2747 0 _1207_.Y
rlabel nsubstratencontact 1336 2888 1336 2888 0 FILL_1__1287_.vdd
rlabel metal1 1324 2642 1356 2658 0 FILL_1__1287_.gnd
rlabel nsubstratencontact 1316 2888 1316 2888 0 FILL_0__1287_.vdd
rlabel metal1 1304 2642 1336 2658 0 FILL_0__1287_.gnd
rlabel metal1 1344 2642 1456 2658 0 _1287_.gnd
rlabel metal1 1344 2882 1456 2898 0 _1287_.vdd
rlabel metal2 1353 2733 1367 2747 0 _1287_.A
rlabel metal2 1373 2753 1387 2767 0 _1287_.B
rlabel metal2 1413 2753 1427 2767 0 _1287_.C
rlabel metal2 1393 2733 1407 2747 0 _1287_.Y
rlabel nsubstratencontact 1484 2888 1484 2888 0 FILL_1__1202_.vdd
rlabel metal1 1464 2642 1496 2658 0 FILL_1__1202_.gnd
rlabel nsubstratencontact 1464 2888 1464 2888 0 FILL_0__1202_.vdd
rlabel metal1 1444 2642 1476 2658 0 FILL_0__1202_.gnd
rlabel metal1 1484 2642 1596 2658 0 _1202_.gnd
rlabel metal1 1484 2882 1596 2898 0 _1202_.vdd
rlabel metal2 1573 2713 1587 2727 0 _1202_.A
rlabel metal2 1553 2733 1567 2747 0 _1202_.B
rlabel metal2 1513 2753 1527 2767 0 _1202_.Y
rlabel nsubstratencontact 1616 2888 1616 2888 0 FILL_1__1205_.vdd
rlabel metal1 1604 2642 1636 2658 0 FILL_1__1205_.gnd
rlabel nsubstratencontact 1596 2888 1596 2888 0 FILL_0__1205_.vdd
rlabel metal1 1584 2642 1616 2658 0 FILL_0__1205_.gnd
rlabel metal1 1624 2642 1716 2658 0 _1205_.gnd
rlabel metal1 1624 2882 1716 2898 0 _1205_.vdd
rlabel metal2 1673 2733 1687 2747 0 _1205_.B
rlabel metal2 1633 2733 1647 2747 0 _1205_.A
rlabel metal2 1653 2713 1667 2727 0 _1205_.Y
rlabel nsubstratencontact 1744 2888 1744 2888 0 FILL_1__1206_.vdd
rlabel metal1 1724 2642 1756 2658 0 FILL_1__1206_.gnd
rlabel nsubstratencontact 1724 2888 1724 2888 0 FILL_0__1206_.vdd
rlabel metal1 1704 2642 1736 2658 0 FILL_0__1206_.gnd
rlabel metal1 1744 2642 1856 2658 0 _1206_.gnd
rlabel metal1 1744 2882 1856 2898 0 _1206_.vdd
rlabel metal2 1833 2733 1847 2747 0 _1206_.A
rlabel metal2 1773 2733 1787 2747 0 _1206_.Y
rlabel metal2 1793 2773 1807 2787 0 _1206_.B
rlabel nsubstratencontact 1904 2888 1904 2888 0 FILL_2__1200_.vdd
rlabel metal1 1884 2642 1916 2658 0 FILL_2__1200_.gnd
rlabel nsubstratencontact 1884 2888 1884 2888 0 FILL_1__1200_.vdd
rlabel metal1 1864 2642 1896 2658 0 FILL_1__1200_.gnd
rlabel nsubstratencontact 1864 2888 1864 2888 0 FILL_0__1200_.vdd
rlabel metal1 1844 2642 1876 2658 0 FILL_0__1200_.gnd
rlabel nsubstratencontact 2016 2888 2016 2888 0 FILL_1__1362_.vdd
rlabel metal1 2004 2642 2036 2658 0 FILL_1__1362_.gnd
rlabel nsubstratencontact 1996 2888 1996 2888 0 FILL_0__1362_.vdd
rlabel metal1 1984 2642 2016 2658 0 FILL_0__1362_.gnd
rlabel metal1 1904 2642 1996 2658 0 _1200_.gnd
rlabel metal1 1904 2882 1996 2898 0 _1200_.vdd
rlabel metal2 1973 2773 1987 2787 0 _1200_.A
rlabel metal2 1933 2773 1947 2787 0 _1200_.B
rlabel metal2 1953 2753 1967 2767 0 _1200_.Y
rlabel nsubstratencontact 2164 2888 2164 2888 0 FILL_1__1333_.vdd
rlabel metal1 2144 2642 2176 2658 0 FILL_1__1333_.gnd
rlabel nsubstratencontact 2144 2888 2144 2888 0 FILL_0__1333_.vdd
rlabel metal1 2124 2642 2156 2658 0 FILL_0__1333_.gnd
rlabel metal1 2024 2642 2136 2658 0 _1362_.gnd
rlabel metal1 2024 2882 2136 2898 0 _1362_.vdd
rlabel metal2 2033 2733 2047 2747 0 _1362_.A
rlabel metal2 2053 2753 2067 2767 0 _1362_.B
rlabel metal2 2093 2753 2107 2767 0 _1362_.C
rlabel metal2 2073 2733 2087 2747 0 _1362_.Y
rlabel nsubstratencontact 2284 2888 2284 2888 0 FILL_0__1232_.vdd
rlabel metal1 2264 2642 2296 2658 0 FILL_0__1232_.gnd
rlabel metal1 2164 2642 2276 2658 0 _1333_.gnd
rlabel metal1 2164 2882 2276 2898 0 _1333_.vdd
rlabel metal2 2253 2733 2267 2747 0 _1333_.A
rlabel metal2 2193 2733 2207 2747 0 _1333_.Y
rlabel metal2 2213 2773 2227 2787 0 _1333_.B
rlabel nsubstratencontact 2304 2888 2304 2888 0 FILL_1__1232_.vdd
rlabel metal1 2284 2642 2316 2658 0 FILL_1__1232_.gnd
rlabel nsubstratencontact 2396 2888 2396 2888 0 FILL_0__1226_.vdd
rlabel metal1 2384 2642 2416 2658 0 FILL_0__1226_.gnd
rlabel metal1 2304 2642 2396 2658 0 _1232_.gnd
rlabel metal1 2304 2882 2396 2898 0 _1232_.vdd
rlabel metal2 2373 2773 2387 2787 0 _1232_.A
rlabel metal2 2333 2773 2347 2787 0 _1232_.B
rlabel metal2 2353 2753 2367 2767 0 _1232_.Y
rlabel nsubstratencontact 2436 2888 2436 2888 0 FILL_2__1226_.vdd
rlabel metal1 2424 2642 2456 2658 0 FILL_2__1226_.gnd
rlabel nsubstratencontact 2416 2888 2416 2888 0 FILL_1__1226_.vdd
rlabel metal1 2404 2642 2436 2658 0 FILL_1__1226_.gnd
rlabel metal1 2444 2642 2536 2658 0 _1226_.gnd
rlabel metal1 2444 2882 2536 2898 0 _1226_.vdd
rlabel metal2 2493 2733 2507 2747 0 _1226_.B
rlabel metal2 2453 2733 2467 2747 0 _1226_.A
rlabel metal2 2473 2713 2487 2727 0 _1226_.Y
rlabel nsubstratencontact 2544 2888 2544 2888 0 FILL_0__1234_.vdd
rlabel metal1 2524 2642 2556 2658 0 FILL_0__1234_.gnd
rlabel nsubstratencontact 2564 2888 2564 2888 0 FILL_1__1234_.vdd
rlabel metal1 2544 2642 2576 2658 0 FILL_1__1234_.gnd
rlabel metal1 2564 2642 2676 2658 0 _1234_.gnd
rlabel metal1 2564 2882 2676 2898 0 _1234_.vdd
rlabel metal2 2653 2753 2667 2767 0 _1234_.A
rlabel metal2 2633 2773 2647 2787 0 _1234_.B
rlabel metal2 2613 2753 2627 2767 0 _1234_.C
rlabel metal2 2593 2773 2607 2787 0 _1234_.Y
rlabel nsubstratencontact 2704 2888 2704 2888 0 FILL_1__1225_.vdd
rlabel metal1 2684 2642 2716 2658 0 FILL_1__1225_.gnd
rlabel nsubstratencontact 2684 2888 2684 2888 0 FILL_0__1225_.vdd
rlabel metal1 2664 2642 2696 2658 0 FILL_0__1225_.gnd
rlabel metal1 2704 2642 2816 2658 0 _1225_.gnd
rlabel metal1 2704 2882 2816 2898 0 _1225_.vdd
rlabel metal2 2793 2733 2807 2747 0 _1225_.A
rlabel metal2 2733 2733 2747 2747 0 _1225_.Y
rlabel metal2 2753 2773 2767 2787 0 _1225_.B
rlabel nsubstratencontact 2856 2888 2856 2888 0 FILL_2__1481_.vdd
rlabel metal1 2844 2642 2876 2658 0 FILL_2__1481_.gnd
rlabel nsubstratencontact 2836 2888 2836 2888 0 FILL_1__1481_.vdd
rlabel metal1 2824 2642 2856 2658 0 FILL_1__1481_.gnd
rlabel nsubstratencontact 2816 2888 2816 2888 0 FILL_0__1481_.vdd
rlabel metal1 2804 2642 2836 2658 0 FILL_0__1481_.gnd
rlabel metal1 2864 2642 2976 2658 0 _1481_.gnd
rlabel metal1 2864 2882 2976 2898 0 _1481_.vdd
rlabel metal2 2873 2733 2887 2747 0 _1481_.A
rlabel metal2 2893 2753 2907 2767 0 _1481_.B
rlabel metal2 2933 2753 2947 2767 0 _1481_.C
rlabel metal2 2913 2733 2927 2747 0 _1481_.Y
rlabel nsubstratencontact 3004 2888 3004 2888 0 FILL_1__1223_.vdd
rlabel metal1 2984 2642 3016 2658 0 FILL_1__1223_.gnd
rlabel nsubstratencontact 2984 2888 2984 2888 0 FILL_0__1223_.vdd
rlabel metal1 2964 2642 2996 2658 0 FILL_0__1223_.gnd
rlabel metal1 3004 2642 3116 2658 0 _1223_.gnd
rlabel metal1 3004 2882 3116 2898 0 _1223_.vdd
rlabel metal2 3093 2753 3107 2767 0 _1223_.A
rlabel metal2 3073 2773 3087 2787 0 _1223_.B
rlabel metal2 3053 2753 3067 2767 0 _1223_.C
rlabel metal2 3033 2773 3047 2787 0 _1223_.Y
rlabel nsubstratencontact 3136 2888 3136 2888 0 FILL_1__1283_.vdd
rlabel metal1 3124 2642 3156 2658 0 FILL_1__1283_.gnd
rlabel nsubstratencontact 3116 2888 3116 2888 0 FILL_0__1283_.vdd
rlabel metal1 3104 2642 3136 2658 0 FILL_0__1283_.gnd
rlabel metal1 3144 2642 3236 2658 0 _1283_.gnd
rlabel metal1 3144 2882 3236 2898 0 _1283_.vdd
rlabel metal2 3153 2773 3167 2787 0 _1283_.A
rlabel metal2 3193 2773 3207 2787 0 _1283_.B
rlabel metal2 3173 2753 3187 2767 0 _1283_.Y
rlabel nsubstratencontact 3264 2888 3264 2888 0 FILL_1__1280_.vdd
rlabel metal1 3244 2642 3276 2658 0 FILL_1__1280_.gnd
rlabel nsubstratencontact 3244 2888 3244 2888 0 FILL_0__1280_.vdd
rlabel metal1 3224 2642 3256 2658 0 FILL_0__1280_.gnd
rlabel metal1 3264 2642 3376 2658 0 _1280_.gnd
rlabel metal1 3264 2882 3376 2898 0 _1280_.vdd
rlabel metal2 3353 2733 3367 2747 0 _1280_.A
rlabel metal2 3333 2753 3347 2767 0 _1280_.B
rlabel metal2 3293 2753 3307 2767 0 _1280_.C
rlabel metal2 3313 2733 3327 2747 0 _1280_.Y
rlabel nsubstratencontact 3404 2888 3404 2888 0 FILL_1__1279_.vdd
rlabel metal1 3384 2642 3416 2658 0 FILL_1__1279_.gnd
rlabel nsubstratencontact 3384 2888 3384 2888 0 FILL_0__1279_.vdd
rlabel metal1 3364 2642 3396 2658 0 FILL_0__1279_.gnd
rlabel metal1 3404 2642 3516 2658 0 _1279_.gnd
rlabel metal1 3404 2882 3516 2898 0 _1279_.vdd
rlabel metal2 3493 2733 3507 2747 0 _1279_.A
rlabel metal2 3433 2733 3447 2747 0 _1279_.Y
rlabel metal2 3453 2773 3467 2787 0 _1279_.B
rlabel nsubstratencontact 3536 2888 3536 2888 0 FILL_1__1175_.vdd
rlabel metal1 3524 2642 3556 2658 0 FILL_1__1175_.gnd
rlabel nsubstratencontact 3516 2888 3516 2888 0 FILL_0__1175_.vdd
rlabel metal1 3504 2642 3536 2658 0 FILL_0__1175_.gnd
rlabel nsubstratencontact 3656 2888 3656 2888 0 FILL_1__1587_.vdd
rlabel metal1 3644 2642 3676 2658 0 FILL_1__1587_.gnd
rlabel nsubstratencontact 3636 2888 3636 2888 0 FILL_0__1587_.vdd
rlabel metal1 3624 2642 3656 2658 0 FILL_0__1587_.gnd
rlabel metal1 3544 2642 3636 2658 0 _1175_.gnd
rlabel metal1 3544 2882 3636 2898 0 _1175_.vdd
rlabel metal2 3593 2733 3607 2747 0 _1175_.B
rlabel metal2 3553 2733 3567 2747 0 _1175_.A
rlabel metal2 3573 2713 3587 2727 0 _1175_.Y
rlabel nsubstratencontact 3796 2888 3796 2888 0 FILL_1__1198_.vdd
rlabel metal1 3784 2642 3816 2658 0 FILL_1__1198_.gnd
rlabel nsubstratencontact 3776 2888 3776 2888 0 FILL_0__1198_.vdd
rlabel metal1 3764 2642 3796 2658 0 FILL_0__1198_.gnd
rlabel metal1 3664 2642 3776 2658 0 _1587_.gnd
rlabel metal1 3664 2882 3776 2898 0 _1587_.vdd
rlabel metal2 3673 2753 3687 2767 0 _1587_.A
rlabel metal2 3693 2773 3707 2787 0 _1587_.B
rlabel metal2 3713 2753 3727 2767 0 _1587_.C
rlabel metal2 3733 2773 3747 2787 0 _1587_.Y
rlabel nsubstratencontact 3924 2888 3924 2888 0 FILL_1__976_.vdd
rlabel metal1 3904 2642 3936 2658 0 FILL_1__976_.gnd
rlabel nsubstratencontact 3904 2888 3904 2888 0 FILL_0__976_.vdd
rlabel metal1 3884 2642 3916 2658 0 FILL_0__976_.gnd
rlabel metal1 3804 2642 3896 2658 0 _1198_.gnd
rlabel metal1 3804 2882 3896 2898 0 _1198_.vdd
rlabel metal2 3813 2773 3827 2787 0 _1198_.A
rlabel metal2 3853 2773 3867 2787 0 _1198_.B
rlabel metal2 3833 2753 3847 2767 0 _1198_.Y
rlabel nsubstratencontact 4024 2888 4024 2888 0 FILL_1__1177_.vdd
rlabel metal1 4004 2642 4036 2658 0 FILL_1__1177_.gnd
rlabel nsubstratencontact 4004 2888 4004 2888 0 FILL_0__1177_.vdd
rlabel metal1 3984 2642 4016 2658 0 FILL_0__1177_.gnd
rlabel metal1 4024 2642 4136 2658 0 _1177_.gnd
rlabel metal1 4024 2882 4136 2898 0 _1177_.vdd
rlabel metal2 4113 2733 4127 2747 0 _1177_.A
rlabel metal2 4093 2753 4107 2767 0 _1177_.B
rlabel metal2 4053 2753 4067 2767 0 _1177_.C
rlabel metal2 4073 2733 4087 2747 0 _1177_.Y
rlabel metal1 3924 2642 3996 2658 0 _976_.gnd
rlabel metal1 3924 2882 3996 2898 0 _976_.vdd
rlabel metal2 3973 2753 3987 2767 0 _976_.A
rlabel metal2 3953 2733 3967 2747 0 _976_.Y
rlabel nsubstratencontact 4156 2888 4156 2888 0 FILL_1__975_.vdd
rlabel metal1 4144 2642 4176 2658 0 FILL_1__975_.gnd
rlabel nsubstratencontact 4276 2888 4276 2888 0 FILL_1__924_.vdd
rlabel metal1 4264 2642 4296 2658 0 FILL_1__924_.gnd
rlabel nsubstratencontact 4136 2888 4136 2888 0 FILL_0__975_.vdd
rlabel metal1 4124 2642 4156 2658 0 FILL_0__975_.gnd
rlabel nsubstratencontact 4256 2888 4256 2888 0 FILL_0__924_.vdd
rlabel metal1 4244 2642 4276 2658 0 FILL_0__924_.gnd
rlabel metal1 4164 2642 4256 2658 0 _975_.gnd
rlabel metal1 4164 2882 4256 2898 0 _975_.vdd
rlabel metal2 4173 2773 4187 2787 0 _975_.A
rlabel metal2 4213 2773 4227 2787 0 _975_.B
rlabel metal2 4193 2753 4207 2767 0 _975_.Y
rlabel metal1 4284 2642 4356 2658 0 _924_.gnd
rlabel metal1 4284 2882 4356 2898 0 _924_.vdd
rlabel metal2 4293 2753 4307 2767 0 _924_.A
rlabel metal2 4313 2733 4327 2747 0 _924_.Y
rlabel nsubstratencontact 4376 2888 4376 2888 0 FILL_1__1176_.vdd
rlabel metal1 4364 2642 4396 2658 0 FILL_1__1176_.gnd
rlabel nsubstratencontact 4356 2888 4356 2888 0 FILL_0__1176_.vdd
rlabel metal1 4344 2642 4376 2658 0 FILL_0__1176_.gnd
rlabel metal1 4384 2642 4456 2658 0 _1176_.gnd
rlabel metal1 4384 2882 4456 2898 0 _1176_.vdd
rlabel metal2 4393 2713 4407 2727 0 _1176_.A
rlabel metal2 4413 2753 4427 2767 0 _1176_.Y
rlabel metal1 4444 2642 4696 2658 0 _1671_.gnd
rlabel metal1 4444 2882 4696 2898 0 _1671_.vdd
rlabel metal2 4593 2733 4607 2747 0 _1671_.D
rlabel metal2 4553 2733 4567 2747 0 _1671_.CLK
rlabel metal2 4473 2733 4487 2747 0 _1671_.Q
rlabel metal1 4984 2642 5096 2658 0 _1605_.gnd
rlabel metal1 4984 2882 5096 2898 0 _1605_.vdd
rlabel metal2 4993 2733 5007 2747 0 _1605_.A
rlabel metal2 5013 2753 5027 2767 0 _1605_.B
rlabel metal2 5053 2753 5067 2767 0 _1605_.C
rlabel metal2 5033 2733 5047 2747 0 _1605_.Y
rlabel metal1 4684 2642 4936 2658 0 _1679_.gnd
rlabel metal1 4684 2882 4936 2898 0 _1679_.vdd
rlabel metal2 4773 2733 4787 2747 0 _1679_.D
rlabel metal2 4813 2733 4827 2747 0 _1679_.CLK
rlabel metal2 4893 2733 4907 2747 0 _1679_.Q
rlabel nsubstratencontact 4936 2888 4936 2888 0 FILL_0__1605_.vdd
rlabel metal1 4924 2642 4956 2658 0 FILL_0__1605_.gnd
rlabel nsubstratencontact 4956 2888 4956 2888 0 FILL_1__1605_.vdd
rlabel metal1 4944 2642 4976 2658 0 FILL_1__1605_.gnd
rlabel nsubstratencontact 4976 2888 4976 2888 0 FILL_2__1605_.vdd
rlabel metal1 4964 2642 4996 2658 0 FILL_2__1605_.gnd
rlabel metal1 5124 2642 5216 2658 0 _1604_.gnd
rlabel metal1 5124 2882 5216 2898 0 _1604_.vdd
rlabel metal2 5133 2773 5147 2787 0 _1604_.A
rlabel metal2 5173 2773 5187 2787 0 _1604_.B
rlabel metal2 5153 2753 5167 2767 0 _1604_.Y
rlabel metal1 5324 2642 5576 2658 0 _1653_.gnd
rlabel metal1 5324 2882 5576 2898 0 _1653_.vdd
rlabel metal2 5473 2733 5487 2747 0 _1653_.D
rlabel metal2 5433 2733 5447 2747 0 _1653_.CLK
rlabel metal2 5353 2733 5367 2747 0 _1653_.Q
rlabel metal1 5244 2642 5336 2658 0 _1686_.gnd
rlabel metal1 5244 2882 5336 2898 0 _1686_.vdd
rlabel metal2 5253 2753 5267 2767 0 _1686_.A
rlabel metal2 5293 2753 5307 2767 0 _1686_.Y
rlabel nsubstratencontact 5096 2888 5096 2888 0 FILL_0__1604_.vdd
rlabel metal1 5084 2642 5116 2658 0 FILL_0__1604_.gnd
rlabel nsubstratencontact 5216 2888 5216 2888 0 FILL_0__1686_.vdd
rlabel metal1 5204 2642 5236 2658 0 FILL_0__1686_.gnd
rlabel nsubstratencontact 5116 2888 5116 2888 0 FILL_1__1604_.vdd
rlabel metal1 5104 2642 5136 2658 0 FILL_1__1604_.gnd
rlabel nsubstratencontact 5236 2888 5236 2888 0 FILL_1__1686_.vdd
rlabel metal1 5224 2642 5256 2658 0 FILL_1__1686_.gnd
rlabel metal1 5604 2642 5716 2658 0 _1599_.gnd
rlabel metal1 5604 2882 5716 2898 0 _1599_.vdd
rlabel metal2 5613 2733 5627 2747 0 _1599_.A
rlabel metal2 5633 2753 5647 2767 0 _1599_.B
rlabel metal2 5673 2753 5687 2767 0 _1599_.C
rlabel metal2 5653 2733 5667 2747 0 _1599_.Y
rlabel nsubstratencontact 5716 2888 5716 2888 0 FILL85650x39750.vdd
rlabel metal1 5704 2642 5736 2658 0 FILL85650x39750.gnd
rlabel nsubstratencontact 5736 2888 5736 2888 0 FILL85950x39750.vdd
rlabel metal1 5724 2642 5756 2658 0 FILL85950x39750.gnd
rlabel nsubstratencontact 5756 2888 5756 2888 0 FILL86250x39750.vdd
rlabel metal1 5744 2642 5776 2658 0 FILL86250x39750.gnd
rlabel nsubstratencontact 5776 2888 5776 2888 0 FILL86550x39750.vdd
rlabel metal1 5764 2642 5796 2658 0 FILL86550x39750.gnd
rlabel nsubstratencontact 5796 2888 5796 2888 0 FILL86850x39750.vdd
rlabel metal1 5784 2642 5816 2658 0 FILL86850x39750.gnd
rlabel nsubstratencontact 5576 2888 5576 2888 0 FILL_0__1599_.vdd
rlabel metal1 5564 2642 5596 2658 0 FILL_0__1599_.gnd
rlabel nsubstratencontact 5596 2888 5596 2888 0 FILL_1__1599_.vdd
rlabel metal1 5584 2642 5616 2658 0 FILL_1__1599_.gnd
rlabel nsubstratencontact 64 2892 64 2892 0 FILL_2__1167_.vdd
rlabel metal1 44 3122 76 3138 0 FILL_2__1167_.gnd
rlabel nsubstratencontact 144 3368 144 3368 0 FILL_1__1190_.vdd
rlabel metal1 124 3122 156 3138 0 FILL_1__1190_.gnd
rlabel nsubstratencontact 44 2892 44 2892 0 FILL_1__1167_.vdd
rlabel metal1 24 3122 56 3138 0 FILL_1__1167_.gnd
rlabel nsubstratencontact 44 3368 44 3368 0 FILL_1__1164_.vdd
rlabel metal1 24 3122 56 3138 0 FILL_1__1164_.gnd
rlabel nsubstratencontact 124 3368 124 3368 0 FILL_0__1190_.vdd
rlabel metal1 104 3122 136 3138 0 FILL_0__1190_.gnd
rlabel nsubstratencontact 24 2892 24 2892 0 FILL_0__1167_.vdd
rlabel metal1 4 3122 36 3138 0 FILL_0__1167_.gnd
rlabel nsubstratencontact 24 3368 24 3368 0 FILL_0__1164_.vdd
rlabel metal1 4 3122 36 3138 0 FILL_0__1164_.gnd
rlabel metal1 64 3122 176 3138 0 _1167_.gnd
rlabel metal1 64 2882 176 2898 0 _1167_.vdd
rlabel metal2 153 3033 167 3047 0 _1167_.A
rlabel metal2 93 3033 107 3047 0 _1167_.Y
rlabel metal2 113 2993 127 3007 0 _1167_.B
rlabel metal1 44 3122 116 3138 0 _1164_.gnd
rlabel metal1 44 3362 116 3378 0 _1164_.vdd
rlabel metal2 93 3193 107 3207 0 _1164_.A
rlabel metal2 73 3233 87 3247 0 _1164_.Y
rlabel nsubstratencontact 216 2892 216 2892 0 FILL_2__1265_.vdd
rlabel metal1 204 3122 236 3138 0 FILL_2__1265_.gnd
rlabel nsubstratencontact 196 2892 196 2892 0 FILL_1__1265_.vdd
rlabel metal1 184 3122 216 3138 0 FILL_1__1265_.gnd
rlabel nsubstratencontact 176 2892 176 2892 0 FILL_0__1265_.vdd
rlabel metal1 164 3122 196 3138 0 FILL_0__1265_.gnd
rlabel nsubstratencontact 264 3368 264 3368 0 FILL_0__1189_.vdd
rlabel metal1 244 3122 276 3138 0 FILL_0__1189_.gnd
rlabel metal1 224 3122 336 3138 0 _1265_.gnd
rlabel metal1 224 2882 336 2898 0 _1265_.vdd
rlabel metal2 233 3013 247 3027 0 _1265_.A
rlabel metal2 253 2993 267 3007 0 _1265_.B
rlabel metal2 273 3013 287 3027 0 _1265_.C
rlabel metal2 293 2993 307 3007 0 _1265_.Y
rlabel metal1 144 3122 256 3138 0 _1190_.gnd
rlabel metal1 144 3362 256 3378 0 _1190_.vdd
rlabel metal2 233 3213 247 3227 0 _1190_.A
rlabel metal2 213 3233 227 3247 0 _1190_.B
rlabel metal2 173 3233 187 3247 0 _1190_.C
rlabel metal2 193 3213 207 3227 0 _1190_.Y
rlabel nsubstratencontact 376 3368 376 3368 0 FILL_1__1567_.vdd
rlabel metal1 364 3122 396 3138 0 FILL_1__1567_.gnd
rlabel nsubstratencontact 356 2892 356 2892 0 FILL_1__1264_.vdd
rlabel metal1 344 3122 376 3138 0 FILL_1__1264_.gnd
rlabel nsubstratencontact 284 3368 284 3368 0 FILL_1__1189_.vdd
rlabel metal1 264 3122 296 3138 0 FILL_1__1189_.gnd
rlabel nsubstratencontact 356 3368 356 3368 0 FILL_0__1567_.vdd
rlabel metal1 344 3122 376 3138 0 FILL_0__1567_.gnd
rlabel nsubstratencontact 336 2892 336 2892 0 FILL_0__1264_.vdd
rlabel metal1 324 3122 356 3138 0 FILL_0__1264_.gnd
rlabel metal1 364 3122 456 3138 0 _1264_.gnd
rlabel metal1 364 2882 456 2898 0 _1264_.vdd
rlabel metal2 373 2993 387 3007 0 _1264_.A
rlabel metal2 413 2993 427 3007 0 _1264_.B
rlabel metal2 393 3013 407 3027 0 _1264_.Y
rlabel metal1 284 3122 356 3138 0 _1189_.gnd
rlabel metal1 284 3362 356 3378 0 _1189_.vdd
rlabel metal2 333 3193 347 3207 0 _1189_.A
rlabel metal2 313 3233 327 3247 0 _1189_.Y
rlabel nsubstratencontact 496 3368 496 3368 0 FILL_1__1568_.vdd
rlabel metal1 484 3122 516 3138 0 FILL_1__1568_.gnd
rlabel nsubstratencontact 484 2892 484 2892 0 FILL_1__1266_.vdd
rlabel metal1 464 3122 496 3138 0 FILL_1__1266_.gnd
rlabel nsubstratencontact 476 3368 476 3368 0 FILL_0__1568_.vdd
rlabel metal1 464 3122 496 3138 0 FILL_0__1568_.gnd
rlabel nsubstratencontact 464 2892 464 2892 0 FILL_0__1266_.vdd
rlabel metal1 444 3122 476 3138 0 FILL_0__1266_.gnd
rlabel metal1 384 3122 476 3138 0 _1567_.gnd
rlabel metal1 384 3362 476 3378 0 _1567_.vdd
rlabel metal2 393 3253 407 3267 0 _1567_.A
rlabel metal2 433 3253 447 3267 0 _1567_.B
rlabel metal2 413 3233 427 3247 0 _1567_.Y
rlabel metal1 484 3122 596 3138 0 _1266_.gnd
rlabel metal1 484 2882 596 2898 0 _1266_.vdd
rlabel metal2 573 3033 587 3047 0 _1266_.A
rlabel metal2 553 3013 567 3027 0 _1266_.B
rlabel metal2 513 3013 527 3027 0 _1266_.C
rlabel metal2 533 3033 547 3047 0 _1266_.Y
rlabel metal1 504 3122 616 3138 0 _1568_.gnd
rlabel metal1 504 3362 616 3378 0 _1568_.vdd
rlabel metal2 513 3233 527 3247 0 _1568_.A
rlabel metal2 533 3193 547 3207 0 _1568_.B
rlabel metal2 553 3233 567 3247 0 _1568_.C
rlabel metal2 573 3213 587 3227 0 _1568_.Y
rlabel nsubstratencontact 616 2892 616 2892 0 FILL_1__1569_.vdd
rlabel metal1 604 3122 636 3138 0 FILL_1__1569_.gnd
rlabel nsubstratencontact 636 3368 636 3368 0 FILL_1__1360_.vdd
rlabel metal1 624 3122 656 3138 0 FILL_1__1360_.gnd
rlabel nsubstratencontact 596 2892 596 2892 0 FILL_0__1569_.vdd
rlabel metal1 584 3122 616 3138 0 FILL_0__1569_.gnd
rlabel nsubstratencontact 616 3368 616 3368 0 FILL_0__1360_.vdd
rlabel metal1 604 3122 636 3138 0 FILL_0__1360_.gnd
rlabel metal1 624 3122 736 3138 0 _1569_.gnd
rlabel metal1 624 2882 736 2898 0 _1569_.vdd
rlabel metal2 633 3033 647 3047 0 _1569_.A
rlabel metal2 653 3013 667 3027 0 _1569_.B
rlabel metal2 693 3013 707 3027 0 _1569_.C
rlabel metal2 673 3033 687 3047 0 _1569_.Y
rlabel nsubstratencontact 756 2892 756 2892 0 FILL_1__1359_.vdd
rlabel metal1 744 3122 776 3138 0 FILL_1__1359_.gnd
rlabel nsubstratencontact 736 2892 736 2892 0 FILL_0__1359_.vdd
rlabel metal1 724 3122 756 3138 0 FILL_0__1359_.gnd
rlabel nsubstratencontact 764 3368 764 3368 0 FILL_0__1357_.vdd
rlabel metal1 744 3122 776 3138 0 FILL_0__1357_.gnd
rlabel metal1 644 3122 756 3138 0 _1360_.gnd
rlabel metal1 644 3362 756 3378 0 _1360_.vdd
rlabel metal2 653 3213 667 3227 0 _1360_.A
rlabel metal2 713 3213 727 3227 0 _1360_.Y
rlabel metal2 693 3253 707 3267 0 _1360_.B
rlabel nsubstratencontact 804 3368 804 3368 0 FILL_2__1357_.vdd
rlabel metal1 784 3122 816 3138 0 FILL_2__1357_.gnd
rlabel nsubstratencontact 784 3368 784 3368 0 FILL_1__1357_.vdd
rlabel metal1 764 3122 796 3138 0 FILL_1__1357_.gnd
rlabel nsubstratencontact 876 2892 876 2892 0 FILL_0__1361_.vdd
rlabel metal1 864 3122 896 3138 0 FILL_0__1361_.gnd
rlabel metal1 764 3122 876 3138 0 _1359_.gnd
rlabel metal1 764 2882 876 2898 0 _1359_.vdd
rlabel metal2 773 3033 787 3047 0 _1359_.A
rlabel metal2 793 3013 807 3027 0 _1359_.B
rlabel metal2 833 3013 847 3027 0 _1359_.C
rlabel metal2 813 3033 827 3047 0 _1359_.Y
rlabel metal1 804 3122 896 3138 0 _1357_.gnd
rlabel metal1 804 3362 896 3378 0 _1357_.vdd
rlabel metal2 873 3253 887 3267 0 _1357_.A
rlabel metal2 833 3253 847 3267 0 _1357_.B
rlabel metal2 853 3233 867 3247 0 _1357_.Y
rlabel nsubstratencontact 896 2892 896 2892 0 FILL_1__1361_.vdd
rlabel metal1 884 3122 916 3138 0 FILL_1__1361_.gnd
rlabel nsubstratencontact 924 3368 924 3368 0 FILL_1__1356_.vdd
rlabel metal1 904 3122 936 3138 0 FILL_1__1356_.gnd
rlabel nsubstratencontact 904 3368 904 3368 0 FILL_0__1356_.vdd
rlabel metal1 884 3122 916 3138 0 FILL_0__1356_.gnd
rlabel nsubstratencontact 1024 2892 1024 2892 0 FILL_0__1269_.vdd
rlabel metal1 1004 3122 1036 3138 0 FILL_0__1269_.gnd
rlabel metal1 904 3122 1016 3138 0 _1361_.gnd
rlabel metal1 904 2882 1016 2898 0 _1361_.vdd
rlabel metal2 913 3033 927 3047 0 _1361_.A
rlabel metal2 933 3013 947 3027 0 _1361_.B
rlabel metal2 973 3013 987 3027 0 _1361_.C
rlabel metal2 953 3033 967 3047 0 _1361_.Y
rlabel metal1 924 3122 1036 3138 0 _1356_.gnd
rlabel metal1 924 3362 1036 3378 0 _1356_.vdd
rlabel metal2 1013 3233 1027 3247 0 _1356_.A
rlabel metal2 993 3253 1007 3267 0 _1356_.B
rlabel metal2 973 3233 987 3247 0 _1356_.C
rlabel metal2 953 3253 967 3267 0 _1356_.Y
rlabel nsubstratencontact 1064 3368 1064 3368 0 FILL_1__1355_.vdd
rlabel metal1 1044 3122 1076 3138 0 FILL_1__1355_.gnd
rlabel nsubstratencontact 1044 2892 1044 2892 0 FILL_1__1269_.vdd
rlabel metal1 1024 3122 1056 3138 0 FILL_1__1269_.gnd
rlabel nsubstratencontact 1144 2892 1144 2892 0 FILL_0__1474_.vdd
rlabel metal1 1124 3122 1156 3138 0 FILL_0__1474_.gnd
rlabel nsubstratencontact 1044 3368 1044 3368 0 FILL_0__1355_.vdd
rlabel metal1 1024 3122 1056 3138 0 FILL_0__1355_.gnd
rlabel metal1 1064 3122 1176 3138 0 _1355_.gnd
rlabel metal1 1064 3362 1176 3378 0 _1355_.vdd
rlabel metal2 1153 3233 1167 3247 0 _1355_.A
rlabel metal2 1133 3253 1147 3267 0 _1355_.B
rlabel metal2 1113 3233 1127 3247 0 _1355_.C
rlabel metal2 1093 3253 1107 3267 0 _1355_.Y
rlabel metal1 1044 3122 1136 3138 0 _1269_.gnd
rlabel metal1 1044 2882 1136 2898 0 _1269_.vdd
rlabel metal2 1113 2993 1127 3007 0 _1269_.A
rlabel metal2 1073 2993 1087 3007 0 _1269_.B
rlabel metal2 1093 3013 1107 3027 0 _1269_.Y
rlabel nsubstratencontact 1184 2892 1184 2892 0 FILL_2__1474_.vdd
rlabel metal1 1164 3122 1196 3138 0 FILL_2__1474_.gnd
rlabel nsubstratencontact 1164 2892 1164 2892 0 FILL_1__1474_.vdd
rlabel metal1 1144 3122 1176 3138 0 FILL_1__1474_.gnd
rlabel nsubstratencontact 1196 3368 1196 3368 0 FILL_1__1347_.vdd
rlabel metal1 1184 3122 1216 3138 0 FILL_1__1347_.gnd
rlabel nsubstratencontact 1176 3368 1176 3368 0 FILL_0__1347_.vdd
rlabel metal1 1164 3122 1196 3138 0 FILL_0__1347_.gnd
rlabel metal1 1184 3122 1276 3138 0 _1474_.gnd
rlabel metal1 1184 2882 1276 2898 0 _1474_.vdd
rlabel metal2 1213 3033 1227 3047 0 _1474_.B
rlabel metal2 1253 3033 1267 3047 0 _1474_.A
rlabel metal2 1233 3053 1247 3067 0 _1474_.Y
rlabel metal1 1204 3122 1316 3138 0 _1347_.gnd
rlabel metal1 1204 3362 1316 3378 0 _1347_.vdd
rlabel metal2 1213 3233 1227 3247 0 _1347_.A
rlabel metal2 1233 3193 1247 3207 0 _1347_.B
rlabel metal2 1253 3233 1267 3247 0 _1347_.C
rlabel metal2 1273 3213 1287 3227 0 _1347_.Y
rlabel nsubstratencontact 1296 2892 1296 2892 0 FILL_1__1351_.vdd
rlabel metal1 1284 3122 1316 3138 0 FILL_1__1351_.gnd
rlabel nsubstratencontact 1344 3368 1344 3368 0 FILL_1__1288_.vdd
rlabel metal1 1324 3122 1356 3138 0 FILL_1__1288_.gnd
rlabel nsubstratencontact 1276 2892 1276 2892 0 FILL_0__1351_.vdd
rlabel metal1 1264 3122 1296 3138 0 FILL_0__1351_.gnd
rlabel nsubstratencontact 1324 3368 1324 3368 0 FILL_0__1288_.vdd
rlabel metal1 1304 3122 1336 3138 0 FILL_0__1288_.gnd
rlabel metal1 1304 3122 1416 3138 0 _1351_.gnd
rlabel metal1 1304 2882 1416 2898 0 _1351_.vdd
rlabel metal2 1313 3033 1327 3047 0 _1351_.A
rlabel metal2 1333 3013 1347 3027 0 _1351_.B
rlabel metal2 1373 3013 1387 3027 0 _1351_.C
rlabel metal2 1353 3033 1367 3047 0 _1351_.Y
rlabel metal1 1344 3122 1416 3138 0 _1288_.gnd
rlabel metal1 1344 3362 1416 3378 0 _1288_.vdd
rlabel metal2 1393 3193 1407 3207 0 _1288_.A
rlabel metal2 1373 3233 1387 3247 0 _1288_.Y
rlabel nsubstratencontact 1444 2892 1444 2892 0 FILL_1__1354_.vdd
rlabel metal1 1424 3122 1456 3138 0 FILL_1__1354_.gnd
rlabel nsubstratencontact 1444 3368 1444 3368 0 FILL_1__1339_.vdd
rlabel metal1 1424 3122 1456 3138 0 FILL_1__1339_.gnd
rlabel nsubstratencontact 1424 2892 1424 2892 0 FILL_0__1354_.vdd
rlabel metal1 1404 3122 1436 3138 0 FILL_0__1354_.gnd
rlabel nsubstratencontact 1424 3368 1424 3368 0 FILL_0__1339_.vdd
rlabel metal1 1404 3122 1436 3138 0 FILL_0__1339_.gnd
rlabel metal1 1444 3122 1556 3138 0 _1354_.gnd
rlabel metal1 1444 2882 1556 2898 0 _1354_.vdd
rlabel metal2 1533 3013 1547 3027 0 _1354_.A
rlabel metal2 1513 2993 1527 3007 0 _1354_.B
rlabel metal2 1493 3013 1507 3027 0 _1354_.C
rlabel metal2 1473 2993 1487 3007 0 _1354_.Y
rlabel metal1 1444 3122 1556 3138 0 _1339_.gnd
rlabel metal1 1444 3362 1556 3378 0 _1339_.vdd
rlabel metal2 1533 3233 1547 3247 0 _1339_.A
rlabel metal2 1513 3253 1527 3267 0 _1339_.B
rlabel metal2 1493 3233 1507 3247 0 _1339_.C
rlabel metal2 1473 3253 1487 3267 0 _1339_.Y
rlabel nsubstratencontact 1604 2892 1604 2892 0 FILL_2__1350_.vdd
rlabel metal1 1584 3122 1616 3138 0 FILL_2__1350_.gnd
rlabel nsubstratencontact 1584 2892 1584 2892 0 FILL_1__1350_.vdd
rlabel metal1 1564 3122 1596 3138 0 FILL_1__1350_.gnd
rlabel nsubstratencontact 1584 3368 1584 3368 0 FILL_1__1348_.vdd
rlabel metal1 1564 3122 1596 3138 0 FILL_1__1348_.gnd
rlabel nsubstratencontact 1564 2892 1564 2892 0 FILL_0__1350_.vdd
rlabel metal1 1544 3122 1576 3138 0 FILL_0__1350_.gnd
rlabel nsubstratencontact 1564 3368 1564 3368 0 FILL_0__1348_.vdd
rlabel metal1 1544 3122 1576 3138 0 FILL_0__1348_.gnd
rlabel metal1 1604 3122 1716 3138 0 _1350_.gnd
rlabel metal1 1604 2882 1716 2898 0 _1350_.vdd
rlabel metal2 1693 3013 1707 3027 0 _1350_.A
rlabel metal2 1673 3053 1687 3067 0 _1350_.B
rlabel metal2 1653 3013 1667 3027 0 _1350_.C
rlabel metal2 1633 3033 1647 3047 0 _1350_.Y
rlabel metal1 1584 3122 1696 3138 0 _1348_.gnd
rlabel metal1 1584 3362 1696 3378 0 _1348_.vdd
rlabel metal2 1673 3233 1687 3247 0 _1348_.A
rlabel metal2 1653 3253 1667 3267 0 _1348_.B
rlabel metal2 1633 3233 1647 3247 0 _1348_.C
rlabel metal2 1613 3253 1627 3267 0 _1348_.Y
rlabel nsubstratencontact 1744 2892 1744 2892 0 FILL_1__1346_.vdd
rlabel metal1 1724 3122 1756 3138 0 FILL_1__1346_.gnd
rlabel nsubstratencontact 1724 3368 1724 3368 0 FILL_1__1342_.vdd
rlabel metal1 1704 3122 1736 3138 0 FILL_1__1342_.gnd
rlabel nsubstratencontact 1724 2892 1724 2892 0 FILL_0__1346_.vdd
rlabel metal1 1704 3122 1736 3138 0 FILL_0__1346_.gnd
rlabel nsubstratencontact 1704 3368 1704 3368 0 FILL_0__1342_.vdd
rlabel metal1 1684 3122 1716 3138 0 FILL_0__1342_.gnd
rlabel metal1 1744 3122 1856 3138 0 _1346_.gnd
rlabel metal1 1744 2882 1856 2898 0 _1346_.vdd
rlabel metal2 1833 3033 1847 3047 0 _1346_.A
rlabel metal2 1813 3013 1827 3027 0 _1346_.B
rlabel metal2 1773 3013 1787 3027 0 _1346_.C
rlabel metal2 1793 3033 1807 3047 0 _1346_.Y
rlabel metal1 1724 3122 1836 3138 0 _1342_.gnd
rlabel metal1 1724 3362 1836 3378 0 _1342_.vdd
rlabel metal2 1813 3233 1827 3247 0 _1342_.A
rlabel metal2 1793 3193 1807 3207 0 _1342_.B
rlabel metal2 1773 3233 1787 3247 0 _1342_.C
rlabel metal2 1753 3213 1767 3227 0 _1342_.Y
rlabel nsubstratencontact 1884 3368 1884 3368 0 FILL_2__1337_.vdd
rlabel metal1 1864 3122 1896 3138 0 FILL_2__1337_.gnd
rlabel nsubstratencontact 1876 2892 1876 2892 0 FILL_1__1349_.vdd
rlabel metal1 1864 3122 1896 3138 0 FILL_1__1349_.gnd
rlabel nsubstratencontact 1864 3368 1864 3368 0 FILL_1__1337_.vdd
rlabel metal1 1844 3122 1876 3138 0 FILL_1__1337_.gnd
rlabel nsubstratencontact 1856 2892 1856 2892 0 FILL_0__1349_.vdd
rlabel metal1 1844 3122 1876 3138 0 FILL_0__1349_.gnd
rlabel nsubstratencontact 1844 3368 1844 3368 0 FILL_0__1337_.vdd
rlabel metal1 1824 3122 1856 3138 0 FILL_0__1337_.gnd
rlabel metal1 1884 3122 1996 3138 0 _1349_.gnd
rlabel metal1 1884 2882 1996 2898 0 _1349_.vdd
rlabel metal2 1893 3033 1907 3047 0 _1349_.A
rlabel metal2 1913 3013 1927 3027 0 _1349_.B
rlabel metal2 1953 3013 1967 3027 0 _1349_.C
rlabel metal2 1933 3033 1947 3047 0 _1349_.Y
rlabel metal1 1884 3122 1976 3138 0 _1337_.gnd
rlabel metal1 1884 3362 1976 3378 0 _1337_.vdd
rlabel metal2 1953 3253 1967 3267 0 _1337_.A
rlabel metal2 1913 3253 1927 3267 0 _1337_.B
rlabel metal2 1933 3233 1947 3247 0 _1337_.Y
rlabel nsubstratencontact 2004 3368 2004 3368 0 FILL_1__1345_.vdd
rlabel metal1 1984 3122 2016 3138 0 FILL_1__1345_.gnd
rlabel nsubstratencontact 2024 2892 2024 2892 0 FILL_1__1344_.vdd
rlabel metal1 2004 3122 2036 3138 0 FILL_1__1344_.gnd
rlabel nsubstratencontact 1984 3368 1984 3368 0 FILL_0__1345_.vdd
rlabel metal1 1964 3122 1996 3138 0 FILL_0__1345_.gnd
rlabel nsubstratencontact 2004 2892 2004 2892 0 FILL_0__1344_.vdd
rlabel metal1 1984 3122 2016 3138 0 FILL_0__1344_.gnd
rlabel metal1 2004 3122 2116 3138 0 _1345_.gnd
rlabel metal1 2004 3362 2116 3378 0 _1345_.vdd
rlabel metal2 2093 3233 2107 3247 0 _1345_.A
rlabel metal2 2073 3193 2087 3207 0 _1345_.B
rlabel metal2 2053 3233 2067 3247 0 _1345_.C
rlabel metal2 2033 3213 2047 3227 0 _1345_.Y
rlabel nsubstratencontact 2044 2892 2044 2892 0 FILL_2__1344_.vdd
rlabel metal1 2024 3122 2056 3138 0 FILL_2__1344_.gnd
rlabel nsubstratencontact 2136 3368 2136 3368 0 FILL_1__1343_.vdd
rlabel metal1 2124 3122 2156 3138 0 FILL_1__1343_.gnd
rlabel nsubstratencontact 2116 3368 2116 3368 0 FILL_0__1343_.vdd
rlabel metal1 2104 3122 2136 3138 0 FILL_0__1343_.gnd
rlabel nsubstratencontact 2164 2892 2164 2892 0 FILL_0__1335_.vdd
rlabel metal1 2144 3122 2176 3138 0 FILL_0__1335_.gnd
rlabel metal1 2044 3122 2156 3138 0 _1344_.gnd
rlabel metal1 2044 2882 2156 2898 0 _1344_.vdd
rlabel metal2 2133 3033 2147 3047 0 _1344_.A
rlabel metal2 2113 3013 2127 3027 0 _1344_.B
rlabel metal2 2073 3013 2087 3027 0 _1344_.C
rlabel metal2 2093 3033 2107 3047 0 _1344_.Y
rlabel metal1 2144 3122 2236 3138 0 _1343_.gnd
rlabel metal1 2144 3362 2236 3378 0 _1343_.vdd
rlabel metal2 2153 3253 2167 3267 0 _1343_.A
rlabel metal2 2193 3253 2207 3267 0 _1343_.B
rlabel metal2 2173 3233 2187 3247 0 _1343_.Y
rlabel nsubstratencontact 2184 2892 2184 2892 0 FILL_1__1335_.vdd
rlabel metal1 2164 3122 2196 3138 0 FILL_1__1335_.gnd
rlabel nsubstratencontact 2264 3368 2264 3368 0 FILL_1__1334_.vdd
rlabel metal1 2244 3122 2276 3138 0 FILL_1__1334_.gnd
rlabel nsubstratencontact 2244 3368 2244 3368 0 FILL_0__1334_.vdd
rlabel metal1 2224 3122 2256 3138 0 FILL_0__1334_.gnd
rlabel metal1 2184 3122 2296 3138 0 _1335_.gnd
rlabel metal1 2184 2882 2296 2898 0 _1335_.vdd
rlabel metal2 2273 3033 2287 3047 0 _1335_.A
rlabel metal2 2253 3013 2267 3027 0 _1335_.B
rlabel metal2 2213 3013 2227 3027 0 _1335_.C
rlabel metal2 2233 3033 2247 3047 0 _1335_.Y
rlabel metal1 2264 3122 2376 3138 0 _1334_.gnd
rlabel metal1 2264 3362 2376 3378 0 _1334_.vdd
rlabel metal2 2353 3213 2367 3227 0 _1334_.A
rlabel metal2 2293 3213 2307 3227 0 _1334_.Y
rlabel metal2 2313 3253 2327 3267 0 _1334_.B
rlabel nsubstratencontact 2344 2892 2344 2892 0 FILL_2__1324_.vdd
rlabel metal1 2324 3122 2356 3138 0 FILL_2__1324_.gnd
rlabel nsubstratencontact 2324 2892 2324 2892 0 FILL_1__1324_.vdd
rlabel metal1 2304 3122 2336 3138 0 FILL_1__1324_.gnd
rlabel nsubstratencontact 2396 3368 2396 3368 0 FILL_1__1323_.vdd
rlabel metal1 2384 3122 2416 3138 0 FILL_1__1323_.gnd
rlabel nsubstratencontact 2304 2892 2304 2892 0 FILL_0__1324_.vdd
rlabel metal1 2284 3122 2316 3138 0 FILL_0__1324_.gnd
rlabel nsubstratencontact 2376 3368 2376 3368 0 FILL_0__1323_.vdd
rlabel metal1 2364 3122 2396 3138 0 FILL_0__1323_.gnd
rlabel metal1 2344 3122 2456 3138 0 _1324_.gnd
rlabel metal1 2344 2882 2456 2898 0 _1324_.vdd
rlabel metal2 2433 3013 2447 3027 0 _1324_.A
rlabel metal2 2413 3053 2427 3067 0 _1324_.B
rlabel metal2 2393 3013 2407 3027 0 _1324_.C
rlabel metal2 2373 3033 2387 3047 0 _1324_.Y
rlabel nsubstratencontact 2484 2892 2484 2892 0 FILL_1__1336_.vdd
rlabel metal1 2464 3122 2496 3138 0 FILL_1__1336_.gnd
rlabel nsubstratencontact 2524 3368 2524 3368 0 FILL_1__1329_.vdd
rlabel metal1 2504 3122 2536 3138 0 FILL_1__1329_.gnd
rlabel nsubstratencontact 2464 2892 2464 2892 0 FILL_0__1336_.vdd
rlabel metal1 2444 3122 2476 3138 0 FILL_0__1336_.gnd
rlabel nsubstratencontact 2504 3368 2504 3368 0 FILL_0__1329_.vdd
rlabel metal1 2484 3122 2516 3138 0 FILL_0__1329_.gnd
rlabel metal1 2484 3122 2596 3138 0 _1336_.gnd
rlabel metal1 2484 2882 2596 2898 0 _1336_.vdd
rlabel metal2 2573 3013 2587 3027 0 _1336_.A
rlabel metal2 2553 3053 2567 3067 0 _1336_.B
rlabel metal2 2533 3013 2547 3027 0 _1336_.C
rlabel metal2 2513 3033 2527 3047 0 _1336_.Y
rlabel metal1 2404 3122 2496 3138 0 _1323_.gnd
rlabel metal1 2404 3362 2496 3378 0 _1323_.vdd
rlabel metal2 2413 3253 2427 3267 0 _1323_.A
rlabel metal2 2453 3253 2467 3267 0 _1323_.B
rlabel metal2 2433 3233 2447 3247 0 _1323_.Y
rlabel metal1 2524 3122 2636 3138 0 _1329_.gnd
rlabel metal1 2524 3362 2636 3378 0 _1329_.vdd
rlabel metal2 2613 3213 2627 3227 0 _1329_.A
rlabel metal2 2593 3233 2607 3247 0 _1329_.B
rlabel metal2 2553 3233 2567 3247 0 _1329_.C
rlabel metal2 2573 3213 2587 3227 0 _1329_.Y
rlabel nsubstratencontact 2664 3368 2664 3368 0 FILL_1__1328_.vdd
rlabel metal1 2644 3122 2676 3138 0 FILL_1__1328_.gnd
rlabel nsubstratencontact 2624 2892 2624 2892 0 FILL_1__1237_.vdd
rlabel metal1 2604 3122 2636 3138 0 FILL_1__1237_.gnd
rlabel nsubstratencontact 2644 3368 2644 3368 0 FILL_0__1328_.vdd
rlabel metal1 2624 3122 2656 3138 0 FILL_0__1328_.gnd
rlabel nsubstratencontact 2604 2892 2604 2892 0 FILL_0__1237_.vdd
rlabel metal1 2584 3122 2616 3138 0 FILL_0__1237_.gnd
rlabel metal1 2664 3122 2776 3138 0 _1328_.gnd
rlabel metal1 2664 3362 2776 3378 0 _1328_.vdd
rlabel metal2 2753 3233 2767 3247 0 _1328_.A
rlabel metal2 2733 3193 2747 3207 0 _1328_.B
rlabel metal2 2713 3233 2727 3247 0 _1328_.C
rlabel metal2 2693 3213 2707 3227 0 _1328_.Y
rlabel metal1 2624 3122 2756 3138 0 _1237_.gnd
rlabel metal1 2624 2882 2756 2898 0 _1237_.vdd
rlabel metal2 2733 3033 2747 3047 0 _1237_.A
rlabel metal2 2713 3013 2727 3027 0 _1237_.B
rlabel metal2 2653 3033 2667 3047 0 _1237_.C
rlabel metal2 2673 3013 2687 3027 0 _1237_.D
rlabel metal2 2693 3033 2707 3047 0 _1237_.Y
rlabel nsubstratencontact 2784 2892 2784 2892 0 FILL_1__1325_.vdd
rlabel metal1 2764 3122 2796 3138 0 FILL_1__1325_.gnd
rlabel nsubstratencontact 2796 3368 2796 3368 0 FILL_1__1222_.vdd
rlabel metal1 2784 3122 2816 3138 0 FILL_1__1222_.gnd
rlabel nsubstratencontact 2764 2892 2764 2892 0 FILL_0__1325_.vdd
rlabel metal1 2744 3122 2776 3138 0 FILL_0__1325_.gnd
rlabel nsubstratencontact 2776 3368 2776 3368 0 FILL_0__1222_.vdd
rlabel metal1 2764 3122 2796 3138 0 FILL_0__1222_.gnd
rlabel metal1 2784 3122 2896 3138 0 _1325_.gnd
rlabel metal1 2784 2882 2896 2898 0 _1325_.vdd
rlabel metal2 2873 3053 2887 3067 0 _1325_.A
rlabel metal2 2853 3033 2867 3047 0 _1325_.B
rlabel metal2 2813 3013 2827 3027 0 _1325_.Y
rlabel metal1 2804 3122 2916 3138 0 _1222_.gnd
rlabel metal1 2804 3362 2916 3378 0 _1222_.vdd
rlabel metal2 2813 3233 2827 3247 0 _1222_.A
rlabel metal2 2833 3253 2847 3267 0 _1222_.B
rlabel metal2 2853 3233 2867 3247 0 _1222_.C
rlabel metal2 2873 3253 2887 3267 0 _1222_.Y
rlabel nsubstratencontact 2916 2892 2916 2892 0 FILL_1__1224_.vdd
rlabel metal1 2904 3122 2936 3138 0 FILL_1__1224_.gnd
rlabel nsubstratencontact 2936 3368 2936 3368 0 FILL_1__1210_.vdd
rlabel metal1 2924 3122 2956 3138 0 FILL_1__1210_.gnd
rlabel nsubstratencontact 2896 2892 2896 2892 0 FILL_0__1224_.vdd
rlabel metal1 2884 3122 2916 3138 0 FILL_0__1224_.gnd
rlabel nsubstratencontact 2916 3368 2916 3368 0 FILL_0__1210_.vdd
rlabel metal1 2904 3122 2936 3138 0 FILL_0__1210_.gnd
rlabel metal1 2924 3122 3016 3138 0 _1224_.gnd
rlabel metal1 2924 2882 3016 2898 0 _1224_.vdd
rlabel metal2 2973 3033 2987 3047 0 _1224_.B
rlabel metal2 2933 3033 2947 3047 0 _1224_.A
rlabel metal2 2953 3053 2967 3067 0 _1224_.Y
rlabel metal1 2944 3122 3056 3138 0 _1210_.gnd
rlabel metal1 2944 3362 3056 3378 0 _1210_.vdd
rlabel metal2 2953 3233 2967 3247 0 _1210_.A
rlabel metal2 2973 3253 2987 3267 0 _1210_.B
rlabel metal2 2993 3233 3007 3247 0 _1210_.C
rlabel metal2 3013 3253 3027 3267 0 _1210_.Y
rlabel nsubstratencontact 3036 2892 3036 2892 0 FILL_1__1220_.vdd
rlabel metal1 3024 3122 3056 3138 0 FILL_1__1220_.gnd
rlabel nsubstratencontact 3016 2892 3016 2892 0 FILL_0__1220_.vdd
rlabel metal1 3004 3122 3036 3138 0 FILL_0__1220_.gnd
rlabel nsubstratencontact 3056 2892 3056 2892 0 FILL_2__1220_.vdd
rlabel metal1 3044 3122 3076 3138 0 FILL_2__1220_.gnd
rlabel nsubstratencontact 3084 3368 3084 3368 0 FILL_1__1149_.vdd
rlabel metal1 3064 3122 3096 3138 0 FILL_1__1149_.gnd
rlabel nsubstratencontact 3164 2892 3164 2892 0 FILL_0__1231_.vdd
rlabel metal1 3144 3122 3176 3138 0 FILL_0__1231_.gnd
rlabel nsubstratencontact 3064 3368 3064 3368 0 FILL_0__1149_.vdd
rlabel metal1 3044 3122 3076 3138 0 FILL_0__1149_.gnd
rlabel metal1 3064 3122 3156 3138 0 _1220_.gnd
rlabel metal1 3064 2882 3156 2898 0 _1220_.vdd
rlabel metal2 3073 2993 3087 3007 0 _1220_.A
rlabel metal2 3113 2993 3127 3007 0 _1220_.B
rlabel metal2 3093 3013 3107 3027 0 _1220_.Y
rlabel metal1 3084 3122 3176 3138 0 _1149_.gnd
rlabel metal1 3084 3362 3176 3378 0 _1149_.vdd
rlabel metal2 3153 3253 3167 3267 0 _1149_.A
rlabel metal2 3113 3253 3127 3267 0 _1149_.B
rlabel metal2 3133 3233 3147 3247 0 _1149_.Y
rlabel nsubstratencontact 3224 3368 3224 3368 0 FILL_2__1174_.vdd
rlabel metal1 3204 3122 3236 3138 0 FILL_2__1174_.gnd
rlabel nsubstratencontact 3184 2892 3184 2892 0 FILL_1__1231_.vdd
rlabel metal1 3164 3122 3196 3138 0 FILL_1__1231_.gnd
rlabel nsubstratencontact 3204 3368 3204 3368 0 FILL_1__1174_.vdd
rlabel metal1 3184 3122 3216 3138 0 FILL_1__1174_.gnd
rlabel nsubstratencontact 3184 3368 3184 3368 0 FILL_0__1174_.vdd
rlabel metal1 3164 3122 3196 3138 0 FILL_0__1174_.gnd
rlabel metal1 3184 3122 3296 3138 0 _1231_.gnd
rlabel metal1 3184 2882 3296 2898 0 _1231_.vdd
rlabel metal2 3273 3033 3287 3047 0 _1231_.A
rlabel metal2 3213 3033 3227 3047 0 _1231_.Y
rlabel metal2 3233 2993 3247 3007 0 _1231_.B
rlabel metal1 3224 3122 3316 3138 0 _1174_.gnd
rlabel metal1 3224 3362 3316 3378 0 _1174_.vdd
rlabel metal2 3293 3253 3307 3267 0 _1174_.A
rlabel metal2 3253 3253 3267 3267 0 _1174_.B
rlabel metal2 3273 3233 3287 3247 0 _1174_.Y
rlabel nsubstratencontact 3336 3368 3336 3368 0 FILL_1__1215_.vdd
rlabel metal1 3324 3122 3356 3138 0 FILL_1__1215_.gnd
rlabel nsubstratencontact 3316 2892 3316 2892 0 FILL_1__1172_.vdd
rlabel metal1 3304 3122 3336 3138 0 FILL_1__1172_.gnd
rlabel nsubstratencontact 3424 3368 3424 3368 0 FILL_0__1219_.vdd
rlabel metal1 3404 3122 3436 3138 0 FILL_0__1219_.gnd
rlabel nsubstratencontact 3316 3368 3316 3368 0 FILL_0__1215_.vdd
rlabel metal1 3304 3122 3336 3138 0 FILL_0__1215_.gnd
rlabel nsubstratencontact 3296 2892 3296 2892 0 FILL_0__1172_.vdd
rlabel metal1 3284 3122 3316 3138 0 FILL_0__1172_.gnd
rlabel metal1 3344 3122 3416 3138 0 _1215_.gnd
rlabel metal1 3344 3362 3416 3378 0 _1215_.vdd
rlabel metal2 3353 3193 3367 3207 0 _1215_.A
rlabel metal2 3373 3233 3387 3247 0 _1215_.Y
rlabel metal1 3324 3122 3436 3138 0 _1172_.gnd
rlabel metal1 3324 2882 3436 2898 0 _1172_.vdd
rlabel metal2 3333 3053 3347 3067 0 _1172_.A
rlabel metal2 3353 3033 3367 3047 0 _1172_.B
rlabel metal2 3393 3013 3407 3027 0 _1172_.Y
rlabel nsubstratencontact 3464 2892 3464 2892 0 FILL_1__1294_.vdd
rlabel metal1 3444 3122 3476 3138 0 FILL_1__1294_.gnd
rlabel nsubstratencontact 3444 3368 3444 3368 0 FILL_1__1219_.vdd
rlabel metal1 3424 3122 3456 3138 0 FILL_1__1219_.gnd
rlabel nsubstratencontact 3444 2892 3444 2892 0 FILL_0__1294_.vdd
rlabel metal1 3424 3122 3456 3138 0 FILL_0__1294_.gnd
rlabel metal1 3464 3122 3576 3138 0 _1294_.gnd
rlabel metal1 3464 2882 3576 2898 0 _1294_.vdd
rlabel metal2 3553 3033 3567 3047 0 _1294_.A
rlabel metal2 3533 3013 3547 3027 0 _1294_.B
rlabel metal2 3493 3013 3507 3027 0 _1294_.C
rlabel metal2 3513 3033 3527 3047 0 _1294_.Y
rlabel metal1 3444 3122 3556 3138 0 _1219_.gnd
rlabel metal1 3444 3362 3556 3378 0 _1219_.vdd
rlabel metal2 3533 3233 3547 3247 0 _1219_.A
rlabel metal2 3513 3253 3527 3267 0 _1219_.B
rlabel metal2 3493 3233 3507 3247 0 _1219_.C
rlabel metal2 3473 3253 3487 3267 0 _1219_.Y
rlabel metal1 3604 3122 3716 3138 0 _1214_.gnd
rlabel metal1 3604 2882 3716 2898 0 _1214_.vdd
rlabel metal2 3693 3033 3707 3047 0 _1214_.A
rlabel metal2 3673 3013 3687 3027 0 _1214_.B
rlabel metal2 3633 3013 3647 3027 0 _1214_.C
rlabel metal2 3653 3033 3667 3047 0 _1214_.Y
rlabel metal1 3584 3122 3696 3138 0 _1297_.gnd
rlabel metal1 3584 3362 3696 3378 0 _1297_.vdd
rlabel metal2 3593 3233 3607 3247 0 _1297_.A
rlabel metal2 3613 3193 3627 3207 0 _1297_.B
rlabel metal2 3633 3233 3647 3247 0 _1297_.C
rlabel metal2 3653 3213 3667 3227 0 _1297_.Y
rlabel nsubstratencontact 3584 2892 3584 2892 0 FILL_0__1214_.vdd
rlabel metal1 3564 3122 3596 3138 0 FILL_0__1214_.gnd
rlabel nsubstratencontact 3556 3368 3556 3368 0 FILL_0__1297_.vdd
rlabel metal1 3544 3122 3576 3138 0 FILL_0__1297_.gnd
rlabel nsubstratencontact 3604 2892 3604 2892 0 FILL_1__1214_.vdd
rlabel metal1 3584 3122 3616 3138 0 FILL_1__1214_.gnd
rlabel nsubstratencontact 3576 3368 3576 3368 0 FILL_1__1297_.vdd
rlabel metal1 3564 3122 3596 3138 0 FILL_1__1297_.gnd
rlabel metal1 3744 3122 3856 3138 0 _1216_.gnd
rlabel metal1 3744 2882 3856 2898 0 _1216_.vdd
rlabel metal2 3833 3053 3847 3067 0 _1216_.A
rlabel metal2 3813 3033 3827 3047 0 _1216_.B
rlabel metal2 3773 3013 3787 3027 0 _1216_.Y
rlabel metal1 3724 3122 3836 3138 0 _1218_.gnd
rlabel metal1 3724 3362 3836 3378 0 _1218_.vdd
rlabel metal2 3813 3213 3827 3227 0 _1218_.A
rlabel metal2 3793 3233 3807 3247 0 _1218_.B
rlabel metal2 3753 3233 3767 3247 0 _1218_.C
rlabel metal2 3773 3213 3787 3227 0 _1218_.Y
rlabel nsubstratencontact 3724 2892 3724 2892 0 FILL_0__1216_.vdd
rlabel metal1 3704 3122 3736 3138 0 FILL_0__1216_.gnd
rlabel nsubstratencontact 3704 3368 3704 3368 0 FILL_0__1218_.vdd
rlabel metal1 3684 3122 3716 3138 0 FILL_0__1218_.gnd
rlabel nsubstratencontact 3744 2892 3744 2892 0 FILL_1__1216_.vdd
rlabel metal1 3724 3122 3756 3138 0 FILL_1__1216_.gnd
rlabel nsubstratencontact 3724 3368 3724 3368 0 FILL_1__1218_.vdd
rlabel metal1 3704 3122 3736 3138 0 FILL_1__1218_.gnd
rlabel nsubstratencontact 3904 2892 3904 2892 0 FILL_2__1213_.vdd
rlabel metal1 3884 3122 3916 3138 0 FILL_2__1213_.gnd
rlabel nsubstratencontact 3856 3368 3856 3368 0 FILL_1__1217_.vdd
rlabel metal1 3844 3122 3876 3138 0 FILL_1__1217_.gnd
rlabel nsubstratencontact 3884 2892 3884 2892 0 FILL_1__1213_.vdd
rlabel metal1 3864 3122 3896 3138 0 FILL_1__1213_.gnd
rlabel nsubstratencontact 4036 2892 4036 2892 0 FILL_1__1212_.vdd
rlabel metal1 4024 3122 4056 3138 0 FILL_1__1212_.gnd
rlabel nsubstratencontact 3836 3368 3836 3368 0 FILL_0__1217_.vdd
rlabel metal1 3824 3122 3856 3138 0 FILL_0__1217_.gnd
rlabel nsubstratencontact 3864 2892 3864 2892 0 FILL_0__1213_.vdd
rlabel metal1 3844 3122 3876 3138 0 FILL_0__1213_.gnd
rlabel nsubstratencontact 4016 2892 4016 2892 0 FILL_0__1212_.vdd
rlabel metal1 4004 3122 4036 3138 0 FILL_0__1212_.gnd
rlabel metal1 3864 3122 3936 3138 0 _1217_.gnd
rlabel metal1 3864 3362 3936 3378 0 _1217_.vdd
rlabel metal2 3873 3193 3887 3207 0 _1217_.A
rlabel metal2 3893 3233 3907 3247 0 _1217_.Y
rlabel metal1 3904 3122 4016 3138 0 _1213_.gnd
rlabel metal1 3904 2882 4016 2898 0 _1213_.vdd
rlabel metal2 3993 3033 4007 3047 0 _1213_.A
rlabel metal2 3933 3033 3947 3047 0 _1213_.Y
rlabel metal2 3953 2993 3967 3007 0 _1213_.B
rlabel metal1 3924 3122 4176 3138 0 _1670_.gnd
rlabel metal1 3924 3362 4176 3378 0 _1670_.vdd
rlabel metal2 4073 3213 4087 3227 0 _1670_.D
rlabel metal2 4033 3213 4047 3227 0 _1670_.CLK
rlabel metal2 3953 3213 3967 3227 0 _1670_.Q
rlabel nsubstratencontact 4196 3368 4196 3368 0 FILL_1__1623_.vdd
rlabel metal1 4184 3122 4216 3138 0 FILL_1__1623_.gnd
rlabel nsubstratencontact 4156 2892 4156 2892 0 FILL_1__1211_.vdd
rlabel metal1 4144 3122 4176 3138 0 FILL_1__1211_.gnd
rlabel nsubstratencontact 4176 3368 4176 3368 0 FILL_0__1623_.vdd
rlabel metal1 4164 3122 4196 3138 0 FILL_0__1623_.gnd
rlabel nsubstratencontact 4136 2892 4136 2892 0 FILL_0__1211_.vdd
rlabel metal1 4124 3122 4156 3138 0 FILL_0__1211_.gnd
rlabel metal1 4204 3122 4316 3138 0 _1623_.gnd
rlabel metal1 4204 3362 4316 3378 0 _1623_.vdd
rlabel metal2 4213 3213 4227 3227 0 _1623_.A
rlabel metal2 4233 3233 4247 3247 0 _1623_.B
rlabel metal2 4273 3233 4287 3247 0 _1623_.C
rlabel metal2 4253 3213 4267 3227 0 _1623_.Y
rlabel metal1 4044 3122 4136 3138 0 _1212_.gnd
rlabel metal1 4044 2882 4136 2898 0 _1212_.vdd
rlabel metal2 4093 3033 4107 3047 0 _1212_.B
rlabel metal2 4053 3033 4067 3047 0 _1212_.A
rlabel metal2 4073 3053 4087 3067 0 _1212_.Y
rlabel metal1 4164 3122 4276 3138 0 _1211_.gnd
rlabel metal1 4164 2882 4276 2898 0 _1211_.vdd
rlabel metal2 4173 3013 4187 3027 0 _1211_.A
rlabel metal2 4193 2993 4207 3007 0 _1211_.B
rlabel metal2 4213 3013 4227 3027 0 _1211_.C
rlabel metal2 4233 2993 4247 3007 0 _1211_.Y
rlabel nsubstratencontact 4556 2892 4556 2892 0 FILL_2__1625_.vdd
rlabel metal1 4544 3122 4576 3138 0 FILL_2__1625_.gnd
rlabel nsubstratencontact 4336 3368 4336 3368 0 FILL_1__1643_.vdd
rlabel metal1 4324 3122 4356 3138 0 FILL_1__1643_.gnd
rlabel nsubstratencontact 4536 2892 4536 2892 0 FILL_1__1625_.vdd
rlabel metal1 4524 3122 4556 3138 0 FILL_1__1625_.gnd
rlabel nsubstratencontact 4316 3368 4316 3368 0 FILL_0__1643_.vdd
rlabel metal1 4304 3122 4336 3138 0 FILL_0__1643_.gnd
rlabel nsubstratencontact 4516 2892 4516 2892 0 FILL_0__1625_.vdd
rlabel metal1 4504 3122 4536 3138 0 FILL_0__1625_.gnd
rlabel metal1 4344 3122 4456 3138 0 _1643_.gnd
rlabel metal1 4344 3362 4456 3378 0 _1643_.vdd
rlabel metal2 4353 3213 4367 3227 0 _1643_.A
rlabel metal2 4373 3233 4387 3247 0 _1643_.B
rlabel metal2 4413 3233 4427 3247 0 _1643_.C
rlabel metal2 4393 3213 4407 3227 0 _1643_.Y
rlabel metal1 4264 3122 4516 3138 0 _1680_.gnd
rlabel metal1 4264 2882 4516 2898 0 _1680_.vdd
rlabel metal2 4353 3033 4367 3047 0 _1680_.D
rlabel metal2 4393 3033 4407 3047 0 _1680_.CLK
rlabel metal2 4473 3033 4487 3047 0 _1680_.Q
rlabel metal1 4444 3122 4696 3138 0 _1669_.gnd
rlabel metal1 4444 3362 4696 3378 0 _1669_.vdd
rlabel metal2 4593 3213 4607 3227 0 _1669_.D
rlabel metal2 4553 3213 4567 3227 0 _1669_.CLK
rlabel metal2 4473 3213 4487 3227 0 _1669_.Q
rlabel nsubstratencontact 4696 2892 4696 2892 0 FILL_1__1641_.vdd
rlabel metal1 4684 3122 4716 3138 0 FILL_1__1641_.gnd
rlabel nsubstratencontact 4716 3368 4716 3368 0 FILL_1__1621_.vdd
rlabel metal1 4704 3122 4736 3138 0 FILL_1__1621_.gnd
rlabel nsubstratencontact 4676 2892 4676 2892 0 FILL_0__1641_.vdd
rlabel metal1 4664 3122 4696 3138 0 FILL_0__1641_.gnd
rlabel nsubstratencontact 4696 3368 4696 3368 0 FILL_0__1621_.vdd
rlabel metal1 4684 3122 4716 3138 0 FILL_0__1621_.gnd
rlabel metal1 4704 3122 4816 3138 0 _1641_.gnd
rlabel metal1 4704 2882 4816 2898 0 _1641_.vdd
rlabel metal2 4713 3033 4727 3047 0 _1641_.A
rlabel metal2 4733 3013 4747 3027 0 _1641_.B
rlabel metal2 4773 3013 4787 3027 0 _1641_.C
rlabel metal2 4753 3033 4767 3047 0 _1641_.Y
rlabel metal1 4564 3122 4676 3138 0 _1625_.gnd
rlabel metal1 4564 2882 4676 2898 0 _1625_.vdd
rlabel metal2 4573 3033 4587 3047 0 _1625_.A
rlabel metal2 4593 3013 4607 3027 0 _1625_.B
rlabel metal2 4633 3013 4647 3027 0 _1625_.C
rlabel metal2 4613 3033 4627 3047 0 _1625_.Y
rlabel metal1 4724 3122 4836 3138 0 _1621_.gnd
rlabel metal1 4724 3362 4836 3378 0 _1621_.vdd
rlabel metal2 4733 3213 4747 3227 0 _1621_.A
rlabel metal2 4753 3233 4767 3247 0 _1621_.B
rlabel metal2 4793 3233 4807 3247 0 _1621_.C
rlabel metal2 4773 3213 4787 3227 0 _1621_.Y
rlabel metal1 4864 3122 4956 3138 0 _1622_.gnd
rlabel metal1 4864 3362 4956 3378 0 _1622_.vdd
rlabel metal2 4933 3253 4947 3267 0 _1622_.A
rlabel metal2 4893 3253 4907 3267 0 _1622_.B
rlabel metal2 4913 3233 4927 3247 0 _1622_.Y
rlabel metal1 4844 3122 4936 3138 0 _1624_.gnd
rlabel metal1 4844 2882 4936 2898 0 _1624_.vdd
rlabel metal2 4913 2993 4927 3007 0 _1624_.A
rlabel metal2 4873 2993 4887 3007 0 _1624_.B
rlabel metal2 4893 3013 4907 3027 0 _1624_.Y
rlabel nsubstratencontact 4844 3368 4844 3368 0 FILL_0__1622_.vdd
rlabel metal1 4824 3122 4856 3138 0 FILL_0__1622_.gnd
rlabel nsubstratencontact 4824 2892 4824 2892 0 FILL_0__1624_.vdd
rlabel metal1 4804 3122 4836 3138 0 FILL_0__1624_.gnd
rlabel nsubstratencontact 4936 2892 4936 2892 0 FILL_0__1640_.vdd
rlabel metal1 4924 3122 4956 3138 0 FILL_0__1640_.gnd
rlabel nsubstratencontact 4864 3368 4864 3368 0 FILL_1__1622_.vdd
rlabel metal1 4844 3122 4876 3138 0 FILL_1__1622_.gnd
rlabel nsubstratencontact 4844 2892 4844 2892 0 FILL_1__1624_.vdd
rlabel metal1 4824 3122 4856 3138 0 FILL_1__1624_.gnd
rlabel metal1 4984 3122 5096 3138 0 _1608_.gnd
rlabel metal1 4984 3362 5096 3378 0 _1608_.vdd
rlabel metal2 5073 3213 5087 3227 0 _1608_.A
rlabel metal2 5053 3233 5067 3247 0 _1608_.B
rlabel metal2 5013 3233 5027 3247 0 _1608_.C
rlabel metal2 5033 3213 5047 3227 0 _1608_.Y
rlabel metal1 4964 3122 5056 3138 0 _1640_.gnd
rlabel metal1 4964 2882 5056 2898 0 _1640_.vdd
rlabel metal2 4973 2993 4987 3007 0 _1640_.A
rlabel metal2 5013 2993 5027 3007 0 _1640_.B
rlabel metal2 4993 3013 5007 3027 0 _1640_.Y
rlabel nsubstratencontact 4964 3368 4964 3368 0 FILL_0__1608_.vdd
rlabel metal1 4944 3122 4976 3138 0 FILL_0__1608_.gnd
rlabel nsubstratencontact 4984 3368 4984 3368 0 FILL_1__1608_.vdd
rlabel metal1 4964 3122 4996 3138 0 FILL_1__1608_.gnd
rlabel nsubstratencontact 4956 2892 4956 2892 0 FILL_1__1640_.vdd
rlabel metal1 4944 3122 4976 3138 0 FILL_1__1640_.gnd
rlabel metal1 5044 3122 5296 3138 0 _1656_.gnd
rlabel metal1 5044 2882 5296 2898 0 _1656_.vdd
rlabel metal2 5133 3033 5147 3047 0 _1656_.D
rlabel metal2 5173 3033 5187 3047 0 _1656_.CLK
rlabel metal2 5253 3033 5267 3047 0 _1656_.Q
rlabel nsubstratencontact 5324 2892 5324 2892 0 FILL_1_CLKBUF1_insert4.vdd
rlabel metal1 5304 3122 5336 3138 0 FILL_1_CLKBUF1_insert4.gnd
rlabel nsubstratencontact 5224 3368 5224 3368 0 FILL_1__1620_.vdd
rlabel metal1 5204 3122 5236 3138 0 FILL_1__1620_.gnd
rlabel nsubstratencontact 5124 3368 5124 3368 0 FILL_1__1606_.vdd
rlabel metal1 5104 3122 5136 3138 0 FILL_1__1606_.gnd
rlabel nsubstratencontact 5304 2892 5304 2892 0 FILL_0_CLKBUF1_insert4.vdd
rlabel metal1 5284 3122 5316 3138 0 FILL_0_CLKBUF1_insert4.gnd
rlabel nsubstratencontact 5204 3368 5204 3368 0 FILL_0__1620_.vdd
rlabel metal1 5184 3122 5216 3138 0 FILL_0__1620_.gnd
rlabel nsubstratencontact 5316 3368 5316 3368 0 FILL_0__1609_.vdd
rlabel metal1 5304 3122 5336 3138 0 FILL_0__1609_.gnd
rlabel nsubstratencontact 5104 3368 5104 3368 0 FILL_0__1606_.vdd
rlabel metal1 5084 3122 5116 3138 0 FILL_0__1606_.gnd
rlabel metal1 5224 3122 5316 3138 0 _1620_.gnd
rlabel metal1 5224 3362 5316 3378 0 _1620_.vdd
rlabel metal2 5293 3253 5307 3267 0 _1620_.A
rlabel metal2 5253 3253 5267 3267 0 _1620_.B
rlabel metal2 5273 3233 5287 3247 0 _1620_.Y
rlabel metal1 5124 3122 5196 3138 0 _1606_.gnd
rlabel metal1 5124 3362 5196 3378 0 _1606_.vdd
rlabel metal2 5173 3193 5187 3207 0 _1606_.A
rlabel metal2 5153 3233 5167 3247 0 _1606_.Y
rlabel nsubstratencontact 5456 3368 5456 3368 0 FILL_2__1611_.vdd
rlabel metal1 5444 3122 5476 3138 0 FILL_2__1611_.gnd
rlabel nsubstratencontact 5436 3368 5436 3368 0 FILL_1__1611_.vdd
rlabel metal1 5424 3122 5456 3138 0 FILL_1__1611_.gnd
rlabel nsubstratencontact 5336 3368 5336 3368 0 FILL_1__1609_.vdd
rlabel metal1 5324 3122 5356 3138 0 FILL_1__1609_.gnd
rlabel nsubstratencontact 5416 3368 5416 3368 0 FILL_0__1611_.vdd
rlabel metal1 5404 3122 5436 3138 0 FILL_0__1611_.gnd
rlabel metal1 5324 3122 5536 3138 0 CLKBUF1_insert4.gnd
rlabel metal1 5324 2882 5536 2898 0 CLKBUF1_insert4.vdd
rlabel metal2 5493 3013 5507 3027 0 CLKBUF1_insert4.A
rlabel metal2 5353 3013 5367 3027 0 CLKBUF1_insert4.Y
rlabel metal1 5464 3122 5576 3138 0 _1611_.gnd
rlabel metal1 5464 3362 5576 3378 0 _1611_.vdd
rlabel metal2 5473 3213 5487 3227 0 _1611_.A
rlabel metal2 5493 3233 5507 3247 0 _1611_.B
rlabel metal2 5533 3233 5547 3247 0 _1611_.C
rlabel metal2 5513 3213 5527 3227 0 _1611_.Y
rlabel metal1 5344 3122 5416 3138 0 _1609_.gnd
rlabel metal1 5344 3362 5416 3378 0 _1609_.vdd
rlabel metal2 5353 3193 5367 3207 0 _1609_.A
rlabel metal2 5373 3233 5387 3247 0 _1609_.Y
rlabel metal1 5524 3122 5776 3138 0 _1657_.gnd
rlabel metal1 5524 2882 5776 2898 0 _1657_.vdd
rlabel metal2 5673 3033 5687 3047 0 _1657_.D
rlabel metal2 5633 3033 5647 3047 0 _1657_.CLK
rlabel metal2 5553 3033 5567 3047 0 _1657_.Q
rlabel nsubstratencontact 5624 3368 5624 3368 0 FILL_2__1598_.vdd
rlabel metal1 5604 3122 5636 3138 0 FILL_2__1598_.gnd
rlabel nsubstratencontact 5604 3368 5604 3368 0 FILL_1__1598_.vdd
rlabel metal1 5584 3122 5616 3138 0 FILL_1__1598_.gnd
rlabel nsubstratencontact 5584 3368 5584 3368 0 FILL_0__1598_.vdd
rlabel metal1 5564 3122 5596 3138 0 FILL_0__1598_.gnd
rlabel metal1 5624 3122 5716 3138 0 _1598_.gnd
rlabel metal1 5624 3362 5716 3378 0 _1598_.vdd
rlabel metal2 5693 3253 5707 3267 0 _1598_.A
rlabel metal2 5653 3253 5667 3267 0 _1598_.B
rlabel metal2 5673 3233 5687 3247 0 _1598_.Y
rlabel nsubstratencontact 5776 3368 5776 3368 0 FILL86550x46950.vdd
rlabel metal1 5764 3122 5796 3138 0 FILL86550x46950.gnd
rlabel nsubstratencontact 5784 2892 5784 2892 0 FILL86550x43350.vdd
rlabel metal1 5764 3122 5796 3138 0 FILL86550x43350.gnd
rlabel nsubstratencontact 5756 3368 5756 3368 0 FILL86250x46950.vdd
rlabel metal1 5744 3122 5776 3138 0 FILL86250x46950.gnd
rlabel nsubstratencontact 5736 3368 5736 3368 0 FILL85950x46950.vdd
rlabel metal1 5724 3122 5756 3138 0 FILL85950x46950.gnd
rlabel nsubstratencontact 5716 3368 5716 3368 0 FILL85650x46950.vdd
rlabel metal1 5704 3122 5736 3138 0 FILL85650x46950.gnd
rlabel nsubstratencontact 5796 3368 5796 3368 0 FILL86850x46950.vdd
rlabel metal1 5784 3122 5816 3138 0 FILL86850x46950.gnd
rlabel nsubstratencontact 5804 2892 5804 2892 0 FILL86850x43350.vdd
rlabel metal1 5784 3122 5816 3138 0 FILL86850x43350.gnd
rlabel nsubstratencontact 44 3372 44 3372 0 FILL_1__1538_.vdd
rlabel metal1 24 3602 56 3618 0 FILL_1__1538_.gnd
rlabel nsubstratencontact 24 3372 24 3372 0 FILL_0__1538_.vdd
rlabel metal1 4 3602 36 3618 0 FILL_0__1538_.gnd
rlabel metal1 44 3602 156 3618 0 _1538_.gnd
rlabel metal1 44 3362 156 3378 0 _1538_.vdd
rlabel metal2 133 3513 147 3527 0 _1538_.A
rlabel metal2 113 3493 127 3507 0 _1538_.B
rlabel metal2 73 3493 87 3507 0 _1538_.C
rlabel metal2 93 3513 107 3527 0 _1538_.Y
rlabel nsubstratencontact 176 3372 176 3372 0 FILL_1__1539_.vdd
rlabel metal1 164 3602 196 3618 0 FILL_1__1539_.gnd
rlabel nsubstratencontact 156 3372 156 3372 0 FILL_0__1539_.vdd
rlabel metal1 144 3602 176 3618 0 FILL_0__1539_.gnd
rlabel metal1 184 3602 296 3618 0 _1539_.gnd
rlabel metal1 184 3362 296 3378 0 _1539_.vdd
rlabel metal2 193 3493 207 3507 0 _1539_.A
rlabel metal2 213 3533 227 3547 0 _1539_.B
rlabel metal2 233 3493 247 3507 0 _1539_.C
rlabel metal2 253 3513 267 3527 0 _1539_.Y
rlabel nsubstratencontact 316 3372 316 3372 0 FILL_1__1529_.vdd
rlabel metal1 304 3602 336 3618 0 FILL_1__1529_.gnd
rlabel nsubstratencontact 296 3372 296 3372 0 FILL_0__1529_.vdd
rlabel metal1 284 3602 316 3618 0 FILL_0__1529_.gnd
rlabel metal1 324 3602 396 3618 0 _1529_.gnd
rlabel metal1 324 3362 396 3378 0 _1529_.vdd
rlabel metal2 333 3533 347 3547 0 _1529_.A
rlabel metal2 353 3493 367 3507 0 _1529_.Y
rlabel nsubstratencontact 416 3372 416 3372 0 FILL_1__1530_.vdd
rlabel metal1 404 3602 436 3618 0 FILL_1__1530_.gnd
rlabel nsubstratencontact 396 3372 396 3372 0 FILL_0__1530_.vdd
rlabel metal1 384 3602 416 3618 0 FILL_0__1530_.gnd
rlabel metal1 424 3602 536 3618 0 _1530_.gnd
rlabel metal1 424 3362 536 3378 0 _1530_.vdd
rlabel metal2 433 3513 447 3527 0 _1530_.A
rlabel metal2 453 3493 467 3507 0 _1530_.B
rlabel metal2 493 3493 507 3507 0 _1530_.C
rlabel metal2 473 3513 487 3527 0 _1530_.Y
rlabel nsubstratencontact 556 3372 556 3372 0 FILL_1__1531_.vdd
rlabel metal1 544 3602 576 3618 0 FILL_1__1531_.gnd
rlabel nsubstratencontact 536 3372 536 3372 0 FILL_0__1531_.vdd
rlabel metal1 524 3602 556 3618 0 FILL_0__1531_.gnd
rlabel metal1 564 3602 676 3618 0 _1531_.gnd
rlabel metal1 564 3362 676 3378 0 _1531_.vdd
rlabel metal2 573 3493 587 3507 0 _1531_.A
rlabel metal2 593 3473 607 3487 0 _1531_.B
rlabel metal2 613 3493 627 3507 0 _1531_.C
rlabel metal2 633 3473 647 3487 0 _1531_.Y
rlabel nsubstratencontact 724 3372 724 3372 0 FILL_2__1363_.vdd
rlabel metal1 704 3602 736 3618 0 FILL_2__1363_.gnd
rlabel nsubstratencontact 704 3372 704 3372 0 FILL_1__1363_.vdd
rlabel metal1 684 3602 716 3618 0 FILL_1__1363_.gnd
rlabel nsubstratencontact 684 3372 684 3372 0 FILL_0__1363_.vdd
rlabel metal1 664 3602 696 3618 0 FILL_0__1363_.gnd
rlabel metal1 724 3602 816 3618 0 _1363_.gnd
rlabel metal1 724 3362 816 3378 0 _1363_.vdd
rlabel metal2 793 3473 807 3487 0 _1363_.A
rlabel metal2 753 3473 767 3487 0 _1363_.B
rlabel metal2 773 3493 787 3507 0 _1363_.Y
rlabel nsubstratencontact 844 3372 844 3372 0 FILL_1__1364_.vdd
rlabel metal1 824 3602 856 3618 0 FILL_1__1364_.gnd
rlabel nsubstratencontact 824 3372 824 3372 0 FILL_0__1364_.vdd
rlabel metal1 804 3602 836 3618 0 FILL_0__1364_.gnd
rlabel metal1 844 3602 936 3618 0 _1364_.gnd
rlabel metal1 844 3362 936 3378 0 _1364_.vdd
rlabel metal2 913 3473 927 3487 0 _1364_.A
rlabel metal2 873 3473 887 3487 0 _1364_.B
rlabel metal2 893 3493 907 3507 0 _1364_.Y
rlabel nsubstratencontact 956 3372 956 3372 0 FILL_1__1523_.vdd
rlabel metal1 944 3602 976 3618 0 FILL_1__1523_.gnd
rlabel nsubstratencontact 936 3372 936 3372 0 FILL_0__1523_.vdd
rlabel metal1 924 3602 956 3618 0 FILL_0__1523_.gnd
rlabel metal1 964 3602 1076 3618 0 _1523_.gnd
rlabel metal1 964 3362 1076 3378 0 _1523_.vdd
rlabel metal2 973 3513 987 3527 0 _1523_.A
rlabel metal2 993 3493 1007 3507 0 _1523_.B
rlabel metal2 1033 3493 1047 3507 0 _1523_.C
rlabel metal2 1013 3513 1027 3527 0 _1523_.Y
rlabel nsubstratencontact 1104 3372 1104 3372 0 FILL_1__1182_.vdd
rlabel metal1 1084 3602 1116 3618 0 FILL_1__1182_.gnd
rlabel nsubstratencontact 1084 3372 1084 3372 0 FILL_0__1182_.vdd
rlabel metal1 1064 3602 1096 3618 0 FILL_0__1182_.gnd
rlabel metal1 1104 3602 1216 3618 0 _1182_.gnd
rlabel metal1 1104 3362 1216 3378 0 _1182_.vdd
rlabel metal2 1193 3493 1207 3507 0 _1182_.A
rlabel metal2 1173 3473 1187 3487 0 _1182_.B
rlabel metal2 1153 3493 1167 3507 0 _1182_.C
rlabel metal2 1133 3473 1147 3487 0 _1182_.Y
rlabel nsubstratencontact 1236 3372 1236 3372 0 FILL_1__1480_.vdd
rlabel metal1 1224 3602 1256 3618 0 FILL_1__1480_.gnd
rlabel nsubstratencontact 1216 3372 1216 3372 0 FILL_0__1480_.vdd
rlabel metal1 1204 3602 1236 3618 0 FILL_0__1480_.gnd
rlabel metal1 1244 3602 1336 3618 0 _1480_.gnd
rlabel metal1 1244 3362 1336 3378 0 _1480_.vdd
rlabel metal2 1253 3473 1267 3487 0 _1480_.A
rlabel metal2 1293 3473 1307 3487 0 _1480_.B
rlabel metal2 1273 3493 1287 3507 0 _1480_.Y
rlabel nsubstratencontact 1364 3372 1364 3372 0 FILL_1__1418_.vdd
rlabel metal1 1344 3602 1376 3618 0 FILL_1__1418_.gnd
rlabel nsubstratencontact 1344 3372 1344 3372 0 FILL_0__1418_.vdd
rlabel metal1 1324 3602 1356 3618 0 FILL_0__1418_.gnd
rlabel metal1 1364 3602 1476 3618 0 _1418_.gnd
rlabel metal1 1364 3362 1476 3378 0 _1418_.vdd
rlabel metal2 1453 3493 1467 3507 0 _1418_.A
rlabel metal2 1433 3473 1447 3487 0 _1418_.B
rlabel metal2 1413 3493 1427 3507 0 _1418_.C
rlabel metal2 1393 3473 1407 3487 0 _1418_.Y
rlabel nsubstratencontact 1496 3372 1496 3372 0 FILL_1__1420_.vdd
rlabel metal1 1484 3602 1516 3618 0 FILL_1__1420_.gnd
rlabel nsubstratencontact 1476 3372 1476 3372 0 FILL_0__1420_.vdd
rlabel metal1 1464 3602 1496 3618 0 FILL_0__1420_.gnd
rlabel metal1 1504 3602 1616 3618 0 _1420_.gnd
rlabel metal1 1504 3362 1616 3378 0 _1420_.vdd
rlabel metal2 1513 3513 1527 3527 0 _1420_.A
rlabel metal2 1533 3493 1547 3507 0 _1420_.B
rlabel metal2 1573 3493 1587 3507 0 _1420_.C
rlabel metal2 1553 3513 1567 3527 0 _1420_.Y
rlabel metal1 1784 3602 1896 3618 0 _1338_.gnd
rlabel metal1 1784 3362 1896 3378 0 _1338_.vdd
rlabel metal2 1873 3493 1887 3507 0 _1338_.A
rlabel metal2 1853 3473 1867 3487 0 _1338_.B
rlabel metal2 1833 3493 1847 3507 0 _1338_.C
rlabel metal2 1813 3473 1827 3487 0 _1338_.Y
rlabel metal1 1924 3602 2036 3618 0 _1369_.gnd
rlabel metal1 1924 3362 2036 3378 0 _1369_.vdd
rlabel metal2 1933 3493 1947 3507 0 _1369_.A
rlabel metal2 1953 3533 1967 3547 0 _1369_.B
rlabel metal2 1973 3493 1987 3507 0 _1369_.C
rlabel metal2 1993 3513 2007 3527 0 _1369_.Y
rlabel metal1 1644 3602 1756 3618 0 _1419_.gnd
rlabel metal1 1644 3362 1756 3378 0 _1419_.vdd
rlabel metal2 1733 3493 1747 3507 0 _1419_.A
rlabel metal2 1713 3533 1727 3547 0 _1419_.B
rlabel metal2 1693 3493 1707 3507 0 _1419_.C
rlabel metal2 1673 3513 1687 3527 0 _1419_.Y
rlabel nsubstratencontact 1764 3372 1764 3372 0 FILL_0__1338_.vdd
rlabel metal1 1744 3602 1776 3618 0 FILL_0__1338_.gnd
rlabel nsubstratencontact 1896 3372 1896 3372 0 FILL_0__1369_.vdd
rlabel metal1 1884 3602 1916 3618 0 FILL_0__1369_.gnd
rlabel nsubstratencontact 1624 3372 1624 3372 0 FILL_0__1419_.vdd
rlabel metal1 1604 3602 1636 3618 0 FILL_0__1419_.gnd
rlabel nsubstratencontact 1784 3372 1784 3372 0 FILL_1__1338_.vdd
rlabel metal1 1764 3602 1796 3618 0 FILL_1__1338_.gnd
rlabel nsubstratencontact 1916 3372 1916 3372 0 FILL_1__1369_.vdd
rlabel metal1 1904 3602 1936 3618 0 FILL_1__1369_.gnd
rlabel nsubstratencontact 1644 3372 1644 3372 0 FILL_1__1419_.vdd
rlabel metal1 1624 3602 1656 3618 0 FILL_1__1419_.gnd
rlabel nsubstratencontact 2064 3372 2064 3372 0 FILL_1__1405_.vdd
rlabel metal1 2044 3602 2076 3618 0 FILL_1__1405_.gnd
rlabel nsubstratencontact 2044 3372 2044 3372 0 FILL_0__1405_.vdd
rlabel metal1 2024 3602 2056 3618 0 FILL_0__1405_.gnd
rlabel metal1 2064 3602 2176 3618 0 _1405_.gnd
rlabel metal1 2064 3362 2176 3378 0 _1405_.vdd
rlabel metal2 2153 3513 2167 3527 0 _1405_.A
rlabel metal2 2133 3493 2147 3507 0 _1405_.B
rlabel metal2 2093 3493 2107 3507 0 _1405_.C
rlabel metal2 2113 3513 2127 3527 0 _1405_.Y
rlabel nsubstratencontact 2216 3372 2216 3372 0 FILL_2__1331_.vdd
rlabel metal1 2204 3602 2236 3618 0 FILL_2__1331_.gnd
rlabel nsubstratencontact 2196 3372 2196 3372 0 FILL_1__1331_.vdd
rlabel metal1 2184 3602 2216 3618 0 FILL_1__1331_.gnd
rlabel nsubstratencontact 2176 3372 2176 3372 0 FILL_0__1331_.vdd
rlabel metal1 2164 3602 2196 3618 0 FILL_0__1331_.gnd
rlabel metal1 2224 3602 2336 3618 0 _1331_.gnd
rlabel metal1 2224 3362 2336 3378 0 _1331_.vdd
rlabel metal2 2233 3513 2247 3527 0 _1331_.A
rlabel metal2 2253 3493 2267 3507 0 _1331_.B
rlabel metal2 2293 3493 2307 3507 0 _1331_.C
rlabel metal2 2273 3513 2287 3527 0 _1331_.Y
rlabel nsubstratencontact 2364 3372 2364 3372 0 FILL_1__1330_.vdd
rlabel metal1 2344 3602 2376 3618 0 FILL_1__1330_.gnd
rlabel nsubstratencontact 2344 3372 2344 3372 0 FILL_0__1330_.vdd
rlabel metal1 2324 3602 2356 3618 0 FILL_0__1330_.gnd
rlabel metal1 2364 3602 2476 3618 0 _1330_.gnd
rlabel metal1 2364 3362 2476 3378 0 _1330_.vdd
rlabel metal2 2453 3493 2467 3507 0 _1330_.A
rlabel metal2 2433 3533 2447 3547 0 _1330_.B
rlabel metal2 2413 3493 2427 3507 0 _1330_.C
rlabel metal2 2393 3513 2407 3527 0 _1330_.Y
rlabel nsubstratencontact 2504 3372 2504 3372 0 FILL_1__1332_.vdd
rlabel metal1 2484 3602 2516 3618 0 FILL_1__1332_.gnd
rlabel nsubstratencontact 2484 3372 2484 3372 0 FILL_0__1332_.vdd
rlabel metal1 2464 3602 2496 3618 0 FILL_0__1332_.gnd
rlabel metal1 2504 3602 2616 3618 0 _1332_.gnd
rlabel metal1 2504 3362 2616 3378 0 _1332_.vdd
rlabel metal2 2593 3513 2607 3527 0 _1332_.A
rlabel metal2 2533 3513 2547 3527 0 _1332_.Y
rlabel metal2 2553 3473 2567 3487 0 _1332_.B
rlabel nsubstratencontact 2636 3372 2636 3372 0 FILL_1__1304_.vdd
rlabel metal1 2624 3602 2656 3618 0 FILL_1__1304_.gnd
rlabel nsubstratencontact 2616 3372 2616 3372 0 FILL_0__1304_.vdd
rlabel metal1 2604 3602 2636 3618 0 FILL_0__1304_.gnd
rlabel metal1 2644 3602 2736 3618 0 _1304_.gnd
rlabel metal1 2644 3362 2736 3378 0 _1304_.vdd
rlabel metal2 2653 3473 2667 3487 0 _1304_.A
rlabel metal2 2693 3473 2707 3487 0 _1304_.B
rlabel metal2 2673 3493 2687 3507 0 _1304_.Y
rlabel nsubstratencontact 2764 3372 2764 3372 0 FILL_1__1327_.vdd
rlabel metal1 2744 3602 2776 3618 0 FILL_1__1327_.gnd
rlabel nsubstratencontact 2744 3372 2744 3372 0 FILL_0__1327_.vdd
rlabel metal1 2724 3602 2756 3618 0 FILL_0__1327_.gnd
rlabel metal1 2764 3602 2876 3618 0 _1327_.gnd
rlabel metal1 2764 3362 2876 3378 0 _1327_.vdd
rlabel metal2 2853 3513 2867 3527 0 _1327_.A
rlabel metal2 2833 3493 2847 3507 0 _1327_.B
rlabel metal2 2793 3493 2807 3507 0 _1327_.C
rlabel metal2 2813 3513 2827 3527 0 _1327_.Y
rlabel nsubstratencontact 2904 3372 2904 3372 0 FILL_1_BUFX2_insert8.vdd
rlabel metal1 2884 3602 2916 3618 0 FILL_1_BUFX2_insert8.gnd
rlabel nsubstratencontact 2884 3372 2884 3372 0 FILL_0_BUFX2_insert8.vdd
rlabel metal1 2864 3602 2896 3618 0 FILL_0_BUFX2_insert8.gnd
rlabel nsubstratencontact 2924 3372 2924 3372 0 FILL_2_BUFX2_insert8.vdd
rlabel metal1 2904 3602 2936 3618 0 FILL_2_BUFX2_insert8.gnd
rlabel nsubstratencontact 3044 3372 3044 3372 0 FILL_1__1300_.vdd
rlabel metal1 3024 3602 3056 3618 0 FILL_1__1300_.gnd
rlabel nsubstratencontact 3024 3372 3024 3372 0 FILL_0__1300_.vdd
rlabel metal1 3004 3602 3036 3618 0 FILL_0__1300_.gnd
rlabel metal1 2924 3602 3016 3618 0 BUFX2_insert8.gnd
rlabel metal1 2924 3362 3016 3378 0 BUFX2_insert8.vdd
rlabel metal2 2993 3513 3007 3527 0 BUFX2_insert8.A
rlabel metal2 2953 3513 2967 3527 0 BUFX2_insert8.Y
rlabel nsubstratencontact 3156 3372 3156 3372 0 FILL_1__1295_.vdd
rlabel metal1 3144 3602 3176 3618 0 FILL_1__1295_.gnd
rlabel nsubstratencontact 3136 3372 3136 3372 0 FILL_0__1295_.vdd
rlabel metal1 3124 3602 3156 3618 0 FILL_0__1295_.gnd
rlabel metal1 3044 3602 3136 3618 0 _1300_.gnd
rlabel metal1 3044 3362 3136 3378 0 _1300_.vdd
rlabel metal2 3113 3473 3127 3487 0 _1300_.A
rlabel metal2 3073 3473 3087 3487 0 _1300_.B
rlabel metal2 3093 3493 3107 3507 0 _1300_.Y
rlabel nsubstratencontact 3284 3372 3284 3372 0 FILL_0__1299_.vdd
rlabel metal1 3264 3602 3296 3618 0 FILL_0__1299_.gnd
rlabel metal1 3164 3602 3276 3618 0 _1295_.gnd
rlabel metal1 3164 3362 3276 3378 0 _1295_.vdd
rlabel metal2 3173 3493 3187 3507 0 _1295_.A
rlabel metal2 3193 3473 3207 3487 0 _1295_.B
rlabel metal2 3213 3493 3227 3507 0 _1295_.C
rlabel metal2 3233 3473 3247 3487 0 _1295_.Y
rlabel nsubstratencontact 3304 3372 3304 3372 0 FILL_1__1299_.vdd
rlabel metal1 3284 3602 3316 3618 0 FILL_1__1299_.gnd
rlabel nsubstratencontact 3424 3372 3424 3372 0 FILL_0__1367_.vdd
rlabel metal1 3404 3602 3436 3618 0 FILL_0__1367_.gnd
rlabel metal1 3304 3602 3416 3618 0 _1299_.gnd
rlabel metal1 3304 3362 3416 3378 0 _1299_.vdd
rlabel metal2 3393 3493 3407 3507 0 _1299_.A
rlabel metal2 3373 3473 3387 3487 0 _1299_.B
rlabel metal2 3353 3493 3367 3507 0 _1299_.C
rlabel metal2 3333 3473 3347 3487 0 _1299_.Y
rlabel nsubstratencontact 3444 3372 3444 3372 0 FILL_1__1367_.vdd
rlabel metal1 3424 3602 3456 3618 0 FILL_1__1367_.gnd
rlabel metal1 3444 3602 3556 3618 0 _1367_.gnd
rlabel metal1 3444 3362 3556 3378 0 _1367_.vdd
rlabel metal2 3533 3513 3547 3527 0 _1367_.A
rlabel metal2 3513 3493 3527 3507 0 _1367_.B
rlabel metal2 3473 3493 3487 3507 0 _1367_.C
rlabel metal2 3493 3513 3507 3527 0 _1367_.Y
rlabel nsubstratencontact 3584 3372 3584 3372 0 FILL_1__1303_.vdd
rlabel metal1 3564 3602 3596 3618 0 FILL_1__1303_.gnd
rlabel nsubstratencontact 3564 3372 3564 3372 0 FILL_0__1303_.vdd
rlabel metal1 3544 3602 3576 3618 0 FILL_0__1303_.gnd
rlabel metal1 3584 3602 3696 3618 0 _1303_.gnd
rlabel metal1 3584 3362 3696 3378 0 _1303_.vdd
rlabel metal2 3673 3513 3687 3527 0 _1303_.A
rlabel metal2 3653 3493 3667 3507 0 _1303_.B
rlabel metal2 3613 3493 3627 3507 0 _1303_.C
rlabel metal2 3633 3513 3647 3527 0 _1303_.Y
rlabel nsubstratencontact 3724 3372 3724 3372 0 FILL_1__1302_.vdd
rlabel metal1 3704 3602 3736 3618 0 FILL_1__1302_.gnd
rlabel nsubstratencontact 3704 3372 3704 3372 0 FILL_0__1302_.vdd
rlabel metal1 3684 3602 3716 3618 0 FILL_0__1302_.gnd
rlabel metal1 3724 3602 3836 3618 0 _1302_.gnd
rlabel metal1 3724 3362 3836 3378 0 _1302_.vdd
rlabel metal2 3813 3513 3827 3527 0 _1302_.A
rlabel metal2 3753 3513 3767 3527 0 _1302_.Y
rlabel metal2 3773 3473 3787 3487 0 _1302_.B
rlabel nsubstratencontact 3856 3372 3856 3372 0 FILL_1__1301_.vdd
rlabel metal1 3844 3602 3876 3618 0 FILL_1__1301_.gnd
rlabel nsubstratencontact 3836 3372 3836 3372 0 FILL_0__1301_.vdd
rlabel metal1 3824 3602 3856 3618 0 FILL_0__1301_.gnd
rlabel metal1 3864 3602 3956 3618 0 _1301_.gnd
rlabel metal1 3864 3362 3956 3378 0 _1301_.vdd
rlabel metal2 3913 3513 3927 3527 0 _1301_.B
rlabel metal2 3873 3513 3887 3527 0 _1301_.A
rlabel metal2 3893 3533 3907 3547 0 _1301_.Y
rlabel nsubstratencontact 4004 3372 4004 3372 0 FILL_2__1298_.vdd
rlabel metal1 3984 3602 4016 3618 0 FILL_2__1298_.gnd
rlabel nsubstratencontact 3984 3372 3984 3372 0 FILL_1__1298_.vdd
rlabel metal1 3964 3602 3996 3618 0 FILL_1__1298_.gnd
rlabel nsubstratencontact 3964 3372 3964 3372 0 FILL_0__1298_.vdd
rlabel metal1 3944 3602 3976 3618 0 FILL_0__1298_.gnd
rlabel metal1 4004 3602 4116 3618 0 _1298_.gnd
rlabel metal1 4004 3362 4116 3378 0 _1298_.vdd
rlabel metal2 4093 3513 4107 3527 0 _1298_.A
rlabel metal2 4073 3493 4087 3507 0 _1298_.B
rlabel metal2 4033 3493 4047 3507 0 _1298_.C
rlabel metal2 4053 3513 4067 3527 0 _1298_.Y
rlabel nsubstratencontact 4136 3372 4136 3372 0 FILL_1__1296_.vdd
rlabel metal1 4124 3602 4156 3618 0 FILL_1__1296_.gnd
rlabel nsubstratencontact 4116 3372 4116 3372 0 FILL_0__1296_.vdd
rlabel metal1 4104 3602 4136 3618 0 FILL_0__1296_.gnd
rlabel metal1 4144 3602 4216 3618 0 _1296_.gnd
rlabel metal1 4144 3362 4216 3378 0 _1296_.vdd
rlabel metal2 4153 3533 4167 3547 0 _1296_.A
rlabel metal2 4173 3493 4187 3507 0 _1296_.Y
rlabel nsubstratencontact 4236 3372 4236 3372 0 FILL_1__1627_.vdd
rlabel metal1 4224 3602 4256 3618 0 FILL_1__1627_.gnd
rlabel nsubstratencontact 4216 3372 4216 3372 0 FILL_0__1627_.vdd
rlabel metal1 4204 3602 4236 3618 0 FILL_0__1627_.gnd
rlabel metal1 4244 3602 4356 3618 0 _1627_.gnd
rlabel metal1 4244 3362 4356 3378 0 _1627_.vdd
rlabel metal2 4253 3513 4267 3527 0 _1627_.A
rlabel metal2 4273 3493 4287 3507 0 _1627_.B
rlabel metal2 4313 3493 4327 3507 0 _1627_.C
rlabel metal2 4293 3513 4307 3527 0 _1627_.Y
rlabel nsubstratencontact 4384 3372 4384 3372 0 FILL_1__1642_.vdd
rlabel metal1 4364 3602 4396 3618 0 FILL_1__1642_.gnd
rlabel nsubstratencontact 4364 3372 4364 3372 0 FILL_0__1642_.vdd
rlabel metal1 4344 3602 4376 3618 0 FILL_0__1642_.gnd
rlabel metal1 4384 3602 4476 3618 0 _1642_.gnd
rlabel metal1 4384 3362 4476 3378 0 _1642_.vdd
rlabel metal2 4453 3473 4467 3487 0 _1642_.A
rlabel metal2 4413 3473 4427 3487 0 _1642_.B
rlabel metal2 4433 3493 4447 3507 0 _1642_.Y
rlabel nsubstratencontact 4496 3372 4496 3372 0 FILL_1__1626_.vdd
rlabel metal1 4484 3602 4516 3618 0 FILL_1__1626_.gnd
rlabel nsubstratencontact 4476 3372 4476 3372 0 FILL_0__1626_.vdd
rlabel metal1 4464 3602 4496 3618 0 FILL_0__1626_.gnd
rlabel metal1 4504 3602 4596 3618 0 _1626_.gnd
rlabel metal1 4504 3362 4596 3378 0 _1626_.vdd
rlabel metal2 4513 3473 4527 3487 0 _1626_.A
rlabel metal2 4553 3473 4567 3487 0 _1626_.B
rlabel metal2 4533 3493 4547 3507 0 _1626_.Y
rlabel metal1 4864 3602 4956 3618 0 _1607_.gnd
rlabel metal1 4864 3362 4956 3378 0 _1607_.vdd
rlabel metal2 4933 3473 4947 3487 0 _1607_.A
rlabel metal2 4893 3473 4907 3487 0 _1607_.B
rlabel metal2 4913 3493 4927 3507 0 _1607_.Y
rlabel metal1 4984 3602 5096 3618 0 _1639_.gnd
rlabel metal1 4984 3362 5096 3378 0 _1639_.vdd
rlabel metal2 5073 3513 5087 3527 0 _1639_.A
rlabel metal2 5053 3493 5067 3507 0 _1639_.B
rlabel metal2 5013 3493 5027 3507 0 _1639_.C
rlabel metal2 5033 3513 5047 3527 0 _1639_.Y
rlabel metal1 4584 3602 4836 3618 0 _1681_.gnd
rlabel metal1 4584 3362 4836 3378 0 _1681_.vdd
rlabel metal2 4733 3513 4747 3527 0 _1681_.D
rlabel metal2 4693 3513 4707 3527 0 _1681_.CLK
rlabel metal2 4613 3513 4627 3527 0 _1681_.Q
rlabel nsubstratencontact 4844 3372 4844 3372 0 FILL_0__1607_.vdd
rlabel metal1 4824 3602 4856 3618 0 FILL_0__1607_.gnd
rlabel nsubstratencontact 4964 3372 4964 3372 0 FILL_0__1639_.vdd
rlabel metal1 4944 3602 4976 3618 0 FILL_0__1639_.gnd
rlabel nsubstratencontact 4864 3372 4864 3372 0 FILL_1__1607_.vdd
rlabel metal1 4844 3602 4876 3618 0 FILL_1__1607_.gnd
rlabel nsubstratencontact 4984 3372 4984 3372 0 FILL_1__1639_.vdd
rlabel metal1 4964 3602 4996 3618 0 FILL_1__1639_.gnd
rlabel metal1 5504 3602 5596 3618 0 _1610_.gnd
rlabel metal1 5504 3362 5596 3378 0 _1610_.vdd
rlabel metal2 5573 3473 5587 3487 0 _1610_.A
rlabel metal2 5533 3473 5547 3487 0 _1610_.B
rlabel metal2 5553 3493 5567 3507 0 _1610_.Y
rlabel metal1 5144 3602 5236 3618 0 _1638_.gnd
rlabel metal1 5144 3362 5236 3378 0 _1638_.vdd
rlabel metal2 5153 3473 5167 3487 0 _1638_.A
rlabel metal2 5193 3473 5207 3487 0 _1638_.B
rlabel metal2 5173 3493 5187 3507 0 _1638_.Y
rlabel metal1 5224 3602 5476 3618 0 _1678_.gnd
rlabel metal1 5224 3362 5476 3378 0 _1678_.vdd
rlabel metal2 5313 3513 5327 3527 0 _1678_.D
rlabel metal2 5353 3513 5367 3527 0 _1678_.CLK
rlabel metal2 5433 3513 5447 3527 0 _1678_.Q
rlabel nsubstratencontact 5484 3372 5484 3372 0 FILL_0__1610_.vdd
rlabel metal1 5464 3602 5496 3618 0 FILL_0__1610_.gnd
rlabel nsubstratencontact 5096 3372 5096 3372 0 FILL_0__1638_.vdd
rlabel metal1 5084 3602 5116 3618 0 FILL_0__1638_.gnd
rlabel nsubstratencontact 5504 3372 5504 3372 0 FILL_1__1610_.vdd
rlabel metal1 5484 3602 5516 3618 0 FILL_1__1610_.gnd
rlabel nsubstratencontact 5116 3372 5116 3372 0 FILL_1__1638_.vdd
rlabel metal1 5104 3602 5136 3618 0 FILL_1__1638_.gnd
rlabel nsubstratencontact 5136 3372 5136 3372 0 FILL_2__1638_.vdd
rlabel metal1 5124 3602 5156 3618 0 FILL_2__1638_.gnd
rlabel metal1 5624 3602 5736 3618 0 _1602_.gnd
rlabel metal1 5624 3362 5736 3378 0 _1602_.vdd
rlabel metal2 5633 3513 5647 3527 0 _1602_.A
rlabel metal2 5653 3493 5667 3507 0 _1602_.B
rlabel metal2 5693 3493 5707 3507 0 _1602_.C
rlabel metal2 5673 3513 5687 3527 0 _1602_.Y
rlabel nsubstratencontact 5744 3372 5744 3372 0 FILL85950x50550.vdd
rlabel metal1 5724 3602 5756 3618 0 FILL85950x50550.gnd
rlabel nsubstratencontact 5764 3372 5764 3372 0 FILL86250x50550.vdd
rlabel metal1 5744 3602 5776 3618 0 FILL86250x50550.gnd
rlabel nsubstratencontact 5784 3372 5784 3372 0 FILL86550x50550.vdd
rlabel metal1 5764 3602 5796 3618 0 FILL86550x50550.gnd
rlabel nsubstratencontact 5804 3372 5804 3372 0 FILL86850x50550.vdd
rlabel metal1 5784 3602 5816 3618 0 FILL86850x50550.gnd
rlabel nsubstratencontact 5596 3372 5596 3372 0 FILL_0__1602_.vdd
rlabel metal1 5584 3602 5616 3618 0 FILL_0__1602_.gnd
rlabel nsubstratencontact 5616 3372 5616 3372 0 FILL_1__1602_.vdd
rlabel metal1 5604 3602 5636 3618 0 FILL_1__1602_.gnd
rlabel nsubstratencontact 44 3848 44 3848 0 FILL_1__1537_.vdd
rlabel metal1 24 3602 56 3618 0 FILL_1__1537_.gnd
rlabel nsubstratencontact 164 3848 164 3848 0 FILL_1__1188_.vdd
rlabel metal1 144 3602 176 3618 0 FILL_1__1188_.gnd
rlabel nsubstratencontact 24 3848 24 3848 0 FILL_0__1537_.vdd
rlabel metal1 4 3602 36 3618 0 FILL_0__1537_.gnd
rlabel nsubstratencontact 144 3848 144 3848 0 FILL_0__1188_.vdd
rlabel metal1 124 3602 156 3618 0 FILL_0__1188_.gnd
rlabel metal1 44 3602 136 3618 0 _1537_.gnd
rlabel metal1 44 3842 136 3858 0 _1537_.vdd
rlabel metal2 113 3733 127 3747 0 _1537_.A
rlabel metal2 73 3733 87 3747 0 _1537_.B
rlabel metal2 93 3713 107 3727 0 _1537_.Y
rlabel metal1 164 3602 276 3618 0 _1188_.gnd
rlabel metal1 164 3842 276 3858 0 _1188_.vdd
rlabel metal2 253 3713 267 3727 0 _1188_.A
rlabel metal2 233 3733 247 3747 0 _1188_.B
rlabel metal2 213 3713 227 3727 0 _1188_.C
rlabel metal2 193 3733 207 3747 0 _1188_.Y
rlabel nsubstratencontact 304 3848 304 3848 0 FILL_1__1184_.vdd
rlabel metal1 284 3602 316 3618 0 FILL_1__1184_.gnd
rlabel nsubstratencontact 284 3848 284 3848 0 FILL_0__1184_.vdd
rlabel metal1 264 3602 296 3618 0 FILL_0__1184_.gnd
rlabel metal1 304 3842 496 3858 0 _1184_.vdd
rlabel metal2 453 3693 467 3707 0 _1184_.A
rlabel metal2 413 3713 427 3727 0 _1184_.B
rlabel metal2 393 3693 407 3707 0 _1184_.C
rlabel metal2 353 3713 367 3727 0 _1184_.Y
rlabel metal1 304 3602 496 3618 0 _1184_.gnd
rlabel nsubstratencontact 524 3848 524 3848 0 FILL_1__1366_.vdd
rlabel metal1 504 3602 536 3618 0 FILL_1__1366_.gnd
rlabel nsubstratencontact 504 3848 504 3848 0 FILL_0__1366_.vdd
rlabel metal1 484 3602 516 3618 0 FILL_0__1366_.gnd
rlabel nsubstratencontact 664 3848 664 3848 0 FILL_1__1365_.vdd
rlabel metal1 644 3602 676 3618 0 FILL_1__1365_.gnd
rlabel nsubstratencontact 644 3848 644 3848 0 FILL_0__1365_.vdd
rlabel metal1 624 3602 656 3618 0 FILL_0__1365_.gnd
rlabel metal1 524 3602 636 3618 0 _1366_.gnd
rlabel metal1 524 3842 636 3858 0 _1366_.vdd
rlabel metal2 613 3693 627 3707 0 _1366_.A
rlabel metal2 593 3713 607 3727 0 _1366_.B
rlabel metal2 553 3713 567 3727 0 _1366_.C
rlabel metal2 573 3693 587 3707 0 _1366_.Y
rlabel nsubstratencontact 776 3848 776 3848 0 FILL_1__1521_.vdd
rlabel metal1 764 3602 796 3618 0 FILL_1__1521_.gnd
rlabel nsubstratencontact 756 3848 756 3848 0 FILL_0__1521_.vdd
rlabel metal1 744 3602 776 3618 0 FILL_0__1521_.gnd
rlabel metal1 784 3602 896 3618 0 _1521_.gnd
rlabel metal1 784 3842 896 3858 0 _1521_.vdd
rlabel metal2 793 3693 807 3707 0 _1521_.A
rlabel metal2 813 3713 827 3727 0 _1521_.B
rlabel metal2 853 3713 867 3727 0 _1521_.C
rlabel metal2 833 3693 847 3707 0 _1521_.Y
rlabel metal1 664 3602 756 3618 0 _1365_.gnd
rlabel metal1 664 3842 756 3858 0 _1365_.vdd
rlabel metal2 733 3733 747 3747 0 _1365_.A
rlabel metal2 693 3733 707 3747 0 _1365_.B
rlabel metal2 713 3713 727 3727 0 _1365_.Y
rlabel nsubstratencontact 944 3848 944 3848 0 FILL_2__1520_.vdd
rlabel metal1 924 3602 956 3618 0 FILL_2__1520_.gnd
rlabel nsubstratencontact 924 3848 924 3848 0 FILL_1__1520_.vdd
rlabel metal1 904 3602 936 3618 0 FILL_1__1520_.gnd
rlabel nsubstratencontact 904 3848 904 3848 0 FILL_0__1520_.vdd
rlabel metal1 884 3602 916 3618 0 FILL_0__1520_.gnd
rlabel metal1 944 3602 1076 3618 0 _1520_.gnd
rlabel metal1 944 3842 1076 3858 0 _1520_.vdd
rlabel metal2 1053 3693 1067 3707 0 _1520_.A
rlabel metal2 1033 3713 1047 3727 0 _1520_.B
rlabel metal2 973 3693 987 3707 0 _1520_.C
rlabel metal2 993 3713 1007 3727 0 _1520_.D
rlabel metal2 1013 3693 1027 3707 0 _1520_.Y
rlabel nsubstratencontact 1096 3848 1096 3848 0 FILL_1__1475_.vdd
rlabel metal1 1084 3602 1116 3618 0 FILL_1__1475_.gnd
rlabel nsubstratencontact 1076 3848 1076 3848 0 FILL_0__1475_.vdd
rlabel metal1 1064 3602 1096 3618 0 FILL_0__1475_.gnd
rlabel metal1 1104 3602 1196 3618 0 _1475_.gnd
rlabel metal1 1104 3842 1196 3858 0 _1475_.vdd
rlabel metal2 1113 3733 1127 3747 0 _1475_.A
rlabel metal2 1153 3733 1167 3747 0 _1475_.B
rlabel metal2 1133 3713 1147 3727 0 _1475_.Y
rlabel nsubstratencontact 1216 3848 1216 3848 0 FILL_1__1526_.vdd
rlabel metal1 1204 3602 1236 3618 0 FILL_1__1526_.gnd
rlabel nsubstratencontact 1196 3848 1196 3848 0 FILL_0__1526_.vdd
rlabel metal1 1184 3602 1216 3618 0 FILL_0__1526_.gnd
rlabel metal1 1224 3602 1336 3618 0 _1526_.gnd
rlabel metal1 1224 3842 1336 3858 0 _1526_.vdd
rlabel metal2 1233 3713 1247 3727 0 _1526_.A
rlabel metal2 1253 3733 1267 3747 0 _1526_.B
rlabel metal2 1273 3713 1287 3727 0 _1526_.C
rlabel metal2 1293 3733 1307 3747 0 _1526_.Y
rlabel nsubstratencontact 1356 3848 1356 3848 0 FILL_1__1476_.vdd
rlabel metal1 1344 3602 1376 3618 0 FILL_1__1476_.gnd
rlabel nsubstratencontact 1336 3848 1336 3848 0 FILL_0__1476_.vdd
rlabel metal1 1324 3602 1356 3618 0 FILL_0__1476_.gnd
rlabel metal1 1364 3602 1476 3618 0 _1476_.gnd
rlabel metal1 1364 3842 1476 3858 0 _1476_.vdd
rlabel metal2 1373 3713 1387 3727 0 _1476_.A
rlabel metal2 1393 3673 1407 3687 0 _1476_.B
rlabel metal2 1413 3713 1427 3727 0 _1476_.C
rlabel metal2 1433 3693 1447 3707 0 _1476_.Y
rlabel nsubstratencontact 1496 3848 1496 3848 0 FILL_1__1478_.vdd
rlabel metal1 1484 3602 1516 3618 0 FILL_1__1478_.gnd
rlabel nsubstratencontact 1476 3848 1476 3848 0 FILL_0__1478_.vdd
rlabel metal1 1464 3602 1496 3618 0 FILL_0__1478_.gnd
rlabel metal1 1504 3602 1616 3618 0 _1478_.gnd
rlabel metal1 1504 3842 1616 3858 0 _1478_.vdd
rlabel metal2 1513 3693 1527 3707 0 _1478_.A
rlabel metal2 1533 3713 1547 3727 0 _1478_.B
rlabel metal2 1573 3713 1587 3727 0 _1478_.C
rlabel metal2 1553 3693 1567 3707 0 _1478_.Y
rlabel nsubstratencontact 1636 3848 1636 3848 0 FILL_1__1423_.vdd
rlabel metal1 1624 3602 1656 3618 0 FILL_1__1423_.gnd
rlabel nsubstratencontact 1616 3848 1616 3848 0 FILL_0__1423_.vdd
rlabel metal1 1604 3602 1636 3618 0 FILL_0__1423_.gnd
rlabel nsubstratencontact 1744 3848 1744 3848 0 FILL_1__1479_.vdd
rlabel metal1 1724 3602 1756 3618 0 FILL_1__1479_.gnd
rlabel nsubstratencontact 1724 3848 1724 3848 0 FILL_0__1479_.vdd
rlabel metal1 1704 3602 1736 3618 0 FILL_0__1479_.gnd
rlabel metal1 1744 3602 1836 3618 0 _1479_.gnd
rlabel metal1 1744 3842 1836 3858 0 _1479_.vdd
rlabel metal2 1813 3733 1827 3747 0 _1479_.A
rlabel metal2 1773 3733 1787 3747 0 _1479_.B
rlabel metal2 1793 3713 1807 3727 0 _1479_.Y
rlabel metal1 1644 3602 1716 3618 0 _1423_.gnd
rlabel metal1 1644 3842 1716 3858 0 _1423_.vdd
rlabel metal2 1653 3673 1667 3687 0 _1423_.A
rlabel metal2 1673 3713 1687 3727 0 _1423_.Y
rlabel nsubstratencontact 1856 3848 1856 3848 0 FILL_1__1424_.vdd
rlabel metal1 1844 3602 1876 3618 0 FILL_1__1424_.gnd
rlabel nsubstratencontact 1836 3848 1836 3848 0 FILL_0__1424_.vdd
rlabel metal1 1824 3602 1856 3618 0 FILL_0__1424_.gnd
rlabel metal1 1864 3602 1956 3618 0 _1424_.gnd
rlabel metal1 1864 3842 1956 3858 0 _1424_.vdd
rlabel metal2 1873 3733 1887 3747 0 _1424_.A
rlabel metal2 1913 3733 1927 3747 0 _1424_.B
rlabel metal2 1893 3713 1907 3727 0 _1424_.Y
rlabel nsubstratencontact 1976 3848 1976 3848 0 FILL_1__1425_.vdd
rlabel metal1 1964 3602 1996 3618 0 FILL_1__1425_.gnd
rlabel nsubstratencontact 1956 3848 1956 3848 0 FILL_0__1425_.vdd
rlabel metal1 1944 3602 1976 3618 0 FILL_0__1425_.gnd
rlabel metal1 1984 3602 2096 3618 0 _1425_.gnd
rlabel metal1 1984 3842 2096 3858 0 _1425_.vdd
rlabel metal2 1993 3673 2007 3687 0 _1425_.A
rlabel metal2 2013 3693 2027 3707 0 _1425_.B
rlabel metal2 2053 3713 2067 3727 0 _1425_.Y
rlabel nsubstratencontact 2116 3848 2116 3848 0 FILL_1__1426_.vdd
rlabel metal1 2104 3602 2136 3618 0 FILL_1__1426_.gnd
rlabel nsubstratencontact 2096 3848 2096 3848 0 FILL_0__1426_.vdd
rlabel metal1 2084 3602 2116 3618 0 FILL_0__1426_.gnd
rlabel metal1 2124 3602 2216 3618 0 _1426_.gnd
rlabel metal1 2124 3842 2216 3858 0 _1426_.vdd
rlabel metal2 2133 3733 2147 3747 0 _1426_.A
rlabel metal2 2173 3733 2187 3747 0 _1426_.B
rlabel metal2 2153 3713 2167 3727 0 _1426_.Y
rlabel nsubstratencontact 2236 3848 2236 3848 0 FILL_1__1078_.vdd
rlabel metal1 2224 3602 2256 3618 0 FILL_1__1078_.gnd
rlabel nsubstratencontact 2216 3848 2216 3848 0 FILL_0__1078_.vdd
rlabel metal1 2204 3602 2236 3618 0 FILL_0__1078_.gnd
rlabel metal1 2244 3602 2356 3618 0 _1078_.gnd
rlabel metal1 2244 3842 2356 3858 0 _1078_.vdd
rlabel metal2 2253 3713 2267 3727 0 _1078_.A
rlabel metal2 2273 3733 2287 3747 0 _1078_.B
rlabel metal2 2293 3713 2307 3727 0 _1078_.C
rlabel metal2 2313 3733 2327 3747 0 _1078_.Y
rlabel nsubstratencontact 2384 3848 2384 3848 0 FILL_1__1079_.vdd
rlabel metal1 2364 3602 2396 3618 0 FILL_1__1079_.gnd
rlabel nsubstratencontact 2364 3848 2364 3848 0 FILL_0__1079_.vdd
rlabel metal1 2344 3602 2376 3618 0 FILL_0__1079_.gnd
rlabel metal1 2384 3602 2496 3618 0 _1079_.gnd
rlabel metal1 2384 3842 2496 3858 0 _1079_.vdd
rlabel metal2 2473 3693 2487 3707 0 _1079_.A
rlabel metal2 2453 3713 2467 3727 0 _1079_.B
rlabel metal2 2413 3713 2427 3727 0 _1079_.C
rlabel metal2 2433 3693 2447 3707 0 _1079_.Y
rlabel nsubstratencontact 2516 3848 2516 3848 0 FILL_1__945_.vdd
rlabel metal1 2504 3602 2536 3618 0 FILL_1__945_.gnd
rlabel nsubstratencontact 2496 3848 2496 3848 0 FILL_0__945_.vdd
rlabel metal1 2484 3602 2516 3618 0 FILL_0__945_.gnd
rlabel metal1 2524 3602 2616 3618 0 _945_.gnd
rlabel metal1 2524 3842 2616 3858 0 _945_.vdd
rlabel metal2 2533 3733 2547 3747 0 _945_.A
rlabel metal2 2573 3733 2587 3747 0 _945_.B
rlabel metal2 2553 3713 2567 3727 0 _945_.Y
rlabel nsubstratencontact 2636 3848 2636 3848 0 FILL_1__1150_.vdd
rlabel metal1 2624 3602 2656 3618 0 FILL_1__1150_.gnd
rlabel nsubstratencontact 2616 3848 2616 3848 0 FILL_0__1150_.vdd
rlabel metal1 2604 3602 2636 3618 0 FILL_0__1150_.gnd
rlabel metal1 2644 3602 2756 3618 0 _1150_.gnd
rlabel metal1 2644 3842 2756 3858 0 _1150_.vdd
rlabel metal2 2653 3693 2667 3707 0 _1150_.A
rlabel metal2 2673 3713 2687 3727 0 _1150_.B
rlabel metal2 2713 3713 2727 3727 0 _1150_.C
rlabel metal2 2693 3693 2707 3707 0 _1150_.Y
rlabel nsubstratencontact 2784 3848 2784 3848 0 FILL_1__1151_.vdd
rlabel metal1 2764 3602 2796 3618 0 FILL_1__1151_.gnd
rlabel nsubstratencontact 2764 3848 2764 3848 0 FILL_0__1151_.vdd
rlabel metal1 2744 3602 2776 3618 0 FILL_0__1151_.gnd
rlabel nsubstratencontact 2884 3848 2884 3848 0 FILL_1__1152_.vdd
rlabel metal1 2864 3602 2896 3618 0 FILL_1__1152_.gnd
rlabel nsubstratencontact 2864 3848 2864 3848 0 FILL_0__1152_.vdd
rlabel metal1 2844 3602 2876 3618 0 FILL_0__1152_.gnd
rlabel metal1 2884 3602 2996 3618 0 _1152_.gnd
rlabel metal1 2884 3842 2996 3858 0 _1152_.vdd
rlabel metal2 2973 3693 2987 3707 0 _1152_.A
rlabel metal2 2953 3713 2967 3727 0 _1152_.B
rlabel metal2 2913 3713 2927 3727 0 _1152_.C
rlabel metal2 2933 3693 2947 3707 0 _1152_.Y
rlabel metal1 2784 3602 2856 3618 0 _1151_.gnd
rlabel metal1 2784 3842 2856 3858 0 _1151_.vdd
rlabel metal2 2833 3673 2847 3687 0 _1151_.A
rlabel metal2 2813 3713 2827 3727 0 _1151_.Y
rlabel nsubstratencontact 3016 3848 3016 3848 0 FILL_1__1171_.vdd
rlabel metal1 3004 3602 3036 3618 0 FILL_1__1171_.gnd
rlabel nsubstratencontact 2996 3848 2996 3848 0 FILL_0__1171_.vdd
rlabel metal1 2984 3602 3016 3618 0 FILL_0__1171_.gnd
rlabel metal1 3024 3602 3116 3618 0 _1171_.gnd
rlabel metal1 3024 3842 3116 3858 0 _1171_.vdd
rlabel metal2 3033 3733 3047 3747 0 _1171_.A
rlabel metal2 3073 3733 3087 3747 0 _1171_.B
rlabel metal2 3053 3713 3067 3727 0 _1171_.Y
rlabel nsubstratencontact 3164 3848 3164 3848 0 FILL_2__1148_.vdd
rlabel metal1 3144 3602 3176 3618 0 FILL_2__1148_.gnd
rlabel nsubstratencontact 3144 3848 3144 3848 0 FILL_1__1148_.vdd
rlabel metal1 3124 3602 3156 3618 0 FILL_1__1148_.gnd
rlabel nsubstratencontact 3124 3848 3124 3848 0 FILL_0__1148_.vdd
rlabel metal1 3104 3602 3136 3618 0 FILL_0__1148_.gnd
rlabel nsubstratencontact 3284 3848 3284 3848 0 FILL_1__1145_.vdd
rlabel metal1 3264 3602 3296 3618 0 FILL_1__1145_.gnd
rlabel nsubstratencontact 3264 3848 3264 3848 0 FILL_0__1145_.vdd
rlabel metal1 3244 3602 3276 3618 0 FILL_0__1145_.gnd
rlabel metal1 3164 3602 3256 3618 0 _1148_.gnd
rlabel metal1 3164 3842 3256 3858 0 _1148_.vdd
rlabel metal2 3233 3733 3247 3747 0 _1148_.A
rlabel metal2 3193 3733 3207 3747 0 _1148_.B
rlabel metal2 3213 3713 3227 3727 0 _1148_.Y
rlabel nsubstratencontact 3376 3848 3376 3848 0 FILL_1__1565_.vdd
rlabel metal1 3364 3602 3396 3618 0 FILL_1__1565_.gnd
rlabel nsubstratencontact 3356 3848 3356 3848 0 FILL_0__1565_.vdd
rlabel metal1 3344 3602 3376 3618 0 FILL_0__1565_.gnd
rlabel metal1 3384 3602 3496 3618 0 _1565_.gnd
rlabel metal1 3384 3842 3496 3858 0 _1565_.vdd
rlabel metal2 3393 3713 3407 3727 0 _1565_.A
rlabel metal2 3413 3733 3427 3747 0 _1565_.B
rlabel metal2 3433 3713 3447 3727 0 _1565_.C
rlabel metal2 3453 3733 3467 3747 0 _1565_.Y
rlabel metal1 3284 3602 3356 3618 0 _1145_.gnd
rlabel metal1 3284 3842 3356 3858 0 _1145_.vdd
rlabel metal2 3333 3673 3347 3687 0 _1145_.A
rlabel metal2 3313 3713 3327 3727 0 _1145_.Y
rlabel nsubstratencontact 3516 3848 3516 3848 0 FILL_1__1292_.vdd
rlabel metal1 3504 3602 3536 3618 0 FILL_1__1292_.gnd
rlabel nsubstratencontact 3496 3848 3496 3848 0 FILL_0__1292_.vdd
rlabel metal1 3484 3602 3516 3618 0 FILL_0__1292_.gnd
rlabel metal1 3524 3602 3596 3618 0 _1292_.gnd
rlabel metal1 3524 3842 3596 3858 0 _1292_.vdd
rlabel metal2 3533 3673 3547 3687 0 _1292_.A
rlabel metal2 3553 3713 3567 3727 0 _1292_.Y
rlabel nsubstratencontact 3756 3848 3756 3848 0 FILL_2__1291_.vdd
rlabel metal1 3744 3602 3776 3618 0 FILL_2__1291_.gnd
rlabel nsubstratencontact 3736 3848 3736 3848 0 FILL_1__1291_.vdd
rlabel metal1 3724 3602 3756 3618 0 FILL_1__1291_.gnd
rlabel nsubstratencontact 3624 3848 3624 3848 0 FILL_1__925_.vdd
rlabel metal1 3604 3602 3636 3618 0 FILL_1__925_.gnd
rlabel nsubstratencontact 3716 3848 3716 3848 0 FILL_0__1291_.vdd
rlabel metal1 3704 3602 3736 3618 0 FILL_0__1291_.gnd
rlabel nsubstratencontact 3604 3848 3604 3848 0 FILL_0__925_.vdd
rlabel metal1 3584 3602 3616 3618 0 FILL_0__925_.gnd
rlabel metal1 3764 3602 3856 3618 0 _1291_.gnd
rlabel metal1 3764 3842 3856 3858 0 _1291_.vdd
rlabel metal2 3773 3733 3787 3747 0 _1291_.A
rlabel metal2 3813 3733 3827 3747 0 _1291_.B
rlabel metal2 3793 3713 3807 3727 0 _1291_.Y
rlabel metal1 3624 3602 3716 3618 0 _925_.gnd
rlabel metal1 3624 3842 3716 3858 0 _925_.vdd
rlabel metal2 3653 3693 3667 3707 0 _925_.B
rlabel metal2 3693 3693 3707 3707 0 _925_.A
rlabel metal2 3673 3673 3687 3687 0 _925_.Y
rlabel nsubstratencontact 3876 3848 3876 3848 0 FILL_1__1077_.vdd
rlabel metal1 3864 3602 3896 3618 0 FILL_1__1077_.gnd
rlabel nsubstratencontact 3984 3848 3984 3848 0 FILL_1__951_.vdd
rlabel metal1 3964 3602 3996 3618 0 FILL_1__951_.gnd
rlabel nsubstratencontact 3856 3848 3856 3848 0 FILL_0__1077_.vdd
rlabel metal1 3844 3602 3876 3618 0 FILL_0__1077_.gnd
rlabel nsubstratencontact 3964 3848 3964 3848 0 FILL_0__951_.vdd
rlabel metal1 3944 3602 3976 3618 0 FILL_0__951_.gnd
rlabel metal1 3884 3602 3956 3618 0 _1077_.gnd
rlabel metal1 3884 3842 3956 3858 0 _1077_.vdd
rlabel metal2 3893 3673 3907 3687 0 _1077_.A
rlabel metal2 3913 3713 3927 3727 0 _1077_.Y
rlabel metal1 3984 3602 4056 3618 0 _951_.gnd
rlabel metal1 3984 3842 4056 3858 0 _951_.vdd
rlabel metal2 4033 3673 4047 3687 0 _951_.A
rlabel metal2 4013 3713 4027 3727 0 _951_.Y
rlabel metal1 4044 3602 4296 3618 0 _1672_.gnd
rlabel metal1 4044 3842 4296 3858 0 _1672_.vdd
rlabel metal2 4193 3693 4207 3707 0 _1672_.D
rlabel metal2 4153 3693 4167 3707 0 _1672_.CLK
rlabel metal2 4073 3693 4087 3707 0 _1672_.Q
rlabel metal1 4484 3602 4576 3618 0 _1493_.gnd
rlabel metal1 4484 3842 4576 3858 0 _1493_.vdd
rlabel metal2 4493 3733 4507 3747 0 _1493_.A
rlabel metal2 4533 3733 4547 3747 0 _1493_.B
rlabel metal2 4513 3713 4527 3727 0 _1493_.Y
rlabel metal1 4324 3602 4456 3618 0 _1548_.gnd
rlabel metal1 4324 3842 4456 3858 0 _1548_.vdd
rlabel metal2 4433 3693 4447 3707 0 _1548_.A
rlabel metal2 4413 3713 4427 3727 0 _1548_.B
rlabel metal2 4353 3693 4367 3707 0 _1548_.C
rlabel metal2 4393 3693 4407 3707 0 _1548_.Y
rlabel metal2 4373 3713 4387 3727 0 _1548_.D
rlabel nsubstratencontact 4456 3848 4456 3848 0 FILL_0__1493_.vdd
rlabel metal1 4444 3602 4476 3618 0 FILL_0__1493_.gnd
rlabel nsubstratencontact 4304 3848 4304 3848 0 FILL_0__1548_.vdd
rlabel metal1 4284 3602 4316 3618 0 FILL_0__1548_.gnd
rlabel nsubstratencontact 4476 3848 4476 3848 0 FILL_1__1493_.vdd
rlabel metal1 4464 3602 4496 3618 0 FILL_1__1493_.gnd
rlabel nsubstratencontact 4324 3848 4324 3848 0 FILL_1__1548_.vdd
rlabel metal1 4304 3602 4336 3618 0 FILL_1__1548_.gnd
rlabel nsubstratencontact 4596 3848 4596 3848 0 FILL_1__1197_.vdd
rlabel metal1 4584 3602 4616 3618 0 FILL_1__1197_.gnd
rlabel nsubstratencontact 4576 3848 4576 3848 0 FILL_0__1197_.vdd
rlabel metal1 4564 3602 4596 3618 0 FILL_0__1197_.gnd
rlabel metal1 4604 3602 4696 3618 0 _1197_.gnd
rlabel metal1 4604 3842 4696 3858 0 _1197_.vdd
rlabel metal2 4653 3693 4667 3707 0 _1197_.B
rlabel metal2 4613 3693 4627 3707 0 _1197_.A
rlabel metal2 4633 3673 4647 3687 0 _1197_.Y
rlabel nsubstratencontact 4716 3848 4716 3848 0 FILL_1__1645_.vdd
rlabel metal1 4704 3602 4736 3618 0 FILL_1__1645_.gnd
rlabel nsubstratencontact 4696 3848 4696 3848 0 FILL_0__1645_.vdd
rlabel metal1 4684 3602 4716 3618 0 FILL_0__1645_.gnd
rlabel metal1 4724 3602 4836 3618 0 _1645_.gnd
rlabel metal1 4724 3842 4836 3858 0 _1645_.vdd
rlabel metal2 4733 3693 4747 3707 0 _1645_.A
rlabel metal2 4753 3713 4767 3727 0 _1645_.B
rlabel metal2 4793 3713 4807 3727 0 _1645_.C
rlabel metal2 4773 3693 4787 3707 0 _1645_.Y
rlabel nsubstratencontact 4856 3848 4856 3848 0 FILL_1__1326_.vdd
rlabel metal1 4844 3602 4876 3618 0 FILL_1__1326_.gnd
rlabel nsubstratencontact 4836 3848 4836 3848 0 FILL_0__1326_.vdd
rlabel metal1 4824 3602 4856 3618 0 FILL_0__1326_.gnd
rlabel metal1 4864 3602 4936 3618 0 _1326_.gnd
rlabel metal1 4864 3842 4936 3858 0 _1326_.vdd
rlabel metal2 4873 3713 4887 3727 0 _1326_.A
rlabel metal2 4893 3693 4907 3707 0 _1326_.Y
rlabel nsubstratencontact 4984 3848 4984 3848 0 FILL_2__1644_.vdd
rlabel metal1 4964 3602 4996 3618 0 FILL_2__1644_.gnd
rlabel nsubstratencontact 4964 3848 4964 3848 0 FILL_1__1644_.vdd
rlabel metal1 4944 3602 4976 3618 0 FILL_1__1644_.gnd
rlabel nsubstratencontact 4944 3848 4944 3848 0 FILL_0__1644_.vdd
rlabel metal1 4924 3602 4956 3618 0 FILL_0__1644_.gnd
rlabel metal1 4984 3602 5076 3618 0 _1644_.gnd
rlabel metal1 4984 3842 5076 3858 0 _1644_.vdd
rlabel metal2 5053 3733 5067 3747 0 _1644_.A
rlabel metal2 5013 3733 5027 3747 0 _1644_.B
rlabel metal2 5033 3713 5047 3727 0 _1644_.Y
rlabel metal1 5104 3602 5176 3618 0 _1196_.gnd
rlabel metal1 5104 3842 5176 3858 0 _1196_.vdd
rlabel metal2 5113 3673 5127 3687 0 _1196_.A
rlabel metal2 5133 3713 5147 3727 0 _1196_.Y
rlabel metal1 5404 3602 5656 3618 0 _1654_.gnd
rlabel metal1 5404 3842 5656 3858 0 _1654_.vdd
rlabel metal2 5553 3693 5567 3707 0 _1654_.D
rlabel metal2 5513 3693 5527 3707 0 _1654_.CLK
rlabel metal2 5433 3693 5447 3707 0 _1654_.Q
rlabel metal1 5204 3602 5416 3618 0 CLKBUF1_insert2.gnd
rlabel metal1 5204 3842 5416 3858 0 CLKBUF1_insert2.vdd
rlabel metal2 5373 3713 5387 3727 0 CLKBUF1_insert2.A
rlabel metal2 5233 3713 5247 3727 0 CLKBUF1_insert2.Y
rlabel nsubstratencontact 5076 3848 5076 3848 0 FILL_0__1196_.vdd
rlabel metal1 5064 3602 5096 3618 0 FILL_0__1196_.gnd
rlabel nsubstratencontact 5184 3848 5184 3848 0 FILL_0_CLKBUF1_insert2.vdd
rlabel metal1 5164 3602 5196 3618 0 FILL_0_CLKBUF1_insert2.gnd
rlabel nsubstratencontact 5096 3848 5096 3848 0 FILL_1__1196_.vdd
rlabel metal1 5084 3602 5116 3618 0 FILL_1__1196_.gnd
rlabel nsubstratencontact 5204 3848 5204 3848 0 FILL_1_CLKBUF1_insert2.vdd
rlabel metal1 5184 3602 5216 3618 0 FILL_1_CLKBUF1_insert2.gnd
rlabel metal1 5684 3602 5776 3618 0 _1636_.gnd
rlabel metal1 5684 3842 5776 3858 0 _1636_.vdd
rlabel metal2 5753 3733 5767 3747 0 _1636_.A
rlabel metal2 5713 3733 5727 3747 0 _1636_.B
rlabel metal2 5733 3713 5747 3727 0 _1636_.Y
rlabel nsubstratencontact 5776 3848 5776 3848 0 FILL86550x54150.vdd
rlabel metal1 5764 3602 5796 3618 0 FILL86550x54150.gnd
rlabel nsubstratencontact 5796 3848 5796 3848 0 FILL86850x54150.vdd
rlabel metal1 5784 3602 5816 3618 0 FILL86850x54150.gnd
rlabel nsubstratencontact 5664 3848 5664 3848 0 FILL_0__1636_.vdd
rlabel metal1 5644 3602 5676 3618 0 FILL_0__1636_.gnd
rlabel nsubstratencontact 5684 3848 5684 3848 0 FILL_1__1636_.vdd
rlabel metal1 5664 3602 5696 3618 0 FILL_1__1636_.gnd
rlabel nsubstratencontact 136 3852 136 3852 0 FILL_1__1011_.vdd
rlabel metal1 124 4082 156 4098 0 FILL_1__1011_.gnd
rlabel nsubstratencontact 44 3852 44 3852 0 FILL_1__965_.vdd
rlabel metal1 24 4082 56 4098 0 FILL_1__965_.gnd
rlabel nsubstratencontact 116 3852 116 3852 0 FILL_0__1011_.vdd
rlabel metal1 104 4082 136 4098 0 FILL_0__1011_.gnd
rlabel nsubstratencontact 24 3852 24 3852 0 FILL_0__965_.vdd
rlabel metal1 4 4082 36 4098 0 FILL_0__965_.gnd
rlabel metal1 44 4082 116 4098 0 _965_.gnd
rlabel metal1 44 3842 116 3858 0 _965_.vdd
rlabel metal2 93 4013 107 4027 0 _965_.A
rlabel metal2 73 3973 87 3987 0 _965_.Y
rlabel nsubstratencontact 156 3852 156 3852 0 FILL_2__1011_.vdd
rlabel metal1 144 4082 176 4098 0 FILL_2__1011_.gnd
rlabel metal1 164 4082 276 4098 0 _1011_.gnd
rlabel metal1 164 3842 276 3858 0 _1011_.vdd
rlabel metal2 173 3993 187 4007 0 _1011_.A
rlabel metal2 193 3973 207 3987 0 _1011_.B
rlabel metal2 233 3973 247 3987 0 _1011_.C
rlabel metal2 213 3993 227 4007 0 _1011_.Y
rlabel nsubstratencontact 304 3852 304 3852 0 FILL_1__968_.vdd
rlabel metal1 284 4082 316 4098 0 FILL_1__968_.gnd
rlabel nsubstratencontact 376 3852 376 3852 0 FILL_0__999_.vdd
rlabel metal1 364 4082 396 4098 0 FILL_0__999_.gnd
rlabel nsubstratencontact 284 3852 284 3852 0 FILL_0__968_.vdd
rlabel metal1 264 4082 296 4098 0 FILL_0__968_.gnd
rlabel metal1 304 4082 376 4098 0 _968_.gnd
rlabel metal1 304 3842 376 3858 0 _968_.vdd
rlabel metal2 353 4013 367 4027 0 _968_.A
rlabel metal2 333 3973 347 3987 0 _968_.Y
rlabel nsubstratencontact 416 3852 416 3852 0 FILL_2__999_.vdd
rlabel metal1 404 4082 436 4098 0 FILL_2__999_.gnd
rlabel nsubstratencontact 396 3852 396 3852 0 FILL_1__999_.vdd
rlabel metal1 384 4082 416 4098 0 FILL_1__999_.gnd
rlabel metal1 424 4082 536 4098 0 _999_.gnd
rlabel metal1 424 3842 536 3858 0 _999_.vdd
rlabel metal2 433 3973 447 3987 0 _999_.A
rlabel metal2 453 4013 467 4027 0 _999_.B
rlabel metal2 473 3973 487 3987 0 _999_.C
rlabel metal2 493 3993 507 4007 0 _999_.Y
rlabel nsubstratencontact 564 3852 564 3852 0 FILL_1__967_.vdd
rlabel metal1 544 4082 576 4098 0 FILL_1__967_.gnd
rlabel nsubstratencontact 544 3852 544 3852 0 FILL_0__967_.vdd
rlabel metal1 524 4082 556 4098 0 FILL_0__967_.gnd
rlabel metal1 564 4082 656 4098 0 _967_.gnd
rlabel metal1 564 3842 656 3858 0 _967_.vdd
rlabel metal2 593 3993 607 4007 0 _967_.B
rlabel metal2 633 3993 647 4007 0 _967_.A
rlabel metal2 613 4013 627 4027 0 _967_.Y
rlabel nsubstratencontact 704 3852 704 3852 0 FILL_2__1180_.vdd
rlabel metal1 684 4082 716 4098 0 FILL_2__1180_.gnd
rlabel nsubstratencontact 684 3852 684 3852 0 FILL_1__1180_.vdd
rlabel metal1 664 4082 696 4098 0 FILL_1__1180_.gnd
rlabel nsubstratencontact 664 3852 664 3852 0 FILL_0__1180_.vdd
rlabel metal1 644 4082 676 4098 0 FILL_0__1180_.gnd
rlabel metal1 704 4082 776 4098 0 _1180_.gnd
rlabel metal1 704 3842 776 3858 0 _1180_.vdd
rlabel metal2 753 4013 767 4027 0 _1180_.A
rlabel metal2 733 3973 747 3987 0 _1180_.Y
rlabel nsubstratencontact 796 3852 796 3852 0 FILL_1__1181_.vdd
rlabel metal1 784 4082 816 4098 0 FILL_1__1181_.gnd
rlabel nsubstratencontact 776 3852 776 3852 0 FILL_0__1181_.vdd
rlabel metal1 764 4082 796 4098 0 FILL_0__1181_.gnd
rlabel metal1 804 4082 916 4098 0 _1181_.gnd
rlabel metal1 804 3842 916 3858 0 _1181_.vdd
rlabel metal2 813 3993 827 4007 0 _1181_.A
rlabel metal2 833 3973 847 3987 0 _1181_.B
rlabel metal2 873 3973 887 3987 0 _1181_.C
rlabel metal2 853 3993 867 4007 0 _1181_.Y
rlabel nsubstratencontact 936 3852 936 3852 0 FILL_1__1168_.vdd
rlabel metal1 924 4082 956 4098 0 FILL_1__1168_.gnd
rlabel nsubstratencontact 1016 3852 1016 3852 0 FILL_0__1170_.vdd
rlabel metal1 1004 4082 1036 4098 0 FILL_0__1170_.gnd
rlabel nsubstratencontact 916 3852 916 3852 0 FILL_0__1168_.vdd
rlabel metal1 904 4082 936 4098 0 FILL_0__1168_.gnd
rlabel metal1 944 4082 1016 4098 0 _1168_.gnd
rlabel metal1 944 3842 1016 3858 0 _1168_.vdd
rlabel metal2 953 4013 967 4027 0 _1168_.A
rlabel metal2 973 3973 987 3987 0 _1168_.Y
rlabel nsubstratencontact 1036 3852 1036 3852 0 FILL_1__1170_.vdd
rlabel metal1 1024 4082 1056 4098 0 FILL_1__1170_.gnd
rlabel nsubstratencontact 1156 3852 1156 3852 0 FILL_0__1525_.vdd
rlabel metal1 1144 4082 1176 4098 0 FILL_0__1525_.gnd
rlabel metal1 1044 4082 1156 4098 0 _1170_.gnd
rlabel metal1 1044 3842 1156 3858 0 _1170_.vdd
rlabel metal2 1053 3973 1067 3987 0 _1170_.A
rlabel metal2 1073 3953 1087 3967 0 _1170_.B
rlabel metal2 1093 3973 1107 3987 0 _1170_.C
rlabel metal2 1113 3953 1127 3967 0 _1170_.Y
rlabel nsubstratencontact 1176 3852 1176 3852 0 FILL_1__1525_.vdd
rlabel metal1 1164 4082 1196 4098 0 FILL_1__1525_.gnd
rlabel nsubstratencontact 1316 3852 1316 3852 0 FILL_0__1422_.vdd
rlabel metal1 1304 4082 1336 4098 0 FILL_0__1422_.gnd
rlabel metal1 1184 4082 1316 4098 0 _1525_.gnd
rlabel metal1 1184 3842 1316 3858 0 _1525_.vdd
rlabel metal2 1193 3993 1207 4007 0 _1525_.A
rlabel metal2 1213 3973 1227 3987 0 _1525_.B
rlabel metal2 1273 3993 1287 4007 0 _1525_.C
rlabel metal2 1253 3973 1267 3987 0 _1525_.D
rlabel metal2 1233 3993 1247 4007 0 _1525_.Y
rlabel nsubstratencontact 1356 3852 1356 3852 0 FILL_2__1422_.vdd
rlabel metal1 1344 4082 1376 4098 0 FILL_2__1422_.gnd
rlabel nsubstratencontact 1336 3852 1336 3852 0 FILL_1__1422_.vdd
rlabel metal1 1324 4082 1356 4098 0 FILL_1__1422_.gnd
rlabel nsubstratencontact 1464 3852 1464 3852 0 FILL_0__1473_.vdd
rlabel metal1 1444 4082 1476 4098 0 FILL_0__1473_.gnd
rlabel metal1 1364 4082 1456 4098 0 _1422_.gnd
rlabel metal1 1364 3842 1456 3858 0 _1422_.vdd
rlabel metal2 1373 3953 1387 3967 0 _1422_.A
rlabel metal2 1413 3953 1427 3967 0 _1422_.B
rlabel metal2 1393 3973 1407 3987 0 _1422_.Y
rlabel nsubstratencontact 1484 3852 1484 3852 0 FILL_1__1473_.vdd
rlabel metal1 1464 4082 1496 4098 0 FILL_1__1473_.gnd
rlabel metal1 1484 4082 1556 4098 0 _1473_.gnd
rlabel metal1 1484 3842 1556 3858 0 _1473_.vdd
rlabel metal2 1533 4013 1547 4027 0 _1473_.A
rlabel metal2 1513 3973 1527 3987 0 _1473_.Y
rlabel nsubstratencontact 1584 3852 1584 3852 0 FILL_1__1524_.vdd
rlabel metal1 1564 4082 1596 4098 0 FILL_1__1524_.gnd
rlabel nsubstratencontact 1564 3852 1564 3852 0 FILL_0__1524_.vdd
rlabel metal1 1544 4082 1576 4098 0 FILL_0__1524_.gnd
rlabel metal1 1584 4082 1676 4098 0 _1524_.gnd
rlabel metal1 1584 3842 1676 3858 0 _1524_.vdd
rlabel metal2 1613 3993 1627 4007 0 _1524_.B
rlabel metal2 1653 3993 1667 4007 0 _1524_.A
rlabel metal2 1633 4013 1647 4027 0 _1524_.Y
rlabel nsubstratencontact 1704 3852 1704 3852 0 FILL_1__1477_.vdd
rlabel metal1 1684 4082 1716 4098 0 FILL_1__1477_.gnd
rlabel nsubstratencontact 1684 3852 1684 3852 0 FILL_0__1477_.vdd
rlabel metal1 1664 4082 1696 4098 0 FILL_0__1477_.gnd
rlabel nsubstratencontact 1776 3852 1776 3852 0 FILL_0__1472_.vdd
rlabel metal1 1764 4082 1796 4098 0 FILL_0__1472_.gnd
rlabel metal1 1704 4082 1776 4098 0 _1477_.gnd
rlabel metal1 1704 3842 1776 3858 0 _1477_.vdd
rlabel metal2 1753 4013 1767 4027 0 _1477_.A
rlabel metal2 1733 3973 1747 3987 0 _1477_.Y
rlabel nsubstratencontact 1796 3852 1796 3852 0 FILL_1__1472_.vdd
rlabel metal1 1784 4082 1816 4098 0 FILL_1__1472_.gnd
rlabel metal1 1804 4082 1916 4098 0 _1472_.gnd
rlabel metal1 1804 3842 1916 3858 0 _1472_.vdd
rlabel metal2 1813 3973 1827 3987 0 _1472_.A
rlabel metal2 1833 3953 1847 3967 0 _1472_.B
rlabel metal2 1853 3973 1867 3987 0 _1472_.C
rlabel metal2 1873 3953 1887 3967 0 _1472_.Y
rlabel nsubstratencontact 1944 3852 1944 3852 0 FILL_1__963_.vdd
rlabel metal1 1924 4082 1956 4098 0 FILL_1__963_.gnd
rlabel nsubstratencontact 1924 3852 1924 3852 0 FILL_0__963_.vdd
rlabel metal1 1904 4082 1936 4098 0 FILL_0__963_.gnd
rlabel metal1 1944 4082 2056 4098 0 _963_.gnd
rlabel metal1 1944 3842 2056 3858 0 _963_.vdd
rlabel metal2 2033 3993 2047 4007 0 _963_.A
rlabel metal2 2013 3973 2027 3987 0 _963_.B
rlabel metal2 1973 3973 1987 3987 0 _963_.C
rlabel metal2 1993 3993 2007 4007 0 _963_.Y
rlabel nsubstratencontact 2104 3852 2104 3852 0 FILL_2__959_.vdd
rlabel metal1 2084 4082 2116 4098 0 FILL_2__959_.gnd
rlabel nsubstratencontact 2084 3852 2084 3852 0 FILL_1__959_.vdd
rlabel metal1 2064 4082 2096 4098 0 FILL_1__959_.gnd
rlabel nsubstratencontact 2064 3852 2064 3852 0 FILL_0__959_.vdd
rlabel metal1 2044 4082 2076 4098 0 FILL_0__959_.gnd
rlabel metal1 2104 4082 2216 4098 0 _959_.gnd
rlabel metal1 2104 3842 2216 3858 0 _959_.vdd
rlabel metal2 2193 3973 2207 3987 0 _959_.A
rlabel metal2 2173 3953 2187 3967 0 _959_.B
rlabel metal2 2153 3973 2167 3987 0 _959_.C
rlabel metal2 2133 3953 2147 3967 0 _959_.Y
rlabel nsubstratencontact 2236 3852 2236 3852 0 FILL_1__928_.vdd
rlabel metal1 2224 4082 2256 4098 0 FILL_1__928_.gnd
rlabel nsubstratencontact 2216 3852 2216 3852 0 FILL_0__928_.vdd
rlabel metal1 2204 4082 2236 4098 0 FILL_0__928_.gnd
rlabel metal1 2244 4082 2356 4098 0 _928_.gnd
rlabel metal1 2244 3842 2356 3858 0 _928_.vdd
rlabel metal2 2253 3973 2267 3987 0 _928_.A
rlabel metal2 2273 3953 2287 3967 0 _928_.B
rlabel metal2 2293 3973 2307 3987 0 _928_.C
rlabel metal2 2313 3953 2327 3967 0 _928_.Y
rlabel nsubstratencontact 2384 3852 2384 3852 0 FILL_1__935_.vdd
rlabel metal1 2364 4082 2396 4098 0 FILL_1__935_.gnd
rlabel nsubstratencontact 2364 3852 2364 3852 0 FILL_0__935_.vdd
rlabel metal1 2344 4082 2376 4098 0 FILL_0__935_.gnd
rlabel metal1 2384 4082 2496 4098 0 _935_.gnd
rlabel metal1 2384 3842 2496 3858 0 _935_.vdd
rlabel metal2 2473 3993 2487 4007 0 _935_.A
rlabel metal2 2453 3973 2467 3987 0 _935_.B
rlabel metal2 2413 3973 2427 3987 0 _935_.C
rlabel metal2 2433 3993 2447 4007 0 _935_.Y
rlabel nsubstratencontact 2524 3852 2524 3852 0 FILL_1__934_.vdd
rlabel metal1 2504 4082 2536 4098 0 FILL_1__934_.gnd
rlabel nsubstratencontact 2504 3852 2504 3852 0 FILL_0__934_.vdd
rlabel metal1 2484 4082 2516 4098 0 FILL_0__934_.gnd
rlabel metal1 2524 4082 2616 4098 0 _934_.gnd
rlabel metal1 2524 3842 2616 3858 0 _934_.vdd
rlabel metal2 2593 3953 2607 3967 0 _934_.A
rlabel metal2 2553 3953 2567 3967 0 _934_.B
rlabel metal2 2573 3973 2587 3987 0 _934_.Y
rlabel nsubstratencontact 2636 3852 2636 3852 0 FILL_1__962_.vdd
rlabel metal1 2624 4082 2656 4098 0 FILL_1__962_.gnd
rlabel nsubstratencontact 2616 3852 2616 3852 0 FILL_0__962_.vdd
rlabel metal1 2604 4082 2636 4098 0 FILL_0__962_.gnd
rlabel metal1 2644 4082 2736 4098 0 _962_.gnd
rlabel metal1 2644 3842 2736 3858 0 _962_.vdd
rlabel metal2 2653 3953 2667 3967 0 _962_.A
rlabel metal2 2693 3953 2707 3967 0 _962_.B
rlabel metal2 2673 3973 2687 3987 0 _962_.Y
rlabel nsubstratencontact 2756 3852 2756 3852 0 FILL_1__1144_.vdd
rlabel metal1 2744 4082 2776 4098 0 FILL_1__1144_.gnd
rlabel nsubstratencontact 2736 3852 2736 3852 0 FILL_0__1144_.vdd
rlabel metal1 2724 4082 2756 4098 0 FILL_0__1144_.gnd
rlabel metal1 2764 4082 2876 4098 0 _1144_.gnd
rlabel metal1 2764 3842 2876 3858 0 _1144_.vdd
rlabel metal2 2773 3973 2787 3987 0 _1144_.A
rlabel metal2 2793 3953 2807 3967 0 _1144_.B
rlabel metal2 2813 3973 2827 3987 0 _1144_.C
rlabel metal2 2833 3953 2847 3967 0 _1144_.Y
rlabel nsubstratencontact 2896 3852 2896 3852 0 FILL_1__1146_.vdd
rlabel metal1 2884 4082 2916 4098 0 FILL_1__1146_.gnd
rlabel nsubstratencontact 2876 3852 2876 3852 0 FILL_0__1146_.vdd
rlabel metal1 2864 4082 2896 4098 0 FILL_0__1146_.gnd
rlabel nsubstratencontact 3044 3852 3044 3852 0 FILL_1__1147_.vdd
rlabel metal1 3024 4082 3056 4098 0 FILL_1__1147_.gnd
rlabel nsubstratencontact 3024 3852 3024 3852 0 FILL_0__1147_.vdd
rlabel metal1 3004 4082 3036 4098 0 FILL_0__1147_.gnd
rlabel metal1 2904 4082 3016 4098 0 _1146_.gnd
rlabel metal1 2904 3842 3016 3858 0 _1146_.vdd
rlabel metal2 2913 3973 2927 3987 0 _1146_.A
rlabel metal2 2933 3953 2947 3967 0 _1146_.B
rlabel metal2 2953 3973 2967 3987 0 _1146_.C
rlabel metal2 2973 3953 2987 3967 0 _1146_.Y
rlabel nsubstratencontact 3144 3852 3144 3852 0 FILL_1__1586_.vdd
rlabel metal1 3124 4082 3156 4098 0 FILL_1__1586_.gnd
rlabel nsubstratencontact 3124 3852 3124 3852 0 FILL_0__1586_.vdd
rlabel metal1 3104 4082 3136 4098 0 FILL_0__1586_.gnd
rlabel metal1 3144 4082 3256 4098 0 _1586_.gnd
rlabel metal1 3144 3842 3256 3858 0 _1586_.vdd
rlabel metal2 3233 3973 3247 3987 0 _1586_.A
rlabel metal2 3213 3953 3227 3967 0 _1586_.B
rlabel metal2 3193 3973 3207 3987 0 _1586_.C
rlabel metal2 3173 3953 3187 3967 0 _1586_.Y
rlabel metal1 3044 4082 3116 4098 0 _1147_.gnd
rlabel metal1 3044 3842 3116 3858 0 _1147_.vdd
rlabel metal2 3093 4013 3107 4027 0 _1147_.A
rlabel metal2 3073 3973 3087 3987 0 _1147_.Y
rlabel nsubstratencontact 3284 3852 3284 3852 0 FILL_1__1581_.vdd
rlabel metal1 3264 4082 3296 4098 0 FILL_1__1581_.gnd
rlabel nsubstratencontact 3264 3852 3264 3852 0 FILL_0__1581_.vdd
rlabel metal1 3244 4082 3276 4098 0 FILL_0__1581_.gnd
rlabel nsubstratencontact 3384 3852 3384 3852 0 FILL_1__1582_.vdd
rlabel metal1 3364 4082 3396 4098 0 FILL_1__1582_.gnd
rlabel nsubstratencontact 3364 3852 3364 3852 0 FILL_0__1582_.vdd
rlabel metal1 3344 4082 3376 4098 0 FILL_0__1582_.gnd
rlabel metal1 3384 4082 3496 4098 0 _1582_.gnd
rlabel metal1 3384 3842 3496 3858 0 _1582_.vdd
rlabel metal2 3473 3993 3487 4007 0 _1582_.A
rlabel metal2 3453 3973 3467 3987 0 _1582_.B
rlabel metal2 3413 3973 3427 3987 0 _1582_.C
rlabel metal2 3433 3993 3447 4007 0 _1582_.Y
rlabel metal1 3284 4082 3356 4098 0 _1581_.gnd
rlabel metal1 3284 3842 3356 3858 0 _1581_.vdd
rlabel metal2 3333 4013 3347 4027 0 _1581_.A
rlabel metal2 3313 3973 3327 3987 0 _1581_.Y
rlabel nsubstratencontact 3516 3852 3516 3852 0 FILL_1__1580_.vdd
rlabel metal1 3504 4082 3536 4098 0 FILL_1__1580_.gnd
rlabel nsubstratencontact 3496 3852 3496 3852 0 FILL_0__1580_.vdd
rlabel metal1 3484 4082 3516 4098 0 FILL_0__1580_.gnd
rlabel metal1 3524 4082 3616 4098 0 _1580_.gnd
rlabel metal1 3524 3842 3616 3858 0 _1580_.vdd
rlabel metal2 3533 3953 3547 3967 0 _1580_.A
rlabel metal2 3573 3953 3587 3967 0 _1580_.B
rlabel metal2 3553 3973 3567 3987 0 _1580_.Y
rlabel nsubstratencontact 3644 3852 3644 3852 0 FILL_1__1578_.vdd
rlabel metal1 3624 4082 3656 4098 0 FILL_1__1578_.gnd
rlabel nsubstratencontact 3624 3852 3624 3852 0 FILL_0__1578_.vdd
rlabel metal1 3604 4082 3636 4098 0 FILL_0__1578_.gnd
rlabel metal1 3644 4082 3756 4098 0 _1578_.gnd
rlabel metal1 3644 3842 3756 3858 0 _1578_.vdd
rlabel metal2 3733 4013 3747 4027 0 _1578_.A
rlabel metal2 3713 3993 3727 4007 0 _1578_.B
rlabel metal2 3673 3973 3687 3987 0 _1578_.Y
rlabel nsubstratencontact 3796 3852 3796 3852 0 FILL_2__1579_.vdd
rlabel metal1 3784 4082 3816 4098 0 FILL_2__1579_.gnd
rlabel nsubstratencontact 3776 3852 3776 3852 0 FILL_1__1579_.vdd
rlabel metal1 3764 4082 3796 4098 0 FILL_1__1579_.gnd
rlabel nsubstratencontact 3756 3852 3756 3852 0 FILL_0__1579_.vdd
rlabel metal1 3744 4082 3776 4098 0 FILL_0__1579_.gnd
rlabel nsubstratencontact 3924 3852 3924 3852 0 FILL_1__1589_.vdd
rlabel metal1 3904 4082 3936 4098 0 FILL_1__1589_.gnd
rlabel nsubstratencontact 3904 3852 3904 3852 0 FILL_0__1589_.vdd
rlabel metal1 3884 4082 3916 4098 0 FILL_0__1589_.gnd
rlabel metal1 3804 4082 3896 4098 0 _1579_.gnd
rlabel metal1 3804 3842 3896 3858 0 _1579_.vdd
rlabel metal2 3813 3953 3827 3967 0 _1579_.A
rlabel metal2 3853 3953 3867 3967 0 _1579_.B
rlabel metal2 3833 3973 3847 3987 0 _1579_.Y
rlabel nsubstratencontact 4044 3852 4044 3852 0 FILL_0__1577_.vdd
rlabel metal1 4024 4082 4056 4098 0 FILL_0__1577_.gnd
rlabel metal1 3924 4082 4036 4098 0 _1589_.gnd
rlabel metal1 3924 3842 4036 3858 0 _1589_.vdd
rlabel metal2 4013 3993 4027 4007 0 _1589_.A
rlabel metal2 3993 3973 4007 3987 0 _1589_.B
rlabel metal2 3953 3973 3967 3987 0 _1589_.C
rlabel metal2 3973 3993 3987 4007 0 _1589_.Y
rlabel nsubstratencontact 4064 3852 4064 3852 0 FILL_1__1577_.vdd
rlabel metal1 4044 4082 4076 4098 0 FILL_1__1577_.gnd
rlabel nsubstratencontact 4176 3852 4176 3852 0 FILL_0__1547_.vdd
rlabel metal1 4164 4082 4196 4098 0 FILL_0__1547_.gnd
rlabel metal1 4064 4082 4176 4098 0 _1577_.gnd
rlabel metal1 4064 3842 4176 3858 0 _1577_.vdd
rlabel metal2 4153 3973 4167 3987 0 _1577_.A
rlabel metal2 4133 4013 4147 4027 0 _1577_.B
rlabel metal2 4113 3973 4127 3987 0 _1577_.C
rlabel metal2 4093 3993 4107 4007 0 _1577_.Y
rlabel nsubstratencontact 4196 3852 4196 3852 0 FILL_1__1547_.vdd
rlabel metal1 4184 4082 4216 4098 0 FILL_1__1547_.gnd
rlabel nsubstratencontact 4296 3852 4296 3852 0 FILL_0__1549_.vdd
rlabel metal1 4284 4082 4316 4098 0 FILL_0__1549_.gnd
rlabel metal1 4204 4082 4296 4098 0 _1547_.gnd
rlabel metal1 4204 3842 4296 3858 0 _1547_.vdd
rlabel metal2 4213 3953 4227 3967 0 _1547_.A
rlabel metal2 4253 3953 4267 3967 0 _1547_.B
rlabel metal2 4233 3973 4247 3987 0 _1547_.Y
rlabel nsubstratencontact 4316 3852 4316 3852 0 FILL_1__1549_.vdd
rlabel metal1 4304 4082 4336 4098 0 FILL_1__1549_.gnd
rlabel metal1 4324 4082 4436 4098 0 _1549_.gnd
rlabel metal1 4324 3842 4436 3858 0 _1549_.vdd
rlabel metal2 4333 3993 4347 4007 0 _1549_.A
rlabel metal2 4353 3973 4367 3987 0 _1549_.B
rlabel metal2 4393 3973 4407 3987 0 _1549_.C
rlabel metal2 4373 3993 4387 4007 0 _1549_.Y
rlabel nsubstratencontact 4456 3852 4456 3852 0 FILL_1__1498_.vdd
rlabel metal1 4444 4082 4476 4098 0 FILL_1__1498_.gnd
rlabel nsubstratencontact 4436 3852 4436 3852 0 FILL_0__1498_.vdd
rlabel metal1 4424 4082 4456 4098 0 FILL_0__1498_.gnd
rlabel metal1 4464 4082 4576 4098 0 _1498_.gnd
rlabel metal1 4464 3842 4576 3858 0 _1498_.vdd
rlabel metal2 4473 3993 4487 4007 0 _1498_.A
rlabel metal2 4493 3973 4507 3987 0 _1498_.B
rlabel metal2 4533 3973 4547 3987 0 _1498_.C
rlabel metal2 4513 3993 4527 4007 0 _1498_.Y
rlabel nsubstratencontact 4596 3852 4596 3852 0 FILL_1__1497_.vdd
rlabel metal1 4584 4082 4616 4098 0 FILL_1__1497_.gnd
rlabel nsubstratencontact 4576 3852 4576 3852 0 FILL_0__1497_.vdd
rlabel metal1 4564 4082 4596 4098 0 FILL_0__1497_.gnd
rlabel metal1 4604 4082 4716 4098 0 _1497_.gnd
rlabel metal1 4604 3842 4716 3858 0 _1497_.vdd
rlabel metal2 4613 4013 4627 4027 0 _1497_.A
rlabel metal2 4633 3993 4647 4007 0 _1497_.B
rlabel metal2 4673 3973 4687 3987 0 _1497_.Y
rlabel nsubstratencontact 4744 3852 4744 3852 0 FILL_1__1499_.vdd
rlabel metal1 4724 4082 4756 4098 0 FILL_1__1499_.gnd
rlabel nsubstratencontact 4724 3852 4724 3852 0 FILL_0__1499_.vdd
rlabel metal1 4704 4082 4736 4098 0 FILL_0__1499_.gnd
rlabel metal1 4744 4082 4836 4098 0 _1499_.gnd
rlabel metal1 4744 3842 4836 3858 0 _1499_.vdd
rlabel metal2 4813 3953 4827 3967 0 _1499_.A
rlabel metal2 4773 3953 4787 3967 0 _1499_.B
rlabel metal2 4793 3973 4807 3987 0 _1499_.Y
rlabel nsubstratencontact 4856 3852 4856 3852 0 FILL_1__1504_.vdd
rlabel metal1 4844 4082 4876 4098 0 FILL_1__1504_.gnd
rlabel nsubstratencontact 4836 3852 4836 3852 0 FILL_0__1504_.vdd
rlabel metal1 4824 4082 4856 4098 0 FILL_0__1504_.gnd
rlabel metal1 4864 4082 4976 4098 0 _1504_.gnd
rlabel metal1 4864 3842 4976 3858 0 _1504_.vdd
rlabel metal2 4873 3973 4887 3987 0 _1504_.A
rlabel metal2 4893 3953 4907 3967 0 _1504_.B
rlabel metal2 4913 3973 4927 3987 0 _1504_.C
rlabel metal2 4933 3953 4947 3967 0 _1504_.Y
rlabel nsubstratencontact 4996 3852 4996 3852 0 FILL_1__1503_.vdd
rlabel metal1 4984 4082 5016 4098 0 FILL_1__1503_.gnd
rlabel nsubstratencontact 4976 3852 4976 3852 0 FILL_0__1503_.vdd
rlabel metal1 4964 4082 4996 4098 0 FILL_0__1503_.gnd
rlabel metal1 5004 4082 5076 4098 0 _1503_.gnd
rlabel metal1 5004 3842 5076 3858 0 _1503_.vdd
rlabel metal2 5013 4013 5027 4027 0 _1503_.A
rlabel metal2 5033 3973 5047 3987 0 _1503_.Y
rlabel metal1 5104 4082 5176 4098 0 _961_.gnd
rlabel metal1 5104 3842 5176 3858 0 _961_.vdd
rlabel metal2 5153 4013 5167 4027 0 _961_.A
rlabel metal2 5133 3973 5147 3987 0 _961_.Y
rlabel metal1 5164 4082 5416 4098 0 _1659_.gnd
rlabel metal1 5164 3842 5416 3858 0 _1659_.vdd
rlabel metal2 5313 3993 5327 4007 0 _1659_.D
rlabel metal2 5273 3993 5287 4007 0 _1659_.CLK
rlabel metal2 5193 3993 5207 4007 0 _1659_.Q
rlabel metal1 5404 4082 5656 4098 0 _1677_.gnd
rlabel metal1 5404 3842 5656 3858 0 _1677_.vdd
rlabel metal2 5553 3993 5567 4007 0 _1677_.D
rlabel metal2 5513 3993 5527 4007 0 _1677_.CLK
rlabel metal2 5433 3993 5447 4007 0 _1677_.Q
rlabel nsubstratencontact 5084 3852 5084 3852 0 FILL_0__961_.vdd
rlabel metal1 5064 4082 5096 4098 0 FILL_0__961_.gnd
rlabel nsubstratencontact 5104 3852 5104 3852 0 FILL_1__961_.vdd
rlabel metal1 5084 4082 5116 4098 0 FILL_1__961_.gnd
rlabel metal1 5684 4082 5796 4098 0 _1637_.gnd
rlabel metal1 5684 3842 5796 3858 0 _1637_.vdd
rlabel metal2 5693 3993 5707 4007 0 _1637_.A
rlabel metal2 5713 3973 5727 3987 0 _1637_.B
rlabel metal2 5753 3973 5767 3987 0 _1637_.C
rlabel metal2 5733 3993 5747 4007 0 _1637_.Y
rlabel nsubstratencontact 5804 3852 5804 3852 0 FILL86850x57750.vdd
rlabel metal1 5784 4082 5816 4098 0 FILL86850x57750.gnd
rlabel nsubstratencontact 5656 3852 5656 3852 0 FILL_0__1637_.vdd
rlabel metal1 5644 4082 5676 4098 0 FILL_0__1637_.gnd
rlabel nsubstratencontact 5676 3852 5676 3852 0 FILL_1__1637_.vdd
rlabel metal1 5664 4082 5696 4098 0 FILL_1__1637_.gnd
rlabel nsubstratencontact 64 4328 64 4328 0 FILL_2__972_.vdd
rlabel metal1 44 4082 76 4098 0 FILL_2__972_.gnd
rlabel nsubstratencontact 44 4328 44 4328 0 FILL_1__972_.vdd
rlabel metal1 24 4082 56 4098 0 FILL_1__972_.gnd
rlabel nsubstratencontact 24 4328 24 4328 0 FILL_0__972_.vdd
rlabel metal1 4 4082 36 4098 0 FILL_0__972_.gnd
rlabel metal1 64 4082 176 4098 0 _972_.gnd
rlabel metal1 64 4322 176 4338 0 _972_.vdd
rlabel metal2 153 4173 167 4187 0 _972_.A
rlabel metal2 133 4193 147 4207 0 _972_.B
rlabel metal2 93 4193 107 4207 0 _972_.C
rlabel metal2 113 4173 127 4187 0 _972_.Y
rlabel nsubstratencontact 204 4328 204 4328 0 FILL_1__969_.vdd
rlabel metal1 184 4082 216 4098 0 FILL_1__969_.gnd
rlabel nsubstratencontact 184 4328 184 4328 0 FILL_0__969_.vdd
rlabel metal1 164 4082 196 4098 0 FILL_0__969_.gnd
rlabel metal1 204 4082 316 4098 0 _969_.gnd
rlabel metal1 204 4322 316 4338 0 _969_.vdd
rlabel metal2 293 4173 307 4187 0 _969_.A
rlabel metal2 273 4193 287 4207 0 _969_.B
rlabel metal2 233 4193 247 4207 0 _969_.C
rlabel metal2 253 4173 267 4187 0 _969_.Y
rlabel nsubstratencontact 364 4328 364 4328 0 FILL_2__966_.vdd
rlabel metal1 344 4082 376 4098 0 FILL_2__966_.gnd
rlabel nsubstratencontact 344 4328 344 4328 0 FILL_1__966_.vdd
rlabel metal1 324 4082 356 4098 0 FILL_1__966_.gnd
rlabel nsubstratencontact 324 4328 324 4328 0 FILL_0__966_.vdd
rlabel metal1 304 4082 336 4098 0 FILL_0__966_.gnd
rlabel metal1 364 4082 476 4098 0 _966_.gnd
rlabel metal1 364 4322 476 4338 0 _966_.vdd
rlabel metal2 453 4193 467 4207 0 _966_.A
rlabel metal2 433 4213 447 4227 0 _966_.B
rlabel metal2 413 4193 427 4207 0 _966_.C
rlabel metal2 393 4213 407 4227 0 _966_.Y
rlabel nsubstratencontact 504 4328 504 4328 0 FILL_1__973_.vdd
rlabel metal1 484 4082 516 4098 0 FILL_1__973_.gnd
rlabel nsubstratencontact 484 4328 484 4328 0 FILL_0__973_.vdd
rlabel metal1 464 4082 496 4098 0 FILL_0__973_.gnd
rlabel metal1 504 4082 616 4098 0 _973_.gnd
rlabel metal1 504 4322 616 4338 0 _973_.vdd
rlabel metal2 593 4193 607 4207 0 _973_.A
rlabel metal2 573 4213 587 4227 0 _973_.B
rlabel metal2 553 4193 567 4207 0 _973_.C
rlabel metal2 533 4213 547 4227 0 _973_.Y
rlabel nsubstratencontact 644 4328 644 4328 0 FILL_1__960_.vdd
rlabel metal1 624 4082 656 4098 0 FILL_1__960_.gnd
rlabel nsubstratencontact 624 4328 624 4328 0 FILL_0__960_.vdd
rlabel metal1 604 4082 636 4098 0 FILL_0__960_.gnd
rlabel nsubstratencontact 764 4328 764 4328 0 FILL_0__1157_.vdd
rlabel metal1 744 4082 776 4098 0 FILL_0__1157_.gnd
rlabel metal1 644 4082 756 4098 0 _960_.gnd
rlabel metal1 644 4322 756 4338 0 _960_.vdd
rlabel metal2 733 4153 747 4167 0 _960_.A
rlabel metal2 713 4173 727 4187 0 _960_.B
rlabel metal2 673 4193 687 4207 0 _960_.Y
rlabel nsubstratencontact 784 4328 784 4328 0 FILL_1__1157_.vdd
rlabel metal1 764 4082 796 4098 0 FILL_1__1157_.gnd
rlabel metal1 784 4082 896 4098 0 _1157_.gnd
rlabel metal1 784 4322 896 4338 0 _1157_.vdd
rlabel metal2 873 4173 887 4187 0 _1157_.A
rlabel metal2 853 4193 867 4207 0 _1157_.B
rlabel metal2 813 4193 827 4207 0 _1157_.C
rlabel metal2 833 4173 847 4187 0 _1157_.Y
rlabel nsubstratencontact 916 4328 916 4328 0 FILL_1__1169_.vdd
rlabel metal1 904 4082 936 4098 0 FILL_1__1169_.gnd
rlabel nsubstratencontact 1024 4328 1024 4328 0 FILL_1__1156_.vdd
rlabel metal1 1004 4082 1036 4098 0 FILL_1__1156_.gnd
rlabel nsubstratencontact 896 4328 896 4328 0 FILL_0__1169_.vdd
rlabel metal1 884 4082 916 4098 0 FILL_0__1169_.gnd
rlabel nsubstratencontact 1004 4328 1004 4328 0 FILL_0__1156_.vdd
rlabel metal1 984 4082 1016 4098 0 FILL_0__1156_.gnd
rlabel metal1 924 4082 996 4098 0 _1169_.gnd
rlabel metal1 924 4322 996 4338 0 _1169_.vdd
rlabel metal2 933 4153 947 4167 0 _1169_.A
rlabel metal2 953 4193 967 4207 0 _1169_.Y
rlabel nsubstratencontact 1144 4328 1144 4328 0 FILL_0__1154_.vdd
rlabel metal1 1124 4082 1156 4098 0 FILL_0__1154_.gnd
rlabel metal1 1024 4082 1136 4098 0 _1156_.gnd
rlabel metal1 1024 4322 1136 4338 0 _1156_.vdd
rlabel metal2 1113 4193 1127 4207 0 _1156_.A
rlabel metal2 1093 4153 1107 4167 0 _1156_.B
rlabel metal2 1073 4193 1087 4207 0 _1156_.C
rlabel metal2 1053 4173 1067 4187 0 _1156_.Y
rlabel nsubstratencontact 1184 4328 1184 4328 0 FILL_2__1154_.vdd
rlabel metal1 1164 4082 1196 4098 0 FILL_2__1154_.gnd
rlabel nsubstratencontact 1164 4328 1164 4328 0 FILL_1__1154_.vdd
rlabel metal1 1144 4082 1176 4098 0 FILL_1__1154_.gnd
rlabel metal1 1184 4082 1296 4098 0 _1154_.gnd
rlabel metal1 1184 4322 1296 4338 0 _1154_.vdd
rlabel metal2 1273 4193 1287 4207 0 _1154_.A
rlabel metal2 1253 4213 1267 4227 0 _1154_.B
rlabel metal2 1233 4193 1247 4207 0 _1154_.C
rlabel metal2 1213 4213 1227 4227 0 _1154_.Y
rlabel nsubstratencontact 1324 4328 1324 4328 0 FILL_1__1517_.vdd
rlabel metal1 1304 4082 1336 4098 0 FILL_1__1517_.gnd
rlabel nsubstratencontact 1304 4328 1304 4328 0 FILL_0__1517_.vdd
rlabel metal1 1284 4082 1316 4098 0 FILL_0__1517_.gnd
rlabel metal1 1324 4082 1416 4098 0 _1517_.gnd
rlabel metal1 1324 4322 1416 4338 0 _1517_.vdd
rlabel metal2 1393 4213 1407 4227 0 _1517_.A
rlabel metal2 1353 4213 1367 4227 0 _1517_.B
rlabel metal2 1373 4193 1387 4207 0 _1517_.Y
rlabel nsubstratencontact 1444 4328 1444 4328 0 FILL_1__1155_.vdd
rlabel metal1 1424 4082 1456 4098 0 FILL_1__1155_.gnd
rlabel nsubstratencontact 1424 4328 1424 4328 0 FILL_0__1155_.vdd
rlabel metal1 1404 4082 1436 4098 0 FILL_0__1155_.gnd
rlabel metal1 1444 4082 1536 4098 0 _1155_.gnd
rlabel metal1 1444 4322 1536 4338 0 _1155_.vdd
rlabel metal2 1513 4213 1527 4227 0 _1155_.A
rlabel metal2 1473 4213 1487 4227 0 _1155_.B
rlabel metal2 1493 4193 1507 4207 0 _1155_.Y
rlabel nsubstratencontact 1564 4328 1564 4328 0 FILL_1__942_.vdd
rlabel metal1 1544 4082 1576 4098 0 FILL_1__942_.gnd
rlabel nsubstratencontact 1544 4328 1544 4328 0 FILL_0__942_.vdd
rlabel metal1 1524 4082 1556 4098 0 FILL_0__942_.gnd
rlabel metal1 1564 4082 1656 4098 0 _942_.gnd
rlabel metal1 1564 4322 1656 4338 0 _942_.vdd
rlabel metal2 1593 4173 1607 4187 0 _942_.B
rlabel metal2 1633 4173 1647 4187 0 _942_.A
rlabel metal2 1613 4153 1627 4167 0 _942_.Y
rlabel nsubstratencontact 1684 4328 1684 4328 0 FILL_1__964_.vdd
rlabel metal1 1664 4082 1696 4098 0 FILL_1__964_.gnd
rlabel nsubstratencontact 1664 4328 1664 4328 0 FILL_0__964_.vdd
rlabel metal1 1644 4082 1676 4098 0 FILL_0__964_.gnd
rlabel metal1 1684 4082 1796 4098 0 _964_.gnd
rlabel metal1 1684 4322 1796 4338 0 _964_.vdd
rlabel metal2 1773 4193 1787 4207 0 _964_.A
rlabel metal2 1753 4213 1767 4227 0 _964_.B
rlabel metal2 1733 4193 1747 4207 0 _964_.C
rlabel metal2 1713 4213 1727 4227 0 _964_.Y
rlabel nsubstratencontact 1824 4328 1824 4328 0 FILL_1__941_.vdd
rlabel metal1 1804 4082 1836 4098 0 FILL_1__941_.gnd
rlabel nsubstratencontact 1804 4328 1804 4328 0 FILL_0__941_.vdd
rlabel metal1 1784 4082 1816 4098 0 FILL_0__941_.gnd
rlabel metal1 1824 4082 1936 4098 0 _941_.gnd
rlabel metal1 1824 4322 1936 4338 0 _941_.vdd
rlabel metal2 1913 4193 1927 4207 0 _941_.A
rlabel metal2 1893 4213 1907 4227 0 _941_.B
rlabel metal2 1873 4193 1887 4207 0 _941_.C
rlabel metal2 1853 4213 1867 4227 0 _941_.Y
rlabel nsubstratencontact 1956 4328 1956 4328 0 FILL_1__958_.vdd
rlabel metal1 1944 4082 1976 4098 0 FILL_1__958_.gnd
rlabel nsubstratencontact 1936 4328 1936 4328 0 FILL_0__958_.vdd
rlabel metal1 1924 4082 1956 4098 0 FILL_0__958_.gnd
rlabel metal1 1964 4082 2076 4098 0 _958_.gnd
rlabel metal1 1964 4322 2076 4338 0 _958_.vdd
rlabel metal2 1973 4193 1987 4207 0 _958_.A
rlabel metal2 1993 4213 2007 4227 0 _958_.B
rlabel metal2 2013 4193 2027 4207 0 _958_.C
rlabel metal2 2033 4213 2047 4227 0 _958_.Y
rlabel nsubstratencontact 2096 4328 2096 4328 0 FILL_1__929_.vdd
rlabel metal1 2084 4082 2116 4098 0 FILL_1__929_.gnd
rlabel nsubstratencontact 2076 4328 2076 4328 0 FILL_0__929_.vdd
rlabel metal1 2064 4082 2096 4098 0 FILL_0__929_.gnd
rlabel metal1 2104 4082 2216 4098 0 _929_.gnd
rlabel metal1 2104 4322 2216 4338 0 _929_.vdd
rlabel metal2 2113 4193 2127 4207 0 _929_.A
rlabel metal2 2133 4213 2147 4227 0 _929_.B
rlabel metal2 2153 4193 2167 4207 0 _929_.C
rlabel metal2 2173 4213 2187 4227 0 _929_.Y
rlabel nsubstratencontact 2244 4328 2244 4328 0 FILL_1__930_.vdd
rlabel metal1 2224 4082 2256 4098 0 FILL_1__930_.gnd
rlabel nsubstratencontact 2224 4328 2224 4328 0 FILL_0__930_.vdd
rlabel metal1 2204 4082 2236 4098 0 FILL_0__930_.gnd
rlabel metal1 2244 4082 2336 4098 0 _930_.gnd
rlabel metal1 2244 4322 2336 4338 0 _930_.vdd
rlabel metal2 2273 4173 2287 4187 0 _930_.B
rlabel metal2 2313 4173 2327 4187 0 _930_.A
rlabel metal2 2293 4153 2307 4167 0 _930_.Y
rlabel nsubstratencontact 2384 4328 2384 4328 0 FILL_2__946_.vdd
rlabel metal1 2364 4082 2396 4098 0 FILL_2__946_.gnd
rlabel nsubstratencontact 2364 4328 2364 4328 0 FILL_1__946_.vdd
rlabel metal1 2344 4082 2376 4098 0 FILL_1__946_.gnd
rlabel nsubstratencontact 2344 4328 2344 4328 0 FILL_0__946_.vdd
rlabel metal1 2324 4082 2356 4098 0 FILL_0__946_.gnd
rlabel metal1 2384 4082 2496 4098 0 _946_.gnd
rlabel metal1 2384 4322 2496 4338 0 _946_.vdd
rlabel metal2 2473 4173 2487 4187 0 _946_.A
rlabel metal2 2453 4193 2467 4207 0 _946_.B
rlabel metal2 2413 4193 2427 4207 0 _946_.C
rlabel metal2 2433 4173 2447 4187 0 _946_.Y
rlabel nsubstratencontact 2524 4328 2524 4328 0 FILL_1__940_.vdd
rlabel metal1 2504 4082 2536 4098 0 FILL_1__940_.gnd
rlabel nsubstratencontact 2504 4328 2504 4328 0 FILL_0__940_.vdd
rlabel metal1 2484 4082 2516 4098 0 FILL_0__940_.gnd
rlabel nsubstratencontact 2544 4328 2544 4328 0 FILL_2__940_.vdd
rlabel metal1 2524 4082 2556 4098 0 FILL_2__940_.gnd
rlabel nsubstratencontact 2656 4328 2656 4328 0 FILL_0__1293_.vdd
rlabel metal1 2644 4082 2676 4098 0 FILL_0__1293_.gnd
rlabel metal1 2544 4082 2656 4098 0 _940_.gnd
rlabel metal1 2544 4322 2656 4338 0 _940_.vdd
rlabel metal2 2633 4193 2647 4207 0 _940_.A
rlabel metal2 2613 4213 2627 4227 0 _940_.B
rlabel metal2 2593 4193 2607 4207 0 _940_.C
rlabel metal2 2573 4213 2587 4227 0 _940_.Y
rlabel nsubstratencontact 2776 4328 2776 4328 0 FILL_1__1527_.vdd
rlabel metal1 2764 4082 2796 4098 0 FILL_1__1527_.gnd
rlabel nsubstratencontact 2676 4328 2676 4328 0 FILL_1__1293_.vdd
rlabel metal1 2664 4082 2696 4098 0 FILL_1__1293_.gnd
rlabel nsubstratencontact 2756 4328 2756 4328 0 FILL_0__1527_.vdd
rlabel metal1 2744 4082 2776 4098 0 FILL_0__1527_.gnd
rlabel metal1 2684 4082 2756 4098 0 _1293_.gnd
rlabel metal1 2684 4322 2756 4338 0 _1293_.vdd
rlabel metal2 2693 4153 2707 4167 0 _1293_.A
rlabel metal2 2713 4193 2727 4207 0 _1293_.Y
rlabel nsubstratencontact 2796 4328 2796 4328 0 FILL_2__1527_.vdd
rlabel metal1 2784 4082 2816 4098 0 FILL_2__1527_.gnd
rlabel metal1 2804 4082 2916 4098 0 _1527_.gnd
rlabel metal1 2804 4322 2916 4338 0 _1527_.vdd
rlabel metal2 2813 4193 2827 4207 0 _1527_.A
rlabel metal2 2833 4213 2847 4227 0 _1527_.B
rlabel metal2 2853 4193 2867 4207 0 _1527_.C
rlabel metal2 2873 4213 2887 4227 0 _1527_.Y
rlabel nsubstratencontact 2936 4328 2936 4328 0 FILL_1__1528_.vdd
rlabel metal1 2924 4082 2956 4098 0 FILL_1__1528_.gnd
rlabel nsubstratencontact 3036 4328 3036 4328 0 FILL_0__1574_.vdd
rlabel metal1 3024 4082 3056 4098 0 FILL_0__1574_.gnd
rlabel nsubstratencontact 2916 4328 2916 4328 0 FILL_0__1528_.vdd
rlabel metal1 2904 4082 2936 4098 0 FILL_0__1528_.gnd
rlabel metal1 2944 4082 3036 4098 0 _1528_.gnd
rlabel metal1 2944 4322 3036 4338 0 _1528_.vdd
rlabel metal2 2953 4213 2967 4227 0 _1528_.A
rlabel metal2 2993 4213 3007 4227 0 _1528_.B
rlabel metal2 2973 4193 2987 4207 0 _1528_.Y
rlabel nsubstratencontact 3056 4328 3056 4328 0 FILL_1__1574_.vdd
rlabel metal1 3044 4082 3076 4098 0 FILL_1__1574_.gnd
rlabel metal1 3064 4082 3176 4098 0 _1574_.gnd
rlabel metal1 3064 4322 3176 4338 0 _1574_.vdd
rlabel metal2 3073 4193 3087 4207 0 _1574_.A
rlabel metal2 3093 4153 3107 4167 0 _1574_.B
rlabel metal2 3113 4193 3127 4207 0 _1574_.C
rlabel metal2 3133 4173 3147 4187 0 _1574_.Y
rlabel nsubstratencontact 3196 4328 3196 4328 0 FILL_1__1562_.vdd
rlabel metal1 3184 4082 3216 4098 0 FILL_1__1562_.gnd
rlabel nsubstratencontact 3176 4328 3176 4328 0 FILL_0__1562_.vdd
rlabel metal1 3164 4082 3196 4098 0 FILL_0__1562_.gnd
rlabel metal1 3204 4082 3316 4098 0 _1562_.gnd
rlabel metal1 3204 4322 3316 4338 0 _1562_.vdd
rlabel metal2 3213 4193 3227 4207 0 _1562_.A
rlabel metal2 3233 4153 3247 4167 0 _1562_.B
rlabel metal2 3253 4193 3267 4207 0 _1562_.C
rlabel metal2 3273 4173 3287 4187 0 _1562_.Y
rlabel nsubstratencontact 3336 4328 3336 4328 0 FILL_1__1564_.vdd
rlabel metal1 3324 4082 3356 4098 0 FILL_1__1564_.gnd
rlabel nsubstratencontact 3316 4328 3316 4328 0 FILL_0__1564_.vdd
rlabel metal1 3304 4082 3336 4098 0 FILL_0__1564_.gnd
rlabel metal1 3344 4082 3456 4098 0 _1564_.gnd
rlabel metal1 3344 4322 3456 4338 0 _1564_.vdd
rlabel metal2 3353 4173 3367 4187 0 _1564_.A
rlabel metal2 3373 4193 3387 4207 0 _1564_.B
rlabel metal2 3413 4193 3427 4207 0 _1564_.C
rlabel metal2 3393 4173 3407 4187 0 _1564_.Y
rlabel nsubstratencontact 3496 4328 3496 4328 0 FILL_2__1585_.vdd
rlabel metal1 3484 4082 3516 4098 0 FILL_2__1585_.gnd
rlabel nsubstratencontact 3476 4328 3476 4328 0 FILL_1__1585_.vdd
rlabel metal1 3464 4082 3496 4098 0 FILL_1__1585_.gnd
rlabel nsubstratencontact 3456 4328 3456 4328 0 FILL_0__1585_.vdd
rlabel metal1 3444 4082 3476 4098 0 FILL_0__1585_.gnd
rlabel metal1 3504 4082 3576 4098 0 _1585_.gnd
rlabel metal1 3504 4322 3576 4338 0 _1585_.vdd
rlabel metal2 3513 4153 3527 4167 0 _1585_.A
rlabel metal2 3533 4193 3547 4207 0 _1585_.Y
rlabel nsubstratencontact 3596 4328 3596 4328 0 FILL_1__1308_.vdd
rlabel metal1 3584 4082 3616 4098 0 FILL_1__1308_.gnd
rlabel nsubstratencontact 3576 4328 3576 4328 0 FILL_0__1308_.vdd
rlabel metal1 3564 4082 3596 4098 0 FILL_0__1308_.gnd
rlabel metal1 3604 4082 3716 4098 0 _1308_.gnd
rlabel metal1 3604 4322 3716 4338 0 _1308_.vdd
rlabel metal2 3613 4193 3627 4207 0 _1308_.A
rlabel metal2 3633 4213 3647 4227 0 _1308_.B
rlabel metal2 3653 4193 3667 4207 0 _1308_.C
rlabel metal2 3673 4213 3687 4227 0 _1308_.Y
rlabel nsubstratencontact 3736 4328 3736 4328 0 FILL_1__1313_.vdd
rlabel metal1 3724 4082 3756 4098 0 FILL_1__1313_.gnd
rlabel nsubstratencontact 3716 4328 3716 4328 0 FILL_0__1313_.vdd
rlabel metal1 3704 4082 3736 4098 0 FILL_0__1313_.gnd
rlabel metal1 3744 4082 3856 4098 0 _1313_.gnd
rlabel metal1 3744 4322 3856 4338 0 _1313_.vdd
rlabel metal2 3753 4193 3767 4207 0 _1313_.A
rlabel metal2 3773 4213 3787 4227 0 _1313_.B
rlabel metal2 3793 4193 3807 4207 0 _1313_.C
rlabel metal2 3813 4213 3827 4227 0 _1313_.Y
rlabel nsubstratencontact 3884 4328 3884 4328 0 FILL_1__922_.vdd
rlabel metal1 3864 4082 3896 4098 0 FILL_1__922_.gnd
rlabel nsubstratencontact 3864 4328 3864 4328 0 FILL_0__922_.vdd
rlabel metal1 3844 4082 3876 4098 0 FILL_0__922_.gnd
rlabel metal1 3884 4082 3976 4098 0 _922_.gnd
rlabel metal1 3884 4322 3976 4338 0 _922_.vdd
rlabel metal2 3953 4213 3967 4227 0 _922_.A
rlabel metal2 3913 4213 3927 4227 0 _922_.B
rlabel metal2 3933 4193 3947 4207 0 _922_.Y
rlabel nsubstratencontact 4024 4328 4024 4328 0 FILL_2__1494_.vdd
rlabel metal1 4004 4082 4036 4098 0 FILL_2__1494_.gnd
rlabel nsubstratencontact 4004 4328 4004 4328 0 FILL_1__1494_.vdd
rlabel metal1 3984 4082 4016 4098 0 FILL_1__1494_.gnd
rlabel nsubstratencontact 3984 4328 3984 4328 0 FILL_0__1494_.vdd
rlabel metal1 3964 4082 3996 4098 0 FILL_0__1494_.gnd
rlabel metal1 4024 4082 4116 4098 0 _1494_.gnd
rlabel metal1 4024 4322 4116 4338 0 _1494_.vdd
rlabel metal2 4093 4213 4107 4227 0 _1494_.A
rlabel metal2 4053 4213 4067 4227 0 _1494_.B
rlabel metal2 4073 4193 4087 4207 0 _1494_.Y
rlabel nsubstratencontact 4144 4328 4144 4328 0 FILL_1__1450_.vdd
rlabel metal1 4124 4082 4156 4098 0 FILL_1__1450_.gnd
rlabel nsubstratencontact 4124 4328 4124 4328 0 FILL_0__1450_.vdd
rlabel metal1 4104 4082 4136 4098 0 FILL_0__1450_.gnd
rlabel metal1 4144 4082 4236 4098 0 _1450_.gnd
rlabel metal1 4144 4322 4236 4338 0 _1450_.vdd
rlabel metal2 4213 4213 4227 4227 0 _1450_.A
rlabel metal2 4173 4213 4187 4227 0 _1450_.B
rlabel metal2 4193 4193 4207 4207 0 _1450_.Y
rlabel nsubstratencontact 4264 4328 4264 4328 0 FILL_1__1495_.vdd
rlabel metal1 4244 4082 4276 4098 0 FILL_1__1495_.gnd
rlabel nsubstratencontact 4244 4328 4244 4328 0 FILL_0__1495_.vdd
rlabel metal1 4224 4082 4256 4098 0 FILL_0__1495_.gnd
rlabel metal1 4264 4082 4376 4098 0 _1495_.gnd
rlabel metal1 4264 4322 4376 4338 0 _1495_.vdd
rlabel metal2 4353 4173 4367 4187 0 _1495_.A
rlabel metal2 4333 4193 4347 4207 0 _1495_.B
rlabel metal2 4293 4193 4307 4207 0 _1495_.C
rlabel metal2 4313 4173 4327 4187 0 _1495_.Y
rlabel nsubstratencontact 4396 4328 4396 4328 0 FILL_1__1451_.vdd
rlabel metal1 4384 4082 4416 4098 0 FILL_1__1451_.gnd
rlabel nsubstratencontact 4376 4328 4376 4328 0 FILL_0__1451_.vdd
rlabel metal1 4364 4082 4396 4098 0 FILL_0__1451_.gnd
rlabel metal1 4404 4082 4516 4098 0 _1451_.gnd
rlabel metal1 4404 4322 4516 4338 0 _1451_.vdd
rlabel metal2 4413 4153 4427 4167 0 _1451_.A
rlabel metal2 4433 4173 4447 4187 0 _1451_.B
rlabel metal2 4473 4193 4487 4207 0 _1451_.Y
rlabel nsubstratencontact 4544 4328 4544 4328 0 FILL_1__1496_.vdd
rlabel metal1 4524 4082 4556 4098 0 FILL_1__1496_.gnd
rlabel nsubstratencontact 4524 4328 4524 4328 0 FILL_0__1496_.vdd
rlabel metal1 4504 4082 4536 4098 0 FILL_0__1496_.gnd
rlabel metal1 4544 4082 4656 4098 0 _1496_.gnd
rlabel metal1 4544 4322 4656 4338 0 _1496_.vdd
rlabel metal2 4633 4173 4647 4187 0 _1496_.A
rlabel metal2 4613 4193 4627 4207 0 _1496_.B
rlabel metal2 4573 4193 4587 4207 0 _1496_.C
rlabel metal2 4593 4173 4607 4187 0 _1496_.Y
rlabel nsubstratencontact 4676 4328 4676 4328 0 FILL_1__1500_.vdd
rlabel metal1 4664 4082 4696 4098 0 FILL_1__1500_.gnd
rlabel nsubstratencontact 4656 4328 4656 4328 0 FILL_0__1500_.vdd
rlabel metal1 4644 4082 4676 4098 0 FILL_0__1500_.gnd
rlabel nsubstratencontact 4696 4328 4696 4328 0 FILL_2__1500_.vdd
rlabel metal1 4684 4082 4716 4098 0 FILL_2__1500_.gnd
rlabel metal1 4704 4082 4816 4098 0 _1500_.gnd
rlabel metal1 4704 4322 4816 4338 0 _1500_.vdd
rlabel metal2 4713 4173 4727 4187 0 _1500_.A
rlabel metal2 4733 4193 4747 4207 0 _1500_.B
rlabel metal2 4773 4193 4787 4207 0 _1500_.C
rlabel metal2 4753 4173 4767 4187 0 _1500_.Y
rlabel nsubstratencontact 4836 4328 4836 4328 0 FILL_1__1545_.vdd
rlabel metal1 4824 4082 4856 4098 0 FILL_1__1545_.gnd
rlabel nsubstratencontact 4816 4328 4816 4328 0 FILL_0__1545_.vdd
rlabel metal1 4804 4082 4836 4098 0 FILL_0__1545_.gnd
rlabel metal1 4844 4082 4936 4098 0 _1545_.gnd
rlabel metal1 4844 4322 4936 4338 0 _1545_.vdd
rlabel metal2 4893 4173 4907 4187 0 _1545_.B
rlabel metal2 4853 4173 4867 4187 0 _1545_.A
rlabel metal2 4873 4153 4887 4167 0 _1545_.Y
rlabel nsubstratencontact 5056 4328 5056 4328 0 FILL_1__1546_.vdd
rlabel metal1 5044 4082 5076 4098 0 FILL_1__1546_.gnd
rlabel nsubstratencontact 4956 4328 4956 4328 0 FILL_1__1544_.vdd
rlabel metal1 4944 4082 4976 4098 0 FILL_1__1544_.gnd
rlabel nsubstratencontact 5036 4328 5036 4328 0 FILL_0__1546_.vdd
rlabel metal1 5024 4082 5056 4098 0 FILL_0__1546_.gnd
rlabel nsubstratencontact 4936 4328 4936 4328 0 FILL_0__1544_.vdd
rlabel metal1 4924 4082 4956 4098 0 FILL_0__1544_.gnd
rlabel metal1 4964 4082 5036 4098 0 _1544_.gnd
rlabel metal1 4964 4322 5036 4338 0 _1544_.vdd
rlabel metal2 4973 4153 4987 4167 0 _1544_.A
rlabel metal2 4993 4193 5007 4207 0 _1544_.Y
rlabel nsubstratencontact 5076 4328 5076 4328 0 FILL_2__1546_.vdd
rlabel metal1 5064 4082 5096 4098 0 FILL_2__1546_.gnd
rlabel metal1 5084 4082 5196 4098 0 _1546_.gnd
rlabel metal1 5084 4322 5196 4338 0 _1546_.vdd
rlabel metal2 5093 4193 5107 4207 0 _1546_.A
rlabel metal2 5113 4153 5127 4167 0 _1546_.B
rlabel metal2 5133 4193 5147 4207 0 _1546_.C
rlabel metal2 5153 4173 5167 4187 0 _1546_.Y
rlabel nsubstratencontact 5216 4328 5216 4328 0 FILL_1__1576_.vdd
rlabel metal1 5204 4082 5236 4098 0 FILL_1__1576_.gnd
rlabel nsubstratencontact 5196 4328 5196 4328 0 FILL_0__1576_.vdd
rlabel metal1 5184 4082 5216 4098 0 FILL_0__1576_.gnd
rlabel metal1 5224 4082 5336 4098 0 _1576_.gnd
rlabel metal1 5224 4322 5336 4338 0 _1576_.vdd
rlabel metal2 5233 4173 5247 4187 0 _1576_.A
rlabel metal2 5253 4193 5267 4207 0 _1576_.B
rlabel metal2 5293 4193 5307 4207 0 _1576_.C
rlabel metal2 5273 4173 5287 4187 0 _1576_.Y
rlabel nsubstratencontact 5356 4328 5356 4328 0 FILL_1__1615_.vdd
rlabel metal1 5344 4082 5376 4098 0 FILL_1__1615_.gnd
rlabel nsubstratencontact 5436 4328 5436 4328 0 FILL_0__1617_.vdd
rlabel metal1 5424 4082 5456 4098 0 FILL_0__1617_.gnd
rlabel nsubstratencontact 5336 4328 5336 4328 0 FILL_0__1615_.vdd
rlabel metal1 5324 4082 5356 4098 0 FILL_0__1615_.gnd
rlabel metal1 5364 4082 5436 4098 0 _1615_.gnd
rlabel metal1 5364 4322 5436 4338 0 _1615_.vdd
rlabel metal2 5373 4153 5387 4167 0 _1615_.A
rlabel metal2 5393 4193 5407 4207 0 _1615_.Y
rlabel nsubstratencontact 5456 4328 5456 4328 0 FILL_1__1617_.vdd
rlabel metal1 5444 4082 5476 4098 0 FILL_1__1617_.gnd
rlabel metal1 5464 4082 5576 4098 0 _1617_.gnd
rlabel metal1 5464 4322 5576 4338 0 _1617_.vdd
rlabel metal2 5473 4173 5487 4187 0 _1617_.A
rlabel metal2 5493 4193 5507 4207 0 _1617_.B
rlabel metal2 5533 4193 5547 4207 0 _1617_.C
rlabel metal2 5513 4173 5527 4187 0 _1617_.Y
rlabel metal1 5564 4082 5816 4098 0 _1658_.gnd
rlabel metal1 5564 4322 5816 4338 0 _1658_.vdd
rlabel metal2 5653 4173 5667 4187 0 _1658_.D
rlabel metal2 5693 4173 5707 4187 0 _1658_.CLK
rlabel metal2 5773 4173 5787 4187 0 _1658_.Q
rlabel nsubstratencontact 44 4332 44 4332 0 FILL_1__998_.vdd
rlabel metal1 24 4562 56 4578 0 FILL_1__998_.gnd
rlabel nsubstratencontact 24 4332 24 4332 0 FILL_0__998_.vdd
rlabel metal1 4 4562 36 4578 0 FILL_0__998_.gnd
rlabel metal1 44 4562 156 4578 0 _998_.gnd
rlabel metal1 44 4322 156 4338 0 _998_.vdd
rlabel metal2 133 4473 147 4487 0 _998_.A
rlabel metal2 113 4453 127 4467 0 _998_.B
rlabel metal2 73 4453 87 4467 0 _998_.C
rlabel metal2 93 4473 107 4487 0 _998_.Y
rlabel nsubstratencontact 184 4332 184 4332 0 FILL_1__970_.vdd
rlabel metal1 164 4562 196 4578 0 FILL_1__970_.gnd
rlabel nsubstratencontact 164 4332 164 4332 0 FILL_0__970_.vdd
rlabel metal1 144 4562 176 4578 0 FILL_0__970_.gnd
rlabel metal1 184 4562 296 4578 0 _970_.gnd
rlabel metal1 184 4322 296 4338 0 _970_.vdd
rlabel metal2 273 4453 287 4467 0 _970_.A
rlabel metal2 253 4433 267 4447 0 _970_.B
rlabel metal2 233 4453 247 4467 0 _970_.C
rlabel metal2 213 4433 227 4447 0 _970_.Y
rlabel nsubstratencontact 316 4332 316 4332 0 FILL_1__990_.vdd
rlabel metal1 304 4562 336 4578 0 FILL_1__990_.gnd
rlabel nsubstratencontact 296 4332 296 4332 0 FILL_0__990_.vdd
rlabel metal1 284 4562 316 4578 0 FILL_0__990_.gnd
rlabel metal1 324 4562 436 4578 0 _990_.gnd
rlabel metal1 324 4322 436 4338 0 _990_.vdd
rlabel metal2 333 4453 347 4467 0 _990_.A
rlabel metal2 353 4493 367 4507 0 _990_.B
rlabel metal2 373 4453 387 4467 0 _990_.C
rlabel metal2 393 4473 407 4487 0 _990_.Y
rlabel nsubstratencontact 484 4332 484 4332 0 FILL_2__992_.vdd
rlabel metal1 464 4562 496 4578 0 FILL_2__992_.gnd
rlabel nsubstratencontact 464 4332 464 4332 0 FILL_1__992_.vdd
rlabel metal1 444 4562 476 4578 0 FILL_1__992_.gnd
rlabel nsubstratencontact 444 4332 444 4332 0 FILL_0__992_.vdd
rlabel metal1 424 4562 456 4578 0 FILL_0__992_.gnd
rlabel metal1 484 4562 596 4578 0 _992_.gnd
rlabel metal1 484 4322 596 4338 0 _992_.vdd
rlabel metal2 573 4473 587 4487 0 _992_.A
rlabel metal2 553 4453 567 4467 0 _992_.B
rlabel metal2 513 4453 527 4467 0 _992_.C
rlabel metal2 533 4473 547 4487 0 _992_.Y
rlabel nsubstratencontact 624 4332 624 4332 0 FILL_1__984_.vdd
rlabel metal1 604 4562 636 4578 0 FILL_1__984_.gnd
rlabel nsubstratencontact 604 4332 604 4332 0 FILL_0__984_.vdd
rlabel metal1 584 4562 616 4578 0 FILL_0__984_.gnd
rlabel metal1 624 4562 736 4578 0 _984_.gnd
rlabel metal1 624 4322 736 4338 0 _984_.vdd
rlabel metal2 713 4473 727 4487 0 _984_.A
rlabel metal2 693 4453 707 4467 0 _984_.B
rlabel metal2 653 4453 667 4467 0 _984_.C
rlabel metal2 673 4473 687 4487 0 _984_.Y
rlabel nsubstratencontact 756 4332 756 4332 0 FILL_1__983_.vdd
rlabel metal1 744 4562 776 4578 0 FILL_1__983_.gnd
rlabel nsubstratencontact 736 4332 736 4332 0 FILL_0__983_.vdd
rlabel metal1 724 4562 756 4578 0 FILL_0__983_.gnd
rlabel nsubstratencontact 856 4332 856 4332 0 FILL_1__1039_.vdd
rlabel metal1 844 4562 876 4578 0 FILL_1__1039_.gnd
rlabel nsubstratencontact 836 4332 836 4332 0 FILL_0__1039_.vdd
rlabel metal1 824 4562 856 4578 0 FILL_0__1039_.gnd
rlabel metal1 864 4562 976 4578 0 _1039_.gnd
rlabel metal1 864 4322 976 4338 0 _1039_.vdd
rlabel metal2 873 4453 887 4467 0 _1039_.A
rlabel metal2 893 4493 907 4507 0 _1039_.B
rlabel metal2 913 4453 927 4467 0 _1039_.C
rlabel metal2 933 4473 947 4487 0 _1039_.Y
rlabel metal1 764 4562 836 4578 0 _983_.gnd
rlabel metal1 764 4322 836 4338 0 _983_.vdd
rlabel metal2 773 4493 787 4507 0 _983_.A
rlabel metal2 793 4453 807 4467 0 _983_.Y
rlabel nsubstratencontact 1004 4332 1004 4332 0 FILL_1__931_.vdd
rlabel metal1 984 4562 1016 4578 0 FILL_1__931_.gnd
rlabel nsubstratencontact 984 4332 984 4332 0 FILL_0__931_.vdd
rlabel metal1 964 4562 996 4578 0 FILL_0__931_.gnd
rlabel metal1 1004 4562 1076 4578 0 _931_.gnd
rlabel metal1 1004 4322 1076 4338 0 _931_.vdd
rlabel metal2 1053 4493 1067 4507 0 _931_.A
rlabel metal2 1033 4453 1047 4467 0 _931_.Y
rlabel nsubstratencontact 1104 4332 1104 4332 0 FILL_1__1143_.vdd
rlabel metal1 1084 4562 1116 4578 0 FILL_1__1143_.gnd
rlabel nsubstratencontact 1084 4332 1084 4332 0 FILL_0__1143_.vdd
rlabel metal1 1064 4562 1096 4578 0 FILL_0__1143_.gnd
rlabel metal1 1104 4562 1216 4578 0 _1143_.gnd
rlabel metal1 1104 4322 1216 4338 0 _1143_.vdd
rlabel metal2 1193 4453 1207 4467 0 _1143_.A
rlabel metal2 1173 4433 1187 4447 0 _1143_.B
rlabel metal2 1153 4453 1167 4467 0 _1143_.C
rlabel metal2 1133 4433 1147 4447 0 _1143_.Y
rlabel nsubstratencontact 1244 4332 1244 4332 0 FILL_1__1130_.vdd
rlabel metal1 1224 4562 1256 4578 0 FILL_1__1130_.gnd
rlabel nsubstratencontact 1224 4332 1224 4332 0 FILL_0__1130_.vdd
rlabel metal1 1204 4562 1236 4578 0 FILL_0__1130_.gnd
rlabel metal1 1244 4562 1356 4578 0 _1130_.gnd
rlabel metal1 1244 4322 1356 4338 0 _1130_.vdd
rlabel metal2 1333 4453 1347 4467 0 _1130_.A
rlabel metal2 1313 4493 1327 4507 0 _1130_.B
rlabel metal2 1293 4453 1307 4467 0 _1130_.C
rlabel metal2 1273 4473 1287 4487 0 _1130_.Y
rlabel nsubstratencontact 1384 4332 1384 4332 0 FILL_1__1129_.vdd
rlabel metal1 1364 4562 1396 4578 0 FILL_1__1129_.gnd
rlabel nsubstratencontact 1364 4332 1364 4332 0 FILL_0__1129_.vdd
rlabel metal1 1344 4562 1376 4578 0 FILL_0__1129_.gnd
rlabel metal1 1384 4562 1456 4578 0 _1129_.gnd
rlabel metal1 1384 4322 1456 4338 0 _1129_.vdd
rlabel metal2 1433 4493 1447 4507 0 _1129_.A
rlabel metal2 1413 4453 1427 4467 0 _1129_.Y
rlabel nsubstratencontact 1476 4332 1476 4332 0 FILL_1__982_.vdd
rlabel metal1 1464 4562 1496 4578 0 FILL_1__982_.gnd
rlabel nsubstratencontact 1456 4332 1456 4332 0 FILL_0__982_.vdd
rlabel metal1 1444 4562 1476 4578 0 FILL_0__982_.gnd
rlabel metal1 1484 4562 1596 4578 0 _982_.gnd
rlabel metal1 1484 4322 1596 4338 0 _982_.vdd
rlabel metal2 1493 4473 1507 4487 0 _982_.A
rlabel metal2 1513 4453 1527 4467 0 _982_.B
rlabel metal2 1553 4453 1567 4467 0 _982_.C
rlabel metal2 1533 4473 1547 4487 0 _982_.Y
rlabel nsubstratencontact 1624 4332 1624 4332 0 FILL_1__977_.vdd
rlabel metal1 1604 4562 1636 4578 0 FILL_1__977_.gnd
rlabel nsubstratencontact 1604 4332 1604 4332 0 FILL_0__977_.vdd
rlabel metal1 1584 4562 1616 4578 0 FILL_0__977_.gnd
rlabel metal1 1624 4562 1716 4578 0 _977_.gnd
rlabel metal1 1624 4322 1716 4338 0 _977_.vdd
rlabel metal2 1693 4433 1707 4447 0 _977_.A
rlabel metal2 1653 4433 1667 4447 0 _977_.B
rlabel metal2 1673 4453 1687 4467 0 _977_.Y
rlabel nsubstratencontact 1744 4332 1744 4332 0 FILL_1__932_.vdd
rlabel metal1 1724 4562 1756 4578 0 FILL_1__932_.gnd
rlabel nsubstratencontact 1724 4332 1724 4332 0 FILL_0__932_.vdd
rlabel metal1 1704 4562 1736 4578 0 FILL_0__932_.gnd
rlabel metal1 1744 4562 1856 4578 0 _932_.gnd
rlabel metal1 1744 4322 1856 4338 0 _932_.vdd
rlabel metal2 1833 4453 1847 4467 0 _932_.A
rlabel metal2 1813 4433 1827 4447 0 _932_.B
rlabel metal2 1793 4453 1807 4467 0 _932_.C
rlabel metal2 1773 4433 1787 4447 0 _932_.Y
rlabel nsubstratencontact 1884 4332 1884 4332 0 FILL_1__981_.vdd
rlabel metal1 1864 4562 1896 4578 0 FILL_1__981_.gnd
rlabel nsubstratencontact 1864 4332 1864 4332 0 FILL_0__981_.vdd
rlabel metal1 1844 4562 1876 4578 0 FILL_0__981_.gnd
rlabel metal1 1884 4562 1976 4578 0 _981_.gnd
rlabel metal1 1884 4322 1976 4338 0 _981_.vdd
rlabel metal2 1913 4473 1927 4487 0 _981_.B
rlabel metal2 1953 4473 1967 4487 0 _981_.A
rlabel metal2 1933 4493 1947 4507 0 _981_.Y
rlabel nsubstratencontact 2004 4332 2004 4332 0 FILL_1__980_.vdd
rlabel metal1 1984 4562 2016 4578 0 FILL_1__980_.gnd
rlabel nsubstratencontact 1984 4332 1984 4332 0 FILL_0__980_.vdd
rlabel metal1 1964 4562 1996 4578 0 FILL_0__980_.gnd
rlabel metal1 2004 4562 2116 4578 0 _980_.gnd
rlabel metal1 2004 4322 2116 4338 0 _980_.vdd
rlabel metal2 2093 4453 2107 4467 0 _980_.A
rlabel metal2 2073 4433 2087 4447 0 _980_.B
rlabel metal2 2053 4453 2067 4467 0 _980_.C
rlabel metal2 2033 4433 2047 4447 0 _980_.Y
rlabel nsubstratencontact 2164 4332 2164 4332 0 FILL_2__979_.vdd
rlabel metal1 2144 4562 2176 4578 0 FILL_2__979_.gnd
rlabel nsubstratencontact 2144 4332 2144 4332 0 FILL_1__979_.vdd
rlabel metal1 2124 4562 2156 4578 0 FILL_1__979_.gnd
rlabel nsubstratencontact 2124 4332 2124 4332 0 FILL_0__979_.vdd
rlabel metal1 2104 4562 2136 4578 0 FILL_0__979_.gnd
rlabel nsubstratencontact 2284 4332 2284 4332 0 FILL_0__1090_.vdd
rlabel metal1 2264 4562 2296 4578 0 FILL_0__1090_.gnd
rlabel metal1 2164 4562 2276 4578 0 _979_.gnd
rlabel metal1 2164 4322 2276 4338 0 _979_.vdd
rlabel metal2 2253 4453 2267 4467 0 _979_.A
rlabel metal2 2233 4433 2247 4447 0 _979_.B
rlabel metal2 2213 4453 2227 4467 0 _979_.C
rlabel metal2 2193 4433 2207 4447 0 _979_.Y
rlabel nsubstratencontact 2304 4332 2304 4332 0 FILL_1__1090_.vdd
rlabel metal1 2284 4562 2316 4578 0 FILL_1__1090_.gnd
rlabel nsubstratencontact 2404 4332 2404 4332 0 FILL_0__1522_.vdd
rlabel metal1 2384 4562 2416 4578 0 FILL_0__1522_.gnd
rlabel metal1 2304 4562 2396 4578 0 _1090_.gnd
rlabel metal1 2304 4322 2396 4338 0 _1090_.vdd
rlabel metal2 2373 4433 2387 4447 0 _1090_.A
rlabel metal2 2333 4433 2347 4447 0 _1090_.B
rlabel metal2 2353 4453 2367 4467 0 _1090_.Y
rlabel nsubstratencontact 2424 4332 2424 4332 0 FILL_1__1522_.vdd
rlabel metal1 2404 4562 2436 4578 0 FILL_1__1522_.gnd
rlabel metal1 2424 4562 2536 4578 0 _1522_.gnd
rlabel metal1 2424 4322 2536 4338 0 _1522_.vdd
rlabel metal2 2513 4453 2527 4467 0 _1522_.A
rlabel metal2 2493 4433 2507 4447 0 _1522_.B
rlabel metal2 2473 4453 2487 4467 0 _1522_.C
rlabel metal2 2453 4433 2467 4447 0 _1522_.Y
rlabel nsubstratencontact 2536 4332 2536 4332 0 FILL_0__1584_.vdd
rlabel metal1 2524 4562 2556 4578 0 FILL_0__1584_.gnd
rlabel nsubstratencontact 2556 4332 2556 4332 0 FILL_1__1584_.vdd
rlabel metal1 2544 4562 2576 4578 0 FILL_1__1584_.gnd
rlabel metal1 2564 4562 2676 4578 0 _1584_.gnd
rlabel metal1 2564 4322 2676 4338 0 _1584_.vdd
rlabel metal2 2573 4453 2587 4467 0 _1584_.A
rlabel metal2 2593 4433 2607 4447 0 _1584_.B
rlabel metal2 2613 4453 2627 4467 0 _1584_.C
rlabel metal2 2633 4433 2647 4447 0 _1584_.Y
rlabel nsubstratencontact 2704 4332 2704 4332 0 FILL_1__1516_.vdd
rlabel metal1 2684 4562 2716 4578 0 FILL_1__1516_.gnd
rlabel nsubstratencontact 2784 4332 2784 4332 0 FILL_0__1583_.vdd
rlabel metal1 2764 4562 2796 4578 0 FILL_0__1583_.gnd
rlabel nsubstratencontact 2684 4332 2684 4332 0 FILL_0__1516_.vdd
rlabel metal1 2664 4562 2696 4578 0 FILL_0__1516_.gnd
rlabel metal1 2704 4562 2776 4578 0 _1516_.gnd
rlabel metal1 2704 4322 2776 4338 0 _1516_.vdd
rlabel metal2 2753 4493 2767 4507 0 _1516_.A
rlabel metal2 2733 4453 2747 4467 0 _1516_.Y
rlabel nsubstratencontact 2804 4332 2804 4332 0 FILL_1__1583_.vdd
rlabel metal1 2784 4562 2816 4578 0 FILL_1__1583_.gnd
rlabel nsubstratencontact 2904 4332 2904 4332 0 FILL_0__1560_.vdd
rlabel metal1 2884 4562 2916 4578 0 FILL_0__1560_.gnd
rlabel metal1 2804 4562 2896 4578 0 _1583_.gnd
rlabel metal1 2804 4322 2896 4338 0 _1583_.vdd
rlabel metal2 2833 4473 2847 4487 0 _1583_.B
rlabel metal2 2873 4473 2887 4487 0 _1583_.A
rlabel metal2 2853 4493 2867 4507 0 _1583_.Y
rlabel nsubstratencontact 2924 4332 2924 4332 0 FILL_1__1560_.vdd
rlabel metal1 2904 4562 2936 4578 0 FILL_1__1560_.gnd
rlabel nsubstratencontact 3044 4332 3044 4332 0 FILL_0__1573_.vdd
rlabel metal1 3024 4562 3056 4578 0 FILL_0__1573_.gnd
rlabel metal1 2924 4562 3036 4578 0 _1560_.gnd
rlabel metal1 2924 4322 3036 4338 0 _1560_.vdd
rlabel metal2 3013 4453 3027 4467 0 _1560_.A
rlabel metal2 2993 4433 3007 4447 0 _1560_.B
rlabel metal2 2973 4453 2987 4467 0 _1560_.C
rlabel metal2 2953 4433 2967 4447 0 _1560_.Y
rlabel nsubstratencontact 3064 4332 3064 4332 0 FILL_1__1573_.vdd
rlabel metal1 3044 4562 3076 4578 0 FILL_1__1573_.gnd
rlabel metal1 3064 4562 3176 4578 0 _1573_.gnd
rlabel metal1 3064 4322 3176 4338 0 _1573_.vdd
rlabel metal2 3153 4453 3167 4467 0 _1573_.A
rlabel metal2 3133 4433 3147 4447 0 _1573_.B
rlabel metal2 3113 4453 3127 4467 0 _1573_.C
rlabel metal2 3093 4433 3107 4447 0 _1573_.Y
rlabel nsubstratencontact 3196 4332 3196 4332 0 FILL_1__1561_.vdd
rlabel metal1 3184 4562 3216 4578 0 FILL_1__1561_.gnd
rlabel nsubstratencontact 3276 4332 3276 4332 0 FILL_0__1575_.vdd
rlabel metal1 3264 4562 3296 4578 0 FILL_0__1575_.gnd
rlabel nsubstratencontact 3176 4332 3176 4332 0 FILL_0__1561_.vdd
rlabel metal1 3164 4562 3196 4578 0 FILL_0__1561_.gnd
rlabel metal1 3204 4562 3276 4578 0 _1561_.gnd
rlabel metal1 3204 4322 3276 4338 0 _1561_.vdd
rlabel metal2 3213 4493 3227 4507 0 _1561_.A
rlabel metal2 3233 4453 3247 4467 0 _1561_.Y
rlabel nsubstratencontact 3296 4332 3296 4332 0 FILL_1__1575_.vdd
rlabel metal1 3284 4562 3316 4578 0 FILL_1__1575_.gnd
rlabel nsubstratencontact 3424 4332 3424 4332 0 FILL_0__1563_.vdd
rlabel metal1 3404 4562 3436 4578 0 FILL_0__1563_.gnd
rlabel metal1 3304 4562 3416 4578 0 _1575_.gnd
rlabel metal1 3304 4322 3416 4338 0 _1575_.vdd
rlabel metal2 3313 4473 3327 4487 0 _1575_.A
rlabel metal2 3333 4453 3347 4467 0 _1575_.B
rlabel metal2 3373 4453 3387 4467 0 _1575_.C
rlabel metal2 3353 4473 3367 4487 0 _1575_.Y
rlabel nsubstratencontact 3444 4332 3444 4332 0 FILL_1__1563_.vdd
rlabel metal1 3424 4562 3456 4578 0 FILL_1__1563_.gnd
rlabel metal1 3444 4562 3556 4578 0 _1563_.gnd
rlabel metal1 3444 4322 3556 4338 0 _1563_.vdd
rlabel metal2 3533 4473 3547 4487 0 _1563_.A
rlabel metal2 3473 4473 3487 4487 0 _1563_.Y
rlabel metal2 3493 4433 3507 4447 0 _1563_.B
rlabel nsubstratencontact 3596 4332 3596 4332 0 FILL_2__1559_.vdd
rlabel metal1 3584 4562 3616 4578 0 FILL_2__1559_.gnd
rlabel nsubstratencontact 3576 4332 3576 4332 0 FILL_1__1559_.vdd
rlabel metal1 3564 4562 3596 4578 0 FILL_1__1559_.gnd
rlabel nsubstratencontact 3556 4332 3556 4332 0 FILL_0__1559_.vdd
rlabel metal1 3544 4562 3576 4578 0 FILL_0__1559_.gnd
rlabel metal1 3604 4562 3696 4578 0 _1559_.gnd
rlabel metal1 3604 4322 3696 4338 0 _1559_.vdd
rlabel metal2 3613 4433 3627 4447 0 _1559_.A
rlabel metal2 3653 4433 3667 4447 0 _1559_.B
rlabel metal2 3633 4453 3647 4467 0 _1559_.Y
rlabel nsubstratencontact 3724 4332 3724 4332 0 FILL_1__1558_.vdd
rlabel metal1 3704 4562 3736 4578 0 FILL_1__1558_.gnd
rlabel nsubstratencontact 3704 4332 3704 4332 0 FILL_0__1558_.vdd
rlabel metal1 3684 4562 3716 4578 0 FILL_0__1558_.gnd
rlabel metal1 3724 4562 3836 4578 0 _1558_.gnd
rlabel metal1 3724 4322 3836 4338 0 _1558_.vdd
rlabel metal2 3813 4493 3827 4507 0 _1558_.A
rlabel metal2 3793 4473 3807 4487 0 _1558_.B
rlabel metal2 3753 4453 3767 4467 0 _1558_.Y
rlabel nsubstratencontact 3856 4332 3856 4332 0 FILL_1__1557_.vdd
rlabel metal1 3844 4562 3876 4578 0 FILL_1__1557_.gnd
rlabel nsubstratencontact 3836 4332 3836 4332 0 FILL_0__1557_.vdd
rlabel metal1 3824 4562 3856 4578 0 FILL_0__1557_.gnd
rlabel metal1 3864 4562 3956 4578 0 _1557_.gnd
rlabel metal1 3864 4322 3956 4338 0 _1557_.vdd
rlabel metal2 3873 4433 3887 4447 0 _1557_.A
rlabel metal2 3913 4433 3927 4447 0 _1557_.B
rlabel metal2 3893 4453 3907 4467 0 _1557_.Y
rlabel nsubstratencontact 3984 4332 3984 4332 0 FILL_1_BUFX2_insert7.vdd
rlabel metal1 3964 4562 3996 4578 0 FILL_1_BUFX2_insert7.gnd
rlabel nsubstratencontact 3964 4332 3964 4332 0 FILL_0_BUFX2_insert7.vdd
rlabel metal1 3944 4562 3976 4578 0 FILL_0_BUFX2_insert7.gnd
rlabel metal1 3984 4562 4076 4578 0 BUFX2_insert7.gnd
rlabel metal1 3984 4322 4076 4338 0 BUFX2_insert7.vdd
rlabel metal2 4053 4473 4067 4487 0 BUFX2_insert7.A
rlabel metal2 4013 4473 4027 4487 0 BUFX2_insert7.Y
rlabel nsubstratencontact 4096 4332 4096 4332 0 FILL_1__921_.vdd
rlabel metal1 4084 4562 4116 4578 0 FILL_1__921_.gnd
rlabel nsubstratencontact 4076 4332 4076 4332 0 FILL_0__921_.vdd
rlabel metal1 4064 4562 4096 4578 0 FILL_0__921_.gnd
rlabel metal1 4104 4562 4216 4578 0 _921_.gnd
rlabel metal1 4104 4322 4216 4338 0 _921_.vdd
rlabel metal2 4113 4473 4127 4487 0 _921_.A
rlabel metal2 4173 4473 4187 4487 0 _921_.Y
rlabel metal2 4153 4433 4167 4447 0 _921_.B
rlabel nsubstratencontact 4244 4332 4244 4332 0 FILL_1__1449_.vdd
rlabel metal1 4224 4562 4256 4578 0 FILL_1__1449_.gnd
rlabel nsubstratencontact 4224 4332 4224 4332 0 FILL_0__1449_.vdd
rlabel metal1 4204 4562 4236 4578 0 FILL_0__1449_.gnd
rlabel metal1 4244 4562 4336 4578 0 _1449_.gnd
rlabel metal1 4244 4322 4336 4338 0 _1449_.vdd
rlabel metal2 4313 4433 4327 4447 0 _1449_.A
rlabel metal2 4273 4433 4287 4447 0 _1449_.B
rlabel metal2 4293 4453 4307 4467 0 _1449_.Y
rlabel nsubstratencontact 4364 4332 4364 4332 0 FILL_1__1452_.vdd
rlabel metal1 4344 4562 4376 4578 0 FILL_1__1452_.gnd
rlabel nsubstratencontact 4344 4332 4344 4332 0 FILL_0__1452_.vdd
rlabel metal1 4324 4562 4356 4578 0 FILL_0__1452_.gnd
rlabel metal1 4364 4562 4476 4578 0 _1452_.gnd
rlabel metal1 4364 4322 4476 4338 0 _1452_.vdd
rlabel metal2 4453 4473 4467 4487 0 _1452_.A
rlabel metal2 4433 4453 4447 4467 0 _1452_.B
rlabel metal2 4393 4453 4407 4467 0 _1452_.C
rlabel metal2 4413 4473 4427 4487 0 _1452_.Y
rlabel nsubstratencontact 4496 4332 4496 4332 0 FILL_1__1453_.vdd
rlabel metal1 4484 4562 4516 4578 0 FILL_1__1453_.gnd
rlabel nsubstratencontact 4476 4332 4476 4332 0 FILL_0__1453_.vdd
rlabel metal1 4464 4562 4496 4578 0 FILL_0__1453_.gnd
rlabel metal1 4504 4562 4596 4578 0 _1453_.gnd
rlabel metal1 4504 4322 4596 4338 0 _1453_.vdd
rlabel metal2 4513 4433 4527 4447 0 _1453_.A
rlabel metal2 4553 4433 4567 4447 0 _1453_.B
rlabel metal2 4533 4453 4547 4467 0 _1453_.Y
rlabel nsubstratencontact 4624 4332 4624 4332 0 FILL_1__1505_.vdd
rlabel metal1 4604 4562 4636 4578 0 FILL_1__1505_.gnd
rlabel nsubstratencontact 4604 4332 4604 4332 0 FILL_0__1505_.vdd
rlabel metal1 4584 4562 4616 4578 0 FILL_0__1505_.gnd
rlabel metal1 4624 4562 4716 4578 0 _1505_.gnd
rlabel metal1 4624 4322 4716 4338 0 _1505_.vdd
rlabel metal2 4693 4433 4707 4447 0 _1505_.A
rlabel metal2 4653 4433 4667 4447 0 _1505_.B
rlabel metal2 4673 4453 4687 4467 0 _1505_.Y
rlabel nsubstratencontact 4736 4332 4736 4332 0 FILL_1__1501_.vdd
rlabel metal1 4724 4562 4756 4578 0 FILL_1__1501_.gnd
rlabel nsubstratencontact 4716 4332 4716 4332 0 FILL_0__1501_.vdd
rlabel metal1 4704 4562 4736 4578 0 FILL_0__1501_.gnd
rlabel metal1 4744 4562 4816 4578 0 _1501_.gnd
rlabel metal1 4744 4322 4816 4338 0 _1501_.vdd
rlabel metal2 4753 4493 4767 4507 0 _1501_.A
rlabel metal2 4773 4453 4787 4467 0 _1501_.Y
rlabel nsubstratencontact 4836 4332 4836 4332 0 FILL_1__1502_.vdd
rlabel metal1 4824 4562 4856 4578 0 FILL_1__1502_.gnd
rlabel nsubstratencontact 4816 4332 4816 4332 0 FILL_0__1502_.vdd
rlabel metal1 4804 4562 4836 4578 0 FILL_0__1502_.gnd
rlabel metal1 4844 4562 4936 4578 0 _1502_.gnd
rlabel metal1 4844 4322 4936 4338 0 _1502_.vdd
rlabel metal2 4853 4433 4867 4447 0 _1502_.A
rlabel metal2 4893 4433 4907 4447 0 _1502_.B
rlabel metal2 4873 4453 4887 4467 0 _1502_.Y
rlabel nsubstratencontact 4956 4332 4956 4332 0 FILL_1__1551_.vdd
rlabel metal1 4944 4562 4976 4578 0 FILL_1__1551_.gnd
rlabel nsubstratencontact 4936 4332 4936 4332 0 FILL_0__1551_.vdd
rlabel metal1 4924 4562 4956 4578 0 FILL_0__1551_.gnd
rlabel metal1 4964 4562 5076 4578 0 _1551_.gnd
rlabel metal1 4964 4322 5076 4338 0 _1551_.vdd
rlabel metal2 4973 4473 4987 4487 0 _1551_.A
rlabel metal2 4993 4453 5007 4467 0 _1551_.B
rlabel metal2 5033 4453 5047 4467 0 _1551_.C
rlabel metal2 5013 4473 5027 4487 0 _1551_.Y
rlabel metal1 5484 4562 5596 4578 0 _1550_.gnd
rlabel metal1 5484 4322 5596 4338 0 _1550_.vdd
rlabel metal2 5493 4493 5507 4507 0 _1550_.A
rlabel metal2 5513 4473 5527 4487 0 _1550_.B
rlabel metal2 5553 4453 5567 4467 0 _1550_.Y
rlabel metal1 5344 4562 5456 4578 0 _1652_.gnd
rlabel metal1 5344 4322 5456 4338 0 _1652_.vdd
rlabel metal2 5353 4473 5367 4487 0 _1652_.A
rlabel metal2 5373 4453 5387 4467 0 _1652_.B
rlabel metal2 5413 4453 5427 4467 0 _1652_.C
rlabel metal2 5393 4473 5407 4487 0 _1652_.Y
rlabel metal1 5064 4562 5316 4578 0 _1684_.gnd
rlabel metal1 5064 4322 5316 4338 0 _1684_.vdd
rlabel metal2 5213 4473 5227 4487 0 _1684_.D
rlabel metal2 5173 4473 5187 4487 0 _1684_.CLK
rlabel metal2 5093 4473 5107 4487 0 _1684_.Q
rlabel nsubstratencontact 5456 4332 5456 4332 0 FILL_0__1550_.vdd
rlabel metal1 5444 4562 5476 4578 0 FILL_0__1550_.gnd
rlabel nsubstratencontact 5316 4332 5316 4332 0 FILL_0__1652_.vdd
rlabel metal1 5304 4562 5336 4578 0 FILL_0__1652_.gnd
rlabel nsubstratencontact 5476 4332 5476 4332 0 FILL_1__1550_.vdd
rlabel metal1 5464 4562 5496 4578 0 FILL_1__1550_.gnd
rlabel nsubstratencontact 5336 4332 5336 4332 0 FILL_1__1652_.vdd
rlabel metal1 5324 4562 5356 4578 0 FILL_1__1652_.gnd
rlabel metal1 5624 4562 5736 4578 0 _1614_.gnd
rlabel metal1 5624 4322 5736 4338 0 _1614_.vdd
rlabel metal2 5713 4473 5727 4487 0 _1614_.A
rlabel metal2 5693 4453 5707 4467 0 _1614_.B
rlabel metal2 5653 4453 5667 4467 0 _1614_.C
rlabel metal2 5673 4473 5687 4487 0 _1614_.Y
rlabel nsubstratencontact 5744 4332 5744 4332 0 FILL85950x64950.vdd
rlabel metal1 5724 4562 5756 4578 0 FILL85950x64950.gnd
rlabel nsubstratencontact 5764 4332 5764 4332 0 FILL86250x64950.vdd
rlabel metal1 5744 4562 5776 4578 0 FILL86250x64950.gnd
rlabel nsubstratencontact 5784 4332 5784 4332 0 FILL86550x64950.vdd
rlabel metal1 5764 4562 5796 4578 0 FILL86550x64950.gnd
rlabel nsubstratencontact 5804 4332 5804 4332 0 FILL86850x64950.vdd
rlabel metal1 5784 4562 5816 4578 0 FILL86850x64950.gnd
rlabel nsubstratencontact 5604 4332 5604 4332 0 FILL_0__1614_.vdd
rlabel metal1 5584 4562 5616 4578 0 FILL_0__1614_.gnd
rlabel nsubstratencontact 5624 4332 5624 4332 0 FILL_1__1614_.vdd
rlabel metal1 5604 4562 5636 4578 0 FILL_1__1614_.gnd
rlabel nsubstratencontact 44 4808 44 4808 0 FILL_1__1034_.vdd
rlabel metal1 24 4562 56 4578 0 FILL_1__1034_.gnd
rlabel nsubstratencontact 24 4808 24 4808 0 FILL_0__1034_.vdd
rlabel metal1 4 4562 36 4578 0 FILL_0__1034_.gnd
rlabel metal1 44 4562 156 4578 0 _1034_.gnd
rlabel metal1 44 4802 156 4818 0 _1034_.vdd
rlabel metal2 133 4673 147 4687 0 _1034_.A
rlabel metal2 113 4633 127 4647 0 _1034_.B
rlabel metal2 93 4673 107 4687 0 _1034_.C
rlabel metal2 73 4653 87 4667 0 _1034_.Y
rlabel nsubstratencontact 184 4808 184 4808 0 FILL_1__974_.vdd
rlabel metal1 164 4562 196 4578 0 FILL_1__974_.gnd
rlabel nsubstratencontact 164 4808 164 4808 0 FILL_0__974_.vdd
rlabel metal1 144 4562 176 4578 0 FILL_0__974_.gnd
rlabel metal1 184 4562 296 4578 0 _974_.gnd
rlabel metal1 184 4802 296 4818 0 _974_.vdd
rlabel metal2 273 4673 287 4687 0 _974_.A
rlabel metal2 253 4693 267 4707 0 _974_.B
rlabel metal2 233 4673 247 4687 0 _974_.C
rlabel metal2 213 4693 227 4707 0 _974_.Y
rlabel nsubstratencontact 316 4808 316 4808 0 FILL_1__989_.vdd
rlabel metal1 304 4562 336 4578 0 FILL_1__989_.gnd
rlabel nsubstratencontact 296 4808 296 4808 0 FILL_0__989_.vdd
rlabel metal1 284 4562 316 4578 0 FILL_0__989_.gnd
rlabel metal1 324 4562 436 4578 0 _989_.gnd
rlabel metal1 324 4802 436 4818 0 _989_.vdd
rlabel metal2 333 4673 347 4687 0 _989_.A
rlabel metal2 353 4633 367 4647 0 _989_.B
rlabel metal2 373 4673 387 4687 0 _989_.C
rlabel metal2 393 4653 407 4667 0 _989_.Y
rlabel nsubstratencontact 456 4808 456 4808 0 FILL_1__993_.vdd
rlabel metal1 444 4562 476 4578 0 FILL_1__993_.gnd
rlabel nsubstratencontact 436 4808 436 4808 0 FILL_0__993_.vdd
rlabel metal1 424 4562 456 4578 0 FILL_0__993_.gnd
rlabel metal1 464 4562 556 4578 0 _993_.gnd
rlabel metal1 464 4802 556 4818 0 _993_.vdd
rlabel metal2 473 4693 487 4707 0 _993_.A
rlabel metal2 513 4693 527 4707 0 _993_.B
rlabel metal2 493 4673 507 4687 0 _993_.Y
rlabel nsubstratencontact 584 4808 584 4808 0 FILL_1__991_.vdd
rlabel metal1 564 4562 596 4578 0 FILL_1__991_.gnd
rlabel nsubstratencontact 564 4808 564 4808 0 FILL_0__991_.vdd
rlabel metal1 544 4562 576 4578 0 FILL_0__991_.gnd
rlabel metal1 584 4562 696 4578 0 _991_.gnd
rlabel metal1 584 4802 696 4818 0 _991_.vdd
rlabel metal2 673 4673 687 4687 0 _991_.A
rlabel metal2 653 4693 667 4707 0 _991_.B
rlabel metal2 633 4673 647 4687 0 _991_.C
rlabel metal2 613 4693 627 4707 0 _991_.Y
rlabel nsubstratencontact 744 4808 744 4808 0 FILL_2__986_.vdd
rlabel metal1 724 4562 756 4578 0 FILL_2__986_.gnd
rlabel nsubstratencontact 724 4808 724 4808 0 FILL_1__986_.vdd
rlabel metal1 704 4562 736 4578 0 FILL_1__986_.gnd
rlabel nsubstratencontact 704 4808 704 4808 0 FILL_0__986_.vdd
rlabel metal1 684 4562 716 4578 0 FILL_0__986_.gnd
rlabel metal1 744 4562 856 4578 0 _986_.gnd
rlabel metal1 744 4802 856 4818 0 _986_.vdd
rlabel metal2 833 4673 847 4687 0 _986_.A
rlabel metal2 813 4693 827 4707 0 _986_.B
rlabel metal2 793 4673 807 4687 0 _986_.C
rlabel metal2 773 4693 787 4707 0 _986_.Y
rlabel nsubstratencontact 876 4808 876 4808 0 FILL_1__978_.vdd
rlabel metal1 864 4562 896 4578 0 FILL_1__978_.gnd
rlabel nsubstratencontact 856 4808 856 4808 0 FILL_0__978_.vdd
rlabel metal1 844 4562 876 4578 0 FILL_0__978_.gnd
rlabel nsubstratencontact 976 4808 976 4808 0 FILL_1__985_.vdd
rlabel metal1 964 4562 996 4578 0 FILL_1__985_.gnd
rlabel nsubstratencontact 956 4808 956 4808 0 FILL_0__985_.vdd
rlabel metal1 944 4562 976 4578 0 FILL_0__985_.gnd
rlabel metal1 984 4562 1056 4578 0 _985_.gnd
rlabel metal1 984 4802 1056 4818 0 _985_.vdd
rlabel metal2 993 4633 1007 4647 0 _985_.A
rlabel metal2 1013 4673 1027 4687 0 _985_.Y
rlabel metal1 884 4562 956 4578 0 _978_.gnd
rlabel metal1 884 4802 956 4818 0 _978_.vdd
rlabel metal2 893 4633 907 4647 0 _978_.A
rlabel metal2 913 4673 927 4687 0 _978_.Y
rlabel nsubstratencontact 1084 4808 1084 4808 0 FILL_1__943_.vdd
rlabel metal1 1064 4562 1096 4578 0 FILL_1__943_.gnd
rlabel nsubstratencontact 1064 4808 1064 4808 0 FILL_0__943_.vdd
rlabel metal1 1044 4562 1076 4578 0 FILL_0__943_.gnd
rlabel metal1 1084 4562 1156 4578 0 _943_.gnd
rlabel metal1 1084 4802 1156 4818 0 _943_.vdd
rlabel metal2 1133 4633 1147 4647 0 _943_.A
rlabel metal2 1113 4673 1127 4687 0 _943_.Y
rlabel nsubstratencontact 1184 4808 1184 4808 0 FILL_1__937_.vdd
rlabel metal1 1164 4562 1196 4578 0 FILL_1__937_.gnd
rlabel nsubstratencontact 1164 4808 1164 4808 0 FILL_0__937_.vdd
rlabel metal1 1144 4562 1176 4578 0 FILL_0__937_.gnd
rlabel metal1 1184 4562 1296 4578 0 _937_.gnd
rlabel metal1 1184 4802 1296 4818 0 _937_.vdd
rlabel metal2 1273 4653 1287 4667 0 _937_.A
rlabel metal2 1253 4673 1267 4687 0 _937_.B
rlabel metal2 1213 4673 1227 4687 0 _937_.C
rlabel metal2 1233 4653 1247 4667 0 _937_.Y
rlabel nsubstratencontact 1316 4808 1316 4808 0 FILL_1__1153_.vdd
rlabel metal1 1304 4562 1336 4578 0 FILL_1__1153_.gnd
rlabel nsubstratencontact 1296 4808 1296 4808 0 FILL_0__1153_.vdd
rlabel metal1 1284 4562 1316 4578 0 FILL_0__1153_.gnd
rlabel metal1 1324 4562 1436 4578 0 _1153_.gnd
rlabel metal1 1324 4802 1436 4818 0 _1153_.vdd
rlabel metal2 1333 4653 1347 4667 0 _1153_.A
rlabel metal2 1353 4673 1367 4687 0 _1153_.B
rlabel metal2 1393 4673 1407 4687 0 _1153_.C
rlabel metal2 1373 4653 1387 4667 0 _1153_.Y
rlabel nsubstratencontact 1456 4808 1456 4808 0 FILL_1__936_.vdd
rlabel metal1 1444 4562 1476 4578 0 FILL_1__936_.gnd
rlabel nsubstratencontact 1436 4808 1436 4808 0 FILL_0__936_.vdd
rlabel metal1 1424 4562 1456 4578 0 FILL_0__936_.gnd
rlabel metal1 1464 4562 1536 4578 0 _936_.gnd
rlabel metal1 1464 4802 1536 4818 0 _936_.vdd
rlabel metal2 1473 4633 1487 4647 0 _936_.A
rlabel metal2 1493 4673 1507 4687 0 _936_.Y
rlabel nsubstratencontact 1556 4808 1556 4808 0 FILL_1__1421_.vdd
rlabel metal1 1544 4562 1576 4578 0 FILL_1__1421_.gnd
rlabel nsubstratencontact 1536 4808 1536 4808 0 FILL_0__1421_.vdd
rlabel metal1 1524 4562 1556 4578 0 FILL_0__1421_.gnd
rlabel metal1 1564 4562 1676 4578 0 _1421_.gnd
rlabel metal1 1564 4802 1676 4818 0 _1421_.vdd
rlabel metal2 1573 4673 1587 4687 0 _1421_.A
rlabel metal2 1593 4693 1607 4707 0 _1421_.B
rlabel metal2 1613 4673 1627 4687 0 _1421_.C
rlabel metal2 1633 4693 1647 4707 0 _1421_.Y
rlabel nsubstratencontact 1704 4808 1704 4808 0 FILL_1__1519_.vdd
rlabel metal1 1684 4562 1716 4578 0 FILL_1__1519_.gnd
rlabel nsubstratencontact 1684 4808 1684 4808 0 FILL_0__1519_.vdd
rlabel metal1 1664 4562 1696 4578 0 FILL_0__1519_.gnd
rlabel metal1 1704 4562 1816 4578 0 _1519_.gnd
rlabel metal1 1704 4802 1816 4818 0 _1519_.vdd
rlabel metal2 1793 4653 1807 4667 0 _1519_.A
rlabel metal2 1773 4673 1787 4687 0 _1519_.B
rlabel metal2 1733 4673 1747 4687 0 _1519_.C
rlabel metal2 1753 4653 1767 4667 0 _1519_.Y
rlabel nsubstratencontact 1844 4808 1844 4808 0 FILL_1__1471_.vdd
rlabel metal1 1824 4562 1856 4578 0 FILL_1__1471_.gnd
rlabel nsubstratencontact 1824 4808 1824 4808 0 FILL_0__1471_.vdd
rlabel metal1 1804 4562 1836 4578 0 FILL_0__1471_.gnd
rlabel metal1 1844 4562 1936 4578 0 _1471_.gnd
rlabel metal1 1844 4802 1936 4818 0 _1471_.vdd
rlabel metal2 1913 4693 1927 4707 0 _1471_.A
rlabel metal2 1873 4693 1887 4707 0 _1471_.B
rlabel metal2 1893 4673 1907 4687 0 _1471_.Y
rlabel nsubstratencontact 1956 4808 1956 4808 0 FILL_1__1518_.vdd
rlabel metal1 1944 4562 1976 4578 0 FILL_1__1518_.gnd
rlabel nsubstratencontact 1936 4808 1936 4808 0 FILL_0__1518_.vdd
rlabel metal1 1924 4562 1956 4578 0 FILL_0__1518_.gnd
rlabel metal1 1964 4562 2076 4578 0 _1518_.gnd
rlabel metal1 1964 4802 2076 4818 0 _1518_.vdd
rlabel metal2 1973 4653 1987 4667 0 _1518_.A
rlabel metal2 1993 4673 2007 4687 0 _1518_.B
rlabel metal2 2033 4673 2047 4687 0 _1518_.C
rlabel metal2 2013 4653 2027 4667 0 _1518_.Y
rlabel nsubstratencontact 2104 4808 2104 4808 0 FILL_1__938_.vdd
rlabel metal1 2084 4562 2116 4578 0 FILL_1__938_.gnd
rlabel nsubstratencontact 2084 4808 2084 4808 0 FILL_0__938_.vdd
rlabel metal1 2064 4562 2096 4578 0 FILL_0__938_.gnd
rlabel metal1 2104 4562 2216 4578 0 _938_.gnd
rlabel metal1 2104 4802 2216 4818 0 _938_.vdd
rlabel metal2 2193 4673 2207 4687 0 _938_.A
rlabel metal2 2173 4693 2187 4707 0 _938_.B
rlabel metal2 2153 4673 2167 4687 0 _938_.C
rlabel metal2 2133 4693 2147 4707 0 _938_.Y
rlabel nsubstratencontact 2244 4808 2244 4808 0 FILL_1_BUFX2_insert6.vdd
rlabel metal1 2224 4562 2256 4578 0 FILL_1_BUFX2_insert6.gnd
rlabel nsubstratencontact 2224 4808 2224 4808 0 FILL_0_BUFX2_insert6.vdd
rlabel metal1 2204 4562 2236 4578 0 FILL_0_BUFX2_insert6.gnd
rlabel metal1 2244 4562 2336 4578 0 BUFX2_insert6.gnd
rlabel metal1 2244 4802 2336 4818 0 BUFX2_insert6.vdd
rlabel metal2 2313 4653 2327 4667 0 BUFX2_insert6.A
rlabel metal2 2273 4653 2287 4667 0 BUFX2_insert6.Y
rlabel nsubstratencontact 2356 4808 2356 4808 0 FILL_1__926_.vdd
rlabel metal1 2344 4562 2376 4578 0 FILL_1__926_.gnd
rlabel nsubstratencontact 2336 4808 2336 4808 0 FILL_0__926_.vdd
rlabel metal1 2324 4562 2356 4578 0 FILL_0__926_.gnd
rlabel metal1 2364 4562 2456 4578 0 _926_.gnd
rlabel metal1 2364 4802 2456 4818 0 _926_.vdd
rlabel metal2 2373 4693 2387 4707 0 _926_.A
rlabel metal2 2413 4693 2427 4707 0 _926_.B
rlabel metal2 2393 4673 2407 4687 0 _926_.Y
rlabel nsubstratencontact 2476 4808 2476 4808 0 FILL_1__952_.vdd
rlabel metal1 2464 4562 2496 4578 0 FILL_1__952_.gnd
rlabel nsubstratencontact 2456 4808 2456 4808 0 FILL_0__952_.vdd
rlabel metal1 2444 4562 2476 4578 0 FILL_0__952_.gnd
rlabel metal1 2484 4562 2576 4578 0 _952_.gnd
rlabel metal1 2484 4802 2576 4818 0 _952_.vdd
rlabel metal2 2493 4693 2507 4707 0 _952_.A
rlabel metal2 2533 4693 2547 4707 0 _952_.B
rlabel metal2 2513 4673 2527 4687 0 _952_.Y
rlabel nsubstratencontact 2604 4808 2604 4808 0 FILL_1_BUFX2_insert10.vdd
rlabel metal1 2584 4562 2616 4578 0 FILL_1_BUFX2_insert10.gnd
rlabel nsubstratencontact 2584 4808 2584 4808 0 FILL_0_BUFX2_insert10.vdd
rlabel metal1 2564 4562 2596 4578 0 FILL_0_BUFX2_insert10.gnd
rlabel metal1 2604 4562 2696 4578 0 BUFX2_insert10.gnd
rlabel metal1 2604 4802 2696 4818 0 BUFX2_insert10.vdd
rlabel metal2 2673 4653 2687 4667 0 BUFX2_insert10.A
rlabel metal2 2633 4653 2647 4667 0 BUFX2_insert10.Y
rlabel nsubstratencontact 2716 4808 2716 4808 0 FILL_1__1317_.vdd
rlabel metal1 2704 4562 2736 4578 0 FILL_1__1317_.gnd
rlabel nsubstratencontact 2696 4808 2696 4808 0 FILL_0__1317_.vdd
rlabel metal1 2684 4562 2716 4578 0 FILL_0__1317_.gnd
rlabel metal1 2724 4562 2836 4578 0 _1317_.gnd
rlabel metal1 2724 4802 2836 4818 0 _1317_.vdd
rlabel metal2 2733 4673 2747 4687 0 _1317_.A
rlabel metal2 2753 4693 2767 4707 0 _1317_.B
rlabel metal2 2773 4673 2787 4687 0 _1317_.C
rlabel metal2 2793 4693 2807 4707 0 _1317_.Y
rlabel nsubstratencontact 2864 4808 2864 4808 0 FILL_1__1321_.vdd
rlabel metal1 2844 4562 2876 4578 0 FILL_1__1321_.gnd
rlabel nsubstratencontact 2844 4808 2844 4808 0 FILL_0__1321_.vdd
rlabel metal1 2824 4562 2856 4578 0 FILL_0__1321_.gnd
rlabel nsubstratencontact 2956 4808 2956 4808 0 FILL_0__1318_.vdd
rlabel metal1 2944 4562 2976 4578 0 FILL_0__1318_.gnd
rlabel metal1 2864 4562 2956 4578 0 _1321_.gnd
rlabel metal1 2864 4802 2956 4818 0 _1321_.vdd
rlabel metal2 2893 4653 2907 4667 0 _1321_.B
rlabel metal2 2933 4653 2947 4667 0 _1321_.A
rlabel metal2 2913 4633 2927 4647 0 _1321_.Y
rlabel nsubstratencontact 2996 4808 2996 4808 0 FILL_2__1318_.vdd
rlabel metal1 2984 4562 3016 4578 0 FILL_2__1318_.gnd
rlabel nsubstratencontact 2976 4808 2976 4808 0 FILL_1__1318_.vdd
rlabel metal1 2964 4562 2996 4578 0 FILL_1__1318_.gnd
rlabel metal1 3004 4562 3136 4578 0 _1318_.gnd
rlabel metal1 3004 4802 3136 4818 0 _1318_.vdd
rlabel metal2 3013 4653 3027 4667 0 _1318_.A
rlabel metal2 3033 4673 3047 4687 0 _1318_.B
rlabel metal2 3093 4653 3107 4667 0 _1318_.C
rlabel metal2 3053 4653 3067 4667 0 _1318_.Y
rlabel metal2 3073 4673 3087 4687 0 _1318_.D
rlabel nsubstratencontact 3164 4808 3164 4808 0 FILL_1__1515_.vdd
rlabel metal1 3144 4562 3176 4578 0 FILL_1__1515_.gnd
rlabel nsubstratencontact 3144 4808 3144 4808 0 FILL_0__1515_.vdd
rlabel metal1 3124 4562 3156 4578 0 FILL_0__1515_.gnd
rlabel nsubstratencontact 3284 4808 3284 4808 0 FILL_1__1322_.vdd
rlabel metal1 3264 4562 3296 4578 0 FILL_1__1322_.gnd
rlabel nsubstratencontact 3264 4808 3264 4808 0 FILL_0__1322_.vdd
rlabel metal1 3244 4562 3276 4578 0 FILL_0__1322_.gnd
rlabel metal1 3164 4562 3256 4578 0 _1515_.gnd
rlabel metal1 3164 4802 3256 4818 0 _1515_.vdd
rlabel metal2 3233 4693 3247 4707 0 _1515_.A
rlabel metal2 3193 4693 3207 4707 0 _1515_.B
rlabel metal2 3213 4673 3227 4687 0 _1515_.Y
rlabel nsubstratencontact 3424 4808 3424 4808 0 FILL_1__1312_.vdd
rlabel metal1 3404 4562 3436 4578 0 FILL_1__1312_.gnd
rlabel nsubstratencontact 3404 4808 3404 4808 0 FILL_0__1312_.vdd
rlabel metal1 3384 4562 3416 4578 0 FILL_0__1312_.gnd
rlabel metal1 3284 4562 3396 4578 0 _1322_.gnd
rlabel metal1 3284 4802 3396 4818 0 _1322_.vdd
rlabel metal2 3373 4673 3387 4687 0 _1322_.A
rlabel metal2 3353 4693 3367 4707 0 _1322_.B
rlabel metal2 3333 4673 3347 4687 0 _1322_.C
rlabel metal2 3313 4693 3327 4707 0 _1322_.Y
rlabel nsubstratencontact 3544 4808 3544 4808 0 FILL_0__1320_.vdd
rlabel metal1 3524 4562 3556 4578 0 FILL_0__1320_.gnd
rlabel metal1 3424 4562 3536 4578 0 _1312_.gnd
rlabel metal1 3424 4802 3536 4818 0 _1312_.vdd
rlabel metal2 3513 4673 3527 4687 0 _1312_.A
rlabel metal2 3493 4633 3507 4647 0 _1312_.B
rlabel metal2 3473 4673 3487 4687 0 _1312_.C
rlabel metal2 3453 4653 3467 4667 0 _1312_.Y
rlabel nsubstratencontact 3564 4808 3564 4808 0 FILL_1__1320_.vdd
rlabel metal1 3544 4562 3576 4578 0 FILL_1__1320_.gnd
rlabel metal1 3564 4562 3676 4578 0 _1320_.gnd
rlabel metal1 3564 4802 3676 4818 0 _1320_.vdd
rlabel metal2 3653 4673 3667 4687 0 _1320_.A
rlabel metal2 3633 4693 3647 4707 0 _1320_.B
rlabel metal2 3613 4673 3627 4687 0 _1320_.C
rlabel metal2 3593 4693 3607 4707 0 _1320_.Y
rlabel nsubstratencontact 3704 4808 3704 4808 0 FILL_1__1316_.vdd
rlabel metal1 3684 4562 3716 4578 0 FILL_1__1316_.gnd
rlabel nsubstratencontact 3684 4808 3684 4808 0 FILL_0__1316_.vdd
rlabel metal1 3664 4562 3696 4578 0 FILL_0__1316_.gnd
rlabel metal1 3704 4562 3816 4578 0 _1316_.gnd
rlabel metal1 3704 4802 3816 4818 0 _1316_.vdd
rlabel metal2 3793 4673 3807 4687 0 _1316_.A
rlabel metal2 3773 4633 3787 4647 0 _1316_.B
rlabel metal2 3753 4673 3767 4687 0 _1316_.C
rlabel metal2 3733 4653 3747 4667 0 _1316_.Y
rlabel nsubstratencontact 3836 4808 3836 4808 0 FILL_1__1319_.vdd
rlabel metal1 3824 4562 3856 4578 0 FILL_1__1319_.gnd
rlabel nsubstratencontact 3816 4808 3816 4808 0 FILL_0__1319_.vdd
rlabel metal1 3804 4562 3836 4578 0 FILL_0__1319_.gnd
rlabel metal1 3844 4562 3956 4578 0 _1319_.gnd
rlabel metal1 3844 4802 3956 4818 0 _1319_.vdd
rlabel metal2 3853 4673 3867 4687 0 _1319_.A
rlabel metal2 3873 4693 3887 4707 0 _1319_.B
rlabel metal2 3893 4673 3907 4687 0 _1319_.C
rlabel metal2 3913 4693 3927 4707 0 _1319_.Y
rlabel nsubstratencontact 3976 4808 3976 4808 0 FILL_1__1315_.vdd
rlabel metal1 3964 4562 3996 4578 0 FILL_1__1315_.gnd
rlabel nsubstratencontact 3956 4808 3956 4808 0 FILL_0__1315_.vdd
rlabel metal1 3944 4562 3976 4578 0 FILL_0__1315_.gnd
rlabel metal1 3984 4562 4096 4578 0 _1315_.gnd
rlabel metal1 3984 4802 4096 4818 0 _1315_.vdd
rlabel metal2 3993 4673 4007 4687 0 _1315_.A
rlabel metal2 4013 4693 4027 4707 0 _1315_.B
rlabel metal2 4033 4673 4047 4687 0 _1315_.C
rlabel metal2 4053 4693 4067 4707 0 _1315_.Y
rlabel nsubstratencontact 4116 4808 4116 4808 0 FILL_1__1306_.vdd
rlabel metal1 4104 4562 4136 4578 0 FILL_1__1306_.gnd
rlabel nsubstratencontact 4096 4808 4096 4808 0 FILL_0__1306_.vdd
rlabel metal1 4084 4562 4116 4578 0 FILL_0__1306_.gnd
rlabel metal1 4124 4562 4196 4578 0 _1306_.gnd
rlabel metal1 4124 4802 4196 4818 0 _1306_.vdd
rlabel metal2 4133 4633 4147 4647 0 _1306_.A
rlabel metal2 4153 4673 4167 4687 0 _1306_.Y
rlabel nsubstratencontact 4224 4808 4224 4808 0 FILL_1__1314_.vdd
rlabel metal1 4204 4562 4236 4578 0 FILL_1__1314_.gnd
rlabel nsubstratencontact 4204 4808 4204 4808 0 FILL_0__1314_.vdd
rlabel metal1 4184 4562 4216 4578 0 FILL_0__1314_.gnd
rlabel metal1 4224 4562 4336 4578 0 _1314_.gnd
rlabel metal1 4224 4802 4336 4818 0 _1314_.vdd
rlabel metal2 4313 4653 4327 4667 0 _1314_.A
rlabel metal2 4253 4653 4267 4667 0 _1314_.Y
rlabel metal2 4273 4693 4287 4707 0 _1314_.B
rlabel nsubstratencontact 4384 4808 4384 4808 0 FILL_2__1305_.vdd
rlabel metal1 4364 4562 4396 4578 0 FILL_2__1305_.gnd
rlabel nsubstratencontact 4364 4808 4364 4808 0 FILL_1__1305_.vdd
rlabel metal1 4344 4562 4376 4578 0 FILL_1__1305_.gnd
rlabel nsubstratencontact 4344 4808 4344 4808 0 FILL_0__1305_.vdd
rlabel metal1 4324 4562 4356 4578 0 FILL_0__1305_.gnd
rlabel metal1 4384 4562 4496 4578 0 _1305_.gnd
rlabel metal1 4384 4802 4496 4818 0 _1305_.vdd
rlabel metal2 4473 4673 4487 4687 0 _1305_.A
rlabel metal2 4453 4693 4467 4707 0 _1305_.B
rlabel metal2 4433 4673 4447 4687 0 _1305_.C
rlabel metal2 4413 4693 4427 4707 0 _1305_.Y
rlabel nsubstratencontact 4516 4808 4516 4808 0 FILL_1__1388_.vdd
rlabel metal1 4504 4562 4536 4578 0 FILL_1__1388_.gnd
rlabel nsubstratencontact 4496 4808 4496 4808 0 FILL_0__1388_.vdd
rlabel metal1 4484 4562 4516 4578 0 FILL_0__1388_.gnd
rlabel metal1 4524 4562 4636 4578 0 _1388_.gnd
rlabel metal1 4524 4802 4636 4818 0 _1388_.vdd
rlabel metal2 4533 4673 4547 4687 0 _1388_.A
rlabel metal2 4553 4693 4567 4707 0 _1388_.B
rlabel metal2 4573 4673 4587 4687 0 _1388_.C
rlabel metal2 4593 4693 4607 4707 0 _1388_.Y
rlabel metal1 4664 4562 4736 4578 0 _1373_.gnd
rlabel metal1 4664 4802 4736 4818 0 _1373_.vdd
rlabel metal2 4673 4633 4687 4647 0 _1373_.A
rlabel metal2 4693 4673 4707 4687 0 _1373_.Y
rlabel metal1 5004 4562 5116 4578 0 _1629_.gnd
rlabel metal1 5004 4802 5116 4818 0 _1629_.vdd
rlabel metal2 5013 4653 5027 4667 0 _1629_.A
rlabel metal2 5033 4673 5047 4687 0 _1629_.B
rlabel metal2 5073 4673 5087 4687 0 _1629_.C
rlabel metal2 5053 4653 5067 4667 0 _1629_.Y
rlabel metal1 4724 4562 4976 4578 0 _1673_.gnd
rlabel metal1 4724 4802 4976 4818 0 _1673_.vdd
rlabel metal2 4873 4653 4887 4667 0 _1673_.D
rlabel metal2 4833 4653 4847 4667 0 _1673_.CLK
rlabel metal2 4753 4653 4767 4667 0 _1673_.Q
rlabel nsubstratencontact 4636 4808 4636 4808 0 FILL_0__1373_.vdd
rlabel metal1 4624 4562 4656 4578 0 FILL_0__1373_.gnd
rlabel nsubstratencontact 4976 4808 4976 4808 0 FILL_0__1629_.vdd
rlabel metal1 4964 4562 4996 4578 0 FILL_0__1629_.gnd
rlabel nsubstratencontact 4656 4808 4656 4808 0 FILL_1__1373_.vdd
rlabel metal1 4644 4562 4676 4578 0 FILL_1__1373_.gnd
rlabel nsubstratencontact 4996 4808 4996 4808 0 FILL_1__1629_.vdd
rlabel metal1 4984 4562 5016 4578 0 FILL_1__1629_.gnd
rlabel nsubstratencontact 5136 4808 5136 4808 0 FILL_1__1628_.vdd
rlabel metal1 5124 4562 5156 4578 0 FILL_1__1628_.gnd
rlabel nsubstratencontact 5116 4808 5116 4808 0 FILL_0__1628_.vdd
rlabel metal1 5104 4562 5136 4578 0 FILL_0__1628_.gnd
rlabel metal1 5144 4562 5236 4578 0 _1628_.gnd
rlabel metal1 5144 4802 5236 4818 0 _1628_.vdd
rlabel metal2 5153 4693 5167 4707 0 _1628_.A
rlabel metal2 5193 4693 5207 4707 0 _1628_.B
rlabel metal2 5173 4673 5187 4687 0 _1628_.Y
rlabel nsubstratencontact 5256 4808 5256 4808 0 FILL_1__1556_.vdd
rlabel metal1 5244 4562 5276 4578 0 FILL_1__1556_.gnd
rlabel nsubstratencontact 5236 4808 5236 4808 0 FILL_0__1556_.vdd
rlabel metal1 5224 4562 5256 4578 0 FILL_0__1556_.gnd
rlabel nsubstratencontact 5376 4808 5376 4808 0 FILL_1__1553_.vdd
rlabel metal1 5364 4562 5396 4578 0 FILL_1__1553_.gnd
rlabel nsubstratencontact 5356 4808 5356 4808 0 FILL_0__1553_.vdd
rlabel metal1 5344 4562 5376 4578 0 FILL_0__1553_.gnd
rlabel metal1 5264 4562 5356 4578 0 _1556_.gnd
rlabel metal1 5264 4802 5356 4818 0 _1556_.vdd
rlabel metal2 5273 4693 5287 4707 0 _1556_.A
rlabel metal2 5313 4693 5327 4707 0 _1556_.B
rlabel metal2 5293 4673 5307 4687 0 _1556_.Y
rlabel nsubstratencontact 5396 4808 5396 4808 0 FILL_2__1553_.vdd
rlabel metal1 5384 4562 5416 4578 0 FILL_2__1553_.gnd
rlabel metal1 5404 4562 5496 4578 0 _1553_.gnd
rlabel metal1 5404 4802 5496 4818 0 _1553_.vdd
rlabel metal2 5413 4693 5427 4707 0 _1553_.A
rlabel metal2 5453 4693 5467 4707 0 _1553_.B
rlabel metal2 5433 4673 5447 4687 0 _1553_.Y
rlabel nsubstratencontact 5516 4808 5516 4808 0 FILL_1__1552_.vdd
rlabel metal1 5504 4562 5536 4578 0 FILL_1__1552_.gnd
rlabel nsubstratencontact 5496 4808 5496 4808 0 FILL_0__1552_.vdd
rlabel metal1 5484 4562 5516 4578 0 FILL_0__1552_.gnd
rlabel metal1 5524 4562 5616 4578 0 _1552_.gnd
rlabel metal1 5524 4802 5616 4818 0 _1552_.vdd
rlabel metal2 5533 4693 5547 4707 0 _1552_.A
rlabel metal2 5573 4693 5587 4707 0 _1552_.B
rlabel metal2 5553 4673 5567 4687 0 _1552_.Y
rlabel metal1 5644 4562 5756 4578 0 _1555_.gnd
rlabel metal1 5644 4802 5756 4818 0 _1555_.vdd
rlabel metal2 5733 4673 5747 4687 0 _1555_.A
rlabel metal2 5713 4693 5727 4707 0 _1555_.B
rlabel metal2 5693 4673 5707 4687 0 _1555_.C
rlabel metal2 5673 4693 5687 4707 0 _1555_.Y
rlabel nsubstratencontact 5756 4808 5756 4808 0 FILL86250x68550.vdd
rlabel metal1 5744 4562 5776 4578 0 FILL86250x68550.gnd
rlabel nsubstratencontact 5776 4808 5776 4808 0 FILL86550x68550.vdd
rlabel metal1 5764 4562 5796 4578 0 FILL86550x68550.gnd
rlabel nsubstratencontact 5796 4808 5796 4808 0 FILL86850x68550.vdd
rlabel metal1 5784 4562 5816 4578 0 FILL86850x68550.gnd
rlabel nsubstratencontact 5624 4808 5624 4808 0 FILL_0__1555_.vdd
rlabel metal1 5604 4562 5636 4578 0 FILL_0__1555_.gnd
rlabel nsubstratencontact 5644 4808 5644 4808 0 FILL_1__1555_.vdd
rlabel metal1 5624 4562 5656 4578 0 FILL_1__1555_.gnd
rlabel nsubstratencontact 44 4812 44 4812 0 FILL_1__994_.vdd
rlabel metal1 24 5042 56 5058 0 FILL_1__994_.gnd
rlabel nsubstratencontact 24 4812 24 4812 0 FILL_0__994_.vdd
rlabel metal1 4 5042 36 5058 0 FILL_0__994_.gnd
rlabel metal1 44 5042 156 5058 0 _994_.gnd
rlabel metal1 44 4802 156 4818 0 _994_.vdd
rlabel metal2 133 4953 147 4967 0 _994_.A
rlabel metal2 113 4933 127 4947 0 _994_.B
rlabel metal2 73 4933 87 4947 0 _994_.C
rlabel metal2 93 4953 107 4967 0 _994_.Y
rlabel nsubstratencontact 184 4812 184 4812 0 FILL_1__988_.vdd
rlabel metal1 164 5042 196 5058 0 FILL_1__988_.gnd
rlabel nsubstratencontact 164 4812 164 4812 0 FILL_0__988_.vdd
rlabel metal1 144 5042 176 5058 0 FILL_0__988_.gnd
rlabel metal1 184 5042 296 5058 0 _988_.gnd
rlabel metal1 184 4802 296 4818 0 _988_.vdd
rlabel metal2 273 4933 287 4947 0 _988_.A
rlabel metal2 253 4913 267 4927 0 _988_.B
rlabel metal2 233 4933 247 4947 0 _988_.C
rlabel metal2 213 4913 227 4927 0 _988_.Y
rlabel nsubstratencontact 316 4812 316 4812 0 FILL_1__1139_.vdd
rlabel metal1 304 5042 336 5058 0 FILL_1__1139_.gnd
rlabel nsubstratencontact 296 4812 296 4812 0 FILL_0__1139_.vdd
rlabel metal1 284 5042 316 5058 0 FILL_0__1139_.gnd
rlabel metal1 324 5042 436 5058 0 _1139_.gnd
rlabel metal1 324 4802 436 4818 0 _1139_.vdd
rlabel metal2 333 4933 347 4947 0 _1139_.A
rlabel metal2 353 4913 367 4927 0 _1139_.B
rlabel metal2 373 4933 387 4947 0 _1139_.C
rlabel metal2 393 4913 407 4927 0 _1139_.Y
rlabel nsubstratencontact 456 4812 456 4812 0 FILL_1__1138_.vdd
rlabel metal1 444 5042 476 5058 0 FILL_1__1138_.gnd
rlabel nsubstratencontact 436 4812 436 4812 0 FILL_0__1138_.vdd
rlabel metal1 424 5042 456 5058 0 FILL_0__1138_.gnd
rlabel metal1 464 5042 576 5058 0 _1138_.gnd
rlabel metal1 464 4802 576 4818 0 _1138_.vdd
rlabel metal2 473 4953 487 4967 0 _1138_.A
rlabel metal2 493 4933 507 4947 0 _1138_.B
rlabel metal2 533 4933 547 4947 0 _1138_.C
rlabel metal2 513 4953 527 4967 0 _1138_.Y
rlabel nsubstratencontact 604 4812 604 4812 0 FILL_1__987_.vdd
rlabel metal1 584 5042 616 5058 0 FILL_1__987_.gnd
rlabel nsubstratencontact 584 4812 584 4812 0 FILL_0__987_.vdd
rlabel metal1 564 5042 596 5058 0 FILL_0__987_.gnd
rlabel metal1 604 5042 696 5058 0 _987_.gnd
rlabel metal1 604 4802 696 4818 0 _987_.vdd
rlabel metal2 673 4913 687 4927 0 _987_.A
rlabel metal2 633 4913 647 4927 0 _987_.B
rlabel metal2 653 4933 667 4947 0 _987_.Y
rlabel nsubstratencontact 724 4812 724 4812 0 FILL_1__957_.vdd
rlabel metal1 704 5042 736 5058 0 FILL_1__957_.gnd
rlabel nsubstratencontact 704 4812 704 4812 0 FILL_0__957_.vdd
rlabel metal1 684 5042 716 5058 0 FILL_0__957_.gnd
rlabel metal1 724 5042 836 5058 0 _957_.gnd
rlabel metal1 724 4802 836 4818 0 _957_.vdd
rlabel metal2 813 4953 827 4967 0 _957_.A
rlabel metal2 793 4933 807 4947 0 _957_.B
rlabel metal2 753 4933 767 4947 0 _957_.C
rlabel metal2 773 4953 787 4967 0 _957_.Y
rlabel nsubstratencontact 864 4812 864 4812 0 FILL_1__949_.vdd
rlabel metal1 844 5042 876 5058 0 FILL_1__949_.gnd
rlabel nsubstratencontact 844 4812 844 4812 0 FILL_0__949_.vdd
rlabel metal1 824 5042 856 5058 0 FILL_0__949_.gnd
rlabel metal1 864 5042 976 5058 0 _949_.gnd
rlabel metal1 864 4802 976 4818 0 _949_.vdd
rlabel metal2 953 4953 967 4967 0 _949_.A
rlabel metal2 933 4933 947 4947 0 _949_.B
rlabel metal2 893 4933 907 4947 0 _949_.C
rlabel metal2 913 4953 927 4967 0 _949_.Y
rlabel nsubstratencontact 1004 4812 1004 4812 0 FILL_1__971_.vdd
rlabel metal1 984 5042 1016 5058 0 FILL_1__971_.gnd
rlabel nsubstratencontact 984 4812 984 4812 0 FILL_0__971_.vdd
rlabel metal1 964 5042 996 5058 0 FILL_0__971_.gnd
rlabel metal1 1004 5042 1116 5058 0 _971_.gnd
rlabel metal1 1004 4802 1116 4818 0 _971_.vdd
rlabel metal2 1093 4933 1107 4947 0 _971_.A
rlabel metal2 1073 4973 1087 4987 0 _971_.B
rlabel metal2 1053 4933 1067 4947 0 _971_.C
rlabel metal2 1033 4953 1047 4967 0 _971_.Y
rlabel nsubstratencontact 1144 4812 1144 4812 0 FILL_1__1131_.vdd
rlabel metal1 1124 5042 1156 5058 0 FILL_1__1131_.gnd
rlabel nsubstratencontact 1124 4812 1124 4812 0 FILL_0__1131_.vdd
rlabel metal1 1104 5042 1136 5058 0 FILL_0__1131_.gnd
rlabel nsubstratencontact 1264 4812 1264 4812 0 FILL_0__948_.vdd
rlabel metal1 1244 5042 1276 5058 0 FILL_0__948_.gnd
rlabel metal1 1144 5042 1256 5058 0 _1131_.gnd
rlabel metal1 1144 4802 1256 4818 0 _1131_.vdd
rlabel metal2 1233 4953 1247 4967 0 _1131_.A
rlabel metal2 1213 4933 1227 4947 0 _1131_.B
rlabel metal2 1173 4933 1187 4947 0 _1131_.C
rlabel metal2 1193 4953 1207 4967 0 _1131_.Y
rlabel nsubstratencontact 1384 4812 1384 4812 0 FILL_1__1417_.vdd
rlabel metal1 1364 5042 1396 5058 0 FILL_1__1417_.gnd
rlabel nsubstratencontact 1284 4812 1284 4812 0 FILL_1__948_.vdd
rlabel metal1 1264 5042 1296 5058 0 FILL_1__948_.gnd
rlabel nsubstratencontact 1364 4812 1364 4812 0 FILL_0__1417_.vdd
rlabel metal1 1344 5042 1376 5058 0 FILL_0__1417_.gnd
rlabel metal1 1384 5042 1476 5058 0 _1417_.gnd
rlabel metal1 1384 4802 1476 4818 0 _1417_.vdd
rlabel metal2 1453 4913 1467 4927 0 _1417_.A
rlabel metal2 1413 4913 1427 4927 0 _1417_.B
rlabel metal2 1433 4933 1447 4947 0 _1417_.Y
rlabel metal1 1284 5042 1356 5058 0 _948_.gnd
rlabel metal1 1284 4802 1356 4818 0 _948_.vdd
rlabel metal2 1333 4973 1347 4987 0 _948_.A
rlabel metal2 1313 4933 1327 4947 0 _948_.Y
rlabel nsubstratencontact 1524 4812 1524 4812 0 FILL_2__1416_.vdd
rlabel metal1 1504 5042 1536 5058 0 FILL_2__1416_.gnd
rlabel nsubstratencontact 1504 4812 1504 4812 0 FILL_1__1416_.vdd
rlabel metal1 1484 5042 1516 5058 0 FILL_1__1416_.gnd
rlabel nsubstratencontact 1484 4812 1484 4812 0 FILL_0__1416_.vdd
rlabel metal1 1464 5042 1496 5058 0 FILL_0__1416_.gnd
rlabel nsubstratencontact 1644 4812 1644 4812 0 FILL_0__1415_.vdd
rlabel metal1 1624 5042 1656 5058 0 FILL_0__1415_.gnd
rlabel metal1 1524 5042 1636 5058 0 _1416_.gnd
rlabel metal1 1524 4802 1636 4818 0 _1416_.vdd
rlabel metal2 1613 4933 1627 4947 0 _1416_.A
rlabel metal2 1593 4913 1607 4927 0 _1416_.B
rlabel metal2 1573 4933 1587 4947 0 _1416_.C
rlabel metal2 1553 4913 1567 4927 0 _1416_.Y
rlabel nsubstratencontact 1664 4812 1664 4812 0 FILL_1__1415_.vdd
rlabel metal1 1644 5042 1676 5058 0 FILL_1__1415_.gnd
rlabel nsubstratencontact 1776 4812 1776 4812 0 FILL_0__1436_.vdd
rlabel metal1 1764 5042 1796 5058 0 FILL_0__1436_.gnd
rlabel metal1 1664 5042 1776 5058 0 _1415_.gnd
rlabel metal1 1664 4802 1776 4818 0 _1415_.vdd
rlabel metal2 1753 4953 1767 4967 0 _1415_.A
rlabel metal2 1733 4933 1747 4947 0 _1415_.B
rlabel metal2 1693 4933 1707 4947 0 _1415_.C
rlabel metal2 1713 4953 1727 4967 0 _1415_.Y
rlabel nsubstratencontact 1796 4812 1796 4812 0 FILL_1__1436_.vdd
rlabel metal1 1784 5042 1816 5058 0 FILL_1__1436_.gnd
rlabel metal1 1804 5042 1916 5058 0 _1436_.gnd
rlabel metal1 1804 4802 1916 4818 0 _1436_.vdd
rlabel metal2 1813 4933 1827 4947 0 _1436_.A
rlabel metal2 1833 4973 1847 4987 0 _1436_.B
rlabel metal2 1853 4933 1867 4947 0 _1436_.C
rlabel metal2 1873 4953 1887 4967 0 _1436_.Y
rlabel nsubstratencontact 1936 4812 1936 4812 0 FILL_1__1467_.vdd
rlabel metal1 1924 5042 1956 5058 0 FILL_1__1467_.gnd
rlabel nsubstratencontact 1916 4812 1916 4812 0 FILL_0__1467_.vdd
rlabel metal1 1904 5042 1936 5058 0 FILL_0__1467_.gnd
rlabel metal1 1944 5042 2036 5058 0 _1467_.gnd
rlabel metal1 1944 4802 2036 4818 0 _1467_.vdd
rlabel metal2 1953 4913 1967 4927 0 _1467_.A
rlabel metal2 1993 4913 2007 4927 0 _1467_.B
rlabel metal2 1973 4933 1987 4947 0 _1467_.Y
rlabel nsubstratencontact 2064 4812 2064 4812 0 FILL_1__1411_.vdd
rlabel metal1 2044 5042 2076 5058 0 FILL_1__1411_.gnd
rlabel nsubstratencontact 2044 4812 2044 4812 0 FILL_0__1411_.vdd
rlabel metal1 2024 5042 2056 5058 0 FILL_0__1411_.gnd
rlabel metal1 2064 5042 2176 5058 0 _1411_.gnd
rlabel metal1 2064 4802 2176 4818 0 _1411_.vdd
rlabel metal2 2153 4933 2167 4947 0 _1411_.A
rlabel metal2 2133 4973 2147 4987 0 _1411_.B
rlabel metal2 2113 4933 2127 4947 0 _1411_.C
rlabel metal2 2093 4953 2107 4967 0 _1411_.Y
rlabel nsubstratencontact 2224 4812 2224 4812 0 FILL_2__1409_.vdd
rlabel metal1 2204 5042 2236 5058 0 FILL_2__1409_.gnd
rlabel nsubstratencontact 2204 4812 2204 4812 0 FILL_1__1409_.vdd
rlabel metal1 2184 5042 2216 5058 0 FILL_1__1409_.gnd
rlabel nsubstratencontact 2184 4812 2184 4812 0 FILL_0__1409_.vdd
rlabel metal1 2164 5042 2196 5058 0 FILL_0__1409_.gnd
rlabel metal1 2224 5042 2296 5058 0 _1409_.gnd
rlabel metal1 2224 4802 2296 4818 0 _1409_.vdd
rlabel metal2 2273 4973 2287 4987 0 _1409_.A
rlabel metal2 2253 4933 2267 4947 0 _1409_.Y
rlabel nsubstratencontact 2324 4812 2324 4812 0 FILL_1__1410_.vdd
rlabel metal1 2304 5042 2336 5058 0 FILL_1__1410_.gnd
rlabel nsubstratencontact 2304 4812 2304 4812 0 FILL_0__1410_.vdd
rlabel metal1 2284 5042 2316 5058 0 FILL_0__1410_.gnd
rlabel metal1 2324 5042 2436 5058 0 _1410_.gnd
rlabel metal1 2324 4802 2436 4818 0 _1410_.vdd
rlabel metal2 2413 4953 2427 4967 0 _1410_.A
rlabel metal2 2393 4933 2407 4947 0 _1410_.B
rlabel metal2 2353 4933 2367 4947 0 _1410_.C
rlabel metal2 2373 4953 2387 4967 0 _1410_.Y
rlabel nsubstratencontact 2464 4812 2464 4812 0 FILL_1__1408_.vdd
rlabel metal1 2444 5042 2476 5058 0 FILL_1__1408_.gnd
rlabel nsubstratencontact 2444 4812 2444 4812 0 FILL_0__1408_.vdd
rlabel metal1 2424 5042 2456 5058 0 FILL_0__1408_.gnd
rlabel metal1 2464 5042 2576 5058 0 _1408_.gnd
rlabel metal1 2464 4802 2576 4818 0 _1408_.vdd
rlabel metal2 2553 4933 2567 4947 0 _1408_.A
rlabel metal2 2533 4913 2547 4927 0 _1408_.B
rlabel metal2 2513 4933 2527 4947 0 _1408_.C
rlabel metal2 2493 4913 2507 4927 0 _1408_.Y
rlabel nsubstratencontact 2604 4812 2604 4812 0 FILL_1__1407_.vdd
rlabel metal1 2584 5042 2616 5058 0 FILL_1__1407_.gnd
rlabel nsubstratencontact 2584 4812 2584 4812 0 FILL_0__1407_.vdd
rlabel metal1 2564 5042 2596 5058 0 FILL_0__1407_.gnd
rlabel metal1 2604 5042 2676 5058 0 _1407_.gnd
rlabel metal1 2604 4802 2676 4818 0 _1407_.vdd
rlabel metal2 2653 4973 2667 4987 0 _1407_.A
rlabel metal2 2633 4933 2647 4947 0 _1407_.Y
rlabel nsubstratencontact 2724 4812 2724 4812 0 FILL_2__1370_.vdd
rlabel metal1 2704 5042 2736 5058 0 FILL_2__1370_.gnd
rlabel nsubstratencontact 2704 4812 2704 4812 0 FILL_1__1370_.vdd
rlabel metal1 2684 5042 2716 5058 0 FILL_1__1370_.gnd
rlabel nsubstratencontact 2684 4812 2684 4812 0 FILL_0__1370_.vdd
rlabel metal1 2664 5042 2696 5058 0 FILL_0__1370_.gnd
rlabel metal1 2724 5042 2816 5058 0 _1370_.gnd
rlabel metal1 2724 4802 2816 4818 0 _1370_.vdd
rlabel metal2 2793 4913 2807 4927 0 _1370_.A
rlabel metal2 2753 4913 2767 4927 0 _1370_.B
rlabel metal2 2773 4933 2787 4947 0 _1370_.Y
rlabel nsubstratencontact 2836 4812 2836 4812 0 FILL_1__1371_.vdd
rlabel metal1 2824 5042 2856 5058 0 FILL_1__1371_.gnd
rlabel nsubstratencontact 2816 4812 2816 4812 0 FILL_0__1371_.vdd
rlabel metal1 2804 5042 2836 5058 0 FILL_0__1371_.gnd
rlabel metal1 2844 5042 2916 5058 0 _1371_.gnd
rlabel metal1 2844 4802 2916 4818 0 _1371_.vdd
rlabel metal2 2853 4973 2867 4987 0 _1371_.A
rlabel metal2 2873 4933 2887 4947 0 _1371_.Y
rlabel nsubstratencontact 2936 4812 2936 4812 0 FILL_1__1380_.vdd
rlabel metal1 2924 5042 2956 5058 0 FILL_1__1380_.gnd
rlabel nsubstratencontact 2916 4812 2916 4812 0 FILL_0__1380_.vdd
rlabel metal1 2904 5042 2936 5058 0 FILL_0__1380_.gnd
rlabel metal1 2944 5042 3056 5058 0 _1380_.gnd
rlabel metal1 2944 4802 3056 4818 0 _1380_.vdd
rlabel metal2 2953 4933 2967 4947 0 _1380_.A
rlabel metal2 2973 4913 2987 4927 0 _1380_.B
rlabel metal2 2993 4933 3007 4947 0 _1380_.C
rlabel metal2 3013 4913 3027 4927 0 _1380_.Y
rlabel nsubstratencontact 3084 4812 3084 4812 0 FILL_1__1379_.vdd
rlabel metal1 3064 5042 3096 5058 0 FILL_1__1379_.gnd
rlabel nsubstratencontact 3064 4812 3064 4812 0 FILL_0__1379_.vdd
rlabel metal1 3044 5042 3076 5058 0 FILL_0__1379_.gnd
rlabel metal1 3084 5042 3196 5058 0 _1379_.gnd
rlabel metal1 3084 4802 3196 4818 0 _1379_.vdd
rlabel metal2 3173 4953 3187 4967 0 _1379_.A
rlabel metal2 3153 4933 3167 4947 0 _1379_.B
rlabel metal2 3113 4933 3127 4947 0 _1379_.C
rlabel metal2 3133 4953 3147 4967 0 _1379_.Y
rlabel nsubstratencontact 3224 4812 3224 4812 0 FILL_1__1377_.vdd
rlabel metal1 3204 5042 3236 5058 0 FILL_1__1377_.gnd
rlabel nsubstratencontact 3204 4812 3204 4812 0 FILL_0__1377_.vdd
rlabel metal1 3184 5042 3216 5058 0 FILL_0__1377_.gnd
rlabel metal1 3224 5042 3336 5058 0 _1377_.gnd
rlabel metal1 3224 4802 3336 4818 0 _1377_.vdd
rlabel metal2 3313 4953 3327 4967 0 _1377_.A
rlabel metal2 3293 4933 3307 4947 0 _1377_.B
rlabel metal2 3253 4933 3267 4947 0 _1377_.C
rlabel metal2 3273 4953 3287 4967 0 _1377_.Y
rlabel nsubstratencontact 3364 4812 3364 4812 0 FILL_1__1378_.vdd
rlabel metal1 3344 5042 3376 5058 0 FILL_1__1378_.gnd
rlabel nsubstratencontact 3344 4812 3344 4812 0 FILL_0__1378_.vdd
rlabel metal1 3324 5042 3356 5058 0 FILL_0__1378_.gnd
rlabel metal1 3364 5042 3476 5058 0 _1378_.gnd
rlabel metal1 3364 4802 3476 4818 0 _1378_.vdd
rlabel metal2 3453 4933 3467 4947 0 _1378_.A
rlabel metal2 3433 4973 3447 4987 0 _1378_.B
rlabel metal2 3413 4933 3427 4947 0 _1378_.C
rlabel metal2 3393 4953 3407 4967 0 _1378_.Y
rlabel nsubstratencontact 3496 4812 3496 4812 0 FILL_1__1309_.vdd
rlabel metal1 3484 5042 3516 5058 0 FILL_1__1309_.gnd
rlabel nsubstratencontact 3476 4812 3476 4812 0 FILL_0__1309_.vdd
rlabel metal1 3464 5042 3496 5058 0 FILL_0__1309_.gnd
rlabel metal1 3504 5042 3616 5058 0 _1309_.gnd
rlabel metal1 3504 4802 3616 4818 0 _1309_.vdd
rlabel metal2 3513 4973 3527 4987 0 _1309_.A
rlabel metal2 3533 4953 3547 4967 0 _1309_.B
rlabel metal2 3573 4933 3587 4947 0 _1309_.Y
rlabel nsubstratencontact 3644 4812 3644 4812 0 FILL_1__1374_.vdd
rlabel metal1 3624 5042 3656 5058 0 FILL_1__1374_.gnd
rlabel nsubstratencontact 3624 4812 3624 4812 0 FILL_0__1374_.vdd
rlabel metal1 3604 5042 3636 5058 0 FILL_0__1374_.gnd
rlabel metal1 3644 5042 3736 5058 0 _1374_.gnd
rlabel metal1 3644 4802 3736 4818 0 _1374_.vdd
rlabel metal2 3673 4953 3687 4967 0 _1374_.B
rlabel metal2 3713 4953 3727 4967 0 _1374_.A
rlabel metal2 3693 4973 3707 4987 0 _1374_.Y
rlabel nsubstratencontact 3764 4812 3764 4812 0 FILL_1__1307_.vdd
rlabel metal1 3744 5042 3776 5058 0 FILL_1__1307_.gnd
rlabel nsubstratencontact 3744 4812 3744 4812 0 FILL_0__1307_.vdd
rlabel metal1 3724 5042 3756 5058 0 FILL_0__1307_.gnd
rlabel metal1 3764 5042 3876 5058 0 _1307_.gnd
rlabel metal1 3764 4802 3876 4818 0 _1307_.vdd
rlabel metal2 3853 4933 3867 4947 0 _1307_.A
rlabel metal2 3833 4913 3847 4927 0 _1307_.B
rlabel metal2 3813 4933 3827 4947 0 _1307_.C
rlabel metal2 3793 4913 3807 4927 0 _1307_.Y
rlabel nsubstratencontact 3904 4812 3904 4812 0 FILL_1__923_.vdd
rlabel metal1 3884 5042 3916 5058 0 FILL_1__923_.gnd
rlabel nsubstratencontact 3884 4812 3884 4812 0 FILL_0__923_.vdd
rlabel metal1 3864 5042 3896 5058 0 FILL_0__923_.gnd
rlabel metal1 3904 5042 3976 5058 0 _923_.gnd
rlabel metal1 3904 4802 3976 4818 0 _923_.vdd
rlabel metal2 3953 4973 3967 4987 0 _923_.A
rlabel metal2 3933 4933 3947 4947 0 _923_.Y
rlabel nsubstratencontact 3996 4812 3996 4812 0 FILL_1__1385_.vdd
rlabel metal1 3984 5042 4016 5058 0 FILL_1__1385_.gnd
rlabel nsubstratencontact 3976 4812 3976 4812 0 FILL_0__1385_.vdd
rlabel metal1 3964 5042 3996 5058 0 FILL_0__1385_.gnd
rlabel metal1 4004 5042 4116 5058 0 _1385_.gnd
rlabel metal1 4004 4802 4116 4818 0 _1385_.vdd
rlabel metal2 4013 4933 4027 4947 0 _1385_.A
rlabel metal2 4033 4913 4047 4927 0 _1385_.B
rlabel metal2 4053 4933 4067 4947 0 _1385_.C
rlabel metal2 4073 4913 4087 4927 0 _1385_.Y
rlabel nsubstratencontact 4136 4812 4136 4812 0 FILL_1__1387_.vdd
rlabel metal1 4124 5042 4156 5058 0 FILL_1__1387_.gnd
rlabel nsubstratencontact 4116 4812 4116 4812 0 FILL_0__1387_.vdd
rlabel metal1 4104 5042 4136 5058 0 FILL_0__1387_.gnd
rlabel metal1 4144 5042 4256 5058 0 _1387_.gnd
rlabel metal1 4144 4802 4256 4818 0 _1387_.vdd
rlabel metal2 4153 4933 4167 4947 0 _1387_.A
rlabel metal2 4173 4913 4187 4927 0 _1387_.B
rlabel metal2 4193 4933 4207 4947 0 _1387_.C
rlabel metal2 4213 4913 4227 4927 0 _1387_.Y
rlabel nsubstratencontact 4284 4812 4284 4812 0 FILL_1__1394_.vdd
rlabel metal1 4264 5042 4296 5058 0 FILL_1__1394_.gnd
rlabel nsubstratencontact 4264 4812 4264 4812 0 FILL_0__1394_.vdd
rlabel metal1 4244 5042 4276 5058 0 FILL_0__1394_.gnd
rlabel metal1 4284 5042 4396 5058 0 _1394_.gnd
rlabel metal1 4284 4802 4396 4818 0 _1394_.vdd
rlabel metal2 4373 4953 4387 4967 0 _1394_.A
rlabel metal2 4313 4953 4327 4967 0 _1394_.Y
rlabel metal2 4333 4913 4347 4927 0 _1394_.B
rlabel nsubstratencontact 4416 4812 4416 4812 0 FILL_1__1389_.vdd
rlabel metal1 4404 5042 4436 5058 0 FILL_1__1389_.gnd
rlabel nsubstratencontact 4396 4812 4396 4812 0 FILL_0__1389_.vdd
rlabel metal1 4384 5042 4416 5058 0 FILL_0__1389_.gnd
rlabel nsubstratencontact 4436 4812 4436 4812 0 FILL_2__1389_.vdd
rlabel metal1 4424 5042 4456 5058 0 FILL_2__1389_.gnd
rlabel metal1 4444 5042 4556 5058 0 _1389_.gnd
rlabel metal1 4444 4802 4556 4818 0 _1389_.vdd
rlabel metal2 4453 4973 4467 4987 0 _1389_.A
rlabel metal2 4473 4953 4487 4967 0 _1389_.B
rlabel metal2 4513 4933 4527 4947 0 _1389_.Y
rlabel nsubstratencontact 4556 4812 4556 4812 0 FILL_0__1393_.vdd
rlabel metal1 4544 5042 4576 5058 0 FILL_0__1393_.gnd
rlabel metal1 4704 5042 4816 5058 0 _1391_.gnd
rlabel metal1 4704 4802 4816 4818 0 _1391_.vdd
rlabel metal2 4793 4953 4807 4967 0 _1391_.A
rlabel metal2 4773 4933 4787 4947 0 _1391_.B
rlabel metal2 4733 4933 4747 4947 0 _1391_.C
rlabel metal2 4753 4953 4767 4967 0 _1391_.Y
rlabel metal1 4584 5042 4676 5058 0 _1393_.gnd
rlabel metal1 4584 4802 4676 4818 0 _1393_.vdd
rlabel metal2 4633 4953 4647 4967 0 _1393_.B
rlabel metal2 4593 4953 4607 4967 0 _1393_.A
rlabel metal2 4613 4973 4627 4987 0 _1393_.Y
rlabel metal1 4804 5042 5056 5058 0 _1676_.gnd
rlabel metal1 4804 4802 5056 4818 0 _1676_.vdd
rlabel metal2 4953 4953 4967 4967 0 _1676_.D
rlabel metal2 4913 4953 4927 4967 0 _1676_.CLK
rlabel metal2 4833 4953 4847 4967 0 _1676_.Q
rlabel nsubstratencontact 4684 4812 4684 4812 0 FILL_0__1391_.vdd
rlabel metal1 4664 5042 4696 5058 0 FILL_0__1391_.gnd
rlabel nsubstratencontact 5056 4812 5056 4812 0 FILL_0__1635_.vdd
rlabel metal1 5044 5042 5076 5058 0 FILL_0__1635_.gnd
rlabel nsubstratencontact 4704 4812 4704 4812 0 FILL_1__1391_.vdd
rlabel metal1 4684 5042 4716 5058 0 FILL_1__1391_.gnd
rlabel nsubstratencontact 4576 4812 4576 4812 0 FILL_1__1393_.vdd
rlabel metal1 4564 5042 4596 5058 0 FILL_1__1393_.gnd
rlabel metal1 5464 5042 5556 5058 0 _1634_.gnd
rlabel metal1 5464 4802 5556 4818 0 _1634_.vdd
rlabel metal2 5533 4913 5547 4927 0 _1634_.A
rlabel metal2 5493 4913 5507 4927 0 _1634_.B
rlabel metal2 5513 4933 5527 4947 0 _1634_.Y
rlabel metal1 5084 5042 5196 5058 0 _1635_.gnd
rlabel metal1 5084 4802 5196 4818 0 _1635_.vdd
rlabel metal2 5093 4953 5107 4967 0 _1635_.A
rlabel metal2 5113 4933 5127 4947 0 _1635_.B
rlabel metal2 5153 4933 5167 4947 0 _1635_.C
rlabel metal2 5133 4953 5147 4967 0 _1635_.Y
rlabel metal1 5184 5042 5436 5058 0 _1683_.gnd
rlabel metal1 5184 4802 5436 4818 0 _1683_.vdd
rlabel metal2 5333 4953 5347 4967 0 _1683_.D
rlabel metal2 5293 4953 5307 4967 0 _1683_.CLK
rlabel metal2 5213 4953 5227 4967 0 _1683_.Q
rlabel nsubstratencontact 5556 4812 5556 4812 0 FILL_0__1616_.vdd
rlabel metal1 5544 5042 5576 5058 0 FILL_0__1616_.gnd
rlabel nsubstratencontact 5444 4812 5444 4812 0 FILL_0__1634_.vdd
rlabel metal1 5424 5042 5456 5058 0 FILL_0__1634_.gnd
rlabel nsubstratencontact 5464 4812 5464 4812 0 FILL_1__1634_.vdd
rlabel metal1 5444 5042 5476 5058 0 FILL_1__1634_.gnd
rlabel nsubstratencontact 5076 4812 5076 4812 0 FILL_1__1635_.vdd
rlabel metal1 5064 5042 5096 5058 0 FILL_1__1635_.gnd
rlabel metal1 5584 5042 5676 5058 0 _1616_.gnd
rlabel metal1 5584 4802 5676 4818 0 _1616_.vdd
rlabel metal2 5593 4913 5607 4927 0 _1616_.A
rlabel metal2 5633 4913 5647 4927 0 _1616_.B
rlabel metal2 5613 4933 5627 4947 0 _1616_.Y
rlabel metal1 5724 5042 5816 5058 0 _1651_.gnd
rlabel metal1 5724 4802 5816 4818 0 _1651_.vdd
rlabel metal2 5733 4913 5747 4927 0 _1651_.A
rlabel metal2 5773 4913 5787 4927 0 _1651_.B
rlabel metal2 5753 4933 5767 4947 0 _1651_.Y
rlabel nsubstratencontact 5676 4812 5676 4812 0 FILL_0__1651_.vdd
rlabel metal1 5664 5042 5696 5058 0 FILL_0__1651_.gnd
rlabel nsubstratencontact 5576 4812 5576 4812 0 FILL_1__1616_.vdd
rlabel metal1 5564 5042 5596 5058 0 FILL_1__1616_.gnd
rlabel nsubstratencontact 5696 4812 5696 4812 0 FILL_1__1651_.vdd
rlabel metal1 5684 5042 5716 5058 0 FILL_1__1651_.gnd
rlabel nsubstratencontact 5716 4812 5716 4812 0 FILL_2__1651_.vdd
rlabel metal1 5704 5042 5736 5058 0 FILL_2__1651_.gnd
rlabel nsubstratencontact 44 5288 44 5288 0 FILL_1__995_.vdd
rlabel metal1 24 5042 56 5058 0 FILL_1__995_.gnd
rlabel nsubstratencontact 24 5288 24 5288 0 FILL_0__995_.vdd
rlabel metal1 4 5042 36 5058 0 FILL_0__995_.gnd
rlabel metal1 44 5042 156 5058 0 _995_.gnd
rlabel metal1 44 5282 156 5298 0 _995_.vdd
rlabel metal2 133 5153 147 5167 0 _995_.A
rlabel metal2 113 5173 127 5187 0 _995_.B
rlabel metal2 93 5153 107 5167 0 _995_.C
rlabel metal2 73 5173 87 5187 0 _995_.Y
rlabel nsubstratencontact 176 5288 176 5288 0 FILL_1__996_.vdd
rlabel metal1 164 5042 196 5058 0 FILL_1__996_.gnd
rlabel nsubstratencontact 156 5288 156 5288 0 FILL_0__996_.vdd
rlabel metal1 144 5042 176 5058 0 FILL_0__996_.gnd
rlabel metal1 184 5042 296 5058 0 _996_.gnd
rlabel metal1 184 5282 296 5298 0 _996_.vdd
rlabel metal2 193 5153 207 5167 0 _996_.A
rlabel metal2 213 5113 227 5127 0 _996_.B
rlabel metal2 233 5153 247 5167 0 _996_.C
rlabel metal2 253 5133 267 5147 0 _996_.Y
rlabel nsubstratencontact 316 5288 316 5288 0 FILL_1__1160_.vdd
rlabel metal1 304 5042 336 5058 0 FILL_1__1160_.gnd
rlabel nsubstratencontact 296 5288 296 5288 0 FILL_0__1160_.vdd
rlabel metal1 284 5042 316 5058 0 FILL_0__1160_.gnd
rlabel metal1 324 5042 396 5058 0 _1160_.gnd
rlabel metal1 324 5282 396 5298 0 _1160_.vdd
rlabel metal2 333 5113 347 5127 0 _1160_.A
rlabel metal2 353 5153 367 5167 0 _1160_.Y
rlabel nsubstratencontact 424 5288 424 5288 0 FILL_1__1159_.vdd
rlabel metal1 404 5042 436 5058 0 FILL_1__1159_.gnd
rlabel nsubstratencontact 404 5288 404 5288 0 FILL_0__1159_.vdd
rlabel metal1 384 5042 416 5058 0 FILL_0__1159_.gnd
rlabel metal1 424 5042 536 5058 0 _1159_.gnd
rlabel metal1 424 5282 536 5298 0 _1159_.vdd
rlabel metal2 513 5153 527 5167 0 _1159_.A
rlabel metal2 493 5173 507 5187 0 _1159_.B
rlabel metal2 473 5153 487 5167 0 _1159_.C
rlabel metal2 453 5173 467 5187 0 _1159_.Y
rlabel nsubstratencontact 556 5288 556 5288 0 FILL_1__1183_.vdd
rlabel metal1 544 5042 576 5058 0 FILL_1__1183_.gnd
rlabel nsubstratencontact 536 5288 536 5288 0 FILL_0__1183_.vdd
rlabel metal1 524 5042 556 5058 0 FILL_0__1183_.gnd
rlabel metal1 564 5042 676 5058 0 _1183_.gnd
rlabel metal1 564 5282 676 5298 0 _1183_.vdd
rlabel metal2 573 5153 587 5167 0 _1183_.A
rlabel metal2 593 5113 607 5127 0 _1183_.B
rlabel metal2 613 5153 627 5167 0 _1183_.C
rlabel metal2 633 5133 647 5147 0 _1183_.Y
rlabel nsubstratencontact 704 5288 704 5288 0 FILL_1__955_.vdd
rlabel metal1 684 5042 716 5058 0 FILL_1__955_.gnd
rlabel nsubstratencontact 684 5288 684 5288 0 FILL_0__955_.vdd
rlabel metal1 664 5042 696 5058 0 FILL_0__955_.gnd
rlabel metal1 704 5042 816 5058 0 _955_.gnd
rlabel metal1 704 5282 816 5298 0 _955_.vdd
rlabel metal2 793 5153 807 5167 0 _955_.A
rlabel metal2 773 5113 787 5127 0 _955_.B
rlabel metal2 753 5153 767 5167 0 _955_.C
rlabel metal2 733 5133 747 5147 0 _955_.Y
rlabel nsubstratencontact 836 5288 836 5288 0 FILL_1__950_.vdd
rlabel metal1 824 5042 856 5058 0 FILL_1__950_.gnd
rlabel nsubstratencontact 816 5288 816 5288 0 FILL_0__950_.vdd
rlabel metal1 804 5042 836 5058 0 FILL_0__950_.gnd
rlabel metal1 844 5042 956 5058 0 _950_.gnd
rlabel metal1 844 5282 956 5298 0 _950_.vdd
rlabel metal2 853 5153 867 5167 0 _950_.A
rlabel metal2 873 5173 887 5187 0 _950_.B
rlabel metal2 893 5153 907 5167 0 _950_.C
rlabel metal2 913 5173 927 5187 0 _950_.Y
rlabel nsubstratencontact 984 5288 984 5288 0 FILL_1__947_.vdd
rlabel metal1 964 5042 996 5058 0 FILL_1__947_.gnd
rlabel nsubstratencontact 964 5288 964 5288 0 FILL_0__947_.vdd
rlabel metal1 944 5042 976 5058 0 FILL_0__947_.gnd
rlabel metal1 984 5042 1096 5058 0 _947_.gnd
rlabel metal1 984 5282 1096 5298 0 _947_.vdd
rlabel metal2 1073 5153 1087 5167 0 _947_.A
rlabel metal2 1053 5173 1067 5187 0 _947_.B
rlabel metal2 1033 5153 1047 5167 0 _947_.C
rlabel metal2 1013 5173 1027 5187 0 _947_.Y
rlabel nsubstratencontact 1116 5288 1116 5288 0 FILL_1__939_.vdd
rlabel metal1 1104 5042 1136 5058 0 FILL_1__939_.gnd
rlabel nsubstratencontact 1096 5288 1096 5288 0 FILL_0__939_.vdd
rlabel metal1 1084 5042 1116 5058 0 FILL_0__939_.gnd
rlabel metal1 1124 5042 1196 5058 0 _939_.gnd
rlabel metal1 1124 5282 1196 5298 0 _939_.vdd
rlabel metal2 1133 5113 1147 5127 0 _939_.A
rlabel metal2 1153 5153 1167 5167 0 _939_.Y
rlabel nsubstratencontact 1224 5288 1224 5288 0 FILL_1__1132_.vdd
rlabel metal1 1204 5042 1236 5058 0 FILL_1__1132_.gnd
rlabel nsubstratencontact 1204 5288 1204 5288 0 FILL_0__1132_.vdd
rlabel metal1 1184 5042 1216 5058 0 FILL_0__1132_.gnd
rlabel metal1 1224 5042 1336 5058 0 _1132_.gnd
rlabel metal1 1224 5282 1336 5298 0 _1132_.vdd
rlabel metal2 1313 5153 1327 5167 0 _1132_.A
rlabel metal2 1293 5173 1307 5187 0 _1132_.B
rlabel metal2 1273 5153 1287 5167 0 _1132_.C
rlabel metal2 1253 5173 1267 5187 0 _1132_.Y
rlabel nsubstratencontact 1384 5288 1384 5288 0 FILL_2__953_.vdd
rlabel metal1 1364 5042 1396 5058 0 FILL_2__953_.gnd
rlabel nsubstratencontact 1364 5288 1364 5288 0 FILL_1__953_.vdd
rlabel metal1 1344 5042 1376 5058 0 FILL_1__953_.gnd
rlabel nsubstratencontact 1344 5288 1344 5288 0 FILL_0__953_.vdd
rlabel metal1 1324 5042 1356 5058 0 FILL_0__953_.gnd
rlabel metal1 1384 5042 1496 5058 0 _953_.gnd
rlabel metal1 1384 5282 1496 5298 0 _953_.vdd
rlabel metal2 1473 5133 1487 5147 0 _953_.A
rlabel metal2 1453 5153 1467 5167 0 _953_.B
rlabel metal2 1413 5153 1427 5167 0 _953_.C
rlabel metal2 1433 5133 1447 5147 0 _953_.Y
rlabel nsubstratencontact 1524 5288 1524 5288 0 FILL_1__1368_.vdd
rlabel metal1 1504 5042 1536 5058 0 FILL_1__1368_.gnd
rlabel nsubstratencontact 1504 5288 1504 5288 0 FILL_0__1368_.vdd
rlabel metal1 1484 5042 1516 5058 0 FILL_0__1368_.gnd
rlabel nsubstratencontact 1624 5288 1624 5288 0 FILL_1__1412_.vdd
rlabel metal1 1604 5042 1636 5058 0 FILL_1__1412_.gnd
rlabel nsubstratencontact 1604 5288 1604 5288 0 FILL_0__1412_.vdd
rlabel metal1 1584 5042 1616 5058 0 FILL_0__1412_.gnd
rlabel metal1 1624 5042 1736 5058 0 _1412_.gnd
rlabel metal1 1624 5282 1736 5298 0 _1412_.vdd
rlabel metal2 1713 5133 1727 5147 0 _1412_.A
rlabel metal2 1693 5153 1707 5167 0 _1412_.B
rlabel metal2 1653 5153 1667 5167 0 _1412_.C
rlabel metal2 1673 5133 1687 5147 0 _1412_.Y
rlabel metal1 1524 5042 1596 5058 0 _1368_.gnd
rlabel metal1 1524 5282 1596 5298 0 _1368_.vdd
rlabel metal2 1573 5113 1587 5127 0 _1368_.A
rlabel metal2 1553 5153 1567 5167 0 _1368_.Y
rlabel nsubstratencontact 1784 5288 1784 5288 0 FILL_2__1435_.vdd
rlabel metal1 1764 5042 1796 5058 0 FILL_2__1435_.gnd
rlabel nsubstratencontact 1764 5288 1764 5288 0 FILL_1__1435_.vdd
rlabel metal1 1744 5042 1776 5058 0 FILL_1__1435_.gnd
rlabel nsubstratencontact 1744 5288 1744 5288 0 FILL_0__1435_.vdd
rlabel metal1 1724 5042 1756 5058 0 FILL_0__1435_.gnd
rlabel metal1 1784 5282 1976 5298 0 _1435_.vdd
rlabel metal2 1933 5133 1947 5147 0 _1435_.A
rlabel metal2 1893 5153 1907 5167 0 _1435_.B
rlabel metal2 1873 5133 1887 5147 0 _1435_.C
rlabel metal2 1833 5153 1847 5167 0 _1435_.Y
rlabel metal1 1784 5042 1976 5058 0 _1435_.gnd
rlabel nsubstratencontact 2004 5288 2004 5288 0 FILL_1__1406_.vdd
rlabel metal1 1984 5042 2016 5058 0 FILL_1__1406_.gnd
rlabel nsubstratencontact 1984 5288 1984 5288 0 FILL_0__1406_.vdd
rlabel metal1 1964 5042 1996 5058 0 FILL_0__1406_.gnd
rlabel metal1 2004 5042 2136 5058 0 _1406_.gnd
rlabel metal1 2004 5282 2136 5298 0 _1406_.vdd
rlabel metal2 2113 5133 2127 5147 0 _1406_.A
rlabel metal2 2093 5153 2107 5167 0 _1406_.B
rlabel metal2 2033 5133 2047 5147 0 _1406_.C
rlabel metal2 2053 5153 2067 5167 0 _1406_.D
rlabel metal2 2073 5133 2087 5147 0 _1406_.Y
rlabel nsubstratencontact 2156 5288 2156 5288 0 FILL_1__1384_.vdd
rlabel metal1 2144 5042 2176 5058 0 FILL_1__1384_.gnd
rlabel nsubstratencontact 2136 5288 2136 5288 0 FILL_0__1384_.vdd
rlabel metal1 2124 5042 2156 5058 0 FILL_0__1384_.gnd
rlabel nsubstratencontact 2284 5288 2284 5288 0 FILL_1__1398_.vdd
rlabel metal1 2264 5042 2296 5058 0 FILL_1__1398_.gnd
rlabel nsubstratencontact 2264 5288 2264 5288 0 FILL_0__1398_.vdd
rlabel metal1 2244 5042 2276 5058 0 FILL_0__1398_.gnd
rlabel metal1 2164 5042 2256 5058 0 _1384_.gnd
rlabel metal1 2164 5282 2256 5298 0 _1384_.vdd
rlabel metal2 2173 5173 2187 5187 0 _1384_.A
rlabel metal2 2213 5173 2227 5187 0 _1384_.B
rlabel metal2 2193 5153 2207 5167 0 _1384_.Y
rlabel nsubstratencontact 2404 5288 2404 5288 0 FILL_0__1397_.vdd
rlabel metal1 2384 5042 2416 5058 0 FILL_0__1397_.gnd
rlabel metal1 2284 5042 2396 5058 0 _1398_.gnd
rlabel metal1 2284 5282 2396 5298 0 _1398_.vdd
rlabel metal2 2373 5153 2387 5167 0 _1398_.A
rlabel metal2 2353 5173 2367 5187 0 _1398_.B
rlabel metal2 2333 5153 2347 5167 0 _1398_.C
rlabel metal2 2313 5173 2327 5187 0 _1398_.Y
rlabel nsubstratencontact 2424 5288 2424 5288 0 FILL_1__1397_.vdd
rlabel metal1 2404 5042 2436 5058 0 FILL_1__1397_.gnd
rlabel metal1 2424 5042 2536 5058 0 _1397_.gnd
rlabel metal1 2424 5282 2536 5298 0 _1397_.vdd
rlabel metal2 2513 5153 2527 5167 0 _1397_.A
rlabel metal2 2493 5113 2507 5127 0 _1397_.B
rlabel metal2 2473 5153 2487 5167 0 _1397_.C
rlabel metal2 2453 5133 2467 5147 0 _1397_.Y
rlabel nsubstratencontact 2544 5288 2544 5288 0 FILL_0__1438_.vdd
rlabel metal1 2524 5042 2556 5058 0 FILL_0__1438_.gnd
rlabel nsubstratencontact 2564 5288 2564 5288 0 FILL_1__1438_.vdd
rlabel metal1 2544 5042 2576 5058 0 FILL_1__1438_.gnd
rlabel nsubstratencontact 2664 5288 2664 5288 0 FILL_1__1437_.vdd
rlabel metal1 2644 5042 2676 5058 0 FILL_1__1437_.gnd
rlabel nsubstratencontact 2644 5288 2644 5288 0 FILL_0__1437_.vdd
rlabel metal1 2624 5042 2656 5058 0 FILL_0__1437_.gnd
rlabel metal1 2564 5042 2636 5058 0 _1438_.gnd
rlabel metal1 2564 5282 2636 5298 0 _1438_.vdd
rlabel metal2 2613 5113 2627 5127 0 _1438_.A
rlabel metal2 2593 5153 2607 5167 0 _1438_.Y
rlabel nsubstratencontact 2784 5288 2784 5288 0 FILL_0__1383_.vdd
rlabel metal1 2764 5042 2796 5058 0 FILL_0__1383_.gnd
rlabel metal1 2664 5042 2776 5058 0 _1437_.gnd
rlabel metal1 2664 5282 2776 5298 0 _1437_.vdd
rlabel metal2 2753 5133 2767 5147 0 _1437_.A
rlabel metal2 2733 5153 2747 5167 0 _1437_.B
rlabel metal2 2693 5153 2707 5167 0 _1437_.C
rlabel metal2 2713 5133 2727 5147 0 _1437_.Y
rlabel nsubstratencontact 2824 5288 2824 5288 0 FILL_2__1383_.vdd
rlabel metal1 2804 5042 2836 5058 0 FILL_2__1383_.gnd
rlabel nsubstratencontact 2804 5288 2804 5288 0 FILL_1__1383_.vdd
rlabel metal1 2784 5042 2816 5058 0 FILL_1__1383_.gnd
rlabel metal1 2824 5042 2936 5058 0 _1383_.gnd
rlabel metal1 2824 5282 2936 5298 0 _1383_.vdd
rlabel metal2 2913 5133 2927 5147 0 _1383_.A
rlabel metal2 2893 5153 2907 5167 0 _1383_.B
rlabel metal2 2853 5153 2867 5167 0 _1383_.C
rlabel metal2 2873 5133 2887 5147 0 _1383_.Y
rlabel nsubstratencontact 2964 5288 2964 5288 0 FILL_1__1382_.vdd
rlabel metal1 2944 5042 2976 5058 0 FILL_1__1382_.gnd
rlabel nsubstratencontact 2944 5288 2944 5288 0 FILL_0__1382_.vdd
rlabel metal1 2924 5042 2956 5058 0 FILL_0__1382_.gnd
rlabel metal1 2964 5042 3076 5058 0 _1382_.gnd
rlabel metal1 2964 5282 3076 5298 0 _1382_.vdd
rlabel metal2 3053 5133 3067 5147 0 _1382_.A
rlabel metal2 2993 5133 3007 5147 0 _1382_.Y
rlabel metal2 3013 5173 3027 5187 0 _1382_.B
rlabel nsubstratencontact 3096 5288 3096 5288 0 FILL_1__1381_.vdd
rlabel metal1 3084 5042 3116 5058 0 FILL_1__1381_.gnd
rlabel nsubstratencontact 3076 5288 3076 5288 0 FILL_0__1381_.vdd
rlabel metal1 3064 5042 3096 5058 0 FILL_0__1381_.gnd
rlabel metal1 3104 5042 3196 5058 0 _1381_.gnd
rlabel metal1 3104 5282 3196 5298 0 _1381_.vdd
rlabel metal2 3153 5133 3167 5147 0 _1381_.B
rlabel metal2 3113 5133 3127 5147 0 _1381_.A
rlabel metal2 3133 5113 3147 5127 0 _1381_.Y
rlabel nsubstratencontact 3244 5288 3244 5288 0 FILL_2__1376_.vdd
rlabel metal1 3224 5042 3256 5058 0 FILL_2__1376_.gnd
rlabel nsubstratencontact 3224 5288 3224 5288 0 FILL_1__1376_.vdd
rlabel metal1 3204 5042 3236 5058 0 FILL_1__1376_.gnd
rlabel nsubstratencontact 3204 5288 3204 5288 0 FILL_0__1376_.vdd
rlabel metal1 3184 5042 3216 5058 0 FILL_0__1376_.gnd
rlabel metal1 3244 5042 3316 5058 0 _1376_.gnd
rlabel metal1 3244 5282 3316 5298 0 _1376_.vdd
rlabel metal2 3293 5113 3307 5127 0 _1376_.A
rlabel metal2 3273 5153 3287 5167 0 _1376_.Y
rlabel nsubstratencontact 3344 5288 3344 5288 0 FILL_1__1372_.vdd
rlabel metal1 3324 5042 3356 5058 0 FILL_1__1372_.gnd
rlabel nsubstratencontact 3324 5288 3324 5288 0 FILL_0__1372_.vdd
rlabel metal1 3304 5042 3336 5058 0 FILL_0__1372_.gnd
rlabel metal1 3344 5042 3436 5058 0 _1372_.gnd
rlabel metal1 3344 5282 3436 5298 0 _1372_.vdd
rlabel metal2 3373 5133 3387 5147 0 _1372_.B
rlabel metal2 3413 5133 3427 5147 0 _1372_.A
rlabel metal2 3393 5113 3407 5127 0 _1372_.Y
rlabel nsubstratencontact 3484 5288 3484 5288 0 FILL_2__1311_.vdd
rlabel metal1 3464 5042 3496 5058 0 FILL_2__1311_.gnd
rlabel nsubstratencontact 3464 5288 3464 5288 0 FILL_1__1311_.vdd
rlabel metal1 3444 5042 3476 5058 0 FILL_1__1311_.gnd
rlabel nsubstratencontact 3444 5288 3444 5288 0 FILL_0__1311_.vdd
rlabel metal1 3424 5042 3456 5058 0 FILL_0__1311_.gnd
rlabel metal1 3484 5042 3596 5058 0 _1311_.gnd
rlabel metal1 3484 5282 3596 5298 0 _1311_.vdd
rlabel metal2 3573 5133 3587 5147 0 _1311_.A
rlabel metal2 3553 5153 3567 5167 0 _1311_.B
rlabel metal2 3513 5153 3527 5167 0 _1311_.C
rlabel metal2 3533 5133 3547 5147 0 _1311_.Y
rlabel nsubstratencontact 3616 5288 3616 5288 0 FILL_1__1375_.vdd
rlabel metal1 3604 5042 3636 5058 0 FILL_1__1375_.gnd
rlabel nsubstratencontact 3596 5288 3596 5288 0 FILL_0__1375_.vdd
rlabel metal1 3584 5042 3616 5058 0 FILL_0__1375_.gnd
rlabel metal1 3624 5042 3716 5058 0 _1375_.gnd
rlabel metal1 3624 5282 3716 5298 0 _1375_.vdd
rlabel metal2 3633 5173 3647 5187 0 _1375_.A
rlabel metal2 3673 5173 3687 5187 0 _1375_.B
rlabel metal2 3653 5153 3667 5167 0 _1375_.Y
rlabel nsubstratencontact 3744 5288 3744 5288 0 FILL_1__1440_.vdd
rlabel metal1 3724 5042 3756 5058 0 FILL_1__1440_.gnd
rlabel nsubstratencontact 3724 5288 3724 5288 0 FILL_0__1440_.vdd
rlabel metal1 3704 5042 3736 5058 0 FILL_0__1440_.gnd
rlabel metal1 3744 5042 3836 5058 0 _1440_.gnd
rlabel metal1 3744 5282 3836 5298 0 _1440_.vdd
rlabel metal2 3813 5173 3827 5187 0 _1440_.A
rlabel metal2 3773 5173 3787 5187 0 _1440_.B
rlabel metal2 3793 5153 3807 5167 0 _1440_.Y
rlabel nsubstratencontact 3884 5288 3884 5288 0 FILL_2__1396_.vdd
rlabel metal1 3864 5042 3896 5058 0 FILL_2__1396_.gnd
rlabel nsubstratencontact 3864 5288 3864 5288 0 FILL_1__1396_.vdd
rlabel metal1 3844 5042 3876 5058 0 FILL_1__1396_.gnd
rlabel nsubstratencontact 3844 5288 3844 5288 0 FILL_0__1396_.vdd
rlabel metal1 3824 5042 3856 5058 0 FILL_0__1396_.gnd
rlabel metal1 3884 5042 3976 5058 0 _1396_.gnd
rlabel metal1 3884 5282 3976 5298 0 _1396_.vdd
rlabel metal2 3953 5173 3967 5187 0 _1396_.A
rlabel metal2 3913 5173 3927 5187 0 _1396_.B
rlabel metal2 3933 5153 3947 5167 0 _1396_.Y
rlabel nsubstratencontact 3996 5288 3996 5288 0 FILL_1__1443_.vdd
rlabel metal1 3984 5042 4016 5058 0 FILL_1__1443_.gnd
rlabel nsubstratencontact 3976 5288 3976 5288 0 FILL_0__1443_.vdd
rlabel metal1 3964 5042 3996 5058 0 FILL_0__1443_.gnd
rlabel metal1 4004 5042 4116 5058 0 _1443_.gnd
rlabel metal1 4004 5282 4116 5298 0 _1443_.vdd
rlabel metal2 4013 5153 4027 5167 0 _1443_.A
rlabel metal2 4033 5173 4047 5187 0 _1443_.B
rlabel metal2 4053 5153 4067 5167 0 _1443_.C
rlabel metal2 4073 5173 4087 5187 0 _1443_.Y
rlabel nsubstratencontact 4144 5288 4144 5288 0 FILL_1__1395_.vdd
rlabel metal1 4124 5042 4156 5058 0 FILL_1__1395_.gnd
rlabel nsubstratencontact 4124 5288 4124 5288 0 FILL_0__1395_.vdd
rlabel metal1 4104 5042 4136 5058 0 FILL_0__1395_.gnd
rlabel metal1 4144 5042 4256 5058 0 _1395_.gnd
rlabel metal1 4144 5282 4256 5298 0 _1395_.vdd
rlabel metal2 4233 5133 4247 5147 0 _1395_.A
rlabel metal2 4213 5153 4227 5167 0 _1395_.B
rlabel metal2 4173 5153 4187 5167 0 _1395_.C
rlabel metal2 4193 5133 4207 5147 0 _1395_.Y
rlabel nsubstratencontact 4296 5288 4296 5288 0 FILL_2__1442_.vdd
rlabel metal1 4284 5042 4316 5058 0 FILL_2__1442_.gnd
rlabel nsubstratencontact 4276 5288 4276 5288 0 FILL_1__1442_.vdd
rlabel metal1 4264 5042 4296 5058 0 FILL_1__1442_.gnd
rlabel nsubstratencontact 4256 5288 4256 5288 0 FILL_0__1442_.vdd
rlabel metal1 4244 5042 4276 5058 0 FILL_0__1442_.gnd
rlabel nsubstratencontact 4416 5288 4416 5288 0 FILL_0__1386_.vdd
rlabel metal1 4404 5042 4436 5058 0 FILL_0__1386_.gnd
rlabel metal1 4304 5042 4416 5058 0 _1442_.gnd
rlabel metal1 4304 5282 4416 5298 0 _1442_.vdd
rlabel metal2 4313 5133 4327 5147 0 _1442_.A
rlabel metal2 4333 5153 4347 5167 0 _1442_.B
rlabel metal2 4373 5153 4387 5167 0 _1442_.C
rlabel metal2 4353 5133 4367 5147 0 _1442_.Y
rlabel nsubstratencontact 4544 5288 4544 5288 0 FILL_1__1392_.vdd
rlabel metal1 4524 5042 4556 5058 0 FILL_1__1392_.gnd
rlabel nsubstratencontact 4436 5288 4436 5288 0 FILL_1__1386_.vdd
rlabel metal1 4424 5042 4456 5058 0 FILL_1__1386_.gnd
rlabel nsubstratencontact 4524 5288 4524 5288 0 FILL_0__1392_.vdd
rlabel metal1 4504 5042 4536 5058 0 FILL_0__1392_.gnd
rlabel metal1 4444 5042 4516 5058 0 _1386_.gnd
rlabel metal1 4444 5282 4516 5298 0 _1386_.vdd
rlabel metal2 4453 5113 4467 5127 0 _1386_.A
rlabel metal2 4473 5153 4487 5167 0 _1386_.Y
rlabel metal1 4544 5042 4656 5058 0 _1392_.gnd
rlabel metal1 4544 5282 4656 5298 0 _1392_.vdd
rlabel metal2 4633 5153 4647 5167 0 _1392_.A
rlabel metal2 4613 5173 4627 5187 0 _1392_.B
rlabel metal2 4593 5153 4607 5167 0 _1392_.C
rlabel metal2 4573 5173 4587 5187 0 _1392_.Y
rlabel metal1 4824 5042 4916 5058 0 _1042_.gnd
rlabel metal1 4824 5282 4916 5298 0 _1042_.vdd
rlabel metal2 4873 5133 4887 5147 0 _1042_.B
rlabel metal2 4833 5133 4847 5147 0 _1042_.A
rlabel metal2 4853 5113 4867 5127 0 _1042_.Y
rlabel metal1 4684 5042 4796 5058 0 _1444_.gnd
rlabel metal1 4684 5282 4796 5298 0 _1444_.vdd
rlabel metal2 4693 5153 4707 5167 0 _1444_.A
rlabel metal2 4713 5113 4727 5127 0 _1444_.B
rlabel metal2 4733 5153 4747 5167 0 _1444_.C
rlabel metal2 4753 5133 4767 5147 0 _1444_.Y
rlabel metal1 4904 5042 5156 5058 0 _1660_.gnd
rlabel metal1 4904 5282 5156 5298 0 _1660_.vdd
rlabel metal2 5053 5133 5067 5147 0 _1660_.D
rlabel metal2 5013 5133 5027 5147 0 _1660_.CLK
rlabel metal2 4933 5133 4947 5147 0 _1660_.Q
rlabel nsubstratencontact 4796 5288 4796 5288 0 FILL_0__1042_.vdd
rlabel metal1 4784 5042 4816 5058 0 FILL_0__1042_.gnd
rlabel nsubstratencontact 4656 5288 4656 5288 0 FILL_0__1444_.vdd
rlabel metal1 4644 5042 4676 5058 0 FILL_0__1444_.gnd
rlabel nsubstratencontact 4816 5288 4816 5288 0 FILL_1__1042_.vdd
rlabel metal1 4804 5042 4836 5058 0 FILL_1__1042_.gnd
rlabel nsubstratencontact 4676 5288 4676 5288 0 FILL_1__1444_.vdd
rlabel metal1 4664 5042 4696 5058 0 FILL_1__1444_.gnd
rlabel nsubstratencontact 5176 5288 5176 5288 0 FILL_1__1619_.vdd
rlabel metal1 5164 5042 5196 5058 0 FILL_1__1619_.gnd
rlabel nsubstratencontact 5156 5288 5156 5288 0 FILL_0__1619_.vdd
rlabel metal1 5144 5042 5176 5058 0 FILL_0__1619_.gnd
rlabel nsubstratencontact 5296 5288 5296 5288 0 FILL_0__1041_.vdd
rlabel metal1 5284 5042 5316 5058 0 FILL_0__1041_.gnd
rlabel metal1 5184 5042 5296 5058 0 _1619_.gnd
rlabel metal1 5184 5282 5296 5298 0 _1619_.vdd
rlabel metal2 5193 5133 5207 5147 0 _1619_.A
rlabel metal2 5213 5153 5227 5167 0 _1619_.B
rlabel metal2 5253 5153 5267 5167 0 _1619_.C
rlabel metal2 5233 5133 5247 5147 0 _1619_.Y
rlabel nsubstratencontact 5416 5288 5416 5288 0 FILL_1__1650_.vdd
rlabel metal1 5404 5042 5436 5058 0 FILL_1__1650_.gnd
rlabel nsubstratencontact 5316 5288 5316 5288 0 FILL_1__1041_.vdd
rlabel metal1 5304 5042 5336 5058 0 FILL_1__1041_.gnd
rlabel nsubstratencontact 5396 5288 5396 5288 0 FILL_0__1650_.vdd
rlabel metal1 5384 5042 5416 5058 0 FILL_0__1650_.gnd
rlabel metal1 5424 5042 5536 5058 0 _1650_.gnd
rlabel metal1 5424 5282 5536 5298 0 _1650_.vdd
rlabel metal2 5433 5133 5447 5147 0 _1650_.A
rlabel metal2 5453 5153 5467 5167 0 _1650_.B
rlabel metal2 5493 5153 5507 5167 0 _1650_.C
rlabel metal2 5473 5133 5487 5147 0 _1650_.Y
rlabel metal1 5324 5042 5396 5058 0 _1041_.gnd
rlabel metal1 5324 5282 5396 5298 0 _1041_.vdd
rlabel metal2 5333 5113 5347 5127 0 _1041_.A
rlabel metal2 5353 5153 5367 5167 0 _1041_.Y
rlabel nsubstratencontact 5564 5288 5564 5288 0 FILL_1__1613_.vdd
rlabel metal1 5544 5042 5576 5058 0 FILL_1__1613_.gnd
rlabel nsubstratencontact 5544 5288 5544 5288 0 FILL_0__1613_.vdd
rlabel metal1 5524 5042 5556 5058 0 FILL_0__1613_.gnd
rlabel metal1 5564 5042 5656 5058 0 _1613_.gnd
rlabel metal1 5564 5282 5656 5298 0 _1613_.vdd
rlabel metal2 5633 5173 5647 5187 0 _1613_.A
rlabel metal2 5593 5173 5607 5187 0 _1613_.B
rlabel metal2 5613 5153 5627 5167 0 _1613_.Y
rlabel metal1 5684 5042 5776 5058 0 _1649_.gnd
rlabel metal1 5684 5282 5776 5298 0 _1649_.vdd
rlabel metal2 5693 5173 5707 5187 0 _1649_.A
rlabel metal2 5733 5173 5747 5187 0 _1649_.B
rlabel metal2 5713 5153 5727 5167 0 _1649_.Y
rlabel nsubstratencontact 5776 5288 5776 5288 0 FILL86550x75750.vdd
rlabel metal1 5764 5042 5796 5058 0 FILL86550x75750.gnd
rlabel nsubstratencontact 5796 5288 5796 5288 0 FILL86850x75750.vdd
rlabel metal1 5784 5042 5816 5058 0 FILL86850x75750.gnd
rlabel nsubstratencontact 5656 5288 5656 5288 0 FILL_0__1649_.vdd
rlabel metal1 5644 5042 5676 5058 0 FILL_0__1649_.gnd
rlabel nsubstratencontact 5676 5288 5676 5288 0 FILL_1__1649_.vdd
rlabel metal1 5664 5042 5696 5058 0 FILL_1__1649_.gnd
rlabel nsubstratencontact 44 5292 44 5292 0 FILL_1__997_.vdd
rlabel metal1 24 5522 56 5538 0 FILL_1__997_.gnd
rlabel nsubstratencontact 24 5292 24 5292 0 FILL_0__997_.vdd
rlabel metal1 4 5522 36 5538 0 FILL_0__997_.gnd
rlabel metal1 44 5522 156 5538 0 _997_.gnd
rlabel metal1 44 5282 156 5298 0 _997_.vdd
rlabel metal2 133 5433 147 5447 0 _997_.A
rlabel metal2 113 5413 127 5427 0 _997_.B
rlabel metal2 73 5413 87 5427 0 _997_.C
rlabel metal2 93 5433 107 5447 0 _997_.Y
rlabel nsubstratencontact 204 5292 204 5292 0 FILL_2__1187_.vdd
rlabel metal1 184 5522 216 5538 0 FILL_2__1187_.gnd
rlabel nsubstratencontact 184 5292 184 5292 0 FILL_1__1187_.vdd
rlabel metal1 164 5522 196 5538 0 FILL_1__1187_.gnd
rlabel nsubstratencontact 164 5292 164 5292 0 FILL_0__1187_.vdd
rlabel metal1 144 5522 176 5538 0 FILL_0__1187_.gnd
rlabel metal1 204 5522 316 5538 0 _1187_.gnd
rlabel metal1 204 5282 316 5298 0 _1187_.vdd
rlabel metal2 293 5413 307 5427 0 _1187_.A
rlabel metal2 273 5393 287 5407 0 _1187_.B
rlabel metal2 253 5413 267 5427 0 _1187_.C
rlabel metal2 233 5393 247 5407 0 _1187_.Y
rlabel nsubstratencontact 344 5292 344 5292 0 FILL_1__1163_.vdd
rlabel metal1 324 5522 356 5538 0 FILL_1__1163_.gnd
rlabel nsubstratencontact 324 5292 324 5292 0 FILL_0__1163_.vdd
rlabel metal1 304 5522 336 5538 0 FILL_0__1163_.gnd
rlabel metal1 344 5522 456 5538 0 _1163_.gnd
rlabel metal1 344 5282 456 5298 0 _1163_.vdd
rlabel metal2 433 5413 447 5427 0 _1163_.A
rlabel metal2 413 5393 427 5407 0 _1163_.B
rlabel metal2 393 5413 407 5427 0 _1163_.C
rlabel metal2 373 5393 387 5407 0 _1163_.Y
rlabel nsubstratencontact 484 5292 484 5292 0 FILL_1__1186_.vdd
rlabel metal1 464 5522 496 5538 0 FILL_1__1186_.gnd
rlabel nsubstratencontact 464 5292 464 5292 0 FILL_0__1186_.vdd
rlabel metal1 444 5522 476 5538 0 FILL_0__1186_.gnd
rlabel metal1 484 5522 596 5538 0 _1186_.gnd
rlabel metal1 484 5282 596 5298 0 _1186_.vdd
rlabel metal2 573 5413 587 5427 0 _1186_.A
rlabel metal2 553 5393 567 5407 0 _1186_.B
rlabel metal2 533 5413 547 5427 0 _1186_.C
rlabel metal2 513 5393 527 5407 0 _1186_.Y
rlabel nsubstratencontact 636 5292 636 5292 0 FILL_2__1141_.vdd
rlabel metal1 624 5522 656 5538 0 FILL_2__1141_.gnd
rlabel nsubstratencontact 616 5292 616 5292 0 FILL_1__1141_.vdd
rlabel metal1 604 5522 636 5538 0 FILL_1__1141_.gnd
rlabel nsubstratencontact 596 5292 596 5292 0 FILL_0__1141_.vdd
rlabel metal1 584 5522 616 5538 0 FILL_0__1141_.gnd
rlabel nsubstratencontact 756 5292 756 5292 0 FILL_0__956_.vdd
rlabel metal1 744 5522 776 5538 0 FILL_0__956_.gnd
rlabel metal1 644 5522 756 5538 0 _1141_.gnd
rlabel metal1 644 5282 756 5298 0 _1141_.vdd
rlabel metal2 653 5413 667 5427 0 _1141_.A
rlabel metal2 673 5393 687 5407 0 _1141_.B
rlabel metal2 693 5413 707 5427 0 _1141_.C
rlabel metal2 713 5393 727 5407 0 _1141_.Y
rlabel nsubstratencontact 776 5292 776 5292 0 FILL_1__956_.vdd
rlabel metal1 764 5522 796 5538 0 FILL_1__956_.gnd
rlabel metal1 784 5522 896 5538 0 _956_.gnd
rlabel metal1 784 5282 896 5298 0 _956_.vdd
rlabel metal2 793 5433 807 5447 0 _956_.A
rlabel metal2 813 5413 827 5427 0 _956_.B
rlabel metal2 853 5413 867 5427 0 _956_.C
rlabel metal2 833 5433 847 5447 0 _956_.Y
rlabel nsubstratencontact 916 5292 916 5292 0 FILL_1__1142_.vdd
rlabel metal1 904 5522 936 5538 0 FILL_1__1142_.gnd
rlabel nsubstratencontact 896 5292 896 5292 0 FILL_0__1142_.vdd
rlabel metal1 884 5522 916 5538 0 FILL_0__1142_.gnd
rlabel metal1 924 5522 1036 5538 0 _1142_.gnd
rlabel metal1 924 5282 1036 5298 0 _1142_.vdd
rlabel metal2 933 5413 947 5427 0 _1142_.A
rlabel metal2 953 5393 967 5407 0 _1142_.B
rlabel metal2 973 5413 987 5427 0 _1142_.C
rlabel metal2 993 5393 1007 5407 0 _1142_.Y
rlabel nsubstratencontact 1064 5292 1064 5292 0 FILL_1__1133_.vdd
rlabel metal1 1044 5522 1076 5538 0 FILL_1__1133_.gnd
rlabel nsubstratencontact 1044 5292 1044 5292 0 FILL_0__1133_.vdd
rlabel metal1 1024 5522 1056 5538 0 FILL_0__1133_.gnd
rlabel metal1 1064 5522 1176 5538 0 _1133_.gnd
rlabel metal1 1064 5282 1176 5298 0 _1133_.vdd
rlabel metal2 1153 5413 1167 5427 0 _1133_.A
rlabel metal2 1133 5453 1147 5467 0 _1133_.B
rlabel metal2 1113 5413 1127 5427 0 _1133_.C
rlabel metal2 1093 5433 1107 5447 0 _1133_.Y
rlabel nsubstratencontact 1196 5292 1196 5292 0 FILL_1__1136_.vdd
rlabel metal1 1184 5522 1216 5538 0 FILL_1__1136_.gnd
rlabel nsubstratencontact 1176 5292 1176 5292 0 FILL_0__1136_.vdd
rlabel metal1 1164 5522 1196 5538 0 FILL_0__1136_.gnd
rlabel metal1 1204 5522 1316 5538 0 _1136_.gnd
rlabel metal1 1204 5282 1316 5298 0 _1136_.vdd
rlabel metal2 1213 5413 1227 5427 0 _1136_.A
rlabel metal2 1233 5393 1247 5407 0 _1136_.B
rlabel metal2 1253 5413 1267 5427 0 _1136_.C
rlabel metal2 1273 5393 1287 5407 0 _1136_.Y
rlabel nsubstratencontact 1356 5292 1356 5292 0 FILL_2__1128_.vdd
rlabel metal1 1344 5522 1376 5538 0 FILL_2__1128_.gnd
rlabel nsubstratencontact 1336 5292 1336 5292 0 FILL_1__1128_.vdd
rlabel metal1 1324 5522 1356 5538 0 FILL_1__1128_.gnd
rlabel nsubstratencontact 1316 5292 1316 5292 0 FILL_0__1128_.vdd
rlabel metal1 1304 5522 1336 5538 0 FILL_0__1128_.gnd
rlabel metal1 1364 5522 1456 5538 0 _1128_.gnd
rlabel metal1 1364 5282 1456 5298 0 _1128_.vdd
rlabel metal2 1413 5433 1427 5447 0 _1128_.B
rlabel metal2 1373 5433 1387 5447 0 _1128_.A
rlabel metal2 1393 5453 1407 5467 0 _1128_.Y
rlabel nsubstratencontact 1484 5292 1484 5292 0 FILL_1__1413_.vdd
rlabel metal1 1464 5522 1496 5538 0 FILL_1__1413_.gnd
rlabel nsubstratencontact 1464 5292 1464 5292 0 FILL_0__1413_.vdd
rlabel metal1 1444 5522 1476 5538 0 FILL_0__1413_.gnd
rlabel metal1 1484 5522 1596 5538 0 _1413_.gnd
rlabel metal1 1484 5282 1596 5298 0 _1413_.vdd
rlabel metal2 1573 5413 1587 5427 0 _1413_.A
rlabel metal2 1553 5393 1567 5407 0 _1413_.B
rlabel metal2 1533 5413 1547 5427 0 _1413_.C
rlabel metal2 1513 5393 1527 5407 0 _1413_.Y
rlabel nsubstratencontact 1616 5292 1616 5292 0 FILL_1__1469_.vdd
rlabel metal1 1604 5522 1636 5538 0 FILL_1__1469_.gnd
rlabel nsubstratencontact 1596 5292 1596 5292 0 FILL_0__1469_.vdd
rlabel metal1 1584 5522 1616 5538 0 FILL_0__1469_.gnd
rlabel metal1 1624 5522 1736 5538 0 _1469_.gnd
rlabel metal1 1624 5282 1736 5298 0 _1469_.vdd
rlabel metal2 1633 5433 1647 5447 0 _1469_.A
rlabel metal2 1653 5413 1667 5427 0 _1469_.B
rlabel metal2 1693 5413 1707 5427 0 _1469_.C
rlabel metal2 1673 5433 1687 5447 0 _1469_.Y
rlabel nsubstratencontact 1764 5292 1764 5292 0 FILL_1__1404_.vdd
rlabel metal1 1744 5522 1776 5538 0 FILL_1__1404_.gnd
rlabel nsubstratencontact 1744 5292 1744 5292 0 FILL_0__1404_.vdd
rlabel metal1 1724 5522 1756 5538 0 FILL_0__1404_.gnd
rlabel metal1 1764 5522 1876 5538 0 _1404_.gnd
rlabel metal1 1764 5282 1876 5298 0 _1404_.vdd
rlabel metal2 1853 5413 1867 5427 0 _1404_.A
rlabel metal2 1833 5393 1847 5407 0 _1404_.B
rlabel metal2 1813 5413 1827 5427 0 _1404_.C
rlabel metal2 1793 5393 1807 5407 0 _1404_.Y
rlabel nsubstratencontact 1904 5292 1904 5292 0 FILL_1__1470_.vdd
rlabel metal1 1884 5522 1916 5538 0 FILL_1__1470_.gnd
rlabel nsubstratencontact 1884 5292 1884 5292 0 FILL_0__1470_.vdd
rlabel metal1 1864 5522 1896 5538 0 FILL_0__1470_.gnd
rlabel nsubstratencontact 2016 5292 2016 5292 0 FILL_0__1466_.vdd
rlabel metal1 2004 5522 2036 5538 0 FILL_0__1466_.gnd
rlabel metal1 1904 5522 2016 5538 0 _1470_.gnd
rlabel metal1 1904 5282 2016 5298 0 _1470_.vdd
rlabel metal2 1993 5413 2007 5427 0 _1470_.A
rlabel metal2 1973 5393 1987 5407 0 _1470_.B
rlabel metal2 1953 5413 1967 5427 0 _1470_.C
rlabel metal2 1933 5393 1947 5407 0 _1470_.Y
rlabel nsubstratencontact 2036 5292 2036 5292 0 FILL_1__1466_.vdd
rlabel metal1 2024 5522 2056 5538 0 FILL_1__1466_.gnd
rlabel nsubstratencontact 2164 5292 2164 5292 0 FILL_1__1402_.vdd
rlabel metal1 2144 5522 2176 5538 0 FILL_1__1402_.gnd
rlabel nsubstratencontact 2144 5292 2144 5292 0 FILL_0__1402_.vdd
rlabel metal1 2124 5522 2156 5538 0 FILL_0__1402_.gnd
rlabel metal1 2044 5522 2136 5538 0 _1466_.gnd
rlabel metal1 2044 5282 2136 5298 0 _1466_.vdd
rlabel metal2 2053 5393 2067 5407 0 _1466_.A
rlabel metal2 2093 5393 2107 5407 0 _1466_.B
rlabel metal2 2073 5413 2087 5427 0 _1466_.Y
rlabel nsubstratencontact 2184 5292 2184 5292 0 FILL_2__1402_.vdd
rlabel metal1 2164 5522 2196 5538 0 FILL_2__1402_.gnd
rlabel nsubstratencontact 2284 5292 2284 5292 0 FILL_1__1401_.vdd
rlabel metal1 2264 5522 2296 5538 0 FILL_1__1401_.gnd
rlabel nsubstratencontact 2264 5292 2264 5292 0 FILL_0__1401_.vdd
rlabel metal1 2244 5522 2276 5538 0 FILL_0__1401_.gnd
rlabel metal1 2184 5522 2256 5538 0 _1402_.gnd
rlabel metal1 2184 5282 2256 5298 0 _1402_.vdd
rlabel metal2 2233 5453 2247 5467 0 _1402_.A
rlabel metal2 2213 5413 2227 5427 0 _1402_.Y
rlabel nsubstratencontact 2396 5292 2396 5292 0 FILL_0__1460_.vdd
rlabel metal1 2384 5522 2416 5538 0 FILL_0__1460_.gnd
rlabel metal1 2284 5522 2396 5538 0 _1401_.gnd
rlabel metal1 2284 5282 2396 5298 0 _1401_.vdd
rlabel metal2 2373 5433 2387 5447 0 _1401_.A
rlabel metal2 2313 5433 2327 5447 0 _1401_.Y
rlabel metal2 2333 5393 2347 5407 0 _1401_.B
rlabel nsubstratencontact 2416 5292 2416 5292 0 FILL_1__1460_.vdd
rlabel metal1 2404 5522 2436 5538 0 FILL_1__1460_.gnd
rlabel metal1 2424 5522 2536 5538 0 _1460_.gnd
rlabel metal1 2424 5282 2536 5298 0 _1460_.vdd
rlabel metal2 2433 5433 2447 5447 0 _1460_.A
rlabel metal2 2453 5413 2467 5427 0 _1460_.B
rlabel metal2 2493 5413 2507 5427 0 _1460_.C
rlabel metal2 2473 5433 2487 5447 0 _1460_.Y
rlabel nsubstratencontact 2544 5292 2544 5292 0 FILL_0__1461_.vdd
rlabel metal1 2524 5522 2556 5538 0 FILL_0__1461_.gnd
rlabel nsubstratencontact 2584 5292 2584 5292 0 FILL_2__1461_.vdd
rlabel metal1 2564 5522 2596 5538 0 FILL_2__1461_.gnd
rlabel nsubstratencontact 2564 5292 2564 5292 0 FILL_1__1461_.vdd
rlabel metal1 2544 5522 2576 5538 0 FILL_1__1461_.gnd
rlabel metal1 2584 5522 2696 5538 0 _1461_.gnd
rlabel metal1 2584 5282 2696 5298 0 _1461_.vdd
rlabel metal2 2673 5413 2687 5427 0 _1461_.A
rlabel metal2 2653 5393 2667 5407 0 _1461_.B
rlabel metal2 2633 5413 2647 5427 0 _1461_.C
rlabel metal2 2613 5393 2627 5407 0 _1461_.Y
rlabel nsubstratencontact 2724 5292 2724 5292 0 FILL_1__1458_.vdd
rlabel metal1 2704 5522 2736 5538 0 FILL_1__1458_.gnd
rlabel nsubstratencontact 2704 5292 2704 5292 0 FILL_0__1458_.vdd
rlabel metal1 2684 5522 2716 5538 0 FILL_0__1458_.gnd
rlabel metal1 2724 5522 2836 5538 0 _1458_.gnd
rlabel metal1 2724 5282 2836 5298 0 _1458_.vdd
rlabel metal2 2813 5413 2827 5427 0 _1458_.A
rlabel metal2 2793 5393 2807 5407 0 _1458_.B
rlabel metal2 2773 5413 2787 5427 0 _1458_.C
rlabel metal2 2753 5393 2767 5407 0 _1458_.Y
rlabel nsubstratencontact 2856 5292 2856 5292 0 FILL_1__1488_.vdd
rlabel metal1 2844 5522 2876 5538 0 FILL_1__1488_.gnd
rlabel nsubstratencontact 2836 5292 2836 5292 0 FILL_0__1488_.vdd
rlabel metal1 2824 5522 2856 5538 0 FILL_0__1488_.gnd
rlabel metal1 2864 5522 2976 5538 0 _1488_.gnd
rlabel metal1 2864 5282 2976 5298 0 _1488_.vdd
rlabel metal2 2873 5433 2887 5447 0 _1488_.A
rlabel metal2 2893 5413 2907 5427 0 _1488_.B
rlabel metal2 2933 5413 2947 5427 0 _1488_.C
rlabel metal2 2913 5433 2927 5447 0 _1488_.Y
rlabel nsubstratencontact 2996 5292 2996 5292 0 FILL_1__1489_.vdd
rlabel metal1 2984 5522 3016 5538 0 FILL_1__1489_.gnd
rlabel nsubstratencontact 2976 5292 2976 5292 0 FILL_0__1489_.vdd
rlabel metal1 2964 5522 2996 5538 0 FILL_0__1489_.gnd
rlabel metal1 3004 5522 3076 5538 0 _1489_.gnd
rlabel metal1 3004 5282 3076 5298 0 _1489_.vdd
rlabel metal2 3013 5453 3027 5467 0 _1489_.A
rlabel metal2 3033 5413 3047 5427 0 _1489_.Y
rlabel nsubstratencontact 3096 5292 3096 5292 0 FILL_1__1513_.vdd
rlabel metal1 3084 5522 3116 5538 0 FILL_1__1513_.gnd
rlabel nsubstratencontact 3076 5292 3076 5292 0 FILL_0__1513_.vdd
rlabel metal1 3064 5522 3096 5538 0 FILL_0__1513_.gnd
rlabel metal1 3104 5522 3196 5538 0 _1513_.gnd
rlabel metal1 3104 5282 3196 5298 0 _1513_.vdd
rlabel metal2 3113 5393 3127 5407 0 _1513_.A
rlabel metal2 3153 5393 3167 5407 0 _1513_.B
rlabel metal2 3133 5413 3147 5427 0 _1513_.Y
rlabel nsubstratencontact 3236 5292 3236 5292 0 FILL_2__1514_.vdd
rlabel metal1 3224 5522 3256 5538 0 FILL_2__1514_.gnd
rlabel nsubstratencontact 3216 5292 3216 5292 0 FILL_1__1514_.vdd
rlabel metal1 3204 5522 3236 5538 0 FILL_1__1514_.gnd
rlabel nsubstratencontact 3196 5292 3196 5292 0 FILL_0__1514_.vdd
rlabel metal1 3184 5522 3216 5538 0 FILL_0__1514_.gnd
rlabel metal1 3244 5522 3356 5538 0 _1514_.gnd
rlabel metal1 3244 5282 3356 5298 0 _1514_.vdd
rlabel metal2 3253 5413 3267 5427 0 _1514_.A
rlabel metal2 3273 5393 3287 5407 0 _1514_.B
rlabel metal2 3293 5413 3307 5427 0 _1514_.C
rlabel metal2 3313 5393 3327 5407 0 _1514_.Y
rlabel nsubstratencontact 3376 5292 3376 5292 0 FILL_1__1512_.vdd
rlabel metal1 3364 5522 3396 5538 0 FILL_1__1512_.gnd
rlabel nsubstratencontact 3356 5292 3356 5292 0 FILL_0__1512_.vdd
rlabel metal1 3344 5522 3376 5538 0 FILL_0__1512_.gnd
rlabel metal1 3384 5522 3476 5538 0 _1512_.gnd
rlabel metal1 3384 5282 3476 5298 0 _1512_.vdd
rlabel metal2 3393 5393 3407 5407 0 _1512_.A
rlabel metal2 3433 5393 3447 5407 0 _1512_.B
rlabel metal2 3413 5413 3427 5427 0 _1512_.Y
rlabel nsubstratencontact 3496 5292 3496 5292 0 FILL_1__1509_.vdd
rlabel metal1 3484 5522 3516 5538 0 FILL_1__1509_.gnd
rlabel nsubstratencontact 3476 5292 3476 5292 0 FILL_0__1509_.vdd
rlabel metal1 3464 5522 3496 5538 0 FILL_0__1509_.gnd
rlabel metal1 3504 5522 3616 5538 0 _1509_.gnd
rlabel metal1 3504 5282 3616 5298 0 _1509_.vdd
rlabel metal2 3513 5453 3527 5467 0 _1509_.A
rlabel metal2 3533 5433 3547 5447 0 _1509_.B
rlabel metal2 3573 5413 3587 5427 0 _1509_.Y
rlabel nsubstratencontact 3644 5292 3644 5292 0 FILL_1__1511_.vdd
rlabel metal1 3624 5522 3656 5538 0 FILL_1__1511_.gnd
rlabel nsubstratencontact 3624 5292 3624 5292 0 FILL_0__1511_.vdd
rlabel metal1 3604 5522 3636 5538 0 FILL_0__1511_.gnd
rlabel metal1 3644 5522 3756 5538 0 _1511_.gnd
rlabel metal1 3644 5282 3756 5298 0 _1511_.vdd
rlabel metal2 3733 5413 3747 5427 0 _1511_.A
rlabel metal2 3713 5393 3727 5407 0 _1511_.B
rlabel metal2 3693 5413 3707 5427 0 _1511_.C
rlabel metal2 3673 5393 3687 5407 0 _1511_.Y
rlabel nsubstratencontact 3784 5292 3784 5292 0 FILL_1__1543_.vdd
rlabel metal1 3764 5522 3796 5538 0 FILL_1__1543_.gnd
rlabel nsubstratencontact 3764 5292 3764 5292 0 FILL_0__1543_.vdd
rlabel metal1 3744 5522 3776 5538 0 FILL_0__1543_.gnd
rlabel metal1 3784 5522 3896 5538 0 _1543_.gnd
rlabel metal1 3784 5282 3896 5298 0 _1543_.vdd
rlabel metal2 3873 5413 3887 5427 0 _1543_.A
rlabel metal2 3853 5453 3867 5467 0 _1543_.B
rlabel metal2 3833 5413 3847 5427 0 _1543_.C
rlabel metal2 3813 5433 3827 5447 0 _1543_.Y
rlabel nsubstratencontact 3916 5292 3916 5292 0 FILL_1__1510_.vdd
rlabel metal1 3904 5522 3936 5538 0 FILL_1__1510_.gnd
rlabel nsubstratencontact 3896 5292 3896 5292 0 FILL_0__1510_.vdd
rlabel metal1 3884 5522 3916 5538 0 FILL_0__1510_.gnd
rlabel nsubstratencontact 4044 5292 4044 5292 0 FILL_1__1491_.vdd
rlabel metal1 4024 5522 4056 5538 0 FILL_1__1491_.gnd
rlabel nsubstratencontact 4024 5292 4024 5292 0 FILL_0__1491_.vdd
rlabel metal1 4004 5522 4036 5538 0 FILL_0__1491_.gnd
rlabel metal1 3924 5522 4016 5538 0 _1510_.gnd
rlabel metal1 3924 5282 4016 5298 0 _1510_.vdd
rlabel metal2 3933 5393 3947 5407 0 _1510_.A
rlabel metal2 3973 5393 3987 5407 0 _1510_.B
rlabel metal2 3953 5413 3967 5427 0 _1510_.Y
rlabel nsubstratencontact 4184 5292 4184 5292 0 FILL_1__1490_.vdd
rlabel metal1 4164 5522 4196 5538 0 FILL_1__1490_.gnd
rlabel nsubstratencontact 4164 5292 4164 5292 0 FILL_0__1490_.vdd
rlabel metal1 4144 5522 4176 5538 0 FILL_0__1490_.gnd
rlabel metal1 4044 5522 4156 5538 0 _1491_.gnd
rlabel metal1 4044 5282 4156 5298 0 _1491_.vdd
rlabel metal2 4133 5433 4147 5447 0 _1491_.A
rlabel metal2 4113 5413 4127 5427 0 _1491_.B
rlabel metal2 4073 5413 4087 5427 0 _1491_.C
rlabel metal2 4093 5433 4107 5447 0 _1491_.Y
rlabel nsubstratencontact 4304 5292 4304 5292 0 FILL_1__1446_.vdd
rlabel metal1 4284 5522 4316 5538 0 FILL_1__1446_.gnd
rlabel nsubstratencontact 4284 5292 4284 5292 0 FILL_0__1446_.vdd
rlabel metal1 4264 5522 4296 5538 0 FILL_0__1446_.gnd
rlabel metal1 4184 5522 4276 5538 0 _1490_.gnd
rlabel metal1 4184 5282 4276 5298 0 _1490_.vdd
rlabel metal2 4253 5393 4267 5407 0 _1490_.A
rlabel metal2 4213 5393 4227 5407 0 _1490_.B
rlabel metal2 4233 5413 4247 5427 0 _1490_.Y
rlabel nsubstratencontact 4416 5292 4416 5292 0 FILL_0__1448_.vdd
rlabel metal1 4404 5522 4436 5538 0 FILL_0__1448_.gnd
rlabel metal1 4304 5522 4416 5538 0 _1446_.gnd
rlabel metal1 4304 5282 4416 5298 0 _1446_.vdd
rlabel metal2 4393 5413 4407 5427 0 _1446_.A
rlabel metal2 4373 5393 4387 5407 0 _1446_.B
rlabel metal2 4353 5413 4367 5427 0 _1446_.C
rlabel metal2 4333 5393 4347 5407 0 _1446_.Y
rlabel nsubstratencontact 4456 5292 4456 5292 0 FILL_2__1448_.vdd
rlabel metal1 4444 5522 4476 5538 0 FILL_2__1448_.gnd
rlabel nsubstratencontact 4436 5292 4436 5292 0 FILL_1__1448_.vdd
rlabel metal1 4424 5522 4456 5538 0 FILL_1__1448_.gnd
rlabel metal1 4464 5522 4576 5538 0 _1448_.gnd
rlabel metal1 4464 5282 4576 5298 0 _1448_.vdd
rlabel metal2 4473 5413 4487 5427 0 _1448_.A
rlabel metal2 4493 5453 4507 5467 0 _1448_.B
rlabel metal2 4513 5413 4527 5427 0 _1448_.C
rlabel metal2 4533 5433 4547 5447 0 _1448_.Y
rlabel metal1 4604 5522 4676 5538 0 _1441_.gnd
rlabel metal1 4604 5282 4676 5298 0 _1441_.vdd
rlabel metal2 4613 5453 4627 5467 0 _1441_.A
rlabel metal2 4633 5413 4647 5427 0 _1441_.Y
rlabel metal1 4704 5522 4816 5538 0 _1445_.gnd
rlabel metal1 4704 5282 4816 5298 0 _1445_.vdd
rlabel metal2 4713 5433 4727 5447 0 _1445_.A
rlabel metal2 4733 5413 4747 5427 0 _1445_.B
rlabel metal2 4773 5413 4787 5427 0 _1445_.C
rlabel metal2 4753 5433 4767 5447 0 _1445_.Y
rlabel metal1 4804 5522 5056 5538 0 _1682_.gnd
rlabel metal1 4804 5282 5056 5298 0 _1682_.vdd
rlabel metal2 4953 5433 4967 5447 0 _1682_.D
rlabel metal2 4913 5433 4927 5447 0 _1682_.CLK
rlabel metal2 4833 5433 4847 5447 0 _1682_.Q
rlabel nsubstratencontact 5056 5292 5056 5292 0 FILL_0__1390_.vdd
rlabel metal1 5044 5522 5076 5538 0 FILL_0__1390_.gnd
rlabel nsubstratencontact 4576 5292 4576 5292 0 FILL_0__1441_.vdd
rlabel metal1 4564 5522 4596 5538 0 FILL_0__1441_.gnd
rlabel nsubstratencontact 4676 5292 4676 5292 0 FILL_0__1445_.vdd
rlabel metal1 4664 5522 4696 5538 0 FILL_0__1445_.gnd
rlabel nsubstratencontact 4596 5292 4596 5292 0 FILL_1__1441_.vdd
rlabel metal1 4584 5522 4616 5538 0 FILL_1__1441_.gnd
rlabel nsubstratencontact 4696 5292 4696 5292 0 FILL_1__1445_.vdd
rlabel metal1 4684 5522 4716 5538 0 FILL_1__1445_.gnd
rlabel metal1 5084 5522 5156 5538 0 _1390_.gnd
rlabel metal1 5084 5282 5156 5298 0 _1390_.vdd
rlabel metal2 5093 5453 5107 5467 0 _1390_.A
rlabel metal2 5113 5413 5127 5427 0 _1390_.Y
rlabel metal1 5424 5522 5536 5538 0 _1633_.gnd
rlabel metal1 5424 5282 5536 5298 0 _1633_.vdd
rlabel metal2 5433 5433 5447 5447 0 _1633_.A
rlabel metal2 5453 5413 5467 5427 0 _1633_.B
rlabel metal2 5493 5413 5507 5427 0 _1633_.C
rlabel metal2 5473 5433 5487 5447 0 _1633_.Y
rlabel metal1 5144 5522 5396 5538 0 _1675_.gnd
rlabel metal1 5144 5282 5396 5298 0 _1675_.vdd
rlabel metal2 5293 5433 5307 5447 0 _1675_.D
rlabel metal2 5253 5433 5267 5447 0 _1675_.CLK
rlabel metal2 5173 5433 5187 5447 0 _1675_.Q
rlabel nsubstratencontact 5536 5292 5536 5292 0 FILL_0__1618_.vdd
rlabel metal1 5524 5522 5556 5538 0 FILL_0__1618_.gnd
rlabel nsubstratencontact 5396 5292 5396 5292 0 FILL_0__1633_.vdd
rlabel metal1 5384 5522 5416 5538 0 FILL_0__1633_.gnd
rlabel nsubstratencontact 5076 5292 5076 5292 0 FILL_1__1390_.vdd
rlabel metal1 5064 5522 5096 5538 0 FILL_1__1390_.gnd
rlabel nsubstratencontact 5556 5292 5556 5292 0 FILL_1__1618_.vdd
rlabel metal1 5544 5522 5576 5538 0 FILL_1__1618_.gnd
rlabel nsubstratencontact 5416 5292 5416 5292 0 FILL_1__1633_.vdd
rlabel metal1 5404 5522 5436 5538 0 FILL_1__1633_.gnd
rlabel metal1 5584 5522 5676 5538 0 _1618_.gnd
rlabel metal1 5584 5282 5676 5298 0 _1618_.vdd
rlabel metal2 5593 5393 5607 5407 0 _1618_.A
rlabel metal2 5633 5393 5647 5407 0 _1618_.B
rlabel metal2 5613 5413 5627 5427 0 _1618_.Y
rlabel metal1 5704 5522 5796 5538 0 _1632_.gnd
rlabel metal1 5704 5282 5796 5298 0 _1632_.vdd
rlabel metal2 5713 5393 5727 5407 0 _1632_.A
rlabel metal2 5753 5393 5767 5407 0 _1632_.B
rlabel metal2 5733 5413 5747 5427 0 _1632_.Y
rlabel nsubstratencontact 5804 5292 5804 5292 0 FILL86850x79350.vdd
rlabel metal1 5784 5522 5816 5538 0 FILL86850x79350.gnd
rlabel nsubstratencontact 5676 5292 5676 5292 0 FILL_0__1632_.vdd
rlabel metal1 5664 5522 5696 5538 0 FILL_0__1632_.gnd
rlabel nsubstratencontact 5696 5292 5696 5292 0 FILL_1__1632_.vdd
rlabel metal1 5684 5522 5716 5538 0 FILL_1__1632_.gnd
rlabel nsubstratencontact 5576 5292 5576 5292 0 FILL_2__1618_.vdd
rlabel metal1 5564 5522 5596 5538 0 FILL_2__1618_.gnd
rlabel nsubstratencontact 44 5768 44 5768 0 FILL_1__1162_.vdd
rlabel metal1 24 5522 56 5538 0 FILL_1__1162_.gnd
rlabel nsubstratencontact 24 5768 24 5768 0 FILL_0__1162_.vdd
rlabel metal1 4 5522 36 5538 0 FILL_0__1162_.gnd
rlabel metal1 44 5522 156 5538 0 _1162_.gnd
rlabel metal1 44 5762 156 5778 0 _1162_.vdd
rlabel metal2 133 5613 147 5627 0 _1162_.A
rlabel metal2 113 5633 127 5647 0 _1162_.B
rlabel metal2 73 5633 87 5647 0 _1162_.C
rlabel metal2 93 5613 107 5627 0 _1162_.Y
rlabel nsubstratencontact 176 5768 176 5768 0 FILL_1__1185_.vdd
rlabel metal1 164 5522 196 5538 0 FILL_1__1185_.gnd
rlabel nsubstratencontact 156 5768 156 5768 0 FILL_0__1185_.vdd
rlabel metal1 144 5522 176 5538 0 FILL_0__1185_.gnd
rlabel metal1 184 5522 296 5538 0 _1185_.gnd
rlabel metal1 184 5762 296 5778 0 _1185_.vdd
rlabel metal2 193 5613 207 5627 0 _1185_.A
rlabel metal2 213 5633 227 5647 0 _1185_.B
rlabel metal2 253 5633 267 5647 0 _1185_.C
rlabel metal2 233 5613 247 5627 0 _1185_.Y
rlabel nsubstratencontact 344 5768 344 5768 0 FILL_2__1161_.vdd
rlabel metal1 324 5522 356 5538 0 FILL_2__1161_.gnd
rlabel nsubstratencontact 324 5768 324 5768 0 FILL_1__1161_.vdd
rlabel metal1 304 5522 336 5538 0 FILL_1__1161_.gnd
rlabel nsubstratencontact 304 5768 304 5768 0 FILL_0__1161_.vdd
rlabel metal1 284 5522 316 5538 0 FILL_0__1161_.gnd
rlabel metal1 344 5522 456 5538 0 _1161_.gnd
rlabel metal1 344 5762 456 5778 0 _1161_.vdd
rlabel metal2 433 5633 447 5647 0 _1161_.A
rlabel metal2 413 5593 427 5607 0 _1161_.B
rlabel metal2 393 5633 407 5647 0 _1161_.C
rlabel metal2 373 5613 387 5627 0 _1161_.Y
rlabel nsubstratencontact 476 5768 476 5768 0 FILL_1__1140_.vdd
rlabel metal1 464 5522 496 5538 0 FILL_1__1140_.gnd
rlabel nsubstratencontact 456 5768 456 5768 0 FILL_0__1140_.vdd
rlabel metal1 444 5522 476 5538 0 FILL_0__1140_.gnd
rlabel metal1 484 5522 596 5538 0 _1140_.gnd
rlabel metal1 484 5762 596 5778 0 _1140_.vdd
rlabel metal2 493 5633 507 5647 0 _1140_.A
rlabel metal2 513 5653 527 5667 0 _1140_.B
rlabel metal2 533 5633 547 5647 0 _1140_.C
rlabel metal2 553 5653 567 5667 0 _1140_.Y
rlabel nsubstratencontact 624 5768 624 5768 0 FILL_1__1158_.vdd
rlabel metal1 604 5522 636 5538 0 FILL_1__1158_.gnd
rlabel nsubstratencontact 604 5768 604 5768 0 FILL_0__1158_.vdd
rlabel metal1 584 5522 616 5538 0 FILL_0__1158_.gnd
rlabel metal1 624 5522 736 5538 0 _1158_.gnd
rlabel metal1 624 5762 736 5778 0 _1158_.vdd
rlabel metal2 713 5613 727 5627 0 _1158_.A
rlabel metal2 693 5633 707 5647 0 _1158_.B
rlabel metal2 653 5633 667 5647 0 _1158_.C
rlabel metal2 673 5613 687 5627 0 _1158_.Y
rlabel nsubstratencontact 764 5768 764 5768 0 FILL_1__954_.vdd
rlabel metal1 744 5522 776 5538 0 FILL_1__954_.gnd
rlabel nsubstratencontact 744 5768 744 5768 0 FILL_0__954_.vdd
rlabel metal1 724 5522 756 5538 0 FILL_0__954_.gnd
rlabel nsubstratencontact 884 5768 884 5768 0 FILL_1__1137_.vdd
rlabel metal1 864 5522 896 5538 0 FILL_1__1137_.gnd
rlabel nsubstratencontact 864 5768 864 5768 0 FILL_0__1137_.vdd
rlabel metal1 844 5522 876 5538 0 FILL_0__1137_.gnd
rlabel metal1 764 5522 856 5538 0 _954_.gnd
rlabel metal1 764 5762 856 5778 0 _954_.vdd
rlabel metal2 833 5653 847 5667 0 _954_.A
rlabel metal2 793 5653 807 5667 0 _954_.B
rlabel metal2 813 5633 827 5647 0 _954_.Y
rlabel nsubstratencontact 1016 5768 1016 5768 0 FILL_1__1135_.vdd
rlabel metal1 1004 5522 1036 5538 0 FILL_1__1135_.gnd
rlabel nsubstratencontact 996 5768 996 5768 0 FILL_0__1135_.vdd
rlabel metal1 984 5522 1016 5538 0 FILL_0__1135_.gnd
rlabel metal1 884 5522 996 5538 0 _1137_.gnd
rlabel metal1 884 5762 996 5778 0 _1137_.vdd
rlabel metal2 973 5633 987 5647 0 _1137_.A
rlabel metal2 953 5593 967 5607 0 _1137_.B
rlabel metal2 933 5633 947 5647 0 _1137_.C
rlabel metal2 913 5613 927 5627 0 _1137_.Y
rlabel nsubstratencontact 1036 5768 1036 5768 0 FILL_2__1135_.vdd
rlabel metal1 1024 5522 1056 5538 0 FILL_2__1135_.gnd
rlabel nsubstratencontact 1144 5768 1144 5768 0 FILL_0__927_.vdd
rlabel metal1 1124 5522 1156 5538 0 FILL_0__927_.gnd
rlabel metal1 1044 5522 1136 5538 0 _1135_.gnd
rlabel metal1 1044 5762 1136 5778 0 _1135_.vdd
rlabel metal2 1093 5613 1107 5627 0 _1135_.B
rlabel metal2 1053 5613 1067 5627 0 _1135_.A
rlabel metal2 1073 5593 1087 5607 0 _1135_.Y
rlabel nsubstratencontact 1184 5768 1184 5768 0 FILL_2__927_.vdd
rlabel metal1 1164 5522 1196 5538 0 FILL_2__927_.gnd
rlabel nsubstratencontact 1164 5768 1164 5768 0 FILL_1__927_.vdd
rlabel metal1 1144 5522 1176 5538 0 FILL_1__927_.gnd
rlabel metal1 1184 5522 1296 5538 0 _927_.gnd
rlabel metal1 1184 5762 1296 5778 0 _927_.vdd
rlabel metal2 1273 5593 1287 5607 0 _927_.A
rlabel metal2 1253 5613 1267 5627 0 _927_.B
rlabel metal2 1213 5633 1227 5647 0 _927_.Y
rlabel nsubstratencontact 1324 5768 1324 5768 0 FILL_1__1134_.vdd
rlabel metal1 1304 5522 1336 5538 0 FILL_1__1134_.gnd
rlabel nsubstratencontact 1304 5768 1304 5768 0 FILL_0__1134_.vdd
rlabel metal1 1284 5522 1316 5538 0 FILL_0__1134_.gnd
rlabel metal1 1324 5522 1436 5538 0 _1134_.gnd
rlabel metal1 1324 5762 1436 5778 0 _1134_.vdd
rlabel metal2 1413 5613 1427 5627 0 _1134_.A
rlabel metal2 1353 5613 1367 5627 0 _1134_.Y
rlabel metal2 1373 5653 1387 5667 0 _1134_.B
rlabel nsubstratencontact 1464 5768 1464 5768 0 FILL_1__1414_.vdd
rlabel metal1 1444 5522 1476 5538 0 FILL_1__1414_.gnd
rlabel nsubstratencontact 1444 5768 1444 5768 0 FILL_0__1414_.vdd
rlabel metal1 1424 5522 1456 5538 0 FILL_0__1414_.gnd
rlabel metal1 1464 5522 1576 5538 0 _1414_.gnd
rlabel metal1 1464 5762 1576 5778 0 _1414_.vdd
rlabel metal2 1553 5633 1567 5647 0 _1414_.A
rlabel metal2 1533 5653 1547 5667 0 _1414_.B
rlabel metal2 1513 5633 1527 5647 0 _1414_.C
rlabel metal2 1493 5653 1507 5667 0 _1414_.Y
rlabel nsubstratencontact 1624 5768 1624 5768 0 FILL_2__1468_.vdd
rlabel metal1 1604 5522 1636 5538 0 FILL_2__1468_.gnd
rlabel nsubstratencontact 1604 5768 1604 5768 0 FILL_1__1468_.vdd
rlabel metal1 1584 5522 1616 5538 0 FILL_1__1468_.gnd
rlabel nsubstratencontact 1584 5768 1584 5768 0 FILL_0__1468_.vdd
rlabel metal1 1564 5522 1596 5538 0 FILL_0__1468_.gnd
rlabel metal1 1624 5522 1736 5538 0 _1468_.gnd
rlabel metal1 1624 5762 1736 5778 0 _1468_.vdd
rlabel metal2 1713 5633 1727 5647 0 _1468_.A
rlabel metal2 1693 5593 1707 5607 0 _1468_.B
rlabel metal2 1673 5633 1687 5647 0 _1468_.C
rlabel metal2 1653 5613 1667 5627 0 _1468_.Y
rlabel nsubstratencontact 1764 5768 1764 5768 0 FILL_1__1403_.vdd
rlabel metal1 1744 5522 1776 5538 0 FILL_1__1403_.gnd
rlabel nsubstratencontact 1744 5768 1744 5768 0 FILL_0__1403_.vdd
rlabel metal1 1724 5522 1756 5538 0 FILL_0__1403_.gnd
rlabel metal1 1764 5522 1876 5538 0 _1403_.gnd
rlabel metal1 1764 5762 1876 5778 0 _1403_.vdd
rlabel metal2 1853 5633 1867 5647 0 _1403_.A
rlabel metal2 1833 5653 1847 5667 0 _1403_.B
rlabel metal2 1813 5633 1827 5647 0 _1403_.C
rlabel metal2 1793 5653 1807 5667 0 _1403_.Y
rlabel nsubstratencontact 1896 5768 1896 5768 0 FILL_1__1399_.vdd
rlabel metal1 1884 5522 1916 5538 0 FILL_1__1399_.gnd
rlabel nsubstratencontact 1876 5768 1876 5768 0 FILL_0__1399_.vdd
rlabel metal1 1864 5522 1896 5538 0 FILL_0__1399_.gnd
rlabel nsubstratencontact 2004 5768 2004 5768 0 FILL_1__1400_.vdd
rlabel metal1 1984 5522 2016 5538 0 FILL_1__1400_.gnd
rlabel nsubstratencontact 1984 5768 1984 5768 0 FILL_0__1400_.vdd
rlabel metal1 1964 5522 1996 5538 0 FILL_0__1400_.gnd
rlabel metal1 2004 5522 2116 5538 0 _1400_.gnd
rlabel metal1 2004 5762 2116 5778 0 _1400_.vdd
rlabel metal2 2093 5613 2107 5627 0 _1400_.A
rlabel metal2 2073 5633 2087 5647 0 _1400_.B
rlabel metal2 2033 5633 2047 5647 0 _1400_.C
rlabel metal2 2053 5613 2067 5627 0 _1400_.Y
rlabel metal1 1904 5522 1976 5538 0 _1399_.gnd
rlabel metal1 1904 5762 1976 5778 0 _1399_.vdd
rlabel metal2 1913 5593 1927 5607 0 _1399_.A
rlabel metal2 1933 5633 1947 5647 0 _1399_.Y
rlabel nsubstratencontact 2136 5768 2136 5768 0 FILL_1__1462_.vdd
rlabel metal1 2124 5522 2156 5538 0 FILL_1__1462_.gnd
rlabel nsubstratencontact 2116 5768 2116 5768 0 FILL_0__1462_.vdd
rlabel metal1 2104 5522 2136 5538 0 FILL_0__1462_.gnd
rlabel metal1 2144 5522 2256 5538 0 _1462_.gnd
rlabel metal1 2144 5762 2256 5778 0 _1462_.vdd
rlabel metal2 2153 5613 2167 5627 0 _1462_.A
rlabel metal2 2173 5633 2187 5647 0 _1462_.B
rlabel metal2 2213 5633 2227 5647 0 _1462_.C
rlabel metal2 2193 5613 2207 5627 0 _1462_.Y
rlabel nsubstratencontact 2276 5768 2276 5768 0 FILL_1__1439_.vdd
rlabel metal1 2264 5522 2296 5538 0 FILL_1__1439_.gnd
rlabel nsubstratencontact 2256 5768 2256 5768 0 FILL_0__1439_.vdd
rlabel metal1 2244 5522 2276 5538 0 FILL_0__1439_.gnd
rlabel nsubstratencontact 2404 5768 2404 5768 0 FILL_0__1464_.vdd
rlabel metal1 2384 5522 2416 5538 0 FILL_0__1464_.gnd
rlabel metal1 2284 5522 2396 5538 0 _1439_.gnd
rlabel metal1 2284 5762 2396 5778 0 _1439_.vdd
rlabel metal2 2293 5633 2307 5647 0 _1439_.A
rlabel metal2 2313 5593 2327 5607 0 _1439_.B
rlabel metal2 2333 5633 2347 5647 0 _1439_.C
rlabel metal2 2353 5613 2367 5627 0 _1439_.Y
rlabel nsubstratencontact 2424 5768 2424 5768 0 FILL_1__1464_.vdd
rlabel metal1 2404 5522 2436 5538 0 FILL_1__1464_.gnd
rlabel nsubstratencontact 2524 5768 2524 5768 0 FILL_0__1465_.vdd
rlabel metal1 2504 5522 2536 5538 0 FILL_0__1465_.gnd
rlabel metal1 2424 5522 2516 5538 0 _1464_.gnd
rlabel metal1 2424 5762 2516 5778 0 _1464_.vdd
rlabel metal2 2493 5653 2507 5667 0 _1464_.A
rlabel metal2 2453 5653 2467 5667 0 _1464_.B
rlabel metal2 2473 5633 2487 5647 0 _1464_.Y
rlabel nsubstratencontact 2544 5768 2544 5768 0 FILL_1__1465_.vdd
rlabel metal1 2524 5522 2556 5538 0 FILL_1__1465_.gnd
rlabel nsubstratencontact 2664 5768 2664 5768 0 FILL_0__1463_.vdd
rlabel metal1 2644 5522 2676 5538 0 FILL_0__1463_.gnd
rlabel metal1 2544 5522 2656 5538 0 _1465_.gnd
rlabel metal1 2544 5762 2656 5778 0 _1465_.vdd
rlabel metal2 2633 5633 2647 5647 0 _1465_.A
rlabel metal2 2613 5653 2627 5667 0 _1465_.B
rlabel metal2 2593 5633 2607 5647 0 _1465_.C
rlabel metal2 2573 5653 2587 5667 0 _1465_.Y
rlabel nsubstratencontact 2684 5768 2684 5768 0 FILL_1__1463_.vdd
rlabel metal1 2664 5522 2696 5538 0 FILL_1__1463_.gnd
rlabel metal1 2684 5522 2796 5538 0 _1463_.gnd
rlabel metal1 2684 5762 2796 5778 0 _1463_.vdd
rlabel metal2 2773 5633 2787 5647 0 _1463_.A
rlabel metal2 2753 5653 2767 5667 0 _1463_.B
rlabel metal2 2733 5633 2747 5647 0 _1463_.C
rlabel metal2 2713 5653 2727 5667 0 _1463_.Y
rlabel nsubstratencontact 2816 5768 2816 5768 0 FILL_1__1459_.vdd
rlabel metal1 2804 5522 2836 5538 0 FILL_1__1459_.gnd
rlabel nsubstratencontact 2796 5768 2796 5768 0 FILL_0__1459_.vdd
rlabel metal1 2784 5522 2816 5538 0 FILL_0__1459_.gnd
rlabel metal1 2824 5522 2916 5538 0 _1459_.gnd
rlabel metal1 2824 5762 2916 5778 0 _1459_.vdd
rlabel metal2 2833 5653 2847 5667 0 _1459_.A
rlabel metal2 2873 5653 2887 5667 0 _1459_.B
rlabel metal2 2853 5633 2867 5647 0 _1459_.Y
rlabel nsubstratencontact 3044 5768 3044 5768 0 FILL_1__1508_.vdd
rlabel metal1 3024 5522 3056 5538 0 FILL_1__1508_.gnd
rlabel nsubstratencontact 2944 5768 2944 5768 0 FILL_1__1492_.vdd
rlabel metal1 2924 5522 2956 5538 0 FILL_1__1492_.gnd
rlabel nsubstratencontact 3024 5768 3024 5768 0 FILL_0__1508_.vdd
rlabel metal1 3004 5522 3036 5538 0 FILL_0__1508_.gnd
rlabel nsubstratencontact 2924 5768 2924 5768 0 FILL_0__1492_.vdd
rlabel metal1 2904 5522 2936 5538 0 FILL_0__1492_.gnd
rlabel metal1 2944 5522 3016 5538 0 _1492_.gnd
rlabel metal1 2944 5762 3016 5778 0 _1492_.vdd
rlabel metal2 2993 5593 3007 5607 0 _1492_.A
rlabel metal2 2973 5633 2987 5647 0 _1492_.Y
rlabel nsubstratencontact 3164 5768 3164 5768 0 FILL_0__1507_.vdd
rlabel metal1 3144 5522 3176 5538 0 FILL_0__1507_.gnd
rlabel metal1 3044 5522 3156 5538 0 _1508_.gnd
rlabel metal1 3044 5762 3156 5778 0 _1508_.vdd
rlabel metal2 3133 5613 3147 5627 0 _1508_.A
rlabel metal2 3113 5633 3127 5647 0 _1508_.B
rlabel metal2 3073 5633 3087 5647 0 _1508_.C
rlabel metal2 3093 5613 3107 5627 0 _1508_.Y
rlabel nsubstratencontact 3204 5768 3204 5768 0 FILL_2__1507_.vdd
rlabel metal1 3184 5522 3216 5538 0 FILL_2__1507_.gnd
rlabel nsubstratencontact 3184 5768 3184 5768 0 FILL_1__1507_.vdd
rlabel metal1 3164 5522 3196 5538 0 FILL_1__1507_.gnd
rlabel metal1 3204 5522 3316 5538 0 _1507_.gnd
rlabel metal1 3204 5762 3316 5778 0 _1507_.vdd
rlabel metal2 3293 5613 3307 5627 0 _1507_.A
rlabel metal2 3233 5613 3247 5627 0 _1507_.Y
rlabel metal2 3253 5653 3267 5667 0 _1507_.B
rlabel nsubstratencontact 3344 5768 3344 5768 0 FILL_1__1506_.vdd
rlabel metal1 3324 5522 3356 5538 0 FILL_1__1506_.gnd
rlabel nsubstratencontact 3324 5768 3324 5768 0 FILL_0__1506_.vdd
rlabel metal1 3304 5522 3336 5538 0 FILL_0__1506_.gnd
rlabel metal1 3344 5522 3436 5538 0 _1506_.gnd
rlabel metal1 3344 5762 3436 5778 0 _1506_.vdd
rlabel metal2 3373 5613 3387 5627 0 _1506_.B
rlabel metal2 3413 5613 3427 5627 0 _1506_.A
rlabel metal2 3393 5593 3407 5607 0 _1506_.Y
rlabel nsubstratencontact 3464 5768 3464 5768 0 FILL_1__1457_.vdd
rlabel metal1 3444 5522 3476 5538 0 FILL_1__1457_.gnd
rlabel nsubstratencontact 3444 5768 3444 5768 0 FILL_0__1457_.vdd
rlabel metal1 3424 5522 3456 5538 0 FILL_0__1457_.gnd
rlabel metal1 3464 5522 3576 5538 0 _1457_.gnd
rlabel metal1 3464 5762 3576 5778 0 _1457_.vdd
rlabel metal2 3553 5633 3567 5647 0 _1457_.A
rlabel metal2 3533 5653 3547 5667 0 _1457_.B
rlabel metal2 3513 5633 3527 5647 0 _1457_.C
rlabel metal2 3493 5653 3507 5667 0 _1457_.Y
rlabel nsubstratencontact 3624 5768 3624 5768 0 FILL_2__1455_.vdd
rlabel metal1 3604 5522 3636 5538 0 FILL_2__1455_.gnd
rlabel nsubstratencontact 3604 5768 3604 5768 0 FILL_1__1455_.vdd
rlabel metal1 3584 5522 3616 5538 0 FILL_1__1455_.gnd
rlabel nsubstratencontact 3584 5768 3584 5768 0 FILL_0__1455_.vdd
rlabel metal1 3564 5522 3596 5538 0 FILL_0__1455_.gnd
rlabel metal1 3624 5522 3696 5538 0 _1455_.gnd
rlabel metal1 3624 5762 3696 5778 0 _1455_.vdd
rlabel metal2 3673 5593 3687 5607 0 _1455_.A
rlabel metal2 3653 5633 3667 5647 0 _1455_.Y
rlabel nsubstratencontact 3724 5768 3724 5768 0 FILL_1__1310_.vdd
rlabel metal1 3704 5522 3736 5538 0 FILL_1__1310_.gnd
rlabel nsubstratencontact 3796 5768 3796 5768 0 FILL_0__1447_.vdd
rlabel metal1 3784 5522 3816 5538 0 FILL_0__1447_.gnd
rlabel nsubstratencontact 3704 5768 3704 5768 0 FILL_0__1310_.vdd
rlabel metal1 3684 5522 3716 5538 0 FILL_0__1310_.gnd
rlabel metal1 3724 5522 3796 5538 0 _1310_.gnd
rlabel metal1 3724 5762 3796 5778 0 _1310_.vdd
rlabel metal2 3773 5593 3787 5607 0 _1310_.A
rlabel metal2 3753 5633 3767 5647 0 _1310_.Y
rlabel nsubstratencontact 3916 5768 3916 5768 0 FILL_1__1454_.vdd
rlabel metal1 3904 5522 3936 5538 0 FILL_1__1454_.gnd
rlabel nsubstratencontact 3816 5768 3816 5768 0 FILL_1__1447_.vdd
rlabel metal1 3804 5522 3836 5538 0 FILL_1__1447_.gnd
rlabel nsubstratencontact 3896 5768 3896 5768 0 FILL_0__1454_.vdd
rlabel metal1 3884 5522 3916 5538 0 FILL_0__1454_.gnd
rlabel metal1 3824 5522 3896 5538 0 _1447_.gnd
rlabel metal1 3824 5762 3896 5778 0 _1447_.vdd
rlabel metal2 3833 5593 3847 5607 0 _1447_.A
rlabel metal2 3853 5633 3867 5647 0 _1447_.Y
rlabel nsubstratencontact 4036 5768 4036 5768 0 FILL_0__1456_.vdd
rlabel metal1 4024 5522 4056 5538 0 FILL_0__1456_.gnd
rlabel metal1 3924 5522 4036 5538 0 _1454_.gnd
rlabel metal1 3924 5762 4036 5778 0 _1454_.vdd
rlabel metal2 3933 5613 3947 5627 0 _1454_.A
rlabel metal2 3953 5633 3967 5647 0 _1454_.B
rlabel metal2 3993 5633 4007 5647 0 _1454_.C
rlabel metal2 3973 5613 3987 5627 0 _1454_.Y
rlabel metal1 4064 5522 4136 5538 0 _1456_.gnd
rlabel metal1 4064 5762 4136 5778 0 _1456_.vdd
rlabel metal2 4073 5593 4087 5607 0 _1456_.A
rlabel metal2 4093 5633 4107 5647 0 _1456_.Y
rlabel metal1 4424 5522 4536 5538 0 _1631_.gnd
rlabel metal1 4424 5762 4536 5778 0 _1631_.vdd
rlabel metal2 4513 5613 4527 5627 0 _1631_.A
rlabel metal2 4493 5633 4507 5647 0 _1631_.B
rlabel metal2 4453 5633 4467 5647 0 _1631_.C
rlabel metal2 4473 5613 4487 5627 0 _1631_.Y
rlabel metal1 4124 5522 4376 5538 0 _1674_.gnd
rlabel metal1 4124 5762 4376 5778 0 _1674_.vdd
rlabel metal2 4273 5613 4287 5627 0 _1674_.D
rlabel metal2 4233 5613 4247 5627 0 _1674_.CLK
rlabel metal2 4153 5613 4167 5627 0 _1674_.Q
rlabel nsubstratencontact 4384 5768 4384 5768 0 FILL_0__1631_.vdd
rlabel metal1 4364 5522 4396 5538 0 FILL_0__1631_.gnd
rlabel nsubstratencontact 4544 5768 4544 5768 0 FILL_0_CLKBUF1_insert3.vdd
rlabel metal1 4524 5522 4556 5538 0 FILL_0_CLKBUF1_insert3.gnd
rlabel nsubstratencontact 4056 5768 4056 5768 0 FILL_1__1456_.vdd
rlabel metal1 4044 5522 4076 5538 0 FILL_1__1456_.gnd
rlabel nsubstratencontact 4404 5768 4404 5768 0 FILL_1__1631_.vdd
rlabel metal1 4384 5522 4416 5538 0 FILL_1__1631_.gnd
rlabel nsubstratencontact 4564 5768 4564 5768 0 FILL_1_CLKBUF1_insert3.vdd
rlabel metal1 4544 5522 4576 5538 0 FILL_1_CLKBUF1_insert3.gnd
rlabel nsubstratencontact 4424 5768 4424 5768 0 FILL_2__1631_.vdd
rlabel metal1 4404 5522 4436 5538 0 FILL_2__1631_.gnd
rlabel nsubstratencontact 4784 5768 4784 5768 0 FILL_0__1646_.vdd
rlabel metal1 4764 5522 4796 5538 0 FILL_0__1646_.gnd
rlabel metal1 4564 5522 4776 5538 0 CLKBUF1_insert3.gnd
rlabel metal1 4564 5762 4776 5778 0 CLKBUF1_insert3.vdd
rlabel metal2 4733 5633 4747 5647 0 CLKBUF1_insert3.A
rlabel metal2 4593 5633 4607 5647 0 CLKBUF1_insert3.Y
rlabel nsubstratencontact 4904 5768 4904 5768 0 FILL_1__1648_.vdd
rlabel metal1 4884 5522 4916 5538 0 FILL_1__1648_.gnd
rlabel nsubstratencontact 4804 5768 4804 5768 0 FILL_1__1646_.vdd
rlabel metal1 4784 5522 4816 5538 0 FILL_1__1646_.gnd
rlabel nsubstratencontact 4884 5768 4884 5768 0 FILL_0__1648_.vdd
rlabel metal1 4864 5522 4896 5538 0 FILL_0__1648_.gnd
rlabel metal1 4904 5522 5016 5538 0 _1648_.gnd
rlabel metal1 4904 5762 5016 5778 0 _1648_.vdd
rlabel metal2 4993 5613 5007 5627 0 _1648_.A
rlabel metal2 4973 5633 4987 5647 0 _1648_.B
rlabel metal2 4933 5633 4947 5647 0 _1648_.C
rlabel metal2 4953 5613 4967 5627 0 _1648_.Y
rlabel metal1 4804 5522 4876 5538 0 _1646_.gnd
rlabel metal1 4804 5762 4876 5778 0 _1646_.vdd
rlabel metal2 4853 5593 4867 5607 0 _1646_.A
rlabel metal2 4833 5633 4847 5647 0 _1646_.Y
rlabel nsubstratencontact 5044 5768 5044 5768 0 FILL_1__1647_.vdd
rlabel metal1 5024 5522 5056 5538 0 FILL_1__1647_.gnd
rlabel nsubstratencontact 5024 5768 5024 5768 0 FILL_0__1647_.vdd
rlabel metal1 5004 5522 5036 5538 0 FILL_0__1647_.gnd
rlabel metal1 5044 5522 5136 5538 0 _1647_.gnd
rlabel metal1 5044 5762 5136 5778 0 _1647_.vdd
rlabel metal2 5113 5653 5127 5667 0 _1647_.A
rlabel metal2 5073 5653 5087 5667 0 _1647_.B
rlabel metal2 5093 5633 5107 5647 0 _1647_.Y
rlabel nsubstratencontact 5156 5768 5156 5768 0 FILL_1__1630_.vdd
rlabel metal1 5144 5522 5176 5538 0 FILL_1__1630_.gnd
rlabel nsubstratencontact 5136 5768 5136 5768 0 FILL_0__1630_.vdd
rlabel metal1 5124 5522 5156 5538 0 FILL_0__1630_.gnd
rlabel metal1 5164 5522 5256 5538 0 _1630_.gnd
rlabel metal1 5164 5762 5256 5778 0 _1630_.vdd
rlabel metal2 5173 5653 5187 5667 0 _1630_.A
rlabel metal2 5213 5653 5227 5667 0 _1630_.B
rlabel metal2 5193 5633 5207 5647 0 _1630_.Y
rlabel nsubstratencontact 5276 5768 5276 5768 0 FILL_1__1724_.vdd
rlabel metal1 5264 5522 5296 5538 0 FILL_1__1724_.gnd
rlabel nsubstratencontact 5256 5768 5256 5768 0 FILL_0__1724_.vdd
rlabel metal1 5244 5522 5276 5538 0 FILL_0__1724_.gnd
rlabel metal1 5284 5522 5396 5538 0 _1724_.gnd
rlabel metal1 5284 5762 5396 5778 0 _1724_.vdd
rlabel metal2 5293 5613 5307 5627 0 _1724_.A
rlabel metal2 5313 5633 5327 5647 0 _1724_.B
rlabel metal2 5353 5633 5367 5647 0 _1724_.C
rlabel metal2 5333 5613 5347 5627 0 _1724_.Y
rlabel nsubstratencontact 5416 5768 5416 5768 0 FILL_1__1727_.vdd
rlabel metal1 5404 5522 5436 5538 0 FILL_1__1727_.gnd
rlabel nsubstratencontact 5396 5768 5396 5768 0 FILL_0__1727_.vdd
rlabel metal1 5384 5522 5416 5538 0 FILL_0__1727_.gnd
rlabel metal1 5424 5522 5496 5538 0 _1727_.gnd
rlabel metal1 5424 5762 5496 5778 0 _1727_.vdd
rlabel metal2 5433 5593 5447 5607 0 _1727_.A
rlabel metal2 5453 5633 5467 5647 0 _1727_.Y
rlabel nsubstratencontact 5516 5768 5516 5768 0 FILL_1__1601_.vdd
rlabel metal1 5504 5522 5536 5538 0 FILL_1__1601_.gnd
rlabel nsubstratencontact 5496 5768 5496 5768 0 FILL_0__1601_.vdd
rlabel metal1 5484 5522 5516 5538 0 FILL_0__1601_.gnd
rlabel metal1 5524 5522 5616 5538 0 _1601_.gnd
rlabel metal1 5524 5762 5616 5778 0 _1601_.vdd
rlabel metal2 5533 5653 5547 5667 0 _1601_.A
rlabel metal2 5573 5653 5587 5667 0 _1601_.B
rlabel metal2 5553 5633 5567 5647 0 _1601_.Y
rlabel metal1 5644 5522 5716 5538 0 _1554_.gnd
rlabel metal1 5644 5762 5716 5778 0 _1554_.vdd
rlabel metal2 5653 5593 5667 5607 0 _1554_.A
rlabel metal2 5673 5633 5687 5647 0 _1554_.Y
rlabel nsubstratencontact 5716 5768 5716 5768 0 FILL85650x82950.vdd
rlabel metal1 5704 5522 5736 5538 0 FILL85650x82950.gnd
rlabel nsubstratencontact 5736 5768 5736 5768 0 FILL85950x82950.vdd
rlabel metal1 5724 5522 5756 5538 0 FILL85950x82950.gnd
rlabel nsubstratencontact 5756 5768 5756 5768 0 FILL86250x82950.vdd
rlabel metal1 5744 5522 5776 5538 0 FILL86250x82950.gnd
rlabel nsubstratencontact 5776 5768 5776 5768 0 FILL86550x82950.vdd
rlabel metal1 5764 5522 5796 5538 0 FILL86550x82950.gnd
rlabel nsubstratencontact 5796 5768 5796 5768 0 FILL86850x82950.vdd
rlabel metal1 5784 5522 5816 5538 0 FILL86850x82950.gnd
rlabel nsubstratencontact 5616 5768 5616 5768 0 FILL_0__1554_.vdd
rlabel metal1 5604 5522 5636 5538 0 FILL_0__1554_.gnd
rlabel nsubstratencontact 5636 5768 5636 5768 0 FILL_1__1554_.vdd
rlabel metal1 5624 5522 5656 5538 0 FILL_1__1554_.gnd
<< end >>
