magic
tech scmos
magscale 1 2
timestamp 1702311544
<< nwell >>
rect -13 154 93 272
<< ntransistor >>
rect 18 14 22 44
rect 38 14 42 54
rect 58 14 62 54
<< ptransistor >>
rect 18 186 22 246
rect 38 166 42 246
rect 58 166 62 246
<< ndiffusion >>
rect 16 14 18 44
rect 22 14 24 44
rect 36 14 38 54
rect 42 14 44 54
rect 56 14 58 54
rect 62 14 64 54
<< pdiffusion >>
rect 16 186 18 246
rect 22 186 24 246
rect 36 168 38 246
rect 24 166 38 168
rect 42 168 44 246
rect 56 168 58 246
rect 42 166 58 168
rect 62 166 64 246
<< ndcontact >>
rect 4 14 16 44
rect 24 14 36 54
rect 44 14 56 54
rect 64 14 76 54
<< pdcontact >>
rect 4 186 16 246
rect 24 168 36 246
rect 44 168 56 246
rect 64 166 76 246
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 254 86 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 58 246 62 250
rect 18 44 22 186
rect 38 164 42 166
rect 58 164 62 166
rect 38 160 62 164
rect 38 155 42 160
rect 38 56 62 60
rect 38 54 42 56
rect 58 54 62 56
rect 18 10 22 14
rect 38 10 42 14
rect 58 10 62 14
<< polycontact >>
rect 6 105 18 117
rect 30 143 42 155
rect 31 60 43 72
<< metal1 >>
rect -6 266 86 268
rect -6 252 86 254
rect 24 246 36 252
rect 64 246 76 252
rect 4 162 12 186
rect 4 156 37 162
rect 30 155 37 156
rect 49 160 56 168
rect 49 154 74 160
rect 3 123 17 137
rect 6 117 17 123
rect 31 72 37 143
rect 66 137 74 154
rect 63 123 77 137
rect 4 60 31 66
rect 66 68 74 123
rect 49 60 74 68
rect 4 44 12 60
rect 49 54 56 60
rect 24 8 36 14
rect 64 8 76 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m1p >>
rect -6 252 86 268
rect 3 123 17 137
rect 63 123 77 137
rect -6 -8 86 8
<< labels >>
rlabel nsubstratencontact 40 260 40 260 0 vdd
port 3 nsew power bidirectional abutment
rlabel psubstratepcontact 40 0 40 0 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 10 131 10 131 0 A
port 1 nsew signal input
rlabel metal1 70 131 70 131 0 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
