magic
tech scmos
timestamp 1555589239
<< checkpaint >>
rect -21 -21 21 21
<< genericcontact >>
rect -1 -1 1 1
<< end >>
