/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module ALU8_Mult(
    inout vdd,
    inout gnd,
    input [7:0] ABCmd_i,
    output [7:0] ACC_o,
    input Flag_i,
    input LoadA_i,
    input LoadB_i,
    input LoadCmd_i,
    input MulH_i,
    input MulL_i,
    input clk,
    input reset
);

wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _873_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _776_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire [7:0] ABCmd_i ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _867_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire LoadA_i ;
wire _388_ ;
wire _600_ ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _864_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _767_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _899_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _861_ ;
wire _441_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _764_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _858_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _896_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _799_ ;
wire _379_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _914_ ;
wire _723_ ;
wire _303_ ;
wire BCD ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _761_ ;
wire _341_ ;
wire clk ;
wire _817_ ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _855_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _893_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _758_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _796_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _852_ ;
wire _432_ ;
wire _908_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _793_ ;
wire _373_ ;
wire _849_ ;
wire _429_ ;
wire _182_ ;
wire _658_ ;
wire _238_ ;
wire _887_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire HC ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _905_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _846_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _884_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _787_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire [3:0] alu_op ;
wire _902_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _805_ ;
wire _65_ ;
wire _614_ ;
wire _843_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _881_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire [7:0] BI ;
wire _784_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _878_ ;
wire _458_ ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _802_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _840_ ;
wire _420_ ;
wire \u_ALU8.AI7  ;
wire _705_ ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _781_ ;
wire _361_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _875_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _778_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire MUL ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _872_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _775_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _869_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _866_ ;
wire _446_ ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _769_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire [7:0] ACC_o ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _634_ ;
wire _214_ ;
wire _863_ ;
wire _443_ ;
wire [7:0] _919_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _766_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _898_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _916_ ;
wire _725_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _895_ ;
wire _475_ ;
wire _284_ ;
wire [7:0] _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _798_ ;
wire _378_ ;
wire _187_ ;
wire _913_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire _816_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _854_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire MulH_i ;
wire _719_ ;
wire _892_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _757_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _795_ ;
wire _375_ ;
wire _184_ ;
wire _889_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _35_ ;
wire _813_ ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _851_ ;
wire _431_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _792_ ;
wire _372_ ;
wire _848_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _886_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _789_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _904_ ;
wire _713_ ;
wire [6:0] ACC ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _845_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _883_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _786_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _901_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire _804_ ;
wire _64_ ;
wire _613_ ;
wire _842_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire Flag_i ;
wire [6:0] AI ;
wire AN ;
wire AV ;
wire AZ ;
wire _783_ ;
wire _363_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire _648_ ;
wire _228_ ;
wire _877_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire LoadB_i ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _645_ ;
wire _225_ ;
wire MUL_bF$buf0 ;
wire MUL_bF$buf1 ;
wire MUL_bF$buf2 ;
wire MUL_bF$buf3 ;
wire MUL_bF$buf4 ;
wire MUL_bF$buf5 ;
wire _874_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _777_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _871_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _774_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _868_ ;
wire _448_ ;
wire LoadCmd_i ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _865_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _768_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _862_ ;
wire _442_ ;
wire _918_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _765_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _859_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _897_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire shr ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _915_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _856_ ;
wire _436_ ;
wire _665_ ;
wire _245_ ;
wire _894_ ;
wire _474_ ;
wire _283_ ;
wire MulL_i ;
wire _759_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _797_ ;
wire _377_ ;
wire _186_ ;
wire _912_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _853_ ;
wire _433_ ;
wire _909_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _891_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _756_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _794_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _888_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _812_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _906_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _791_ ;
wire _371_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _885_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _788_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _903_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire _806_ ;
wire _66_ ;
wire _615_ ;
wire _844_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _882_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire CI ;
wire CO ;
wire _785_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _879_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _497_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _612_ ;
wire reset ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _782_ ;
wire _362_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _876_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire alu_op_2_bF$buf0 ;
wire alu_op_2_bF$buf1 ;
wire alu_op_2_bF$buf2 ;
wire alu_op_2_bF$buf3 ;
wire _779_ ;
wire _359_ ;

FILL FILL_0__1241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1402_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1677_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_18_),
    .CLK(clk_bF$buf2),
    .Q(BI[0])
);

NAND3X1 _1257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_343_),
    .B(_344_),
    .C(_345_),
    .Y(_349_)
);

FILL FILL_0__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1211_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_574_),
    .B(_571_),
    .C(_712_),
    .Y(_575_)
);

NAND2X1 _1066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf5),
    .B(AI[6]),
    .Y(_158_)
);

FILL FILL_0__1526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1020_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_384_),
    .B(_134_),
    .C(_385_),
    .Y(_386_)
);

FILL FILL_0__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_477_),
    .B(_478_),
    .Y(_479_)
);

FILL FILL_0__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1182_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(ABCmd_i[1]),
    .Y(_683_)
);

NAND3X1 _932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf4),
    .B(BI[2]),
    .C(AI[1]),
    .Y(_724_)
);

FILL FILL_1__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[1]),
    .B(_289_),
    .Y(_290_)
);

FILL FILL_0__1238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_801_),
    .B(_790_),
    .Y(_802_)
);

OAI21X1 _1410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_316_),
    .B(_499_),
    .C(_486_),
    .Y(_500_)
);

FILL FILL_1__1572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1208_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_58_),
    .B(_61_),
    .C(_49_),
    .Y(_62_)
);

FILL FILL_1__1381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1085_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_586_),
    .B(_591_),
    .C(_585_),
    .Y(_592_)
);

FILL FILL_1__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_873_),
    .B(_898_),
    .C(_903_),
    .Y(_904_)
);

NAND3X1 _1313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[5]),
    .B(_399_),
    .C(_713_),
    .Y(_404_)
);

FILL FILL_1__1895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1055_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .B(_626_),
    .C(_712_),
    .Y(_629_)
);

NAND3X1 _1122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_146_),
    .B(_213_),
    .C(_209_),
    .Y(_214_)
);

FILL FILL_1__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__926_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf4),
    .B(BI[1]),
    .C(AI[2]),
    .Y(_721_)
);

OAI21X1 _1771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_743_),
    .B(_745_),
    .C(_746_),
    .Y(_747_)
);

OAI21X1 _1351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_438_),
    .B(_441_),
    .C(_377_),
    .Y(_442_)
);

FILL FILL_1__1093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__920_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(_798_),
    .C(_796_),
    .Y(_799_)
);

INVX1 _1407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_),
    .Y(_497_)
);

FILL FILL_1__1569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1149_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_665_),
    .B(_664_),
    .Y(_666_)
);

INVX1 _1160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_251_),
    .Y(_252_)
);

FILL FILL_1__942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[0]),
    .B(LoadB_i),
    .Y(_703_)
);

OR2X2 _1216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_168_),
    .B(_303_),
    .Y(_308_)
);

FILL FILL_0__964_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_50_),
    .B(_51_),
    .Y(_59_)
);

FILL FILL_1__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_830_),
    .Y(_834_)
);

OAI21X1 _1445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_401_),
    .B(_135_),
    .C(_533_),
    .Y(_534_)
);

NAND2X1 _1025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_115_),
    .B(_116_),
    .Y(_117_)
);

FILL FILL_1__1187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__980_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1674_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_15_),
    .CLK(clk_bF$buf1),
    .Q(AI[5])
);

AOI21X1 _1254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_345_),
    .B(_344_),
    .C(_343_),
    .Y(_346_)
);

FILL FILL_0__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AV),
    .Y(_572_)
);

INVX1 _1063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_154_),
    .Y(_155_)
);

FILL FILL_0__1523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1103_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .B(_624_),
    .C(_625_),
    .Y(_626_)
);

NAND3X1 _1119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_205_),
    .C(_206_),
    .Y(_211_)
);

INVX1 _1292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_382_),
    .Y(_383_)
);

FILL FILL_0__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf3),
    .B(BI[3]),
    .C(_858_),
    .Y(_744_)
);

NAND3X1 _1348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_429_),
    .B(_422_),
    .C(_432_),
    .Y(_439_)
);

FILL FILL_0__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1302_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_405_),
    .B(_134_),
    .C(_634_),
    .Y(_663_)
);

OAI21X1 _1157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_247_),
    .B(_248_),
    .C(_246_),
    .Y(_249_)
);

FILL FILL_1__939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86550x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1111_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_475_),
    .Y(_476_)
);

FILL FILL_0__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_207_),
    .B(_186_),
    .C(_206_),
    .Y(_287_)
);

FILL FILL_1__977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _1289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_329_),
    .B(_330_),
    .C(_301_),
    .Y(_380_)
);

FILL FILL_0__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1082_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_182_),
    .Y(_589_)
);

FILL FILL_1__1243_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_188_),
    .B(_189_),
    .C(_187_),
    .Y(_190_)
);

FILL FILL_0__1558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_870_),
    .B(_862_),
    .C(BI[0]),
    .Y(_901_)
);

INVX1 _1310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[5]),
    .Y(_401_)
);

FILL FILL_1__1892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__923_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[3]),
    .B(_717_),
    .Y(_718_)
);

FILL FILL_1__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_868_),
    .B(_791_),
    .C(_795_),
    .D(_794_),
    .Y(_796_)
);

NAND3X1 _1404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_490_),
    .B(_493_),
    .C(_459_),
    .Y(_494_)
);

FILL FILL_1__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadA_i),
    .B(_480_),
    .C(_701_),
    .Y(_16_)
);

AND2X2 _1213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_168_),
    .B(_303_),
    .Y(_305_)
);

FILL FILL_0__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf4),
    .B(BI[2]),
    .C(AI[3]),
    .Y(_56_)
);

FILL FILL_1__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_830_),
    .B(_790_),
    .Y(_831_)
);

OAI21X1 _1442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_475_),
    .B(_484_),
    .C(_479_),
    .Y(_531_)
);

OAI21X1 _1022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_111_),
    .B(_113_),
    .C(_108_),
    .Y(_114_)
);

FILL FILL_1__1184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1079_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1671_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_12_),
    .CLK(clk_bF$buf3),
    .Q(AI[2])
);

INVX1 _1251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_286_),
    .Y(_343_)
);

FILL FILL_0__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_876_),
    .Y(_898_)
);

NAND3X1 _1307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf3),
    .B(AI[5]),
    .C(BI[4]),
    .Y(_398_)
);

FILL FILL_1__1889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1049_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_262_),
    .B(_273_),
    .Y(_569_)
);

NOR2X1 _1060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_150_),
    .B(_151_),
    .Y(_152_)
);

FILL FILL_0__1520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1291_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(_616_),
    .C(_623_),
    .Y(_0_[4])
);

NAND3X1 _1116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_205_),
    .B(_206_),
    .C(_207_),
    .Y(_208_)
);

FILL FILL_1__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL85950x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_862_),
    .B(BI[3]),
    .C(_740_),
    .D(_863_),
    .Y(_741_)
);

AOI21X1 _1345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_434_),
    .B(_435_),
    .C(_395_),
    .Y(_436_)
);

FILL FILL_1__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_614_),
    .C(_659_),
    .Y(_660_)
);

NAND3X1 _1154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_244_),
    .B(_245_),
    .C(_235_),
    .Y(_246_)
);

FILL FILL_1__936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_471_),
    .B(_472_),
    .C(_460_),
    .Y(_473_)
);

FILL FILL_0__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1003_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_799_),
    .B(_816_),
    .C(_815_),
    .Y(_828_)
);

AOI21X1 _1439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_491_),
    .B(_488_),
    .C(_487_),
    .Y(_528_)
);

NOR2X1 _1019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .B(_110_),
    .Y(_111_)
);

AOI21X1 _1192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_209_),
    .B(_146_),
    .C(_216_),
    .Y(_284_)
);

FILL FILL_1__974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1668_ (
    .gnd(gnd),
    .vdd(vdd),
    .R(_1_),
    .S(vdd),
    .D(_0_[7]),
    .CLK(clk_bF$buf4),
    .Q(_919_[7])
);

AOI21X1 _1248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .B(_331_),
    .C(_300_),
    .Y(_340_)
);

FILL FILL_0__996_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_55_),
    .B(_57_),
    .C(_59_),
    .Y(_91_)
);

FILL FILL_0__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1202_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_919_[7]),
    .Y(ACC_o[7])
);

INVX1 _1477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_560_),
    .Y(_566_)
);

AOI21X1 _1057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_100_),
    .B(_97_),
    .C(_94_),
    .Y(_149_)
);

FILL FILL_0__1517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1011_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_286_),
    .B(_341_),
    .C(_376_),
    .Y(_377_)
);

FILL FILL86850x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1240_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .B(_102_),
    .C(_122_),
    .Y(_187_)
);

FILL FILL_0__1555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__920_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf3),
    .Y(_715_)
);

FILL FILL_1__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_280_),
    .Y(_281_)
);

FILL FILL_0__1649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1229_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[6]),
    .B(_792_),
    .Y(_793_)
);

AND2X2 _1401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_473_),
    .B(_470_),
    .Y(_491_)
);

FILL FILL_1__1563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1619_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[5]),
    .B(LoadA_i),
    .Y(_700_)
);

NAND3X1 _1210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf2),
    .B(AI[3]),
    .C(BI[5]),
    .Y(_302_)
);

INVX1 _961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .Y(_53_)
);

FILL FILL_1__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1237_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf0),
    .B(_858_),
    .C(_894_),
    .Y(_895_)
);

NAND2X1 _1304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_390_),
    .B(_394_),
    .Y(_395_)
);

FILL FILL_1__1886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CO),
    .B(_364_),
    .C(_365_),
    .Y(_621_)
);

NAND3X1 _1113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_189_),
    .B(_187_),
    .C(_188_),
    .Y(_205_)
);

FILL FILL_1__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1344_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(shr),
    .B(AI[4]),
    .Y(_738_)
);

AOI21X1 _1342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_426_),
    .B(_428_),
    .C(_423_),
    .Y(_433_)
);

FILL FILL_1__1084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1399_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_784_),
    .B(_787_),
    .C(_783_),
    .Y(_790_)
);

OAI21X1 _1571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_655_),
    .B(_654_),
    .C(_656_),
    .Y(_657_)
);

INVX1 _1151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_242_),
    .Y(_243_)
);

FILL FILL_1__933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1611_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadA_i),
    .B(_387_),
    .C(_698_),
    .Y(_13_)
);

OAI21X1 _1207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .B(_298_),
    .C(_290_),
    .Y(_299_)
);

FILL FILL_0__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf4),
    .B(BI[1]),
    .C(AI[4]),
    .Y(_50_)
);

FILL FILL_1__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1369_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_461_),
    .B(_469_),
    .C(_467_),
    .Y(_470_)
);

FILL FILL_0__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_825_),
    .B(_822_),
    .Y(AZ)
);

AOI21X1 _1436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_457_),
    .B(_505_),
    .C(_524_),
    .Y(_525_)
);

INVX1 _1016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_107_),
    .Y(_108_)
);

FILL FILL_1__1598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1665_ (
    .gnd(gnd),
    .vdd(vdd),
    .R(_1_),
    .S(vdd),
    .D(_0_[4]),
    .CLK(clk_bF$buf4),
    .Q(_919_[4])
);

NAND3X1 _1245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_332_),
    .B(_336_),
    .C(_287_),
    .Y(_337_)
);

FILL FILL_0__993_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_86_),
    .B(_80_),
    .C(_48_),
    .Y(_88_)
);

FILL FILL_0__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_919_[4]),
    .Y(ACC_o[4])
);

NOR2X1 _1474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_360_),
    .B(_448_),
    .Y(_563_)
);

INVX1 _1054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_132_),
    .Y(_146_)
);

FILL FILL_0__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_373_),
    .B(_371_),
    .Y(_374_)
);

FILL FILL_0__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1323_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_735_),
    .Y(ACC[2])
);

NAND3X1 _1339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_422_),
    .B(_429_),
    .C(_381_),
    .Y(_430_)
);

NAND2X1 _1092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_181_),
    .B(_183_),
    .Y(_184_)
);

FILL FILL_0__1552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_653_),
    .B(_357_),
    .C(_281_),
    .Y(_654_)
);

NAND2X1 _1148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .B(_239_),
    .Y(_240_)
);

FILL FILL_0__1608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_751_),
    .B(_771_),
    .C(_757_),
    .Y(HC)
);

OAI21X1 _1377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_462_),
    .B(_407_),
    .C(_466_),
    .Y(_467_)
);

FILL FILL_0__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MulH_i),
    .Y(_712_)
);

FILL FILL_1__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_719_),
    .B(_87_),
    .C(_232_),
    .Y(_278_)
);

FILL FILL_1__968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL85950x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1234_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_167_),
    .B(_171_),
    .C(_175_),
    .Y(_181_)
);

FILL FILL_0__1549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf0),
    .B(BI[1]),
    .C(_858_),
    .Y(_892_)
);

NOR2X1 _1301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_391_),
    .B(_388_),
    .Y(_392_)
);

FILL FILL_1__1883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x32550 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_275_),
    .B(_252_),
    .C(_274_),
    .Y(_618_)
);

NAND3X1 _1110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_191_),
    .B(_201_),
    .C(_200_),
    .Y(_202_)
);

FILL FILL_1__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_784_),
    .B(_787_),
    .Y(_788_)
);

FILL FILL_1__1557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[2]),
    .B(LoadA_i),
    .Y(_697_)
);

NAND3X1 _1204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_291_),
    .B(_295_),
    .C(_294_),
    .Y(_296_)
);

FILL FILL_0__952_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_39_),
    .B(_41_),
    .C(_29_),
    .Y(_47_)
);

FILL FILL_1__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_801_),
    .B(_790_),
    .Y(_823_)
);

NAND2X1 _1433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(_522_),
    .Y(_523_)
);

OAI21X1 _1013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_94_),
    .B(_95_),
    .C(_96_),
    .Y(_105_)
);

FILL FILL_1__1595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1662_ (
    .gnd(gnd),
    .vdd(vdd),
    .R(_1_),
    .S(vdd),
    .D(_0_[1]),
    .CLK(clk_bF$buf4),
    .Q(_919_[1])
);

NAND3X1 _1242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(_326_),
    .C(_328_),
    .Y(_334_)
);

FILL FILL_0__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_84_),
    .B(_83_),
    .Y(_85_)
);

FILL FILL_0__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[0]),
    .B(_888_),
    .Y(_889_)
);

BUFX2 _1891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_919_[1]),
    .Y(ACC_o[1])
);

NAND2X1 _1471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_556_),
    .Y(_560_)
);

NAND2X1 _1051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_142_),
    .B(_139_),
    .Y(_143_)
);

FILL FILL_0__1511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1109_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_603_),
    .B(_614_),
    .C(_613_),
    .Y(_615_)
);

NAND3X1 _1107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_192_),
    .B(_198_),
    .C(_195_),
    .Y(_199_)
);

FILL FILL_1__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_267_),
    .B(_370_),
    .C(MulL_i),
    .Y(_371_)
);

FILL FILL_0__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1320_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918_),
    .B(_727_),
    .C(_732_),
    .Y(_733_)
);

AOI21X1 _1336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_323_),
    .B(_325_),
    .C(_424_),
    .Y(_427_)
);

FILL FILL_1__1498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MulH_i),
    .B(_647_),
    .C(_651_),
    .Y(_652_)
);

INVX1 _1145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_236_),
    .Y(_237_)
);

FILL FILL_1__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_730_),
    .B(_911_),
    .Y(_769_)
);

NOR2X1 _1374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_715_),
    .B(_463_),
    .Y(_464_)
);

FILL FILL_0__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_250_),
    .B(_234_),
    .C(_249_),
    .Y(_275_)
);

FILL FILL_1__965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1659_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_8_),
    .CLK(clk_bF$buf2),
    .Q(BCD)
);

OAI21X1 _1239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_329_),
    .B(_330_),
    .C(_328_),
    .Y(_331_)
);

FILL FILL_0__987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL85950x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1613_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CO),
    .B(_855_),
    .Y(_856_)
);

AOI21X1 _1468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_490_),
    .B(_493_),
    .C(_495_),
    .Y(_557_)
);

NAND3X1 _1048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .B(_127_),
    .C(_126_),
    .Y(_140_)
);

FILL FILL_0__1508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1002_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .Y(_869_)
);

NAND2X1 _1277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(_368_),
    .Y(_369_)
);

FILL FILL_0__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86550x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1231_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_161_),
    .B(_177_),
    .C(_165_),
    .Y(_178_)
);

FILL FILL_0__1546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1393_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_784_),
    .Y(_785_)
);

FILL FILL_1__1554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1029_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadA_i),
    .B(_43_),
    .C(_695_),
    .Y(_10_)
);

AOI22X1 _1201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_116_),
    .B(_174_),
    .C(_171_),
    .D(_167_),
    .Y(_293_)
);

NAND2X1 _952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf0),
    .B(BI[4]),
    .Y(_44_)
);

FILL FILL_1__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1419_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ACC[0]),
    .B(_770_),
    .Y(_820_)
);

NOR2X1 _1430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Flag_i),
    .B(ACC[2]),
    .Y(_520_)
);

NAND3X1 _1010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_91_),
    .B(_98_),
    .C(_101_),
    .Y(_102_)
);

FILL FILL_1__1592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1228_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_58_),
    .B(_61_),
    .C(_49_),
    .Y(_82_)
);

FILL FILL_2__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1296_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[1]),
    .B(BI[1]),
    .C(_864_),
    .Y(_886_)
);

FILL FILL_1__1877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86250x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_560_),
    .B(_512_),
    .Y(_612_)
);

NAND2X1 _1104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[1]),
    .B(_134_),
    .Y(_196_)
);

FILL FILL_1__1686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _1753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_729_),
    .B(_728_),
    .S(_918_),
    .Y(_730_)
);

AND2X2 _1333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_318_),
    .B(_320_),
    .Y(_424_)
);

FILL FILL_1__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf3),
    .B(BI[5]),
    .C(_781_),
    .Y(_782_)
);

AOI21X1 _1562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_614_),
    .C(_603_),
    .Y(_649_)
);

NAND3X1 _1142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_42_),
    .B(_228_),
    .C(_227_),
    .Y(_234_)
);

FILL FILL_1__924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1199_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(ABCmd_i[7]),
    .Y(_694_)
);

FILL FILL_0__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_34_),
    .B(_40_),
    .C(_30_),
    .Y(_41_)
);

OAI21X1 _1791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(_765_),
    .C(_763_),
    .Y(_766_)
);

INVX1 _1371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_460_),
    .Y(_461_)
);

FILL FILL_0__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_805_),
    .B(_806_),
    .C(_817_),
    .Y(_818_)
);

AND2X2 _1427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_264_),
    .B(_269_),
    .Y(_517_)
);

OR2X2 _1007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_92_),
    .B(_93_),
    .Y(_99_)
);

FILL FILL_1__1589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1169_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_246_),
    .Y(_272_)
);

FILL FILL_1__962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1656_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5_),
    .CLK(clk_bF$buf3),
    .Q(alu_op[3])
);

OAI21X1 _1236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_184_),
    .B(_179_),
    .C(_165_),
    .Y(_328_)
);

FILL FILL_0__984_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_78_),
    .B(_76_),
    .Y(_79_)
);

FILL FILL_1__1398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1610_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_850_),
    .B(_819_),
    .C(_818_),
    .Y(_853_)
);

NAND3X1 _1465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_526_),
    .B(_552_),
    .C(_553_),
    .Y(_554_)
);

NAND2X1 _1045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_136_),
    .B(_132_),
    .Y(_137_)
);

FILL FILL_0__1505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[0]),
    .B(alu_op[1]),
    .Y(_866_)
);

OAI21X1 _1274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(HC),
    .B(_364_),
    .C(_365_),
    .Y(_366_)
);

FILL FILL_0__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1314_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_116_),
    .B(_174_),
    .Y(_175_)
);

FILL FILL_0__1543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_644_),
    .B(_645_),
    .Y(_646_)
);

NAND3X1 _1139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_66_),
    .B(_62_),
    .C(_85_),
    .Y(_231_)
);

FILL FILL_0__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1513_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_762_),
    .B(_761_),
    .C(_758_),
    .Y(_763_)
);

INVX1 _1368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_457_),
    .Y(_458_)
);

FILL FILL_0__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL85950x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[0]),
    .Y(_680_)
);

OAI21X1 _1177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_268_),
    .B(_67_),
    .C(_263_),
    .Y(_269_)
);

FILL FILL_1__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1293_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_876_),
    .B(_874_),
    .Y(_883_)
);

FILL FILL_1__1874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_453_),
    .B(_359_),
    .C(_608_),
    .Y(_609_)
);

AOI21X1 _1101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108_),
    .B(_112_),
    .C(_111_),
    .Y(_193_)
);

FILL FILL_1__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf1),
    .B(BI[2]),
    .C(_726_),
    .Y(_727_)
);

AOI21X1 _1330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_409_),
    .B(_413_),
    .C(_420_),
    .Y(_421_)
);

FILL FILL86550x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1387_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[5]),
    .B(_776_),
    .C(_868_),
    .Y(_779_)
);

FILL FILL_1__1548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1196_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BCD),
    .Y(_692_)
);

FILL FILL_0__943_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_36_),
    .B(_37_),
    .C(_32_),
    .Y(_38_)
);

FILL FILL_1__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(_814_),
    .C(_812_),
    .Y(_815_)
);

NAND2X1 _1424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_513_),
    .B(_456_),
    .Y(_514_)
);

NAND3X1 _1004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf1),
    .B(BI[2]),
    .C(AI[4]),
    .Y(_96_)
);

FILL FILL_1__1586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1166_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1653_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2_),
    .CLK(clk_bF$buf3),
    .Q(alu_op[0])
);

OAI21X1 _1233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_316_),
    .B(_317_),
    .C(_313_),
    .Y(_325_)
);

FILL FILL_0__981_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .B(_75_),
    .C(_70_),
    .Y(_76_)
);

FILL FILL_1__1395_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(shr),
    .B(_859_),
    .C(_879_),
    .Y(_881_)
);

NAND2X1 _1882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_848_),
    .B(_849_),
    .Y(_850_)
);

OAI21X1 _1462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_489_),
    .B(_474_),
    .C(_492_),
    .Y(_551_)
);

NOR2X1 _1042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_715_),
    .B(_133_),
    .Y(_134_)
);

FILL FILL_0__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1099_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_525_),
    .B(_555_),
    .C(_605_),
    .Y(_606_)
);

NAND2X1 _1691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[0]),
    .B(_862_),
    .Y(_863_)
);

NOR2X1 _1271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ACC[0]),
    .B(Flag_i),
    .Y(_363_)
);

FILL FILL_0__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1082_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[2]),
    .B(_914_),
    .C(_868_),
    .Y(_917_)
);

OAI21X1 _1327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_417_),
    .B(_26_),
    .C(_314_),
    .Y(_418_)
);

FILL FILL_1__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_110_),
    .B(_168_),
    .C(_171_),
    .Y(_172_)
);

FILL FILL_0__1540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_642_),
    .B(_640_),
    .Y(_643_)
);

NAND3X1 _1136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_222_),
    .B(_223_),
    .C(_224_),
    .Y(_228_)
);

FILL FILL_1__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[4]),
    .B(_759_),
    .Y(_760_)
);

NAND2X1 _1365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_442_),
    .B(_454_),
    .Y(_455_)
);

FILL FILL_0__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86250x64950 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_627_),
    .B(AN),
    .C(MulH_i),
    .Y(_679_)
);

NAND2X1 _1174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .B(_717_),
    .Y(_266_)
);

FILL FILL_1__956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL85950x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1604_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_845_),
    .B(_846_),
    .Y(_847_)
);

NAND2X1 _1459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_543_),
    .B(_546_),
    .Y(_548_)
);

AOI21X1 _1039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_70_),
    .B(_74_),
    .C(_73_),
    .Y(_131_)
);

FILL FILL_1__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1413_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(shr),
    .B(_859_),
    .Y(_860_)
);

NAND2X1 _1268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_351_),
    .B(_347_),
    .Y(_360_)
);

FILL FILL_0__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1222_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_584_),
    .B(_581_),
    .Y(_585_)
);

INVX1 _1077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[4]),
    .Y(_169_)
);

FILL FILL_0__1537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86550x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_864_),
    .B(BI[5]),
    .Y(_776_)
);

FILL FILL_1__1545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(shr),
    .Y(_690_)
);

FILL FILL_0__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_34_),
    .Y(_35_)
);

FILL FILL_1__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1249_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_811_),
    .B(_810_),
    .C(_807_),
    .Y(_812_)
);

NAND3X1 _1421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .B(_506_),
    .C(_510_),
    .Y(_511_)
);

NAND3X1 _1001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf1),
    .B(BI[0]),
    .C(AI[6]),
    .Y(_93_)
);

FILL FILL_1__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1219_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadB_i),
    .B(_133_),
    .C(_710_),
    .Y(_24_)
);

NAND3X1 _1230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_319_),
    .B(_312_),
    .C(_321_),
    .Y(_322_)
);

NOR2X1 _981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_71_),
    .B(_72_),
    .Y(_73_)
);

FILL FILL_1__1392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1287_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(_876_),
    .C(_874_),
    .Y(_878_)
);

FILL FILL_1__1868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_601_),
    .Y(_603_)
);

FILL FILL_1__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[0]),
    .B(_913_),
    .Y(_914_)
);

AOI21X1 _1324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_326_),
    .B(_324_),
    .C(_414_),
    .Y(_415_)
);

FILL FILL_1__1486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_633_),
    .B(_639_),
    .Y(_640_)
);

AOI21X1 _1133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_224_),
    .B(_223_),
    .C(_222_),
    .Y(_225_)
);

FILL FILL_1__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CI),
    .Y(_688_)
);

FILL FILL_0__937_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_),
    .B(_748_),
    .C(_756_),
    .Y(_757_)
);

OAI21X1 _1362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_449_),
    .B(_452_),
    .C(_374_),
    .Y(_0_[1])
);

FILL FILL_0__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1402_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU8.AI7 ),
    .B(_808_),
    .Y(_809_)
);

NAND3X1 _1418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_439_),
    .B(_445_),
    .C(_507_),
    .Y(_508_)
);

NOR2X1 _1591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .B(_354_),
    .Y(_676_)
);

NAND2X1 _1171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_242_),
    .B(_240_),
    .Y(_263_)
);

FILL FILL_1__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1211_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[5]),
    .B(LoadB_i),
    .Y(_709_)
);

NAND2X1 _1227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_313_),
    .B(_318_),
    .Y(_319_)
);

FILL FILL_0__975_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_69_),
    .Y(_70_)
);

FILL FILL_1__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1601_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_842_),
    .B(_816_),
    .Y(_844_)
);

INVX1 _1456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_542_),
    .Y(_545_)
);

NAND3X1 _1036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_102_),
    .B(_106_),
    .C(_123_),
    .Y(_128_)
);

FILL FILL_1__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1410_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf1),
    .Y(_857_)
);

NAND3X1 _1265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .B(_258_),
    .C(_256_),
    .Y(_357_)
);

FILL FILL_0__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1076_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[6]),
    .B(_405_),
    .Y(_582_)
);

NAND3X1 _1074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf5),
    .B(BI[5]),
    .C(AI[2]),
    .Y(_166_)
);

FILL FILL_0__1534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86250x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL),
    .Y(MUL_bF$buf5)
);

BUFX2 BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL),
    .Y(MUL_bF$buf4)
);

BUFX2 BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL),
    .Y(MUL_bF$buf3)
);

BUFX2 BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL),
    .Y(MUL_bF$buf2)
);

BUFX2 BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL),
    .Y(MUL_bF$buf1)
);

FILL FILL_0__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_749_),
    .B(_750_),
    .C(_753_),
    .Y(_754_)
);

OAI21X1 _1359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_360_),
    .B(_359_),
    .C(_351_),
    .Y(_450_)
);

FILL FILL_0__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_658_),
    .B(_673_),
    .Y(_0_[6])
);

INVX1 _1168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_247_),
    .Y(_260_)
);

FILL FILL_0__1628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1381_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_768_),
    .B(_773_),
    .Y(ACC[4])
);

FILL FILL_1__1542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1122_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_413_),
    .B(_416_),
    .C(_486_),
    .Y(_487_)
);

FILL FILL_2__1611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1190_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf0),
    .B(BI[0]),
    .C(AI[4]),
    .Y(_32_)
);

FILL FILL_1__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1284_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .B(alu_op_2_bF$buf1),
    .C(_858_),
    .Y(_875_)
);

FILL FILL_1__1865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1093_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_596_),
    .B(_599_),
    .Y(_600_)
);

FILL FILL_1__1254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86550x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1149_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_910_),
    .B(_905_),
    .C(_906_),
    .Y(_911_)
);

NOR2X1 _1321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_408_),
    .B(_316_),
    .Y(_412_)
);

FILL FILL_1__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1119_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_592_),
    .B(_636_),
    .Y(_637_)
);

AOI21X1 _1130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_27_),
    .C(_722_),
    .Y(_222_)
);

FILL FILL_1__1292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1187_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[3]),
    .Y(_686_)
);

FILL FILL_0__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_724_),
    .B(_28_),
    .C(_723_),
    .Y(_29_)
);

FILL FILL_1__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x68550 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_786_),
    .B(_783_),
    .C(_800_),
    .Y(_806_)
);

OAI21X1 _1415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_496_),
    .B(_501_),
    .C(_459_),
    .Y(_505_)
);

FILL FILL_1__1577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[4]),
    .B(LoadB_i),
    .Y(_707_)
);

NOR2X1 _1224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_314_),
    .B(_315_),
    .Y(_316_)
);

FILL FILL_0__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf5),
    .B(AI[0]),
    .Y(_67_)
);

FILL FILL_1__1386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AN),
    .B(_839_),
    .C(_840_),
    .Y(_841_)
);

NAND2X1 _1453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_541_),
    .B(_540_),
    .Y(_542_)
);

AOI21X1 _1033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_120_),
    .B(_124_),
    .C(_90_),
    .Y(_125_)
);

FILL FILL_1__1195_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_593_),
    .B(_546_),
    .Y(_597_)
);

DFFPOSX1 _1682_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_23_),
    .CLK(clk_bF$buf1),
    .Q(BI[5])
);

INVX1 _1262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_218_),
    .Y(_354_)
);

FILL FILL_0__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1302_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_908_),
    .B(_897_),
    .Y(_909_)
);

OAI22X1 _1318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_316_),
    .B(_408_),
    .C(_407_),
    .D(_403_),
    .Y(_409_)
);

OAI21X1 _1491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_529_),
    .B(_578_),
    .C(_532_),
    .Y(_579_)
);

NAND3X1 _1071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_159_),
    .B(_155_),
    .C(_157_),
    .Y(_163_)
);

FILL FILL_0__1531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1111_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU8.AI7 ),
    .B(_289_),
    .Y(_634_)
);

AOI21X1 _1127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_217_),
    .B(_214_),
    .C(_145_),
    .Y(_219_)
);

FILL FILL_1__1289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1501_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_751_),
    .Y(ACC[3])
);

NAND3X1 _1356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_445_),
    .B(_446_),
    .C(_444_),
    .Y(_447_)
);

FILL FILL_1__1098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1310_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_661_),
    .Y(_671_)
);

INVX1 _1165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .Y(_257_)
);

FILL FILL_1__947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__969_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_477_),
    .B(_478_),
    .Y(_484_)
);

FILL FILL_0__1854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1404_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1679_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_20_),
    .CLK(clk_bF$buf3),
    .Q(BI[2])
);

NAND3X1 _1259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_349_),
    .B(_350_),
    .C(_348_),
    .Y(_351_)
);

FILL FILL_0__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_528_),
    .B(_548_),
    .C(_554_),
    .Y(_576_)
);

NAND3X1 _1068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_159_),
    .B(_154_),
    .C(_157_),
    .Y(_160_)
);

FILL FILL_2__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1281_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_868_),
    .B(_871_),
    .Y(_872_)
);

FILL FILL_1__1862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1022_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_307_),
    .B(_310_),
    .C(_304_),
    .Y(_388_)
);

FILL FILL_0__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86550x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1184_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf2),
    .Y(_684_)
);

FILL FILL_0__931_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf2),
    .B(BI[1]),
    .Y(_26_)
);

FILL FILL_1__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_803_),
    .B(_802_),
    .Y(_804_)
);

OAI21X1 _1412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_496_),
    .B(_501_),
    .C(_495_),
    .Y(_502_)
);

FILL FILL_1__1574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1049_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadB_i),
    .B(_268_),
    .C(_705_),
    .Y(_20_)
);

AOI21X1 _1221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_159_),
    .B(_155_),
    .C(_152_),
    .Y(_313_)
);

OAI21X1 _972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_59_),
    .B(_60_),
    .C(_57_),
    .Y(_64_)
);

FILL FILL_1__1383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1019_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_826_),
    .B(_827_),
    .C(_838_),
    .Y(CO)
);

NAND2X1 _1450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU8.AI7 ),
    .B(_713_),
    .Y(_539_)
);

AOI21X1 _1030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_101_),
    .B(_98_),
    .C(_91_),
    .Y(_122_)
);

FILL FILL_1__1192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1087_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_546_),
    .B(_593_),
    .Y(_594_)
);

FILL FILL_1__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(_893_),
    .C(_891_),
    .Y(_906_)
);

NAND3X1 _1315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[3]),
    .B(_398_),
    .C(_405_),
    .Y(_406_)
);

FILL FILL_1__1897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1546_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_581_),
    .Y(_631_)
);

AOI21X1 _1124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_204_),
    .B(_208_),
    .C(_147_),
    .Y(_216_)
);

FILL FILL86850x54150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__928_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_736_),
    .B(_737_),
    .C(_748_),
    .Y(_749_)
);

OAI21X1 _1353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_343_),
    .B(_443_),
    .C(_337_),
    .Y(_444_)
);

FILL FILL_1__1095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_800_),
    .Y(_801_)
);

INVX1 _1409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_413_),
    .Y(_499_)
);

OAI21X1 _1582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_661_),
    .B(_660_),
    .C(_667_),
    .Y(_668_)
);

OAI21X1 _1162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_253_),
    .C(_719_),
    .Y(_254_)
);

FILL FILL_1__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1202_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[1]),
    .B(LoadB_i),
    .Y(_704_)
);

OAI21X1 _1218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_309_),
    .B(_54_),
    .C(_168_),
    .Y(_310_)
);

FILL FILL_0__966_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_59_),
    .B(_60_),
    .C(_56_),
    .Y(_61_)
);

OAI21X1 _1391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_480_),
    .B(_44_),
    .C(_478_),
    .Y(_481_)
);

FILL FILL_0__1851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1011_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_832_),
    .Y(_836_)
);

INVX1 _1447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_535_),
    .Y(_536_)
);

NAND2X1 _1027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_118_),
    .B(_114_),
    .Y(_119_)
);

FILL FILL_1__1189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1676_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_17_),
    .CLK(clk_bF$buf1),
    .Q(\u_ALU8.AI7 )
);

OAI21X1 _1256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_132_),
    .B(_215_),
    .C(_213_),
    .Y(_348_)
);

FILL FILL_0__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1210_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Flag_i),
    .B(_572_),
    .C(_573_),
    .Y(_574_)
);

OR2X2 _1065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_150_),
    .B(_151_),
    .Y(_157_)
);

FILL FILL_0__1525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1105_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_302_),
    .B(_305_),
    .C(_308_),
    .Y(_385_)
);

FILL FILL_0__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_663_),
    .B(_662_),
    .Y(_665_)
);

FILL FILL_0_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_234_),
    .B(_249_),
    .C(_250_),
    .Y(_251_)
);

FILL FILL_0__1619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1113_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf3),
    .B(\u_ALU8.AI7 ),
    .C(BI[3]),
    .Y(_478_)
);

FILL FILL_0__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1181_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[1]),
    .Y(_682_)
);

INVX1 _931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_722_),
    .Y(_723_)
);

FILL FILL_1__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1342_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_715_),
    .B(_288_),
    .Y(_289_)
);

FILL FILL_1__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86550x32550 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .Y(_591_)
);

FILL FILL_1__1245_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_868_),
    .B(_871_),
    .C(_902_),
    .Y(_903_)
);

AOI21X1 _1312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_400_),
    .B(_402_),
    .C(_397_),
    .Y(_403_)
);

FILL FILL_1__1894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1369_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_627_),
    .B(ACC[5]),
    .Y(_628_)
);

NAND3X1 _1121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_211_),
    .B(_210_),
    .C(_212_),
    .Y(_213_)
);

FILL FILL_1__1283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x75750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf2),
    .B(BI[0]),
    .C(AI[3]),
    .Y(_720_)
);

FILL FILL_1__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1339_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(_745_),
    .C(_743_),
    .Y(_746_)
);

AOI21X1 _1350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_440_),
    .B(_439_),
    .C(_378_),
    .Y(_441_)
);

FILL FILL_1__1092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf2),
    .B(BI[6]),
    .C(_797_),
    .Y(_798_)
);

AOI22X1 _1406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470_),
    .B(_473_),
    .C(_492_),
    .D(_488_),
    .Y(_496_)
);

FILL FILL_1__1568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__941_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadA_i),
    .B(_417_),
    .C(_702_),
    .Y(_17_)
);

INVX1 _1215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_302_),
    .Y(_307_)
);

FILL FILL_0__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_55_),
    .B(_57_),
    .C(_52_),
    .Y(_58_)
);

FILL FILL_1__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1866_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_829_),
    .B(_832_),
    .C(_831_),
    .Y(_833_)
);

AOI21X1 _1444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_476_),
    .B(_481_),
    .C(_483_),
    .Y(_533_)
);

INVX1 _1024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_110_),
    .Y(_116_)
);

FILL FILL_1__1186_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1673_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_14_),
    .CLK(clk_bF$buf2),
    .Q(AI[4])
);

OAI21X1 _1253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_339_),
    .B(_340_),
    .C(_287_),
    .Y(_345_)
);

FILL FILL86250x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _1729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[1]),
    .B(_869_),
    .S(alu_op[0]),
    .Y(_900_)
);

OR2X2 _1309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_398_),
    .B(_399_),
    .Y(_400_)
);

AOI21X1 _1482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_270_),
    .B(_569_),
    .C(_570_),
    .Y(_571_)
);

NAND3X1 _1062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf1),
    .B(BI[2]),
    .C(AI[5]),
    .Y(_154_)
);

FILL FILL_0__1522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .B(_624_),
    .C(MulL_i),
    .Y(_625_)
);

OAI21X1 _1118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .B(_125_),
    .C(_141_),
    .Y(_210_)
);

NAND2X1 _1291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[2]),
    .B(_289_),
    .Y(_382_)
);

FILL FILL_0__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_742_),
    .B(_741_),
    .C(_738_),
    .Y(_743_)
);

AOI21X1 _1347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_430_),
    .B(_437_),
    .C(_379_),
    .Y(_438_)
);

FILL FILL_1__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_592_),
    .B(_636_),
    .C(_642_),
    .Y(_662_)
);

AOI21X1 _1156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .B(_245_),
    .C(_244_),
    .Y(_248_)
);

FILL FILL_1__938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL85650x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf3),
    .B(AI[5]),
    .C(BI[5]),
    .Y(_475_)
);

FILL FILL_0__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1005_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_191_),
    .B(_285_),
    .C(_200_),
    .Y(_286_)
);

FILL FILL_1__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86250x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1204_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_561_),
    .B(_567_),
    .Y(_568_)
);

NAND3X1 _1059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf5),
    .B(BI[0]),
    .C(\u_ALU8.AI7 ),
    .Y(_151_)
);

FILL FILL_0__1519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1013_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_378_),
    .Y(_379_)
);

FILL FILL_0__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1081_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_417_),
    .B(_182_),
    .C(_587_),
    .Y(_588_)
);

FILL FILL_1__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_161_),
    .B(_165_),
    .C(_184_),
    .Y(_189_)
);

FILL FILL_2__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__922_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_715_),
    .B(_716_),
    .Y(_717_)
);

FILL FILL_1__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[6]),
    .B(_792_),
    .C(_868_),
    .Y(_795_)
);

NAND3X1 _1403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_492_),
    .B(_488_),
    .C(_491_),
    .Y(_493_)
);

FILL FILL_1__1565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1145_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[6]),
    .B(LoadA_i),
    .Y(_701_)
);

NOR2X1 _1212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_168_),
    .B(_303_),
    .Y(_304_)
);

FILL FILL_0__960_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_53_),
    .B(_54_),
    .C(_50_),
    .Y(_55_)
);

FILL FILL_1__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1269_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_816_),
    .B(_800_),
    .Y(_830_)
);

INVX1 _1441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_529_),
    .Y(_530_)
);

INVX1 _1021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .Y(_113_)
);

FILL FILL_1__1183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1670_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_11_),
    .CLK(clk_bF$buf0),
    .Q(AI[1])
);

AOI21X1 _1250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_337_),
    .B(_341_),
    .C(_286_),
    .Y(_342_)
);

FILL FILL_0__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_896_),
    .B(_884_),
    .Y(_897_)
);

INVX1 _1306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_396_),
    .Y(_397_)
);

FILL FILL_1__1888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x28950 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(_622_),
    .Y(_623_)
);

AND2X2 _1115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_199_),
    .B(_202_),
    .Y(_207_)
);

FILL FILL_1__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1277_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[3]),
    .B(_739_),
    .Y(_740_)
);

OAI21X1 _1344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_424_),
    .B(_330_),
    .C(_414_),
    .Y(_435_)
);

FILL FILL_1__1086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_601_),
    .B(_602_),
    .C(_650_),
    .Y(_659_)
);

OAI21X1 _1153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_722_),
    .B(_28_),
    .C(_724_),
    .Y(_245_)
);

FILL FILL_1__935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1613_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadA_i),
    .B(_463_),
    .C(_699_),
    .Y(_14_)
);

AOI21X1 _1209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_161_),
    .B(_177_),
    .C(_180_),
    .Y(_301_)
);

FILL FILL_0__957_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_468_),
    .B(_465_),
    .Y(_472_)
);

FILL FILL_0__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BCD),
    .B(_824_),
    .Y(_827_)
);

INVX1 _1438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_526_),
    .Y(_527_)
);

NAND3X1 _1018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf1),
    .B(BI[3]),
    .C(AI[3]),
    .Y(_110_)
);

OAI21X1 _1191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .B(_282_),
    .C(_218_),
    .Y(_283_)
);

FILL FILL_1__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1667_ (
    .gnd(gnd),
    .vdd(vdd),
    .R(_1_),
    .S(vdd),
    .D(_0_[6]),
    .CLK(clk_bF$buf4),
    .Q(_919_[6])
);

AOI21X1 _1247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_334_),
    .B(_335_),
    .C(_333_),
    .Y(_339_)
);

FILL FILL_0__995_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_82_),
    .C(_62_),
    .Y(_90_)
);

FILL FILL_0__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1201_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_919_[6]),
    .Y(ACC_o[6])
);

AOI21X1 _1476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_564_),
    .B(_455_),
    .C(_512_),
    .Y(_565_)
);

OAI21X1 _1056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_121_),
    .B(_123_),
    .C(_106_),
    .Y(_148_)
);

FILL FILL_0__1516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1010_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_338_),
    .B(_375_),
    .Y(_376_)
);

FILL FILL_0__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_185_),
    .C(_148_),
    .Y(_186_)
);

FILL FILL_0__1554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1104_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_772_),
    .B(HC),
    .Y(_773_)
);

OAI21X1 _1379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_463_),
    .B(_135_),
    .C(_468_),
    .Y(_469_)
);

FILL FILL_0__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1172_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[0]),
    .B(_713_),
    .Y(_714_)
);

FILL FILL_1__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1333_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .B(_255_),
    .C(_279_),
    .Y(_280_)
);

FILL FILL_2__1402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_864_),
    .B(BI[6]),
    .Y(_792_)
);

OAI21X1 _1400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .B(_489_),
    .C(_474_),
    .Y(_490_)
);

FILL FILL_1__1562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1618_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_50_),
    .B(_51_),
    .Y(_52_)
);

FILL FILL_1__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1305_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_893_),
    .Y(_894_)
);

OAI21X1 _1303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_392_),
    .B(_393_),
    .C(_382_),
    .Y(_394_)
);

FILL FILL86250x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Flag_i),
    .B(ACC[4]),
    .Y(_620_)
);

OAI21X1 _1112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_186_),
    .C(_203_),
    .Y(_204_)
);

FILL FILL86850x82950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1169_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_911_),
    .B(_730_),
    .Y(_737_)
);

OAI21X1 _1341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_300_),
    .B(_431_),
    .C(_334_),
    .Y(_432_)
);

FILL FILL_1__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1398_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_789_),
    .Y(ACC[5])
);

FILL FILL_1__1559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1139_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ACC[6]),
    .B(_627_),
    .Y(_656_)
);

OAI21X1 _1150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_716_),
    .B(_26_),
    .C(_236_),
    .Y(_242_)
);

FILL FILL_1__932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1610_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[3]),
    .B(LoadA_i),
    .Y(_698_)
);

AND2X2 _1206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_293_),
    .B(_292_),
    .Y(_298_)
);

FILL FILL_0__954_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_30_),
    .B(_40_),
    .C(_35_),
    .Y(_49_)
);

FILL FILL_1__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1017_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_824_),
    .B(AN),
    .Y(_825_)
);

NOR3X1 _1435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_496_),
    .B(_501_),
    .C(_459_),
    .Y(_524_)
);

NAND3X1 _1015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf1),
    .B(BI[5]),
    .C(AI[1]),
    .Y(_107_)
);

FILL FILL_1__1597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1246_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1664_ (
    .gnd(gnd),
    .vdd(vdd),
    .R(_1_),
    .S(vdd),
    .D(_0_[3]),
    .CLK(clk_bF$buf4),
    .Q(_919_[3])
);

NAND3X1 _1244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_333_),
    .B(_335_),
    .C(_334_),
    .Y(_336_)
);

FILL FILL_0__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_80_),
    .B(_86_),
    .C(_48_),
    .Y(_87_)
);

FILL FILL_0__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x14550 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_919_[3]),
    .Y(ACC_o[3])
);

INVX1 _1473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_511_),
    .Y(_562_)
);

INVX1 _1053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .Y(_145_)
);

FILL FILL_0__1513_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .Y(_617_)
);

OAI21X1 _1109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_716_),
    .B(_135_),
    .C(_193_),
    .Y(_201_)
);

AOI21X1 _1282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_372_),
    .B(_365_),
    .C(MulH_i),
    .Y(_373_)
);

FILL FILL_0__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1322_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_731_),
    .B(_734_),
    .Y(_735_)
);

NAND3X1 _1338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_428_),
    .B(_423_),
    .C(_426_),
    .Y(_429_)
);

OAI21X1 _1091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_725_),
    .B(_182_),
    .C(_172_),
    .Y(_183_)
);

FILL FILL_0__1551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(_356_),
    .Y(_653_)
);

INVX1 _1147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_238_),
    .Y(_239_)
);

FILL FILL_1__929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL85650x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1101_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BCD),
    .B(_770_),
    .Y(_771_)
);

INVX1 _1376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_465_),
    .Y(_466_)
);

FILL FILL_0__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1330_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_253_),
    .C(_220_),
    .Y(_277_)
);

FILL FILL_1__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[0]),
    .B(_869_),
    .C(_870_),
    .Y(_871_)
);

AND2X2 _1279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_266_),
    .B(_265_),
    .Y(_370_)
);

FILL FILL_0__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .B(_156_),
    .C(_149_),
    .Y(_180_)
);

FILL FILL_2__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887_),
    .B(_890_),
    .C(_885_),
    .Y(_891_)
);

NAND2X1 _1300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[6]),
    .B(_384_),
    .Y(_391_)
);

FILL FILL_1__1882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86250x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86550x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1395_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(HC),
    .B(_772_),
    .C(_774_),
    .Y(_787_)
);

FILL FILL_1__1556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1625_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadA_i),
    .B(_716_),
    .C(_696_),
    .Y(_11_)
);

OAI21X1 _1203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_725_),
    .B(_135_),
    .C(_293_),
    .Y(_295_)
);

FILL FILL_0__951_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_45_),
    .B(_719_),
    .Y(_46_)
);

FILL FILL_1__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1365_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_821_),
    .B(ACC[4]),
    .Y(_822_)
);

OAI21X1 _1432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_520_),
    .B(_521_),
    .C(_519_),
    .Y(_522_)
);

NAND3X1 _1012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_100_),
    .B(_97_),
    .C(_99_),
    .Y(_104_)
);

FILL FILL_1__1594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1661_ (
    .gnd(gnd),
    .vdd(vdd),
    .R(_1_),
    .S(vdd),
    .D(_0_[0]),
    .CLK(clk_bF$buf4),
    .Q(_919_[0])
);

AND2X2 _1241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_296_),
    .B(_299_),
    .Y(_333_)
);

OAI21X1 _992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .B(_75_),
    .C(_69_),
    .Y(_84_)
);

FILL FILL_0__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[1]),
    .Y(_888_)
);

FILL FILL_1__1879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_919_[0]),
    .Y(ACC_o[0])
);

NAND3X1 _1470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_550_),
    .B(_554_),
    .C(_558_),
    .Y(_559_)
);

NAND3X1 _1050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .B(_141_),
    .C(_140_),
    .Y(_142_)
);

FILL FILL_0__1510_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_283_),
    .B(_612_),
    .C(_563_),
    .Y(_614_)
);

NAND2X1 _1106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_193_),
    .B(_197_),
    .Y(_198_)
);

FILL FILL_1__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1337_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(_727_),
    .C(_918_),
    .Y(_732_)
);

OAI21X1 _1335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_424_),
    .B(_330_),
    .C(_425_),
    .Y(_426_)
);

FILL FILL_1__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1566_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_648_),
    .B(_649_),
    .C(_650_),
    .Y(_651_)
);

NAND3X1 _1144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf0),
    .B(BI[0]),
    .C(AI[2]),
    .Y(_236_)
);

FILL FILL_1__926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_),
    .B(_757_),
    .C(_767_),
    .Y(_768_)
);

INVX1 _1373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[4]),
    .Y(_463_)
);

FILL FILL_0__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1413_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_818_),
    .B(_819_),
    .Y(AN)
);

OAI21X1 _1429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_267_),
    .B(_517_),
    .C(_518_),
    .Y(_519_)
);

NAND3X1 _1009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_100_),
    .B(_96_),
    .C(_99_),
    .Y(_101_)
);

NAND3X1 _1182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_262_),
    .C(_273_),
    .Y(_274_)
);

FILL FILL_1__964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1658_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_7_),
    .CLK(clk_bF$buf2),
    .Q(shr)
);

AOI21X1 _1238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_321_),
    .B(_319_),
    .C(_312_),
    .Y(_330_)
);

FILL FILL_0__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_64_),
    .B(_65_),
    .C(_63_),
    .Y(_81_)
);

FILL FILL_0__1871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1612_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853_),
    .B(_852_),
    .Y(_855_)
);

NAND2X1 _1467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_525_),
    .B(_555_),
    .Y(_556_)
);

OAI21X1 _1047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_125_),
    .C(_138_),
    .Y(_139_)
);

FILL FILL_0__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1001_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(shr),
    .Y(_868_)
);

OAI21X1 _1276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_363_),
    .B(_366_),
    .C(_367_),
    .Y(_368_)
);

FILL FILL_0__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_173_),
    .Y(_177_)
);

FILL FILL_0__1545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(_680_),
    .C(_681_),
    .Y(_2_)
);

INVX1 _1179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_270_),
    .Y(_271_)
);

FILL FILL_2__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1392_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_780_),
    .B(_782_),
    .C(_783_),
    .Y(_784_)
);

FILL FILL_1__1553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1609_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[0]),
    .B(LoadA_i),
    .Y(_695_)
);

NAND2X1 _1200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[2]),
    .B(_134_),
    .Y(_292_)
);

INVX1 _951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[0]),
    .Y(_43_)
);

FILL FILL_1__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86250x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1295_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(shr),
    .B(AI[2]),
    .Y(_885_)
);

FILL FILL_1__1876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1036_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_351_),
    .B(_448_),
    .C(_447_),
    .Y(_611_)
);

OAI21X1 _1103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_716_),
    .B(_135_),
    .C(_194_),
    .Y(_195_)
);

FILL FILL_1__1685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf0),
    .B(_858_),
    .C(_728_),
    .Y(_729_)
);

AND2X2 _1332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_394_),
    .B(_390_),
    .Y(_423_)
);

FILL FILL_1__1494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86550x68550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf3),
    .B(BI[5]),
    .C(_858_),
    .Y(_781_)
);

INVX1 _1561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .Y(_648_)
);

NAND3X1 _1141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .B(_87_),
    .C(_232_),
    .Y(_233_)
);

FILL FILL_1__923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1198_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(_692_),
    .C(_693_),
    .Y(_8_)
);

FILL FILL_0__945_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_38_),
    .Y(_40_)
);

FILL FILL_1__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf2),
    .B(BI[4]),
    .C(_764_),
    .Y(_765_)
);

NAND2X1 _1370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[7]),
    .B(_384_),
    .Y(_460_)
);

FILL FILL_0__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1410_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_816_),
    .Y(_817_)
);

NAND2X1 _1426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_514_),
    .B(_515_),
    .Y(_516_)
);

OAI21X1 _1006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_94_),
    .B(_95_),
    .C(_97_),
    .Y(_98_)
);

FILL FILL_1__1588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x21750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1655_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4_),
    .CLK(clk_bF$buf3),
    .Q(alu_op[2])
);

NAND3X1 _1235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(_326_),
    .C(_301_),
    .Y(_327_)
);

FILL FILL_0__983_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_69_),
    .B(_74_),
    .C(_77_),
    .Y(_78_)
);

FILL FILL_1__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_843_),
    .B(_844_),
    .C(_851_),
    .Y(_852_)
);

NAND2X1 _1464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_548_),
    .B(_528_),
    .Y(_553_)
);

OAI21X1 _1044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_43_),
    .B(_135_),
    .C(_131_),
    .Y(_136_)
);

FILL FILL_0__1504_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .B(_864_),
    .Y(_865_)
);

INVX2 _1273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MulL_i),
    .Y(_365_)
);

FILL FILL_0__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1313_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf1),
    .B(BI[2]),
    .C(_858_),
    .Y(_726_)
);

OAI21X1 _1329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_312_),
    .B(_419_),
    .C(_324_),
    .Y(_420_)
);

INVX1 _1082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_168_),
    .Y(_174_)
);

FILL FILL_0__1542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_643_),
    .B(_630_),
    .Y(_645_)
);

OAI21X1 _1138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_81_),
    .B(_82_),
    .C(_79_),
    .Y(_230_)
);

FILL FILL_0__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1512_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[4]),
    .B(_759_),
    .C(_868_),
    .Y(_762_)
);

OAI21X1 _1367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_382_),
    .B(_393_),
    .C(_386_),
    .Y(_457_)
);

FILL FILL_0__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1321_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX4 _1596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(reset),
    .Y(_1_)
);

INVX1 _1176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .Y(_268_)
);

FILL FILL_1__958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1224_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_586_),
    .B(_585_),
    .Y(_587_)
);

OAI21X1 _1079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_169_),
    .B(_37_),
    .C(_170_),
    .Y(_171_)
);

FILL FILL_0__1539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1292_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882_),
    .Y(ACC[0])
);

FILL FILL86250x46950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1509_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_556_),
    .B(_607_),
    .C(_454_),
    .D(_442_),
    .Y(_608_)
);

INVX1 _1100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_191_),
    .Y(_192_)
);

FILL FILL_1__1262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x3750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1386_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_862_),
    .B(BI[5]),
    .C(_777_),
    .D(_863_),
    .Y(_778_)
);

FILL FILL_1__1547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1195_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(_690_),
    .C(_691_),
    .Y(_7_)
);

FILL FILL_0__942_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf2),
    .B(AI[3]),
    .Y(_37_)
);

FILL FILL_1__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1356_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf2),
    .B(BI[7]),
    .C(_813_),
    .Y(_814_)
);

INVX1 _1423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_512_),
    .Y(_513_)
);

AND2X2 _1003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_92_),
    .B(_93_),
    .Y(_95_)
);

FILL FILL_1__1585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1165_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadB_i),
    .B(_288_),
    .C(_711_),
    .Y(_25_)
);

NAND2X1 _1232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .B(_318_),
    .Y(_324_)
);

FILL FILL_0__980_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_74_),
    .Y(_75_)
);

FILL FILL_1__1394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1289_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_879_),
    .B(_861_),
    .Y(_880_)
);

OR2X2 _1881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_847_),
    .B(\u_ALU8.AI7 ),
    .Y(_849_)
);

NAND3X1 _1461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_527_),
    .B(_549_),
    .C(_547_),
    .Y(_550_)
);

INVX1 _1041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[6]),
    .Y(_133_)
);

FILL FILL_0__1501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1098_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_556_),
    .B(_508_),
    .Y(_605_)
);

FILL FILL86550x54150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[1]),
    .Y(_862_)
);

NAND2X1 _1270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_353_),
    .B(_361_),
    .Y(_362_)
);

FILL FILL_0__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1310_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_862_),
    .B(BI[2]),
    .C(_915_),
    .D(_863_),
    .Y(_916_)
);

INVX2 _1326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU8.AI7 ),
    .Y(_417_)
);

FILL FILL_1__1488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_641_),
    .B(_638_),
    .C(_637_),
    .Y(_642_)
);

NOR2X1 _1135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .B(_226_),
    .Y(_227_)
);

FILL FILL_1__1297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__939_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_864_),
    .B(BI[4]),
    .Y(_759_)
);

NAND2X1 _1364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_447_),
    .B(_351_),
    .Y(_454_)
);

FILL FILL_0__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__933_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_676_),
    .B(_358_),
    .C(_677_),
    .Y(_678_)
);

NAND2X1 _1173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[1]),
    .B(_68_),
    .Y(_265_)
);

FILL FILL_1__955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[6]),
    .B(LoadB_i),
    .Y(_710_)
);

OAI21X1 _1229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_316_),
    .B(_317_),
    .C(_320_),
    .Y(_321_)
);

FILL FILL_0__977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1603_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(_812_),
    .Y(_846_)
);

NAND3X1 _1458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_543_),
    .B(_546_),
    .C(_528_),
    .Y(_547_)
);

NAND2X1 _1038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[6]),
    .B(_68_),
    .Y(_130_)
);

FILL FILL_1__993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_857_),
    .B(_858_),
    .C(CI),
    .Y(_859_)
);

AOI21X1 _1267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_355_),
    .B(_358_),
    .C(_354_),
    .Y(_359_)
);

FILL FILL_0__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .B(_540_),
    .C(_583_),
    .Y(_584_)
);

NAND3X1 _1076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf5),
    .B(AI[4]),
    .C(BI[4]),
    .Y(_168_)
);

FILL FILL_0__1536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL85950x82950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1383_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(shr),
    .B(AI[6]),
    .Y(_775_)
);

FILL FILL_1__1544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1124_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_488_),
    .Y(_489_)
);

FILL FILL_0__1859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1192_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(_688_),
    .C(_689_),
    .Y(_6_)
);

NOR2X1 _942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_32_),
    .B(_33_),
    .Y(_34_)
);

FILL FILL_1__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU8.AI7 ),
    .B(_808_),
    .C(_868_),
    .Y(_811_)
);

OAI21X1 _1420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_379_),
    .B(_509_),
    .C(_439_),
    .Y(_510_)
);

NAND3X1 _1000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf1),
    .B(BI[1]),
    .C(AI[5]),
    .Y(_92_)
);

FILL FILL_1__1582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86250x32550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1218_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf4),
    .B(BI[3]),
    .C(AI[2]),
    .Y(_72_)
);

FILL FILL_1__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1286_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf3),
    .B(_858_),
    .Y(_877_)
);

FILL FILL_1__1867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1095_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_576_),
    .B(_596_),
    .C(_599_),
    .Y(_602_)
);

FILL FILL_1__1256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86550x75750 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .Y(_913_)
);

NAND2X1 _1323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_413_),
    .B(_409_),
    .Y(_414_)
);

FILL FILL_1__1485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1065_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_637_),
    .Y(_639_)
);

NAND3X1 _1132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_30_),
    .B(_38_),
    .C(_35_),
    .Y(_224_)
);

FILL FILL_1__1294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1189_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(_686_),
    .C(_687_),
    .Y(_5_)
);

FILL FILL_0__936_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_30_),
    .Y(_31_)
);

INVX1 _1781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_746_),
    .Y(_756_)
);

OAI21X1 _1361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_451_),
    .B(_450_),
    .C(MulH_i),
    .Y(_452_)
);

FILL FILL_0__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1592_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_864_),
    .B(BI[7]),
    .Y(_808_)
);

NAND2X1 _1417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .B(_506_),
    .Y(_507_)
);

FILL FILL_1__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1159_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(_674_),
    .Y(_675_)
);

NAND3X1 _1170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_246_),
    .B(_260_),
    .C(_261_),
    .Y(_262_)
);

FILL FILL_1__952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1210_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[5]),
    .Y(_708_)
);

NOR2X1 _1226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_316_),
    .B(_317_),
    .Y(_318_)
);

FILL FILL_0__974_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[5]),
    .B(_68_),
    .Y(_69_)
);

FILL FILL_1__1388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1600_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_816_),
    .B(_842_),
    .Y(_843_)
);

INVX1 _1455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_537_),
    .Y(_544_)
);

OAI21X1 _1035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_122_),
    .B(_121_),
    .C(_119_),
    .Y(_127_)
);

FILL FILL_1__1197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__990_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1684_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_25_),
    .CLK(clk_bF$buf2),
    .Q(BI[7])
);

NAND2X1 _1264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .B(_258_),
    .Y(_356_)
);

FILL FILL_0__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1304_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[5]),
    .B(_289_),
    .Y(_581_)
);

NAND3X1 _1073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_164_),
    .B(_162_),
    .C(_163_),
    .Y(_165_)
);

FILL FILL_0__1533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1113_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_582_),
    .B(_634_),
    .C(_635_),
    .Y(_636_)
);

INVX1 _1129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_724_),
    .Y(_221_)
);

FILL FILL_0__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1503_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_735_),
    .B(_909_),
    .C(_752_),
    .Y(_753_)
);

AOI21X1 _1358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_353_),
    .B(_351_),
    .C(_448_),
    .Y(_449_)
);

FILL FILL_0__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1312_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MulH_i),
    .B(_672_),
    .C(_668_),
    .Y(_673_)
);

AND2X2 _1167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_258_),
    .B(_144_),
    .Y(_259_)
);

FILL FILL_1__949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1121_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_485_),
    .B(_482_),
    .Y(_486_)
);

FILL FILL_0__1856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1283_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_867_),
    .B(_872_),
    .C(_873_),
    .Y(_874_)
);

FILL FILL_1__1864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .B(_389_),
    .C(_386_),
    .Y(_390_)
);

FILL FILL_0__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1092_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_579_),
    .B(_598_),
    .C(_597_),
    .Y(_599_)
);

FILL FILL_1__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_893_),
    .B(_891_),
    .Y(_910_)
);

NAND3X1 _1320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_397_),
    .B(_402_),
    .C(_400_),
    .Y(_411_)
);

FILL FILL_1__1482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1186_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(_684_),
    .C(_685_),
    .Y(_4_)
);

FILL FILL_0__933_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_27_),
    .Y(_28_)
);

FILL FILL_1__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1416_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_799_),
    .Y(_805_)
);

NAND3X1 _1414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_490_),
    .B(_493_),
    .C(_495_),
    .Y(_504_)
);

FILL FILL_1__1576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1156_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadB_i),
    .B(_309_),
    .C(_706_),
    .Y(_21_)
);

NAND3X1 _1223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf5),
    .B(\u_ALU8.AI7 ),
    .C(BI[1]),
    .Y(_315_)
);

FILL FILL_0__971_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_63_),
    .B(_65_),
    .C(_64_),
    .Y(_66_)
);

FILL FILL_1__1385_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_833_),
    .B(_837_),
    .Y(_840_)
);

OAI21X1 _1452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_417_),
    .B(_44_),
    .C(_538_),
    .Y(_541_)
);

OAI21X1 _1032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_122_),
    .B(_121_),
    .C(_123_),
    .Y(_124_)
);

FILL FILL_0_CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_594_),
    .B(_595_),
    .C(_580_),
    .Y(_596_)
);

DFFPOSX1 _1681_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_22_),
    .CLK(clk_bF$buf0),
    .Q(BI[4])
);

NAND2X1 _1261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_352_),
    .B(_283_),
    .Y(_353_)
);

FILL FILL_0__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1301_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_905_),
    .B(_907_),
    .Y(_908_)
);

NAND3X1 _1317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf0),
    .B(\u_ALU8.AI7 ),
    .C(BI[2]),
    .Y(_408_)
);

FILL FILL_1__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1059_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_534_),
    .B(_532_),
    .Y(_578_)
);

OAI21X1 _1070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .B(_95_),
    .C(_99_),
    .Y(_162_)
);

FILL FILL_0__1530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1110_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_631_),
    .B(_583_),
    .C(_632_),
    .Y(_633_)
);

NAND3X1 _1126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_145_),
    .B(_214_),
    .C(_217_),
    .Y(_218_)
);

FILL FILL_1__1288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1500_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_750_),
    .B(_749_),
    .Y(_751_)
);

NAND3X1 _1355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_379_),
    .B(_437_),
    .C(_430_),
    .Y(_446_)
);

FILL FILL_1__1097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_606_),
    .B(_669_),
    .C(_609_),
    .Y(_670_)
);

INVX1 _1164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .Y(_256_)
);

FILL FILL_1__946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__968_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_477_),
    .B(_478_),
    .Y(_483_)
);

FILL FILL_0__1853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1013_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_837_),
    .B(_833_),
    .Y(_838_)
);

NAND2X1 _1449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[5]),
    .B(_405_),
    .Y(_538_)
);

AOI21X1 _1029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_104_),
    .B(_105_),
    .C(_103_),
    .Y(_121_)
);

FILL FILL_1__984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1678_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_19_),
    .CLK(clk_bF$buf0),
    .Q(BI[1])
);

NAND3X1 _1258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_286_),
    .B(_341_),
    .C(_337_),
    .Y(_350_)
);

FILL FILL_0__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(_568_),
    .C(_575_),
    .Y(_0_[3])
);

OAI21X1 _1067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_36_),
    .B(_158_),
    .C(_151_),
    .Y(_159_)
);

FILL FILL_0__1527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1021_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[3]),
    .Y(_387_)
);

FILL FILL_0__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1183_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(_682_),
    .C(_683_),
    .Y(_3_)
);

FILL FILL_0__930_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[2]),
    .Y(_725_)
);

FILL FILL_1__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1344_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_290_),
    .Y(_291_)
);

FILL FILL_2__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_783_),
    .B(_800_),
    .C(_786_),
    .Y(_803_)
);

AOI21X1 _1411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_500_),
    .C(_474_),
    .Y(_501_)
);

FILL FILL_1__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[2]),
    .B(LoadB_i),
    .Y(_705_)
);

NAND2X1 _1220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_306_),
    .B(_311_),
    .Y(_312_)
);

AOI21X1 _971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_31_),
    .B(_38_),
    .C(_34_),
    .Y(_63_)
);

FILL FILL_1__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1086_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_592_),
    .B(_588_),
    .Y(_593_)
);

FILL FILL_1__1247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86550x82950 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_874_),
    .B(_899_),
    .C(_904_),
    .D(_860_),
    .Y(_905_)
);

AND2X2 _1314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf3),
    .B(AI[6]),
    .Y(_405_)
);

FILL FILL_1__1896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_579_),
    .B(_598_),
    .C(_594_),
    .Y(_630_)
);

AOI21X1 _1123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_212_),
    .B(_211_),
    .C(_210_),
    .Y(_215_)
);

FILL FILL_1__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__927_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_747_),
    .Y(_748_)
);

AOI21X1 _1352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_332_),
    .B(_336_),
    .C(_287_),
    .Y(_443_)
);

FILL FILL_1__1094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_796_),
    .B(_798_),
    .C(_799_),
    .Y(_800_)
);

NAND3X1 _1408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .B(_413_),
    .C(_497_),
    .Y(_498_)
);

INVX1 _1581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_666_),
    .Y(_667_)
);

AOI21X1 _1161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_230_),
    .B(_231_),
    .C(_229_),
    .Y(_253_)
);

FILL FILL_1__943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1201_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadB_i),
    .B(_53_),
    .C(_703_),
    .Y(_18_)
);

INVX1 _1217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[3]),
    .Y(_309_)
);

FILL FILL_0__965_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_55_),
    .Y(_60_)
);

FILL FILL_1__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1379_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[6]),
    .Y(_480_)
);

FILL FILL_0__1850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1010_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_786_),
    .B(_783_),
    .C(_834_),
    .Y(_835_)
);

NAND3X1 _1446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_530_),
    .B(_534_),
    .C(_532_),
    .Y(_535_)
);

NAND3X1 _1026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_107_),
    .B(_112_),
    .C(_117_),
    .Y(_118_)
);

FILL FILL_1__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1400_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1675_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_16_),
    .CLK(clk_bF$buf1),
    .Q(AI[6])
);

OAI21X1 _1255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_346_),
    .B(_342_),
    .C(_284_),
    .Y(_347_)
);

FILL FILL_0__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Flag_i),
    .B(ACC[3]),
    .C(_365_),
    .Y(_573_)
);

OAI21X1 _1064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_152_),
    .B(_153_),
    .C(_155_),
    .Y(_156_)
);

FILL FILL86850x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1104_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_37_),
    .Y(_384_)
);

FILL FILL_0__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1333_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf3),
    .B(BI[3]),
    .C(_744_),
    .Y(_745_)
);

OAI21X1 _1349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_433_),
    .B(_436_),
    .C(_381_),
    .Y(_440_)
);

FILL FILL_0__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1303_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_662_),
    .B(_663_),
    .Y(_664_)
);

OAI21X1 _1158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_225_),
    .B(_47_),
    .C(_46_),
    .Y(_250_)
);

FILL FILL_0__1618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1112_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf3),
    .B(AI[6]),
    .C(BI[4]),
    .Y(_477_)
);

FILL FILL_0__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_720_),
    .B(_721_),
    .Y(_722_)
);

FILL FILL_1__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1341_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[7]),
    .Y(_288_)
);

FILL FILL_1__978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1150_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL),
    .Y(MUL_bF$buf0)
);

BUFX2 BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[2]),
    .Y(alu_op_2_bF$buf3)
);

BUFX2 BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[2]),
    .Y(alu_op_2_bF$buf2)
);

BUFX2 BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[2]),
    .Y(alu_op_2_bF$buf1)
);

BUFX2 BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[2]),
    .Y(alu_op_2_bF$buf0)
);

FILL FILL_0__1885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1083_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU8.AI7 ),
    .B(_589_),
    .Y(_590_)
);

FILL FILL_1__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[7]),
    .B(_68_),
    .Y(_191_)
);

FILL FILL_0__1559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1139_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_901_),
    .B(_900_),
    .Y(_902_)
);

OAI21X1 _1311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_401_),
    .B(_44_),
    .C(_399_),
    .Y(_402_)
);

FILL FILL_1__1893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1109_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Flag_i),
    .B(MulL_i),
    .Y(_627_)
);

OAI21X1 _1120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_186_),
    .C(_207_),
    .Y(_212_)
);

FILL FILL_1__1282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__924_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_718_),
    .B(_714_),
    .Y(_719_)
);

FILL FILL_1__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1091_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf2),
    .B(BI[6]),
    .C(_858_),
    .Y(_797_)
);

OAI21X1 _1405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_395_),
    .B(_421_),
    .C(_426_),
    .Y(_495_)
);

FILL FILL_1__1567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__940_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[7]),
    .B(LoadA_i),
    .Y(_702_)
);

OAI21X1 _1214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_304_),
    .B(_305_),
    .C(_302_),
    .Y(_306_)
);

FILL FILL_0__962_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_56_),
    .Y(_57_)
);

FILL FILL_1__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_870_),
    .B(_868_),
    .Y(_832_)
);

NAND3X1 _1443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[5]),
    .B(_134_),
    .C(_531_),
    .Y(_532_)
);

INVX1 _1023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .Y(_115_)
);

FILL FILL_1__1185_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1672_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_13_),
    .CLK(clk_bF$buf0),
    .Q(AI[3])
);

NAND3X1 _1252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_332_),
    .B(_336_),
    .C(_338_),
    .Y(_344_)
);

FILL FILL_0__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1063_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf0),
    .B(_858_),
    .C(_898_),
    .Y(_899_)
);

NAND3X1 _1308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf0),
    .B(AI[6]),
    .C(BI[3]),
    .Y(_399_)
);

OAI21X1 _1481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_270_),
    .B(_569_),
    .C(MulL_i),
    .Y(_570_)
);

AND2X2 _1061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_150_),
    .B(_151_),
    .Y(_153_)
);

FILL FILL_0__1521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1101_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(_279_),
    .Y(_624_)
);

NAND3X1 _1117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_208_),
    .B(_204_),
    .C(_147_),
    .Y(_209_)
);

FILL FILL_1__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1279_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_333_),
    .B(_335_),
    .C(_380_),
    .Y(_381_)
);

FILL FILL_2__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1330_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[3]),
    .B(_739_),
    .C(_868_),
    .Y(_742_)
);

OAI21X1 _1346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_436_),
    .B(_433_),
    .C(_432_),
    .Y(_437_)
);

FILL FILL_1__1088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1300_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_646_),
    .C(_645_),
    .Y(_661_)
);

NAND2X1 _1155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[3]),
    .B(_68_),
    .Y(_247_)
);

FILL FILL_1__937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__959_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470_),
    .B(_473_),
    .Y(_474_)
);

FILL FILL_0__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_197_),
    .B(_194_),
    .Y(_285_)
);

FILL FILL_1__975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x43350 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1669_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_10_),
    .CLK(clk_bF$buf0),
    .Q(AI[0])
);

OAI21X1 _1249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_339_),
    .B(_340_),
    .C(_338_),
    .Y(_341_)
);

FILL FILL_0__997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_562_),
    .B(_565_),
    .C(_566_),
    .Y(_567_)
);

NAND3X1 _1058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf5),
    .B(BI[1]),
    .C(AI[6]),
    .Y(_150_)
);

FILL FILL_0__1518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_290_),
    .B(_298_),
    .C(_294_),
    .Y(_378_)
);

FILL FILL_0__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1241_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_180_),
    .B(_179_),
    .C(_177_),
    .Y(_188_)
);

FILL FILL_0__1556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__921_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[1]),
    .Y(_716_)
);

FILL FILL_1__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1335_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_862_),
    .B(BI[6]),
    .C(_793_),
    .D(_863_),
    .Y(_794_)
);

INVX1 _1402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .Y(_492_)
);

FILL FILL_1__1564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1039_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadA_i),
    .B(_401_),
    .C(_700_),
    .Y(_15_)
);

NAND3X1 _1211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf5),
    .B(AI[5]),
    .C(BI[3]),
    .Y(_303_)
);

NAND2X1 _962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf2),
    .B(AI[5]),
    .Y(_54_)
);

FILL FILL_1__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1009_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_828_),
    .Y(_829_)
);

NAND2X1 _1440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[7]),
    .B(_464_),
    .Y(_529_)
);

OAI21X1 _1020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_725_),
    .B(_44_),
    .C(_110_),
    .Y(_112_)
);

FILL FILL_1__1182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1238_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _1725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_895_),
    .B(_894_),
    .S(_891_),
    .Y(_896_)
);

NAND3X1 _1305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf3),
    .B(AI[4]),
    .C(BI[5]),
    .Y(_396_)
);

FILL FILL_1__1887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86250x68550 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_620_),
    .B(_621_),
    .C(_619_),
    .Y(_622_)
);

NAND3X1 _1114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_185_),
    .C(_148_),
    .Y(_206_)
);

FILL FILL_1__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1276_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_864_),
    .B(BI[3]),
    .Y(_739_)
);

NAND2X1 _1343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_427_),
    .B(_425_),
    .Y(_434_)
);

FILL FILL_1__1085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1154_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU8.AI7 ),
    .Y(_791_)
);

NAND2X1 _1572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(_657_),
    .Y(_658_)
);

OAI21X1 _1152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_241_),
    .B(_243_),
    .C(_240_),
    .Y(_244_)
);

FILL FILL_1__934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1383_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[4]),
    .B(LoadA_i),
    .Y(_699_)
);

NAND2X1 _1208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_299_),
    .B(_296_),
    .Y(_300_)
);

FILL FILL_0__956_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf2),
    .B(BI[0]),
    .C(AI[5]),
    .Y(_51_)
);

NOR2X1 _1381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_465_),
    .B(_468_),
    .Y(_471_)
);

FILL FILL_0__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1001_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_819_),
    .B(_818_),
    .Y(_826_)
);

OAI21X1 _1437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_460_),
    .B(_472_),
    .C(_467_),
    .Y(_526_)
);

NAND3X1 _1017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf1),
    .B(BI[4]),
    .C(AI[2]),
    .Y(_109_)
);

FILL FILL_1__1599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1179_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_256_),
    .B(_281_),
    .C(_259_),
    .Y(_282_)
);

FILL FILL_1__972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1666_ (
    .gnd(gnd),
    .vdd(vdd),
    .R(_1_),
    .S(vdd),
    .D(_0_[5]),
    .CLK(clk_bF$buf3),
    .Q(_919_[5])
);

AOI21X1 _1246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_205_),
    .C(_190_),
    .Y(_338_)
);

FILL FILL_0__994_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_719_),
    .B(_88_),
    .C(_87_),
    .Y(_89_)
);

FILL FILL_0__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x64950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1200_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _1895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_919_[5]),
    .Y(ACC_o[5])
);

NAND2X1 _1475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_283_),
    .B(_563_),
    .Y(_564_)
);

AOI21X1 _1055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_138_),
    .B(_140_),
    .C(_129_),
    .Y(_147_)
);

FILL FILL_0__1515_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_332_),
    .B(_336_),
    .Y(_375_)
);

FILL FILL_0__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_180_),
    .B(_179_),
    .C(_184_),
    .Y(_185_)
);

FILL FILL_0__1553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_280_),
    .B(_356_),
    .C(MulL_i),
    .Y(_655_)
);

NAND2X1 _1149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .B(_68_),
    .Y(_241_)
);

FILL FILL_0__1609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1103_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_767_),
    .Y(_772_)
);

AOI21X1 _1378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_397_),
    .B(_402_),
    .C(_462_),
    .Y(_468_)
);

FILL FILL_0__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1171_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf3),
    .B(BI[4]),
    .Y(_713_)
);

FILL FILL_1__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1332_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_251_),
    .B(_278_),
    .C(_277_),
    .Y(_279_)
);

FILL FILL_1__969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86550x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1235_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf0),
    .B(BI[1]),
    .C(_892_),
    .Y(_893_)
);

AND2X2 _1302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_388_),
    .B(_391_),
    .Y(_393_)
);

FILL FILL_1__1884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1359_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MulL_i),
    .B(_618_),
    .C(_617_),
    .Y(_619_)
);

NAND2X1 _1111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_202_),
    .B(_199_),
    .Y(_203_)
);

FILL FILL_1__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1329_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_732_),
    .Y(_736_)
);

AOI21X1 _1340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(_326_),
    .C(_328_),
    .Y(_431_)
);

FILL FILL_1__1082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1397_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_786_),
    .B(_788_),
    .Y(_789_)
);

FILL FILL_1__1558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1207_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadA_i),
    .B(_725_),
    .C(_697_),
    .Y(_12_)
);

NOR2X1 _1205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_292_),
    .B(_293_),
    .Y(_297_)
);

FILL FILL_0__953_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_46_),
    .B(_47_),
    .C(_42_),
    .Y(_48_)
);

FILL FILL_1__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1367_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_806_),
    .B(_823_),
    .C(_789_),
    .Y(_824_)
);

OAI21X1 _1434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(_516_),
    .C(_523_),
    .Y(_0_[2])
);

NAND3X1 _1014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_104_),
    .B(_105_),
    .C(_103_),
    .Y(_106_)
);

FILL FILL_1__1596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1176_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _1663_ (
    .gnd(gnd),
    .vdd(vdd),
    .R(_1_),
    .S(vdd),
    .D(_0_[2]),
    .CLK(clk_bF$buf4),
    .Q(_919_[2])
);

OAI21X1 _1243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_329_),
    .B(_330_),
    .C(_301_),
    .Y(_335_)
);

FILL FILL_0__991_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_81_),
    .B(_82_),
    .C(_85_),
    .Y(_86_)
);

FILL FILL_0__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1474_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[1]),
    .B(_889_),
    .C(_868_),
    .Y(_890_)
);

BUFX2 _1892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_919_[2]),
    .Y(ACC_o[2])
);

NAND3X1 _1472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_511_),
    .B(_560_),
    .C(_514_),
    .Y(_561_)
);

NAND2X1 _1052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .B(_143_),
    .Y(_144_)
);

FILL FILL_0__1512_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_615_),
    .B(_610_),
    .Y(_616_)
);

NAND2X1 _1108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_197_),
    .B(_194_),
    .Y(_200_)
);

MUX2X1 _1281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AN),
    .B(ACC[1]),
    .S(Flag_i),
    .Y(_372_)
);

FILL FILL_0__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1321_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_906_),
    .B(_733_),
    .C(_897_),
    .Y(_734_)
);

NAND2X1 _1337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_414_),
    .B(_427_),
    .Y(_428_)
);

FILL FILL_1__1499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1079_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf0),
    .B(BI[5]),
    .Y(_182_)
);

FILL FILL_0__1550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_629_),
    .B(_652_),
    .Y(_0_[5])
);

NAND3X1 _1146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf0),
    .B(BI[1]),
    .C(AI[1]),
    .Y(_238_)
);

FILL FILL_1__928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1100_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_769_),
    .B(_737_),
    .C(_909_),
    .Y(_770_)
);

NAND2X1 _1375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[6]),
    .B(_464_),
    .Y(_465_)
);

FILL FILL_0__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1415_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _1184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_275_),
    .B(_274_),
    .C(_252_),
    .Y(_276_)
);

FILL FILL_1__966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1614_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_854_),
    .B(_856_),
    .Y(AV)
);

OAI21X1 _1469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_458_),
    .B(_557_),
    .C(_504_),
    .Y(_558_)
);

NAND3X1 _1049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_120_),
    .B(_124_),
    .C(_90_),
    .Y(_141_)
);

FILL FILL_0__1509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1003_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[0]),
    .Y(_870_)
);

OAI21X1 _1278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(_362_),
    .C(_369_),
    .Y(_0_[0])
);

FILL FILL_0__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1232_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_163_),
    .B(_164_),
    .C(_162_),
    .Y(_179_)
);

FILL FILL85650x82950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1394_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_774_),
    .B(_768_),
    .C(_785_),
    .Y(_786_)
);

FILL FILL_1__1555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[1]),
    .B(LoadA_i),
    .Y(_696_)
);

OR2X2 _1202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_293_),
    .B(_292_),
    .Y(_294_)
);

FILL FILL_0__950_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_43_),
    .B(_44_),
    .C(_718_),
    .Y(_45_)
);

FILL FILL_1__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1259_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_751_),
    .B(_820_),
    .Y(_821_)
);

OAI21X1 _1431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AZ),
    .B(_364_),
    .C(_365_),
    .Y(_521_)
);

OAI21X1 _1011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_56_),
    .B(_60_),
    .C(_52_),
    .Y(_103_)
);

FILL FILL_1__1593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1229_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1660_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_9_),
    .CLK(clk_bF$buf1),
    .Q(MUL)
);

NAND3X1 _1240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_300_),
    .B(_331_),
    .C(_327_),
    .Y(_332_)
);

NAND3X1 _991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_74_),
    .B(_77_),
    .C(_70_),
    .Y(_83_)
);

FILL FILL_0__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1297_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_862_),
    .B(BI[1]),
    .C(_886_),
    .D(_863_),
    .Y(_887_)
);

FILL FILL_1__1878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1527_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_556_),
    .B(_607_),
    .C(_612_),
    .D(_611_),
    .Y(_613_)
);

INVX1 _1105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_196_),
    .Y(_197_)
);

FILL FILL_1__1687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1267_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_730_),
    .B(_911_),
    .Y(_731_)
);

AND2X2 _1334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_409_),
    .B(_413_),
    .Y(_425_)
);

FILL FILL_1__1496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1076_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_645_),
    .B(_644_),
    .Y(_650_)
);

NAND3X1 _1143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_27_),
    .C(_723_),
    .Y(_235_)
);

FILL FILL_1__925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(_715_),
    .C(_694_),
    .Y(_9_)
);

FILL FILL_0__947_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_763_),
    .B(_765_),
    .C(_766_),
    .Y(_767_)
);

NOR2X1 _1372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_398_),
    .B(_399_),
    .Y(_462_)
);

FILL FILL_0__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1412_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_799_),
    .B(_816_),
    .C(_802_),
    .Y(_819_)
);

NOR2X1 _1428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(_271_),
    .Y(_518_)
);

OAI21X1 _1008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_36_),
    .B(_54_),
    .C(_93_),
    .Y(_100_)
);

OAI21X1 _1181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_248_),
    .B(_272_),
    .C(_247_),
    .Y(_273_)
);

FILL FILL_1__963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1657_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6_),
    .CLK(clk_bF$buf3),
    .Q(CI)
);

AOI22X1 _1237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_306_),
    .B(_311_),
    .C(_324_),
    .D(_325_),
    .Y(_329_)
);

FILL FILL_0__985_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_66_),
    .B(_62_),
    .C(_79_),
    .Y(_80_)
);

FILL FILL_1__1399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1611_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_852_),
    .B(_853_),
    .C(_841_),
    .Y(_854_)
);

NAND2X1 _1466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_554_),
    .B(_550_),
    .Y(_555_)
);

INVX1 _1046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .Y(_138_)
);

FILL FILL_0__1506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1000_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .B(_866_),
    .C(_863_),
    .D(_865_),
    .Y(_867_)
);

NAND3X1 _1275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .B(MulL_i),
    .C(_68_),
    .Y(_367_)
);

FILL FILL_0__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1315_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_166_),
    .B(_171_),
    .C(_175_),
    .Y(_176_)
);

FILL FILL_0__1544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1514_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf3),
    .B(BI[4]),
    .C(_858_),
    .Y(_764_)
);

AOI21X1 _1369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_423_),
    .B(_428_),
    .C(_415_),
    .Y(_459_)
);

FILL FILL_0__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1323_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[0]),
    .B(LoadCmd_i),
    .Y(_681_)
);

NAND3X1 _1178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_267_),
    .B(_269_),
    .C(_264_),
    .Y(_270_)
);

FILL FILL_0__1638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1391_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(_782_),
    .C(_780_),
    .Y(_783_)
);

FILL FILL_1__1552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1608_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_41_),
    .B(_29_),
    .C(_39_),
    .Y(_42_)
);

FILL FILL_1__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1294_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_861_),
    .B(_883_),
    .C(_878_),
    .Y(_884_)
);

FILL FILL_1__1875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1035_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .B(_606_),
    .C(_609_),
    .Y(_610_)
);

INVX1 _1102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_193_),
    .Y(_194_)
);

FILL FILL_1__1264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1159_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_727_),
    .Y(_728_)
);

OAI21X1 _1331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .B(_421_),
    .C(_395_),
    .Y(_422_)
);

FILL FILL_1__1493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1388_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_779_),
    .B(_778_),
    .C(_775_),
    .Y(_780_)
);

FILL FILL_1__1549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1129_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_646_),
    .C(_610_),
    .Y(_647_)
);

NAND3X1 _1140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_231_),
    .B(_230_),
    .C(_229_),
    .Y(_232_)
);

FILL FILL_1__922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1197_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(ABCmd_i[6]),
    .Y(_693_)
);

FILL FILL_0__944_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_31_),
    .B(_38_),
    .C(_35_),
    .Y(_39_)
);

FILL FILL_1__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1180_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_812_),
    .B(_814_),
    .C(_815_),
    .Y(_816_)
);

OR2X2 _1425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_456_),
    .B(_513_),
    .Y(_515_)
);

INVX1 _1005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .Y(_97_)
);

FILL FILL_1__1587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__960_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1654_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3_),
    .CLK(clk_bF$buf2),
    .Q(alu_op[1])
);

NAND3X1 _1234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_324_),
    .B(_325_),
    .C(_323_),
    .Y(_326_)
);

FILL FILL_0__982_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .Y(_77_)
);

FILL FILL_1__1396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1885_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_850_),
    .Y(_851_)
);

NAND3X1 _1463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_543_),
    .B(_546_),
    .C(_551_),
    .Y(_552_)
);

INVX4 _1043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134_),
    .Y(_135_)
);

FILL FILL_0__1503_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_525_),
    .B(_555_),
    .C(_511_),
    .Y(_607_)
);

INVX2 _1692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[0]),
    .Y(_864_)
);

INVX1 _1272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Flag_i),
    .Y(_364_)
);

FILL FILL_0__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1312_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_917_),
    .B(_916_),
    .C(_912_),
    .Y(_918_)
);

AOI21X1 _1328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .B(_418_),
    .C(_320_),
    .Y(_419_)
);

NAND2X1 _1081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_167_),
    .B(_172_),
    .Y(_173_)
);

FILL FILL_2__1559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_630_),
    .B(_643_),
    .Y(_644_)
);

AOI21X1 _1137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_227_),
    .B(_228_),
    .C(_225_),
    .Y(_229_)
);

FILL FILL_1__1299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1511_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_862_),
    .B(BI[4]),
    .C(_760_),
    .D(_863_),
    .Y(_761_)
);

OAI21X1 _1366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_453_),
    .B(_359_),
    .C(_455_),
    .Y(_456_)
);

FILL FILL_0__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1320_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_678_),
    .B(_679_),
    .C(_668_),
    .D(_675_),
    .Y(_0_[7])
);

NOR2X1 _1175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_265_),
    .B(_266_),
    .Y(_267_)
);

FILL FILL_1__957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86550x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1414_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_860_),
    .Y(_861_)
);

NAND2X1 _1269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_360_),
    .B(_359_),
    .Y(_361_)
);

FILL FILL_0__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1223_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_288_),
    .B(_54_),
    .C(_584_),
    .Y(_586_)
);

NAND3X1 _1078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf2),
    .B(BI[3]),
    .C(AI[4]),
    .Y(_170_)
);

FILL FILL_0__1538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x79350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1291_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(_880_),
    .Y(_882_)
);

FILL FILL_1__1872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1385_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[5]),
    .B(_776_),
    .Y(_777_)
);

FILL FILL_1__1546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1194_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(ABCmd_i[5]),
    .Y(_691_)
);

FILL FILL_0__941_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[1]),
    .Y(_36_)
);

FILL FILL_1__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1004_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op_2_bF$buf2),
    .B(BI[7]),
    .C(_858_),
    .Y(_813_)
);

NAND2X1 _1422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_511_),
    .B(_508_),
    .Y(_512_)
);

NOR2X1 _1002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_92_),
    .B(_93_),
    .Y(_94_)
);

FILL FILL_1__1584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86250x82950 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[7]),
    .B(LoadB_i),
    .Y(_711_)
);

AND2X2 _1231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .B(_306_),
    .Y(_323_)
);

OAI21X1 _982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_716_),
    .B(_44_),
    .C(_72_),
    .Y(_74_)
);

FILL FILL_1__1393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1288_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_874_),
    .B(_876_),
    .C(_878_),
    .Y(_879_)
);

FILL FILL85950x64950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1029_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU8.AI7 ),
    .B(_847_),
    .Y(_848_)
);

OAI21X1 _1460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .B(_501_),
    .C(_548_),
    .Y(_549_)
);

OR2X2 _1040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_131_),
    .B(_130_),
    .Y(_132_)
);

FILL FILL_0__1500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1097_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_603_),
    .Y(_604_)
);

FILL FILL_1__1258_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[2]),
    .B(_914_),
    .Y(_915_)
);

OR2X2 _1325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_314_),
    .B(_315_),
    .Y(_416_)
);

FILL FILL_1__1487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1067_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_633_),
    .Y(_641_)
);

AND2X2 _1134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_718_),
    .B(_714_),
    .Y(_226_)
);

FILL FILL_1__1296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__938_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(shr),
    .B(AI[5]),
    .Y(_758_)
);

NAND2X1 _1363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_352_),
    .B(_451_),
    .Y(_453_)
);

FILL FILL_0__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1174_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_862_),
    .B(BI[7]),
    .C(_809_),
    .D(_863_),
    .Y(_810_)
);

AOI21X1 _1419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_422_),
    .B(_429_),
    .C(_432_),
    .Y(_509_)
);

AOI21X1 _1592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_676_),
    .B(_358_),
    .C(_365_),
    .Y(_677_)
);

OR2X2 _1172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_241_),
    .Y(_264_)
);

FILL FILL_1__954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1212_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadB_i),
    .B(_708_),
    .C(_709_),
    .Y(_23_)
);

OAI21X1 _1228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_153_),
    .B(_154_),
    .C(_157_),
    .Y(_320_)
);

FILL FILL_0__976_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf4),
    .B(BI[4]),
    .C(AI[1]),
    .Y(_71_)
);

FILL FILL_2__1879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1602_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_814_),
    .Y(_845_)
);

NAND3X1 _1457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_535_),
    .B(_545_),
    .C(_544_),
    .Y(_546_)
);

AOI21X1 _1037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_127_),
    .B(_128_),
    .C(_126_),
    .Y(_129_)
);

FILL FILL_1__1199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1411_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX4 _1686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[3]),
    .Y(_858_)
);

OAI21X1 _1266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_280_),
    .B(_356_),
    .C(_357_),
    .Y(_358_)
);

FILL FILL_0__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL85950x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_538_),
    .B(_539_),
    .C(_582_),
    .Y(_583_)
);

INVX1 _1075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_166_),
    .Y(_167_)
);

FILL FILL_0__1535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1314_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_582_),
    .B(_634_),
    .C(_665_),
    .Y(_674_)
);

INVX1 _1169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_248_),
    .Y(_261_)
);

FILL FILL_0__1629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1382_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_766_),
    .Y(_774_)
);

FILL FILL_1__1543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1123_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .B(_486_),
    .C(_413_),
    .Y(_488_)
);

FILL FILL_0__1858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1191_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(ABCmd_i[4]),
    .Y(_689_)
);

NAND3X1 _941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf4),
    .B(BI[1]),
    .C(AI[3]),
    .Y(_33_)
);

FILL FILL_1__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1285_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .B(alu_op_2_bF$buf1),
    .C(_875_),
    .Y(_876_)
);

FILL FILL_1__1866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1094_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_577_),
    .B(_600_),
    .Y(_601_)
);

FILL FILL_1__1255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1324_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(shr),
    .B(AI[3]),
    .Y(_912_)
);

NAND3X1 _1322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(_412_),
    .C(_411_),
    .Y(_413_)
);

FILL FILL_1__1484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1379_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .B(_587_),
    .C(_636_),
    .Y(_638_)
);

OAI21X1 _1131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_34_),
    .B(_40_),
    .C(_31_),
    .Y(_223_)
);

FILL FILL_1__1293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1188_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(ABCmd_i[3]),
    .Y(_687_)
);

FILL FILL_0__935_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf4),
    .B(BI[2]),
    .C(AI[2]),
    .Y(_30_)
);

FILL FILL_1__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1349_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_732_),
    .B(_731_),
    .Y(_755_)
);

AND2X2 _1360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_442_),
    .B(_447_),
    .Y(_451_)
);

FILL FILL_0__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1400_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(shr),
    .B(CI),
    .Y(_807_)
);

NAND3X1 _1416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_457_),
    .B(_504_),
    .C(_505_),
    .Y(_506_)
);

FILL FILL_1__1578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL85950x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadB_i),
    .B(_169_),
    .C(_707_),
    .Y(_22_)
);

AND2X2 _1225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_314_),
    .B(_315_),
    .Y(_317_)
);

FILL FILL_0__973_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_67_),
    .Y(_68_)
);

FILL FILL_1__1387_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_790_),
    .B(_801_),
    .C(_805_),
    .Y(_842_)
);

OAI21X1 _1454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_537_),
    .B(_536_),
    .C(_542_),
    .Y(_543_)
);

AOI21X1 _1034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_79_),
    .B(_66_),
    .C(_81_),
    .Y(_126_)
);

FILL FILL_1__1196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1265_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1683_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_24_),
    .CLK(clk_bF$buf1),
    .Q(BI[6])
);

INVX1 _1263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .Y(_355_)
);

FILL FILL_0__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1494_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_909_),
    .Y(ACC[1])
);

NAND3X1 _1319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_396_),
    .B(_404_),
    .C(_406_),
    .Y(_410_)
);

INVX1 _1492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_579_),
    .Y(_580_)
);

OAI21X1 _1072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_152_),
    .B(_153_),
    .C(_154_),
    .Y(_164_)
);

FILL FILL_0__1532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1112_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_288_),
    .B(_158_),
    .C(_417_),
    .D(_135_),
    .Y(_635_)
);

NOR2X1 _1128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_714_),
    .B(_718_),
    .Y(_220_)
);

FILL FILL_0__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1502_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BCD),
    .Y(_752_)
);

NAND2X1 _1357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_447_),
    .B(_442_),
    .Y(_448_)
);

FILL FILL_1__1099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1311_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_671_),
    .B(_666_),
    .C(_670_),
    .Y(_672_)
);

NAND3X1 _1166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_139_),
    .B(_142_),
    .C(_257_),
    .Y(_258_)
);

FILL FILL_1__948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86550x43350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1120_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf0)
);

OAI21X1 _1395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_483_),
    .B(_484_),
    .C(_475_),
    .Y(_485_)
);

FILL FILL_0__1855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1214_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_576_),
    .Y(_577_)
);

NAND3X1 _1069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_149_),
    .B(_156_),
    .C(_160_),
    .Y(_161_)
);

FILL FILL_0__1529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1282_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[1]),
    .B(shr),
    .Y(_873_)
);

FILL FILL_1__1863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1023_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_387_),
    .B(_135_),
    .C(_388_),
    .Y(_389_)
);

FILL FILL_0__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1091_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_546_),
    .B(_593_),
    .Y(_598_)
);

FILL FILL_1__1252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1185_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCmd_i),
    .B(ABCmd_i[2]),
    .Y(_685_)
);

FILL FILL_0__932_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_725_),
    .B(_26_),
    .C(_720_),
    .Y(_27_)
);

FILL FILL_1__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86850x18150 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_804_),
    .Y(ACC[6])
);

NAND3X1 _1413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_458_),
    .B(_502_),
    .C(_494_),
    .Y(_503_)
);

FILL FILL_1__1575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__999_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABCmd_i[3]),
    .B(LoadB_i),
    .Y(_706_)
);

NAND3X1 _1222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MUL_bF$buf2),
    .B(AI[6]),
    .C(BI[2]),
    .Y(_314_)
);

FILL FILL_0__970_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_55_),
    .B(_56_),
    .C(_52_),
    .Y(_65_)
);

FILL FILL_1__1384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1279_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_804_),
    .B(_789_),
    .C(_752_),
    .Y(_839_)
);

OR2X2 _1451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_538_),
    .B(_539_),
    .Y(_540_)
);

AND2X2 _1031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114_),
    .B(_118_),
    .Y(_123_)
);

FILL FILL_1__1193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1088_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_593_),
    .B(_546_),
    .Y(_595_)
);

FILL FILL_1__1249_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1680_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_21_),
    .CLK(clk_bF$buf0),
    .Q(BI[3])
);

AND2X2 _1260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_347_),
    .B(_351_),
    .Y(_352_)
);

FILL FILL_0__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1300_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_891_),
    .B(_893_),
    .C(_906_),
    .Y(_907_)
);

AOI21X1 _1316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_404_),
    .B(_406_),
    .C(_396_),
    .Y(_407_)
);

FILL FILL_1__1478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1058_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .B(_540_),
    .Y(_632_)
);

OAI21X1 _1125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_215_),
    .B(_216_),
    .C(_132_),
    .Y(_217_)
);

FILL FILL_1__1287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__929_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_732_),
    .B(_747_),
    .C(_731_),
    .Y(_750_)
);

NAND3X1 _1354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_378_),
    .B(_439_),
    .C(_440_),
    .Y(_445_)
);

FILL FILL_1__1096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1585_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_646_),
    .B(_603_),
    .Y(_669_)
);

NAND3X1 _1163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_233_),
    .B(_252_),
    .C(_254_),
    .Y(_255_)
);

FILL FILL_1__945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1203_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadB_i),
    .B(_36_),
    .C(_704_),
    .Y(_19_)
);

NAND3X1 _1219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_307_),
    .B(_310_),
    .C(_308_),
    .Y(_311_)
);

FILL FILL_0__967_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_476_),
    .B(_481_),
    .C(_479_),
    .Y(_482_)
);

FILL FILL_0__1852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL86550x64950 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_828_),
    .B(_835_),
    .C(_836_),
    .Y(_837_)
);

AOI21X1 _1448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_532_),
    .B(_534_),
    .C(_530_),
    .Y(_537_)
);

NAND3X1 _1028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_102_),
    .B(_119_),
    .C(_106_),
    .Y(_120_)
);

FILL FILL_1__983_ (
    .gnd(gnd),
    .vdd(vdd)
);

endmodule
