#--------------------------------------------------
# LEF file for Route & Via Rile
#  Ported from osu050 by GoodKook@gmail.com
#

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

USEMINSPACING OBS ON ;
USEMINSPACING PIN OFF ;
CLEARANCEMEASURE EUCLIDEAN ;

MANUFACTURINGGRID 0.15 ;

LAYER nwell
  TYPE	MASTERSLICE ;
END nwell

LAYER nactive
  TYPE	MASTERSLICE ;
END nactive

LAYER pactive
  TYPE	MASTERSLICE ;
END pactive

LAYER poly
  TYPE	MASTERSLICE ;
END poly

LAYER cc
  TYPE	CUT ;
  SPACING	0.6 ;
END cc

LAYER metal1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		3.0 ;
  OFFSET	1.5 ;
  WIDTH	    0.9 ;   # ETRI050 Rule: WIDTH=0.8
  SPACING	0.9 ;   # ETRI050 Rule: SPACING=0.8(1.0 for Width >10um)
  RESISTANCE	RPERSQ 0.09 ;
  CAPACITANCE	CPERSQDIST 3.2e-05 ;
END metal1

LAYER via1
  TYPE	CUT ;
  SPACING	0.9 ;
END via1

LAYER metal2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		3.0 ;
  OFFSET	1.5 ;
  WIDTH		1.05 ;  # ETRI050 Rule: WIDTH=1.0
  SPACING	0.9 ;   # ETRI050 Rule: SPACING=1.0(1.2 for Width >10um)
  RESISTANCE	RPERSQ 0.09 ;
  CAPACITANCE	CPERSQDIST 1.6e-05 ;
END metal2

LAYER via2
  TYPE	CUT ;
  SPACING	0.9 ;
END via2

LAYER metal3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		3.0 ;
  OFFSET	1.5 ;
  WIDTH		1.2 ;   # ETRI050 Rule: WIDTH=1.2
  SPACING	0.9 ;   # ETRI050 Rule: SPACING=1.0(1.2 for Width >10um)
  RESISTANCE	RPERSQ 0.05 ;
  CAPACITANCE	CPERSQDIST 1e-05 ;
END metal3

SPACING
  SAMENET cc   via1	0.900 ;
  SAMENET via1 via2	0.900 ;
END SPACING

VIA M2_M1 DEFAULT
  LAYER metal1 ;
    RECT -1.050 -1.050 1.050 1.050 ;
  LAYER via1 ;
    RECT -0.450 -0.450 0.450 0.450 ;
  LAYER metal2 ;
    RECT -1.050 -1.050 1.050 1.050 ;
END M2_M1

VIA M3_M2 DEFAULT
  LAYER metal2 ;
    RECT -1.050 -1.050 1.050 1.050 ;
  LAYER via2 ;
    RECT -0.450 -0.450 0.450 0.450 ;
  LAYER metal3 ;
    RECT -1.050 -1.050 1.050 1.050 ;
END M3_M2


VIARULE viagen21 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER via1 ;
#    RECT -1.05 -1.05 1.05 1.05 ;
    RECT -0.450 -0.450 0.450 0.450 ;
    SPACING 0.9 BY 0.9 ;
END viagen21

VIARULE viagen32 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER via2 ;
#    RECT -1.05 -1.05 1.05 1.05 ;
    RECT -0.450 -0.450 0.450 0.450 ;
    SPACING 0.9 BY 0.9 ;
END viagen32

VIARULE TURN1 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
  LAYER metal1 ;
    DIRECTION VERTICAL ;
END TURN1

VIARULE TURN2 GENERATE
  LAYER metal2 ;
    DIRECTION HORIZONTAL ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
END TURN2

VIARULE TURN3 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
  LAYER metal3 ;
    DIRECTION VERTICAL ;
END TURN3

SITE  corner
    CLASS	PAD ;
    SYMMETRY	R90 Y ;
    SIZE	300.000 BY 300.000 ;
END  corner

SITE  IO
    CLASS	PAD ;
    SYMMETRY	Y ;
    SIZE	90.000 BY 300.000 ;
END  IO

SITE  core
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	3.000 BY 30.000 ;
END  core

# =====================================================================
#  Core MACROS
# =====================================================================
MACRO AND2X1
  CLASS CORE ;
  FOREIGN AND2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 15.450 2.550 17.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.450 12.450 11.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 15.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 27.900 2.850 33.750 ;
        RECT 4.050 27.900 5.850 33.750 ;
        RECT 7.050 27.900 8.850 33.750 ;
        RECT 10.050 27.900 11.850 33.750 ;
        RECT 0.450 13.350 2.550 15.450 ;
        RECT 0.600 11.550 2.400 13.350 ;
        RECT 4.200 10.350 5.250 27.900 ;
        RECT 6.450 16.350 8.550 18.450 ;
        RECT 10.200 16.650 11.250 27.900 ;
        RECT 6.600 14.550 8.400 16.350 ;
        RECT 9.450 14.550 11.550 16.650 ;
        RECT 6.750 10.350 8.550 10.800 ;
        RECT 1.050 9.000 8.550 10.350 ;
        RECT 1.050 2.250 2.850 9.000 ;
        RECT 5.250 2.250 7.050 8.100 ;
        RECT 10.200 6.300 11.250 14.550 ;
        RECT 8.550 5.100 11.250 6.300 ;
        RECT 8.550 2.250 10.350 5.100 ;
      LAYER metal2 ;
        RECT 6.450 16.350 8.550 17.250 ;
        RECT 9.450 15.750 11.550 16.650 ;
        RECT 0.450 13.350 2.550 14.250 ;
  END
END AND2X1
MACRO AND2X2
  CLASS CORE ;
  FOREIGN AND2X2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 12.450 2.550 14.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.450 12.450 11.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 15.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 27.900 2.850 33.750 ;
        RECT 4.050 27.900 5.850 33.750 ;
        RECT 0.600 16.650 2.400 18.450 ;
        RECT 0.450 14.550 2.550 16.650 ;
        RECT 4.200 10.800 5.400 27.900 ;
        RECT 7.650 21.900 9.450 33.750 ;
        RECT 10.650 21.900 12.450 33.750 ;
        RECT 6.450 16.350 8.550 18.450 ;
        RECT 10.650 16.650 11.850 21.900 ;
        RECT 6.600 14.550 8.400 16.350 ;
        RECT 9.450 14.550 11.850 16.650 ;
        RECT 1.050 9.600 8.550 10.800 ;
        RECT 1.050 2.250 2.850 9.600 ;
        RECT 6.750 9.000 8.550 9.600 ;
        RECT 10.650 8.100 11.850 14.550 ;
        RECT 5.550 2.250 7.350 8.100 ;
        RECT 8.550 6.600 11.850 8.100 ;
        RECT 8.550 2.250 10.350 6.600 ;
      LAYER metal2 ;
        RECT 0.450 15.750 2.550 16.650 ;
        RECT 6.450 16.350 8.550 17.250 ;
        RECT 9.450 15.750 11.550 16.650 ;
  END
END AND2X2
MACRO AOI21X1
  CLASS CORE ;
  FOREIGN AOI21X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 15.450 2.550 17.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 9.450 5.550 11.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.450 15.450 8.550 17.550 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.450 12.450 11.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 15.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 22.800 2.850 33.750 ;
        RECT 4.050 23.700 5.850 33.750 ;
        RECT 7.050 22.800 8.850 33.750 ;
        RECT 1.050 21.900 8.850 22.800 ;
        RECT 10.050 21.900 11.850 33.750 ;
        RECT 10.200 16.650 11.400 21.900 ;
        RECT 0.450 13.350 2.550 15.450 ;
        RECT 3.600 13.650 5.400 15.450 ;
        RECT 0.600 11.550 2.400 13.350 ;
        RECT 3.450 11.550 5.550 13.650 ;
        RECT 6.450 13.350 8.550 15.450 ;
        RECT 9.450 14.550 11.550 16.650 ;
        RECT 6.600 11.550 8.400 13.350 ;
        RECT 10.200 8.100 11.400 14.550 ;
        RECT 1.500 2.250 3.300 8.100 ;
        RECT 5.700 6.450 11.400 8.100 ;
        RECT 5.700 2.250 7.500 6.450 ;
        RECT 9.000 2.250 10.800 5.100 ;
      LAYER metal2 ;
        RECT 9.750 15.750 11.550 16.650 ;
        RECT 0.450 13.350 2.550 14.250 ;
        RECT 3.450 12.750 5.550 13.650 ;
        RECT 6.450 13.350 8.250 14.250 ;
  END
END AOI21X1
MACRO AOI22X1
  CLASS CORE ;
  FOREIGN AOI22X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 12.450 2.550 14.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 12.450 12.450 14.550 14.550 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.450 12.450 8.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 18.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 18.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 23.100 2.850 33.750 ;
        RECT 4.050 24.000 5.850 33.750 ;
        RECT 7.050 33.000 14.850 33.750 ;
        RECT 7.050 23.100 8.850 33.000 ;
        RECT 1.050 22.200 8.850 23.100 ;
        RECT 10.050 21.900 11.850 32.100 ;
        RECT 13.050 21.900 14.850 33.000 ;
        RECT 9.900 21.000 11.700 21.900 ;
        RECT 7.650 20.100 11.700 21.000 ;
        RECT 0.750 16.650 2.550 18.450 ;
        RECT 7.650 16.650 8.550 20.100 ;
        RECT 12.600 16.650 14.400 18.450 ;
        RECT 0.450 14.550 2.550 16.650 ;
        RECT 3.450 13.350 5.550 15.450 ;
        RECT 3.750 11.550 5.550 13.350 ;
        RECT 6.450 14.550 8.550 16.650 ;
        RECT 6.450 8.100 7.500 14.550 ;
        RECT 9.450 13.350 11.550 15.450 ;
        RECT 12.450 14.550 14.550 16.650 ;
        RECT 9.450 11.550 11.250 13.350 ;
        RECT 1.500 2.250 3.300 8.100 ;
        RECT 5.700 2.250 7.500 8.100 ;
        RECT 9.900 2.250 11.700 8.100 ;
      LAYER metal2 ;
        RECT 0.450 15.750 2.250 16.650 ;
        RECT 6.750 15.750 8.250 16.650 ;
        RECT 12.750 15.750 14.550 16.650 ;
        RECT 3.750 13.350 5.250 14.250 ;
        RECT 9.750 13.350 11.250 14.250 ;
  END
END AOI22X1
MACRO BUFX2
  CLASS CORE ;
  FOREIGN BUFX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 12.450 2.550 14.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.450 12.450 8.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 12.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 12.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 27.900 2.850 33.750 ;
        RECT 1.050 21.000 2.250 27.900 ;
        RECT 4.350 21.900 6.150 33.750 ;
        RECT 7.350 21.900 9.150 33.750 ;
        RECT 1.050 20.100 6.750 21.000 ;
        RECT 4.500 19.200 6.750 20.100 ;
        RECT 0.600 16.650 2.400 18.450 ;
        RECT 0.450 14.550 2.550 16.650 ;
        RECT 4.500 10.800 5.550 19.200 ;
        RECT 7.650 16.650 8.850 21.900 ;
        RECT 6.450 14.550 8.850 16.650 ;
        RECT 4.500 9.900 6.750 10.800 ;
        RECT 1.650 9.000 6.750 9.900 ;
        RECT 1.650 5.100 2.850 9.000 ;
        RECT 7.650 8.100 8.850 14.550 ;
        RECT 1.050 2.250 2.850 5.100 ;
        RECT 4.350 2.250 6.150 8.100 ;
        RECT 7.350 2.250 9.150 8.100 ;
      LAYER metal2 ;
        RECT 0.450 15.750 2.550 16.650 ;
        RECT 6.450 15.750 8.550 16.650 ;
  END
END BUFX2
MACRO BUFX4
  CLASS CORE ;
  FOREIGN BUFX4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 12.450 2.550 14.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.450 12.450 11.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 16.050 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 16.200 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 21.000 2.850 33.750 ;
        RECT 4.350 21.900 6.150 33.750 ;
        RECT 7.350 21.900 9.150 33.750 ;
        RECT 10.350 21.900 12.150 33.750 ;
        RECT 1.050 20.100 6.900 21.000 ;
        RECT 5.100 19.200 6.900 20.100 ;
        RECT 0.600 16.650 2.400 18.450 ;
        RECT 0.450 14.550 2.550 16.650 ;
        RECT 5.100 10.800 6.300 19.200 ;
        RECT 7.800 16.650 8.850 21.900 ;
        RECT 7.800 14.550 11.550 16.650 ;
        RECT 5.100 9.900 6.900 10.800 ;
        RECT 1.050 9.000 6.900 9.900 ;
        RECT 1.050 6.600 2.250 9.000 ;
        RECT 7.800 8.100 8.850 14.550 ;
        RECT 1.050 2.250 2.850 6.600 ;
        RECT 4.350 2.250 6.150 8.100 ;
        RECT 7.350 2.250 9.150 8.100 ;
        RECT 10.350 2.250 12.150 8.100 ;
      LAYER metal2 ;
        RECT 0.450 15.750 2.550 16.650 ;
        RECT 9.450 15.750 11.550 16.650 ;
  END
END BUFX4
MACRO CLKBUF1
  CLASS CORE ;
  FOREIGN CLKBUF1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 24.450 15.450 26.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 30.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 30.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 21.900 2.850 33.750 ;
        RECT 4.050 21.000 5.850 33.750 ;
        RECT 7.050 21.900 8.850 33.750 ;
        RECT 10.050 21.000 11.850 33.750 ;
        RECT 13.050 21.900 14.850 33.750 ;
        RECT 16.050 21.000 17.850 33.750 ;
        RECT 19.050 21.900 20.850 33.750 ;
        RECT 22.050 21.000 23.850 33.750 ;
        RECT 25.050 21.900 26.850 33.750 ;
        RECT 4.050 19.800 7.950 21.000 ;
        RECT 10.050 19.800 13.800 21.000 ;
        RECT 16.050 19.800 19.800 21.000 ;
        RECT 22.050 19.800 24.750 21.000 ;
        RECT 3.450 13.350 5.550 15.450 ;
        RECT 3.600 11.550 5.400 13.350 ;
        RECT 6.750 12.900 7.950 19.800 ;
        RECT 12.600 12.900 13.800 19.800 ;
        RECT 18.600 12.900 19.800 19.800 ;
        RECT 23.700 15.450 24.750 19.800 ;
        RECT 23.700 13.350 26.550 15.450 ;
        RECT 6.750 11.100 10.800 12.900 ;
        RECT 12.600 11.100 16.800 12.900 ;
        RECT 18.600 11.100 22.800 12.900 ;
        RECT 6.750 10.200 7.950 11.100 ;
        RECT 12.600 10.200 13.800 11.100 ;
        RECT 18.600 10.200 19.800 11.100 ;
        RECT 23.700 10.200 24.750 13.350 ;
        RECT 3.900 9.000 7.950 10.200 ;
        RECT 10.050 9.000 13.800 10.200 ;
        RECT 15.900 9.000 19.800 10.200 ;
        RECT 21.900 9.150 24.750 10.200 ;
        RECT 21.900 9.000 24.600 9.150 ;
        RECT 3.900 8.100 5.700 9.000 ;
        RECT 1.050 2.250 2.850 8.100 ;
        RECT 4.050 2.250 5.850 8.100 ;
        RECT 7.050 2.250 8.850 8.100 ;
        RECT 10.050 2.250 11.850 9.000 ;
        RECT 15.900 8.100 17.700 9.000 ;
        RECT 21.900 8.100 23.700 9.000 ;
        RECT 13.050 2.250 14.850 8.100 ;
        RECT 16.050 2.250 17.850 8.100 ;
        RECT 19.050 2.250 20.850 8.100 ;
        RECT 22.050 2.250 23.850 8.100 ;
        RECT 25.050 2.250 26.850 8.100 ;
      LAYER metal2 ;
        RECT 3.450 13.350 5.550 14.250 ;
        RECT 24.450 13.350 26.550 14.250 ;
  END
END CLKBUF1
MACRO CLKBUF2
  CLASS CORE ;
  FOREIGN CLKBUF2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 42.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 36.450 15.450 38.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 42.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 42.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 21.900 2.850 33.750 ;
        RECT 4.050 21.900 5.850 33.750 ;
        RECT 7.050 21.900 8.850 33.750 ;
        RECT 10.050 21.900 11.850 33.750 ;
        RECT 13.050 21.900 14.850 33.750 ;
        RECT 3.900 21.000 5.700 21.900 ;
        RECT 9.900 21.000 11.700 21.900 ;
        RECT 16.050 21.000 17.850 33.750 ;
        RECT 19.050 21.900 20.850 33.750 ;
        RECT 22.050 21.900 23.850 33.750 ;
        RECT 25.050 21.900 26.850 33.750 ;
        RECT 21.900 21.000 23.700 21.900 ;
        RECT 28.050 21.000 29.850 33.750 ;
        RECT 31.050 21.900 32.850 33.750 ;
        RECT 34.050 21.900 35.850 33.750 ;
        RECT 37.050 21.900 38.850 33.750 ;
        RECT 33.900 21.000 35.700 21.900 ;
        RECT 3.900 19.800 7.950 21.000 ;
        RECT 9.900 19.800 13.800 21.000 ;
        RECT 16.050 19.800 19.800 21.000 ;
        RECT 21.900 19.800 26.100 21.000 ;
        RECT 28.050 19.800 31.200 21.000 ;
        RECT 33.900 19.800 37.200 21.000 ;
        RECT 3.450 13.350 5.550 15.450 ;
        RECT 3.600 11.550 5.400 13.350 ;
        RECT 6.750 12.900 7.950 19.800 ;
        RECT 12.600 12.900 13.800 19.800 ;
        RECT 18.600 12.900 19.800 19.800 ;
        RECT 24.900 12.900 26.100 19.800 ;
        RECT 30.000 12.900 31.200 19.800 ;
        RECT 36.000 15.450 37.200 19.800 ;
        RECT 36.000 13.350 38.550 15.450 ;
        RECT 6.750 11.100 10.800 12.900 ;
        RECT 12.600 11.100 16.800 12.900 ;
        RECT 18.600 11.100 22.800 12.900 ;
        RECT 24.900 11.100 28.800 12.900 ;
        RECT 30.000 11.100 34.800 12.900 ;
        RECT 6.750 10.200 7.950 11.100 ;
        RECT 12.600 10.200 13.800 11.100 ;
        RECT 18.600 10.200 19.800 11.100 ;
        RECT 24.900 10.200 26.100 11.100 ;
        RECT 30.000 10.200 31.200 11.100 ;
        RECT 36.000 10.200 37.200 13.350 ;
        RECT 4.050 9.000 7.950 10.200 ;
        RECT 10.050 9.000 13.800 10.200 ;
        RECT 16.050 9.000 19.800 10.200 ;
        RECT 21.900 9.000 26.100 10.200 ;
        RECT 28.050 9.000 31.200 10.200 ;
        RECT 34.050 9.000 37.200 10.200 ;
        RECT 1.050 2.250 2.850 8.100 ;
        RECT 4.050 2.250 5.850 9.000 ;
        RECT 7.050 2.250 8.850 8.100 ;
        RECT 10.050 2.250 11.850 9.000 ;
        RECT 13.050 2.250 14.850 8.100 ;
        RECT 16.050 2.250 17.850 9.000 ;
        RECT 21.900 8.100 23.700 9.000 ;
        RECT 19.050 2.250 20.850 8.100 ;
        RECT 22.050 2.250 23.850 8.100 ;
        RECT 25.050 2.250 26.850 8.100 ;
        RECT 28.050 2.250 29.850 9.000 ;
        RECT 31.050 2.250 32.850 8.100 ;
        RECT 34.050 2.250 35.850 9.000 ;
        RECT 37.050 2.250 38.850 8.100 ;
      LAYER metal2 ;
        RECT 3.450 13.350 5.550 14.250 ;
        RECT 36.450 13.350 38.550 14.250 ;
  END
END CLKBUF2
MACRO CLKBUF3
  CLASS CORE ;
  FOREIGN CLKBUF3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 54.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 48.450 15.450 50.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 54.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 55.200 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 21.900 2.850 33.750 ;
        RECT 4.050 21.000 5.850 33.750 ;
        RECT 7.050 21.900 8.850 33.750 ;
        RECT 10.050 21.000 11.850 33.750 ;
        RECT 13.050 21.900 14.850 33.750 ;
        RECT 16.050 21.000 17.850 33.750 ;
        RECT 19.050 21.900 20.850 33.750 ;
        RECT 22.050 21.000 23.850 33.750 ;
        RECT 25.050 21.900 26.850 33.750 ;
        RECT 28.050 21.000 29.850 33.750 ;
        RECT 31.050 21.900 32.850 33.750 ;
        RECT 34.050 21.000 35.850 33.750 ;
        RECT 37.050 21.900 38.850 33.750 ;
        RECT 40.050 21.000 41.850 33.750 ;
        RECT 43.050 21.900 44.850 33.750 ;
        RECT 46.050 21.000 47.850 33.750 ;
        RECT 49.050 21.900 50.850 33.750 ;
        RECT 4.050 19.800 7.800 21.000 ;
        RECT 10.050 19.800 13.800 21.000 ;
        RECT 16.050 19.800 19.800 21.000 ;
        RECT 22.050 19.800 26.100 21.000 ;
        RECT 28.050 19.800 31.200 21.000 ;
        RECT 34.050 19.800 37.800 21.000 ;
        RECT 40.050 19.800 42.900 21.000 ;
        RECT 46.050 19.800 49.050 21.000 ;
        RECT 3.450 13.350 5.550 15.450 ;
        RECT 3.600 11.550 5.400 13.350 ;
        RECT 6.750 12.900 7.800 19.800 ;
        RECT 12.600 12.900 13.800 19.800 ;
        RECT 18.600 12.900 19.800 19.800 ;
        RECT 24.900 12.900 26.100 19.800 ;
        RECT 30.000 12.900 31.200 19.800 ;
        RECT 36.600 12.900 37.800 19.800 ;
        RECT 41.700 12.900 42.900 19.800 ;
        RECT 47.850 15.450 49.050 19.800 ;
        RECT 47.850 13.350 50.550 15.450 ;
        RECT 6.750 11.100 10.800 12.900 ;
        RECT 12.600 11.100 16.800 12.900 ;
        RECT 18.600 11.100 22.800 12.900 ;
        RECT 24.900 11.100 28.800 12.900 ;
        RECT 30.000 11.100 34.800 12.900 ;
        RECT 36.600 11.100 40.800 12.900 ;
        RECT 41.700 11.100 46.800 12.900 ;
        RECT 6.750 10.200 7.800 11.100 ;
        RECT 12.600 10.200 13.800 11.100 ;
        RECT 18.600 10.200 19.800 11.100 ;
        RECT 24.900 10.200 26.100 11.100 ;
        RECT 30.000 10.200 31.200 11.100 ;
        RECT 36.600 10.200 37.800 11.100 ;
        RECT 41.700 10.200 42.900 11.100 ;
        RECT 47.850 10.200 49.050 13.350 ;
        RECT 4.050 9.000 7.800 10.200 ;
        RECT 10.050 9.000 13.800 10.200 ;
        RECT 16.050 9.000 19.800 10.200 ;
        RECT 22.050 9.000 26.100 10.200 ;
        RECT 28.050 9.000 31.200 10.200 ;
        RECT 34.050 9.000 37.800 10.200 ;
        RECT 40.050 9.000 42.900 10.200 ;
        RECT 45.900 9.000 49.050 10.200 ;
        RECT 1.050 2.250 2.850 8.100 ;
        RECT 4.050 2.250 5.850 9.000 ;
        RECT 7.050 2.250 8.850 8.100 ;
        RECT 10.050 2.250 11.850 9.000 ;
        RECT 13.050 2.250 14.850 8.100 ;
        RECT 16.050 2.250 17.850 9.000 ;
        RECT 19.050 2.250 20.850 8.100 ;
        RECT 22.050 2.250 23.850 9.000 ;
        RECT 25.050 2.250 26.850 8.100 ;
        RECT 28.050 2.250 29.850 9.000 ;
        RECT 31.050 2.250 32.850 8.100 ;
        RECT 34.050 2.250 35.850 9.000 ;
        RECT 37.050 2.250 38.850 8.100 ;
        RECT 40.050 2.250 41.850 9.000 ;
        RECT 45.900 8.100 47.700 9.000 ;
        RECT 43.050 2.250 44.850 8.100 ;
        RECT 46.050 2.250 47.850 8.100 ;
        RECT 49.050 2.250 50.850 8.100 ;
      LAYER metal2 ;
        RECT 3.450 13.350 5.550 14.250 ;
        RECT 48.450 13.350 50.550 14.250 ;
  END
END CLKBUF3
MACRO DFFNEGX1
  CLASS CORE ;
  FOREIGN DFFNEGX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 12.450 5.550 14.550 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal2 ;
        RECT 15.450 12.450 17.550 14.550 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 30.450 12.450 32.550 14.550 ;
    END
  END Q
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 36.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 36.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 21.300 2.850 33.750 ;
        RECT 4.050 27.900 5.850 33.750 ;
        RECT 8.850 29.550 10.650 33.750 ;
        RECT 7.050 27.900 10.650 29.550 ;
        RECT 13.650 27.900 15.450 33.750 ;
        RECT 7.050 27.300 8.700 27.900 ;
        RECT 6.600 25.200 8.700 27.300 ;
        RECT 16.650 27.000 18.450 33.750 ;
        RECT 20.400 27.900 22.200 33.750 ;
        RECT 24.750 27.900 26.550 33.750 ;
        RECT 29.250 30.900 31.050 33.750 ;
        RECT 9.750 24.300 11.550 27.000 ;
        RECT 12.750 25.200 19.350 27.000 ;
        RECT 24.450 25.800 26.550 27.900 ;
        RECT 9.600 22.200 11.700 24.300 ;
        RECT 20.250 22.200 27.150 24.000 ;
        RECT 20.250 21.300 21.150 22.200 ;
        RECT 1.050 20.100 21.150 21.300 ;
        RECT 32.250 21.900 34.050 33.750 ;
        RECT 1.050 8.100 1.950 20.100 ;
        RECT 7.950 19.500 9.750 20.100 ;
        RECT 14.550 18.600 16.350 19.200 ;
        RECT 3.600 16.650 5.400 18.450 ;
        RECT 6.600 17.400 16.350 18.600 ;
        RECT 24.450 18.000 26.550 18.600 ;
        RECT 29.550 18.000 31.350 18.600 ;
        RECT 3.450 14.550 5.550 16.650 ;
        RECT 6.600 16.500 8.700 17.400 ;
        RECT 24.450 16.800 31.350 18.000 ;
        RECT 24.450 16.500 26.550 16.800 ;
        RECT 9.600 11.400 11.700 13.200 ;
        RECT 32.250 12.450 33.450 21.900 ;
        RECT 15.450 11.400 17.550 12.450 ;
        RECT 30.450 12.150 33.450 12.450 ;
        RECT 3.000 10.200 23.850 11.400 ;
        RECT 27.150 10.350 33.450 12.150 ;
        RECT 3.000 9.600 4.800 10.200 ;
        RECT 7.950 9.000 9.750 10.200 ;
        RECT 22.050 8.700 23.850 10.200 ;
        RECT 32.250 8.100 33.450 10.350 ;
        RECT 1.050 2.250 2.850 8.100 ;
        RECT 6.600 6.000 8.700 8.100 ;
        RECT 12.750 7.200 14.550 7.800 ;
        RECT 12.750 6.000 17.850 7.200 ;
        RECT 7.050 5.100 8.700 6.000 ;
        RECT 16.650 5.100 17.850 6.000 ;
        RECT 4.050 2.250 5.850 5.100 ;
        RECT 7.050 4.050 10.650 5.100 ;
        RECT 8.850 2.250 10.650 4.050 ;
        RECT 13.350 2.250 15.150 5.100 ;
        RECT 16.650 2.250 18.450 5.100 ;
        RECT 20.250 2.250 22.050 5.100 ;
        RECT 24.450 4.200 26.550 7.200 ;
        RECT 24.750 2.250 26.550 4.200 ;
        RECT 29.250 2.250 31.050 5.100 ;
        RECT 32.250 2.250 34.050 8.100 ;
      LAYER metal2 ;
        RECT 6.600 25.200 8.700 27.300 ;
        RECT 24.450 25.800 26.550 27.900 ;
        RECT 7.200 18.600 8.250 25.200 ;
        RECT 9.600 22.200 11.700 24.300 ;
        RECT 3.450 15.750 5.550 16.650 ;
        RECT 6.600 16.500 8.700 18.600 ;
        RECT 7.200 8.100 8.250 16.500 ;
        RECT 10.200 13.200 11.400 22.200 ;
        RECT 24.900 18.600 26.100 25.800 ;
        RECT 24.450 16.500 26.550 18.600 ;
        RECT 9.600 11.100 11.700 13.200 ;
        RECT 15.450 10.350 17.550 11.250 ;
        RECT 6.600 6.000 8.700 8.100 ;
        RECT 24.900 7.200 26.100 16.500 ;
        RECT 30.450 10.350 32.550 11.250 ;
        RECT 24.450 5.100 26.550 7.200 ;
  END
END DFFNEGX1
MACRO DFFPOSX1
  CLASS CORE ;
  FOREIGN DFFPOSX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 12.450 12.450 14.550 14.550 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal2 ;
        RECT 18.450 12.450 20.550 14.550 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 30.450 12.450 32.550 14.550 ;
    END
  END Q
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 36.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 36.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.650 21.900 3.450 33.750 ;
        RECT 4.650 27.900 6.450 33.750 ;
        RECT 9.750 27.900 11.550 33.750 ;
        RECT 14.550 27.900 16.350 33.750 ;
        RECT 10.050 27.000 11.250 27.900 ;
        RECT 17.550 27.000 19.350 33.750 ;
        RECT 21.450 27.900 23.250 33.750 ;
        RECT 25.650 27.900 27.450 33.750 ;
        RECT 30.150 30.900 31.950 33.750 ;
        RECT 6.450 24.900 11.250 27.000 ;
        RECT 13.650 25.200 20.550 27.000 ;
        RECT 25.650 25.800 29.550 27.900 ;
        RECT 10.050 24.000 11.250 24.900 ;
        RECT 22.950 24.300 24.750 24.900 ;
        RECT 10.050 22.800 17.550 24.000 ;
        RECT 15.750 22.200 17.550 22.800 ;
        RECT 18.450 23.400 24.750 24.300 ;
        RECT 1.650 21.300 12.750 21.900 ;
        RECT 18.450 21.300 19.350 23.400 ;
        RECT 22.950 23.100 24.750 23.400 ;
        RECT 25.650 23.100 28.350 24.900 ;
        RECT 25.650 22.200 26.550 23.100 ;
        RECT 1.650 20.700 19.350 21.300 ;
        RECT 1.650 8.100 2.550 20.700 ;
        RECT 10.950 20.400 19.350 20.700 ;
        RECT 20.550 21.300 26.550 22.200 ;
        RECT 27.450 21.300 29.550 22.200 ;
        RECT 33.150 21.900 34.950 33.750 ;
        RECT 10.950 20.100 12.750 20.400 ;
        RECT 20.550 16.650 21.450 21.300 ;
        RECT 27.450 20.100 31.650 21.300 ;
        RECT 30.750 18.300 32.550 20.100 ;
        RECT 12.450 15.600 14.550 16.650 ;
        RECT 3.600 13.650 5.400 15.450 ;
        RECT 6.600 14.550 14.550 15.600 ;
        RECT 18.450 14.550 21.450 16.650 ;
        RECT 6.600 13.800 8.400 14.550 ;
        RECT 4.500 12.900 5.400 13.650 ;
        RECT 9.600 12.900 11.400 13.500 ;
        RECT 4.500 11.700 11.400 12.900 ;
        RECT 10.350 10.500 11.400 11.700 ;
        RECT 20.550 10.500 21.450 14.550 ;
        RECT 30.450 14.250 32.550 14.550 ;
        RECT 28.650 12.450 32.550 14.250 ;
        RECT 33.750 12.450 34.950 21.900 ;
        RECT 10.350 9.600 21.450 10.500 ;
        RECT 30.450 10.350 34.950 12.450 ;
        RECT 10.350 8.700 11.400 9.600 ;
        RECT 20.550 9.300 21.450 9.600 ;
        RECT 1.650 2.250 3.450 8.100 ;
        RECT 6.450 6.000 8.550 8.100 ;
        RECT 10.050 6.900 11.850 8.700 ;
        RECT 13.350 7.950 15.150 8.700 ;
        RECT 13.350 6.900 18.300 7.950 ;
        RECT 20.550 7.500 22.350 9.300 ;
        RECT 33.750 8.100 34.950 10.350 ;
        RECT 27.450 7.200 29.550 8.100 ;
        RECT 7.500 5.100 8.550 6.000 ;
        RECT 17.250 5.100 18.300 6.900 ;
        RECT 25.800 6.000 29.550 7.200 ;
        RECT 25.800 5.100 26.850 6.000 ;
        RECT 4.650 2.250 6.450 5.100 ;
        RECT 7.500 4.200 11.250 5.100 ;
        RECT 9.450 2.250 11.250 4.200 ;
        RECT 13.950 2.250 15.750 5.100 ;
        RECT 17.250 2.250 19.050 5.100 ;
        RECT 21.150 2.250 22.950 5.100 ;
        RECT 25.350 2.250 27.150 5.100 ;
        RECT 29.850 2.250 31.650 5.100 ;
        RECT 33.150 2.250 34.950 8.100 ;
      LAYER metal2 ;
        RECT 6.450 24.900 8.550 27.000 ;
        RECT 27.450 25.800 29.550 27.900 ;
        RECT 6.900 8.100 8.100 24.900 ;
        RECT 27.750 22.200 28.950 25.800 ;
        RECT 27.450 20.100 29.550 22.200 ;
        RECT 12.450 15.750 14.550 16.650 ;
        RECT 18.450 15.750 20.550 16.650 ;
        RECT 27.750 8.100 28.950 20.100 ;
        RECT 30.450 10.350 32.550 11.250 ;
        RECT 6.450 6.000 8.550 8.100 ;
        RECT 27.450 6.000 29.550 8.100 ;
  END
END DFFPOSX1
MACRO DFFSR
  CLASS CORE ;
  FOREIGN DFFSR ;
  ORIGIN 0.000 0.000 ;
  SIZE 72.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END R
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END S
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 27.450 9.450 29.550 11.550 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 54.450 15.450 56.550 17.550 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 66.450 15.450 68.550 17.550 ;
    END
  END Q
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 72.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 72.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.200 27.900 3.000 33.750 ;
        RECT 4.200 27.900 6.000 33.750 ;
        RECT 7.200 27.900 9.000 33.750 ;
        RECT 4.200 27.000 5.250 27.900 ;
        RECT 1.200 26.100 5.250 27.000 ;
        RECT 1.200 12.600 2.400 26.100 ;
        RECT 10.200 25.200 12.000 33.750 ;
        RECT 13.200 30.450 15.000 33.750 ;
        RECT 16.350 30.900 18.750 33.750 ;
        RECT 19.650 30.900 21.750 33.750 ;
        RECT 22.800 30.900 24.750 33.750 ;
        RECT 16.350 29.550 17.550 30.900 ;
        RECT 19.650 29.550 20.550 30.900 ;
        RECT 22.800 29.550 24.000 30.900 ;
        RECT 15.450 27.450 17.550 29.550 ;
        RECT 18.450 27.450 20.550 29.550 ;
        RECT 21.450 27.900 24.000 29.550 ;
        RECT 25.950 27.900 27.750 33.750 ;
        RECT 29.700 27.900 31.500 33.750 ;
        RECT 32.700 27.900 34.500 33.750 ;
        RECT 21.450 27.450 23.550 27.900 ;
        RECT 30.150 27.000 31.500 27.900 ;
        RECT 35.700 27.000 37.500 33.750 ;
        RECT 39.450 30.900 41.250 33.750 ;
        RECT 30.150 25.350 32.550 27.000 ;
        RECT 5.700 24.150 23.400 25.200 ;
        RECT 30.450 24.900 32.550 25.350 ;
        RECT 34.500 26.700 37.500 27.000 ;
        RECT 34.500 24.900 38.400 26.700 ;
        RECT 5.700 23.400 7.500 24.150 ;
        RECT 18.450 22.650 20.550 23.250 ;
        RECT 9.000 21.450 20.550 22.650 ;
        RECT 21.450 23.100 23.400 24.150 ;
        RECT 39.600 23.850 40.950 30.900 ;
        RECT 42.450 27.450 44.250 33.750 ;
        RECT 45.450 30.900 47.250 33.750 ;
        RECT 45.600 29.700 47.100 30.900 ;
        RECT 45.600 27.600 47.700 29.700 ;
        RECT 49.200 27.900 51.000 33.750 ;
        RECT 42.450 26.550 44.550 27.450 ;
        RECT 52.200 27.000 54.000 33.750 ;
        RECT 55.200 27.900 57.000 33.750 ;
        RECT 58.200 27.900 60.000 33.750 ;
        RECT 61.200 27.900 63.000 33.750 ;
        RECT 64.950 27.900 66.750 33.750 ;
        RECT 67.950 27.900 69.750 33.750 ;
        RECT 49.350 26.550 51.150 27.000 ;
        RECT 42.450 25.350 51.150 26.550 ;
        RECT 52.200 25.800 57.900 27.000 ;
        RECT 49.350 25.200 51.150 25.350 ;
        RECT 56.100 25.200 57.900 25.800 ;
        RECT 58.800 23.850 60.000 27.900 ;
        RECT 39.450 23.100 41.550 23.850 ;
        RECT 21.450 21.750 41.550 23.100 ;
        RECT 45.450 22.950 62.850 23.850 ;
        RECT 45.450 21.750 47.550 22.950 ;
        RECT 9.000 20.850 10.800 21.450 ;
        RECT 18.450 21.150 20.550 21.450 ;
        RECT 48.450 20.850 60.750 22.050 ;
        RECT 21.450 19.950 49.500 20.850 ;
        RECT 58.950 20.250 60.750 20.850 ;
        RECT 9.750 19.650 49.500 19.950 ;
        RECT 9.450 19.050 23.400 19.650 ;
        RECT 3.450 16.350 5.550 18.450 ;
        RECT 9.450 17.850 13.350 19.050 ;
        RECT 30.450 18.150 45.000 18.750 ;
        RECT 9.450 17.550 11.550 17.850 ;
        RECT 14.250 16.950 21.000 17.850 ;
        RECT 3.600 14.550 5.400 16.350 ;
        RECT 14.250 14.550 15.450 16.950 ;
        RECT 3.600 13.500 15.450 14.550 ;
        RECT 17.250 14.250 19.050 16.050 ;
        RECT 19.950 15.450 21.000 16.950 ;
        RECT 21.900 17.550 45.000 18.150 ;
        RECT 21.900 16.950 32.550 17.550 ;
        RECT 21.900 16.350 23.700 16.950 ;
        RECT 30.450 16.650 32.550 16.950 ;
        RECT 34.650 15.750 36.750 16.050 ;
        RECT 43.200 15.750 45.000 17.550 ;
        RECT 46.350 16.500 53.400 18.300 ;
        RECT 19.950 14.550 31.950 15.450 ;
        RECT 1.200 11.700 16.500 12.600 ;
        RECT 1.200 8.100 2.400 11.700 ;
        RECT 5.400 10.200 7.200 10.800 ;
        RECT 5.400 9.000 13.800 10.200 ;
        RECT 12.300 8.100 13.800 9.000 ;
        RECT 1.200 2.250 3.000 8.100 ;
        RECT 6.600 2.250 8.400 8.100 ;
        RECT 12.000 2.250 13.800 8.100 ;
        RECT 15.450 8.550 16.500 11.700 ;
        RECT 18.000 10.800 19.050 14.250 ;
        RECT 25.650 11.850 29.550 13.650 ;
        RECT 27.450 11.550 29.550 11.850 ;
        RECT 30.900 13.050 31.950 14.550 ;
        RECT 32.850 13.950 36.750 15.750 ;
        RECT 46.350 14.850 47.250 16.500 ;
        RECT 54.450 15.600 56.550 19.650 ;
        RECT 37.650 13.800 47.250 14.850 ;
        RECT 48.300 14.550 56.550 15.600 ;
        RECT 37.650 13.050 38.550 13.800 ;
        RECT 30.900 11.700 38.550 13.050 ;
        RECT 48.300 12.750 49.350 14.550 ;
        RECT 39.450 11.700 49.350 12.750 ;
        RECT 52.800 11.700 60.600 13.500 ;
        RECT 20.550 10.800 22.350 11.250 ;
        RECT 39.450 10.800 40.500 11.700 ;
        RECT 18.000 10.350 22.350 10.800 ;
        RECT 18.000 9.600 25.650 10.350 ;
        RECT 20.550 9.450 25.650 9.600 ;
        RECT 15.450 6.450 17.550 8.550 ;
        RECT 18.450 6.450 20.550 8.550 ;
        RECT 21.450 6.450 23.550 8.550 ;
        RECT 24.750 8.100 25.650 9.450 ;
        RECT 33.600 9.000 40.500 10.800 ;
        RECT 41.400 9.000 48.150 10.800 ;
        RECT 52.800 8.100 54.300 11.700 ;
        RECT 61.650 8.100 62.850 22.950 ;
        RECT 24.750 6.750 28.800 8.100 ;
        RECT 30.450 7.800 32.550 8.100 ;
        RECT 16.200 5.100 17.550 6.450 ;
        RECT 19.200 5.100 20.550 6.450 ;
        RECT 22.200 5.100 23.550 6.450 ;
        RECT 27.000 6.300 28.800 6.750 ;
        RECT 29.700 6.000 32.550 7.800 ;
        RECT 34.650 7.800 36.750 8.100 ;
        RECT 34.650 6.000 37.500 7.800 ;
        RECT 16.200 2.250 18.000 5.100 ;
        RECT 19.200 2.250 21.000 5.100 ;
        RECT 22.200 2.250 24.000 5.100 ;
        RECT 25.200 2.250 27.000 5.100 ;
        RECT 29.700 2.250 31.500 6.000 ;
        RECT 32.700 2.250 34.500 5.100 ;
        RECT 35.700 2.250 37.500 6.000 ;
        RECT 39.450 6.000 41.550 8.100 ;
        RECT 42.450 6.000 44.550 8.100 ;
        RECT 45.450 6.000 47.550 8.100 ;
        RECT 50.100 6.900 54.300 8.100 ;
        RECT 39.450 2.250 41.250 6.000 ;
        RECT 42.450 2.250 44.250 6.000 ;
        RECT 45.450 2.250 47.250 6.000 ;
        RECT 50.100 2.250 51.900 6.900 ;
        RECT 55.650 2.250 57.450 8.100 ;
        RECT 61.050 2.250 62.850 8.100 ;
        RECT 64.950 15.450 66.450 27.900 ;
        RECT 64.950 13.350 68.550 15.450 ;
        RECT 64.950 5.100 66.450 13.350 ;
        RECT 64.950 2.250 66.750 5.100 ;
        RECT 67.950 2.250 69.750 5.100 ;
      LAYER metal2 ;
        RECT 15.450 27.450 17.550 29.550 ;
        RECT 18.450 27.450 20.550 29.550 ;
        RECT 21.450 27.450 23.550 29.550 ;
        RECT 45.600 27.600 47.700 29.700 ;
        RECT 9.450 18.750 11.550 19.650 ;
        RECT 3.450 16.350 5.550 17.250 ;
        RECT 16.050 8.550 17.250 27.450 ;
        RECT 19.050 23.250 20.250 27.450 ;
        RECT 18.450 21.150 20.550 23.250 ;
        RECT 19.050 8.550 20.250 21.150 ;
        RECT 22.050 8.550 23.250 27.450 ;
        RECT 30.450 24.900 32.550 27.000 ;
        RECT 34.500 24.900 36.600 27.000 ;
        RECT 42.450 25.350 44.550 27.450 ;
        RECT 30.750 18.750 31.950 24.900 ;
        RECT 30.450 16.650 32.550 18.750 ;
        RECT 27.450 12.750 29.550 13.650 ;
        RECT 15.450 6.450 17.550 8.550 ;
        RECT 18.450 6.450 20.550 8.550 ;
        RECT 21.450 6.450 23.550 8.550 ;
        RECT 30.750 8.100 31.950 16.650 ;
        RECT 34.950 16.050 36.150 24.900 ;
        RECT 39.450 21.750 41.550 23.850 ;
        RECT 34.650 13.950 36.750 16.050 ;
        RECT 34.950 8.100 36.150 13.950 ;
        RECT 39.900 8.100 41.100 21.750 ;
        RECT 43.050 8.100 44.250 25.350 ;
        RECT 45.750 23.850 46.950 27.600 ;
        RECT 45.450 21.750 47.550 23.850 ;
        RECT 45.750 8.100 46.950 21.750 ;
        RECT 54.450 18.750 56.550 19.650 ;
        RECT 66.450 13.350 68.550 14.250 ;
        RECT 30.450 6.000 32.550 8.100 ;
        RECT 34.650 6.000 36.750 8.100 ;
        RECT 39.450 6.000 41.550 8.100 ;
        RECT 42.450 6.000 44.550 8.100 ;
        RECT 45.450 6.000 47.550 8.100 ;
  END
END DFFSR
MACRO FAX1
  CLASS CORE ;
  FOREIGN FAX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 45.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.900 12.900 5.100 15.450 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 30.900 12.900 32.100 15.450 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.900 17.550 8.100 20.100 ;
    END
  END C
  PIN YS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 36.900 12.900 38.100 15.450 ;
    END
  END YS
  PIN YC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 39.900 17.550 41.100 20.100 ;
    END
  END YC
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 45.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 45.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 25.800 2.700 36.750 ;
        RECT 3.900 27.000 5.700 36.750 ;
        RECT 6.900 27.000 8.700 36.750 ;
        RECT 6.900 25.800 8.250 27.000 ;
        RECT 9.900 26.100 11.700 36.750 ;
        RECT 0.900 24.900 8.250 25.800 ;
        RECT 9.450 24.000 11.550 26.100 ;
        RECT 14.400 24.900 16.200 36.750 ;
        RECT 17.400 27.000 19.200 36.750 ;
        RECT 20.400 27.900 22.200 36.750 ;
        RECT 23.400 27.000 25.200 36.750 ;
        RECT 17.400 26.100 25.200 27.000 ;
        RECT 26.400 24.000 28.350 36.750 ;
        RECT 32.700 30.900 34.500 36.750 ;
        RECT 35.700 32.250 37.500 36.750 ;
        RECT 35.400 30.900 37.500 32.250 ;
        RECT 39.300 30.900 41.100 36.750 ;
        RECT 42.300 30.900 44.100 36.750 ;
        RECT 21.450 21.900 23.550 24.000 ;
        RECT 24.450 21.900 28.350 24.000 ;
        RECT 35.400 23.400 36.300 30.900 ;
        RECT 37.500 26.400 39.600 26.550 ;
        RECT 37.500 24.600 41.400 26.400 ;
        RECT 37.500 24.450 39.600 24.600 ;
        RECT 42.300 23.400 43.500 30.900 ;
        RECT 35.400 22.500 38.250 23.400 ;
        RECT 21.900 21.300 23.550 21.900 ;
        RECT 21.900 19.500 23.700 21.300 ;
        RECT 27.450 21.150 28.350 21.900 ;
        RECT 27.450 20.250 36.300 21.150 ;
        RECT 34.500 19.350 36.300 20.250 ;
        RECT 3.000 17.550 4.800 19.350 ;
        RECT 19.800 17.700 21.600 18.300 ;
        RECT 25.800 17.700 27.600 18.450 ;
        RECT 19.800 17.550 27.600 17.700 ;
        RECT 3.450 15.450 5.550 17.550 ;
        RECT 6.450 16.500 27.600 17.550 ;
        RECT 28.800 17.550 30.600 18.450 ;
        RECT 37.350 17.550 38.250 22.500 ;
        RECT 39.450 22.200 43.500 23.400 ;
        RECT 39.450 17.550 40.650 22.200 ;
        RECT 6.450 15.750 10.350 16.500 ;
        RECT 6.450 15.450 8.550 15.750 ;
        RECT 28.800 15.600 32.550 17.550 ;
        RECT 3.600 11.700 5.100 15.450 ;
        RECT 17.400 14.550 32.550 15.600 ;
        RECT 36.450 15.450 38.550 17.550 ;
        RECT 39.450 15.450 41.550 17.550 ;
        RECT 6.000 13.650 7.800 14.550 ;
        RECT 11.400 13.650 13.200 14.550 ;
        RECT 17.400 13.650 19.200 14.550 ;
        RECT 6.000 12.600 19.200 13.650 ;
        RECT 22.050 11.700 29.700 12.600 ;
        RECT 3.600 10.800 23.250 11.700 ;
        RECT 28.500 10.800 33.900 11.700 ;
        RECT 14.400 9.900 16.200 10.800 ;
        RECT 0.900 7.200 8.100 8.100 ;
        RECT 9.450 7.800 11.550 9.900 ;
        RECT 24.450 8.700 27.450 10.800 ;
        RECT 32.100 9.750 33.900 10.800 ;
        RECT 0.900 2.250 2.700 7.200 ;
        RECT 3.900 2.250 5.700 6.300 ;
        RECT 6.900 2.250 8.700 7.200 ;
        RECT 9.900 6.900 11.550 7.800 ;
        RECT 9.900 2.250 11.700 6.900 ;
        RECT 14.400 2.250 16.200 7.500 ;
        RECT 17.400 6.900 25.200 7.800 ;
        RECT 17.400 2.250 19.200 6.900 ;
        RECT 20.400 2.250 22.200 6.000 ;
        RECT 23.400 2.250 25.200 6.900 ;
        RECT 26.400 6.600 27.450 8.700 ;
        RECT 37.350 7.200 38.250 15.450 ;
        RECT 26.400 2.250 28.350 6.600 ;
        RECT 36.000 6.000 38.250 7.200 ;
        RECT 36.000 5.100 36.900 6.000 ;
        RECT 39.450 5.100 40.500 15.450 ;
        RECT 32.700 2.250 34.500 5.100 ;
        RECT 35.700 2.250 37.500 5.100 ;
        RECT 39.300 2.250 41.100 5.100 ;
        RECT 42.300 2.250 44.100 5.100 ;
      LAYER metal2 ;
        RECT 37.500 26.100 39.600 26.550 ;
        RECT 9.450 25.200 39.600 26.100 ;
        RECT 9.450 24.000 11.550 25.200 ;
        RECT 3.450 16.650 5.550 17.550 ;
        RECT 6.450 15.450 8.550 16.350 ;
        RECT 10.050 9.900 10.950 24.000 ;
        RECT 21.450 21.900 23.550 25.200 ;
        RECT 37.500 24.450 39.600 25.200 ;
        RECT 24.450 21.900 26.550 24.000 ;
        RECT 25.050 10.800 26.250 21.900 ;
        RECT 30.450 16.650 32.550 17.550 ;
        RECT 36.450 16.650 38.550 17.550 ;
        RECT 39.450 15.450 41.550 16.350 ;
        RECT 9.450 7.800 11.550 9.900 ;
        RECT 24.450 8.700 26.550 10.800 ;
  END
END FAX1
MACRO FILL
  CLASS CORE ;
  FOREIGN FILL ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 3.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 3.900 1.200 ;
    END
  END gnd
END FILL
MACRO HAX1
  CLASS CORE ;
  FOREIGN HAX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.900 12.900 2.100 15.450 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 15.900 17.550 17.100 20.100 ;
    END
  END B
  PIN YS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 21.900 12.900 23.100 15.450 ;
    END
  END YS
  PIN YC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.900 17.550 11.100 20.100 ;
    END
  END YC
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 30.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 30.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 30.900 2.700 36.750 ;
        RECT 3.900 31.500 5.700 36.750 ;
        RECT 1.200 30.600 2.700 30.900 ;
        RECT 6.900 30.900 8.700 36.750 ;
        RECT 10.500 30.900 12.300 36.750 ;
        RECT 13.500 30.900 15.300 36.750 ;
        RECT 6.900 30.600 8.100 30.900 ;
        RECT 1.200 29.700 8.100 30.600 ;
        RECT 7.050 17.850 8.100 29.700 ;
        RECT 0.450 17.400 2.550 17.550 ;
        RECT 0.450 15.450 4.350 17.400 ;
        RECT 6.450 15.750 8.550 17.850 ;
        RECT 10.500 17.550 11.550 30.900 ;
        RECT 16.500 24.900 18.300 36.750 ;
        RECT 20.700 30.900 22.500 36.750 ;
        RECT 23.700 30.900 25.500 36.750 ;
        RECT 16.650 22.950 17.550 24.900 ;
        RECT 16.650 22.050 19.950 22.950 ;
        RECT 9.450 15.450 11.550 17.550 ;
        RECT 15.450 15.450 17.550 17.550 ;
        RECT 2.850 12.150 4.200 15.450 ;
        RECT 6.000 14.550 7.800 14.850 ;
        RECT 15.600 14.550 17.400 15.450 ;
        RECT 6.000 13.650 17.400 14.550 ;
        RECT 18.600 14.250 19.950 22.050 ;
        RECT 23.700 17.550 24.600 30.900 ;
        RECT 21.450 15.450 24.600 17.550 ;
        RECT 6.000 13.050 7.800 13.650 ;
        RECT 18.600 13.350 22.200 14.250 ;
        RECT 18.600 12.150 20.400 12.450 ;
        RECT 2.850 11.100 20.400 12.150 ;
        RECT 18.600 10.650 20.400 11.100 ;
        RECT 21.300 10.650 22.200 13.350 ;
        RECT 23.700 12.450 24.600 15.450 ;
        RECT 23.700 11.550 28.200 12.450 ;
        RECT 5.100 9.900 8.550 10.200 ;
        RECT 5.100 8.100 11.550 9.900 ;
        RECT 21.300 9.750 23.400 10.650 ;
        RECT 17.850 8.850 23.400 9.750 ;
        RECT 17.850 8.100 19.650 8.850 ;
        RECT 0.900 2.250 2.700 8.100 ;
        RECT 5.100 2.250 6.900 8.100 ;
        RECT 8.700 4.950 10.800 7.200 ;
        RECT 8.700 2.250 10.500 4.950 ;
        RECT 11.700 2.250 13.500 5.100 ;
        RECT 14.700 3.000 16.500 8.100 ;
        RECT 17.700 3.900 19.500 8.100 ;
        RECT 20.700 3.000 22.500 7.500 ;
        RECT 27.300 5.100 28.200 11.550 ;
        RECT 14.700 2.250 22.500 3.000 ;
        RECT 24.300 2.250 26.100 5.100 ;
        RECT 27.300 2.250 29.100 5.100 ;
      LAYER metal2 ;
        RECT 0.450 16.650 2.550 17.550 ;
        RECT 6.450 15.750 8.550 17.850 ;
        RECT 21.450 16.650 23.550 17.550 ;
        RECT 6.900 10.200 7.950 15.750 ;
        RECT 9.450 15.450 11.550 16.350 ;
        RECT 15.450 15.450 17.550 16.350 ;
        RECT 6.450 8.100 8.550 10.200 ;
        RECT 10.200 7.200 11.400 15.450 ;
        RECT 8.700 5.100 11.400 7.200 ;
  END
END HAX1
MACRO INVX1
  CLASS CORE ;
  FOREIGN INVX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 9.450 2.550 11.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 9.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 9.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 27.900 2.850 33.750 ;
        RECT 4.050 27.900 5.850 33.750 ;
        RECT 3.900 15.450 5.100 27.900 ;
        RECT 0.600 13.650 2.400 15.450 ;
        RECT 0.450 11.550 2.550 13.650 ;
        RECT 3.450 13.350 5.550 15.450 ;
        RECT 3.900 5.100 5.100 13.350 ;
        RECT 1.050 2.250 2.850 5.100 ;
        RECT 4.050 2.250 5.850 5.100 ;
      LAYER metal2 ;
        RECT 0.450 12.750 2.550 13.650 ;
        RECT 3.450 13.350 5.550 14.250 ;
  END
END INVX1
MACRO INVX2
  CLASS CORE ;
  FOREIGN INVX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 15.450 2.550 17.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 12.450 5.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 9.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 9.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 21.900 2.850 33.750 ;
        RECT 4.050 21.900 5.850 33.750 ;
        RECT 3.900 16.650 5.100 21.900 ;
        RECT 0.450 13.350 2.550 15.450 ;
        RECT 3.450 14.550 5.550 16.650 ;
        RECT 0.600 11.550 2.400 13.350 ;
        RECT 3.900 8.100 5.100 14.550 ;
        RECT 1.050 2.250 2.850 8.100 ;
        RECT 4.050 2.250 5.850 8.100 ;
      LAYER metal2 ;
        RECT 3.750 15.750 5.550 16.650 ;
        RECT 0.450 13.350 2.250 14.250 ;
  END
END INVX2
MACRO INVX4
  CLASS CORE ;
  FOREIGN INVX4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 15.450 2.550 17.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.450 15.450 8.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 12.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 12.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 21.900 2.850 33.750 ;
        RECT 4.050 21.900 5.850 33.750 ;
        RECT 7.050 21.900 8.850 33.750 ;
        RECT 4.350 15.450 5.700 21.900 ;
        RECT 0.450 13.350 2.550 15.450 ;
        RECT 4.350 13.350 8.550 15.450 ;
        RECT 0.600 11.550 2.400 13.350 ;
        RECT 4.350 8.100 5.700 13.350 ;
        RECT 1.050 2.250 2.850 8.100 ;
        RECT 4.050 2.250 5.850 8.100 ;
        RECT 7.050 2.250 8.850 8.100 ;
      LAYER metal2 ;
        RECT 0.450 13.350 2.550 14.250 ;
        RECT 6.450 13.350 8.550 14.250 ;
  END
END INVX4
MACRO INVX8
  CLASS CORE ;
  FOREIGN INVX8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 12.450 5.550 14.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.450 12.450 11.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 18.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 18.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 21.900 2.850 33.750 ;
        RECT 4.050 21.000 5.850 33.750 ;
        RECT 7.050 21.900 8.850 33.750 ;
        RECT 10.050 21.900 11.850 33.750 ;
        RECT 13.050 21.900 14.850 33.750 ;
        RECT 10.050 21.000 11.250 21.900 ;
        RECT 4.050 20.100 11.250 21.000 ;
        RECT 3.600 16.650 5.400 18.450 ;
        RECT 10.050 16.650 11.250 20.100 ;
        RECT 3.450 14.550 5.550 16.650 ;
        RECT 9.450 14.550 11.550 16.650 ;
        RECT 10.050 10.200 11.250 14.550 ;
        RECT 4.050 9.000 11.250 10.200 ;
        RECT 4.050 8.100 5.250 9.000 ;
        RECT 10.050 8.100 11.250 9.000 ;
        RECT 1.050 2.250 2.850 8.100 ;
        RECT 4.050 2.250 5.850 8.100 ;
        RECT 7.050 2.250 8.850 8.100 ;
        RECT 10.050 2.250 11.850 8.100 ;
        RECT 13.050 2.250 14.850 8.100 ;
      LAYER metal2 ;
        RECT 3.450 15.750 5.550 16.650 ;
        RECT 9.450 15.750 11.550 16.650 ;
  END
END INVX8
MACRO LATCH
  CLASS CORE ;
  FOREIGN LATCH ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 12.900 20.550 14.100 23.100 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.900 14.550 5.100 17.100 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 15.900 12.900 17.100 15.450 ;
    END
  END Q
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 21.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 21.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.200 24.900 3.000 36.750 ;
        RECT 4.200 24.900 6.000 36.750 ;
        RECT 9.300 30.900 11.250 36.750 ;
        RECT 9.450 28.800 11.550 30.900 ;
        RECT 15.000 24.900 16.800 36.750 ;
        RECT 18.000 24.900 19.800 36.750 ;
        RECT 1.200 21.300 2.400 24.900 ;
        RECT 9.450 24.000 11.550 24.900 ;
        RECT 9.450 22.800 17.400 24.000 ;
        RECT 15.600 22.200 17.400 22.800 ;
        RECT 1.200 20.400 9.900 21.300 ;
        RECT 1.200 8.100 2.400 20.400 ;
        RECT 8.100 19.500 9.900 20.400 ;
        RECT 5.100 18.450 6.900 19.350 ;
        RECT 11.700 18.450 14.550 20.550 ;
        RECT 5.100 17.550 12.750 18.450 ;
        RECT 18.600 17.550 19.800 24.900 ;
        RECT 15.450 17.250 19.800 17.550 ;
        RECT 13.650 15.450 19.800 17.250 ;
        RECT 9.900 14.550 11.700 14.850 ;
        RECT 3.450 13.050 11.700 14.550 ;
        RECT 3.450 12.450 5.550 13.050 ;
        RECT 3.300 10.650 5.100 12.450 ;
        RECT 8.550 9.900 9.600 13.050 ;
        RECT 8.550 8.100 10.350 9.900 ;
        RECT 18.600 8.100 19.800 15.450 ;
        RECT 1.200 2.250 3.000 8.100 ;
        RECT 9.450 5.100 11.550 7.200 ;
        RECT 4.200 2.250 6.000 5.100 ;
        RECT 9.300 2.250 11.400 5.100 ;
        RECT 15.000 2.250 16.800 8.100 ;
        RECT 18.000 2.250 19.800 8.100 ;
      LAYER metal2 ;
        RECT 9.450 28.800 11.550 30.900 ;
        RECT 9.600 24.900 10.800 28.800 ;
        RECT 9.450 22.800 11.550 24.900 ;
        RECT 3.450 12.450 5.550 13.350 ;
        RECT 9.600 7.200 10.800 22.800 ;
        RECT 12.450 18.450 14.550 19.350 ;
        RECT 15.450 16.650 17.550 17.550 ;
        RECT 9.450 5.100 11.550 7.200 ;
  END
END LATCH
MACRO MUX2X1
  CLASS CORE ;
  FOREIGN MUX2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 12.450 12.450 14.550 14.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 12.450 5.550 14.550 ;
    END
  END B
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 15.450 2.550 17.550 ;
    END
  END S
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 18.750 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 18.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 26.700 2.850 32.700 ;
        RECT 4.050 26.700 5.850 33.750 ;
        RECT 1.950 21.600 2.850 26.700 ;
        RECT 8.550 23.400 10.350 32.700 ;
        RECT 8.550 22.500 10.650 23.400 ;
        RECT 1.950 20.700 8.100 21.600 ;
        RECT 3.750 16.650 5.550 18.450 ;
        RECT 0.450 13.350 2.550 15.450 ;
        RECT 3.450 14.550 5.550 16.650 ;
        RECT 6.750 18.000 8.100 20.700 ;
        RECT 6.750 16.200 8.550 18.000 ;
        RECT 0.750 11.550 2.550 13.350 ;
        RECT 6.750 10.500 8.100 16.200 ;
        RECT 9.750 15.450 10.650 22.500 ;
        RECT 13.050 21.900 14.850 33.750 ;
        RECT 12.600 16.650 14.400 18.450 ;
        RECT 9.450 13.350 11.550 15.450 ;
        RECT 12.450 14.550 14.550 16.650 ;
        RECT 1.800 9.600 8.100 10.500 ;
        RECT 1.800 6.300 2.850 9.600 ;
        RECT 9.750 8.700 10.650 13.350 ;
        RECT 8.550 7.800 10.650 8.700 ;
        RECT 1.050 3.300 2.850 6.300 ;
        RECT 4.050 2.250 5.850 6.300 ;
        RECT 8.550 3.300 10.350 7.800 ;
        RECT 13.050 2.250 14.850 9.300 ;
      LAYER metal2 ;
        RECT 3.750 15.750 5.550 16.650 ;
        RECT 12.750 15.750 14.550 16.650 ;
        RECT 0.450 13.350 2.250 14.250 ;
        RECT 9.450 13.350 11.250 14.250 ;
  END
END MUX2X1
MACRO NAND2X1
  CLASS CORE ;
  FOREIGN NAND2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 12.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 12.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 27.900 2.850 33.750 ;
        RECT 4.050 27.900 5.850 33.750 ;
        RECT 7.050 27.900 8.850 33.750 ;
        RECT 4.050 19.650 5.250 27.900 ;
        RECT 0.450 16.350 2.550 18.450 ;
        RECT 3.450 17.550 5.550 19.650 ;
        RECT 0.600 14.550 2.400 16.350 ;
        RECT 4.050 10.200 5.250 17.550 ;
        RECT 6.450 16.350 8.550 18.450 ;
        RECT 6.600 14.550 8.400 16.350 ;
        RECT 4.050 9.300 7.650 10.200 ;
        RECT 1.350 2.250 3.150 8.100 ;
        RECT 5.850 2.250 7.650 9.300 ;
      LAYER metal2 ;
        RECT 3.750 18.750 5.250 19.650 ;
        RECT 0.450 16.350 2.250 17.250 ;
        RECT 6.750 16.350 8.550 17.250 ;
  END
END NAND2X1
MACRO NAND3X1
  CLASS CORE ;
  FOREIGN NAND3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 15.450 2.550 17.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.450 15.450 8.550 17.550 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 15.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 27.900 2.850 33.750 ;
        RECT 4.050 27.900 5.850 33.750 ;
        RECT 7.050 28.500 8.850 33.750 ;
        RECT 4.200 27.600 5.850 27.900 ;
        RECT 10.050 27.900 11.850 33.750 ;
        RECT 10.050 27.600 11.250 27.900 ;
        RECT 4.200 26.700 11.250 27.600 ;
        RECT 3.600 22.650 5.400 24.450 ;
        RECT 0.600 19.650 2.400 21.450 ;
        RECT 3.450 20.550 5.550 22.650 ;
        RECT 6.750 19.650 8.550 21.450 ;
        RECT 0.450 17.550 2.550 19.650 ;
        RECT 6.450 17.550 8.550 19.650 ;
        RECT 10.200 18.450 11.250 26.700 ;
        RECT 9.450 16.350 11.550 18.450 ;
        RECT 9.900 12.150 11.100 16.350 ;
        RECT 1.200 2.250 3.000 11.100 ;
        RECT 6.600 10.500 11.100 12.150 ;
        RECT 6.600 2.250 8.400 10.500 ;
      LAYER metal2 ;
        RECT 3.450 21.750 5.550 22.650 ;
        RECT 0.450 18.750 2.250 19.650 ;
        RECT 6.750 18.750 8.250 19.650 ;
        RECT 9.750 16.350 11.550 17.250 ;
  END
END NAND3X1
MACRO NOR2X1
  CLASS CORE ;
  FOREIGN NOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 12.450 2.550 14.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.450 12.450 8.550 14.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 9.450 5.550 11.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 12.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 12.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 21.900 2.850 33.750 ;
        RECT 5.250 21.900 7.050 33.750 ;
        RECT 4.500 20.850 7.050 21.900 ;
        RECT 0.600 16.650 2.400 18.450 ;
        RECT 0.450 14.550 2.550 16.650 ;
        RECT 4.500 13.650 5.550 20.850 ;
        RECT 6.600 16.650 8.400 18.450 ;
        RECT 6.450 14.550 8.550 16.650 ;
        RECT 3.450 11.550 5.550 13.650 ;
        RECT 4.500 5.100 5.550 11.550 ;
        RECT 1.050 2.250 2.850 5.100 ;
        RECT 4.050 2.250 5.850 5.100 ;
        RECT 7.050 2.250 8.850 5.100 ;
      LAYER metal2 ;
        RECT 0.450 15.750 2.550 16.650 ;
        RECT 6.450 15.750 8.550 16.650 ;
        RECT 3.750 12.750 5.250 13.650 ;
  END
END NOR2X1
MACRO NOR3X1
  CLASS CORE ;
  FOREIGN NOR3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 12.450 5.550 14.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 12.450 12.450 14.550 14.550 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 18.450 15.450 20.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 27.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 27.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 24.000 2.850 33.750 ;
        RECT 4.050 24.900 5.850 33.750 ;
        RECT 7.050 33.000 14.850 33.750 ;
        RECT 7.050 24.000 8.850 33.000 ;
        RECT 1.050 23.100 8.850 24.000 ;
        RECT 10.050 24.300 11.850 32.100 ;
        RECT 13.050 25.200 14.850 33.000 ;
        RECT 16.650 33.000 24.450 33.750 ;
        RECT 16.650 24.300 18.450 33.000 ;
        RECT 10.050 23.400 18.450 24.300 ;
        RECT 19.650 24.300 21.450 32.100 ;
        RECT 19.650 21.900 20.850 24.300 ;
        RECT 22.650 23.700 24.450 33.000 ;
        RECT 17.400 20.700 20.850 21.900 ;
        RECT 3.600 16.650 5.400 18.450 ;
        RECT 12.600 16.650 14.400 18.450 ;
        RECT 3.450 14.550 5.550 16.650 ;
        RECT 9.450 13.350 11.550 15.450 ;
        RECT 12.450 14.550 14.550 16.650 ;
        RECT 17.400 15.450 18.600 20.700 ;
        RECT 17.400 13.350 20.550 15.450 ;
        RECT 9.600 11.550 11.400 13.350 ;
        RECT 17.400 6.900 18.600 13.350 ;
        RECT 7.800 6.000 18.600 6.900 ;
        RECT 7.800 5.100 8.850 6.000 ;
        RECT 13.800 5.100 14.850 6.000 ;
        RECT 3.750 2.250 5.850 5.100 ;
        RECT 7.050 2.250 8.850 5.100 ;
        RECT 10.050 2.250 11.850 5.100 ;
        RECT 13.050 2.250 14.850 5.100 ;
      LAYER metal2 ;
        RECT 3.450 15.750 5.550 16.650 ;
        RECT 12.750 15.750 14.550 16.650 ;
        RECT 9.450 13.350 11.250 14.250 ;
        RECT 18.450 13.350 20.550 14.250 ;
  END
END NOR3X1
MACRO OAI21X1
  CLASS CORE ;
  FOREIGN OAI21X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 12.450 2.550 14.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.450 12.450 8.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 15.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.800 21.900 3.600 33.750 ;
        RECT 6.000 21.900 7.800 33.750 ;
        RECT 9.300 27.900 11.100 33.750 ;
        RECT 0.600 16.650 2.400 18.450 ;
        RECT 6.450 16.650 7.650 21.900 ;
        RECT 9.450 19.650 11.250 21.450 ;
        RECT 9.450 17.550 11.550 19.650 ;
        RECT 0.450 14.550 2.550 16.650 ;
        RECT 3.450 13.350 5.550 15.450 ;
        RECT 6.450 14.550 8.550 16.650 ;
        RECT 3.600 11.550 5.400 13.350 ;
        RECT 7.350 11.250 8.550 14.550 ;
        RECT 7.500 10.200 11.250 11.250 ;
        RECT 1.050 7.200 8.850 8.550 ;
        RECT 1.050 2.250 2.850 7.200 ;
        RECT 4.050 2.250 5.850 6.300 ;
        RECT 7.050 2.250 8.850 7.200 ;
        RECT 10.050 8.100 11.250 10.200 ;
        RECT 10.050 2.250 11.850 8.100 ;
      LAYER metal2 ;
        RECT 9.450 18.750 11.550 19.650 ;
        RECT 0.450 15.750 2.250 16.650 ;
        RECT 6.750 15.750 8.250 16.650 ;
        RECT 3.750 13.350 5.250 14.250 ;
  END
END OAI21X1
MACRO OAI22X1
  CLASS CORE ;
  FOREIGN OAI22X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 12.450 2.550 14.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 12.450 12.450 14.550 14.550 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.450 12.450 8.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 18.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 18.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 21.900 2.850 33.750 ;
        RECT 5.550 21.900 8.850 33.750 ;
        RECT 11.550 21.900 13.350 33.750 ;
        RECT 0.600 16.650 2.400 18.450 ;
        RECT 7.050 16.650 8.250 21.900 ;
        RECT 12.450 16.650 14.250 18.450 ;
        RECT 0.450 14.550 2.550 16.650 ;
        RECT 3.450 13.350 5.550 15.450 ;
        RECT 6.450 14.550 8.550 16.650 ;
        RECT 3.600 11.550 5.400 13.350 ;
        RECT 6.900 10.650 8.100 14.550 ;
        RECT 9.450 13.350 11.550 15.450 ;
        RECT 12.450 14.550 14.550 16.650 ;
        RECT 9.000 11.550 10.800 13.350 ;
        RECT 6.900 9.600 11.250 10.650 ;
        RECT 1.050 7.500 8.850 8.400 ;
        RECT 10.350 8.100 11.250 9.600 ;
        RECT 1.050 2.250 2.850 7.500 ;
        RECT 4.050 2.250 5.850 6.600 ;
        RECT 7.050 3.000 8.850 7.500 ;
        RECT 10.050 3.900 11.850 8.100 ;
        RECT 13.050 3.000 14.850 8.100 ;
        RECT 7.050 2.250 14.850 3.000 ;
      LAYER metal2 ;
        RECT 0.450 15.750 2.250 16.650 ;
        RECT 6.750 15.750 8.250 16.650 ;
        RECT 12.750 15.750 14.550 16.650 ;
        RECT 3.750 13.350 5.250 14.250 ;
        RECT 9.750 13.350 11.250 14.250 ;
  END
END OAI22X1
MACRO OR2X1
  CLASS CORE ;
  FOREIGN OR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 9.450 2.550 11.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 12.450 5.550 14.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.450 12.450 11.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 34.800 15.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 21.000 2.850 33.750 ;
        RECT 5.550 21.900 7.350 33.750 ;
        RECT 8.850 27.900 10.650 33.750 ;
        RECT 8.850 27.000 11.550 27.900 ;
        RECT 1.050 20.100 9.450 21.000 ;
        RECT 7.350 19.200 9.450 20.100 ;
        RECT 0.600 13.650 2.400 15.450 ;
        RECT 0.450 11.550 2.550 13.650 ;
        RECT 3.450 10.350 5.550 12.450 ;
        RECT 3.600 8.550 5.400 10.350 ;
        RECT 7.350 8.400 8.550 19.200 ;
        RECT 10.350 12.450 11.550 27.000 ;
        RECT 9.450 10.350 11.850 12.450 ;
        RECT 7.350 7.500 9.750 8.400 ;
        RECT 4.350 6.600 9.750 7.500 ;
        RECT 4.350 5.100 5.250 6.600 ;
        RECT 10.650 5.100 11.850 10.350 ;
        RECT 1.050 2.250 2.850 5.100 ;
        RECT 4.050 2.250 5.850 5.100 ;
        RECT 7.050 2.250 8.850 5.100 ;
        RECT 10.050 2.250 11.850 5.100 ;
      LAYER metal2 ;
        RECT 0.450 12.750 2.250 13.650 ;
        RECT 3.750 10.350 5.550 11.250 ;
        RECT 9.450 10.350 11.550 11.250 ;
  END
END OR2X1
MACRO OR2X2
  CLASS CORE ;
  FOREIGN OR2X2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 36.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.450 9.450 2.550 11.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 3.450 12.450 5.550 14.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 34.800 15.900 37.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 21.900 2.850 33.750 ;
        RECT 5.550 22.050 7.350 33.750 ;
        RECT 8.550 23.400 10.350 33.750 ;
        RECT 8.550 22.050 10.950 23.400 ;
        RECT 1.050 20.700 2.250 21.900 ;
        RECT 6.450 20.700 8.250 21.150 ;
        RECT 1.050 19.500 8.250 20.700 ;
        RECT 6.450 19.350 8.250 19.500 ;
        RECT 3.600 16.650 5.400 18.450 ;
        RECT 0.600 13.650 2.400 15.450 ;
        RECT 3.450 14.550 5.550 16.650 ;
        RECT 0.450 11.550 2.550 13.650 ;
        RECT 7.200 11.100 8.100 19.350 ;
        RECT 9.600 15.450 10.950 22.050 ;
        RECT 9.450 13.350 11.550 15.450 ;
        RECT 6.450 10.200 8.250 11.100 ;
        RECT 4.950 9.300 8.250 10.200 ;
        RECT 4.950 5.100 5.850 9.300 ;
        RECT 10.500 8.100 11.550 13.350 ;
        RECT 1.050 2.250 2.850 5.100 ;
        RECT 4.050 2.250 5.850 5.100 ;
        RECT 7.050 2.250 8.850 5.100 ;
        RECT 10.050 2.250 11.850 8.100 ;
      LAYER metal2 ;
        RECT 3.450 15.750 5.550 16.650 ;
        RECT 0.450 12.750 2.250 13.650 ;
        RECT 9.450 13.350 11.550 14.250 ;
  END
END OR2X2
MACRO TBUFX1
  CLASS CORE ;
  FOREIGN TBUFX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 11.400 17.550 12.600 20.100 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.900 17.550 2.100 20.100 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 6.900 17.550 8.100 20.100 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 16.050 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 16.050 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.200 30.900 3.000 36.750 ;
        RECT 4.200 30.900 6.000 36.750 ;
        RECT 5.100 23.550 6.000 30.900 ;
        RECT 7.500 24.900 9.300 36.750 ;
        RECT 12.000 24.900 13.800 36.750 ;
        RECT 5.100 21.750 6.900 23.550 ;
        RECT 1.200 17.550 3.000 19.200 ;
        RECT 0.900 15.450 3.000 17.550 ;
        RECT 5.100 5.100 6.000 21.750 ;
        RECT 7.950 17.550 9.000 24.900 ;
        RECT 10.800 17.550 12.600 19.200 ;
        RECT 6.900 15.450 9.000 17.550 ;
        RECT 10.500 15.450 12.600 17.550 ;
        RECT 7.950 8.100 9.000 15.450 ;
        RECT 1.200 2.250 3.000 5.100 ;
        RECT 4.200 2.250 6.000 5.100 ;
        RECT 7.500 2.250 9.300 8.100 ;
        RECT 12.000 2.250 13.800 8.100 ;
      LAYER metal2 ;
        RECT 0.900 15.450 3.000 16.200 ;
        RECT 6.900 15.450 9.000 16.350 ;
        RECT 10.500 15.450 12.600 16.350 ;
  END
END TBUFX1
MACRO TBUFX2
  CLASS CORE ;
  FOREIGN TBUFX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 15.900 17.550 17.100 20.100 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.900 17.550 2.100 20.100 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.900 17.550 11.100 20.100 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 22.050 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 22.050 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 24.900 2.400 36.750 ;
        RECT 3.600 24.900 5.400 36.750 ;
        RECT 6.600 36.000 14.400 36.750 ;
        RECT 6.600 24.900 8.400 36.000 ;
        RECT 9.600 24.900 11.400 35.100 ;
        RECT 12.600 26.100 14.400 36.000 ;
        RECT 15.600 27.000 17.400 36.750 ;
        RECT 18.600 26.100 20.400 36.750 ;
        RECT 12.600 24.900 20.400 26.100 ;
        RECT 4.500 22.950 5.400 24.900 ;
        RECT 4.500 21.150 6.300 22.950 ;
        RECT 0.900 15.450 3.000 17.550 ;
        RECT 1.500 13.650 3.300 15.450 ;
        RECT 4.500 8.100 5.400 21.150 ;
        RECT 9.600 17.550 10.500 24.900 ;
        RECT 9.600 15.450 11.700 17.550 ;
        RECT 15.600 15.450 17.700 17.550 ;
        RECT 9.600 8.100 10.500 15.450 ;
        RECT 15.900 13.650 17.700 15.450 ;
        RECT 12.600 8.100 19.800 9.000 ;
        RECT 0.600 2.250 2.400 8.100 ;
        RECT 3.600 2.250 5.400 8.100 ;
        RECT 6.600 3.000 8.400 8.100 ;
        RECT 9.600 3.900 11.400 8.100 ;
        RECT 12.600 3.000 14.400 8.100 ;
        RECT 6.600 2.250 14.400 3.000 ;
        RECT 15.600 2.250 17.400 7.200 ;
        RECT 18.600 2.250 20.400 8.100 ;
      LAYER metal2 ;
        RECT 0.900 15.450 3.000 16.350 ;
        RECT 9.600 15.450 11.700 16.350 ;
        RECT 15.600 15.450 17.700 16.350 ;
  END
END TBUFX2
MACRO XNOR2X1
  CLASS CORE ;
  FOREIGN XNOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.900 15.300 3.000 17.400 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15.450 15.300 17.550 17.400 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.900 18.300 12.000 20.400 ;
    END
    PORT
      LAYER metal1 ;
        RECT 9.900 9.600 12.000 11.700 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 21.900 40.200 ;
        RECT 3.900 27.000 5.700 37.800 ;
        RECT 12.600 27.000 14.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3.900 1.200 5.700 7.200 ;
        RECT 12.600 1.200 14.400 7.200 ;
        RECT -0.900 -1.200 21.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 25.800 2.700 36.900 ;
        RECT 8.400 25.800 10.200 36.900 ;
        RECT 15.900 26.100 17.700 36.900 ;
        RECT 0.900 24.600 5.700 25.800 ;
        RECT 8.400 24.900 11.700 25.800 ;
        RECT 3.600 23.700 5.700 24.600 ;
        RECT 3.600 22.800 9.000 23.700 ;
        RECT 7.200 21.450 9.000 22.800 ;
        RECT 10.500 21.450 11.700 24.900 ;
        RECT 12.600 24.900 17.700 26.100 ;
        RECT 12.600 24.000 14.700 24.900 ;
        RECT 7.200 20.700 8.850 21.450 ;
        RECT 5.700 17.700 7.500 19.500 ;
        RECT 15.600 18.450 17.400 19.200 ;
        RECT 5.700 15.600 7.800 17.700 ;
        RECT 4.050 14.250 7.800 14.700 ;
        RECT 1.200 13.500 7.800 14.250 ;
        RECT 5.700 12.600 7.800 13.500 ;
        RECT 8.850 12.750 9.750 17.250 ;
        RECT 10.800 15.600 12.600 17.250 ;
        RECT 10.650 13.500 12.750 15.600 ;
        RECT 3.150 10.500 5.250 11.100 ;
        RECT 6.150 10.800 7.950 12.600 ;
        RECT 0.900 9.000 5.250 10.500 ;
        RECT 13.200 9.300 15.300 11.400 ;
        RECT 0.900 8.100 2.400 9.000 ;
        RECT 0.900 2.100 2.700 8.100 ;
        RECT 8.850 7.500 9.900 8.550 ;
        RECT 13.200 8.100 17.700 9.300 ;
        RECT 8.100 2.100 9.900 7.500 ;
        RECT 15.900 2.100 17.700 8.100 ;
      LAYER metal2 ;
        RECT 3.600 23.700 5.700 25.800 ;
        RECT 12.600 24.000 14.700 26.100 ;
        RECT 3.900 11.100 4.800 23.700 ;
        RECT 5.700 17.400 7.800 17.700 ;
        RECT 13.650 17.400 14.550 24.000 ;
        RECT 5.700 16.500 14.550 17.400 ;
        RECT 5.700 15.600 7.800 16.500 ;
        RECT 10.650 14.700 12.750 15.600 ;
        RECT 5.700 13.500 12.750 14.700 ;
        RECT 5.700 12.600 7.800 13.500 ;
        RECT 13.650 11.400 14.550 16.500 ;
        RECT 3.150 9.000 5.250 11.100 ;
        RECT 13.200 9.300 15.300 11.400 ;
  END
END XNOR2X1
MACRO XOR2X1
  CLASS CORE ;
  FOREIGN XOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.900 15.450 3.000 17.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15.450 15.450 17.550 17.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.600 18.300 11.700 20.400 ;
    END
    PORT
      LAYER metal1 ;
        RECT 9.600 9.600 11.700 11.700 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 21.750 40.200 ;
        RECT 3.900 27.000 5.700 37.800 ;
        RECT 12.900 27.000 14.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3.900 1.200 5.700 7.200 ;
        RECT 12.900 1.200 14.700 7.200 ;
        RECT -0.900 -1.200 21.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 25.800 2.700 36.900 ;
        RECT 0.900 24.900 5.400 25.800 ;
        RECT 8.400 24.900 10.200 36.900 ;
        RECT 15.900 26.100 17.700 36.900 ;
        RECT 3.300 22.800 5.400 24.900 ;
        RECT 9.000 23.400 10.200 24.900 ;
        RECT 12.900 24.900 17.700 26.100 ;
        RECT 12.900 24.000 15.000 24.900 ;
        RECT 9.000 22.500 10.500 23.400 ;
        RECT 9.600 21.450 10.500 22.500 ;
        RECT 6.600 21.000 8.550 21.300 ;
        RECT 4.800 19.200 8.550 21.000 ;
        RECT 15.600 18.600 17.400 19.350 ;
        RECT 6.000 17.400 7.800 18.000 ;
        RECT 4.050 16.200 7.800 17.400 ;
        RECT 0.900 13.650 2.700 14.400 ;
        RECT 6.000 12.900 7.800 14.700 ;
        RECT 5.700 10.800 7.800 12.900 ;
        RECT 8.700 12.750 9.750 17.250 ;
        RECT 11.100 14.700 12.900 16.500 ;
        RECT 10.650 12.750 12.750 14.700 ;
        RECT 1.500 9.900 7.800 10.800 ;
        RECT 1.500 8.100 2.700 9.900 ;
        RECT 12.900 9.000 15.000 10.200 ;
        RECT 8.700 8.100 9.900 8.550 ;
        RECT 12.900 8.100 17.700 9.000 ;
        RECT 0.900 2.100 2.700 8.100 ;
        RECT 8.400 2.100 10.200 8.100 ;
        RECT 15.900 2.100 17.700 8.100 ;
      LAYER metal2 ;
        RECT 3.300 22.800 5.400 24.900 ;
        RECT 12.900 24.000 15.000 26.100 ;
        RECT 4.200 13.800 5.100 22.800 ;
        RECT 6.600 19.200 8.700 21.300 ;
        RECT 7.800 16.800 8.700 19.200 ;
        RECT 13.500 16.800 14.550 24.000 ;
        RECT 7.800 15.600 14.550 16.800 ;
        RECT 10.650 13.800 12.750 14.700 ;
        RECT 4.200 12.600 12.750 13.800 ;
        RECT 5.700 10.800 7.800 12.600 ;
        RECT 13.650 10.200 14.550 15.600 ;
        RECT 12.900 8.100 15.000 10.200 ;
  END
END XOR2X1
END LIBRARY
