magic
tech scmos
magscale 1 2
timestamp 1728340007
<< nwell >>
rect -13 134 252 252
rect -13 132 52 134
<< ntransistor >>
rect 21 14 25 54
rect 41 14 45 34
rect 53 14 57 34
rect 73 14 77 34
rect 83 14 87 34
rect 105 14 109 34
rect 149 14 153 34
rect 159 14 163 34
rect 179 14 183 34
rect 189 14 193 34
rect 209 14 213 54
<< ptransistor >>
rect 21 146 25 226
rect 41 186 45 226
rect 53 186 57 226
rect 73 186 77 226
rect 85 186 89 226
rect 105 186 109 226
rect 150 186 154 226
rect 159 186 163 226
rect 179 206 183 226
rect 189 206 193 226
rect 209 146 213 226
<< ndiffusion >>
rect 19 14 21 54
rect 25 34 36 54
rect 198 34 209 54
rect 25 14 27 34
rect 39 14 41 34
rect 45 14 53 34
rect 57 14 59 34
rect 71 14 73 34
rect 77 14 83 34
rect 87 14 89 34
rect 101 14 105 34
rect 109 14 111 34
rect 147 14 149 34
rect 153 14 159 34
rect 163 14 165 34
rect 177 14 179 34
rect 183 14 189 34
rect 193 14 195 34
rect 207 14 209 34
rect 213 14 215 54
<< pdiffusion >>
rect 19 146 21 226
rect 25 186 27 226
rect 39 186 41 226
rect 45 186 53 226
rect 57 186 59 226
rect 71 186 73 226
rect 77 186 85 226
rect 89 186 91 226
rect 103 186 105 226
rect 109 186 111 226
rect 148 186 150 226
rect 154 186 159 226
rect 163 206 165 226
rect 177 206 179 226
rect 183 206 189 226
rect 193 206 195 226
rect 207 206 209 226
rect 163 186 173 206
rect 25 146 36 186
rect 198 146 209 206
rect 213 146 215 226
<< ndcontact >>
rect 7 14 19 54
rect 27 14 39 34
rect 59 14 71 34
rect 89 14 101 34
rect 111 14 123 34
rect 135 14 147 34
rect 165 14 177 34
rect 195 14 207 34
rect 215 14 227 54
<< pdcontact >>
rect 7 146 19 226
rect 27 186 39 226
rect 59 186 71 226
rect 91 186 103 226
rect 111 186 123 226
rect 136 186 148 226
rect 165 206 177 226
rect 195 206 207 226
rect 215 146 227 226
<< psubstratepcontact >>
rect -6 -6 246 6
<< nsubstratencontact >>
rect -6 234 246 246
<< polysilicon >>
rect 21 226 25 230
rect 41 226 45 230
rect 53 226 57 230
rect 73 226 77 230
rect 85 226 89 230
rect 105 226 109 230
rect 150 226 154 230
rect 159 226 163 230
rect 179 226 183 230
rect 189 226 193 230
rect 209 226 213 230
rect 21 137 25 146
rect 12 131 25 137
rect 12 76 16 131
rect 41 123 45 186
rect 53 142 57 186
rect 73 180 77 186
rect 85 180 89 186
rect 65 130 77 134
rect 36 111 45 123
rect 12 64 20 76
rect 21 54 25 64
rect 41 34 45 111
rect 53 34 57 60
rect 73 34 77 130
rect 85 54 89 168
rect 105 128 109 186
rect 150 182 154 186
rect 83 52 89 54
rect 83 40 85 52
rect 83 34 87 40
rect 105 34 109 116
rect 117 180 154 182
rect 129 178 154 180
rect 159 174 163 186
rect 117 42 121 168
rect 157 167 163 174
rect 135 50 139 148
rect 157 70 161 167
rect 179 160 183 206
rect 181 148 183 160
rect 189 139 193 206
rect 159 60 161 70
rect 181 134 193 139
rect 181 81 185 134
rect 159 58 183 60
rect 147 54 183 58
rect 135 46 163 50
rect 117 38 153 42
rect 149 34 153 38
rect 159 34 163 46
rect 179 34 183 54
rect 189 34 193 69
rect 209 54 213 146
rect 21 10 25 14
rect 41 10 45 14
rect 53 10 57 14
rect 73 10 77 14
rect 83 10 87 14
rect 105 10 109 14
rect 149 10 153 14
rect 159 10 163 14
rect 179 10 183 14
rect 189 10 193 14
rect 209 10 213 14
<< polycontact >>
rect 65 168 77 180
rect 85 168 97 180
rect 53 130 65 142
rect 24 111 36 123
rect 20 64 32 76
rect 53 60 65 72
rect 97 116 109 128
rect 85 40 97 52
rect 117 168 129 180
rect 135 148 147 160
rect 169 148 181 160
rect 147 58 159 70
rect 197 112 209 124
rect 181 69 193 81
<< metal1 >>
rect -6 246 246 248
rect -6 232 246 234
rect 27 226 39 232
rect 91 226 103 232
rect 136 226 148 232
rect 195 226 207 232
rect 47 186 59 197
rect 165 186 177 206
rect 47 182 58 186
rect 111 180 123 186
rect 97 168 117 180
rect 65 162 77 168
rect 147 148 169 160
rect 7 142 19 146
rect 135 142 141 148
rect 7 134 53 142
rect 7 54 13 134
rect 65 134 141 142
rect 58 116 97 124
rect 177 112 197 120
rect 32 74 64 76
rect 215 83 223 146
rect 78 74 103 76
rect 32 72 103 74
rect 32 68 53 72
rect 65 69 103 72
rect 117 70 159 76
rect 117 69 147 70
rect 65 68 147 69
rect 193 69 203 81
rect 217 69 223 83
rect 215 54 223 69
rect 97 40 119 48
rect 47 34 58 40
rect 111 34 119 40
rect 47 27 59 34
rect 163 28 165 34
rect 27 8 39 14
rect 89 8 101 14
rect 135 8 147 14
rect 195 8 207 14
rect -6 6 246 8
rect -6 -8 246 -6
<< m2contact >>
rect 44 168 58 182
rect 163 172 177 186
rect 64 148 78 162
rect 23 97 37 111
rect 44 110 58 124
rect 163 110 177 124
rect 64 74 78 88
rect 103 69 117 83
rect 203 69 217 83
rect 44 40 58 54
rect 163 34 177 48
<< metal2 >>
rect 48 124 55 168
rect 23 83 37 97
rect 48 54 55 110
rect 68 88 76 148
rect 166 124 174 172
rect 103 83 117 97
rect 166 48 174 110
rect 203 83 217 97
<< m1p >>
rect -6 232 246 248
rect -6 -8 246 8
<< m2p >>
rect 23 83 37 97
rect 103 83 117 97
rect 203 83 217 97
<< labels >>
rlabel metal1 -6 -8 246 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 -6 232 246 248 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal2 23 83 37 97 0 D
port 0 nsew signal input
rlabel metal2 103 83 117 97 0 CLK
port 1 nsew clock input
rlabel metal2 203 83 217 97 0 Q
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 240 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
