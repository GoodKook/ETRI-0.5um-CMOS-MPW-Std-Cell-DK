magic
tech scmos
magscale 1 6
timestamp 1727178243
<< checkpaint >>
rect 8700 8700 29300 29300
<< metal1 >>
rect 28080 28027 29160 28040
rect 28080 28009 28941 28027
rect 28959 28009 28977 28027
rect 28995 28009 29013 28027
rect 29031 28009 29049 28027
rect 29067 28009 29085 28027
rect 29103 28009 29121 28027
rect 29139 28009 29160 28027
rect 28080 27991 29160 28009
rect 28080 27973 28941 27991
rect 28959 27973 28977 27991
rect 28995 27973 29013 27991
rect 29031 27973 29049 27991
rect 29067 27973 29085 27991
rect 29103 27973 29121 27991
rect 29139 27973 29160 27991
rect 28080 27955 29160 27973
rect 28080 27937 28941 27955
rect 28959 27937 28977 27955
rect 28995 27937 29013 27955
rect 29031 27937 29049 27955
rect 29067 27937 29085 27955
rect 29103 27937 29121 27955
rect 29139 27937 29160 27955
rect 28080 27919 29160 27937
rect 28080 27901 28941 27919
rect 28959 27901 28977 27919
rect 28995 27901 29013 27919
rect 29031 27901 29049 27919
rect 29067 27901 29085 27919
rect 29103 27901 29121 27919
rect 29139 27901 29160 27919
rect 28080 27883 29160 27901
rect 28080 27865 28941 27883
rect 28959 27865 28977 27883
rect 28995 27865 29013 27883
rect 29031 27865 29049 27883
rect 29067 27865 29085 27883
rect 29103 27865 29121 27883
rect 29139 27865 29160 27883
rect 28080 27847 29160 27865
rect 28080 27829 28941 27847
rect 28959 27829 28977 27847
rect 28995 27829 29013 27847
rect 29031 27829 29049 27847
rect 29067 27829 29085 27847
rect 29103 27829 29121 27847
rect 29139 27829 29160 27847
rect 28080 27811 29160 27829
rect 28080 27793 28941 27811
rect 28959 27793 28977 27811
rect 28995 27793 29013 27811
rect 29031 27793 29049 27811
rect 29067 27793 29085 27811
rect 29103 27793 29121 27811
rect 29139 27793 29160 27811
rect 8840 27757 9800 27780
rect 8840 27739 8861 27757
rect 8879 27739 8897 27757
rect 8915 27739 8933 27757
rect 8951 27739 8969 27757
rect 8987 27739 9005 27757
rect 9023 27739 9041 27757
rect 9059 27739 9800 27757
rect 8840 27721 9800 27739
rect 8840 27703 8861 27721
rect 8879 27703 8897 27721
rect 8915 27703 8933 27721
rect 8951 27703 8969 27721
rect 8987 27703 9005 27721
rect 9023 27703 9041 27721
rect 9059 27703 9800 27721
rect 8840 27685 9800 27703
rect 8840 27667 8861 27685
rect 8879 27667 8897 27685
rect 8915 27667 8933 27685
rect 8951 27667 8969 27685
rect 8987 27667 9005 27685
rect 9023 27667 9041 27685
rect 9059 27667 9800 27685
rect 8840 27649 9800 27667
rect 8840 27631 8861 27649
rect 8879 27631 8897 27649
rect 8915 27631 8933 27649
rect 8951 27631 8969 27649
rect 8987 27631 9005 27649
rect 9023 27631 9041 27649
rect 9059 27631 9800 27649
rect 8840 27613 9800 27631
rect 8840 27595 8861 27613
rect 8879 27595 8897 27613
rect 8915 27595 8933 27613
rect 8951 27595 8969 27613
rect 8987 27595 9005 27613
rect 9023 27595 9041 27613
rect 9059 27595 9800 27613
rect 8840 27577 9800 27595
rect 8840 27559 8861 27577
rect 8879 27559 8897 27577
rect 8915 27559 8933 27577
rect 8951 27559 8969 27577
rect 8987 27559 9005 27577
rect 9023 27559 9041 27577
rect 9059 27559 9800 27577
rect 8840 27541 9800 27559
rect 8840 27523 8861 27541
rect 8879 27523 8897 27541
rect 8915 27523 8933 27541
rect 8951 27523 8969 27541
rect 8987 27523 9005 27541
rect 9023 27523 9041 27541
rect 9059 27523 9800 27541
rect 8840 27505 9800 27523
rect 8840 27487 8861 27505
rect 8879 27487 8897 27505
rect 8915 27487 8933 27505
rect 8951 27487 8969 27505
rect 8987 27487 9005 27505
rect 9023 27487 9041 27505
rect 9059 27487 9800 27505
rect 8840 27469 9800 27487
rect 8840 27451 8861 27469
rect 8879 27451 8897 27469
rect 8915 27451 8933 27469
rect 8951 27451 8969 27469
rect 8987 27451 9005 27469
rect 9023 27451 9041 27469
rect 9059 27451 9800 27469
rect 8840 27433 9800 27451
rect 8840 27415 8861 27433
rect 8879 27415 8897 27433
rect 8915 27415 8933 27433
rect 8951 27415 8969 27433
rect 8987 27415 9005 27433
rect 9023 27415 9041 27433
rect 9059 27415 9800 27433
rect 8840 27397 9800 27415
rect 8840 27379 8861 27397
rect 8879 27379 8897 27397
rect 8915 27379 8933 27397
rect 8951 27379 8969 27397
rect 8987 27379 9005 27397
rect 9023 27379 9041 27397
rect 9059 27379 9800 27397
rect 8840 27361 9800 27379
rect 8840 27343 8861 27361
rect 8879 27343 8897 27361
rect 8915 27343 8933 27361
rect 8951 27343 8969 27361
rect 8987 27343 9005 27361
rect 9023 27343 9041 27361
rect 9059 27343 9800 27361
rect 8840 27325 9800 27343
rect 8840 27307 8861 27325
rect 8879 27307 8897 27325
rect 8915 27307 8933 27325
rect 8951 27307 8969 27325
rect 8987 27307 9005 27325
rect 9023 27307 9041 27325
rect 9059 27307 9800 27325
rect 8840 27289 9800 27307
rect 8840 27271 8861 27289
rect 8879 27271 8897 27289
rect 8915 27271 8933 27289
rect 8951 27271 8969 27289
rect 8987 27271 9005 27289
rect 9023 27271 9041 27289
rect 9059 27271 9800 27289
rect 8840 27253 9800 27271
rect 8840 27235 8861 27253
rect 8879 27235 8897 27253
rect 8915 27235 8933 27253
rect 8951 27235 8969 27253
rect 8987 27235 9005 27253
rect 9023 27235 9041 27253
rect 9059 27235 9800 27253
rect 8840 27217 9800 27235
rect 8840 27199 8861 27217
rect 8879 27199 8897 27217
rect 8915 27199 8933 27217
rect 8951 27199 8969 27217
rect 8987 27199 9005 27217
rect 9023 27199 9041 27217
rect 9059 27199 9800 27217
rect 8840 27181 9800 27199
rect 8840 27163 8861 27181
rect 8879 27163 8897 27181
rect 8915 27163 8933 27181
rect 8951 27163 8969 27181
rect 8987 27163 9005 27181
rect 9023 27163 9041 27181
rect 9059 27163 9800 27181
rect 8840 27145 9800 27163
rect 8840 27127 8861 27145
rect 8879 27127 8897 27145
rect 8915 27127 8933 27145
rect 8951 27127 8969 27145
rect 8987 27127 9005 27145
rect 9023 27127 9041 27145
rect 9059 27127 9800 27145
rect 8840 27109 9800 27127
rect 8840 27091 8861 27109
rect 8879 27091 8897 27109
rect 8915 27091 8933 27109
rect 8951 27091 8969 27109
rect 8987 27091 9005 27109
rect 9023 27091 9041 27109
rect 9059 27091 9800 27109
rect 8840 27073 9800 27091
rect 8840 27055 8861 27073
rect 8879 27055 8897 27073
rect 8915 27055 8933 27073
rect 8951 27055 8969 27073
rect 8987 27055 9005 27073
rect 9023 27055 9041 27073
rect 9059 27055 9800 27073
rect 8840 27037 9800 27055
rect 8840 27019 8861 27037
rect 8879 27019 8897 27037
rect 8915 27019 8933 27037
rect 8951 27019 8969 27037
rect 8987 27019 9005 27037
rect 9023 27019 9041 27037
rect 9059 27019 9800 27037
rect 8840 27001 9800 27019
rect 8840 26983 8861 27001
rect 8879 26983 8897 27001
rect 8915 26983 8933 27001
rect 8951 26983 8969 27001
rect 8987 26983 9005 27001
rect 9023 26983 9041 27001
rect 9059 26983 9800 27001
rect 8840 26965 9800 26983
rect 8840 26947 8861 26965
rect 8879 26947 8897 26965
rect 8915 26947 8933 26965
rect 8951 26947 8969 26965
rect 8987 26947 9005 26965
rect 9023 26947 9041 26965
rect 9059 26947 9800 26965
rect 8840 26929 9800 26947
rect 8840 26911 8861 26929
rect 8879 26911 8897 26929
rect 8915 26911 8933 26929
rect 8951 26911 8969 26929
rect 8987 26911 9005 26929
rect 9023 26911 9041 26929
rect 9059 26911 9800 26929
rect 8840 26893 9800 26911
rect 8840 26875 8861 26893
rect 8879 26875 8897 26893
rect 8915 26875 8933 26893
rect 8951 26875 8969 26893
rect 8987 26875 9005 26893
rect 9023 26875 9041 26893
rect 9059 26875 9800 26893
rect 8840 26857 9800 26875
rect 8840 26839 8861 26857
rect 8879 26839 8897 26857
rect 8915 26839 8933 26857
rect 8951 26839 8969 26857
rect 8987 26839 9005 26857
rect 9023 26839 9041 26857
rect 9059 26839 9800 26857
rect 8840 26821 9800 26839
rect 8840 26803 8861 26821
rect 8879 26803 8897 26821
rect 8915 26803 8933 26821
rect 8951 26803 8969 26821
rect 8987 26803 9005 26821
rect 9023 26803 9041 26821
rect 9059 26803 9800 26821
rect 8840 26785 9800 26803
rect 8840 26767 8861 26785
rect 8879 26767 8897 26785
rect 8915 26767 8933 26785
rect 8951 26767 8969 26785
rect 8987 26767 9005 26785
rect 9023 26767 9041 26785
rect 9059 26767 9800 26785
rect 8840 26749 9800 26767
rect 8840 26731 8861 26749
rect 8879 26731 8897 26749
rect 8915 26731 8933 26749
rect 8951 26731 8969 26749
rect 8987 26731 9005 26749
rect 9023 26731 9041 26749
rect 9059 26731 9800 26749
rect 8840 26713 9800 26731
rect 8840 26695 8861 26713
rect 8879 26695 8897 26713
rect 8915 26695 8933 26713
rect 8951 26695 8969 26713
rect 8987 26695 9005 26713
rect 9023 26695 9041 26713
rect 9059 26695 9800 26713
rect 8840 26677 9800 26695
rect 8840 26659 8861 26677
rect 8879 26659 8897 26677
rect 8915 26659 8933 26677
rect 8951 26659 8969 26677
rect 8987 26659 9005 26677
rect 9023 26659 9041 26677
rect 9059 26659 9800 26677
rect 8840 26641 9800 26659
rect 8840 26623 8861 26641
rect 8879 26623 8897 26641
rect 8915 26623 8933 26641
rect 8951 26623 8969 26641
rect 8987 26623 9005 26641
rect 9023 26623 9041 26641
rect 9059 26623 9800 26641
rect 8840 26605 9800 26623
rect 8840 26587 8861 26605
rect 8879 26587 8897 26605
rect 8915 26587 8933 26605
rect 8951 26587 8969 26605
rect 8987 26587 9005 26605
rect 9023 26587 9041 26605
rect 9059 26587 9800 26605
rect 8840 26569 9800 26587
rect 8840 26551 8861 26569
rect 8879 26551 8897 26569
rect 8915 26551 8933 26569
rect 8951 26551 8969 26569
rect 8987 26551 9005 26569
rect 9023 26551 9041 26569
rect 9059 26551 9800 26569
rect 8840 26533 9800 26551
rect 8840 26515 8861 26533
rect 8879 26515 8897 26533
rect 8915 26515 8933 26533
rect 8951 26515 8969 26533
rect 8987 26515 9005 26533
rect 9023 26515 9041 26533
rect 9059 26515 9800 26533
rect 8840 26497 9800 26515
rect 8840 26479 8861 26497
rect 8879 26479 8897 26497
rect 8915 26479 8933 26497
rect 8951 26479 8969 26497
rect 8987 26479 9005 26497
rect 9023 26479 9041 26497
rect 9059 26479 9800 26497
rect 8840 26461 9800 26479
rect 8840 26443 8861 26461
rect 8879 26443 8897 26461
rect 8915 26443 8933 26461
rect 8951 26443 8969 26461
rect 8987 26443 9005 26461
rect 9023 26443 9041 26461
rect 9059 26443 9800 26461
rect 8840 26420 9800 26443
rect 28080 27775 29160 27793
rect 28080 27757 28941 27775
rect 28959 27757 28977 27775
rect 28995 27757 29013 27775
rect 29031 27757 29049 27775
rect 29067 27757 29085 27775
rect 29103 27757 29121 27775
rect 29139 27757 29160 27775
rect 28080 27739 29160 27757
rect 28080 27721 28941 27739
rect 28959 27721 28977 27739
rect 28995 27721 29013 27739
rect 29031 27721 29049 27739
rect 29067 27721 29085 27739
rect 29103 27721 29121 27739
rect 29139 27721 29160 27739
rect 28080 27703 29160 27721
rect 28080 27685 28941 27703
rect 28959 27685 28977 27703
rect 28995 27685 29013 27703
rect 29031 27685 29049 27703
rect 29067 27685 29085 27703
rect 29103 27685 29121 27703
rect 29139 27685 29160 27703
rect 28080 27667 29160 27685
rect 28080 27649 28941 27667
rect 28959 27649 28977 27667
rect 28995 27649 29013 27667
rect 29031 27649 29049 27667
rect 29067 27649 29085 27667
rect 29103 27649 29121 27667
rect 29139 27649 29160 27667
rect 28080 27631 29160 27649
rect 28080 27613 28941 27631
rect 28959 27613 28977 27631
rect 28995 27613 29013 27631
rect 29031 27613 29049 27631
rect 29067 27613 29085 27631
rect 29103 27613 29121 27631
rect 29139 27613 29160 27631
rect 28080 27595 29160 27613
rect 28080 27577 28941 27595
rect 28959 27577 28977 27595
rect 28995 27577 29013 27595
rect 29031 27577 29049 27595
rect 29067 27577 29085 27595
rect 29103 27577 29121 27595
rect 29139 27577 29160 27595
rect 28080 27559 29160 27577
rect 28080 27541 28941 27559
rect 28959 27541 28977 27559
rect 28995 27541 29013 27559
rect 29031 27541 29049 27559
rect 29067 27541 29085 27559
rect 29103 27541 29121 27559
rect 29139 27541 29160 27559
rect 28080 27523 29160 27541
rect 28080 27505 28941 27523
rect 28959 27505 28977 27523
rect 28995 27505 29013 27523
rect 29031 27505 29049 27523
rect 29067 27505 29085 27523
rect 29103 27505 29121 27523
rect 29139 27505 29160 27523
rect 28080 27487 29160 27505
rect 28080 27469 28941 27487
rect 28959 27469 28977 27487
rect 28995 27469 29013 27487
rect 29031 27469 29049 27487
rect 29067 27469 29085 27487
rect 29103 27469 29121 27487
rect 29139 27469 29160 27487
rect 28080 27451 29160 27469
rect 28080 27433 28941 27451
rect 28959 27433 28977 27451
rect 28995 27433 29013 27451
rect 29031 27433 29049 27451
rect 29067 27433 29085 27451
rect 29103 27433 29121 27451
rect 29139 27433 29160 27451
rect 28080 27415 29160 27433
rect 28080 27397 28941 27415
rect 28959 27397 28977 27415
rect 28995 27397 29013 27415
rect 29031 27397 29049 27415
rect 29067 27397 29085 27415
rect 29103 27397 29121 27415
rect 29139 27397 29160 27415
rect 28080 27379 29160 27397
rect 28080 27361 28941 27379
rect 28959 27361 28977 27379
rect 28995 27361 29013 27379
rect 29031 27361 29049 27379
rect 29067 27361 29085 27379
rect 29103 27361 29121 27379
rect 29139 27361 29160 27379
rect 28080 27343 29160 27361
rect 28080 27325 28941 27343
rect 28959 27325 28977 27343
rect 28995 27325 29013 27343
rect 29031 27325 29049 27343
rect 29067 27325 29085 27343
rect 29103 27325 29121 27343
rect 29139 27325 29160 27343
rect 28080 27307 29160 27325
rect 28080 27289 28941 27307
rect 28959 27289 28977 27307
rect 28995 27289 29013 27307
rect 29031 27289 29049 27307
rect 29067 27289 29085 27307
rect 29103 27289 29121 27307
rect 29139 27289 29160 27307
rect 28080 27271 29160 27289
rect 28080 27253 28941 27271
rect 28959 27253 28977 27271
rect 28995 27253 29013 27271
rect 29031 27253 29049 27271
rect 29067 27253 29085 27271
rect 29103 27253 29121 27271
rect 29139 27253 29160 27271
rect 28080 27235 29160 27253
rect 28080 27217 28941 27235
rect 28959 27217 28977 27235
rect 28995 27217 29013 27235
rect 29031 27217 29049 27235
rect 29067 27217 29085 27235
rect 29103 27217 29121 27235
rect 29139 27217 29160 27235
rect 28080 27199 29160 27217
rect 28080 27181 28941 27199
rect 28959 27181 28977 27199
rect 28995 27181 29013 27199
rect 29031 27181 29049 27199
rect 29067 27181 29085 27199
rect 29103 27181 29121 27199
rect 29139 27181 29160 27199
rect 28080 27163 29160 27181
rect 28080 27145 28941 27163
rect 28959 27145 28977 27163
rect 28995 27145 29013 27163
rect 29031 27145 29049 27163
rect 29067 27145 29085 27163
rect 29103 27145 29121 27163
rect 29139 27145 29160 27163
rect 28080 27127 29160 27145
rect 28080 27109 28941 27127
rect 28959 27109 28977 27127
rect 28995 27109 29013 27127
rect 29031 27109 29049 27127
rect 29067 27109 29085 27127
rect 29103 27109 29121 27127
rect 29139 27109 29160 27127
rect 28080 27091 29160 27109
rect 28080 27073 28941 27091
rect 28959 27073 28977 27091
rect 28995 27073 29013 27091
rect 29031 27073 29049 27091
rect 29067 27073 29085 27091
rect 29103 27073 29121 27091
rect 29139 27073 29160 27091
rect 28080 27055 29160 27073
rect 28080 27037 28941 27055
rect 28959 27037 28977 27055
rect 28995 27037 29013 27055
rect 29031 27037 29049 27055
rect 29067 27037 29085 27055
rect 29103 27037 29121 27055
rect 29139 27037 29160 27055
rect 28080 27019 29160 27037
rect 28080 27001 28941 27019
rect 28959 27001 28977 27019
rect 28995 27001 29013 27019
rect 29031 27001 29049 27019
rect 29067 27001 29085 27019
rect 29103 27001 29121 27019
rect 29139 27001 29160 27019
rect 28080 26983 29160 27001
rect 28080 26965 28941 26983
rect 28959 26965 28977 26983
rect 28995 26965 29013 26983
rect 29031 26965 29049 26983
rect 29067 26965 29085 26983
rect 29103 26965 29121 26983
rect 29139 26965 29160 26983
rect 28080 26947 29160 26965
rect 28080 26929 28941 26947
rect 28959 26929 28977 26947
rect 28995 26929 29013 26947
rect 29031 26929 29049 26947
rect 29067 26929 29085 26947
rect 29103 26929 29121 26947
rect 29139 26929 29160 26947
rect 28080 26911 29160 26929
rect 28080 26893 28941 26911
rect 28959 26893 28977 26911
rect 28995 26893 29013 26911
rect 29031 26893 29049 26911
rect 29067 26893 29085 26911
rect 29103 26893 29121 26911
rect 29139 26893 29160 26911
rect 28080 26875 29160 26893
rect 28080 26857 28941 26875
rect 28959 26857 28977 26875
rect 28995 26857 29013 26875
rect 29031 26857 29049 26875
rect 29067 26857 29085 26875
rect 29103 26857 29121 26875
rect 29139 26857 29160 26875
rect 28080 26839 29160 26857
rect 28080 26821 28941 26839
rect 28959 26821 28977 26839
rect 28995 26821 29013 26839
rect 29031 26821 29049 26839
rect 29067 26821 29085 26839
rect 29103 26821 29121 26839
rect 29139 26821 29160 26839
rect 28080 26803 29160 26821
rect 28080 26785 28941 26803
rect 28959 26785 28977 26803
rect 28995 26785 29013 26803
rect 29031 26785 29049 26803
rect 29067 26785 29085 26803
rect 29103 26785 29121 26803
rect 29139 26785 29160 26803
rect 28080 26767 29160 26785
rect 28080 26749 28941 26767
rect 28959 26749 28977 26767
rect 28995 26749 29013 26767
rect 29031 26749 29049 26767
rect 29067 26749 29085 26767
rect 29103 26749 29121 26767
rect 29139 26749 29160 26767
rect 28080 26731 29160 26749
rect 28080 26713 28941 26731
rect 28959 26713 28977 26731
rect 28995 26713 29013 26731
rect 29031 26713 29049 26731
rect 29067 26713 29085 26731
rect 29103 26713 29121 26731
rect 29139 26713 29160 26731
rect 28080 26695 29160 26713
rect 28080 26677 28941 26695
rect 28959 26677 28977 26695
rect 28995 26677 29013 26695
rect 29031 26677 29049 26695
rect 29067 26677 29085 26695
rect 29103 26677 29121 26695
rect 29139 26677 29160 26695
rect 28080 26659 29160 26677
rect 28080 26641 28941 26659
rect 28959 26641 28977 26659
rect 28995 26641 29013 26659
rect 29031 26641 29049 26659
rect 29067 26641 29085 26659
rect 29103 26641 29121 26659
rect 29139 26641 29160 26659
rect 28080 26623 29160 26641
rect 28080 26605 28941 26623
rect 28959 26605 28977 26623
rect 28995 26605 29013 26623
rect 29031 26605 29049 26623
rect 29067 26605 29085 26623
rect 29103 26605 29121 26623
rect 29139 26605 29160 26623
rect 28080 26587 29160 26605
rect 28080 26569 28941 26587
rect 28959 26569 28977 26587
rect 28995 26569 29013 26587
rect 29031 26569 29049 26587
rect 29067 26569 29085 26587
rect 29103 26569 29121 26587
rect 29139 26569 29160 26587
rect 28080 26551 29160 26569
rect 28080 26533 28941 26551
rect 28959 26533 28977 26551
rect 28995 26533 29013 26551
rect 29031 26533 29049 26551
rect 29067 26533 29085 26551
rect 29103 26533 29121 26551
rect 29139 26533 29160 26551
rect 28080 26515 29160 26533
rect 28080 26497 28941 26515
rect 28959 26497 28977 26515
rect 28995 26497 29013 26515
rect 29031 26497 29049 26515
rect 29067 26497 29085 26515
rect 29103 26497 29121 26515
rect 29139 26497 29160 26515
rect 28080 26479 29160 26497
rect 28080 26461 28941 26479
rect 28959 26461 28977 26479
rect 28995 26461 29013 26479
rect 29031 26461 29049 26479
rect 29067 26461 29085 26479
rect 29103 26461 29121 26479
rect 29139 26461 29160 26479
rect 28080 26443 29160 26461
rect 28080 26425 28941 26443
rect 28959 26425 28977 26443
rect 28995 26425 29013 26443
rect 29031 26425 29049 26443
rect 29067 26425 29085 26443
rect 29103 26425 29121 26443
rect 29139 26425 29160 26443
rect 28080 26407 29160 26425
rect 28080 26389 28941 26407
rect 28959 26389 28977 26407
rect 28995 26389 29013 26407
rect 29031 26389 29049 26407
rect 29067 26389 29085 26407
rect 29103 26389 29121 26407
rect 29139 26389 29160 26407
rect 28080 26371 29160 26389
rect 28080 26353 28941 26371
rect 28959 26353 28977 26371
rect 28995 26353 29013 26371
rect 29031 26353 29049 26371
rect 29067 26353 29085 26371
rect 29103 26353 29121 26371
rect 29139 26353 29160 26371
rect 28080 26335 29160 26353
rect 28080 26317 28941 26335
rect 28959 26317 28977 26335
rect 28995 26317 29013 26335
rect 29031 26317 29049 26335
rect 29067 26317 29085 26335
rect 29103 26317 29121 26335
rect 29139 26317 29160 26335
rect 28080 26299 29160 26317
rect 28080 26281 28941 26299
rect 28959 26281 28977 26299
rect 28995 26281 29013 26299
rect 29031 26281 29049 26299
rect 29067 26281 29085 26299
rect 29103 26281 29121 26299
rect 29139 26281 29160 26299
rect 28080 26263 29160 26281
rect 28080 26245 28941 26263
rect 28959 26245 28977 26263
rect 28995 26245 29013 26263
rect 29031 26245 29049 26263
rect 29067 26245 29085 26263
rect 29103 26245 29121 26263
rect 29139 26245 29160 26263
rect 28080 26227 29160 26245
rect 28080 26209 28941 26227
rect 28959 26209 28977 26227
rect 28995 26209 29013 26227
rect 29031 26209 29049 26227
rect 29067 26209 29085 26227
rect 29103 26209 29121 26227
rect 29139 26209 29160 26227
rect 28080 26191 29160 26209
rect 28080 26173 28941 26191
rect 28959 26173 28977 26191
rect 28995 26173 29013 26191
rect 29031 26173 29049 26191
rect 29067 26173 29085 26191
rect 29103 26173 29121 26191
rect 29139 26173 29160 26191
rect 28080 26160 29160 26173
rect 8840 11547 9800 11560
rect 8840 11529 8861 11547
rect 8879 11529 8897 11547
rect 8915 11529 8933 11547
rect 8951 11529 8969 11547
rect 8987 11529 9005 11547
rect 9023 11529 9041 11547
rect 9059 11529 9800 11547
rect 8840 11511 9800 11529
rect 8840 11493 8861 11511
rect 8879 11493 8897 11511
rect 8915 11493 8933 11511
rect 8951 11493 8969 11511
rect 8987 11493 9005 11511
rect 9023 11493 9041 11511
rect 9059 11493 9800 11511
rect 8840 11475 9800 11493
rect 8840 11457 8861 11475
rect 8879 11457 8897 11475
rect 8915 11457 8933 11475
rect 8951 11457 8969 11475
rect 8987 11457 9005 11475
rect 9023 11457 9041 11475
rect 9059 11457 9800 11475
rect 8840 11439 9800 11457
rect 8840 11421 8861 11439
rect 8879 11421 8897 11439
rect 8915 11421 8933 11439
rect 8951 11421 8969 11439
rect 8987 11421 9005 11439
rect 9023 11421 9041 11439
rect 9059 11421 9800 11439
rect 8840 11403 9800 11421
rect 8840 11385 8861 11403
rect 8879 11385 8897 11403
rect 8915 11385 8933 11403
rect 8951 11385 8969 11403
rect 8987 11385 9005 11403
rect 9023 11385 9041 11403
rect 9059 11385 9800 11403
rect 8840 11367 9800 11385
rect 8840 11349 8861 11367
rect 8879 11349 8897 11367
rect 8915 11349 8933 11367
rect 8951 11349 8969 11367
rect 8987 11349 9005 11367
rect 9023 11349 9041 11367
rect 9059 11349 9800 11367
rect 8840 11331 9800 11349
rect 8840 11313 8861 11331
rect 8879 11313 8897 11331
rect 8915 11313 8933 11331
rect 8951 11313 8969 11331
rect 8987 11313 9005 11331
rect 9023 11313 9041 11331
rect 9059 11313 9800 11331
rect 8840 11295 9800 11313
rect 8840 11277 8861 11295
rect 8879 11277 8897 11295
rect 8915 11277 8933 11295
rect 8951 11277 8969 11295
rect 8987 11277 9005 11295
rect 9023 11277 9041 11295
rect 9059 11277 9800 11295
rect 8840 11259 9800 11277
rect 8840 11241 8861 11259
rect 8879 11241 8897 11259
rect 8915 11241 8933 11259
rect 8951 11241 8969 11259
rect 8987 11241 9005 11259
rect 9023 11241 9041 11259
rect 9059 11241 9800 11259
rect 8840 11223 9800 11241
rect 8840 11205 8861 11223
rect 8879 11205 8897 11223
rect 8915 11205 8933 11223
rect 8951 11205 8969 11223
rect 8987 11205 9005 11223
rect 9023 11205 9041 11223
rect 9059 11205 9800 11223
rect 8840 11187 9800 11205
rect 8840 11169 8861 11187
rect 8879 11169 8897 11187
rect 8915 11169 8933 11187
rect 8951 11169 8969 11187
rect 8987 11169 9005 11187
rect 9023 11169 9041 11187
rect 9059 11169 9800 11187
rect 8840 11151 9800 11169
rect 8840 11133 8861 11151
rect 8879 11133 8897 11151
rect 8915 11133 8933 11151
rect 8951 11133 8969 11151
rect 8987 11133 9005 11151
rect 9023 11133 9041 11151
rect 9059 11133 9800 11151
rect 8840 11115 9800 11133
rect 8840 11097 8861 11115
rect 8879 11097 8897 11115
rect 8915 11097 8933 11115
rect 8951 11097 8969 11115
rect 8987 11097 9005 11115
rect 9023 11097 9041 11115
rect 9059 11097 9800 11115
rect 8840 11079 9800 11097
rect 8840 11061 8861 11079
rect 8879 11061 8897 11079
rect 8915 11061 8933 11079
rect 8951 11061 8969 11079
rect 8987 11061 9005 11079
rect 9023 11061 9041 11079
rect 9059 11061 9800 11079
rect 8840 11043 9800 11061
rect 8840 11025 8861 11043
rect 8879 11025 8897 11043
rect 8915 11025 8933 11043
rect 8951 11025 8969 11043
rect 8987 11025 9005 11043
rect 9023 11025 9041 11043
rect 9059 11025 9800 11043
rect 8840 11007 9800 11025
rect 8840 10989 8861 11007
rect 8879 10989 8897 11007
rect 8915 10989 8933 11007
rect 8951 10989 8969 11007
rect 8987 10989 9005 11007
rect 9023 10989 9041 11007
rect 9059 10989 9800 11007
rect 8840 10971 9800 10989
rect 8840 10953 8861 10971
rect 8879 10953 8897 10971
rect 8915 10953 8933 10971
rect 8951 10953 8969 10971
rect 8987 10953 9005 10971
rect 9023 10953 9041 10971
rect 9059 10953 9800 10971
rect 8840 10935 9800 10953
rect 8840 10917 8861 10935
rect 8879 10917 8897 10935
rect 8915 10917 8933 10935
rect 8951 10917 8969 10935
rect 8987 10917 9005 10935
rect 9023 10917 9041 10935
rect 9059 10917 9800 10935
rect 8840 10899 9800 10917
rect 8840 10881 8861 10899
rect 8879 10881 8897 10899
rect 8915 10881 8933 10899
rect 8951 10881 8969 10899
rect 8987 10881 9005 10899
rect 9023 10881 9041 10899
rect 9059 10881 9800 10899
rect 8840 10863 9800 10881
rect 8840 10845 8861 10863
rect 8879 10845 8897 10863
rect 8915 10845 8933 10863
rect 8951 10845 8969 10863
rect 8987 10845 9005 10863
rect 9023 10845 9041 10863
rect 9059 10845 9800 10863
rect 8840 10827 9800 10845
rect 8840 10809 8861 10827
rect 8879 10809 8897 10827
rect 8915 10809 8933 10827
rect 8951 10809 8969 10827
rect 8987 10809 9005 10827
rect 9023 10809 9041 10827
rect 9059 10809 9800 10827
rect 8840 10791 9800 10809
rect 8840 10773 8861 10791
rect 8879 10773 8897 10791
rect 8915 10773 8933 10791
rect 8951 10773 8969 10791
rect 8987 10773 9005 10791
rect 9023 10773 9041 10791
rect 9059 10773 9800 10791
rect 8840 10755 9800 10773
rect 8840 10737 8861 10755
rect 8879 10737 8897 10755
rect 8915 10737 8933 10755
rect 8951 10737 8969 10755
rect 8987 10737 9005 10755
rect 9023 10737 9041 10755
rect 9059 10737 9800 10755
rect 8840 10719 9800 10737
rect 8840 10701 8861 10719
rect 8879 10701 8897 10719
rect 8915 10701 8933 10719
rect 8951 10701 8969 10719
rect 8987 10701 9005 10719
rect 9023 10701 9041 10719
rect 9059 10701 9800 10719
rect 8840 10683 9800 10701
rect 8840 10665 8861 10683
rect 8879 10665 8897 10683
rect 8915 10665 8933 10683
rect 8951 10665 8969 10683
rect 8987 10665 9005 10683
rect 9023 10665 9041 10683
rect 9059 10665 9800 10683
rect 8840 10647 9800 10665
rect 8840 10629 8861 10647
rect 8879 10629 8897 10647
rect 8915 10629 8933 10647
rect 8951 10629 8969 10647
rect 8987 10629 9005 10647
rect 9023 10629 9041 10647
rect 9059 10629 9800 10647
rect 8840 10611 9800 10629
rect 8840 10593 8861 10611
rect 8879 10593 8897 10611
rect 8915 10593 8933 10611
rect 8951 10593 8969 10611
rect 8987 10593 9005 10611
rect 9023 10593 9041 10611
rect 9059 10593 9800 10611
rect 8840 10575 9800 10593
rect 8840 10557 8861 10575
rect 8879 10557 8897 10575
rect 8915 10557 8933 10575
rect 8951 10557 8969 10575
rect 8987 10557 9005 10575
rect 9023 10557 9041 10575
rect 9059 10557 9800 10575
rect 8840 10539 9800 10557
rect 8840 10521 8861 10539
rect 8879 10521 8897 10539
rect 8915 10521 8933 10539
rect 8951 10521 8969 10539
rect 8987 10521 9005 10539
rect 9023 10521 9041 10539
rect 9059 10521 9800 10539
rect 8840 10503 9800 10521
rect 8840 10485 8861 10503
rect 8879 10485 8897 10503
rect 8915 10485 8933 10503
rect 8951 10485 8969 10503
rect 8987 10485 9005 10503
rect 9023 10485 9041 10503
rect 9059 10485 9800 10503
rect 8840 10467 9800 10485
rect 8840 10449 8861 10467
rect 8879 10449 8897 10467
rect 8915 10449 8933 10467
rect 8951 10449 8969 10467
rect 8987 10449 9005 10467
rect 9023 10449 9041 10467
rect 9059 10449 9800 10467
rect 8840 10431 9800 10449
rect 8840 10413 8861 10431
rect 8879 10413 8897 10431
rect 8915 10413 8933 10431
rect 8951 10413 8969 10431
rect 8987 10413 9005 10431
rect 9023 10413 9041 10431
rect 9059 10413 9800 10431
rect 8840 10395 9800 10413
rect 8840 10377 8861 10395
rect 8879 10377 8897 10395
rect 8915 10377 8933 10395
rect 8951 10377 8969 10395
rect 8987 10377 9005 10395
rect 9023 10377 9041 10395
rect 9059 10377 9800 10395
rect 8840 10359 9800 10377
rect 8840 10341 8861 10359
rect 8879 10341 8897 10359
rect 8915 10341 8933 10359
rect 8951 10341 8969 10359
rect 8987 10341 9005 10359
rect 9023 10341 9041 10359
rect 9059 10341 9800 10359
rect 8840 10323 9800 10341
rect 8840 10305 8861 10323
rect 8879 10305 8897 10323
rect 8915 10305 8933 10323
rect 8951 10305 8969 10323
rect 8987 10305 9005 10323
rect 9023 10305 9041 10323
rect 9059 10305 9800 10323
rect 8840 10287 9800 10305
rect 8840 10269 8861 10287
rect 8879 10269 8897 10287
rect 8915 10269 8933 10287
rect 8951 10269 8969 10287
rect 8987 10269 9005 10287
rect 9023 10269 9041 10287
rect 9059 10269 9800 10287
rect 8840 10251 9800 10269
rect 8840 10233 8861 10251
rect 8879 10233 8897 10251
rect 8915 10233 8933 10251
rect 8951 10233 8969 10251
rect 8987 10233 9005 10251
rect 9023 10233 9041 10251
rect 9059 10233 9800 10251
rect 8840 10220 9800 10233
<< m2contact >>
rect 28941 28009 28959 28027
rect 28977 28009 28995 28027
rect 29013 28009 29031 28027
rect 29049 28009 29067 28027
rect 29085 28009 29103 28027
rect 29121 28009 29139 28027
rect 28941 27973 28959 27991
rect 28977 27973 28995 27991
rect 29013 27973 29031 27991
rect 29049 27973 29067 27991
rect 29085 27973 29103 27991
rect 29121 27973 29139 27991
rect 28941 27937 28959 27955
rect 28977 27937 28995 27955
rect 29013 27937 29031 27955
rect 29049 27937 29067 27955
rect 29085 27937 29103 27955
rect 29121 27937 29139 27955
rect 28941 27901 28959 27919
rect 28977 27901 28995 27919
rect 29013 27901 29031 27919
rect 29049 27901 29067 27919
rect 29085 27901 29103 27919
rect 29121 27901 29139 27919
rect 28941 27865 28959 27883
rect 28977 27865 28995 27883
rect 29013 27865 29031 27883
rect 29049 27865 29067 27883
rect 29085 27865 29103 27883
rect 29121 27865 29139 27883
rect 28941 27829 28959 27847
rect 28977 27829 28995 27847
rect 29013 27829 29031 27847
rect 29049 27829 29067 27847
rect 29085 27829 29103 27847
rect 29121 27829 29139 27847
rect 28941 27793 28959 27811
rect 28977 27793 28995 27811
rect 29013 27793 29031 27811
rect 29049 27793 29067 27811
rect 29085 27793 29103 27811
rect 29121 27793 29139 27811
rect 8861 27739 8879 27757
rect 8897 27739 8915 27757
rect 8933 27739 8951 27757
rect 8969 27739 8987 27757
rect 9005 27739 9023 27757
rect 9041 27739 9059 27757
rect 8861 27703 8879 27721
rect 8897 27703 8915 27721
rect 8933 27703 8951 27721
rect 8969 27703 8987 27721
rect 9005 27703 9023 27721
rect 9041 27703 9059 27721
rect 8861 27667 8879 27685
rect 8897 27667 8915 27685
rect 8933 27667 8951 27685
rect 8969 27667 8987 27685
rect 9005 27667 9023 27685
rect 9041 27667 9059 27685
rect 8861 27631 8879 27649
rect 8897 27631 8915 27649
rect 8933 27631 8951 27649
rect 8969 27631 8987 27649
rect 9005 27631 9023 27649
rect 9041 27631 9059 27649
rect 8861 27595 8879 27613
rect 8897 27595 8915 27613
rect 8933 27595 8951 27613
rect 8969 27595 8987 27613
rect 9005 27595 9023 27613
rect 9041 27595 9059 27613
rect 8861 27559 8879 27577
rect 8897 27559 8915 27577
rect 8933 27559 8951 27577
rect 8969 27559 8987 27577
rect 9005 27559 9023 27577
rect 9041 27559 9059 27577
rect 8861 27523 8879 27541
rect 8897 27523 8915 27541
rect 8933 27523 8951 27541
rect 8969 27523 8987 27541
rect 9005 27523 9023 27541
rect 9041 27523 9059 27541
rect 8861 27487 8879 27505
rect 8897 27487 8915 27505
rect 8933 27487 8951 27505
rect 8969 27487 8987 27505
rect 9005 27487 9023 27505
rect 9041 27487 9059 27505
rect 8861 27451 8879 27469
rect 8897 27451 8915 27469
rect 8933 27451 8951 27469
rect 8969 27451 8987 27469
rect 9005 27451 9023 27469
rect 9041 27451 9059 27469
rect 8861 27415 8879 27433
rect 8897 27415 8915 27433
rect 8933 27415 8951 27433
rect 8969 27415 8987 27433
rect 9005 27415 9023 27433
rect 9041 27415 9059 27433
rect 8861 27379 8879 27397
rect 8897 27379 8915 27397
rect 8933 27379 8951 27397
rect 8969 27379 8987 27397
rect 9005 27379 9023 27397
rect 9041 27379 9059 27397
rect 8861 27343 8879 27361
rect 8897 27343 8915 27361
rect 8933 27343 8951 27361
rect 8969 27343 8987 27361
rect 9005 27343 9023 27361
rect 9041 27343 9059 27361
rect 8861 27307 8879 27325
rect 8897 27307 8915 27325
rect 8933 27307 8951 27325
rect 8969 27307 8987 27325
rect 9005 27307 9023 27325
rect 9041 27307 9059 27325
rect 8861 27271 8879 27289
rect 8897 27271 8915 27289
rect 8933 27271 8951 27289
rect 8969 27271 8987 27289
rect 9005 27271 9023 27289
rect 9041 27271 9059 27289
rect 8861 27235 8879 27253
rect 8897 27235 8915 27253
rect 8933 27235 8951 27253
rect 8969 27235 8987 27253
rect 9005 27235 9023 27253
rect 9041 27235 9059 27253
rect 8861 27199 8879 27217
rect 8897 27199 8915 27217
rect 8933 27199 8951 27217
rect 8969 27199 8987 27217
rect 9005 27199 9023 27217
rect 9041 27199 9059 27217
rect 8861 27163 8879 27181
rect 8897 27163 8915 27181
rect 8933 27163 8951 27181
rect 8969 27163 8987 27181
rect 9005 27163 9023 27181
rect 9041 27163 9059 27181
rect 8861 27127 8879 27145
rect 8897 27127 8915 27145
rect 8933 27127 8951 27145
rect 8969 27127 8987 27145
rect 9005 27127 9023 27145
rect 9041 27127 9059 27145
rect 8861 27091 8879 27109
rect 8897 27091 8915 27109
rect 8933 27091 8951 27109
rect 8969 27091 8987 27109
rect 9005 27091 9023 27109
rect 9041 27091 9059 27109
rect 8861 27055 8879 27073
rect 8897 27055 8915 27073
rect 8933 27055 8951 27073
rect 8969 27055 8987 27073
rect 9005 27055 9023 27073
rect 9041 27055 9059 27073
rect 8861 27019 8879 27037
rect 8897 27019 8915 27037
rect 8933 27019 8951 27037
rect 8969 27019 8987 27037
rect 9005 27019 9023 27037
rect 9041 27019 9059 27037
rect 8861 26983 8879 27001
rect 8897 26983 8915 27001
rect 8933 26983 8951 27001
rect 8969 26983 8987 27001
rect 9005 26983 9023 27001
rect 9041 26983 9059 27001
rect 8861 26947 8879 26965
rect 8897 26947 8915 26965
rect 8933 26947 8951 26965
rect 8969 26947 8987 26965
rect 9005 26947 9023 26965
rect 9041 26947 9059 26965
rect 8861 26911 8879 26929
rect 8897 26911 8915 26929
rect 8933 26911 8951 26929
rect 8969 26911 8987 26929
rect 9005 26911 9023 26929
rect 9041 26911 9059 26929
rect 8861 26875 8879 26893
rect 8897 26875 8915 26893
rect 8933 26875 8951 26893
rect 8969 26875 8987 26893
rect 9005 26875 9023 26893
rect 9041 26875 9059 26893
rect 8861 26839 8879 26857
rect 8897 26839 8915 26857
rect 8933 26839 8951 26857
rect 8969 26839 8987 26857
rect 9005 26839 9023 26857
rect 9041 26839 9059 26857
rect 8861 26803 8879 26821
rect 8897 26803 8915 26821
rect 8933 26803 8951 26821
rect 8969 26803 8987 26821
rect 9005 26803 9023 26821
rect 9041 26803 9059 26821
rect 8861 26767 8879 26785
rect 8897 26767 8915 26785
rect 8933 26767 8951 26785
rect 8969 26767 8987 26785
rect 9005 26767 9023 26785
rect 9041 26767 9059 26785
rect 8861 26731 8879 26749
rect 8897 26731 8915 26749
rect 8933 26731 8951 26749
rect 8969 26731 8987 26749
rect 9005 26731 9023 26749
rect 9041 26731 9059 26749
rect 8861 26695 8879 26713
rect 8897 26695 8915 26713
rect 8933 26695 8951 26713
rect 8969 26695 8987 26713
rect 9005 26695 9023 26713
rect 9041 26695 9059 26713
rect 8861 26659 8879 26677
rect 8897 26659 8915 26677
rect 8933 26659 8951 26677
rect 8969 26659 8987 26677
rect 9005 26659 9023 26677
rect 9041 26659 9059 26677
rect 8861 26623 8879 26641
rect 8897 26623 8915 26641
rect 8933 26623 8951 26641
rect 8969 26623 8987 26641
rect 9005 26623 9023 26641
rect 9041 26623 9059 26641
rect 8861 26587 8879 26605
rect 8897 26587 8915 26605
rect 8933 26587 8951 26605
rect 8969 26587 8987 26605
rect 9005 26587 9023 26605
rect 9041 26587 9059 26605
rect 8861 26551 8879 26569
rect 8897 26551 8915 26569
rect 8933 26551 8951 26569
rect 8969 26551 8987 26569
rect 9005 26551 9023 26569
rect 9041 26551 9059 26569
rect 8861 26515 8879 26533
rect 8897 26515 8915 26533
rect 8933 26515 8951 26533
rect 8969 26515 8987 26533
rect 9005 26515 9023 26533
rect 9041 26515 9059 26533
rect 8861 26479 8879 26497
rect 8897 26479 8915 26497
rect 8933 26479 8951 26497
rect 8969 26479 8987 26497
rect 9005 26479 9023 26497
rect 9041 26479 9059 26497
rect 8861 26443 8879 26461
rect 8897 26443 8915 26461
rect 8933 26443 8951 26461
rect 8969 26443 8987 26461
rect 9005 26443 9023 26461
rect 9041 26443 9059 26461
rect 28941 27757 28959 27775
rect 28977 27757 28995 27775
rect 29013 27757 29031 27775
rect 29049 27757 29067 27775
rect 29085 27757 29103 27775
rect 29121 27757 29139 27775
rect 28941 27721 28959 27739
rect 28977 27721 28995 27739
rect 29013 27721 29031 27739
rect 29049 27721 29067 27739
rect 29085 27721 29103 27739
rect 29121 27721 29139 27739
rect 28941 27685 28959 27703
rect 28977 27685 28995 27703
rect 29013 27685 29031 27703
rect 29049 27685 29067 27703
rect 29085 27685 29103 27703
rect 29121 27685 29139 27703
rect 28941 27649 28959 27667
rect 28977 27649 28995 27667
rect 29013 27649 29031 27667
rect 29049 27649 29067 27667
rect 29085 27649 29103 27667
rect 29121 27649 29139 27667
rect 28941 27613 28959 27631
rect 28977 27613 28995 27631
rect 29013 27613 29031 27631
rect 29049 27613 29067 27631
rect 29085 27613 29103 27631
rect 29121 27613 29139 27631
rect 28941 27577 28959 27595
rect 28977 27577 28995 27595
rect 29013 27577 29031 27595
rect 29049 27577 29067 27595
rect 29085 27577 29103 27595
rect 29121 27577 29139 27595
rect 28941 27541 28959 27559
rect 28977 27541 28995 27559
rect 29013 27541 29031 27559
rect 29049 27541 29067 27559
rect 29085 27541 29103 27559
rect 29121 27541 29139 27559
rect 28941 27505 28959 27523
rect 28977 27505 28995 27523
rect 29013 27505 29031 27523
rect 29049 27505 29067 27523
rect 29085 27505 29103 27523
rect 29121 27505 29139 27523
rect 28941 27469 28959 27487
rect 28977 27469 28995 27487
rect 29013 27469 29031 27487
rect 29049 27469 29067 27487
rect 29085 27469 29103 27487
rect 29121 27469 29139 27487
rect 28941 27433 28959 27451
rect 28977 27433 28995 27451
rect 29013 27433 29031 27451
rect 29049 27433 29067 27451
rect 29085 27433 29103 27451
rect 29121 27433 29139 27451
rect 28941 27397 28959 27415
rect 28977 27397 28995 27415
rect 29013 27397 29031 27415
rect 29049 27397 29067 27415
rect 29085 27397 29103 27415
rect 29121 27397 29139 27415
rect 28941 27361 28959 27379
rect 28977 27361 28995 27379
rect 29013 27361 29031 27379
rect 29049 27361 29067 27379
rect 29085 27361 29103 27379
rect 29121 27361 29139 27379
rect 28941 27325 28959 27343
rect 28977 27325 28995 27343
rect 29013 27325 29031 27343
rect 29049 27325 29067 27343
rect 29085 27325 29103 27343
rect 29121 27325 29139 27343
rect 28941 27289 28959 27307
rect 28977 27289 28995 27307
rect 29013 27289 29031 27307
rect 29049 27289 29067 27307
rect 29085 27289 29103 27307
rect 29121 27289 29139 27307
rect 28941 27253 28959 27271
rect 28977 27253 28995 27271
rect 29013 27253 29031 27271
rect 29049 27253 29067 27271
rect 29085 27253 29103 27271
rect 29121 27253 29139 27271
rect 28941 27217 28959 27235
rect 28977 27217 28995 27235
rect 29013 27217 29031 27235
rect 29049 27217 29067 27235
rect 29085 27217 29103 27235
rect 29121 27217 29139 27235
rect 28941 27181 28959 27199
rect 28977 27181 28995 27199
rect 29013 27181 29031 27199
rect 29049 27181 29067 27199
rect 29085 27181 29103 27199
rect 29121 27181 29139 27199
rect 28941 27145 28959 27163
rect 28977 27145 28995 27163
rect 29013 27145 29031 27163
rect 29049 27145 29067 27163
rect 29085 27145 29103 27163
rect 29121 27145 29139 27163
rect 28941 27109 28959 27127
rect 28977 27109 28995 27127
rect 29013 27109 29031 27127
rect 29049 27109 29067 27127
rect 29085 27109 29103 27127
rect 29121 27109 29139 27127
rect 28941 27073 28959 27091
rect 28977 27073 28995 27091
rect 29013 27073 29031 27091
rect 29049 27073 29067 27091
rect 29085 27073 29103 27091
rect 29121 27073 29139 27091
rect 28941 27037 28959 27055
rect 28977 27037 28995 27055
rect 29013 27037 29031 27055
rect 29049 27037 29067 27055
rect 29085 27037 29103 27055
rect 29121 27037 29139 27055
rect 28941 27001 28959 27019
rect 28977 27001 28995 27019
rect 29013 27001 29031 27019
rect 29049 27001 29067 27019
rect 29085 27001 29103 27019
rect 29121 27001 29139 27019
rect 28941 26965 28959 26983
rect 28977 26965 28995 26983
rect 29013 26965 29031 26983
rect 29049 26965 29067 26983
rect 29085 26965 29103 26983
rect 29121 26965 29139 26983
rect 28941 26929 28959 26947
rect 28977 26929 28995 26947
rect 29013 26929 29031 26947
rect 29049 26929 29067 26947
rect 29085 26929 29103 26947
rect 29121 26929 29139 26947
rect 28941 26893 28959 26911
rect 28977 26893 28995 26911
rect 29013 26893 29031 26911
rect 29049 26893 29067 26911
rect 29085 26893 29103 26911
rect 29121 26893 29139 26911
rect 28941 26857 28959 26875
rect 28977 26857 28995 26875
rect 29013 26857 29031 26875
rect 29049 26857 29067 26875
rect 29085 26857 29103 26875
rect 29121 26857 29139 26875
rect 28941 26821 28959 26839
rect 28977 26821 28995 26839
rect 29013 26821 29031 26839
rect 29049 26821 29067 26839
rect 29085 26821 29103 26839
rect 29121 26821 29139 26839
rect 28941 26785 28959 26803
rect 28977 26785 28995 26803
rect 29013 26785 29031 26803
rect 29049 26785 29067 26803
rect 29085 26785 29103 26803
rect 29121 26785 29139 26803
rect 28941 26749 28959 26767
rect 28977 26749 28995 26767
rect 29013 26749 29031 26767
rect 29049 26749 29067 26767
rect 29085 26749 29103 26767
rect 29121 26749 29139 26767
rect 28941 26713 28959 26731
rect 28977 26713 28995 26731
rect 29013 26713 29031 26731
rect 29049 26713 29067 26731
rect 29085 26713 29103 26731
rect 29121 26713 29139 26731
rect 28941 26677 28959 26695
rect 28977 26677 28995 26695
rect 29013 26677 29031 26695
rect 29049 26677 29067 26695
rect 29085 26677 29103 26695
rect 29121 26677 29139 26695
rect 28941 26641 28959 26659
rect 28977 26641 28995 26659
rect 29013 26641 29031 26659
rect 29049 26641 29067 26659
rect 29085 26641 29103 26659
rect 29121 26641 29139 26659
rect 28941 26605 28959 26623
rect 28977 26605 28995 26623
rect 29013 26605 29031 26623
rect 29049 26605 29067 26623
rect 29085 26605 29103 26623
rect 29121 26605 29139 26623
rect 28941 26569 28959 26587
rect 28977 26569 28995 26587
rect 29013 26569 29031 26587
rect 29049 26569 29067 26587
rect 29085 26569 29103 26587
rect 29121 26569 29139 26587
rect 28941 26533 28959 26551
rect 28977 26533 28995 26551
rect 29013 26533 29031 26551
rect 29049 26533 29067 26551
rect 29085 26533 29103 26551
rect 29121 26533 29139 26551
rect 28941 26497 28959 26515
rect 28977 26497 28995 26515
rect 29013 26497 29031 26515
rect 29049 26497 29067 26515
rect 29085 26497 29103 26515
rect 29121 26497 29139 26515
rect 28941 26461 28959 26479
rect 28977 26461 28995 26479
rect 29013 26461 29031 26479
rect 29049 26461 29067 26479
rect 29085 26461 29103 26479
rect 29121 26461 29139 26479
rect 28941 26425 28959 26443
rect 28977 26425 28995 26443
rect 29013 26425 29031 26443
rect 29049 26425 29067 26443
rect 29085 26425 29103 26443
rect 29121 26425 29139 26443
rect 28941 26389 28959 26407
rect 28977 26389 28995 26407
rect 29013 26389 29031 26407
rect 29049 26389 29067 26407
rect 29085 26389 29103 26407
rect 29121 26389 29139 26407
rect 28941 26353 28959 26371
rect 28977 26353 28995 26371
rect 29013 26353 29031 26371
rect 29049 26353 29067 26371
rect 29085 26353 29103 26371
rect 29121 26353 29139 26371
rect 28941 26317 28959 26335
rect 28977 26317 28995 26335
rect 29013 26317 29031 26335
rect 29049 26317 29067 26335
rect 29085 26317 29103 26335
rect 29121 26317 29139 26335
rect 28941 26281 28959 26299
rect 28977 26281 28995 26299
rect 29013 26281 29031 26299
rect 29049 26281 29067 26299
rect 29085 26281 29103 26299
rect 29121 26281 29139 26299
rect 28941 26245 28959 26263
rect 28977 26245 28995 26263
rect 29013 26245 29031 26263
rect 29049 26245 29067 26263
rect 29085 26245 29103 26263
rect 29121 26245 29139 26263
rect 28941 26209 28959 26227
rect 28977 26209 28995 26227
rect 29013 26209 29031 26227
rect 29049 26209 29067 26227
rect 29085 26209 29103 26227
rect 29121 26209 29139 26227
rect 28941 26173 28959 26191
rect 28977 26173 28995 26191
rect 29013 26173 29031 26191
rect 29049 26173 29067 26191
rect 29085 26173 29103 26191
rect 29121 26173 29139 26191
rect 8861 11529 8879 11547
rect 8897 11529 8915 11547
rect 8933 11529 8951 11547
rect 8969 11529 8987 11547
rect 9005 11529 9023 11547
rect 9041 11529 9059 11547
rect 8861 11493 8879 11511
rect 8897 11493 8915 11511
rect 8933 11493 8951 11511
rect 8969 11493 8987 11511
rect 9005 11493 9023 11511
rect 9041 11493 9059 11511
rect 8861 11457 8879 11475
rect 8897 11457 8915 11475
rect 8933 11457 8951 11475
rect 8969 11457 8987 11475
rect 9005 11457 9023 11475
rect 9041 11457 9059 11475
rect 8861 11421 8879 11439
rect 8897 11421 8915 11439
rect 8933 11421 8951 11439
rect 8969 11421 8987 11439
rect 9005 11421 9023 11439
rect 9041 11421 9059 11439
rect 8861 11385 8879 11403
rect 8897 11385 8915 11403
rect 8933 11385 8951 11403
rect 8969 11385 8987 11403
rect 9005 11385 9023 11403
rect 9041 11385 9059 11403
rect 8861 11349 8879 11367
rect 8897 11349 8915 11367
rect 8933 11349 8951 11367
rect 8969 11349 8987 11367
rect 9005 11349 9023 11367
rect 9041 11349 9059 11367
rect 8861 11313 8879 11331
rect 8897 11313 8915 11331
rect 8933 11313 8951 11331
rect 8969 11313 8987 11331
rect 9005 11313 9023 11331
rect 9041 11313 9059 11331
rect 8861 11277 8879 11295
rect 8897 11277 8915 11295
rect 8933 11277 8951 11295
rect 8969 11277 8987 11295
rect 9005 11277 9023 11295
rect 9041 11277 9059 11295
rect 8861 11241 8879 11259
rect 8897 11241 8915 11259
rect 8933 11241 8951 11259
rect 8969 11241 8987 11259
rect 9005 11241 9023 11259
rect 9041 11241 9059 11259
rect 8861 11205 8879 11223
rect 8897 11205 8915 11223
rect 8933 11205 8951 11223
rect 8969 11205 8987 11223
rect 9005 11205 9023 11223
rect 9041 11205 9059 11223
rect 8861 11169 8879 11187
rect 8897 11169 8915 11187
rect 8933 11169 8951 11187
rect 8969 11169 8987 11187
rect 9005 11169 9023 11187
rect 9041 11169 9059 11187
rect 8861 11133 8879 11151
rect 8897 11133 8915 11151
rect 8933 11133 8951 11151
rect 8969 11133 8987 11151
rect 9005 11133 9023 11151
rect 9041 11133 9059 11151
rect 8861 11097 8879 11115
rect 8897 11097 8915 11115
rect 8933 11097 8951 11115
rect 8969 11097 8987 11115
rect 9005 11097 9023 11115
rect 9041 11097 9059 11115
rect 8861 11061 8879 11079
rect 8897 11061 8915 11079
rect 8933 11061 8951 11079
rect 8969 11061 8987 11079
rect 9005 11061 9023 11079
rect 9041 11061 9059 11079
rect 8861 11025 8879 11043
rect 8897 11025 8915 11043
rect 8933 11025 8951 11043
rect 8969 11025 8987 11043
rect 9005 11025 9023 11043
rect 9041 11025 9059 11043
rect 8861 10989 8879 11007
rect 8897 10989 8915 11007
rect 8933 10989 8951 11007
rect 8969 10989 8987 11007
rect 9005 10989 9023 11007
rect 9041 10989 9059 11007
rect 8861 10953 8879 10971
rect 8897 10953 8915 10971
rect 8933 10953 8951 10971
rect 8969 10953 8987 10971
rect 9005 10953 9023 10971
rect 9041 10953 9059 10971
rect 8861 10917 8879 10935
rect 8897 10917 8915 10935
rect 8933 10917 8951 10935
rect 8969 10917 8987 10935
rect 9005 10917 9023 10935
rect 9041 10917 9059 10935
rect 8861 10881 8879 10899
rect 8897 10881 8915 10899
rect 8933 10881 8951 10899
rect 8969 10881 8987 10899
rect 9005 10881 9023 10899
rect 9041 10881 9059 10899
rect 8861 10845 8879 10863
rect 8897 10845 8915 10863
rect 8933 10845 8951 10863
rect 8969 10845 8987 10863
rect 9005 10845 9023 10863
rect 9041 10845 9059 10863
rect 8861 10809 8879 10827
rect 8897 10809 8915 10827
rect 8933 10809 8951 10827
rect 8969 10809 8987 10827
rect 9005 10809 9023 10827
rect 9041 10809 9059 10827
rect 8861 10773 8879 10791
rect 8897 10773 8915 10791
rect 8933 10773 8951 10791
rect 8969 10773 8987 10791
rect 9005 10773 9023 10791
rect 9041 10773 9059 10791
rect 8861 10737 8879 10755
rect 8897 10737 8915 10755
rect 8933 10737 8951 10755
rect 8969 10737 8987 10755
rect 9005 10737 9023 10755
rect 9041 10737 9059 10755
rect 8861 10701 8879 10719
rect 8897 10701 8915 10719
rect 8933 10701 8951 10719
rect 8969 10701 8987 10719
rect 9005 10701 9023 10719
rect 9041 10701 9059 10719
rect 8861 10665 8879 10683
rect 8897 10665 8915 10683
rect 8933 10665 8951 10683
rect 8969 10665 8987 10683
rect 9005 10665 9023 10683
rect 9041 10665 9059 10683
rect 8861 10629 8879 10647
rect 8897 10629 8915 10647
rect 8933 10629 8951 10647
rect 8969 10629 8987 10647
rect 9005 10629 9023 10647
rect 9041 10629 9059 10647
rect 8861 10593 8879 10611
rect 8897 10593 8915 10611
rect 8933 10593 8951 10611
rect 8969 10593 8987 10611
rect 9005 10593 9023 10611
rect 9041 10593 9059 10611
rect 8861 10557 8879 10575
rect 8897 10557 8915 10575
rect 8933 10557 8951 10575
rect 8969 10557 8987 10575
rect 9005 10557 9023 10575
rect 9041 10557 9059 10575
rect 8861 10521 8879 10539
rect 8897 10521 8915 10539
rect 8933 10521 8951 10539
rect 8969 10521 8987 10539
rect 9005 10521 9023 10539
rect 9041 10521 9059 10539
rect 8861 10485 8879 10503
rect 8897 10485 8915 10503
rect 8933 10485 8951 10503
rect 8969 10485 8987 10503
rect 9005 10485 9023 10503
rect 9041 10485 9059 10503
rect 8861 10449 8879 10467
rect 8897 10449 8915 10467
rect 8933 10449 8951 10467
rect 8969 10449 8987 10467
rect 9005 10449 9023 10467
rect 9041 10449 9059 10467
rect 8861 10413 8879 10431
rect 8897 10413 8915 10431
rect 8933 10413 8951 10431
rect 8969 10413 8987 10431
rect 9005 10413 9023 10431
rect 9041 10413 9059 10431
rect 8861 10377 8879 10395
rect 8897 10377 8915 10395
rect 8933 10377 8951 10395
rect 8969 10377 8987 10395
rect 9005 10377 9023 10395
rect 9041 10377 9059 10395
rect 8861 10341 8879 10359
rect 8897 10341 8915 10359
rect 8933 10341 8951 10359
rect 8969 10341 8987 10359
rect 9005 10341 9023 10359
rect 9041 10341 9059 10359
rect 8861 10305 8879 10323
rect 8897 10305 8915 10323
rect 8933 10305 8951 10323
rect 8969 10305 8987 10323
rect 9005 10305 9023 10323
rect 9041 10305 9059 10323
rect 8861 10269 8879 10287
rect 8897 10269 8915 10287
rect 8933 10269 8951 10287
rect 8969 10269 8987 10287
rect 9005 10269 9023 10287
rect 9041 10269 9059 10287
rect 8861 10233 8879 10251
rect 8897 10233 8915 10251
rect 8933 10233 8951 10251
rect 8969 10233 8987 10251
rect 9005 10233 9023 10251
rect 9041 10233 9059 10251
<< metal2 >>
rect 11960 29003 12040 29180
rect 11960 28985 11973 29003
rect 11991 28985 12009 29003
rect 12027 28985 12040 29003
rect 11960 28967 12040 28985
rect 11960 28949 11973 28967
rect 11991 28949 12009 28967
rect 12027 28949 12040 28967
rect 11960 28931 12040 28949
rect 11960 28913 11973 28931
rect 11991 28913 12009 28931
rect 12027 28913 12040 28931
rect 11960 28895 12040 28913
rect 11960 28877 11973 28895
rect 11991 28877 12009 28895
rect 12027 28877 12040 28895
rect 11960 28860 12040 28877
rect 12400 28923 12480 28940
rect 12400 28905 12413 28923
rect 12431 28905 12449 28923
rect 12467 28905 12480 28923
rect 12400 28887 12480 28905
rect 12400 28869 12413 28887
rect 12431 28869 12449 28887
rect 12467 28869 12480 28887
rect 12400 28851 12480 28869
rect 12400 28833 12413 28851
rect 12431 28833 12449 28851
rect 12467 28833 12480 28851
rect 12400 28815 12480 28833
rect 12400 28797 12413 28815
rect 12431 28797 12449 28815
rect 12467 28797 12480 28815
rect 12400 28220 12480 28797
rect 14660 28380 14740 29180
rect 17360 28500 17440 29180
rect 20060 28620 20140 29180
rect 22760 28740 22840 29180
rect 25460 28740 25540 29180
rect 22760 28719 22940 28740
rect 22760 28701 22787 28719
rect 22805 28701 22823 28719
rect 22841 28701 22859 28719
rect 22877 28701 22895 28719
rect 22913 28701 22940 28719
rect 22760 28680 22940 28701
rect 24040 28719 24220 28740
rect 24040 28701 24067 28719
rect 24085 28701 24103 28719
rect 24121 28701 24139 28719
rect 24157 28701 24175 28719
rect 24193 28701 24220 28719
rect 24040 28680 24220 28701
rect 20060 28599 22000 28620
rect 20060 28581 21847 28599
rect 21865 28581 21883 28599
rect 21901 28581 21919 28599
rect 21937 28581 21955 28599
rect 21973 28581 22000 28599
rect 20060 28560 22000 28581
rect 23900 28599 24080 28620
rect 23900 28581 23927 28599
rect 23945 28581 23963 28599
rect 23981 28581 23999 28599
rect 24017 28581 24035 28599
rect 24053 28581 24080 28599
rect 23900 28560 24080 28581
rect 17360 28479 17540 28500
rect 17360 28461 17387 28479
rect 17405 28461 17423 28479
rect 17441 28461 17459 28479
rect 17477 28461 17495 28479
rect 17513 28461 17540 28479
rect 17360 28440 17540 28461
rect 19420 28479 20620 28500
rect 19420 28461 19447 28479
rect 19465 28461 19483 28479
rect 19501 28461 19519 28479
rect 19537 28461 19555 28479
rect 19573 28461 20620 28479
rect 19420 28440 20620 28461
rect 14660 28359 14840 28380
rect 14660 28341 14687 28359
rect 14705 28341 14723 28359
rect 14741 28341 14759 28359
rect 14777 28341 14795 28359
rect 14813 28341 14840 28359
rect 14660 28320 14840 28341
rect 17180 28359 18820 28380
rect 17180 28341 17207 28359
rect 17225 28341 17243 28359
rect 17261 28341 17279 28359
rect 17297 28341 17315 28359
rect 17333 28341 18820 28359
rect 17180 28320 18820 28341
rect 18760 28220 18820 28320
rect 20560 28220 20620 28440
rect 24020 28220 24080 28560
rect 24160 28220 24220 28680
rect 24460 28719 24640 28740
rect 24460 28701 24487 28719
rect 24505 28701 24523 28719
rect 24541 28701 24559 28719
rect 24577 28701 24595 28719
rect 24613 28701 24640 28719
rect 24460 28680 24640 28701
rect 25360 28719 25540 28740
rect 25360 28701 25387 28719
rect 25405 28701 25423 28719
rect 25441 28701 25459 28719
rect 25477 28701 25495 28719
rect 25513 28701 25540 28719
rect 25360 28680 25540 28701
rect 24460 28220 24520 28680
rect 28160 28620 28240 29180
rect 24580 28599 25740 28620
rect 24580 28581 25587 28599
rect 25605 28581 25623 28599
rect 25641 28581 25659 28599
rect 25677 28581 25695 28599
rect 25713 28581 25740 28599
rect 24580 28560 25740 28581
rect 28060 28599 28240 28620
rect 28060 28581 28087 28599
rect 28105 28581 28123 28599
rect 28141 28581 28159 28599
rect 28177 28581 28195 28599
rect 28213 28581 28240 28599
rect 28060 28560 28240 28581
rect 24580 28220 24660 28560
rect 28920 28027 29180 28040
rect 28920 28009 28941 28027
rect 28959 28009 28977 28027
rect 28995 28009 29013 28027
rect 29031 28009 29049 28027
rect 29067 28009 29085 28027
rect 29103 28009 29121 28027
rect 29139 28009 29180 28027
rect 28920 27991 29180 28009
rect 28920 27973 28941 27991
rect 28959 27973 28977 27991
rect 28995 27973 29013 27991
rect 29031 27973 29049 27991
rect 29067 27973 29085 27991
rect 29103 27973 29121 27991
rect 29139 27973 29180 27991
rect 28920 27955 29180 27973
rect 28920 27937 28941 27955
rect 28959 27937 28977 27955
rect 28995 27937 29013 27955
rect 29031 27937 29049 27955
rect 29067 27937 29085 27955
rect 29103 27937 29121 27955
rect 29139 27937 29180 27955
rect 28920 27919 29180 27937
rect 28920 27901 28941 27919
rect 28959 27901 28977 27919
rect 28995 27901 29013 27919
rect 29031 27901 29049 27919
rect 29067 27901 29085 27919
rect 29103 27901 29121 27919
rect 29139 27901 29180 27919
rect 28920 27883 29180 27901
rect 28920 27865 28941 27883
rect 28959 27865 28977 27883
rect 28995 27865 29013 27883
rect 29031 27865 29049 27883
rect 29067 27865 29085 27883
rect 29103 27865 29121 27883
rect 29139 27865 29180 27883
rect 28920 27847 29180 27865
rect 28920 27829 28941 27847
rect 28959 27829 28977 27847
rect 28995 27829 29013 27847
rect 29031 27829 29049 27847
rect 29067 27829 29085 27847
rect 29103 27829 29121 27847
rect 29139 27829 29180 27847
rect 28920 27811 29180 27829
rect 28920 27793 28941 27811
rect 28959 27793 28977 27811
rect 28995 27793 29013 27811
rect 29031 27793 29049 27811
rect 29067 27793 29085 27811
rect 29103 27793 29121 27811
rect 29139 27793 29180 27811
rect 8820 27757 9080 27780
rect 8820 27739 8861 27757
rect 8879 27739 8897 27757
rect 8915 27739 8933 27757
rect 8951 27739 8969 27757
rect 8987 27739 9005 27757
rect 9023 27739 9041 27757
rect 9059 27739 9080 27757
rect 8820 27721 9080 27739
rect 8820 27703 8861 27721
rect 8879 27703 8897 27721
rect 8915 27703 8933 27721
rect 8951 27703 8969 27721
rect 8987 27703 9005 27721
rect 9023 27703 9041 27721
rect 9059 27703 9080 27721
rect 8820 27685 9080 27703
rect 8820 27667 8861 27685
rect 8879 27667 8897 27685
rect 8915 27667 8933 27685
rect 8951 27667 8969 27685
rect 8987 27667 9005 27685
rect 9023 27667 9041 27685
rect 9059 27667 9080 27685
rect 8820 27649 9080 27667
rect 8820 27631 8861 27649
rect 8879 27631 8897 27649
rect 8915 27631 8933 27649
rect 8951 27631 8969 27649
rect 8987 27631 9005 27649
rect 9023 27631 9041 27649
rect 9059 27631 9080 27649
rect 8820 27613 9080 27631
rect 8820 27595 8861 27613
rect 8879 27595 8897 27613
rect 8915 27595 8933 27613
rect 8951 27595 8969 27613
rect 8987 27595 9005 27613
rect 9023 27595 9041 27613
rect 9059 27595 9080 27613
rect 8820 27577 9080 27595
rect 8820 27559 8861 27577
rect 8879 27559 8897 27577
rect 8915 27559 8933 27577
rect 8951 27559 8969 27577
rect 8987 27559 9005 27577
rect 9023 27559 9041 27577
rect 9059 27559 9080 27577
rect 8820 27541 9080 27559
rect 8820 27523 8861 27541
rect 8879 27523 8897 27541
rect 8915 27523 8933 27541
rect 8951 27523 8969 27541
rect 8987 27523 9005 27541
rect 9023 27523 9041 27541
rect 9059 27523 9080 27541
rect 8820 27505 9080 27523
rect 8820 27487 8861 27505
rect 8879 27487 8897 27505
rect 8915 27487 8933 27505
rect 8951 27487 8969 27505
rect 8987 27487 9005 27505
rect 9023 27487 9041 27505
rect 9059 27487 9080 27505
rect 8820 27469 9080 27487
rect 8820 27451 8861 27469
rect 8879 27451 8897 27469
rect 8915 27451 8933 27469
rect 8951 27451 8969 27469
rect 8987 27451 9005 27469
rect 9023 27451 9041 27469
rect 9059 27451 9080 27469
rect 8820 27433 9080 27451
rect 8820 27415 8861 27433
rect 8879 27415 8897 27433
rect 8915 27415 8933 27433
rect 8951 27415 8969 27433
rect 8987 27415 9005 27433
rect 9023 27415 9041 27433
rect 9059 27415 9080 27433
rect 8820 27397 9080 27415
rect 8820 27379 8861 27397
rect 8879 27379 8897 27397
rect 8915 27379 8933 27397
rect 8951 27379 8969 27397
rect 8987 27379 9005 27397
rect 9023 27379 9041 27397
rect 9059 27379 9080 27397
rect 8820 27361 9080 27379
rect 8820 27343 8861 27361
rect 8879 27343 8897 27361
rect 8915 27343 8933 27361
rect 8951 27343 8969 27361
rect 8987 27343 9005 27361
rect 9023 27343 9041 27361
rect 9059 27343 9080 27361
rect 8820 27325 9080 27343
rect 8820 27307 8861 27325
rect 8879 27307 8897 27325
rect 8915 27307 8933 27325
rect 8951 27307 8969 27325
rect 8987 27307 9005 27325
rect 9023 27307 9041 27325
rect 9059 27307 9080 27325
rect 8820 27289 9080 27307
rect 8820 27271 8861 27289
rect 8879 27271 8897 27289
rect 8915 27271 8933 27289
rect 8951 27271 8969 27289
rect 8987 27271 9005 27289
rect 9023 27271 9041 27289
rect 9059 27271 9080 27289
rect 8820 27253 9080 27271
rect 8820 27235 8861 27253
rect 8879 27235 8897 27253
rect 8915 27235 8933 27253
rect 8951 27235 8969 27253
rect 8987 27235 9005 27253
rect 9023 27235 9041 27253
rect 9059 27235 9080 27253
rect 8820 27217 9080 27235
rect 8820 27199 8861 27217
rect 8879 27199 8897 27217
rect 8915 27199 8933 27217
rect 8951 27199 8969 27217
rect 8987 27199 9005 27217
rect 9023 27199 9041 27217
rect 9059 27199 9080 27217
rect 8820 27181 9080 27199
rect 8820 27163 8861 27181
rect 8879 27163 8897 27181
rect 8915 27163 8933 27181
rect 8951 27163 8969 27181
rect 8987 27163 9005 27181
rect 9023 27163 9041 27181
rect 9059 27163 9080 27181
rect 8820 27145 9080 27163
rect 8820 27127 8861 27145
rect 8879 27127 8897 27145
rect 8915 27127 8933 27145
rect 8951 27127 8969 27145
rect 8987 27127 9005 27145
rect 9023 27127 9041 27145
rect 9059 27127 9080 27145
rect 8820 27109 9080 27127
rect 8820 27091 8861 27109
rect 8879 27091 8897 27109
rect 8915 27091 8933 27109
rect 8951 27091 8969 27109
rect 8987 27091 9005 27109
rect 9023 27091 9041 27109
rect 9059 27091 9080 27109
rect 8820 27073 9080 27091
rect 8820 27055 8861 27073
rect 8879 27055 8897 27073
rect 8915 27055 8933 27073
rect 8951 27055 8969 27073
rect 8987 27055 9005 27073
rect 9023 27055 9041 27073
rect 9059 27055 9080 27073
rect 8820 27037 9080 27055
rect 8820 27019 8861 27037
rect 8879 27019 8897 27037
rect 8915 27019 8933 27037
rect 8951 27019 8969 27037
rect 8987 27019 9005 27037
rect 9023 27019 9041 27037
rect 9059 27019 9080 27037
rect 8820 27001 9080 27019
rect 8820 26983 8861 27001
rect 8879 26983 8897 27001
rect 8915 26983 8933 27001
rect 8951 26983 8969 27001
rect 8987 26983 9005 27001
rect 9023 26983 9041 27001
rect 9059 26983 9080 27001
rect 8820 26965 9080 26983
rect 8820 26947 8861 26965
rect 8879 26947 8897 26965
rect 8915 26947 8933 26965
rect 8951 26947 8969 26965
rect 8987 26947 9005 26965
rect 9023 26947 9041 26965
rect 9059 26947 9080 26965
rect 8820 26929 9080 26947
rect 8820 26911 8861 26929
rect 8879 26911 8897 26929
rect 8915 26911 8933 26929
rect 8951 26911 8969 26929
rect 8987 26911 9005 26929
rect 9023 26911 9041 26929
rect 9059 26911 9080 26929
rect 8820 26893 9080 26911
rect 8820 26875 8861 26893
rect 8879 26875 8897 26893
rect 8915 26875 8933 26893
rect 8951 26875 8969 26893
rect 8987 26875 9005 26893
rect 9023 26875 9041 26893
rect 9059 26875 9080 26893
rect 8820 26857 9080 26875
rect 8820 26839 8861 26857
rect 8879 26839 8897 26857
rect 8915 26839 8933 26857
rect 8951 26839 8969 26857
rect 8987 26839 9005 26857
rect 9023 26839 9041 26857
rect 9059 26839 9080 26857
rect 8820 26821 9080 26839
rect 8820 26803 8861 26821
rect 8879 26803 8897 26821
rect 8915 26803 8933 26821
rect 8951 26803 8969 26821
rect 8987 26803 9005 26821
rect 9023 26803 9041 26821
rect 9059 26803 9080 26821
rect 8820 26785 9080 26803
rect 8820 26767 8861 26785
rect 8879 26767 8897 26785
rect 8915 26767 8933 26785
rect 8951 26767 8969 26785
rect 8987 26767 9005 26785
rect 9023 26767 9041 26785
rect 9059 26767 9080 26785
rect 8820 26749 9080 26767
rect 8820 26731 8861 26749
rect 8879 26731 8897 26749
rect 8915 26731 8933 26749
rect 8951 26731 8969 26749
rect 8987 26731 9005 26749
rect 9023 26731 9041 26749
rect 9059 26731 9080 26749
rect 8820 26713 9080 26731
rect 8820 26695 8861 26713
rect 8879 26695 8897 26713
rect 8915 26695 8933 26713
rect 8951 26695 8969 26713
rect 8987 26695 9005 26713
rect 9023 26695 9041 26713
rect 9059 26695 9080 26713
rect 8820 26677 9080 26695
rect 8820 26659 8861 26677
rect 8879 26659 8897 26677
rect 8915 26659 8933 26677
rect 8951 26659 8969 26677
rect 8987 26659 9005 26677
rect 9023 26659 9041 26677
rect 9059 26659 9080 26677
rect 8820 26641 9080 26659
rect 8820 26623 8861 26641
rect 8879 26623 8897 26641
rect 8915 26623 8933 26641
rect 8951 26623 8969 26641
rect 8987 26623 9005 26641
rect 9023 26623 9041 26641
rect 9059 26623 9080 26641
rect 8820 26605 9080 26623
rect 8820 26587 8861 26605
rect 8879 26587 8897 26605
rect 8915 26587 8933 26605
rect 8951 26587 8969 26605
rect 8987 26587 9005 26605
rect 9023 26587 9041 26605
rect 9059 26587 9080 26605
rect 8820 26569 9080 26587
rect 8820 26551 8861 26569
rect 8879 26551 8897 26569
rect 8915 26551 8933 26569
rect 8951 26551 8969 26569
rect 8987 26551 9005 26569
rect 9023 26551 9041 26569
rect 9059 26551 9080 26569
rect 8820 26533 9080 26551
rect 8820 26515 8861 26533
rect 8879 26515 8897 26533
rect 8915 26515 8933 26533
rect 8951 26515 8969 26533
rect 8987 26515 9005 26533
rect 9023 26515 9041 26533
rect 9059 26515 9080 26533
rect 8820 26497 9080 26515
rect 8820 26479 8861 26497
rect 8879 26479 8897 26497
rect 8915 26479 8933 26497
rect 8951 26479 8969 26497
rect 8987 26479 9005 26497
rect 9023 26479 9041 26497
rect 9059 26479 9080 26497
rect 8820 26461 9080 26479
rect 8820 26443 8861 26461
rect 8879 26443 8897 26461
rect 8915 26443 8933 26461
rect 8951 26443 8969 26461
rect 8987 26443 9005 26461
rect 9023 26443 9041 26461
rect 9059 26443 9080 26461
rect 8820 26420 9080 26443
rect 28920 27775 29180 27793
rect 28920 27757 28941 27775
rect 28959 27757 28977 27775
rect 28995 27757 29013 27775
rect 29031 27757 29049 27775
rect 29067 27757 29085 27775
rect 29103 27757 29121 27775
rect 29139 27757 29180 27775
rect 28920 27739 29180 27757
rect 28920 27721 28941 27739
rect 28959 27721 28977 27739
rect 28995 27721 29013 27739
rect 29031 27721 29049 27739
rect 29067 27721 29085 27739
rect 29103 27721 29121 27739
rect 29139 27721 29180 27739
rect 28920 27703 29180 27721
rect 28920 27685 28941 27703
rect 28959 27685 28977 27703
rect 28995 27685 29013 27703
rect 29031 27685 29049 27703
rect 29067 27685 29085 27703
rect 29103 27685 29121 27703
rect 29139 27685 29180 27703
rect 28920 27667 29180 27685
rect 28920 27649 28941 27667
rect 28959 27649 28977 27667
rect 28995 27649 29013 27667
rect 29031 27649 29049 27667
rect 29067 27649 29085 27667
rect 29103 27649 29121 27667
rect 29139 27649 29180 27667
rect 28920 27631 29180 27649
rect 28920 27613 28941 27631
rect 28959 27613 28977 27631
rect 28995 27613 29013 27631
rect 29031 27613 29049 27631
rect 29067 27613 29085 27631
rect 29103 27613 29121 27631
rect 29139 27613 29180 27631
rect 28920 27595 29180 27613
rect 28920 27577 28941 27595
rect 28959 27577 28977 27595
rect 28995 27577 29013 27595
rect 29031 27577 29049 27595
rect 29067 27577 29085 27595
rect 29103 27577 29121 27595
rect 29139 27577 29180 27595
rect 28920 27559 29180 27577
rect 28920 27541 28941 27559
rect 28959 27541 28977 27559
rect 28995 27541 29013 27559
rect 29031 27541 29049 27559
rect 29067 27541 29085 27559
rect 29103 27541 29121 27559
rect 29139 27541 29180 27559
rect 28920 27523 29180 27541
rect 28920 27505 28941 27523
rect 28959 27505 28977 27523
rect 28995 27505 29013 27523
rect 29031 27505 29049 27523
rect 29067 27505 29085 27523
rect 29103 27505 29121 27523
rect 29139 27505 29180 27523
rect 28920 27487 29180 27505
rect 28920 27469 28941 27487
rect 28959 27469 28977 27487
rect 28995 27469 29013 27487
rect 29031 27469 29049 27487
rect 29067 27469 29085 27487
rect 29103 27469 29121 27487
rect 29139 27469 29180 27487
rect 28920 27451 29180 27469
rect 28920 27433 28941 27451
rect 28959 27433 28977 27451
rect 28995 27433 29013 27451
rect 29031 27433 29049 27451
rect 29067 27433 29085 27451
rect 29103 27433 29121 27451
rect 29139 27433 29180 27451
rect 28920 27415 29180 27433
rect 28920 27397 28941 27415
rect 28959 27397 28977 27415
rect 28995 27397 29013 27415
rect 29031 27397 29049 27415
rect 29067 27397 29085 27415
rect 29103 27397 29121 27415
rect 29139 27397 29180 27415
rect 28920 27379 29180 27397
rect 28920 27361 28941 27379
rect 28959 27361 28977 27379
rect 28995 27361 29013 27379
rect 29031 27361 29049 27379
rect 29067 27361 29085 27379
rect 29103 27361 29121 27379
rect 29139 27361 29180 27379
rect 28920 27343 29180 27361
rect 28920 27325 28941 27343
rect 28959 27325 28977 27343
rect 28995 27325 29013 27343
rect 29031 27325 29049 27343
rect 29067 27325 29085 27343
rect 29103 27325 29121 27343
rect 29139 27325 29180 27343
rect 28920 27307 29180 27325
rect 28920 27289 28941 27307
rect 28959 27289 28977 27307
rect 28995 27289 29013 27307
rect 29031 27289 29049 27307
rect 29067 27289 29085 27307
rect 29103 27289 29121 27307
rect 29139 27289 29180 27307
rect 28920 27271 29180 27289
rect 28920 27253 28941 27271
rect 28959 27253 28977 27271
rect 28995 27253 29013 27271
rect 29031 27253 29049 27271
rect 29067 27253 29085 27271
rect 29103 27253 29121 27271
rect 29139 27253 29180 27271
rect 28920 27235 29180 27253
rect 28920 27217 28941 27235
rect 28959 27217 28977 27235
rect 28995 27217 29013 27235
rect 29031 27217 29049 27235
rect 29067 27217 29085 27235
rect 29103 27217 29121 27235
rect 29139 27217 29180 27235
rect 28920 27199 29180 27217
rect 28920 27181 28941 27199
rect 28959 27181 28977 27199
rect 28995 27181 29013 27199
rect 29031 27181 29049 27199
rect 29067 27181 29085 27199
rect 29103 27181 29121 27199
rect 29139 27181 29180 27199
rect 28920 27163 29180 27181
rect 28920 27145 28941 27163
rect 28959 27145 28977 27163
rect 28995 27145 29013 27163
rect 29031 27145 29049 27163
rect 29067 27145 29085 27163
rect 29103 27145 29121 27163
rect 29139 27145 29180 27163
rect 28920 27127 29180 27145
rect 28920 27109 28941 27127
rect 28959 27109 28977 27127
rect 28995 27109 29013 27127
rect 29031 27109 29049 27127
rect 29067 27109 29085 27127
rect 29103 27109 29121 27127
rect 29139 27109 29180 27127
rect 28920 27091 29180 27109
rect 28920 27073 28941 27091
rect 28959 27073 28977 27091
rect 28995 27073 29013 27091
rect 29031 27073 29049 27091
rect 29067 27073 29085 27091
rect 29103 27073 29121 27091
rect 29139 27073 29180 27091
rect 28920 27055 29180 27073
rect 28920 27037 28941 27055
rect 28959 27037 28977 27055
rect 28995 27037 29013 27055
rect 29031 27037 29049 27055
rect 29067 27037 29085 27055
rect 29103 27037 29121 27055
rect 29139 27037 29180 27055
rect 28920 27019 29180 27037
rect 28920 27001 28941 27019
rect 28959 27001 28977 27019
rect 28995 27001 29013 27019
rect 29031 27001 29049 27019
rect 29067 27001 29085 27019
rect 29103 27001 29121 27019
rect 29139 27001 29180 27019
rect 28920 26983 29180 27001
rect 28920 26965 28941 26983
rect 28959 26965 28977 26983
rect 28995 26965 29013 26983
rect 29031 26965 29049 26983
rect 29067 26965 29085 26983
rect 29103 26965 29121 26983
rect 29139 26965 29180 26983
rect 28920 26947 29180 26965
rect 28920 26929 28941 26947
rect 28959 26929 28977 26947
rect 28995 26929 29013 26947
rect 29031 26929 29049 26947
rect 29067 26929 29085 26947
rect 29103 26929 29121 26947
rect 29139 26929 29180 26947
rect 28920 26911 29180 26929
rect 28920 26893 28941 26911
rect 28959 26893 28977 26911
rect 28995 26893 29013 26911
rect 29031 26893 29049 26911
rect 29067 26893 29085 26911
rect 29103 26893 29121 26911
rect 29139 26893 29180 26911
rect 28920 26875 29180 26893
rect 28920 26857 28941 26875
rect 28959 26857 28977 26875
rect 28995 26857 29013 26875
rect 29031 26857 29049 26875
rect 29067 26857 29085 26875
rect 29103 26857 29121 26875
rect 29139 26857 29180 26875
rect 28920 26839 29180 26857
rect 28920 26821 28941 26839
rect 28959 26821 28977 26839
rect 28995 26821 29013 26839
rect 29031 26821 29049 26839
rect 29067 26821 29085 26839
rect 29103 26821 29121 26839
rect 29139 26821 29180 26839
rect 28920 26803 29180 26821
rect 28920 26785 28941 26803
rect 28959 26785 28977 26803
rect 28995 26785 29013 26803
rect 29031 26785 29049 26803
rect 29067 26785 29085 26803
rect 29103 26785 29121 26803
rect 29139 26785 29180 26803
rect 28920 26767 29180 26785
rect 28920 26749 28941 26767
rect 28959 26749 28977 26767
rect 28995 26749 29013 26767
rect 29031 26749 29049 26767
rect 29067 26749 29085 26767
rect 29103 26749 29121 26767
rect 29139 26749 29180 26767
rect 28920 26731 29180 26749
rect 28920 26713 28941 26731
rect 28959 26713 28977 26731
rect 28995 26713 29013 26731
rect 29031 26713 29049 26731
rect 29067 26713 29085 26731
rect 29103 26713 29121 26731
rect 29139 26713 29180 26731
rect 28920 26695 29180 26713
rect 28920 26677 28941 26695
rect 28959 26677 28977 26695
rect 28995 26677 29013 26695
rect 29031 26677 29049 26695
rect 29067 26677 29085 26695
rect 29103 26677 29121 26695
rect 29139 26677 29180 26695
rect 28920 26659 29180 26677
rect 28920 26641 28941 26659
rect 28959 26641 28977 26659
rect 28995 26641 29013 26659
rect 29031 26641 29049 26659
rect 29067 26641 29085 26659
rect 29103 26641 29121 26659
rect 29139 26641 29180 26659
rect 28920 26623 29180 26641
rect 28920 26605 28941 26623
rect 28959 26605 28977 26623
rect 28995 26605 29013 26623
rect 29031 26605 29049 26623
rect 29067 26605 29085 26623
rect 29103 26605 29121 26623
rect 29139 26605 29180 26623
rect 28920 26587 29180 26605
rect 28920 26569 28941 26587
rect 28959 26569 28977 26587
rect 28995 26569 29013 26587
rect 29031 26569 29049 26587
rect 29067 26569 29085 26587
rect 29103 26569 29121 26587
rect 29139 26569 29180 26587
rect 28920 26551 29180 26569
rect 28920 26533 28941 26551
rect 28959 26533 28977 26551
rect 28995 26533 29013 26551
rect 29031 26533 29049 26551
rect 29067 26533 29085 26551
rect 29103 26533 29121 26551
rect 29139 26533 29180 26551
rect 28920 26515 29180 26533
rect 28920 26497 28941 26515
rect 28959 26497 28977 26515
rect 28995 26497 29013 26515
rect 29031 26497 29049 26515
rect 29067 26497 29085 26515
rect 29103 26497 29121 26515
rect 29139 26497 29180 26515
rect 28920 26479 29180 26497
rect 28920 26461 28941 26479
rect 28959 26461 28977 26479
rect 28995 26461 29013 26479
rect 29031 26461 29049 26479
rect 29067 26461 29085 26479
rect 29103 26461 29121 26479
rect 29139 26461 29180 26479
rect 28920 26443 29180 26461
rect 28920 26425 28941 26443
rect 28959 26425 28977 26443
rect 28995 26425 29013 26443
rect 29031 26425 29049 26443
rect 29067 26425 29085 26443
rect 29103 26425 29121 26443
rect 29139 26425 29180 26443
rect 28920 26407 29180 26425
rect 28920 26389 28941 26407
rect 28959 26389 28977 26407
rect 28995 26389 29013 26407
rect 29031 26389 29049 26407
rect 29067 26389 29085 26407
rect 29103 26389 29121 26407
rect 29139 26389 29180 26407
rect 28920 26371 29180 26389
rect 28920 26353 28941 26371
rect 28959 26353 28977 26371
rect 28995 26353 29013 26371
rect 29031 26353 29049 26371
rect 29067 26353 29085 26371
rect 29103 26353 29121 26371
rect 29139 26353 29180 26371
rect 28920 26335 29180 26353
rect 28920 26317 28941 26335
rect 28959 26317 28977 26335
rect 28995 26317 29013 26335
rect 29031 26317 29049 26335
rect 29067 26317 29085 26335
rect 29103 26317 29121 26335
rect 29139 26317 29180 26335
rect 28920 26299 29180 26317
rect 28920 26281 28941 26299
rect 28959 26281 28977 26299
rect 28995 26281 29013 26299
rect 29031 26281 29049 26299
rect 29067 26281 29085 26299
rect 29103 26281 29121 26299
rect 29139 26281 29180 26299
rect 28920 26263 29180 26281
rect 28920 26245 28941 26263
rect 28959 26245 28977 26263
rect 28995 26245 29013 26263
rect 29031 26245 29049 26263
rect 29067 26245 29085 26263
rect 29103 26245 29121 26263
rect 29139 26245 29180 26263
rect 28920 26227 29180 26245
rect 28920 26209 28941 26227
rect 28959 26209 28977 26227
rect 28995 26209 29013 26227
rect 29031 26209 29049 26227
rect 29067 26209 29085 26227
rect 29103 26209 29121 26227
rect 29139 26209 29180 26227
rect 28920 26191 29180 26209
rect 28920 26173 28941 26191
rect 28959 26173 28977 26191
rect 28995 26173 29013 26191
rect 29031 26173 29049 26191
rect 29067 26173 29085 26191
rect 29103 26173 29121 26191
rect 29139 26173 29180 26191
rect 28920 26160 29180 26173
rect 28860 23813 28920 23840
rect 28860 23795 28881 23813
rect 28899 23795 28920 23813
rect 28860 23777 28920 23795
rect 28860 23759 28881 23777
rect 28899 23759 28920 23777
rect 28860 23741 28920 23759
rect 28860 23723 28881 23741
rect 28899 23723 28920 23741
rect 28860 23705 28920 23723
rect 28860 23687 28881 23705
rect 28899 23687 28920 23705
rect 28860 23380 28920 23687
rect 8820 23260 9260 23340
rect 28860 23300 29180 23380
rect 9200 22393 9260 23260
rect 9200 22375 9221 22393
rect 9239 22375 9260 22393
rect 9200 22357 9260 22375
rect 9200 22339 9221 22357
rect 9239 22339 9260 22357
rect 9200 22321 9260 22339
rect 9200 22303 9221 22321
rect 9239 22303 9260 22321
rect 9200 22285 9260 22303
rect 9200 22267 9221 22285
rect 9239 22267 9260 22285
rect 9200 22240 9260 22267
rect 28660 21893 28720 21920
rect 28660 21875 28681 21893
rect 28699 21875 28720 21893
rect 28660 21857 28720 21875
rect 28660 21839 28681 21857
rect 28699 21839 28720 21857
rect 28660 21821 28720 21839
rect 28660 21803 28681 21821
rect 28699 21803 28720 21821
rect 28660 21785 28720 21803
rect 28660 21767 28681 21785
rect 28699 21767 28720 21785
rect 9320 21293 9380 21320
rect 9320 21275 9341 21293
rect 9359 21275 9380 21293
rect 9320 21257 9380 21275
rect 9320 21239 9341 21257
rect 9359 21239 9380 21257
rect 9320 21221 9380 21239
rect 9320 21203 9341 21221
rect 9359 21203 9380 21221
rect 9320 21185 9380 21203
rect 9320 21167 9341 21185
rect 9359 21167 9380 21185
rect 9200 20713 9260 20740
rect 9200 20695 9221 20713
rect 9239 20695 9260 20713
rect 9200 20677 9260 20695
rect 9200 20659 9221 20677
rect 9239 20659 9260 20677
rect 9200 20641 9260 20659
rect 9200 20640 9221 20641
rect 8820 20623 9221 20640
rect 9239 20623 9260 20641
rect 8820 20605 9260 20623
rect 8820 20587 9221 20605
rect 9239 20587 9260 20605
rect 8820 20560 9260 20587
rect 9320 19593 9380 21167
rect 28660 20680 28720 21767
rect 28660 20600 29180 20680
rect 9320 19575 9341 19593
rect 9359 19575 9380 19593
rect 9320 19557 9380 19575
rect 9320 19539 9341 19557
rect 9359 19539 9380 19557
rect 9320 19521 9380 19539
rect 9320 19503 9341 19521
rect 9359 19503 9380 19521
rect 9320 19485 9380 19503
rect 9320 19467 9341 19485
rect 9359 19467 9380 19485
rect 9320 19440 9380 19467
rect 28540 20233 28600 20260
rect 28540 20215 28561 20233
rect 28579 20215 28600 20233
rect 28540 20197 28600 20215
rect 28540 20179 28561 20197
rect 28579 20179 28600 20197
rect 28540 20161 28600 20179
rect 28540 20143 28561 20161
rect 28579 20143 28600 20161
rect 28540 20125 28600 20143
rect 28540 20107 28561 20125
rect 28579 20107 28600 20125
rect 9440 19113 9500 19140
rect 9440 19095 9461 19113
rect 9479 19095 9500 19113
rect 9440 19077 9500 19095
rect 9440 19059 9461 19077
rect 9479 19059 9500 19077
rect 9440 19041 9500 19059
rect 9440 19023 9461 19041
rect 9479 19023 9500 19041
rect 9440 19005 9500 19023
rect 9440 18987 9461 19005
rect 9479 18987 9500 19005
rect 9320 18013 9380 18040
rect 9320 17995 9341 18013
rect 9359 17995 9380 18013
rect 9320 17977 9380 17995
rect 9320 17959 9341 17977
rect 9359 17959 9380 17977
rect 9320 17941 9380 17959
rect 9320 17940 9341 17941
rect 8820 17923 9341 17940
rect 9359 17923 9380 17941
rect 8820 17905 9380 17923
rect 8820 17887 9341 17905
rect 9359 17887 9380 17905
rect 8820 17860 9380 17887
rect 9440 17673 9500 18987
rect 28540 17980 28600 20107
rect 28540 17900 29180 17980
rect 9440 17655 9461 17673
rect 9479 17655 9500 17673
rect 9440 17637 9500 17655
rect 9440 17619 9461 17637
rect 9479 17619 9500 17637
rect 9440 17601 9500 17619
rect 9440 17583 9461 17601
rect 9479 17583 9500 17601
rect 9440 17565 9500 17583
rect 9440 17547 9461 17565
rect 9479 17547 9500 17565
rect 9440 17520 9500 17547
rect 28420 17633 28480 17660
rect 28420 17615 28441 17633
rect 28459 17615 28480 17633
rect 28420 17597 28480 17615
rect 28420 17579 28441 17597
rect 28459 17579 28480 17597
rect 28420 17561 28480 17579
rect 28420 17543 28441 17561
rect 28459 17543 28480 17561
rect 28420 17525 28480 17543
rect 28420 17507 28441 17525
rect 28459 17507 28480 17525
rect 9560 16653 9620 16680
rect 9560 16635 9581 16653
rect 9599 16635 9620 16653
rect 9560 16617 9620 16635
rect 9560 16599 9581 16617
rect 9599 16599 9620 16617
rect 9560 16581 9620 16599
rect 9560 16563 9581 16581
rect 9599 16563 9620 16581
rect 9560 16545 9620 16563
rect 9560 16527 9581 16545
rect 9599 16527 9620 16545
rect 9440 15313 9500 15340
rect 9440 15295 9461 15313
rect 9479 15295 9500 15313
rect 9440 15277 9500 15295
rect 9440 15259 9461 15277
rect 9479 15259 9500 15277
rect 9440 15241 9500 15259
rect 9440 15240 9461 15241
rect 8820 15223 9461 15240
rect 9479 15223 9500 15241
rect 8820 15205 9500 15223
rect 8820 15187 9461 15205
rect 9479 15187 9500 15205
rect 8820 15160 9500 15187
rect 9560 15013 9620 16527
rect 28420 15280 28480 17507
rect 28420 15200 29180 15280
rect 9560 14995 9581 15013
rect 9599 14995 9620 15013
rect 9560 14977 9620 14995
rect 9560 14959 9581 14977
rect 9599 14959 9620 14977
rect 9560 14941 9620 14959
rect 9560 14923 9581 14941
rect 9599 14923 9620 14941
rect 9560 14905 9620 14923
rect 9560 14887 9581 14905
rect 9599 14887 9620 14905
rect 9560 14860 9620 14887
rect 9560 12613 9620 12640
rect 9560 12595 9581 12613
rect 9599 12595 9620 12613
rect 9560 12577 9620 12595
rect 9560 12559 9581 12577
rect 9599 12559 9620 12577
rect 9560 12541 9620 12559
rect 9560 12540 9581 12541
rect 8820 12523 9581 12540
rect 9599 12523 9620 12541
rect 8820 12505 9620 12523
rect 8820 12487 9581 12505
rect 9599 12487 9620 12505
rect 8820 12460 9620 12487
rect 28420 12561 29180 12580
rect 28420 12543 28441 12561
rect 28459 12543 29180 12561
rect 28420 12525 29180 12543
rect 28420 12507 28441 12525
rect 28459 12507 29180 12525
rect 28420 12500 29180 12507
rect 28420 12489 28480 12500
rect 28420 12471 28441 12489
rect 28459 12471 28480 12489
rect 28420 12453 28480 12471
rect 28420 12435 28441 12453
rect 28459 12435 28480 12453
rect 28420 12417 28480 12435
rect 28420 12399 28441 12417
rect 28459 12399 28480 12417
rect 28420 12380 28480 12399
rect 28560 12013 29180 12040
rect 28560 11995 28581 12013
rect 28599 11995 29180 12013
rect 28560 11977 29180 11995
rect 28560 11959 28581 11977
rect 28599 11960 29180 11977
rect 28599 11959 28620 11960
rect 28560 11941 28620 11959
rect 28560 11923 28581 11941
rect 28599 11923 28620 11941
rect 28560 11905 28620 11923
rect 28560 11887 28581 11905
rect 28599 11887 28620 11905
rect 28560 11860 28620 11887
rect 8840 11547 9080 11560
rect 8840 11529 8861 11547
rect 8879 11529 8897 11547
rect 8915 11529 8933 11547
rect 8951 11529 8969 11547
rect 8987 11529 9005 11547
rect 9023 11529 9041 11547
rect 9059 11529 9080 11547
rect 8840 11511 9080 11529
rect 8840 11493 8861 11511
rect 8879 11493 8897 11511
rect 8915 11493 8933 11511
rect 8951 11493 8969 11511
rect 8987 11493 9005 11511
rect 9023 11493 9041 11511
rect 9059 11493 9080 11511
rect 8840 11475 9080 11493
rect 8840 11457 8861 11475
rect 8879 11457 8897 11475
rect 8915 11457 8933 11475
rect 8951 11457 8969 11475
rect 8987 11457 9005 11475
rect 9023 11457 9041 11475
rect 9059 11457 9080 11475
rect 8840 11439 9080 11457
rect 8840 11421 8861 11439
rect 8879 11421 8897 11439
rect 8915 11421 8933 11439
rect 8951 11421 8969 11439
rect 8987 11421 9005 11439
rect 9023 11421 9041 11439
rect 9059 11421 9080 11439
rect 8840 11403 9080 11421
rect 8840 11385 8861 11403
rect 8879 11385 8897 11403
rect 8915 11385 8933 11403
rect 8951 11385 8969 11403
rect 8987 11385 9005 11403
rect 9023 11385 9041 11403
rect 9059 11385 9080 11403
rect 8840 11367 9080 11385
rect 8840 11349 8861 11367
rect 8879 11349 8897 11367
rect 8915 11349 8933 11367
rect 8951 11349 8969 11367
rect 8987 11349 9005 11367
rect 9023 11349 9041 11367
rect 9059 11349 9080 11367
rect 8840 11331 9080 11349
rect 8840 11313 8861 11331
rect 8879 11313 8897 11331
rect 8915 11313 8933 11331
rect 8951 11313 8969 11331
rect 8987 11313 9005 11331
rect 9023 11313 9041 11331
rect 9059 11313 9080 11331
rect 8840 11295 9080 11313
rect 8840 11277 8861 11295
rect 8879 11277 8897 11295
rect 8915 11277 8933 11295
rect 8951 11277 8969 11295
rect 8987 11277 9005 11295
rect 9023 11277 9041 11295
rect 9059 11277 9080 11295
rect 8840 11259 9080 11277
rect 8840 11241 8861 11259
rect 8879 11241 8897 11259
rect 8915 11241 8933 11259
rect 8951 11241 8969 11259
rect 8987 11241 9005 11259
rect 9023 11241 9041 11259
rect 9059 11241 9080 11259
rect 8840 11223 9080 11241
rect 8840 11205 8861 11223
rect 8879 11205 8897 11223
rect 8915 11205 8933 11223
rect 8951 11205 8969 11223
rect 8987 11205 9005 11223
rect 9023 11205 9041 11223
rect 9059 11205 9080 11223
rect 8840 11187 9080 11205
rect 8840 11169 8861 11187
rect 8879 11169 8897 11187
rect 8915 11169 8933 11187
rect 8951 11169 8969 11187
rect 8987 11169 9005 11187
rect 9023 11169 9041 11187
rect 9059 11169 9080 11187
rect 8840 11151 9080 11169
rect 8840 11133 8861 11151
rect 8879 11133 8897 11151
rect 8915 11133 8933 11151
rect 8951 11133 8969 11151
rect 8987 11133 9005 11151
rect 9023 11133 9041 11151
rect 9059 11133 9080 11151
rect 8840 11115 9080 11133
rect 8840 11097 8861 11115
rect 8879 11097 8897 11115
rect 8915 11097 8933 11115
rect 8951 11097 8969 11115
rect 8987 11097 9005 11115
rect 9023 11097 9041 11115
rect 9059 11097 9080 11115
rect 8840 11079 9080 11097
rect 8840 11061 8861 11079
rect 8879 11061 8897 11079
rect 8915 11061 8933 11079
rect 8951 11061 8969 11079
rect 8987 11061 9005 11079
rect 9023 11061 9041 11079
rect 9059 11061 9080 11079
rect 8840 11043 9080 11061
rect 8840 11025 8861 11043
rect 8879 11025 8897 11043
rect 8915 11025 8933 11043
rect 8951 11025 8969 11043
rect 8987 11025 9005 11043
rect 9023 11025 9041 11043
rect 9059 11025 9080 11043
rect 8840 11007 9080 11025
rect 8840 10989 8861 11007
rect 8879 10989 8897 11007
rect 8915 10989 8933 11007
rect 8951 10989 8969 11007
rect 8987 10989 9005 11007
rect 9023 10989 9041 11007
rect 9059 10989 9080 11007
rect 8840 10971 9080 10989
rect 8840 10953 8861 10971
rect 8879 10953 8897 10971
rect 8915 10953 8933 10971
rect 8951 10953 8969 10971
rect 8987 10953 9005 10971
rect 9023 10953 9041 10971
rect 9059 10953 9080 10971
rect 8840 10935 9080 10953
rect 8840 10917 8861 10935
rect 8879 10917 8897 10935
rect 8915 10917 8933 10935
rect 8951 10917 8969 10935
rect 8987 10917 9005 10935
rect 9023 10917 9041 10935
rect 9059 10917 9080 10935
rect 8840 10899 9080 10917
rect 8840 10881 8861 10899
rect 8879 10881 8897 10899
rect 8915 10881 8933 10899
rect 8951 10881 8969 10899
rect 8987 10881 9005 10899
rect 9023 10881 9041 10899
rect 9059 10881 9080 10899
rect 8840 10863 9080 10881
rect 8840 10845 8861 10863
rect 8879 10845 8897 10863
rect 8915 10845 8933 10863
rect 8951 10845 8969 10863
rect 8987 10845 9005 10863
rect 9023 10845 9041 10863
rect 9059 10845 9080 10863
rect 8840 10827 9080 10845
rect 8840 10809 8861 10827
rect 8879 10809 8897 10827
rect 8915 10809 8933 10827
rect 8951 10809 8969 10827
rect 8987 10809 9005 10827
rect 9023 10809 9041 10827
rect 9059 10809 9080 10827
rect 8840 10791 9080 10809
rect 8840 10773 8861 10791
rect 8879 10773 8897 10791
rect 8915 10773 8933 10791
rect 8951 10773 8969 10791
rect 8987 10773 9005 10791
rect 9023 10773 9041 10791
rect 9059 10773 9080 10791
rect 8840 10755 9080 10773
rect 8840 10737 8861 10755
rect 8879 10737 8897 10755
rect 8915 10737 8933 10755
rect 8951 10737 8969 10755
rect 8987 10737 9005 10755
rect 9023 10737 9041 10755
rect 9059 10737 9080 10755
rect 8840 10719 9080 10737
rect 8840 10701 8861 10719
rect 8879 10701 8897 10719
rect 8915 10701 8933 10719
rect 8951 10701 8969 10719
rect 8987 10701 9005 10719
rect 9023 10701 9041 10719
rect 9059 10701 9080 10719
rect 8840 10683 9080 10701
rect 8840 10665 8861 10683
rect 8879 10665 8897 10683
rect 8915 10665 8933 10683
rect 8951 10665 8969 10683
rect 8987 10665 9005 10683
rect 9023 10665 9041 10683
rect 9059 10665 9080 10683
rect 8840 10647 9080 10665
rect 8840 10629 8861 10647
rect 8879 10629 8897 10647
rect 8915 10629 8933 10647
rect 8951 10629 8969 10647
rect 8987 10629 9005 10647
rect 9023 10629 9041 10647
rect 9059 10629 9080 10647
rect 8840 10611 9080 10629
rect 8840 10593 8861 10611
rect 8879 10593 8897 10611
rect 8915 10593 8933 10611
rect 8951 10593 8969 10611
rect 8987 10593 9005 10611
rect 9023 10593 9041 10611
rect 9059 10593 9080 10611
rect 8840 10575 9080 10593
rect 8840 10557 8861 10575
rect 8879 10557 8897 10575
rect 8915 10557 8933 10575
rect 8951 10557 8969 10575
rect 8987 10557 9005 10575
rect 9023 10557 9041 10575
rect 9059 10557 9080 10575
rect 8840 10539 9080 10557
rect 8840 10521 8861 10539
rect 8879 10521 8897 10539
rect 8915 10521 8933 10539
rect 8951 10521 8969 10539
rect 8987 10521 9005 10539
rect 9023 10521 9041 10539
rect 9059 10521 9080 10539
rect 8840 10503 9080 10521
rect 8840 10485 8861 10503
rect 8879 10485 8897 10503
rect 8915 10485 8933 10503
rect 8951 10485 8969 10503
rect 8987 10485 9005 10503
rect 9023 10485 9041 10503
rect 9059 10485 9080 10503
rect 8840 10467 9080 10485
rect 8840 10449 8861 10467
rect 8879 10449 8897 10467
rect 8915 10449 8933 10467
rect 8951 10449 8969 10467
rect 8987 10449 9005 10467
rect 9023 10449 9041 10467
rect 9059 10449 9080 10467
rect 8840 10431 9080 10449
rect 8840 10413 8861 10431
rect 8879 10413 8897 10431
rect 8915 10413 8933 10431
rect 8951 10413 8969 10431
rect 8987 10413 9005 10431
rect 9023 10413 9041 10431
rect 9059 10413 9080 10431
rect 8840 10395 9080 10413
rect 8840 10377 8861 10395
rect 8879 10377 8897 10395
rect 8915 10377 8933 10395
rect 8951 10377 8969 10395
rect 8987 10377 9005 10395
rect 9023 10377 9041 10395
rect 9059 10377 9080 10395
rect 8840 10359 9080 10377
rect 8840 10341 8861 10359
rect 8879 10341 8897 10359
rect 8915 10341 8933 10359
rect 8951 10341 8969 10359
rect 8987 10341 9005 10359
rect 9023 10341 9041 10359
rect 9059 10341 9080 10359
rect 8840 10323 9080 10341
rect 8840 10305 8861 10323
rect 8879 10305 8897 10323
rect 8915 10305 8933 10323
rect 8951 10305 8969 10323
rect 8987 10305 9005 10323
rect 9023 10305 9041 10323
rect 9059 10305 9080 10323
rect 8840 10287 9080 10305
rect 8840 10269 8861 10287
rect 8879 10269 8897 10287
rect 8915 10269 8933 10287
rect 8951 10269 8969 10287
rect 8987 10269 9005 10287
rect 9023 10269 9041 10287
rect 9059 10269 9080 10287
rect 8840 10251 9080 10269
rect 8840 10233 8861 10251
rect 8879 10233 8897 10251
rect 8915 10233 8933 10251
rect 8951 10233 8969 10251
rect 8987 10233 9005 10251
rect 9023 10233 9041 10251
rect 9059 10233 9080 10251
rect 8840 10220 9080 10233
rect 10240 9080 10320 10060
rect 11020 9200 11100 10060
rect 11440 9320 11520 10080
rect 12820 9440 12900 10060
rect 15640 9560 15720 10060
rect 18760 9680 18840 10060
rect 20140 9800 20220 10060
rect 20440 9920 20520 10060
rect 20440 9899 23340 9920
rect 20440 9881 23187 9899
rect 23205 9881 23223 9899
rect 23241 9881 23259 9899
rect 23277 9881 23295 9899
rect 23313 9881 23340 9899
rect 20440 9860 23340 9881
rect 25680 9899 28620 9920
rect 25680 9881 25707 9899
rect 25725 9881 25743 9899
rect 25761 9881 25779 9899
rect 25797 9881 25815 9899
rect 25833 9881 28467 9899
rect 28485 9881 28503 9899
rect 28521 9881 28539 9899
rect 28557 9881 28575 9899
rect 28593 9881 28620 9899
rect 25680 9860 28620 9881
rect 20140 9779 20320 9800
rect 20140 9761 20167 9779
rect 20185 9761 20203 9779
rect 20221 9761 20239 9779
rect 20257 9761 20275 9779
rect 20293 9761 20320 9779
rect 20140 9740 20320 9761
rect 23000 9779 25660 9800
rect 23000 9761 23027 9779
rect 23045 9761 23063 9779
rect 23081 9761 23099 9779
rect 23117 9761 23135 9779
rect 23153 9761 25507 9779
rect 25525 9761 25543 9779
rect 25561 9761 25579 9779
rect 25597 9761 25615 9779
rect 25633 9761 25660 9779
rect 23000 9740 25660 9761
rect 28060 9779 28240 9800
rect 28060 9761 28087 9779
rect 28105 9761 28123 9779
rect 28141 9761 28159 9779
rect 28177 9761 28195 9779
rect 28213 9761 28240 9779
rect 28060 9740 28240 9761
rect 18760 9659 18940 9680
rect 18760 9641 18787 9659
rect 18805 9641 18823 9659
rect 18841 9641 18859 9659
rect 18877 9641 18895 9659
rect 18913 9641 18940 9659
rect 18760 9620 18940 9641
rect 20380 9659 23000 9680
rect 20380 9641 20407 9659
rect 20425 9641 20443 9659
rect 20461 9641 20479 9659
rect 20497 9641 20515 9659
rect 20533 9641 22847 9659
rect 22865 9641 22883 9659
rect 22901 9641 22919 9659
rect 22937 9641 22955 9659
rect 22973 9641 23000 9659
rect 20380 9620 23000 9641
rect 25360 9659 25540 9680
rect 25360 9641 25387 9659
rect 25405 9641 25423 9659
rect 25441 9641 25459 9659
rect 25477 9641 25495 9659
rect 25513 9641 25540 9659
rect 25360 9620 25540 9641
rect 15640 9539 19160 9560
rect 15640 9521 19007 9539
rect 19025 9521 19043 9539
rect 19061 9521 19079 9539
rect 19097 9521 19115 9539
rect 19133 9521 19160 9539
rect 15640 9500 19160 9521
rect 22660 9539 22840 9560
rect 22660 9521 22687 9539
rect 22705 9521 22723 9539
rect 22741 9521 22759 9539
rect 22777 9521 22795 9539
rect 22813 9521 22840 9539
rect 22660 9500 22840 9521
rect 12820 9419 14800 9440
rect 12820 9401 14647 9419
rect 14665 9401 14683 9419
rect 14701 9401 14719 9419
rect 14737 9401 14755 9419
rect 14773 9401 14800 9419
rect 12820 9380 14800 9401
rect 17800 9419 17980 9440
rect 17800 9401 17827 9419
rect 17845 9401 17863 9419
rect 17881 9401 17899 9419
rect 17917 9401 17935 9419
rect 17953 9401 17980 9419
rect 17800 9380 17980 9401
rect 11440 9299 13100 9320
rect 11440 9281 12947 9299
rect 12965 9281 12983 9299
rect 13001 9281 13019 9299
rect 13037 9281 13055 9299
rect 13073 9281 13100 9299
rect 11440 9260 13100 9281
rect 15100 9299 15280 9320
rect 15100 9281 15127 9299
rect 15145 9281 15163 9299
rect 15181 9281 15199 9299
rect 15217 9281 15235 9299
rect 15253 9281 15280 9299
rect 15100 9260 15280 9281
rect 11020 9179 11200 9200
rect 11020 9161 11047 9179
rect 11065 9161 11083 9179
rect 11101 9161 11119 9179
rect 11137 9161 11155 9179
rect 11173 9161 11200 9179
rect 11020 9140 11200 9161
rect 12400 9179 12580 9200
rect 12400 9161 12427 9179
rect 12445 9161 12463 9179
rect 12481 9161 12499 9179
rect 12517 9161 12535 9179
rect 12553 9161 12580 9179
rect 12400 9140 12580 9161
rect 9800 9020 10320 9080
rect 9800 8820 9880 9020
rect 12500 8820 12580 9140
rect 15200 8820 15280 9260
rect 17900 8820 17980 9380
rect 22760 8820 22840 9500
rect 25460 8820 25540 9620
rect 28160 8820 28240 9740
<< m3contact >>
rect 11973 28985 11991 29003
rect 12009 28985 12027 29003
rect 11973 28949 11991 28967
rect 12009 28949 12027 28967
rect 11973 28913 11991 28931
rect 12009 28913 12027 28931
rect 11973 28877 11991 28895
rect 12009 28877 12027 28895
rect 12413 28905 12431 28923
rect 12449 28905 12467 28923
rect 12413 28869 12431 28887
rect 12449 28869 12467 28887
rect 12413 28833 12431 28851
rect 12449 28833 12467 28851
rect 12413 28797 12431 28815
rect 12449 28797 12467 28815
rect 22787 28701 22805 28719
rect 22823 28701 22841 28719
rect 22859 28701 22877 28719
rect 22895 28701 22913 28719
rect 24067 28701 24085 28719
rect 24103 28701 24121 28719
rect 24139 28701 24157 28719
rect 24175 28701 24193 28719
rect 21847 28581 21865 28599
rect 21883 28581 21901 28599
rect 21919 28581 21937 28599
rect 21955 28581 21973 28599
rect 23927 28581 23945 28599
rect 23963 28581 23981 28599
rect 23999 28581 24017 28599
rect 24035 28581 24053 28599
rect 17387 28461 17405 28479
rect 17423 28461 17441 28479
rect 17459 28461 17477 28479
rect 17495 28461 17513 28479
rect 19447 28461 19465 28479
rect 19483 28461 19501 28479
rect 19519 28461 19537 28479
rect 19555 28461 19573 28479
rect 14687 28341 14705 28359
rect 14723 28341 14741 28359
rect 14759 28341 14777 28359
rect 14795 28341 14813 28359
rect 17207 28341 17225 28359
rect 17243 28341 17261 28359
rect 17279 28341 17297 28359
rect 17315 28341 17333 28359
rect 24487 28701 24505 28719
rect 24523 28701 24541 28719
rect 24559 28701 24577 28719
rect 24595 28701 24613 28719
rect 25387 28701 25405 28719
rect 25423 28701 25441 28719
rect 25459 28701 25477 28719
rect 25495 28701 25513 28719
rect 25587 28581 25605 28599
rect 25623 28581 25641 28599
rect 25659 28581 25677 28599
rect 25695 28581 25713 28599
rect 28087 28581 28105 28599
rect 28123 28581 28141 28599
rect 28159 28581 28177 28599
rect 28195 28581 28213 28599
rect 28881 23795 28899 23813
rect 28881 23759 28899 23777
rect 28881 23723 28899 23741
rect 28881 23687 28899 23705
rect 9221 22375 9239 22393
rect 9221 22339 9239 22357
rect 9221 22303 9239 22321
rect 9221 22267 9239 22285
rect 28681 21875 28699 21893
rect 28681 21839 28699 21857
rect 28681 21803 28699 21821
rect 28681 21767 28699 21785
rect 9341 21275 9359 21293
rect 9341 21239 9359 21257
rect 9341 21203 9359 21221
rect 9341 21167 9359 21185
rect 9221 20695 9239 20713
rect 9221 20659 9239 20677
rect 9221 20623 9239 20641
rect 9221 20587 9239 20605
rect 9341 19575 9359 19593
rect 9341 19539 9359 19557
rect 9341 19503 9359 19521
rect 9341 19467 9359 19485
rect 28561 20215 28579 20233
rect 28561 20179 28579 20197
rect 28561 20143 28579 20161
rect 28561 20107 28579 20125
rect 9461 19095 9479 19113
rect 9461 19059 9479 19077
rect 9461 19023 9479 19041
rect 9461 18987 9479 19005
rect 9341 17995 9359 18013
rect 9341 17959 9359 17977
rect 9341 17923 9359 17941
rect 9341 17887 9359 17905
rect 9461 17655 9479 17673
rect 9461 17619 9479 17637
rect 9461 17583 9479 17601
rect 9461 17547 9479 17565
rect 28441 17615 28459 17633
rect 28441 17579 28459 17597
rect 28441 17543 28459 17561
rect 28441 17507 28459 17525
rect 9581 16635 9599 16653
rect 9581 16599 9599 16617
rect 9581 16563 9599 16581
rect 9581 16527 9599 16545
rect 9461 15295 9479 15313
rect 9461 15259 9479 15277
rect 9461 15223 9479 15241
rect 9461 15187 9479 15205
rect 9581 14995 9599 15013
rect 9581 14959 9599 14977
rect 9581 14923 9599 14941
rect 9581 14887 9599 14905
rect 9581 12595 9599 12613
rect 9581 12559 9599 12577
rect 9581 12523 9599 12541
rect 9581 12487 9599 12505
rect 28441 12543 28459 12561
rect 28441 12507 28459 12525
rect 28441 12471 28459 12489
rect 28441 12435 28459 12453
rect 28441 12399 28459 12417
rect 28581 11995 28599 12013
rect 28581 11959 28599 11977
rect 28581 11923 28599 11941
rect 28581 11887 28599 11905
rect 23187 9881 23205 9899
rect 23223 9881 23241 9899
rect 23259 9881 23277 9899
rect 23295 9881 23313 9899
rect 25707 9881 25725 9899
rect 25743 9881 25761 9899
rect 25779 9881 25797 9899
rect 25815 9881 25833 9899
rect 28467 9881 28485 9899
rect 28503 9881 28521 9899
rect 28539 9881 28557 9899
rect 28575 9881 28593 9899
rect 20167 9761 20185 9779
rect 20203 9761 20221 9779
rect 20239 9761 20257 9779
rect 20275 9761 20293 9779
rect 23027 9761 23045 9779
rect 23063 9761 23081 9779
rect 23099 9761 23117 9779
rect 23135 9761 23153 9779
rect 25507 9761 25525 9779
rect 25543 9761 25561 9779
rect 25579 9761 25597 9779
rect 25615 9761 25633 9779
rect 28087 9761 28105 9779
rect 28123 9761 28141 9779
rect 28159 9761 28177 9779
rect 28195 9761 28213 9779
rect 18787 9641 18805 9659
rect 18823 9641 18841 9659
rect 18859 9641 18877 9659
rect 18895 9641 18913 9659
rect 20407 9641 20425 9659
rect 20443 9641 20461 9659
rect 20479 9641 20497 9659
rect 20515 9641 20533 9659
rect 22847 9641 22865 9659
rect 22883 9641 22901 9659
rect 22919 9641 22937 9659
rect 22955 9641 22973 9659
rect 25387 9641 25405 9659
rect 25423 9641 25441 9659
rect 25459 9641 25477 9659
rect 25495 9641 25513 9659
rect 19007 9521 19025 9539
rect 19043 9521 19061 9539
rect 19079 9521 19097 9539
rect 19115 9521 19133 9539
rect 22687 9521 22705 9539
rect 22723 9521 22741 9539
rect 22759 9521 22777 9539
rect 22795 9521 22813 9539
rect 14647 9401 14665 9419
rect 14683 9401 14701 9419
rect 14719 9401 14737 9419
rect 14755 9401 14773 9419
rect 17827 9401 17845 9419
rect 17863 9401 17881 9419
rect 17899 9401 17917 9419
rect 17935 9401 17953 9419
rect 12947 9281 12965 9299
rect 12983 9281 13001 9299
rect 13019 9281 13037 9299
rect 13055 9281 13073 9299
rect 15127 9281 15145 9299
rect 15163 9281 15181 9299
rect 15199 9281 15217 9299
rect 15235 9281 15253 9299
rect 11047 9161 11065 9179
rect 11083 9161 11101 9179
rect 11119 9161 11137 9179
rect 11155 9161 11173 9179
rect 12427 9161 12445 9179
rect 12463 9161 12481 9179
rect 12499 9161 12517 9179
rect 12535 9161 12553 9179
<< metal3 >>
rect 11960 29003 12040 29020
rect 11960 28985 11973 29003
rect 11991 28985 12009 29003
rect 12027 28985 12040 29003
rect 11960 28967 12040 28985
rect 11960 28949 11973 28967
rect 11991 28949 12009 28967
rect 12027 28949 12040 28967
rect 11960 28940 12040 28949
rect 11960 28931 12480 28940
rect 11960 28913 11973 28931
rect 11991 28913 12009 28931
rect 12027 28923 12480 28931
rect 12027 28913 12413 28923
rect 11960 28905 12413 28913
rect 12431 28905 12449 28923
rect 12467 28905 12480 28923
rect 11960 28895 12480 28905
rect 11960 28877 11973 28895
rect 11991 28877 12009 28895
rect 12027 28887 12480 28895
rect 12027 28877 12413 28887
rect 11960 28869 12413 28877
rect 12431 28869 12449 28887
rect 12467 28869 12480 28887
rect 11960 28860 12480 28869
rect 12400 28851 12480 28860
rect 12400 28833 12413 28851
rect 12431 28833 12449 28851
rect 12467 28833 12480 28851
rect 12400 28815 12480 28833
rect 12400 28797 12413 28815
rect 12431 28797 12449 28815
rect 12467 28797 12480 28815
rect 12400 28780 12480 28797
rect 22760 28719 24220 28740
rect 22760 28701 22787 28719
rect 22805 28701 22823 28719
rect 22841 28701 22859 28719
rect 22877 28701 22895 28719
rect 22913 28701 24067 28719
rect 24085 28701 24103 28719
rect 24121 28701 24139 28719
rect 24157 28701 24175 28719
rect 24193 28701 24220 28719
rect 22760 28680 24220 28701
rect 24460 28719 25540 28740
rect 24460 28701 24487 28719
rect 24505 28701 24523 28719
rect 24541 28701 24559 28719
rect 24577 28701 24595 28719
rect 24613 28701 25387 28719
rect 25405 28701 25423 28719
rect 25441 28701 25459 28719
rect 25477 28701 25495 28719
rect 25513 28701 25540 28719
rect 24460 28680 25540 28701
rect 21820 28599 24080 28620
rect 21820 28581 21847 28599
rect 21865 28581 21883 28599
rect 21901 28581 21919 28599
rect 21937 28581 21955 28599
rect 21973 28581 23927 28599
rect 23945 28581 23963 28599
rect 23981 28581 23999 28599
rect 24017 28581 24035 28599
rect 24053 28581 24080 28599
rect 21820 28560 24080 28581
rect 25560 28599 28240 28620
rect 25560 28581 25587 28599
rect 25605 28581 25623 28599
rect 25641 28581 25659 28599
rect 25677 28581 25695 28599
rect 25713 28581 28087 28599
rect 28105 28581 28123 28599
rect 28141 28581 28159 28599
rect 28177 28581 28195 28599
rect 28213 28581 28240 28599
rect 25560 28560 28240 28581
rect 17360 28479 19600 28500
rect 17360 28461 17387 28479
rect 17405 28461 17423 28479
rect 17441 28461 17459 28479
rect 17477 28461 17495 28479
rect 17513 28461 19447 28479
rect 19465 28461 19483 28479
rect 19501 28461 19519 28479
rect 19537 28461 19555 28479
rect 19573 28461 19600 28479
rect 17360 28440 19600 28461
rect 14660 28359 17360 28380
rect 14660 28341 14687 28359
rect 14705 28341 14723 28359
rect 14741 28341 14759 28359
rect 14777 28341 14795 28359
rect 14813 28341 17207 28359
rect 17225 28341 17243 28359
rect 17261 28341 17279 28359
rect 17297 28341 17315 28359
rect 17333 28341 17360 28359
rect 14660 28320 17360 28341
rect 28020 23813 28920 23840
rect 28020 23795 28881 23813
rect 28899 23795 28920 23813
rect 28020 23777 28920 23795
rect 28020 23760 28881 23777
rect 28860 23759 28881 23760
rect 28899 23759 28920 23777
rect 28860 23741 28920 23759
rect 28860 23723 28881 23741
rect 28899 23723 28920 23741
rect 28860 23705 28920 23723
rect 28860 23687 28881 23705
rect 28899 23687 28920 23705
rect 28860 23660 28920 23687
rect 28020 23040 28720 23120
rect 9200 22393 9260 22420
rect 9200 22375 9221 22393
rect 9239 22375 9260 22393
rect 9200 22357 9260 22375
rect 9200 22339 9221 22357
rect 9239 22339 9260 22357
rect 9200 22321 9260 22339
rect 9200 22303 9221 22321
rect 9239 22303 9260 22321
rect 9200 22285 9260 22303
rect 9200 22267 9221 22285
rect 9239 22267 9260 22285
rect 9200 21740 9260 22267
rect 28020 22200 28600 22260
rect 9200 21660 9920 21740
rect 9200 21520 9920 21600
rect 9200 20713 9260 21520
rect 9320 21293 9920 21320
rect 9320 21275 9341 21293
rect 9359 21275 9920 21293
rect 9320 21257 9920 21275
rect 9320 21239 9341 21257
rect 9359 21240 9920 21257
rect 9359 21239 9380 21240
rect 9320 21221 9380 21239
rect 9320 21203 9341 21221
rect 9359 21203 9380 21221
rect 9320 21185 9380 21203
rect 9320 21167 9341 21185
rect 9359 21167 9380 21185
rect 9320 21140 9380 21167
rect 9200 20695 9221 20713
rect 9239 20695 9260 20713
rect 9200 20677 9260 20695
rect 9200 20659 9221 20677
rect 9239 20659 9260 20677
rect 9200 20641 9260 20659
rect 9200 20623 9221 20641
rect 9239 20623 9260 20641
rect 9200 20605 9260 20623
rect 9200 20587 9221 20605
rect 9239 20587 9260 20605
rect 9200 20560 9260 20587
rect 28540 20233 28600 22200
rect 28660 21893 28720 23040
rect 28660 21875 28681 21893
rect 28699 21875 28720 21893
rect 28660 21857 28720 21875
rect 28660 21839 28681 21857
rect 28699 21839 28720 21857
rect 28660 21821 28720 21839
rect 28660 21803 28681 21821
rect 28699 21803 28720 21821
rect 28660 21785 28720 21803
rect 28660 21767 28681 21785
rect 28699 21767 28720 21785
rect 28660 21740 28720 21767
rect 28540 20215 28561 20233
rect 28579 20215 28600 20233
rect 28540 20197 28600 20215
rect 28540 20179 28561 20197
rect 28579 20179 28600 20197
rect 28540 20161 28600 20179
rect 28540 20143 28561 20161
rect 28579 20143 28600 20161
rect 28540 20125 28600 20143
rect 28540 20107 28561 20125
rect 28579 20107 28600 20125
rect 28540 20080 28600 20107
rect 28020 19860 28480 19920
rect 9320 19593 9380 19620
rect 9320 19575 9341 19593
rect 9359 19575 9380 19593
rect 9320 19557 9380 19575
rect 9320 19539 9341 19557
rect 9359 19539 9380 19557
rect 9320 19521 9380 19539
rect 9320 19503 9341 19521
rect 9359 19503 9380 19521
rect 9320 19485 9380 19503
rect 9320 19467 9341 19485
rect 9359 19467 9380 19485
rect 9320 18013 9380 19467
rect 9440 19113 9920 19140
rect 9440 19095 9461 19113
rect 9479 19095 9920 19113
rect 9440 19077 9920 19095
rect 9440 19059 9461 19077
rect 9479 19060 9920 19077
rect 9479 19059 9500 19060
rect 9440 19041 9500 19059
rect 9440 19023 9461 19041
rect 9479 19023 9500 19041
rect 9440 19005 9500 19023
rect 9440 18987 9461 19005
rect 9479 18987 9500 19005
rect 9440 18960 9500 18987
rect 9320 17995 9341 18013
rect 9359 17995 9380 18013
rect 9320 17977 9380 17995
rect 9320 17959 9341 17977
rect 9359 17959 9380 17977
rect 9320 17941 9380 17959
rect 9320 17923 9341 17941
rect 9359 17923 9380 17941
rect 9320 17905 9380 17923
rect 9320 17887 9341 17905
rect 9359 17887 9380 17905
rect 9320 17860 9380 17887
rect 9440 17673 9500 17700
rect 9440 17655 9461 17673
rect 9479 17655 9500 17673
rect 9440 17637 9500 17655
rect 9440 17619 9461 17637
rect 9479 17619 9500 17637
rect 9440 17601 9500 17619
rect 9440 17583 9461 17601
rect 9479 17583 9500 17601
rect 9440 17565 9500 17583
rect 9440 17547 9461 17565
rect 9479 17547 9500 17565
rect 9440 15313 9500 17547
rect 28420 17633 28480 19860
rect 28420 17615 28441 17633
rect 28459 17615 28480 17633
rect 28420 17597 28480 17615
rect 28420 17579 28441 17597
rect 28459 17579 28480 17597
rect 28420 17561 28480 17579
rect 28420 17543 28441 17561
rect 28459 17543 28480 17561
rect 28420 17525 28480 17543
rect 28420 17507 28441 17525
rect 28459 17507 28480 17525
rect 28420 17480 28480 17507
rect 9560 16653 9920 16680
rect 9560 16635 9581 16653
rect 9599 16635 9920 16653
rect 9560 16617 9920 16635
rect 9560 16599 9581 16617
rect 9599 16600 9920 16617
rect 9599 16599 9620 16600
rect 9560 16581 9620 16599
rect 9560 16563 9581 16581
rect 9599 16563 9620 16581
rect 9560 16545 9620 16563
rect 9560 16527 9581 16545
rect 9599 16527 9620 16545
rect 9560 16500 9620 16527
rect 9440 15295 9461 15313
rect 9479 15295 9500 15313
rect 9440 15277 9500 15295
rect 9440 15259 9461 15277
rect 9479 15259 9500 15277
rect 9440 15241 9500 15259
rect 9440 15223 9461 15241
rect 9479 15223 9500 15241
rect 9440 15205 9500 15223
rect 9440 15187 9461 15205
rect 9479 15187 9500 15205
rect 9440 15160 9500 15187
rect 9560 15013 9620 15040
rect 9560 14995 9581 15013
rect 9599 14995 9620 15013
rect 9560 14977 9620 14995
rect 9560 14959 9581 14977
rect 9599 14959 9620 14977
rect 9560 14941 9620 14959
rect 9560 14923 9581 14941
rect 9599 14923 9620 14941
rect 9560 14905 9620 14923
rect 9560 14887 9581 14905
rect 9599 14887 9620 14905
rect 9560 12613 9620 14887
rect 9560 12595 9581 12613
rect 9599 12595 9620 12613
rect 9560 12577 9620 12595
rect 9560 12559 9581 12577
rect 9599 12559 9620 12577
rect 9560 12541 9620 12559
rect 9560 12523 9581 12541
rect 9599 12523 9620 12541
rect 9560 12505 9620 12523
rect 9560 12487 9581 12505
rect 9599 12487 9620 12505
rect 9560 12460 9620 12487
rect 28420 12561 28480 12580
rect 28420 12543 28441 12561
rect 28459 12543 28480 12561
rect 28420 12525 28480 12543
rect 28420 12507 28441 12525
rect 28459 12507 28480 12525
rect 28420 12489 28480 12507
rect 28420 12471 28441 12489
rect 28459 12471 28480 12489
rect 28420 12453 28480 12471
rect 28420 12435 28441 12453
rect 28459 12435 28480 12453
rect 28420 12417 28480 12435
rect 28420 12399 28441 12417
rect 28459 12399 28480 12417
rect 28420 11340 28480 12399
rect 28020 11280 28480 11340
rect 28560 12013 28620 12040
rect 28560 11995 28581 12013
rect 28599 11995 28620 12013
rect 28560 11977 28620 11995
rect 28560 11959 28581 11977
rect 28599 11959 28620 11977
rect 28560 11941 28620 11959
rect 28560 11923 28581 11941
rect 28599 11923 28620 11941
rect 28560 11905 28620 11923
rect 28560 11887 28581 11905
rect 28599 11887 28620 11905
rect 28560 9920 28620 11887
rect 23160 9899 25860 9920
rect 23160 9881 23187 9899
rect 23205 9881 23223 9899
rect 23241 9881 23259 9899
rect 23277 9881 23295 9899
rect 23313 9881 25707 9899
rect 25725 9881 25743 9899
rect 25761 9881 25779 9899
rect 25797 9881 25815 9899
rect 25833 9881 25860 9899
rect 23160 9860 25860 9881
rect 28440 9899 28620 9920
rect 28440 9881 28467 9899
rect 28485 9881 28503 9899
rect 28521 9881 28539 9899
rect 28557 9881 28575 9899
rect 28593 9881 28620 9899
rect 28440 9860 28620 9881
rect 20140 9779 23180 9800
rect 20140 9761 20167 9779
rect 20185 9761 20203 9779
rect 20221 9761 20239 9779
rect 20257 9761 20275 9779
rect 20293 9761 23027 9779
rect 23045 9761 23063 9779
rect 23081 9761 23099 9779
rect 23117 9761 23135 9779
rect 23153 9761 23180 9779
rect 20140 9740 23180 9761
rect 25480 9779 28240 9800
rect 25480 9761 25507 9779
rect 25525 9761 25543 9779
rect 25561 9761 25579 9779
rect 25597 9761 25615 9779
rect 25633 9761 28087 9779
rect 28105 9761 28123 9779
rect 28141 9761 28159 9779
rect 28177 9761 28195 9779
rect 28213 9761 28240 9779
rect 25480 9740 28240 9761
rect 18760 9659 20560 9680
rect 18760 9641 18787 9659
rect 18805 9641 18823 9659
rect 18841 9641 18859 9659
rect 18877 9641 18895 9659
rect 18913 9641 20407 9659
rect 20425 9641 20443 9659
rect 20461 9641 20479 9659
rect 20497 9641 20515 9659
rect 20533 9641 20560 9659
rect 18760 9620 20560 9641
rect 22820 9659 25540 9680
rect 22820 9641 22847 9659
rect 22865 9641 22883 9659
rect 22901 9641 22919 9659
rect 22937 9641 22955 9659
rect 22973 9641 25387 9659
rect 25405 9641 25423 9659
rect 25441 9641 25459 9659
rect 25477 9641 25495 9659
rect 25513 9641 25540 9659
rect 22820 9620 25540 9641
rect 18980 9539 22840 9560
rect 18980 9521 19007 9539
rect 19025 9521 19043 9539
rect 19061 9521 19079 9539
rect 19097 9521 19115 9539
rect 19133 9521 22687 9539
rect 22705 9521 22723 9539
rect 22741 9521 22759 9539
rect 22777 9521 22795 9539
rect 22813 9521 22840 9539
rect 18980 9500 22840 9521
rect 14620 9419 17980 9440
rect 14620 9401 14647 9419
rect 14665 9401 14683 9419
rect 14701 9401 14719 9419
rect 14737 9401 14755 9419
rect 14773 9401 17827 9419
rect 17845 9401 17863 9419
rect 17881 9401 17899 9419
rect 17917 9401 17935 9419
rect 17953 9401 17980 9419
rect 14620 9380 17980 9401
rect 12920 9299 15280 9320
rect 12920 9281 12947 9299
rect 12965 9281 12983 9299
rect 13001 9281 13019 9299
rect 13037 9281 13055 9299
rect 13073 9281 15127 9299
rect 15145 9281 15163 9299
rect 15181 9281 15199 9299
rect 15217 9281 15235 9299
rect 15253 9281 15280 9299
rect 12920 9260 15280 9281
rect 11020 9179 12580 9200
rect 11020 9161 11047 9179
rect 11065 9161 11083 9179
rect 11101 9161 11119 9179
rect 11137 9161 11155 9179
rect 11173 9161 12427 9179
rect 12445 9161 12463 9179
rect 12481 9161 12499 9179
rect 12517 9161 12535 9179
rect 12553 9161 12580 9179
rect 11020 9140 12580 9161
<< end >>
