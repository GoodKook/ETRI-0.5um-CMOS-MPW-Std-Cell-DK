magic
tech scmos
magscale 1 2
timestamp 1726541006
<< nwell >>
rect -12 154 132 272
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 60 14 64 54
rect 80 14 84 54
<< ptransistor >>
rect 20 166 24 246
rect 30 166 34 246
rect 60 166 64 246
rect 70 166 74 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 44 40 54
rect 24 14 26 44
rect 38 14 40 44
rect 44 14 46 54
rect 58 14 60 54
rect 64 26 66 54
rect 78 26 80 54
rect 64 14 80 26
rect 84 14 86 54
<< pdiffusion >>
rect 18 166 20 246
rect 24 166 30 246
rect 34 166 36 246
rect 58 166 60 246
rect 64 166 70 246
rect 74 166 76 246
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 44
rect 46 14 58 54
rect 66 26 78 54
rect 86 14 98 54
<< pdcontact >>
rect 6 166 18 246
rect 36 166 58 246
rect 76 166 88 246
<< psubstratepcontact >>
rect -6 -6 126 6
<< nsubstratencontact >>
rect -6 254 126 266
<< polysilicon >>
rect 20 246 24 250
rect 30 246 34 250
rect 60 246 64 250
rect 70 246 74 250
rect 20 162 24 166
rect 10 158 24 162
rect 30 162 34 166
rect 30 158 44 162
rect 10 128 16 158
rect 10 82 16 116
rect 40 102 44 158
rect 36 90 44 102
rect 10 76 24 82
rect 20 54 24 76
rect 40 54 44 90
rect 60 54 64 166
rect 70 162 74 166
rect 70 158 88 162
rect 84 128 88 158
rect 84 82 88 116
rect 80 76 88 82
rect 80 54 84 76
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
rect 80 10 84 14
<< polycontact >>
rect 4 116 16 128
rect 24 90 36 102
rect 84 116 96 128
rect 64 90 76 102
<< metal1 >>
rect -6 266 126 268
rect -6 252 126 254
rect 6 246 18 252
rect 76 246 88 252
rect 44 116 52 166
rect 43 86 50 102
rect 44 72 52 86
rect 44 64 74 72
rect 6 54 58 56
rect 68 54 74 64
rect 18 50 46 54
rect 58 14 86 20
rect 26 8 38 14
rect -6 6 126 8
rect -6 -8 126 -6
<< m2contact >>
rect 3 102 17 116
rect 23 102 37 116
rect 43 102 57 116
rect 63 102 77 116
rect 83 102 97 116
<< metal2 >>
rect 26 116 34 134
rect 66 116 74 134
rect 6 86 14 102
rect 46 86 54 102
rect 86 86 94 102
<< m1p >>
rect -6 252 126 268
rect -6 -8 126 8
<< m2p >>
rect 26 118 34 134
rect 66 118 74 134
rect 6 86 14 100
rect 46 86 54 100
rect 86 86 94 100
<< labels >>
rlabel metal1 -6 252 106 268 0 vdd
port 6 nsew power bidirectional abutment
rlabel metal1 -6 -8 106 8 0 gnd
port 7 nsew ground bidirectional abutment
rlabel metal2 10 90 10 90 1 A
port 1 n signal input
rlabel metal2 30 130 30 130 1 B
port 2 n signal input
rlabel metal2 50 88 50 88 5 Y
port 5 n signal output
rlabel metal2 70 130 70 130 1 D
port 4 n signal input
rlabel metal2 90 90 90 90 1 C
port 3 n signal input
<< properties >>
string FIXED_BBOX 0 0 120 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
