magic
tech scmos
magscale 1 30
timestamp 1725401611
<< checkpaint >>
rect 18300 186927 44800 197000
rect 13915 181835 44800 186927
rect 46919 186419 142100 190000
rect 46919 181835 143266 186419
rect 6771 176042 185015 181835
rect 6771 175958 328570 176042
rect 205 167042 328570 175958
rect 205 160774 185015 167042
rect 6771 143081 185015 160774
rect 0 142100 185015 143081
rect 0 102896 190000 142100
rect -13866 102380 190000 102896
rect -25613 89180 190000 102380
rect -24170 89077 190000 89180
rect -17472 83925 190000 89077
rect 0 47900 190000 83925
rect 6771 46919 190000 47900
rect 6771 32547 185015 46919
rect 6771 31724 186496 32547
rect -4457 10781 186496 31724
rect -4457 8670 185015 10781
rect -4457 7765 35955 8670
rect 205 1458 35955 7765
rect -600 -600 630 630
rect 46919 0 142100 8670
<< electrode >>
rect 91900 143200 111200 143800
<< genericcontact >>
rect 91900 143200 92900 143800
rect 110300 143200 111200 143800
<< metal1 >>
rect 89900 143200 92900 143800
rect 110300 143200 112900 143800
rect 139700 103800 145300 113200
rect 44700 91600 51100 98400
<< m2contact >>
rect 89500 143200 89900 143800
rect 112900 143200 113800 143800
rect 145300 103800 145800 113200
rect 44200 91600 44700 98400
<< metal2 >>
rect 59800 141300 60200 145900
rect 73300 142000 73700 145900
rect 86800 142700 87200 145900
rect 89500 143800 89900 145900
rect 48200 130200 48500 139700
rect 90800 137300 91100 139700
rect 96200 137300 96500 140400
rect 97400 137300 97700 141100
rect 106400 137300 106700 141800
rect 113800 139200 114200 145900
rect 113800 138900 117500 139200
rect 127300 138900 127700 145900
rect 117200 137300 117500 138900
rect 121700 138600 127700 138900
rect 140800 138600 141200 145900
rect 121700 137300 122000 138600
rect 125900 137300 126200 138000
rect 44100 129800 48500 130200
rect 142400 130000 145900 130400
rect 44100 116300 47600 116700
rect 143000 116500 145900 116900
rect 44100 102800 47600 103200
rect 143000 89500 145900 89900
rect 44100 75800 48300 76200
rect 142400 76000 145900 76400
rect 44100 62300 49000 62700
rect 141300 62500 145900 62900
rect 100100 53700 100400 54200
rect 103700 53100 104000 54300
rect 44100 48800 49700 49200
rect 59800 44100 60200 53100
rect 106700 52500 107000 54300
rect 73300 44100 73700 52500
rect 108200 51900 108500 54300
rect 86800 44100 87200 51900
rect 100300 44100 100700 51300
rect 110600 51200 110900 54300
rect 112400 51200 112700 54300
rect 114200 51800 114500 54300
rect 116000 52600 116300 54300
rect 103000 44100 103400 50600
rect 116500 44100 117000 50600
rect 130000 44100 130400 51200
rect 142100 49400 142500 52000
rect 142100 49000 145900 49400
<< m3contact >>
rect 86800 142100 87200 142700
rect 73300 141400 73700 142000
rect 106400 141800 106700 142400
rect 59800 140700 60200 141300
rect 97400 141100 97700 141700
rect 96200 140400 96500 141000
rect 48200 139700 48500 140300
rect 90800 139700 91100 140300
rect 125900 138000 126500 138300
rect 140800 138000 141200 138600
rect 141800 130000 142400 130400
rect 47600 116300 48200 116700
rect 142400 116500 143000 116900
rect 47600 102800 48200 103200
rect 142400 89500 143000 89900
rect 48300 75800 48900 76200
rect 141800 76000 142400 76400
rect 49000 62300 49600 62700
rect 140700 62500 141300 62900
rect 59800 53100 60200 53700
rect 99800 53400 100400 53700
rect 49700 48800 50300 49200
rect 73300 52500 73700 53100
rect 86800 51900 87200 52500
rect 106400 52200 107000 52500
rect 100300 51300 100700 51900
rect 107900 51600 108500 51900
rect 103000 50600 103400 51200
rect 110300 50900 110900 51200
rect 116000 52300 116600 52600
rect 142100 52000 142500 52600
rect 114200 51500 114800 51800
rect 130000 51200 130400 51800
rect 112400 50900 113000 51200
rect 116500 50600 117000 51200
<< metal3 >>
rect 87200 142100 106400 142400
rect 73700 141400 97400 141700
rect 60200 140700 96200 141000
rect 48500 140000 90800 140300
rect 126500 138000 140800 138300
rect 47900 107500 48200 116300
rect 141800 113200 142100 130000
rect 140300 112900 142100 113200
rect 47900 107200 50900 107500
rect 47900 106600 50900 106900
rect 47900 103200 48200 106600
rect 48600 104200 50900 104500
rect 48600 76200 48900 104200
rect 49300 103600 50900 103900
rect 49300 62700 49600 103600
rect 142400 103300 142700 116500
rect 50000 103000 50900 103300
rect 140300 103000 142700 103300
rect 50000 49200 50300 103000
rect 140300 102100 142700 102400
rect 140300 99400 142100 99700
rect 141800 76400 142100 99400
rect 142400 89900 142700 102100
rect 140300 68200 141000 68500
rect 140700 62900 141000 68200
rect 60200 53400 99800 53700
rect 73700 52800 104000 53100
rect 87200 52200 106400 52500
rect 116600 52300 142100 52600
rect 100700 51600 107900 51900
rect 114800 51500 130000 51800
rect 103400 50900 110300 51200
rect 113000 50900 116500 51200
use PIC  CIN_0
timestamp 1537935238
transform 1 0 129500 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_1
timestamp 1537935238
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_2
timestamp 1537935238
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_3
timestamp 1537935238
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_4
timestamp 1537935238
transform 1 0 48500 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_5
timestamp 1537935238
transform 0 1 18900 -1 0 141500
box -100 -9150 12100 25300
use PIC  CLK
timestamp 1537935238
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use POB8  CLK_OUT
timestamp 1537935238
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use fir_pe_Core  fir_pe_Core_0
timestamp 1725247039
transform 1 0 51960 0 1 54510
box -1110 -360 88410 82845
use PVSS  GND
timestamp 1537935238
transform 0 -1 171100 1 0 102500
box 0 -9150 12000 25300
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/pads_ETRI050
timestamp 1719894731
transform 0 -1 171100 -1 0 75646
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_1
timestamp 1719894731
transform 0 -1 171100 -1 0 62146
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_2
timestamp 1719894731
transform 0 -1 171100 -1 0 102646
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_3
timestamp 1719894731
transform 0 -1 171100 -1 0 89146
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_4
timestamp 1719894731
transform 0 -1 171100 -1 0 129646
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_5
timestamp 1719894731
transform 0 -1 171100 -1 0 116146
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_6
timestamp 1719894731
transform 1 0 73845 0 1 18900
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_7
timestamp 1719894731
transform 1 0 60345 0 1 18900
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_8
timestamp 1719894731
transform 1 0 100845 0 1 18900
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_9
timestamp 1719894731
transform 1 0 87345 0 1 18900
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_10
timestamp 1719894731
transform 1 0 127845 0 1 18900
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_11
timestamp 1719894731
transform 1 0 114345 0 1 18900
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_12
timestamp 1719894731
transform 0 1 18900 -1 0 75655
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_13
timestamp 1719894731
transform 0 1 18900 -1 0 62155
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_14
timestamp 1719894731
transform 0 1 18900 -1 0 102655
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_15
timestamp 1719894731
transform 0 1 18900 -1 0 89155
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_16
timestamp 1719894731
transform 1 0 73845 0 -1 171099
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_17
timestamp 1719894731
transform 0 1 18900 -1 0 116155
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_18
timestamp 1719894731
transform 0 1 18900 -1 0 129655
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_19
timestamp 1719894731
transform 1 0 60345 0 -1 171099
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_20
timestamp 1719894731
transform 1 0 100845 0 -1 171099
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_21
timestamp 1719894731
transform 1 0 87345 0 -1 171099
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_22
timestamp 1719894731
transform 1 0 127845 0 -1 171099
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_23
timestamp 1719894731
transform 1 0 114345 0 -1 171099
box 0 0 1800 25050
use IOFILLER50  IOFILLER50_0
timestamp 1537935238
transform 1 0 43585 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1537935238
transform 1 0 141465 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1537935238
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1537935238
transform 1 0 43585 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1537935238
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1537935238
transform 0 1 18900 -1 0 146415
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1537935238
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1537935238
transform 0 -1 171100 -1 0 146415
box -35 0 5035 25060
use MY_LOGO  MY_LOGO_0
timestamp 1724157349
transform 1 0 158160 0 1 11865
box 60 75 7170 3015
use PCORNER  PCORNER_0
timestamp 1537935238
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1537935238
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1537935238
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1537935238
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
use PIC  RDY
timestamp 1537935238
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use PVDD  VDD
timestamp 1537935238
transform 0 1 18900 -1 0 101000
box 0 -9150 12000 25300
use POB8  VLD
timestamp 1537935238
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use PIC  XIN_0
timestamp 1537935238
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use PIC  XIN_1
timestamp 1537935238
transform 0 1 18900 -1 0 74000
box -100 -9150 12100 25300
use PIC  XIN_2
timestamp 1537935238
transform 0 1 18900 -1 0 87500
box -100 -9150 12100 25300
use PIC  XIN_3
timestamp 1537935238
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use POB8  XOUT_0
timestamp 1537935238
transform 0 -1 171100 1 0 75500
box -100 -9150 12100 25300
use POB8  XOUT_1
timestamp 1537935238
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
use POB8  XOUT_2
timestamp 1537935238
transform 0 -1 171100 1 0 89000
box -100 -9150 12100 25300
use POB8  XOUT_3
timestamp 1537935238
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
use PIC  YIN_0
timestamp 1537935238
transform 1 0 48500 0 1 18900
box -100 -9150 12100 25300
use PIC  YIN_1
timestamp 1537935238
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use PIC  YIN_2
timestamp 1537935238
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use PIC  YIN_3
timestamp 1537935238
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use POB8  YOUT_0
timestamp 1537935238
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use POB8  YOUT_1
timestamp 1537935238
transform 1 0 129500 0 1 18900
box -100 -9150 12100 25300
use POB8  YOUT_2
timestamp 1537935238
transform 0 -1 171100 1 0 48500
box -100 -9150 12100 25300
use POB8  YOUT_3
timestamp 1537935238
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
<< end >>
