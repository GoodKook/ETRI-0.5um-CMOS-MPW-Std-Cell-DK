magic
tech scmos
magscale 1 2
timestamp 1702316108
<< nwell >>
rect -13 154 153 272
<< ntransistor >>
rect 18 14 22 54
rect 58 14 62 54
rect 78 14 82 54
rect 98 14 102 54
rect 118 14 122 54
<< ptransistor >>
rect 18 166 22 246
rect 58 166 62 246
rect 78 166 82 246
rect 98 166 102 246
rect 118 166 122 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 14 24 54
rect 56 14 58 54
rect 62 26 64 54
rect 76 26 78 54
rect 62 14 78 26
rect 82 14 84 54
rect 96 14 98 54
rect 102 48 118 54
rect 102 14 104 48
rect 116 14 118 48
rect 122 14 124 54
<< pdiffusion >>
rect 16 166 18 246
rect 22 166 24 246
rect 56 166 58 246
rect 62 234 78 246
rect 62 166 64 234
rect 76 166 78 234
rect 82 166 84 246
rect 96 166 98 246
rect 102 242 118 246
rect 102 180 104 242
rect 116 180 118 242
rect 102 166 118 180
rect 122 166 124 246
<< ndcontact >>
rect 4 14 16 54
rect 24 14 36 54
rect 44 14 56 54
rect 64 26 76 54
rect 84 14 96 54
rect 104 14 116 48
rect 124 14 136 54
<< pdcontact >>
rect 4 166 16 246
rect 24 166 36 246
rect 44 166 56 246
rect 64 166 76 234
rect 84 166 96 246
rect 104 180 116 242
rect 124 166 136 246
<< psubstratepcontact >>
rect -7 -6 147 6
<< nsubstratencontact >>
rect -7 254 147 266
<< polysilicon >>
rect 18 246 22 250
rect 58 246 62 250
rect 78 246 82 250
rect 98 246 102 250
rect 118 246 122 250
rect 18 60 22 166
rect 58 164 62 166
rect 78 164 82 166
rect 38 160 82 164
rect 98 164 102 166
rect 118 164 122 166
rect 98 160 122 164
rect 38 148 42 160
rect 118 60 122 160
rect 18 56 82 60
rect 18 54 22 56
rect 58 54 62 56
rect 78 54 82 56
rect 98 56 122 60
rect 98 54 102 56
rect 118 54 122 56
rect 18 10 22 14
rect 58 10 62 14
rect 78 10 82 14
rect 98 10 102 14
rect 118 10 122 14
<< polycontact >>
rect 6 105 18 117
rect 30 136 42 148
rect 122 105 134 117
<< metal1 >>
rect -7 266 147 268
rect -7 252 147 254
rect 4 246 16 252
rect 56 240 84 246
rect 104 242 116 252
rect 96 166 124 174
rect 30 148 36 166
rect 3 123 17 137
rect 6 117 17 123
rect 66 137 74 166
rect 30 54 36 136
rect 63 123 77 137
rect 123 123 137 137
rect 66 54 74 123
rect 123 117 134 123
rect 84 54 132 60
rect 56 14 84 20
rect 4 8 16 14
rect 104 8 116 14
rect -7 6 147 8
rect -7 -8 147 -6
<< m1p >>
rect -7 252 147 268
rect 3 123 17 137
rect 63 123 77 137
rect 123 123 137 137
rect -7 -8 147 8
<< labels >>
rlabel nsubstratencontact 70 260 70 260 0 vdd
port 4 nsew power bidirectional abutment
rlabel psubstratepcontact 70 0 70 0 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 10 130 10 130 0 EN
port 2 nsew signal input
rlabel metal1 70 131 70 131 0 Y
port 3 nsew signal output
rlabel metal1 131 130 131 130 0 A
port 1 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 140 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
