VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ALU_wrapper
  CLASS BLOCK ;
  FOREIGN ALU_wrapper ;
  ORIGIN 6.000 6.000 ;
  SIZE 783.000 BY 735.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 4.800 686.700 6.600 694.800 ;
        RECT 13.800 686.700 15.600 691.800 ;
        RECT 31.800 686.700 33.600 691.800 ;
        RECT 43.800 686.700 45.600 690.600 ;
        RECT 53.400 686.700 55.200 691.800 ;
        RECT 73.800 686.700 75.600 691.800 ;
        RECT 83.700 686.700 85.500 690.600 ;
        RECT 91.200 686.700 93.000 693.600 ;
        RECT 103.800 686.700 105.600 691.800 ;
        RECT 110.400 686.700 112.200 690.600 ;
        RECT 125.400 686.700 127.200 691.800 ;
        RECT 134.400 686.700 136.200 694.800 ;
        RECT 148.800 686.700 150.600 691.800 ;
        RECT 158.700 686.700 160.500 693.600 ;
        RECT 170.700 686.700 172.500 690.600 ;
        RECT 178.200 686.700 180.000 693.600 ;
        RECT 188.400 686.700 190.200 691.800 ;
        RECT 208.500 686.700 210.300 693.600 ;
        RECT 217.800 686.700 219.600 690.600 ;
        RECT 223.800 687.600 225.600 690.600 ;
        RECT 224.400 686.700 225.600 687.600 ;
        RECT 232.800 686.700 234.600 690.600 ;
        RECT 247.800 686.700 249.600 691.800 ;
        RECT 254.400 686.700 256.200 690.600 ;
        RECT 260.400 686.700 262.200 690.600 ;
        RECT 271.800 686.700 273.600 690.600 ;
        RECT 278.400 686.700 280.200 691.800 ;
        RECT 290.400 686.700 292.200 690.600 ;
        RECT 296.400 686.700 298.200 690.600 ;
        RECT 305.700 686.700 307.500 690.600 ;
        RECT 313.200 686.700 315.000 693.600 ;
        RECT 320.400 686.700 322.200 691.800 ;
        RECT 337.800 686.700 339.600 693.600 ;
        RECT 343.800 686.700 345.600 693.600 ;
        RECT 347.700 686.700 349.500 693.600 ;
        RECT 364.800 686.700 366.600 693.600 ;
        RECT 373.200 686.700 375.000 693.600 ;
        RECT 383.400 686.700 385.200 691.800 ;
        RECT 395.700 686.700 397.500 693.600 ;
        RECT 410.400 686.700 412.200 690.600 ;
        RECT 427.800 686.700 429.600 693.600 ;
        RECT 434.700 686.700 436.500 693.600 ;
        RECT 447.150 686.700 448.950 690.600 ;
        RECT 456.450 686.700 458.250 690.600 ;
        RECT 463.350 686.700 465.150 690.600 ;
        RECT 472.350 686.700 474.150 690.600 ;
        RECT 484.800 686.700 486.600 693.600 ;
        RECT 490.800 686.700 492.600 693.600 ;
        RECT 496.800 686.700 498.600 693.600 ;
        RECT 502.800 686.700 504.600 693.600 ;
        RECT 508.800 686.700 510.600 693.600 ;
        RECT 515.400 686.700 517.200 691.800 ;
        RECT 538.500 686.700 540.300 693.600 ;
        RECT 545.850 686.700 547.650 690.600 ;
        RECT 554.850 686.700 556.650 690.600 ;
        RECT 561.750 686.700 563.550 690.600 ;
        RECT 571.050 686.700 572.850 690.600 ;
        RECT 578.400 686.700 580.200 693.600 ;
        RECT 584.400 686.700 586.200 693.600 ;
        RECT 590.400 686.700 592.200 693.600 ;
        RECT 596.400 686.700 598.200 693.600 ;
        RECT 602.400 686.700 604.200 693.600 ;
        RECT 610.200 686.700 612.000 690.600 ;
        RECT 622.500 686.700 624.300 693.600 ;
        RECT 645.000 686.700 646.800 690.600 ;
        RECT 652.500 686.700 654.300 690.600 ;
        RECT 671.100 686.700 672.900 693.600 ;
        RECT 683.700 686.700 685.500 690.600 ;
        RECT 691.200 686.700 693.000 693.600 ;
        RECT 697.200 686.700 699.000 690.600 ;
        RECT 709.500 686.700 711.300 693.600 ;
        RECT 732.000 686.700 733.800 690.600 ;
        RECT 739.500 686.700 741.300 690.600 ;
        RECT 758.100 686.700 759.900 693.600 ;
        RECT 771.300 686.700 780.300 722.700 ;
        RECT 0.600 684.300 780.300 686.700 ;
        RECT 10.500 677.400 12.300 684.300 ;
        RECT 25.800 679.200 27.600 684.300 ;
        RECT 32.700 677.400 34.500 684.300 ;
        RECT 55.500 674.400 57.300 684.300 ;
        RECT 67.500 677.400 69.300 684.300 ;
        RECT 82.500 677.400 84.300 684.300 ;
        RECT 94.800 679.200 96.600 684.300 ;
        RECT 101.400 680.400 103.200 684.300 ;
        RECT 107.400 680.400 109.200 684.300 ;
        RECT 121.800 679.200 123.600 684.300 ;
        RECT 128.700 677.400 130.500 684.300 ;
        RECT 151.800 679.200 153.600 684.300 ;
        RECT 160.800 680.400 162.600 684.300 ;
        RECT 166.800 680.400 168.600 684.300 ;
        RECT 181.800 679.200 183.600 684.300 ;
        RECT 196.800 679.200 198.600 684.300 ;
        RECT 208.800 680.400 210.600 684.300 ;
        RECT 220.800 679.200 222.600 684.300 ;
        RECT 228.000 677.400 229.800 684.300 ;
        RECT 236.400 677.400 238.200 684.300 ;
        RECT 259.500 674.400 261.300 684.300 ;
        RECT 271.500 677.400 273.300 684.300 ;
        RECT 286.800 679.200 288.600 684.300 ;
        RECT 293.700 677.400 295.500 684.300 ;
        RECT 316.500 674.400 318.300 684.300 ;
        RECT 328.500 677.400 330.300 684.300 ;
        RECT 337.800 677.400 339.600 684.300 ;
        RECT 346.200 677.400 348.000 684.300 ;
        RECT 358.800 679.200 360.600 684.300 ;
        RECT 365.700 677.400 367.500 684.300 ;
        RECT 380.400 680.400 382.200 684.300 ;
        RECT 386.400 680.400 388.200 684.300 ;
        RECT 392.400 680.400 394.200 684.300 ;
        RECT 404.700 677.400 406.500 684.300 ;
        RECT 416.400 680.400 418.200 684.300 ;
        RECT 433.500 677.400 435.300 684.300 ;
        RECT 437.400 680.400 439.200 684.300 ;
        RECT 457.800 679.200 459.600 684.300 ;
        RECT 467.850 680.400 469.650 684.300 ;
        RECT 476.850 680.400 478.650 684.300 ;
        RECT 483.750 680.400 485.550 684.300 ;
        RECT 493.050 680.400 494.850 684.300 ;
        RECT 503.400 679.200 505.200 684.300 ;
        RECT 515.700 677.400 517.500 684.300 ;
        RECT 527.400 680.400 529.200 684.300 ;
        RECT 539.400 679.200 541.200 684.300 ;
        RECT 559.500 677.400 561.300 684.300 ;
        RECT 567.150 680.400 568.950 684.300 ;
        RECT 576.450 680.400 578.250 684.300 ;
        RECT 583.350 680.400 585.150 684.300 ;
        RECT 592.350 680.400 594.150 684.300 ;
        RECT 607.500 677.400 609.300 684.300 ;
        RECT 613.200 680.400 615.000 684.300 ;
        RECT 625.500 677.400 627.300 684.300 ;
        RECT 648.000 680.400 649.800 684.300 ;
        RECT 655.500 680.400 657.300 684.300 ;
        RECT 674.100 677.400 675.900 684.300 ;
        RECT 686.700 677.400 688.500 684.300 ;
        RECT 706.800 679.200 708.600 684.300 ;
        RECT 718.800 680.400 720.600 684.300 ;
        RECT 724.800 680.400 726.600 684.300 ;
        RECT 739.500 674.400 741.300 684.300 ;
        RECT 746.400 680.400 748.200 684.300 ;
        RECT 755.400 680.400 757.200 684.300 ;
        RECT 4.800 614.700 6.600 618.600 ;
        RECT 10.800 614.700 12.600 618.600 ;
        RECT 18.900 614.700 20.700 621.600 ;
        RECT 37.500 614.700 39.300 621.600 ;
        RECT 41.700 614.700 43.500 624.600 ;
        RECT 59.400 614.700 61.200 618.600 ;
        RECT 69.000 614.700 70.800 621.600 ;
        RECT 76.500 614.700 78.300 618.600 ;
        RECT 88.800 614.700 90.600 618.600 ;
        RECT 100.800 614.700 102.600 619.800 ;
        RECT 115.800 614.700 117.600 619.800 ;
        RECT 125.700 614.700 127.500 618.600 ;
        RECT 133.200 614.700 135.000 621.600 ;
        RECT 148.800 614.700 150.600 619.800 ;
        RECT 163.800 614.700 165.600 619.800 ;
        RECT 178.800 614.700 180.600 619.800 ;
        RECT 188.700 614.700 190.500 621.600 ;
        RECT 205.800 614.700 207.600 621.600 ;
        RECT 214.200 614.700 216.000 621.600 ;
        RECT 225.300 614.700 227.100 621.600 ;
        RECT 241.500 614.700 243.300 621.600 ;
        RECT 253.800 614.700 255.600 619.800 ;
        RECT 261.000 614.700 262.800 621.600 ;
        RECT 269.400 614.700 271.200 621.600 ;
        RECT 278.700 614.700 280.500 621.600 ;
        RECT 295.800 614.700 297.600 621.600 ;
        RECT 307.800 614.700 309.600 619.800 ;
        RECT 319.800 614.700 321.600 618.600 ;
        RECT 331.500 614.700 333.300 621.600 ;
        RECT 341.400 614.700 343.200 619.800 ;
        RECT 350.400 614.700 352.200 622.800 ;
        RECT 362.700 614.700 364.500 621.600 ;
        RECT 371.700 614.700 373.500 621.600 ;
        RECT 391.800 614.700 393.600 619.800 ;
        RECT 406.500 614.700 408.300 621.600 ;
        RECT 416.850 614.700 418.650 618.600 ;
        RECT 425.850 614.700 427.650 618.600 ;
        RECT 432.750 614.700 434.550 618.600 ;
        RECT 442.050 614.700 443.850 618.600 ;
        RECT 460.800 614.700 462.600 619.800 ;
        RECT 467.700 614.700 469.500 621.600 ;
        RECT 482.850 614.700 484.650 618.600 ;
        RECT 491.850 614.700 493.650 618.600 ;
        RECT 498.750 614.700 500.550 618.600 ;
        RECT 508.050 614.700 509.850 618.600 ;
        RECT 518.700 614.700 520.500 621.600 ;
        RECT 538.500 614.700 540.300 621.600 ;
        RECT 550.800 614.700 552.600 619.800 ;
        RECT 565.500 614.700 567.300 621.600 ;
        RECT 577.800 614.700 579.600 619.800 ;
        RECT 587.700 614.700 589.500 621.600 ;
        RECT 599.400 614.700 601.200 619.800 ;
        RECT 615.150 614.700 616.950 618.600 ;
        RECT 624.450 614.700 626.250 618.600 ;
        RECT 631.350 614.700 633.150 618.600 ;
        RECT 640.350 614.700 642.150 618.600 ;
        RECT 652.800 614.700 654.600 618.600 ;
        RECT 658.800 615.600 660.600 618.600 ;
        RECT 659.400 614.700 660.600 615.600 ;
        RECT 670.800 614.700 672.600 619.800 ;
        RECT 685.800 614.700 687.600 619.800 ;
        RECT 703.800 614.700 705.600 620.100 ;
        RECT 710.400 614.700 712.200 618.600 ;
        RECT 724.800 614.700 726.600 621.600 ;
        RECT 733.200 614.700 735.000 621.600 ;
        RECT 740.400 614.700 742.200 618.600 ;
        RECT 757.800 614.700 759.600 619.800 ;
        RECT 771.300 614.700 780.300 684.300 ;
        RECT 0.600 612.300 780.300 614.700 ;
        RECT 8.400 607.200 10.200 612.300 ;
        RECT 28.800 608.400 30.600 612.300 ;
        RECT 35.400 607.200 37.200 612.300 ;
        RECT 58.500 605.400 60.300 612.300 ;
        RECT 65.700 602.400 67.500 612.300 ;
        RECT 83.700 608.400 85.500 612.300 ;
        RECT 91.200 605.400 93.000 612.300 ;
        RECT 100.800 608.400 102.600 612.300 ;
        RECT 104.700 605.400 106.500 612.300 ;
        RECT 116.400 608.400 118.200 612.300 ;
        RECT 130.500 605.400 132.300 612.300 ;
        RECT 143.700 605.400 145.500 612.300 ;
        RECT 160.500 605.400 162.300 612.300 ;
        RECT 166.800 608.400 168.600 612.300 ;
        RECT 172.800 608.400 174.600 612.300 ;
        RECT 181.800 608.400 183.600 612.300 ;
        RECT 185.700 605.400 187.500 612.300 ;
        RECT 205.800 607.200 207.600 612.300 ;
        RECT 213.000 605.400 214.800 612.300 ;
        RECT 221.400 605.400 223.200 612.300 ;
        RECT 230.700 605.400 232.500 612.300 ;
        RECT 248.400 607.200 250.200 612.300 ;
        RECT 270.300 605.400 272.100 612.300 ;
        RECT 289.500 602.400 291.300 612.300 ;
        RECT 301.800 607.200 303.600 612.300 ;
        RECT 308.400 608.400 310.200 612.300 ;
        RECT 314.400 608.400 316.200 612.300 ;
        RECT 328.800 608.400 330.600 612.300 ;
        RECT 335.400 607.200 337.200 612.300 ;
        RECT 347.400 608.400 349.200 612.300 ;
        RECT 364.800 608.400 366.600 612.300 ;
        RECT 368.400 608.400 370.200 612.300 ;
        RECT 381.150 608.400 382.950 612.300 ;
        RECT 390.450 608.400 392.250 612.300 ;
        RECT 397.350 608.400 399.150 612.300 ;
        RECT 406.350 608.400 408.150 612.300 ;
        RECT 416.850 608.400 418.650 612.300 ;
        RECT 425.850 608.400 427.650 612.300 ;
        RECT 432.750 608.400 434.550 612.300 ;
        RECT 442.050 608.400 443.850 612.300 ;
        RECT 449.700 605.400 451.500 612.300 ;
        RECT 469.800 607.200 471.600 612.300 ;
        RECT 476.400 608.400 478.200 612.300 ;
        RECT 490.500 605.400 492.300 612.300 ;
        RECT 502.500 605.400 504.300 612.300 ;
        RECT 520.500 605.400 522.300 612.300 ;
        RECT 532.800 607.200 534.600 612.300 ;
        RECT 542.850 608.400 544.650 612.300 ;
        RECT 551.850 608.400 553.650 612.300 ;
        RECT 558.750 608.400 560.550 612.300 ;
        RECT 568.050 608.400 569.850 612.300 ;
        RECT 579.150 608.400 580.950 612.300 ;
        RECT 588.450 608.400 590.250 612.300 ;
        RECT 595.350 608.400 597.150 612.300 ;
        RECT 604.350 608.400 606.150 612.300 ;
        RECT 616.800 608.400 618.600 612.300 ;
        RECT 628.500 605.400 630.300 612.300 ;
        RECT 635.700 605.400 637.500 612.300 ;
        RECT 649.800 608.400 651.600 612.300 ;
        RECT 655.800 608.400 657.600 612.300 ;
        RECT 660.000 605.400 661.800 612.300 ;
        RECT 667.500 608.400 669.300 612.300 ;
        RECT 677.400 607.200 679.200 612.300 ;
        RECT 694.800 608.400 696.600 612.300 ;
        RECT 698.400 608.400 700.200 612.300 ;
        RECT 704.400 608.400 706.200 612.300 ;
        RECT 710.400 608.400 712.200 612.300 ;
        RECT 722.400 608.400 724.200 612.300 ;
        RECT 728.400 608.400 730.200 612.300 ;
        RECT 737.400 607.200 739.200 612.300 ;
        RECT 750.000 605.400 751.800 612.300 ;
        RECT 757.500 608.400 759.300 612.300 ;
        RECT 7.500 542.700 9.300 549.600 ;
        RECT 25.800 542.700 27.600 547.800 ;
        RECT 35.400 542.700 37.200 547.800 ;
        RECT 50.700 542.700 52.500 546.600 ;
        RECT 58.200 542.700 60.000 549.600 ;
        RECT 65.400 542.700 67.200 547.800 ;
        RECT 78.000 542.700 79.800 549.600 ;
        RECT 85.500 542.700 87.300 546.600 ;
        RECT 100.800 542.700 102.600 547.800 ;
        RECT 115.800 542.700 117.600 547.800 ;
        RECT 128.400 542.700 130.200 547.800 ;
        RECT 148.800 542.700 150.600 547.800 ;
        RECT 158.700 542.700 160.500 546.600 ;
        RECT 166.200 542.700 168.000 549.600 ;
        RECT 173.400 542.700 175.200 547.800 ;
        RECT 193.500 542.700 195.300 549.600 ;
        RECT 199.800 542.700 201.600 546.600 ;
        RECT 205.800 542.700 207.600 546.600 ;
        RECT 220.500 542.700 222.300 549.600 ;
        RECT 232.800 542.700 234.600 547.800 ;
        RECT 240.000 542.700 241.800 549.600 ;
        RECT 248.400 542.700 250.200 549.600 ;
        RECT 257.700 542.700 259.500 549.600 ;
        RECT 275.400 542.700 277.200 547.800 ;
        RECT 294.300 542.700 296.100 549.600 ;
        RECT 307.800 542.700 309.600 549.600 ;
        RECT 314.400 542.700 316.200 547.800 ;
        RECT 331.500 542.700 333.300 549.600 ;
        RECT 341.850 542.700 343.650 546.600 ;
        RECT 350.850 542.700 352.650 546.600 ;
        RECT 357.750 542.700 359.550 546.600 ;
        RECT 367.050 542.700 368.850 546.600 ;
        RECT 374.400 542.700 376.200 546.600 ;
        RECT 386.400 542.700 388.200 547.800 ;
        RECT 401.700 542.700 403.500 549.600 ;
        RECT 421.800 542.700 423.600 547.800 ;
        RECT 434.400 542.700 436.200 547.800 ;
        RECT 454.500 542.700 456.300 549.600 ;
        RECT 462.150 542.700 463.950 546.600 ;
        RECT 471.450 542.700 473.250 546.600 ;
        RECT 478.350 542.700 480.150 546.600 ;
        RECT 487.350 542.700 489.150 546.600 ;
        RECT 500.700 542.700 502.500 549.600 ;
        RECT 514.500 542.700 516.300 549.600 ;
        RECT 526.500 542.700 528.300 549.600 ;
        RECT 536.850 542.700 538.650 546.600 ;
        RECT 545.850 542.700 547.650 546.600 ;
        RECT 552.750 542.700 554.550 546.600 ;
        RECT 562.050 542.700 563.850 546.600 ;
        RECT 572.700 542.700 574.500 549.600 ;
        RECT 592.800 542.700 594.600 547.800 ;
        RECT 599.400 542.700 601.200 546.600 ;
        RECT 605.400 542.700 607.200 546.600 ;
        RECT 617.400 542.700 619.200 547.800 ;
        RECT 629.400 542.700 631.200 546.600 ;
        RECT 646.800 542.700 648.600 546.600 ;
        RECT 653.700 542.700 655.500 549.600 ;
        RECT 665.400 542.700 667.200 546.600 ;
        RECT 671.400 542.700 673.200 546.600 ;
        RECT 678.000 542.700 679.800 549.600 ;
        RECT 686.400 542.700 688.200 549.600 ;
        RECT 698.400 542.700 700.200 547.800 ;
        RECT 710.700 542.700 712.500 552.600 ;
        RECT 727.800 542.700 729.600 549.600 ;
        RECT 733.800 542.700 735.600 549.600 ;
        RECT 744.900 542.700 746.700 549.600 ;
        RECT 771.300 542.700 780.300 612.300 ;
        RECT 0.600 540.300 780.300 542.700 ;
        RECT 10.500 533.400 12.300 540.300 ;
        RECT 23.700 536.400 25.500 540.300 ;
        RECT 31.200 533.400 33.000 540.300 ;
        RECT 43.800 536.400 45.600 540.300 ;
        RECT 55.800 535.200 57.600 540.300 ;
        RECT 70.500 533.400 72.300 540.300 ;
        RECT 82.800 535.200 84.600 540.300 ;
        RECT 97.800 535.200 99.600 540.300 ;
        RECT 104.700 533.400 106.500 540.300 ;
        RECT 117.000 533.400 118.800 540.300 ;
        RECT 124.500 536.400 126.300 540.300 ;
        RECT 136.800 536.400 138.600 540.300 ;
        RECT 143.700 536.400 145.500 540.300 ;
        RECT 151.200 533.400 153.000 540.300 ;
        RECT 155.400 536.400 157.200 540.300 ;
        RECT 165.000 533.400 166.800 540.300 ;
        RECT 172.500 536.400 174.300 540.300 ;
        RECT 185.400 535.200 187.200 540.300 ;
        RECT 200.400 536.400 202.200 540.300 ;
        RECT 206.400 536.400 208.200 540.300 ;
        RECT 212.400 536.400 214.200 540.300 ;
        RECT 218.400 536.400 220.200 540.300 ;
        RECT 226.800 536.400 228.600 540.300 ;
        RECT 232.800 536.400 234.600 540.300 ;
        RECT 237.000 533.400 238.800 540.300 ;
        RECT 245.400 533.400 247.200 540.300 ;
        RECT 254.700 533.400 256.500 540.300 ;
        RECT 273.300 533.400 275.100 540.300 ;
        RECT 289.800 535.200 291.600 540.300 ;
        RECT 297.000 533.400 298.800 540.300 ;
        RECT 305.400 533.400 307.200 540.300 ;
        RECT 317.700 533.400 319.500 540.300 ;
        RECT 333.900 533.400 335.700 540.300 ;
        RECT 347.400 535.200 349.200 540.300 ;
        RECT 362.400 536.400 364.200 540.300 ;
        RECT 368.400 536.400 370.200 540.300 ;
        RECT 382.800 535.200 384.600 540.300 ;
        RECT 389.700 533.400 391.500 540.300 ;
        RECT 412.800 535.200 414.600 540.300 ;
        RECT 419.400 536.400 421.200 540.300 ;
        RECT 428.700 533.400 430.500 540.300 ;
        RECT 443.700 536.400 445.500 540.300 ;
        RECT 451.200 533.400 453.000 540.300 ;
        RECT 458.400 535.200 460.200 540.300 ;
        RECT 470.700 533.400 472.500 540.300 ;
        RECT 485.850 536.400 487.650 540.300 ;
        RECT 494.850 536.400 496.650 540.300 ;
        RECT 501.750 536.400 503.550 540.300 ;
        RECT 511.050 536.400 512.850 540.300 ;
        RECT 521.400 535.200 523.200 540.300 ;
        RECT 533.700 533.400 535.500 540.300 ;
        RECT 548.700 533.400 550.500 540.300 ;
        RECT 560.400 535.200 562.200 540.300 ;
        RECT 575.850 536.400 577.650 540.300 ;
        RECT 584.850 536.400 586.650 540.300 ;
        RECT 591.750 536.400 593.550 540.300 ;
        RECT 601.050 536.400 602.850 540.300 ;
        RECT 614.400 535.200 616.200 540.300 ;
        RECT 626.700 533.400 628.500 540.300 ;
        RECT 641.700 533.400 643.500 540.300 ;
        RECT 653.700 533.400 655.500 540.300 ;
        RECT 665.700 533.400 667.500 540.300 ;
        RECT 679.800 533.400 681.600 540.300 ;
        RECT 685.800 533.400 687.600 540.300 ;
        RECT 691.800 533.400 693.600 540.300 ;
        RECT 697.800 533.400 699.600 540.300 ;
        RECT 703.800 533.400 705.600 540.300 ;
        RECT 712.800 536.400 714.600 540.300 ;
        RECT 716.400 536.400 718.200 540.300 ;
        RECT 722.400 536.400 724.200 540.300 ;
        RECT 728.700 533.400 730.500 540.300 ;
        RECT 743.400 536.400 745.200 540.300 ;
        RECT 757.500 533.400 759.300 540.300 ;
        RECT 10.800 470.700 12.600 474.600 ;
        RECT 22.500 470.700 24.300 477.600 ;
        RECT 32.700 470.700 34.500 474.600 ;
        RECT 40.200 470.700 42.000 477.600 ;
        RECT 55.500 470.700 57.300 480.600 ;
        RECT 67.500 470.700 69.300 477.600 ;
        RECT 71.700 470.700 73.500 480.600 ;
        RECT 89.400 470.700 91.200 475.800 ;
        RECT 109.500 470.700 111.300 477.600 ;
        RECT 121.800 470.700 123.600 475.800 ;
        RECT 134.400 470.700 136.200 475.800 ;
        RECT 154.800 470.700 156.600 475.800 ;
        RECT 169.800 470.700 171.600 475.800 ;
        RECT 176.400 470.700 178.200 474.600 ;
        RECT 188.700 470.700 190.500 474.600 ;
        RECT 196.200 470.700 198.000 477.600 ;
        RECT 200.700 470.700 202.500 477.600 ;
        RECT 215.400 470.700 217.200 474.600 ;
        RECT 227.400 470.700 229.200 476.100 ;
        RECT 253.800 470.700 255.600 475.800 ;
        RECT 265.800 470.700 267.600 474.600 ;
        RECT 271.800 470.700 273.600 474.600 ;
        RECT 280.800 470.700 282.600 474.600 ;
        RECT 286.800 470.700 288.600 474.600 ;
        RECT 295.800 470.700 297.600 477.600 ;
        RECT 304.200 470.700 306.000 477.600 ;
        RECT 311.850 470.700 313.650 474.600 ;
        RECT 320.850 470.700 322.650 474.600 ;
        RECT 327.750 470.700 329.550 474.600 ;
        RECT 337.050 470.700 338.850 474.600 ;
        RECT 347.700 470.700 349.500 477.600 ;
        RECT 356.700 470.700 358.500 477.600 ;
        RECT 376.800 470.700 378.600 475.800 ;
        RECT 394.800 470.700 396.600 475.800 ;
        RECT 408.300 470.700 410.100 477.600 ;
        RECT 421.800 470.700 423.600 477.600 ;
        RECT 428.850 470.700 430.650 474.600 ;
        RECT 437.850 470.700 439.650 474.600 ;
        RECT 444.750 470.700 446.550 474.600 ;
        RECT 454.050 470.700 455.850 474.600 ;
        RECT 463.800 470.700 465.600 477.600 ;
        RECT 469.800 470.700 471.600 477.600 ;
        RECT 475.800 470.700 477.600 477.600 ;
        RECT 481.800 470.700 483.600 477.600 ;
        RECT 487.800 470.700 489.600 477.600 ;
        RECT 499.800 470.700 501.600 475.800 ;
        RECT 511.800 470.700 513.600 474.600 ;
        RECT 515.700 470.700 517.500 477.600 ;
        RECT 530.700 470.700 532.500 474.600 ;
        RECT 538.200 470.700 540.000 477.600 ;
        RECT 553.500 470.700 555.300 480.600 ;
        RECT 557.400 470.700 559.200 474.600 ;
        RECT 563.400 470.700 565.200 474.600 ;
        RECT 569.700 470.700 571.500 477.600 ;
        RECT 582.000 470.700 583.800 477.600 ;
        RECT 590.400 470.700 592.200 477.600 ;
        RECT 607.500 470.700 609.300 477.600 ;
        RECT 614.400 470.700 616.200 474.600 ;
        RECT 620.400 470.700 622.200 474.600 ;
        RECT 631.800 470.700 633.600 474.600 ;
        RECT 641.400 470.700 643.200 475.800 ;
        RECT 664.800 470.700 666.600 476.100 ;
        RECT 671.400 470.700 673.200 474.600 ;
        RECT 677.400 470.700 679.200 474.600 ;
        RECT 683.700 470.700 685.500 477.600 ;
        RECT 703.800 470.700 705.600 475.800 ;
        RECT 713.400 470.700 715.200 475.800 ;
        RECT 725.400 470.700 727.200 474.600 ;
        RECT 731.400 470.700 733.200 474.600 ;
        RECT 745.800 470.700 747.600 474.600 ;
        RECT 751.800 471.600 753.600 474.600 ;
        RECT 752.400 470.700 753.600 471.600 ;
        RECT 759.900 470.700 761.700 477.600 ;
        RECT 771.300 470.700 780.300 540.300 ;
        RECT 0.600 468.300 780.300 470.700 ;
        RECT 7.800 464.400 9.600 468.300 ;
        RECT 19.800 463.200 21.600 468.300 ;
        RECT 30.900 461.400 32.700 468.300 ;
        RECT 55.500 458.400 57.300 468.300 ;
        RECT 59.400 464.400 61.200 468.300 ;
        RECT 73.800 464.400 75.600 468.300 ;
        RECT 80.700 458.400 82.500 468.300 ;
        RECT 98.400 464.400 100.200 468.300 ;
        RECT 115.500 461.400 117.300 468.300 ;
        RECT 119.700 458.400 121.500 468.300 ;
        RECT 137.400 464.400 139.200 468.300 ;
        RECT 149.400 463.200 151.200 468.300 ;
        RECT 164.700 458.400 166.500 468.300 ;
        RECT 181.800 464.400 183.600 468.300 ;
        RECT 187.800 464.400 189.600 468.300 ;
        RECT 191.400 464.400 193.200 468.300 ;
        RECT 197.400 464.400 199.200 468.300 ;
        RECT 206.700 461.400 208.500 468.300 ;
        RECT 218.400 464.400 220.200 468.300 ;
        RECT 224.400 464.400 226.200 468.300 ;
        RECT 230.400 464.400 232.200 468.300 ;
        RECT 236.400 464.400 238.200 468.300 ;
        RECT 246.900 461.400 248.700 468.300 ;
        RECT 259.800 464.400 261.600 468.300 ;
        RECT 265.800 464.400 267.600 468.300 ;
        RECT 272.400 464.400 274.200 468.300 ;
        RECT 278.400 464.400 280.200 468.300 ;
        RECT 287.400 464.400 289.200 468.300 ;
        RECT 296.700 461.400 298.500 468.300 ;
        RECT 308.400 464.400 310.200 468.300 ;
        RECT 318.000 461.400 319.800 468.300 ;
        RECT 326.400 461.400 328.200 468.300 ;
        RECT 336.000 461.400 337.800 468.300 ;
        RECT 343.500 464.400 345.300 468.300 ;
        RECT 353.700 464.400 355.500 468.300 ;
        RECT 361.200 461.400 363.000 468.300 ;
        RECT 368.850 464.400 370.650 468.300 ;
        RECT 377.850 464.400 379.650 468.300 ;
        RECT 384.750 464.400 386.550 468.300 ;
        RECT 394.050 464.400 395.850 468.300 ;
        RECT 407.700 464.400 409.500 468.300 ;
        RECT 415.200 461.400 417.000 468.300 ;
        RECT 422.400 463.200 424.200 468.300 ;
        RECT 436.800 461.400 438.600 468.300 ;
        RECT 442.800 461.400 444.600 468.300 ;
        RECT 448.800 461.400 450.600 468.300 ;
        RECT 454.800 461.400 456.600 468.300 ;
        RECT 460.800 461.400 462.600 468.300 ;
        RECT 475.500 461.400 477.300 468.300 ;
        RECT 487.500 461.400 489.300 468.300 ;
        RECT 499.500 461.400 501.300 468.300 ;
        RECT 503.700 458.400 505.500 468.300 ;
        RECT 529.500 458.400 531.300 468.300 ;
        RECT 541.800 464.400 543.600 468.300 ;
        RECT 556.800 463.200 558.600 468.300 ;
        RECT 563.400 464.400 565.200 468.300 ;
        RECT 575.400 463.200 577.200 468.300 ;
        RECT 601.500 458.400 603.300 468.300 ;
        RECT 608.700 464.400 610.500 468.300 ;
        RECT 616.200 461.400 618.000 468.300 ;
        RECT 625.800 461.400 627.600 468.300 ;
        RECT 634.200 461.400 636.000 468.300 ;
        RECT 646.500 461.400 648.300 468.300 ;
        RECT 650.400 464.400 652.200 468.300 ;
        RECT 662.400 463.200 664.200 468.300 ;
        RECT 685.500 458.400 687.300 468.300 ;
        RECT 697.800 464.400 699.600 468.300 ;
        RECT 702.000 461.400 703.800 468.300 ;
        RECT 709.500 464.400 711.300 468.300 ;
        RECT 719.400 464.400 721.200 468.300 ;
        RECT 725.400 464.400 727.200 468.300 ;
        RECT 734.400 467.400 735.600 468.300 ;
        RECT 734.400 464.400 736.200 467.400 ;
        RECT 740.400 464.400 742.200 468.300 ;
        RECT 752.400 463.200 754.200 468.300 ;
        RECT 7.800 398.700 9.600 402.600 ;
        RECT 19.800 398.700 21.600 403.800 ;
        RECT 32.400 398.700 34.200 403.800 ;
        RECT 55.500 398.700 57.300 405.600 ;
        RECT 70.500 398.700 72.300 408.600 ;
        RECT 74.700 398.700 76.500 408.600 ;
        RECT 97.500 398.700 99.300 405.600 ;
        RECT 101.700 398.700 103.500 408.600 ;
        RECT 124.500 398.700 126.300 405.600 ;
        RECT 135.900 398.700 137.700 405.600 ;
        RECT 149.400 398.700 151.200 403.800 ;
        RECT 161.700 398.700 163.500 405.600 ;
        RECT 173.700 398.700 175.500 408.600 ;
        RECT 188.700 398.700 190.500 405.600 ;
        RECT 203.400 398.700 205.200 402.600 ;
        RECT 215.400 398.700 217.200 403.800 ;
        RECT 230.400 398.700 232.200 403.800 ;
        RECT 245.400 398.700 247.200 402.600 ;
        RECT 254.700 398.700 256.500 405.600 ;
        RECT 269.400 398.700 271.200 403.800 ;
        RECT 284.700 398.700 286.500 402.600 ;
        RECT 292.200 398.700 294.000 405.600 ;
        RECT 307.800 398.700 309.600 403.800 ;
        RECT 322.800 398.700 324.600 403.800 ;
        RECT 337.800 398.700 339.600 403.800 ;
        RECT 344.700 398.700 346.500 405.600 ;
        RECT 359.700 398.700 361.500 402.600 ;
        RECT 367.200 398.700 369.000 405.600 ;
        RECT 379.800 398.700 381.600 403.800 ;
        RECT 391.800 398.700 393.600 405.600 ;
        RECT 397.800 398.700 399.600 405.600 ;
        RECT 406.800 398.700 408.600 405.600 ;
        RECT 415.200 398.700 417.000 405.600 ;
        RECT 419.400 398.700 421.200 402.600 ;
        RECT 431.700 398.700 433.500 405.600 ;
        RECT 445.500 398.700 447.300 405.600 ;
        RECT 463.500 398.700 465.300 405.600 ;
        RECT 472.800 398.700 474.600 402.600 ;
        RECT 484.800 398.700 486.600 403.800 ;
        RECT 505.800 398.700 507.600 402.600 ;
        RECT 511.800 398.700 513.900 402.600 ;
        RECT 529.800 398.700 531.600 403.800 ;
        RECT 536.400 398.700 538.200 402.600 ;
        RECT 548.700 398.700 550.500 405.600 ;
        RECT 571.500 398.700 573.300 408.600 ;
        RECT 578.700 398.700 580.500 402.600 ;
        RECT 586.200 398.700 588.000 405.600 ;
        RECT 598.800 398.700 600.600 403.800 ;
        RECT 608.400 398.700 610.200 403.800 ;
        RECT 631.500 398.700 633.300 408.600 ;
        RECT 636.000 398.700 637.800 405.600 ;
        RECT 643.500 398.700 645.300 402.600 ;
        RECT 651.000 398.700 652.800 405.600 ;
        RECT 659.400 398.700 661.200 405.600 ;
        RECT 676.500 398.700 678.300 405.600 ;
        RECT 683.700 398.700 685.500 402.600 ;
        RECT 691.200 398.700 693.000 405.600 ;
        RECT 695.700 398.700 697.500 408.600 ;
        RECT 713.700 398.700 715.500 402.600 ;
        RECT 721.200 398.700 723.000 405.600 ;
        RECT 725.700 398.700 727.500 408.600 ;
        RECT 740.700 398.700 742.500 408.600 ;
        RECT 771.300 398.700 780.300 468.300 ;
        RECT 0.600 396.300 780.300 398.700 ;
        RECT 7.800 392.400 9.600 396.300 ;
        RECT 14.400 395.400 15.600 396.300 ;
        RECT 13.800 392.400 15.600 395.400 ;
        RECT 25.500 389.400 27.300 396.300 ;
        RECT 32.700 389.400 34.500 396.300 ;
        RECT 44.400 392.400 46.200 396.300 ;
        RECT 61.800 391.200 63.600 396.300 ;
        RECT 73.800 392.400 75.600 396.300 ;
        RECT 81.000 389.400 82.800 396.300 ;
        RECT 88.500 392.400 90.300 396.300 ;
        RECT 95.700 386.400 97.500 396.300 ;
        RECT 110.700 386.400 112.500 396.300 ;
        RECT 130.800 392.400 132.600 396.300 ;
        RECT 142.800 392.400 144.600 396.300 ;
        RECT 149.400 395.400 150.600 396.300 ;
        RECT 148.800 392.400 150.600 395.400 ;
        RECT 152.700 386.400 154.500 396.300 ;
        RECT 181.800 392.400 183.600 396.300 ;
        RECT 187.800 392.400 189.900 396.300 ;
        RECT 194.400 392.400 196.200 396.300 ;
        RECT 209.400 391.200 211.200 396.300 ;
        RECT 224.400 391.200 226.200 396.300 ;
        RECT 242.700 392.400 244.500 396.300 ;
        RECT 250.200 389.400 252.000 396.300 ;
        RECT 262.800 391.200 264.600 396.300 ;
        RECT 274.800 389.400 276.600 396.300 ;
        RECT 283.200 389.400 285.000 396.300 ;
        RECT 295.800 392.400 297.600 396.300 ;
        RECT 303.150 392.400 304.950 396.300 ;
        RECT 312.450 392.400 314.250 396.300 ;
        RECT 319.350 392.400 321.150 396.300 ;
        RECT 328.350 392.400 330.150 396.300 ;
        RECT 338.700 392.400 340.500 396.300 ;
        RECT 346.200 389.400 348.000 396.300 ;
        RECT 358.800 389.400 360.600 396.300 ;
        RECT 367.200 389.400 369.000 396.300 ;
        RECT 376.800 392.400 378.600 396.300 ;
        RECT 383.850 392.400 385.650 396.300 ;
        RECT 392.850 392.400 394.650 396.300 ;
        RECT 399.750 392.400 401.550 396.300 ;
        RECT 409.050 392.400 410.850 396.300 ;
        RECT 419.850 392.400 421.650 396.300 ;
        RECT 428.850 392.400 430.650 396.300 ;
        RECT 435.750 392.400 437.550 396.300 ;
        RECT 445.050 392.400 446.850 396.300 ;
        RECT 460.800 391.200 462.600 396.300 ;
        RECT 470.700 392.400 472.500 396.300 ;
        RECT 478.200 389.400 480.000 396.300 ;
        RECT 482.700 386.400 484.500 396.300 ;
        RECT 500.400 392.400 502.200 396.300 ;
        RECT 516.900 389.400 518.700 396.300 ;
        RECT 532.800 392.400 534.600 396.300 ;
        RECT 547.500 386.400 549.300 396.300 ;
        RECT 565.500 386.400 567.300 396.300 ;
        RECT 577.800 391.200 579.600 396.300 ;
        RECT 590.400 391.200 592.200 396.300 ;
        RECT 602.400 392.400 604.200 396.300 ;
        RECT 622.500 386.400 624.300 396.300 ;
        RECT 626.700 386.400 628.500 396.300 ;
        RECT 652.500 386.400 654.300 396.300 ;
        RECT 661.800 392.400 663.600 396.300 ;
        RECT 673.800 391.200 675.600 396.300 ;
        RECT 686.700 392.400 688.500 396.300 ;
        RECT 694.200 389.400 696.000 396.300 ;
        RECT 709.500 386.400 711.300 396.300 ;
        RECT 719.400 391.200 721.200 396.300 ;
        RECT 736.800 392.400 738.600 396.300 ;
        RECT 743.400 391.200 745.200 396.300 ;
        RECT 10.800 326.700 12.600 330.600 ;
        RECT 17.400 326.700 19.200 331.800 ;
        RECT 34.800 326.700 36.600 330.600 ;
        RECT 40.800 327.600 42.600 330.600 ;
        RECT 41.400 326.700 42.600 327.600 ;
        RECT 51.900 326.700 53.700 333.600 ;
        RECT 62.700 326.700 64.500 336.600 ;
        RECT 77.700 326.700 79.500 336.600 ;
        RECT 95.400 326.700 97.200 331.800 ;
        RECT 121.500 326.700 123.300 336.600 ;
        RECT 125.400 326.700 127.200 330.600 ;
        RECT 135.000 326.700 136.800 333.600 ;
        RECT 142.500 326.700 144.300 330.600 ;
        RECT 152.400 326.700 154.200 331.800 ;
        RECT 172.800 326.700 174.600 330.600 ;
        RECT 181.800 326.700 183.600 330.600 ;
        RECT 187.800 326.700 189.600 330.600 ;
        RECT 196.800 326.700 198.600 330.600 ;
        RECT 203.700 326.700 205.500 330.600 ;
        RECT 211.200 326.700 213.000 333.600 ;
        RECT 215.400 326.700 217.200 330.600 ;
        RECT 221.400 326.700 223.200 330.600 ;
        RECT 232.800 326.700 234.600 333.600 ;
        RECT 241.200 326.700 243.000 333.600 ;
        RECT 250.800 326.700 252.600 330.600 ;
        RECT 258.150 326.700 259.950 330.600 ;
        RECT 267.450 326.700 269.250 330.600 ;
        RECT 274.350 326.700 276.150 330.600 ;
        RECT 283.350 326.700 285.150 330.600 ;
        RECT 293.700 326.700 295.500 333.600 ;
        RECT 313.800 326.700 315.600 331.800 ;
        RECT 325.800 326.700 327.600 333.600 ;
        RECT 334.200 326.700 336.000 333.600 ;
        RECT 343.800 326.700 345.600 330.600 ;
        RECT 351.150 326.700 352.950 330.600 ;
        RECT 360.450 326.700 362.250 330.600 ;
        RECT 367.350 326.700 369.150 330.600 ;
        RECT 376.350 326.700 378.150 330.600 ;
        RECT 390.900 326.700 392.700 333.600 ;
        RECT 412.500 326.700 414.300 333.600 ;
        RECT 424.800 326.700 426.600 330.600 ;
        RECT 431.400 326.700 433.200 331.800 ;
        RECT 451.500 326.700 453.300 333.600 ;
        RECT 463.800 326.700 465.600 330.600 ;
        RECT 467.700 326.700 469.500 333.600 ;
        RECT 479.400 326.700 481.200 330.600 ;
        RECT 485.400 326.700 487.200 330.600 ;
        RECT 505.500 326.700 507.300 336.600 ;
        RECT 517.800 326.700 519.600 331.800 ;
        RECT 527.400 326.700 529.200 331.800 ;
        RECT 540.000 326.700 541.800 333.600 ;
        RECT 547.500 326.700 549.300 330.600 ;
        RECT 562.800 326.700 564.600 331.800 ;
        RECT 583.800 326.700 585.600 330.600 ;
        RECT 589.800 326.700 591.900 330.600 ;
        RECT 596.400 326.700 598.200 330.600 ;
        RECT 608.700 326.700 610.500 330.600 ;
        RECT 616.200 326.700 618.000 333.600 ;
        RECT 623.700 326.700 625.500 336.600 ;
        RECT 641.400 326.700 643.200 331.800 ;
        RECT 656.700 326.700 658.500 330.600 ;
        RECT 664.200 326.700 666.000 333.600 ;
        RECT 679.500 326.700 681.300 336.600 ;
        RECT 697.500 326.700 699.300 336.600 ;
        RECT 715.500 326.700 717.300 336.600 ;
        RECT 730.800 326.700 732.600 331.800 ;
        RECT 740.400 326.700 742.200 331.800 ;
        RECT 752.700 326.700 754.500 336.600 ;
        RECT 771.300 326.700 780.300 396.300 ;
        RECT 0.600 324.300 780.300 326.700 ;
        RECT 10.800 320.400 12.600 324.300 ;
        RECT 22.500 317.400 24.300 324.300 ;
        RECT 26.700 317.400 28.500 324.300 ;
        RECT 41.700 314.400 43.500 324.300 ;
        RECT 56.700 317.400 58.500 324.300 ;
        RECT 76.800 319.200 78.600 324.300 ;
        RECT 83.700 317.400 85.500 324.300 ;
        RECT 95.400 323.400 96.600 324.300 ;
        RECT 95.400 320.400 97.200 323.400 ;
        RECT 101.400 320.400 103.200 324.300 ;
        RECT 121.500 317.400 123.300 324.300 ;
        RECT 136.500 314.400 138.300 324.300 ;
        RECT 140.400 320.400 142.200 324.300 ;
        RECT 146.400 320.400 148.200 324.300 ;
        RECT 158.700 320.400 160.500 324.300 ;
        RECT 166.200 317.400 168.000 324.300 ;
        RECT 176.700 320.400 178.500 324.300 ;
        RECT 184.200 317.400 186.000 324.300 ;
        RECT 191.400 319.200 193.200 324.300 ;
        RECT 203.700 317.400 205.500 324.300 ;
        RECT 216.000 317.400 217.800 324.300 ;
        RECT 224.400 317.400 226.200 324.300 ;
        RECT 237.000 317.400 238.800 324.300 ;
        RECT 244.500 320.400 246.300 324.300 ;
        RECT 259.800 319.200 261.600 324.300 ;
        RECT 269.400 319.200 271.200 324.300 ;
        RECT 281.400 320.400 283.200 324.300 ;
        RECT 301.500 314.400 303.300 324.300 ;
        RECT 307.800 320.400 309.600 324.300 ;
        RECT 313.800 320.400 315.600 324.300 ;
        RECT 320.400 319.200 322.200 324.300 ;
        RECT 335.700 317.400 337.500 324.300 ;
        RECT 347.700 317.400 349.500 324.300 ;
        RECT 359.700 317.400 361.500 324.300 ;
        RECT 375.900 317.400 377.700 324.300 ;
        RECT 392.700 317.400 394.500 324.300 ;
        RECT 404.700 317.400 406.500 324.300 ;
        RECT 421.800 319.200 423.600 324.300 ;
        RECT 439.500 317.400 441.300 324.300 ;
        RECT 443.400 320.400 445.200 324.300 ;
        RECT 452.700 314.400 454.500 324.300 ;
        RECT 467.700 317.400 469.500 324.300 ;
        RECT 479.700 314.400 481.500 324.300 ;
        RECT 502.500 317.400 504.300 324.300 ;
        RECT 510.900 317.400 512.700 324.300 ;
        RECT 529.500 317.400 531.300 324.300 ;
        RECT 536.700 320.400 538.500 324.300 ;
        RECT 544.200 317.400 546.000 324.300 ;
        RECT 556.500 317.400 558.300 324.300 ;
        RECT 571.500 314.400 573.300 324.300 ;
        RECT 575.400 320.400 577.200 324.300 ;
        RECT 592.800 319.200 594.600 324.300 ;
        RECT 605.400 319.200 607.200 324.300 ;
        RECT 623.700 320.400 625.500 324.300 ;
        RECT 631.200 317.400 633.000 324.300 ;
        RECT 649.500 314.400 651.300 324.300 ;
        RECT 664.500 314.400 666.300 324.300 ;
        RECT 671.700 320.400 673.500 324.300 ;
        RECT 679.200 317.400 681.000 324.300 ;
        RECT 697.500 314.400 699.300 324.300 ;
        RECT 701.700 317.400 703.500 324.300 ;
        RECT 724.500 314.400 726.300 324.300 ;
        RECT 729.000 317.400 730.800 324.300 ;
        RECT 736.500 320.400 738.300 324.300 ;
        RECT 747.000 317.400 748.800 324.300 ;
        RECT 754.500 320.400 756.300 324.300 ;
        RECT 10.800 254.700 12.600 259.800 ;
        RECT 25.500 254.700 27.300 261.600 ;
        RECT 32.700 254.700 34.500 264.600 ;
        RECT 55.500 254.700 57.300 261.600 ;
        RECT 59.700 254.700 61.500 264.600 ;
        RECT 77.700 254.700 79.500 258.600 ;
        RECT 85.200 254.700 87.000 261.600 ;
        RECT 92.700 254.700 94.500 261.600 ;
        RECT 109.800 254.700 111.600 258.600 ;
        RECT 115.800 254.700 117.600 258.600 ;
        RECT 127.800 254.700 129.600 259.800 ;
        RECT 137.400 254.700 139.200 260.100 ;
        RECT 155.700 254.700 157.500 258.600 ;
        RECT 163.200 254.700 165.000 261.600 ;
        RECT 167.400 254.700 169.200 258.600 ;
        RECT 173.400 254.700 175.200 258.600 ;
        RECT 179.400 254.700 181.200 258.600 ;
        RECT 185.400 254.700 187.200 258.600 ;
        RECT 194.700 254.700 196.500 261.600 ;
        RECT 206.700 254.700 208.500 261.600 ;
        RECT 221.700 254.700 223.500 261.600 ;
        RECT 233.700 254.700 235.500 261.600 ;
        RECT 245.400 254.700 247.200 261.600 ;
        RECT 260.700 254.700 262.500 258.600 ;
        RECT 268.200 254.700 270.000 261.600 ;
        RECT 280.500 254.700 282.300 261.600 ;
        RECT 289.800 254.700 291.600 261.600 ;
        RECT 295.800 254.700 297.600 261.600 ;
        RECT 299.400 254.700 301.200 261.600 ;
        RECT 313.800 254.700 315.600 261.600 ;
        RECT 320.700 254.700 322.500 261.600 ;
        RECT 340.500 254.700 342.300 264.600 ;
        RECT 352.500 254.700 354.300 261.600 ;
        RECT 362.700 254.700 364.500 258.600 ;
        RECT 370.200 254.700 372.000 261.600 ;
        RECT 374.700 254.700 376.500 261.600 ;
        RECT 389.700 254.700 391.500 261.600 ;
        RECT 405.300 254.700 407.100 261.600 ;
        RECT 413.400 254.700 415.200 261.600 ;
        RECT 428.700 254.700 430.500 261.600 ;
        RECT 444.300 254.700 446.100 261.600 ;
        RECT 456.900 254.700 458.700 261.600 ;
        RECT 475.800 254.700 477.600 261.600 ;
        RECT 484.200 254.700 486.000 261.600 ;
        RECT 495.300 254.700 497.100 261.600 ;
        RECT 503.700 254.700 505.500 261.600 ;
        RECT 518.400 254.700 520.200 259.800 ;
        RECT 530.700 254.700 532.500 261.600 ;
        RECT 545.400 254.700 547.200 259.800 ;
        RECT 557.400 254.700 559.200 258.600 ;
        RECT 563.400 254.700 565.200 258.600 ;
        RECT 572.700 254.700 574.500 261.600 ;
        RECT 589.500 254.700 591.300 261.600 ;
        RECT 594.000 254.700 595.800 261.600 ;
        RECT 602.400 254.700 604.200 261.600 ;
        RECT 616.800 254.700 618.600 258.600 ;
        RECT 622.800 254.700 624.600 258.600 ;
        RECT 626.700 254.700 628.500 261.600 ;
        RECT 649.500 254.700 651.300 261.600 ;
        RECT 656.400 254.700 658.200 259.800 ;
        RECT 668.400 254.700 670.200 258.600 ;
        RECT 680.700 254.700 682.500 258.600 ;
        RECT 688.200 254.700 690.000 261.600 ;
        RECT 697.800 254.700 699.600 258.600 ;
        RECT 704.400 254.700 706.200 259.800 ;
        RECT 719.400 254.700 721.200 259.800 ;
        RECT 742.500 254.700 744.300 264.600 ;
        RECT 746.700 254.700 748.500 264.600 ;
        RECT 771.300 254.700 780.300 324.300 ;
        RECT 0.600 252.300 780.300 254.700 ;
        RECT 10.800 248.400 12.600 252.300 ;
        RECT 17.400 251.400 18.600 252.300 ;
        RECT 16.800 248.400 18.600 251.400 ;
        RECT 28.500 245.400 30.300 252.300 ;
        RECT 37.800 248.400 39.600 252.300 ;
        RECT 44.400 251.400 45.600 252.300 ;
        RECT 43.800 248.400 45.600 251.400 ;
        RECT 58.800 247.200 60.600 252.300 ;
        RECT 70.800 248.400 72.600 252.300 ;
        RECT 74.700 242.400 76.500 252.300 ;
        RECT 97.500 245.400 99.300 252.300 ;
        RECT 109.500 245.400 111.300 252.300 ;
        RECT 113.400 248.400 115.200 252.300 ;
        RECT 119.400 248.400 121.200 252.300 ;
        RECT 128.400 246.900 130.200 252.300 ;
        RECT 143.400 248.400 145.200 252.300 ;
        RECT 149.400 248.400 151.200 252.300 ;
        RECT 163.800 248.400 165.600 252.300 ;
        RECT 172.800 248.400 174.600 252.300 ;
        RECT 178.800 248.400 180.600 252.300 ;
        RECT 184.800 248.400 186.600 252.300 ;
        RECT 188.700 245.400 190.500 252.300 ;
        RECT 205.800 245.400 207.600 252.300 ;
        RECT 214.200 245.400 216.000 252.300 ;
        RECT 225.900 245.400 227.700 252.300 ;
        RECT 236.700 245.400 238.500 252.300 ;
        RECT 256.800 247.200 258.600 252.300 ;
        RECT 274.800 247.200 276.600 252.300 ;
        RECT 288.300 245.400 290.100 252.300 ;
        RECT 300.000 245.400 301.800 252.300 ;
        RECT 308.400 245.400 310.200 252.300 ;
        RECT 322.500 245.400 324.300 252.300 ;
        RECT 333.900 245.400 335.700 252.300 ;
        RECT 349.500 245.400 351.300 252.300 ;
        RECT 361.800 245.400 363.600 252.300 ;
        RECT 369.900 245.400 371.700 252.300 ;
        RECT 387.900 245.400 389.700 252.300 ;
        RECT 398.700 245.400 400.500 252.300 ;
        RECT 418.800 247.200 420.600 252.300 ;
        RECT 425.700 245.400 427.500 252.300 ;
        RECT 445.800 247.200 447.600 252.300 ;
        RECT 466.500 242.400 468.300 252.300 ;
        RECT 470.700 245.400 472.500 252.300 ;
        RECT 490.800 247.200 492.600 252.300 ;
        RECT 505.500 245.400 507.300 252.300 ;
        RECT 509.400 248.400 511.200 252.300 ;
        RECT 519.000 245.400 520.800 252.300 ;
        RECT 527.400 245.400 529.200 252.300 ;
        RECT 542.400 247.200 544.200 252.300 ;
        RECT 554.700 242.400 556.500 252.300 ;
        RECT 580.500 245.400 582.300 252.300 ;
        RECT 586.800 248.400 588.600 252.300 ;
        RECT 592.800 248.400 594.600 252.300 ;
        RECT 607.500 245.400 609.300 252.300 ;
        RECT 611.400 251.400 612.600 252.300 ;
        RECT 611.400 248.400 613.200 251.400 ;
        RECT 617.400 248.400 619.200 252.300 ;
        RECT 632.700 248.400 634.500 252.300 ;
        RECT 640.200 245.400 642.000 252.300 ;
        RECT 652.500 245.400 654.300 252.300 ;
        RECT 660.900 245.400 662.700 252.300 ;
        RECT 672.000 245.400 673.800 252.300 ;
        RECT 680.400 245.400 682.200 252.300 ;
        RECT 697.800 247.200 699.600 252.300 ;
        RECT 707.400 247.200 709.200 252.300 ;
        RECT 719.700 242.400 721.500 252.300 ;
        RECT 737.700 242.400 739.500 252.300 ;
        RECT 766.500 242.400 768.300 252.300 ;
        RECT 10.800 182.700 12.600 187.800 ;
        RECT 22.800 182.700 24.600 186.600 ;
        RECT 29.400 182.700 31.200 187.800 ;
        RECT 41.700 182.700 43.500 192.600 ;
        RECT 64.800 182.700 66.600 186.600 ;
        RECT 71.700 182.700 73.500 186.600 ;
        RECT 79.200 182.700 81.000 189.600 ;
        RECT 83.700 182.700 85.500 189.600 ;
        RECT 106.800 182.700 108.600 187.800 ;
        RECT 118.800 182.700 120.600 186.600 ;
        RECT 124.800 182.700 126.600 186.600 ;
        RECT 133.800 182.700 135.600 186.600 ;
        RECT 144.300 182.700 146.100 189.600 ;
        RECT 155.400 182.700 157.200 187.800 ;
        RECT 169.800 182.700 171.600 186.600 ;
        RECT 175.800 182.700 177.600 186.600 ;
        RECT 182.400 182.700 184.200 188.100 ;
        RECT 197.700 182.700 199.500 189.600 ;
        RECT 209.700 182.700 211.500 189.600 ;
        RECT 221.700 182.700 223.500 189.600 ;
        RECT 234.000 182.700 235.800 189.600 ;
        RECT 242.400 182.700 244.200 189.600 ;
        RECT 254.700 182.700 256.500 186.600 ;
        RECT 262.200 182.700 264.000 189.600 ;
        RECT 277.500 182.700 279.300 192.600 ;
        RECT 281.700 182.700 283.500 189.600 ;
        RECT 296.700 182.700 298.500 189.600 ;
        RECT 312.900 182.700 314.700 189.600 ;
        RECT 331.500 182.700 333.300 189.600 ;
        RECT 346.800 182.700 348.600 187.800 ;
        RECT 353.700 182.700 355.500 192.600 ;
        RECT 376.800 182.700 378.600 187.800 ;
        RECT 385.800 182.700 387.600 186.600 ;
        RECT 391.800 182.700 393.600 186.600 ;
        RECT 398.700 182.700 400.500 186.600 ;
        RECT 406.200 182.700 408.000 189.600 ;
        RECT 412.800 182.700 414.600 186.600 ;
        RECT 418.800 182.700 420.600 186.600 ;
        RECT 430.500 182.700 432.300 189.600 ;
        RECT 443.400 182.700 445.200 187.800 ;
        RECT 463.500 182.700 465.300 189.600 ;
        RECT 467.700 182.700 469.500 192.600 ;
        RECT 485.400 182.700 487.200 187.800 ;
        RECT 500.400 182.700 502.200 187.800 ;
        RECT 515.400 182.700 517.200 186.600 ;
        RECT 524.400 182.700 526.200 186.600 ;
        RECT 533.700 182.700 535.500 192.600 ;
        RECT 556.500 182.700 558.300 189.600 ;
        RECT 564.900 182.700 566.700 189.600 ;
        RECT 576.000 182.700 577.800 189.600 ;
        RECT 584.400 182.700 586.200 189.600 ;
        RECT 600.900 182.700 602.700 189.600 ;
        RECT 614.400 182.700 616.200 187.800 ;
        RECT 626.400 182.700 628.200 186.600 ;
        RECT 635.700 182.700 637.500 189.600 ;
        RECT 647.700 182.700 649.500 192.600 ;
        RECT 666.000 182.700 667.800 189.600 ;
        RECT 673.500 182.700 675.300 186.600 ;
        RECT 680.700 182.700 682.500 192.600 ;
        RECT 696.000 182.700 697.800 189.600 ;
        RECT 703.500 182.700 705.300 186.600 ;
        RECT 713.400 182.700 715.200 187.800 ;
        RECT 725.700 182.700 727.500 192.600 ;
        RECT 740.700 182.700 742.500 192.600 ;
        RECT 763.800 182.700 765.600 187.800 ;
        RECT 771.300 182.700 780.300 252.300 ;
        RECT 0.600 180.300 780.300 182.700 ;
        RECT 7.800 176.400 9.600 180.300 ;
        RECT 13.800 176.400 15.600 180.300 ;
        RECT 17.400 179.400 18.600 180.300 ;
        RECT 17.400 176.400 19.200 179.400 ;
        RECT 23.400 176.400 25.200 180.300 ;
        RECT 46.500 170.400 48.300 180.300 ;
        RECT 50.400 176.400 52.200 180.300 ;
        RECT 62.400 175.200 64.200 180.300 ;
        RECT 79.800 176.400 81.600 180.300 ;
        RECT 86.400 179.400 87.600 180.300 ;
        RECT 85.800 176.400 87.600 179.400 ;
        RECT 89.700 173.400 91.500 180.300 ;
        RECT 115.500 170.400 117.300 180.300 ;
        RECT 127.800 176.400 129.600 180.300 ;
        RECT 136.800 176.400 138.600 180.300 ;
        RECT 148.500 173.400 150.300 180.300 ;
        RECT 160.800 176.400 162.600 180.300 ;
        RECT 167.400 175.200 169.200 180.300 ;
        RECT 187.800 175.200 189.600 180.300 ;
        RECT 197.400 176.400 199.200 180.300 ;
        RECT 206.400 176.400 208.200 180.300 ;
        RECT 216.000 173.400 217.800 180.300 ;
        RECT 223.500 176.400 225.300 180.300 ;
        RECT 233.700 170.400 235.500 180.300 ;
        RECT 259.500 170.400 261.300 180.300 ;
        RECT 263.400 176.400 265.200 180.300 ;
        RECT 269.400 176.400 271.200 180.300 ;
        RECT 280.800 176.400 282.600 180.300 ;
        RECT 295.800 175.200 297.600 180.300 ;
        RECT 302.400 176.400 304.200 180.300 ;
        RECT 316.800 176.400 318.600 180.300 ;
        RECT 320.700 170.400 322.500 180.300 ;
        RECT 343.500 173.400 345.300 180.300 ;
        RECT 347.400 176.400 349.200 180.300 ;
        RECT 367.800 175.200 369.600 180.300 ;
        RECT 379.800 173.400 381.600 180.300 ;
        RECT 388.200 173.400 390.000 180.300 ;
        RECT 396.900 173.400 398.700 180.300 ;
        RECT 415.800 176.400 417.600 180.300 ;
        RECT 425.400 175.200 427.200 180.300 ;
        RECT 445.500 173.400 447.300 180.300 ;
        RECT 452.400 176.400 454.200 180.300 ;
        RECT 458.400 176.400 460.200 180.300 ;
        RECT 464.700 173.400 466.500 180.300 ;
        RECT 481.800 173.400 483.600 180.300 ;
        RECT 490.200 173.400 492.000 180.300 ;
        RECT 494.700 170.400 496.500 180.300 ;
        RECT 512.400 176.400 514.200 180.300 ;
        RECT 524.700 173.400 526.500 180.300 ;
        RECT 544.500 173.400 546.300 180.300 ;
        RECT 559.500 170.400 561.300 180.300 ;
        RECT 574.800 175.200 576.600 180.300 ;
        RECT 592.500 170.400 594.300 180.300 ;
        RECT 597.000 173.400 598.800 180.300 ;
        RECT 604.500 176.400 606.300 180.300 ;
        RECT 614.400 175.200 616.200 180.300 ;
        RECT 631.800 176.400 633.600 180.300 ;
        RECT 646.800 175.200 648.600 180.300 ;
        RECT 661.800 175.200 663.600 180.300 ;
        RECT 671.700 170.400 673.500 180.300 ;
        RECT 690.000 173.400 691.800 180.300 ;
        RECT 697.500 176.400 699.300 180.300 ;
        RECT 707.400 175.200 709.200 180.300 ;
        RECT 725.700 176.400 727.500 180.300 ;
        RECT 733.200 173.400 735.000 180.300 ;
        RECT 751.500 170.400 753.300 180.300 ;
        RECT 7.800 110.700 9.600 114.600 ;
        RECT 16.800 110.700 18.600 114.600 ;
        RECT 31.500 110.700 33.300 120.600 ;
        RECT 39.000 110.700 40.800 117.600 ;
        RECT 46.500 110.700 48.300 114.600 ;
        RECT 61.500 110.700 63.300 117.600 ;
        RECT 73.800 110.700 75.600 115.800 ;
        RECT 80.400 110.700 82.200 114.600 ;
        RECT 86.400 110.700 88.200 114.600 ;
        RECT 103.500 110.700 105.300 120.600 ;
        RECT 115.500 110.700 117.300 117.600 ;
        RECT 127.500 110.700 129.300 117.600 ;
        RECT 136.800 110.700 138.600 117.600 ;
        RECT 148.500 110.700 150.300 117.600 ;
        RECT 163.500 110.700 165.300 117.600 ;
        RECT 178.500 110.700 180.300 117.600 ;
        RECT 190.800 110.700 192.600 115.800 ;
        RECT 207.300 110.700 209.100 117.600 ;
        RECT 223.500 110.700 225.300 117.600 ;
        RECT 232.800 110.700 234.600 114.600 ;
        RECT 247.800 110.700 249.600 116.100 ;
        RECT 262.500 110.700 264.300 117.600 ;
        RECT 270.000 110.700 271.800 117.600 ;
        RECT 277.500 110.700 279.300 114.600 ;
        RECT 292.800 110.700 294.600 115.800 ;
        RECT 299.400 110.700 301.200 114.600 ;
        RECT 305.400 110.700 307.200 114.600 ;
        RECT 319.500 110.700 321.300 117.600 ;
        RECT 323.700 110.700 325.500 117.600 ;
        RECT 340.800 110.700 342.600 114.600 ;
        RECT 346.800 110.700 348.600 114.600 ;
        RECT 350.700 110.700 352.500 117.600 ;
        RECT 370.500 110.700 372.300 117.600 ;
        RECT 374.700 110.700 376.500 117.600 ;
        RECT 389.700 110.700 391.500 114.600 ;
        RECT 397.200 110.700 399.000 117.600 ;
        RECT 401.700 110.700 403.500 120.600 ;
        RECT 430.500 110.700 432.300 120.600 ;
        RECT 445.800 110.700 447.600 115.800 ;
        RECT 455.700 110.700 457.500 114.600 ;
        RECT 463.200 110.700 465.000 117.600 ;
        RECT 473.700 110.700 475.500 114.600 ;
        RECT 481.200 110.700 483.000 117.600 ;
        RECT 493.500 110.700 495.300 117.600 ;
        RECT 497.400 110.700 499.200 114.600 ;
        RECT 514.800 110.700 516.600 115.800 ;
        RECT 529.800 110.700 531.600 115.800 ;
        RECT 539.400 110.700 541.200 115.800 ;
        RECT 551.700 110.700 553.500 120.600 ;
        RECT 569.700 110.700 571.500 120.600 ;
        RECT 589.800 110.700 591.600 117.600 ;
        RECT 598.200 110.700 600.000 117.600 ;
        RECT 602.700 110.700 604.500 120.600 ;
        RECT 617.700 110.700 619.500 120.600 ;
        RECT 633.000 110.700 634.800 117.600 ;
        RECT 640.500 110.700 642.300 114.600 ;
        RECT 653.700 110.700 655.500 114.600 ;
        RECT 661.200 110.700 663.000 117.600 ;
        RECT 665.700 110.700 667.500 120.600 ;
        RECT 691.500 110.700 693.300 120.600 ;
        RECT 698.400 110.700 700.200 115.800 ;
        RECT 713.700 110.700 715.500 114.600 ;
        RECT 721.200 110.700 723.000 117.600 ;
        RECT 725.700 110.700 727.500 120.600 ;
        RECT 746.700 110.700 748.500 114.600 ;
        RECT 754.200 110.700 756.000 117.600 ;
        RECT 771.300 110.700 780.300 180.300 ;
        RECT 0.600 108.300 780.300 110.700 ;
        RECT 16.500 98.400 18.300 108.300 ;
        RECT 23.400 103.200 25.200 108.300 ;
        RECT 35.700 98.400 37.500 108.300 ;
        RECT 53.400 103.200 55.200 108.300 ;
        RECT 68.400 104.400 70.200 108.300 ;
        RECT 77.700 98.400 79.500 108.300 ;
        RECT 103.800 103.200 105.600 108.300 ;
        RECT 110.400 104.400 112.200 108.300 ;
        RECT 125.700 104.400 127.500 108.300 ;
        RECT 133.200 101.400 135.000 108.300 ;
        RECT 142.800 104.400 144.600 108.300 ;
        RECT 149.400 107.400 150.600 108.300 ;
        RECT 148.800 104.400 150.600 107.400 ;
        RECT 155.700 104.400 157.500 108.300 ;
        RECT 163.200 101.400 165.000 108.300 ;
        RECT 181.500 98.400 183.300 108.300 ;
        RECT 191.400 103.200 193.200 108.300 ;
        RECT 203.400 104.400 205.200 108.300 ;
        RECT 212.700 101.400 214.500 108.300 ;
        RECT 224.700 98.400 226.500 108.300 ;
        RECT 241.800 104.400 243.600 108.300 ;
        RECT 247.800 104.400 249.600 108.300 ;
        RECT 256.800 104.400 258.600 108.300 ;
        RECT 263.400 107.400 264.600 108.300 ;
        RECT 262.800 104.400 264.600 107.400 ;
        RECT 277.500 98.400 279.300 108.300 ;
        RECT 287.700 104.400 289.500 108.300 ;
        RECT 295.200 101.400 297.000 108.300 ;
        RECT 299.700 98.400 301.500 108.300 ;
        RECT 322.800 103.200 324.600 108.300 ;
        RECT 332.700 104.400 334.500 108.300 ;
        RECT 340.200 101.400 342.000 108.300 ;
        RECT 354.300 101.400 356.100 108.300 ;
        RECT 363.000 101.400 364.800 108.300 ;
        RECT 371.400 101.400 373.200 108.300 ;
        RECT 380.700 98.400 382.500 108.300 ;
        RECT 406.500 98.400 408.300 108.300 ;
        RECT 411.000 101.400 412.800 108.300 ;
        RECT 418.500 104.400 420.300 108.300 ;
        RECT 430.800 101.400 432.600 108.300 ;
        RECT 439.200 101.400 441.000 108.300 ;
        RECT 446.700 98.400 448.500 108.300 ;
        RECT 464.700 104.400 466.500 108.300 ;
        RECT 472.200 101.400 474.000 108.300 ;
        RECT 481.800 104.400 483.600 108.300 ;
        RECT 496.500 98.400 498.300 108.300 ;
        RECT 511.800 103.200 513.600 108.300 ;
        RECT 529.500 98.400 531.300 108.300 ;
        RECT 536.700 104.400 538.500 108.300 ;
        RECT 544.200 101.400 546.000 108.300 ;
        RECT 551.700 104.400 553.500 108.300 ;
        RECT 559.200 101.400 561.000 108.300 ;
        RECT 563.700 98.400 565.500 108.300 ;
        RECT 578.400 104.400 580.200 108.300 ;
        RECT 590.400 104.400 592.200 108.300 ;
        RECT 610.500 101.400 612.300 108.300 ;
        RECT 618.900 101.400 620.700 108.300 ;
        RECT 632.700 104.400 634.500 108.300 ;
        RECT 640.200 101.400 642.000 108.300 ;
        RECT 652.800 103.200 654.600 108.300 ;
        RECT 665.400 103.200 667.200 108.300 ;
        RECT 680.400 103.200 682.200 108.300 ;
        RECT 692.700 98.400 694.500 108.300 ;
        RECT 710.700 98.400 712.500 108.300 ;
        RECT 728.700 104.400 730.500 108.300 ;
        RECT 736.200 101.400 738.000 108.300 ;
        RECT 740.700 98.400 742.500 108.300 ;
        RECT 10.500 38.700 12.300 45.600 ;
        RECT 25.500 38.700 27.300 48.600 ;
        RECT 32.400 38.700 34.200 43.800 ;
        RECT 52.500 38.700 54.300 45.600 ;
        RECT 64.800 38.700 66.600 42.600 ;
        RECT 68.700 38.700 70.500 48.600 ;
        RECT 91.800 38.700 93.600 42.600 ;
        RECT 97.800 39.600 99.600 42.600 ;
        RECT 98.400 38.700 99.600 39.600 ;
        RECT 102.000 38.700 103.800 45.600 ;
        RECT 109.500 38.700 111.300 42.600 ;
        RECT 119.400 38.700 121.200 43.800 ;
        RECT 139.500 38.700 141.300 45.600 ;
        RECT 143.700 38.700 145.500 48.600 ;
        RECT 172.500 38.700 174.300 48.600 ;
        RECT 187.500 38.700 189.300 48.600 ;
        RECT 191.400 38.700 193.200 42.600 ;
        RECT 200.700 38.700 202.500 45.600 ;
        RECT 212.700 38.700 214.500 48.600 ;
        RECT 227.700 38.700 229.500 45.600 ;
        RECT 243.900 38.700 245.700 45.600 ;
        RECT 265.500 38.700 267.300 45.600 ;
        RECT 272.400 38.700 274.200 42.600 ;
        RECT 278.400 38.700 280.200 42.600 ;
        RECT 295.500 38.700 297.300 48.600 ;
        RECT 307.800 38.700 309.600 43.800 ;
        RECT 318.000 38.700 319.800 45.600 ;
        RECT 325.500 38.700 327.300 42.600 ;
        RECT 343.500 38.700 345.300 48.600 ;
        RECT 350.700 38.700 352.500 48.600 ;
        RECT 370.800 38.700 372.600 42.600 ;
        RECT 374.700 38.700 376.500 48.600 ;
        RECT 389.700 38.700 391.500 48.600 ;
        RECT 410.400 38.700 412.200 43.800 ;
        RECT 423.000 38.700 424.800 45.600 ;
        RECT 430.500 38.700 432.300 42.600 ;
        RECT 440.400 38.700 442.200 43.800 ;
        RECT 452.700 38.700 454.500 48.600 ;
        RECT 478.500 38.700 480.300 48.600 ;
        RECT 485.700 38.700 487.500 48.600 ;
        RECT 501.000 38.700 502.800 45.600 ;
        RECT 508.500 38.700 510.300 42.600 ;
        RECT 515.700 38.700 517.500 48.600 ;
        RECT 533.400 38.700 535.200 43.800 ;
        RECT 545.700 38.700 547.500 48.600 ;
        RECT 563.400 38.700 565.200 43.800 ;
        RECT 578.700 38.700 580.500 45.600 ;
        RECT 590.400 38.700 592.200 42.600 ;
        RECT 596.400 38.700 598.200 42.600 ;
        RECT 607.800 38.700 609.600 42.600 ;
        RECT 613.800 38.700 615.600 42.600 ;
        RECT 625.800 38.700 627.600 43.800 ;
        RECT 635.700 38.700 637.500 45.600 ;
        RECT 647.400 38.700 649.200 42.600 ;
        RECT 659.400 38.700 661.200 43.800 ;
        RECT 674.700 38.700 676.500 42.600 ;
        RECT 682.200 38.700 684.000 45.600 ;
        RECT 689.700 38.700 691.500 42.600 ;
        RECT 697.200 38.700 699.000 45.600 ;
        RECT 701.700 38.700 703.500 48.600 ;
        RECT 730.500 38.700 732.300 48.600 ;
        RECT 734.700 38.700 736.500 48.600 ;
        RECT 750.000 38.700 751.800 45.600 ;
        RECT 757.500 38.700 759.300 42.600 ;
        RECT 771.300 38.700 780.300 108.300 ;
        RECT 0.600 36.300 780.300 38.700 ;
        RECT 4.800 32.400 6.600 36.300 ;
        RECT 10.800 32.400 12.600 36.300 ;
        RECT 18.900 29.400 20.700 36.300 ;
        RECT 35.400 31.200 37.200 36.300 ;
        RECT 54.300 29.400 56.100 36.300 ;
        RECT 70.500 29.400 72.300 36.300 ;
        RECT 75.000 29.400 76.800 36.300 ;
        RECT 83.400 29.400 85.200 36.300 ;
        RECT 92.700 26.400 94.500 36.300 ;
        RECT 110.700 32.400 112.500 36.300 ;
        RECT 118.200 29.400 120.000 36.300 ;
        RECT 122.700 26.400 124.500 36.300 ;
        RECT 145.800 31.200 147.600 36.300 ;
        RECT 155.400 31.200 157.200 36.300 ;
        RECT 173.400 31.200 175.200 36.300 ;
        RECT 185.700 26.400 187.500 36.300 ;
        RECT 200.700 26.400 202.500 36.300 ;
        RECT 226.800 31.200 228.600 36.300 ;
        RECT 236.700 32.400 238.500 36.300 ;
        RECT 244.200 29.400 246.000 36.300 ;
        RECT 248.700 26.400 250.500 36.300 ;
        RECT 264.000 29.400 265.800 36.300 ;
        RECT 271.500 32.400 273.300 36.300 ;
        RECT 281.400 31.200 283.200 36.300 ;
        RECT 293.700 26.400 295.500 36.300 ;
        RECT 314.700 32.400 316.500 36.300 ;
        RECT 322.200 29.400 324.000 36.300 ;
        RECT 329.700 26.400 331.500 36.300 ;
        RECT 352.800 31.200 354.600 36.300 ;
        RECT 362.400 31.200 364.200 36.300 ;
        RECT 377.100 32.400 379.200 36.300 ;
        RECT 383.400 32.400 385.200 36.300 ;
        RECT 407.400 31.200 409.200 36.300 ;
        RECT 425.700 32.400 427.500 36.300 ;
        RECT 433.200 29.400 435.000 36.300 ;
        RECT 444.300 29.400 446.100 36.300 ;
        RECT 460.800 29.400 462.600 36.300 ;
        RECT 469.200 29.400 471.000 36.300 ;
        RECT 473.700 29.400 475.500 36.300 ;
        RECT 493.800 31.200 495.600 36.300 ;
        RECT 507.300 29.400 509.100 36.300 ;
        RECT 520.800 32.400 522.600 36.300 ;
        RECT 526.800 32.400 528.600 36.300 ;
        RECT 533.400 31.200 535.200 36.300 ;
        RECT 548.400 32.400 550.200 36.300 ;
        RECT 557.700 26.400 559.500 36.300 ;
        RECT 577.800 32.400 579.600 36.300 ;
        RECT 584.400 35.400 585.600 36.300 ;
        RECT 583.800 32.400 585.600 35.400 ;
        RECT 595.500 29.400 597.300 36.300 ;
        RECT 607.500 29.400 609.300 36.300 ;
        RECT 622.500 26.400 624.300 36.300 ;
        RECT 626.700 26.400 628.500 36.300 ;
        RECT 641.700 29.400 643.500 36.300 ;
        RECT 664.500 26.400 666.300 36.300 ;
        RECT 671.400 32.400 673.200 36.300 ;
        RECT 683.700 26.400 685.500 36.300 ;
        RECT 698.700 29.400 700.500 36.300 ;
        RECT 713.400 31.200 715.200 36.300 ;
        RECT 733.800 31.200 735.600 36.300 ;
        RECT 743.400 31.200 745.200 36.300 ;
        RECT 771.300 0.300 780.300 36.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.300 720.300 770.400 722.700 ;
        RECT -9.300 650.700 -0.300 720.300 ;
        RECT 4.800 707.400 6.600 720.300 ;
        RECT 13.800 712.200 15.600 720.300 ;
        RECT 26.400 713.400 28.200 720.300 ;
        RECT 33.900 707.400 35.700 720.300 ;
        RECT 43.800 713.400 45.600 720.300 ;
        RECT 51.300 707.400 53.100 720.300 ;
        RECT 58.800 713.400 60.600 720.300 ;
        RECT 68.400 713.400 70.200 720.300 ;
        RECT 75.900 707.400 77.700 720.300 ;
        RECT 88.800 709.200 90.600 720.300 ;
        RECT 98.400 713.400 100.200 720.300 ;
        RECT 105.900 707.400 107.700 720.300 ;
        RECT 110.400 713.400 112.200 720.300 ;
        RECT 125.400 712.200 127.200 720.300 ;
        RECT 134.400 707.400 136.200 720.300 ;
        RECT 143.400 713.400 145.200 720.300 ;
        RECT 150.900 707.400 152.700 720.300 ;
        RECT 158.700 707.400 160.500 720.300 ;
        RECT 175.800 709.200 177.600 720.300 ;
        RECT 186.300 707.400 188.100 720.300 ;
        RECT 193.800 713.400 195.600 720.300 ;
        RECT 202.800 713.400 204.600 720.300 ;
        RECT 208.800 713.400 210.600 720.300 ;
        RECT 219.300 707.550 221.100 720.300 ;
        RECT 232.800 713.400 234.600 720.300 ;
        RECT 242.400 713.400 244.200 720.300 ;
        RECT 249.900 707.400 251.700 720.300 ;
        RECT 254.400 707.400 256.200 720.300 ;
        RECT 271.800 713.400 273.600 720.300 ;
        RECT 276.300 707.400 278.100 720.300 ;
        RECT 283.800 713.400 285.600 720.300 ;
        RECT 290.400 707.400 292.200 720.300 ;
        RECT 310.800 709.200 312.600 720.300 ;
        RECT 318.300 707.400 320.100 720.300 ;
        RECT 325.800 713.400 327.600 720.300 ;
        RECT 337.800 707.400 339.600 720.300 ;
        RECT 343.800 707.400 345.600 720.300 ;
        RECT 347.400 713.400 349.200 720.300 ;
        RECT 353.400 713.400 355.200 720.300 ;
        RECT 370.800 709.500 372.600 720.300 ;
        RECT 381.300 707.400 383.100 720.300 ;
        RECT 388.800 713.400 390.600 720.300 ;
        RECT 395.400 713.400 397.200 720.300 ;
        RECT 401.400 713.400 403.200 720.300 ;
        RECT 410.400 713.400 412.200 720.300 ;
        RECT 427.800 707.400 429.600 720.300 ;
        RECT 434.700 707.400 436.500 720.300 ;
        RECT 447.150 713.400 448.950 720.300 ;
        RECT 457.350 713.400 459.150 720.300 ;
        RECT 463.950 713.400 465.750 720.300 ;
        RECT 472.650 716.400 474.450 720.300 ;
        RECT 484.800 707.400 486.600 720.300 ;
        RECT 490.800 707.400 492.600 720.300 ;
        RECT 496.800 707.400 498.600 720.300 ;
        RECT 502.800 707.400 504.600 720.300 ;
        RECT 508.800 707.400 510.600 720.300 ;
        RECT 513.300 707.400 515.100 720.300 ;
        RECT 520.800 713.400 522.600 720.300 ;
        RECT 532.800 713.400 534.600 720.300 ;
        RECT 538.800 713.400 540.600 720.300 ;
        RECT 545.550 716.400 547.350 720.300 ;
        RECT 554.250 713.400 556.050 720.300 ;
        RECT 560.850 713.400 562.650 720.300 ;
        RECT 571.050 713.400 572.850 720.300 ;
        RECT 578.400 707.400 580.200 720.300 ;
        RECT 584.400 707.400 586.200 720.300 ;
        RECT 590.400 707.400 592.200 720.300 ;
        RECT 596.400 707.400 598.200 720.300 ;
        RECT 602.400 707.400 604.200 720.300 ;
        RECT 610.200 713.400 612.000 720.300 ;
        RECT 616.800 713.400 618.600 720.300 ;
        RECT 622.800 713.400 624.600 720.300 ;
        RECT 628.800 713.400 630.600 720.300 ;
        RECT 645.000 713.400 646.800 720.300 ;
        RECT 651.900 713.400 653.700 720.300 ;
        RECT 664.500 718.050 666.300 720.300 ;
        RECT 664.500 715.950 666.600 718.050 ;
        RECT 670.500 713.400 672.300 720.300 ;
        RECT 676.500 713.400 678.300 720.300 ;
        RECT 688.800 709.200 690.600 720.300 ;
        RECT 697.200 713.400 699.000 720.300 ;
        RECT 703.800 713.400 705.600 720.300 ;
        RECT 709.800 713.400 711.600 720.300 ;
        RECT 715.800 713.400 717.600 720.300 ;
        RECT 732.000 713.400 733.800 720.300 ;
        RECT 738.900 713.400 740.700 720.300 ;
        RECT 751.500 718.050 753.300 720.300 ;
        RECT 751.500 715.950 753.600 718.050 ;
        RECT 757.500 713.400 759.300 720.300 ;
        RECT 763.500 713.400 765.300 720.300 ;
        RECT 4.800 650.700 6.600 657.600 ;
        RECT 10.800 650.700 12.600 657.600 ;
        RECT 20.400 650.700 22.200 657.600 ;
        RECT 27.900 650.700 29.700 663.600 ;
        RECT 32.400 650.700 34.200 657.600 ;
        RECT 38.400 650.700 40.200 657.600 ;
        RECT 49.800 650.700 51.600 657.000 ;
        RECT 55.800 650.700 57.600 657.600 ;
        RECT 61.800 650.700 63.600 657.600 ;
        RECT 67.800 650.700 69.600 657.600 ;
        RECT 76.800 650.700 78.600 657.600 ;
        RECT 82.800 650.700 84.600 657.600 ;
        RECT 89.400 650.700 91.200 657.600 ;
        RECT 96.900 650.700 98.700 663.600 ;
        RECT 101.400 650.700 103.200 663.600 ;
        RECT 116.400 650.700 118.200 657.600 ;
        RECT 123.900 650.700 125.700 663.600 ;
        RECT 128.400 650.700 130.200 657.600 ;
        RECT 134.400 650.700 136.200 657.600 ;
        RECT 146.400 650.700 148.200 657.600 ;
        RECT 153.900 650.700 155.700 663.600 ;
        RECT 166.800 650.700 168.600 663.600 ;
        RECT 176.400 650.700 178.200 657.600 ;
        RECT 183.900 650.700 185.700 663.600 ;
        RECT 191.400 650.700 193.200 657.600 ;
        RECT 198.900 650.700 200.700 663.600 ;
        RECT 208.800 650.700 210.600 657.600 ;
        RECT 215.400 650.700 217.200 657.600 ;
        RECT 222.900 650.700 224.700 663.600 ;
        RECT 230.400 650.700 232.200 661.500 ;
        RECT 253.800 650.700 255.600 657.000 ;
        RECT 259.800 650.700 261.600 657.600 ;
        RECT 265.800 650.700 267.600 657.600 ;
        RECT 271.800 650.700 273.600 657.600 ;
        RECT 281.400 650.700 283.200 657.600 ;
        RECT 288.900 650.700 290.700 663.600 ;
        RECT 293.400 650.700 295.200 657.600 ;
        RECT 299.400 650.700 301.200 657.600 ;
        RECT 310.800 650.700 312.600 657.000 ;
        RECT 316.800 650.700 318.600 657.600 ;
        RECT 322.800 650.700 324.600 657.600 ;
        RECT 328.800 650.700 330.600 657.600 ;
        RECT 343.800 650.700 345.600 661.500 ;
        RECT 353.400 650.700 355.200 657.600 ;
        RECT 360.900 650.700 362.700 663.600 ;
        RECT 365.400 650.700 367.200 657.600 ;
        RECT 371.400 650.700 373.200 657.600 ;
        RECT 380.400 650.700 382.200 663.600 ;
        RECT 392.400 650.700 394.200 657.600 ;
        RECT 404.400 650.700 406.200 657.600 ;
        RECT 410.400 650.700 412.200 657.600 ;
        RECT 416.400 650.700 418.200 657.600 ;
        RECT 427.800 650.700 429.600 657.600 ;
        RECT 433.800 650.700 435.600 657.600 ;
        RECT 437.400 650.700 439.200 657.600 ;
        RECT 452.400 650.700 454.200 657.600 ;
        RECT 459.900 650.700 461.700 663.600 ;
        RECT 467.550 650.700 469.350 654.600 ;
        RECT 476.250 650.700 478.050 657.600 ;
        RECT 482.850 650.700 484.650 657.600 ;
        RECT 493.050 650.700 494.850 657.600 ;
        RECT 501.300 650.700 503.100 663.600 ;
        RECT 508.800 650.700 510.600 657.600 ;
        RECT 515.400 650.700 517.200 657.600 ;
        RECT 521.400 650.700 523.200 657.600 ;
        RECT 527.400 650.700 529.200 657.600 ;
        RECT 537.300 650.700 539.100 663.600 ;
        RECT 544.800 650.700 546.600 657.600 ;
        RECT 553.800 650.700 555.600 657.600 ;
        RECT 559.800 650.700 561.600 657.600 ;
        RECT 567.150 650.700 568.950 657.600 ;
        RECT 577.350 650.700 579.150 657.600 ;
        RECT 583.950 650.700 585.750 657.600 ;
        RECT 592.650 650.700 594.450 654.600 ;
        RECT 601.800 650.700 603.600 657.600 ;
        RECT 607.800 650.700 609.600 657.600 ;
        RECT 613.200 650.700 615.000 657.600 ;
        RECT 619.800 650.700 621.600 657.600 ;
        RECT 625.800 650.700 627.600 657.600 ;
        RECT 631.800 650.700 633.600 657.600 ;
        RECT 648.000 650.700 649.800 657.600 ;
        RECT 654.900 650.700 656.700 657.600 ;
        RECT 667.500 650.700 669.300 655.050 ;
        RECT 673.500 650.700 675.300 657.600 ;
        RECT 679.500 650.700 681.300 657.600 ;
        RECT 686.400 650.700 688.200 657.600 ;
        RECT 692.400 650.700 694.200 657.600 ;
        RECT 701.400 650.700 703.200 657.600 ;
        RECT 708.900 650.700 710.700 663.600 ;
        RECT 724.800 650.700 726.600 663.600 ;
        RECT 733.800 650.700 735.600 657.000 ;
        RECT 739.800 650.700 741.600 657.600 ;
        RECT 746.400 650.700 748.200 657.600 ;
        RECT 755.400 650.700 757.200 657.600 ;
        RECT -9.300 648.300 770.400 650.700 ;
        RECT -9.300 578.700 -0.300 648.300 ;
        RECT 10.800 635.400 12.600 648.300 ;
        RECT 14.400 641.400 16.200 648.300 ;
        RECT 21.000 635.400 22.800 648.300 ;
        RECT 31.800 641.400 33.600 648.300 ;
        RECT 37.800 641.400 39.600 648.300 ;
        RECT 41.400 641.400 43.200 648.300 ;
        RECT 47.400 642.000 49.200 648.300 ;
        RECT 59.400 641.400 61.200 648.300 ;
        RECT 71.400 637.200 73.200 648.300 ;
        RECT 88.800 641.400 90.600 648.300 ;
        RECT 95.400 641.400 97.200 648.300 ;
        RECT 102.900 635.400 104.700 648.300 ;
        RECT 110.400 641.400 112.200 648.300 ;
        RECT 117.900 635.400 119.700 648.300 ;
        RECT 130.800 637.200 132.600 648.300 ;
        RECT 143.400 641.400 145.200 648.300 ;
        RECT 150.900 635.400 152.700 648.300 ;
        RECT 158.400 641.400 160.200 648.300 ;
        RECT 165.900 635.400 167.700 648.300 ;
        RECT 173.400 641.400 175.200 648.300 ;
        RECT 180.900 635.400 182.700 648.300 ;
        RECT 188.400 641.400 190.200 648.300 ;
        RECT 194.400 641.400 196.200 648.300 ;
        RECT 211.800 637.500 213.600 648.300 ;
        RECT 223.200 635.400 225.000 648.300 ;
        RECT 229.800 641.400 231.600 648.300 ;
        RECT 235.800 641.400 237.600 648.300 ;
        RECT 241.800 641.400 243.600 648.300 ;
        RECT 248.400 641.400 250.200 648.300 ;
        RECT 255.900 635.400 257.700 648.300 ;
        RECT 263.400 637.500 265.200 648.300 ;
        RECT 278.400 641.400 280.200 648.300 ;
        RECT 284.400 641.400 286.200 648.300 ;
        RECT 295.800 635.400 297.600 648.300 ;
        RECT 302.400 641.400 304.200 648.300 ;
        RECT 309.900 635.400 311.700 648.300 ;
        RECT 319.800 641.400 321.600 648.300 ;
        RECT 325.800 641.400 327.600 648.300 ;
        RECT 331.800 641.400 333.600 648.300 ;
        RECT 341.400 640.200 343.200 648.300 ;
        RECT 350.400 635.400 352.200 648.300 ;
        RECT 362.700 635.400 364.500 648.300 ;
        RECT 371.400 641.400 373.200 648.300 ;
        RECT 377.400 641.400 379.200 648.300 ;
        RECT 386.400 641.400 388.200 648.300 ;
        RECT 393.900 635.400 395.700 648.300 ;
        RECT 406.500 635.400 408.300 648.300 ;
        RECT 416.550 644.400 418.350 648.300 ;
        RECT 425.250 641.400 427.050 648.300 ;
        RECT 431.850 641.400 433.650 648.300 ;
        RECT 442.050 641.400 443.850 648.300 ;
        RECT 455.400 641.400 457.200 648.300 ;
        RECT 462.900 635.400 464.700 648.300 ;
        RECT 467.400 641.400 469.200 648.300 ;
        RECT 473.400 641.400 475.200 648.300 ;
        RECT 482.550 644.400 484.350 648.300 ;
        RECT 491.250 641.400 493.050 648.300 ;
        RECT 497.850 641.400 499.650 648.300 ;
        RECT 508.050 641.400 509.850 648.300 ;
        RECT 518.700 635.400 520.500 648.300 ;
        RECT 532.800 641.400 534.600 648.300 ;
        RECT 538.800 641.400 540.600 648.300 ;
        RECT 545.400 641.400 547.200 648.300 ;
        RECT 552.900 635.400 554.700 648.300 ;
        RECT 559.800 641.400 561.600 648.300 ;
        RECT 565.800 641.400 567.600 648.300 ;
        RECT 572.400 641.400 574.200 648.300 ;
        RECT 579.900 635.400 581.700 648.300 ;
        RECT 587.700 635.400 589.500 648.300 ;
        RECT 597.300 635.400 599.100 648.300 ;
        RECT 604.800 641.400 606.600 648.300 ;
        RECT 615.150 641.400 616.950 648.300 ;
        RECT 625.350 641.400 627.150 648.300 ;
        RECT 631.950 641.400 633.750 648.300 ;
        RECT 640.650 644.400 642.450 648.300 ;
        RECT 654.300 635.550 656.100 648.300 ;
        RECT 665.400 641.400 667.200 648.300 ;
        RECT 672.900 635.400 674.700 648.300 ;
        RECT 676.950 646.950 679.050 648.300 ;
        RECT 680.400 641.400 682.200 648.300 ;
        RECT 687.900 635.400 689.700 648.300 ;
        RECT 696.300 635.400 698.100 648.300 ;
        RECT 706.800 635.400 708.600 648.300 ;
        RECT 710.400 641.400 712.200 648.300 ;
        RECT 730.800 637.500 732.600 648.300 ;
        RECT 740.400 641.400 742.200 648.300 ;
        RECT 752.400 641.400 754.200 648.300 ;
        RECT 759.900 635.400 761.700 648.300 ;
        RECT 6.300 578.700 8.100 591.600 ;
        RECT 13.800 578.700 15.600 585.600 ;
        RECT 28.800 578.700 30.600 585.600 ;
        RECT 33.300 578.700 35.100 591.600 ;
        RECT 40.800 578.700 42.600 585.600 ;
        RECT 52.800 578.700 54.600 585.600 ;
        RECT 58.800 578.700 60.600 585.600 ;
        RECT 65.400 578.700 67.200 585.600 ;
        RECT 71.400 578.700 73.200 585.000 ;
        RECT 88.800 578.700 90.600 589.800 ;
        RECT 100.800 578.700 102.600 585.600 ;
        RECT 104.400 578.700 106.200 585.600 ;
        RECT 110.400 578.700 112.200 585.600 ;
        RECT 116.400 578.700 118.200 585.600 ;
        RECT 130.500 578.700 132.300 591.600 ;
        RECT 143.700 578.700 145.500 591.600 ;
        RECT 154.800 578.700 156.600 585.600 ;
        RECT 160.800 578.700 162.600 585.600 ;
        RECT 172.800 578.700 174.600 591.600 ;
        RECT 181.800 578.700 183.600 585.600 ;
        RECT 185.400 578.700 187.200 585.600 ;
        RECT 191.400 578.700 193.200 585.600 ;
        RECT 200.400 578.700 202.200 585.600 ;
        RECT 207.900 578.700 209.700 591.600 ;
        RECT 215.400 578.700 217.200 589.500 ;
        RECT 230.400 578.700 232.200 585.600 ;
        RECT 236.400 578.700 238.200 585.600 ;
        RECT 246.300 578.700 248.100 591.600 ;
        RECT 253.800 578.700 255.600 585.600 ;
        RECT 268.200 578.700 270.000 591.600 ;
        RECT 274.800 578.700 276.600 585.600 ;
        RECT 283.800 578.700 285.600 585.000 ;
        RECT 289.800 578.700 291.600 585.600 ;
        RECT 296.400 578.700 298.200 585.600 ;
        RECT 303.900 578.700 305.700 591.600 ;
        RECT 308.400 578.700 310.200 591.600 ;
        RECT 328.800 578.700 330.600 585.600 ;
        RECT 333.300 578.700 335.100 591.600 ;
        RECT 340.800 578.700 342.600 585.600 ;
        RECT 347.400 578.700 349.200 585.600 ;
        RECT 364.800 578.700 366.600 585.600 ;
        RECT 368.400 578.700 370.200 585.600 ;
        RECT 381.150 578.700 382.950 585.600 ;
        RECT 391.350 578.700 393.150 585.600 ;
        RECT 397.950 578.700 399.750 585.600 ;
        RECT 406.650 578.700 408.450 582.600 ;
        RECT 416.550 578.700 418.350 582.600 ;
        RECT 425.250 578.700 427.050 585.600 ;
        RECT 431.850 578.700 433.650 585.600 ;
        RECT 442.050 578.700 443.850 585.600 ;
        RECT 449.400 578.700 451.200 585.600 ;
        RECT 455.400 578.700 457.200 585.600 ;
        RECT 464.400 578.700 466.200 585.600 ;
        RECT 471.900 578.700 473.700 591.600 ;
        RECT 476.400 578.700 478.200 585.600 ;
        RECT 490.500 578.700 492.300 591.600 ;
        RECT 502.500 578.700 504.300 591.600 ;
        RECT 514.800 578.700 516.600 585.600 ;
        RECT 520.800 578.700 522.600 585.600 ;
        RECT 527.400 578.700 529.200 585.600 ;
        RECT 534.900 578.700 536.700 591.600 ;
        RECT 542.550 578.700 544.350 582.600 ;
        RECT 551.250 578.700 553.050 585.600 ;
        RECT 557.850 578.700 559.650 585.600 ;
        RECT 568.050 578.700 569.850 585.600 ;
        RECT 579.150 578.700 580.950 585.600 ;
        RECT 589.350 578.700 591.150 585.600 ;
        RECT 595.950 578.700 597.750 585.600 ;
        RECT 604.650 578.700 606.450 582.600 ;
        RECT 616.800 578.700 618.600 585.600 ;
        RECT 628.500 578.700 630.300 591.600 ;
        RECT 635.400 578.700 637.200 585.600 ;
        RECT 641.400 578.700 643.200 585.600 ;
        RECT 655.800 578.700 657.600 591.600 ;
        RECT 662.400 578.700 664.200 589.800 ;
        RECT 675.300 578.700 677.100 591.600 ;
        RECT 682.800 578.700 684.600 585.600 ;
        RECT 694.800 578.700 696.600 585.600 ;
        RECT 698.400 578.700 700.200 591.600 ;
        RECT 710.400 578.700 712.200 585.600 ;
        RECT 722.400 578.700 724.200 591.600 ;
        RECT 735.300 578.700 737.100 591.600 ;
        RECT 742.800 578.700 744.600 585.600 ;
        RECT 752.400 578.700 754.200 589.800 ;
        RECT -9.300 576.300 770.400 578.700 ;
        RECT -9.300 506.700 -0.300 576.300 ;
        RECT 7.500 563.400 9.300 576.300 ;
        RECT 20.400 569.400 22.200 576.300 ;
        RECT 27.900 563.400 29.700 576.300 ;
        RECT 33.300 563.400 35.100 576.300 ;
        RECT 40.800 569.400 42.600 576.300 ;
        RECT 55.800 565.200 57.600 576.300 ;
        RECT 63.300 563.400 65.100 576.300 ;
        RECT 70.800 569.400 72.600 576.300 ;
        RECT 80.400 565.200 82.200 576.300 ;
        RECT 95.400 569.400 97.200 576.300 ;
        RECT 102.900 563.400 104.700 576.300 ;
        RECT 110.400 569.400 112.200 576.300 ;
        RECT 117.900 563.400 119.700 576.300 ;
        RECT 126.300 563.400 128.100 576.300 ;
        RECT 133.800 569.400 135.600 576.300 ;
        RECT 143.400 569.400 145.200 576.300 ;
        RECT 150.900 563.400 152.700 576.300 ;
        RECT 163.800 565.200 165.600 576.300 ;
        RECT 171.300 563.400 173.100 576.300 ;
        RECT 178.800 569.400 180.600 576.300 ;
        RECT 187.800 569.400 189.600 576.300 ;
        RECT 193.800 569.400 195.600 576.300 ;
        RECT 205.800 563.400 207.600 576.300 ;
        RECT 214.800 569.400 216.600 576.300 ;
        RECT 220.800 569.400 222.600 576.300 ;
        RECT 227.400 569.400 229.200 576.300 ;
        RECT 234.900 563.400 236.700 576.300 ;
        RECT 242.400 565.500 244.200 576.300 ;
        RECT 257.400 569.400 259.200 576.300 ;
        RECT 263.400 569.400 265.200 576.300 ;
        RECT 273.300 563.400 275.100 576.300 ;
        RECT 280.800 569.400 282.600 576.300 ;
        RECT 292.200 563.400 294.000 576.300 ;
        RECT 298.800 569.400 300.600 576.300 ;
        RECT 307.800 563.400 309.600 576.300 ;
        RECT 312.300 563.400 314.100 576.300 ;
        RECT 319.800 569.400 321.600 576.300 ;
        RECT 331.500 563.400 333.300 576.300 ;
        RECT 341.550 572.400 343.350 576.300 ;
        RECT 350.250 569.400 352.050 576.300 ;
        RECT 356.850 569.400 358.650 576.300 ;
        RECT 367.050 569.400 368.850 576.300 ;
        RECT 374.400 569.400 376.200 576.300 ;
        RECT 384.300 563.400 386.100 576.300 ;
        RECT 391.800 569.400 393.600 576.300 ;
        RECT 401.400 569.400 403.200 576.300 ;
        RECT 407.400 569.400 409.200 576.300 ;
        RECT 416.400 569.400 418.200 576.300 ;
        RECT 423.900 563.400 425.700 576.300 ;
        RECT 432.300 563.400 434.100 576.300 ;
        RECT 439.800 569.400 441.600 576.300 ;
        RECT 448.800 569.400 450.600 576.300 ;
        RECT 454.800 569.400 456.600 576.300 ;
        RECT 462.150 569.400 463.950 576.300 ;
        RECT 472.350 569.400 474.150 576.300 ;
        RECT 478.950 569.400 480.750 576.300 ;
        RECT 487.650 572.400 489.450 576.300 ;
        RECT 500.700 563.400 502.500 576.300 ;
        RECT 514.500 563.400 516.300 576.300 ;
        RECT 526.500 563.400 528.300 576.300 ;
        RECT 536.550 572.400 538.350 576.300 ;
        RECT 545.250 569.400 547.050 576.300 ;
        RECT 551.850 569.400 553.650 576.300 ;
        RECT 562.050 569.400 563.850 576.300 ;
        RECT 572.700 563.400 574.500 576.300 ;
        RECT 587.400 569.400 589.200 576.300 ;
        RECT 594.900 563.400 596.700 576.300 ;
        RECT 599.400 563.400 601.200 576.300 ;
        RECT 615.300 563.400 617.100 576.300 ;
        RECT 622.800 569.400 624.600 576.300 ;
        RECT 629.400 569.400 631.200 576.300 ;
        RECT 646.800 569.400 648.600 576.300 ;
        RECT 653.400 569.400 655.200 576.300 ;
        RECT 659.400 569.400 661.200 576.300 ;
        RECT 665.400 563.400 667.200 576.300 ;
        RECT 680.400 565.500 682.200 576.300 ;
        RECT 696.300 563.400 698.100 576.300 ;
        RECT 703.800 569.400 705.600 576.300 ;
        RECT 710.400 569.400 712.200 576.300 ;
        RECT 716.400 570.000 718.200 576.300 ;
        RECT 727.800 563.400 729.600 576.300 ;
        RECT 733.800 563.400 735.600 576.300 ;
        RECT 740.400 569.400 742.200 576.300 ;
        RECT 747.000 563.400 748.800 576.300 ;
        RECT 10.500 506.700 12.300 519.600 ;
        RECT 28.800 506.700 30.600 517.800 ;
        RECT 43.800 506.700 45.600 513.600 ;
        RECT 50.400 506.700 52.200 513.600 ;
        RECT 57.900 506.700 59.700 519.600 ;
        RECT 64.800 506.700 66.600 513.600 ;
        RECT 70.800 506.700 72.600 513.600 ;
        RECT 77.400 506.700 79.200 513.600 ;
        RECT 84.900 506.700 86.700 519.600 ;
        RECT 92.400 506.700 94.200 513.600 ;
        RECT 99.900 506.700 101.700 519.600 ;
        RECT 104.400 506.700 106.200 513.600 ;
        RECT 110.400 506.700 112.200 513.600 ;
        RECT 119.400 506.700 121.200 517.800 ;
        RECT 136.800 506.700 138.600 513.600 ;
        RECT 148.800 506.700 150.600 517.800 ;
        RECT 155.400 506.700 157.200 513.600 ;
        RECT 167.400 506.700 169.200 517.800 ;
        RECT 183.300 506.700 185.100 519.600 ;
        RECT 190.800 506.700 192.600 513.600 ;
        RECT 200.400 506.700 202.200 519.600 ;
        RECT 212.400 506.700 214.200 519.600 ;
        RECT 232.800 506.700 234.600 519.600 ;
        RECT 239.400 506.700 241.200 517.500 ;
        RECT 254.400 506.700 256.200 513.600 ;
        RECT 260.400 506.700 262.200 513.600 ;
        RECT 271.200 506.700 273.000 519.600 ;
        RECT 277.800 506.700 279.600 513.600 ;
        RECT 284.400 506.700 286.200 513.600 ;
        RECT 291.900 506.700 293.700 519.600 ;
        RECT 299.400 506.700 301.200 517.500 ;
        RECT 317.400 506.700 319.200 513.600 ;
        RECT 323.400 506.700 325.200 513.600 ;
        RECT 329.400 506.700 331.200 513.600 ;
        RECT 336.000 506.700 337.800 519.600 ;
        RECT 345.300 506.700 347.100 519.600 ;
        RECT 352.800 506.700 354.600 513.600 ;
        RECT 362.400 506.700 364.200 519.600 ;
        RECT 377.400 506.700 379.200 513.600 ;
        RECT 384.900 506.700 386.700 519.600 ;
        RECT 389.400 506.700 391.200 513.600 ;
        RECT 395.400 506.700 397.200 513.600 ;
        RECT 407.400 506.700 409.200 513.600 ;
        RECT 414.900 506.700 416.700 519.600 ;
        RECT 419.400 506.700 421.200 513.600 ;
        RECT 428.400 506.700 430.200 513.600 ;
        RECT 434.400 506.700 436.200 513.600 ;
        RECT 448.800 506.700 450.600 517.800 ;
        RECT 456.300 506.700 458.100 519.600 ;
        RECT 463.800 506.700 465.600 513.600 ;
        RECT 470.400 506.700 472.200 513.600 ;
        RECT 476.400 506.700 478.200 513.600 ;
        RECT 485.550 506.700 487.350 510.600 ;
        RECT 494.250 506.700 496.050 513.600 ;
        RECT 500.850 506.700 502.650 513.600 ;
        RECT 511.050 506.700 512.850 513.600 ;
        RECT 519.300 506.700 521.100 519.600 ;
        RECT 526.800 506.700 528.600 513.600 ;
        RECT 533.400 506.700 535.200 513.600 ;
        RECT 539.400 506.700 541.200 513.600 ;
        RECT 548.700 506.700 550.500 519.600 ;
        RECT 558.300 506.700 560.100 519.600 ;
        RECT 565.800 506.700 567.600 513.600 ;
        RECT 575.550 506.700 577.350 510.600 ;
        RECT 584.250 506.700 586.050 513.600 ;
        RECT 590.850 506.700 592.650 513.600 ;
        RECT 601.050 506.700 602.850 513.600 ;
        RECT 612.300 506.700 614.100 519.600 ;
        RECT 619.800 506.700 621.600 513.600 ;
        RECT 626.400 506.700 628.200 513.600 ;
        RECT 632.400 506.700 634.200 513.600 ;
        RECT 641.700 506.700 643.500 519.600 ;
        RECT 653.400 506.700 655.200 513.600 ;
        RECT 659.400 506.700 661.200 513.600 ;
        RECT 665.400 506.700 667.200 513.600 ;
        RECT 671.400 506.700 673.200 513.600 ;
        RECT 679.800 506.700 681.600 519.600 ;
        RECT 685.800 506.700 687.600 519.600 ;
        RECT 691.800 506.700 693.600 519.600 ;
        RECT 697.800 506.700 699.600 519.600 ;
        RECT 703.800 506.700 705.600 519.600 ;
        RECT 712.800 506.700 714.600 513.600 ;
        RECT 716.400 506.700 718.200 519.600 ;
        RECT 728.400 506.700 730.200 513.600 ;
        RECT 734.400 506.700 736.200 513.600 ;
        RECT 743.400 506.700 745.200 513.600 ;
        RECT 757.500 506.700 759.300 519.600 ;
        RECT -9.300 504.300 770.400 506.700 ;
        RECT -9.300 434.700 -0.300 504.300 ;
        RECT 10.800 497.400 12.600 504.300 ;
        RECT 16.800 497.400 18.600 504.300 ;
        RECT 22.800 497.400 24.600 504.300 ;
        RECT 37.800 493.200 39.600 504.300 ;
        RECT 49.800 498.000 51.600 504.300 ;
        RECT 55.800 497.400 57.600 504.300 ;
        RECT 61.800 497.400 63.600 504.300 ;
        RECT 67.800 497.400 69.600 504.300 ;
        RECT 71.400 497.400 73.200 504.300 ;
        RECT 77.400 498.000 79.200 504.300 ;
        RECT 87.300 491.400 89.100 504.300 ;
        RECT 94.800 497.400 96.600 504.300 ;
        RECT 103.800 497.400 105.600 504.300 ;
        RECT 109.800 497.400 111.600 504.300 ;
        RECT 116.400 497.400 118.200 504.300 ;
        RECT 123.900 491.400 125.700 504.300 ;
        RECT 132.300 491.400 134.100 504.300 ;
        RECT 139.800 497.400 141.600 504.300 ;
        RECT 149.400 497.400 151.200 504.300 ;
        RECT 156.900 491.400 158.700 504.300 ;
        RECT 164.400 497.400 166.200 504.300 ;
        RECT 171.900 491.400 173.700 504.300 ;
        RECT 176.400 497.400 178.200 504.300 ;
        RECT 193.800 493.200 195.600 504.300 ;
        RECT 200.400 497.400 202.200 504.300 ;
        RECT 206.400 497.400 208.200 504.300 ;
        RECT 215.400 497.400 217.200 504.300 ;
        RECT 224.400 491.400 226.200 504.300 ;
        RECT 234.900 491.400 236.700 504.300 ;
        RECT 248.400 497.400 250.200 504.300 ;
        RECT 255.900 491.400 257.700 504.300 ;
        RECT 271.800 491.400 273.600 504.300 ;
        RECT 286.800 491.400 288.600 504.300 ;
        RECT 301.800 493.500 303.600 504.300 ;
        RECT 311.550 500.400 313.350 504.300 ;
        RECT 320.250 497.400 322.050 504.300 ;
        RECT 326.850 497.400 328.650 504.300 ;
        RECT 337.050 497.400 338.850 504.300 ;
        RECT 347.700 491.400 349.500 504.300 ;
        RECT 356.400 497.400 358.200 504.300 ;
        RECT 362.400 497.400 364.200 504.300 ;
        RECT 371.400 497.400 373.200 504.300 ;
        RECT 378.900 491.400 380.700 504.300 ;
        RECT 389.400 497.400 391.200 504.300 ;
        RECT 396.900 491.400 398.700 504.300 ;
        RECT 406.200 491.400 408.000 504.300 ;
        RECT 412.800 497.400 414.600 504.300 ;
        RECT 421.800 491.400 423.600 504.300 ;
        RECT 428.550 500.400 430.350 504.300 ;
        RECT 437.250 497.400 439.050 504.300 ;
        RECT 443.850 497.400 445.650 504.300 ;
        RECT 454.050 497.400 455.850 504.300 ;
        RECT 463.800 491.400 465.600 504.300 ;
        RECT 469.800 491.400 471.600 504.300 ;
        RECT 475.800 491.400 477.600 504.300 ;
        RECT 481.800 491.400 483.600 504.300 ;
        RECT 487.800 491.400 489.600 504.300 ;
        RECT 494.400 497.400 496.200 504.300 ;
        RECT 501.900 491.400 503.700 504.300 ;
        RECT 511.800 497.400 513.600 504.300 ;
        RECT 515.400 497.400 517.200 504.300 ;
        RECT 521.400 497.400 523.200 504.300 ;
        RECT 535.800 493.200 537.600 504.300 ;
        RECT 547.800 498.000 549.600 504.300 ;
        RECT 553.800 497.400 555.600 504.300 ;
        RECT 557.400 491.400 559.200 504.300 ;
        RECT 569.400 497.400 571.200 504.300 ;
        RECT 575.400 497.400 577.200 504.300 ;
        RECT 584.400 493.500 586.200 504.300 ;
        RECT 601.800 497.400 603.600 504.300 ;
        RECT 607.800 497.400 609.600 504.300 ;
        RECT 614.400 491.400 616.200 504.300 ;
        RECT 631.800 497.400 633.600 504.300 ;
        RECT 639.300 491.400 641.100 504.300 ;
        RECT 646.800 497.400 648.600 504.300 ;
        RECT 657.300 491.400 659.100 504.300 ;
        RECT 667.800 491.400 669.600 504.300 ;
        RECT 671.400 491.400 673.200 504.300 ;
        RECT 683.400 497.400 685.200 504.300 ;
        RECT 689.400 497.400 691.200 504.300 ;
        RECT 698.400 497.400 700.200 504.300 ;
        RECT 705.900 491.400 707.700 504.300 ;
        RECT 711.300 491.400 713.100 504.300 ;
        RECT 718.800 497.400 720.600 504.300 ;
        RECT 725.400 491.400 727.200 504.300 ;
        RECT 747.300 491.550 749.100 504.300 ;
        RECT 755.400 497.400 757.200 504.300 ;
        RECT 762.000 491.400 763.800 504.300 ;
        RECT 7.800 434.700 9.600 441.600 ;
        RECT 14.400 434.700 16.200 441.600 ;
        RECT 21.900 434.700 23.700 447.600 ;
        RECT 26.400 434.700 28.200 441.600 ;
        RECT 33.000 434.700 34.800 447.600 ;
        RECT 49.800 434.700 51.600 441.000 ;
        RECT 55.800 434.700 57.600 441.600 ;
        RECT 59.400 434.700 61.200 441.600 ;
        RECT 73.800 434.700 75.600 441.600 ;
        RECT 80.400 434.700 82.200 441.600 ;
        RECT 86.400 434.700 88.200 441.000 ;
        RECT 98.400 434.700 100.200 441.600 ;
        RECT 109.800 434.700 111.600 441.600 ;
        RECT 115.800 434.700 117.600 441.600 ;
        RECT 119.400 434.700 121.200 441.600 ;
        RECT 125.400 434.700 127.200 441.000 ;
        RECT 137.400 434.700 139.200 441.600 ;
        RECT 147.300 434.700 149.100 447.600 ;
        RECT 154.800 434.700 156.600 441.600 ;
        RECT 164.400 434.700 166.200 441.600 ;
        RECT 170.400 434.700 172.200 441.000 ;
        RECT 187.800 434.700 189.600 447.600 ;
        RECT 191.400 434.700 193.200 447.600 ;
        RECT 206.400 434.700 208.200 441.600 ;
        RECT 212.400 434.700 214.200 441.600 ;
        RECT 218.400 434.700 220.200 447.600 ;
        RECT 230.400 434.700 232.200 447.600 ;
        RECT 242.400 434.700 244.200 441.600 ;
        RECT 249.000 434.700 250.800 447.600 ;
        RECT 265.800 434.700 267.600 447.600 ;
        RECT 272.400 434.700 274.200 447.600 ;
        RECT 287.400 434.700 289.200 441.600 ;
        RECT 296.400 434.700 298.200 441.600 ;
        RECT 302.400 434.700 304.200 441.600 ;
        RECT 308.400 434.700 310.200 441.600 ;
        RECT 320.400 434.700 322.200 445.500 ;
        RECT 338.400 434.700 340.200 445.800 ;
        RECT 358.800 434.700 360.600 445.800 ;
        RECT 368.550 434.700 370.350 438.600 ;
        RECT 377.250 434.700 379.050 441.600 ;
        RECT 383.850 434.700 385.650 441.600 ;
        RECT 394.050 434.700 395.850 441.600 ;
        RECT 412.800 434.700 414.600 445.800 ;
        RECT 420.300 434.700 422.100 447.600 ;
        RECT 427.800 434.700 429.600 441.600 ;
        RECT 436.800 434.700 438.600 447.600 ;
        RECT 442.800 434.700 444.600 447.600 ;
        RECT 448.800 434.700 450.600 447.600 ;
        RECT 454.800 434.700 456.600 447.600 ;
        RECT 460.800 434.700 462.600 447.600 ;
        RECT 469.800 434.700 471.600 441.600 ;
        RECT 475.800 434.700 477.600 441.600 ;
        RECT 481.800 434.700 483.600 441.600 ;
        RECT 487.800 434.700 489.600 441.600 ;
        RECT 493.800 434.700 495.600 441.600 ;
        RECT 499.800 434.700 501.600 441.600 ;
        RECT 503.400 434.700 505.200 441.600 ;
        RECT 509.400 434.700 511.200 441.000 ;
        RECT 523.800 434.700 525.600 441.000 ;
        RECT 529.800 434.700 531.600 441.600 ;
        RECT 541.800 434.700 543.600 441.600 ;
        RECT 551.400 434.700 553.200 441.600 ;
        RECT 558.900 434.700 560.700 447.600 ;
        RECT 563.400 434.700 565.200 441.600 ;
        RECT 573.300 434.700 575.100 447.600 ;
        RECT 580.800 434.700 582.600 441.600 ;
        RECT 595.800 434.700 597.600 441.000 ;
        RECT 601.800 434.700 603.600 441.600 ;
        RECT 613.800 434.700 615.600 445.800 ;
        RECT 631.800 434.700 633.600 445.500 ;
        RECT 640.800 434.700 642.600 441.600 ;
        RECT 646.800 434.700 648.600 441.600 ;
        RECT 650.400 434.700 652.200 441.600 ;
        RECT 660.300 434.700 662.100 447.600 ;
        RECT 667.800 434.700 669.600 441.600 ;
        RECT 679.800 434.700 681.600 441.000 ;
        RECT 685.800 434.700 687.600 441.600 ;
        RECT 697.800 434.700 699.600 441.600 ;
        RECT 704.400 434.700 706.200 445.800 ;
        RECT 719.400 434.700 721.200 447.600 ;
        RECT 738.900 434.700 740.700 447.450 ;
        RECT 750.300 434.700 752.100 447.600 ;
        RECT 757.800 434.700 759.600 441.600 ;
        RECT -9.300 432.300 770.400 434.700 ;
        RECT -9.300 362.700 -0.300 432.300 ;
        RECT 7.800 425.400 9.600 432.300 ;
        RECT 14.400 425.400 16.200 432.300 ;
        RECT 21.900 419.400 23.700 432.300 ;
        RECT 30.300 419.400 32.100 432.300 ;
        RECT 37.800 425.400 39.600 432.300 ;
        RECT 49.800 425.400 51.600 432.300 ;
        RECT 55.800 425.400 57.600 432.300 ;
        RECT 64.800 426.000 66.600 432.300 ;
        RECT 70.800 425.400 72.600 432.300 ;
        RECT 74.400 425.400 76.200 432.300 ;
        RECT 80.400 426.000 82.200 432.300 ;
        RECT 91.800 425.400 93.600 432.300 ;
        RECT 97.800 425.400 99.600 432.300 ;
        RECT 101.400 425.400 103.200 432.300 ;
        RECT 107.400 426.000 109.200 432.300 ;
        RECT 118.800 425.400 120.600 432.300 ;
        RECT 124.800 425.400 126.600 432.300 ;
        RECT 131.400 425.400 133.200 432.300 ;
        RECT 138.000 419.400 139.800 432.300 ;
        RECT 147.300 419.400 149.100 432.300 ;
        RECT 154.800 425.400 156.600 432.300 ;
        RECT 161.400 425.400 163.200 432.300 ;
        RECT 167.400 425.400 169.200 432.300 ;
        RECT 173.400 425.400 175.200 432.300 ;
        RECT 179.400 426.000 181.200 432.300 ;
        RECT 188.400 425.400 190.200 432.300 ;
        RECT 194.400 425.400 196.200 432.300 ;
        RECT 203.400 425.400 205.200 432.300 ;
        RECT 213.300 419.400 215.100 432.300 ;
        RECT 220.800 425.400 222.600 432.300 ;
        RECT 228.300 419.400 230.100 432.300 ;
        RECT 235.800 425.400 237.600 432.300 ;
        RECT 245.400 425.400 247.200 432.300 ;
        RECT 254.400 425.400 256.200 432.300 ;
        RECT 260.400 425.400 262.200 432.300 ;
        RECT 267.300 419.400 269.100 432.300 ;
        RECT 274.800 425.400 276.600 432.300 ;
        RECT 289.800 421.200 291.600 432.300 ;
        RECT 302.400 425.400 304.200 432.300 ;
        RECT 309.900 419.400 311.700 432.300 ;
        RECT 317.400 425.400 319.200 432.300 ;
        RECT 324.900 419.400 326.700 432.300 ;
        RECT 332.400 425.400 334.200 432.300 ;
        RECT 339.900 419.400 341.700 432.300 ;
        RECT 344.400 425.400 346.200 432.300 ;
        RECT 350.400 425.400 352.200 432.300 ;
        RECT 364.800 421.200 366.600 432.300 ;
        RECT 374.400 425.400 376.200 432.300 ;
        RECT 381.900 419.400 383.700 432.300 ;
        RECT 391.800 419.400 393.600 432.300 ;
        RECT 397.800 419.400 399.600 432.300 ;
        RECT 412.800 421.500 414.600 432.300 ;
        RECT 419.400 425.400 421.200 432.300 ;
        RECT 431.700 419.400 433.500 432.300 ;
        RECT 445.500 419.400 447.300 432.300 ;
        RECT 457.800 425.400 459.600 432.300 ;
        RECT 463.800 425.400 465.600 432.300 ;
        RECT 472.800 425.400 474.600 432.300 ;
        RECT 479.400 425.400 481.200 432.300 ;
        RECT 486.900 419.400 488.700 432.300 ;
        RECT 511.800 422.400 513.600 432.300 ;
        RECT 524.400 425.400 526.200 432.300 ;
        RECT 531.900 419.400 533.700 432.300 ;
        RECT 536.400 425.400 538.200 432.300 ;
        RECT 548.700 419.400 550.500 432.300 ;
        RECT 565.800 426.000 567.600 432.300 ;
        RECT 571.800 425.400 573.600 432.300 ;
        RECT 583.800 421.200 585.600 432.300 ;
        RECT 593.400 425.400 595.200 432.300 ;
        RECT 600.900 419.400 602.700 432.300 ;
        RECT 606.300 419.400 608.100 432.300 ;
        RECT 613.800 425.400 615.600 432.300 ;
        RECT 625.800 426.000 627.600 432.300 ;
        RECT 631.800 425.400 633.600 432.300 ;
        RECT 638.400 421.200 640.200 432.300 ;
        RECT 653.400 421.500 655.200 432.300 ;
        RECT 670.800 425.400 672.600 432.300 ;
        RECT 676.800 425.400 678.600 432.300 ;
        RECT 688.800 421.200 690.600 432.300 ;
        RECT 695.400 425.400 697.200 432.300 ;
        RECT 701.400 426.000 703.200 432.300 ;
        RECT 718.800 421.200 720.600 432.300 ;
        RECT 725.400 425.400 727.200 432.300 ;
        RECT 731.400 426.000 733.200 432.300 ;
        RECT 740.400 425.400 742.200 432.300 ;
        RECT 746.400 426.000 748.200 432.300 ;
        RECT 9.300 362.700 11.100 375.450 ;
        RECT 19.800 362.700 21.600 369.600 ;
        RECT 25.800 362.700 27.600 369.600 ;
        RECT 32.400 362.700 34.200 369.600 ;
        RECT 38.400 362.700 40.200 369.600 ;
        RECT 44.400 362.700 46.200 369.600 ;
        RECT 56.400 362.700 58.200 369.600 ;
        RECT 63.900 362.700 65.700 375.600 ;
        RECT 73.800 362.700 75.600 369.600 ;
        RECT 83.400 362.700 85.200 373.800 ;
        RECT 95.400 362.700 97.200 369.600 ;
        RECT 101.400 362.700 103.200 369.000 ;
        RECT 110.400 362.700 112.200 369.600 ;
        RECT 116.400 362.700 118.200 369.000 ;
        RECT 130.800 362.700 132.600 369.600 ;
        RECT 144.300 362.700 146.100 375.450 ;
        RECT 152.400 362.700 154.200 369.600 ;
        RECT 158.400 362.700 160.200 369.000 ;
        RECT 187.800 362.700 189.600 372.600 ;
        RECT 194.400 362.700 196.200 369.600 ;
        RECT 207.300 362.700 209.100 375.600 ;
        RECT 214.800 362.700 216.600 369.600 ;
        RECT 222.300 362.700 224.100 375.600 ;
        RECT 229.800 362.700 231.600 369.600 ;
        RECT 247.800 362.700 249.600 373.800 ;
        RECT 257.400 362.700 259.200 369.600 ;
        RECT 264.900 362.700 266.700 375.600 ;
        RECT 280.800 362.700 282.600 373.500 ;
        RECT 295.800 362.700 297.600 369.600 ;
        RECT 303.150 362.700 304.950 369.600 ;
        RECT 313.350 362.700 315.150 369.600 ;
        RECT 319.950 362.700 321.750 369.600 ;
        RECT 328.650 362.700 330.450 366.600 ;
        RECT 343.800 362.700 345.600 373.800 ;
        RECT 364.800 362.700 366.600 373.500 ;
        RECT 376.800 362.700 378.600 369.600 ;
        RECT 383.550 362.700 385.350 366.600 ;
        RECT 392.250 362.700 394.050 369.600 ;
        RECT 398.850 362.700 400.650 369.600 ;
        RECT 409.050 362.700 410.850 369.600 ;
        RECT 419.550 362.700 421.350 366.600 ;
        RECT 428.250 362.700 430.050 369.600 ;
        RECT 434.850 362.700 436.650 369.600 ;
        RECT 445.050 362.700 446.850 369.600 ;
        RECT 455.400 362.700 457.200 369.600 ;
        RECT 462.900 362.700 464.700 375.600 ;
        RECT 475.800 362.700 477.600 373.800 ;
        RECT 482.400 362.700 484.200 369.600 ;
        RECT 488.400 362.700 490.200 369.000 ;
        RECT 500.400 362.700 502.200 369.600 ;
        RECT 512.400 362.700 514.200 369.600 ;
        RECT 519.000 362.700 520.800 375.600 ;
        RECT 532.800 362.700 534.600 369.600 ;
        RECT 541.800 362.700 543.600 369.000 ;
        RECT 547.800 362.700 549.600 369.600 ;
        RECT 559.800 362.700 561.600 369.000 ;
        RECT 565.800 362.700 567.600 369.600 ;
        RECT 572.400 362.700 574.200 369.600 ;
        RECT 579.900 362.700 581.700 375.600 ;
        RECT 588.300 362.700 590.100 375.600 ;
        RECT 595.800 362.700 597.600 369.600 ;
        RECT 602.400 362.700 604.200 369.600 ;
        RECT 616.800 362.700 618.600 369.000 ;
        RECT 622.800 362.700 624.600 369.600 ;
        RECT 626.400 362.700 628.200 369.600 ;
        RECT 632.400 362.700 634.200 369.000 ;
        RECT 646.800 362.700 648.600 369.000 ;
        RECT 652.800 362.700 654.600 369.600 ;
        RECT 661.800 362.700 663.600 369.600 ;
        RECT 668.400 362.700 670.200 369.600 ;
        RECT 675.900 362.700 677.700 375.600 ;
        RECT 691.800 362.700 693.600 373.800 ;
        RECT 703.800 362.700 705.600 369.000 ;
        RECT 709.800 362.700 711.600 369.600 ;
        RECT 717.300 362.700 719.100 375.600 ;
        RECT 724.800 362.700 726.600 369.600 ;
        RECT 736.800 362.700 738.600 369.600 ;
        RECT 741.300 362.700 743.100 375.600 ;
        RECT 748.800 362.700 750.600 369.600 ;
        RECT -9.300 360.300 770.400 362.700 ;
        RECT -9.300 290.700 -0.300 360.300 ;
        RECT 10.800 353.400 12.600 360.300 ;
        RECT 15.300 347.400 17.100 360.300 ;
        RECT 22.800 353.400 24.600 360.300 ;
        RECT 36.300 347.550 38.100 360.300 ;
        RECT 47.400 353.400 49.200 360.300 ;
        RECT 54.000 347.400 55.800 360.300 ;
        RECT 62.400 353.400 64.200 360.300 ;
        RECT 68.400 354.000 70.200 360.300 ;
        RECT 77.400 353.400 79.200 360.300 ;
        RECT 83.400 354.000 85.200 360.300 ;
        RECT 93.300 347.400 95.100 360.300 ;
        RECT 100.800 353.400 102.600 360.300 ;
        RECT 115.800 354.000 117.600 360.300 ;
        RECT 121.800 353.400 123.600 360.300 ;
        RECT 125.400 353.400 127.200 360.300 ;
        RECT 137.400 349.200 139.200 360.300 ;
        RECT 150.300 347.400 152.100 360.300 ;
        RECT 157.800 353.400 159.600 360.300 ;
        RECT 172.800 353.400 174.600 360.300 ;
        RECT 187.800 347.400 189.600 360.300 ;
        RECT 196.800 353.400 198.600 360.300 ;
        RECT 208.800 349.200 210.600 360.300 ;
        RECT 215.400 347.400 217.200 360.300 ;
        RECT 238.800 349.500 240.600 360.300 ;
        RECT 250.800 353.400 252.600 360.300 ;
        RECT 258.150 353.400 259.950 360.300 ;
        RECT 268.350 353.400 270.150 360.300 ;
        RECT 274.950 353.400 276.750 360.300 ;
        RECT 283.650 356.400 285.450 360.300 ;
        RECT 293.700 347.400 295.500 360.300 ;
        RECT 308.400 353.400 310.200 360.300 ;
        RECT 315.900 347.400 317.700 360.300 ;
        RECT 331.800 349.500 333.600 360.300 ;
        RECT 343.800 353.400 345.600 360.300 ;
        RECT 351.150 353.400 352.950 360.300 ;
        RECT 361.350 353.400 363.150 360.300 ;
        RECT 367.950 353.400 369.750 360.300 ;
        RECT 376.650 356.400 378.450 360.300 ;
        RECT 386.400 353.400 388.200 360.300 ;
        RECT 393.000 347.400 394.800 360.300 ;
        RECT 406.800 353.400 408.600 360.300 ;
        RECT 412.800 353.400 414.600 360.300 ;
        RECT 424.800 353.400 426.600 360.300 ;
        RECT 429.300 347.400 431.100 360.300 ;
        RECT 436.800 353.400 438.600 360.300 ;
        RECT 445.800 353.400 447.600 360.300 ;
        RECT 451.800 353.400 453.600 360.300 ;
        RECT 463.800 353.400 465.600 360.300 ;
        RECT 467.400 353.400 469.200 360.300 ;
        RECT 473.400 353.400 475.200 360.300 ;
        RECT 479.400 347.400 481.200 360.300 ;
        RECT 499.800 354.000 501.600 360.300 ;
        RECT 505.800 353.400 507.600 360.300 ;
        RECT 512.400 353.400 514.200 360.300 ;
        RECT 519.900 347.400 521.700 360.300 ;
        RECT 525.300 347.400 527.100 360.300 ;
        RECT 532.800 353.400 534.600 360.300 ;
        RECT 542.400 349.200 544.200 360.300 ;
        RECT 557.400 353.400 559.200 360.300 ;
        RECT 564.900 347.400 566.700 360.300 ;
        RECT 589.800 350.400 591.600 360.300 ;
        RECT 596.400 353.400 598.200 360.300 ;
        RECT 613.800 349.200 615.600 360.300 ;
        RECT 623.400 353.400 625.200 360.300 ;
        RECT 629.400 354.000 631.200 360.300 ;
        RECT 639.300 347.400 641.100 360.300 ;
        RECT 646.800 353.400 648.600 360.300 ;
        RECT 661.800 349.200 663.600 360.300 ;
        RECT 673.800 354.000 675.600 360.300 ;
        RECT 679.800 353.400 681.600 360.300 ;
        RECT 691.800 354.000 693.600 360.300 ;
        RECT 697.800 353.400 699.600 360.300 ;
        RECT 709.800 354.000 711.600 360.300 ;
        RECT 715.800 353.400 717.600 360.300 ;
        RECT 725.400 353.400 727.200 360.300 ;
        RECT 732.900 347.400 734.700 360.300 ;
        RECT 738.300 347.400 740.100 360.300 ;
        RECT 745.800 353.400 747.600 360.300 ;
        RECT 752.400 353.400 754.200 360.300 ;
        RECT 758.400 354.000 760.200 360.300 ;
        RECT 10.800 290.700 12.600 297.600 ;
        RECT 16.800 290.700 18.600 297.600 ;
        RECT 22.800 290.700 24.600 297.600 ;
        RECT 26.400 290.700 28.200 297.600 ;
        RECT 32.400 290.700 34.200 297.600 ;
        RECT 41.400 290.700 43.200 297.600 ;
        RECT 47.400 290.700 49.200 297.000 ;
        RECT 56.400 290.700 58.200 297.600 ;
        RECT 62.400 290.700 64.200 297.600 ;
        RECT 71.400 290.700 73.200 297.600 ;
        RECT 78.900 290.700 80.700 303.600 ;
        RECT 83.400 290.700 85.200 297.600 ;
        RECT 89.400 290.700 91.200 297.600 ;
        RECT 99.900 290.700 101.700 303.450 ;
        RECT 115.800 290.700 117.600 297.600 ;
        RECT 121.800 290.700 123.600 297.600 ;
        RECT 130.800 290.700 132.600 297.000 ;
        RECT 136.800 290.700 138.600 297.600 ;
        RECT 140.400 290.700 142.200 303.600 ;
        RECT 163.800 290.700 165.600 301.800 ;
        RECT 181.800 290.700 183.600 301.800 ;
        RECT 189.300 290.700 191.100 303.600 ;
        RECT 196.800 290.700 198.600 297.600 ;
        RECT 203.400 290.700 205.200 297.600 ;
        RECT 209.400 290.700 211.200 297.600 ;
        RECT 218.400 290.700 220.200 301.500 ;
        RECT 239.400 290.700 241.200 301.800 ;
        RECT 254.400 290.700 256.200 297.600 ;
        RECT 261.900 290.700 263.700 303.600 ;
        RECT 267.300 290.700 269.100 303.600 ;
        RECT 274.800 290.700 276.600 297.600 ;
        RECT 281.400 290.700 283.200 297.600 ;
        RECT 295.800 290.700 297.600 297.000 ;
        RECT 301.800 290.700 303.600 297.600 ;
        RECT 313.800 290.700 315.600 303.600 ;
        RECT 318.300 290.700 320.100 303.600 ;
        RECT 325.800 290.700 327.600 297.600 ;
        RECT 335.700 290.700 337.500 303.600 ;
        RECT 347.400 290.700 349.200 297.600 ;
        RECT 353.400 290.700 355.200 297.600 ;
        RECT 359.400 290.700 361.200 297.600 ;
        RECT 365.400 290.700 367.200 297.600 ;
        RECT 371.400 290.700 373.200 297.600 ;
        RECT 378.000 290.700 379.800 303.600 ;
        RECT 392.700 290.700 394.500 303.600 ;
        RECT 404.700 290.700 406.500 303.600 ;
        RECT 416.400 290.700 418.200 297.600 ;
        RECT 423.900 290.700 425.700 303.600 ;
        RECT 433.800 290.700 435.600 297.600 ;
        RECT 439.800 290.700 441.600 297.600 ;
        RECT 443.400 290.700 445.200 297.600 ;
        RECT 452.400 290.700 454.200 297.600 ;
        RECT 458.400 290.700 460.200 297.000 ;
        RECT 467.400 290.700 469.200 297.600 ;
        RECT 473.400 290.700 475.200 297.600 ;
        RECT 479.400 290.700 481.200 297.600 ;
        RECT 485.400 290.700 487.200 297.000 ;
        RECT 496.800 290.700 498.600 297.600 ;
        RECT 502.800 290.700 504.600 297.600 ;
        RECT 506.400 290.700 508.200 297.600 ;
        RECT 513.000 290.700 514.800 303.600 ;
        RECT 523.800 290.700 525.600 297.600 ;
        RECT 529.800 290.700 531.600 297.600 ;
        RECT 541.800 290.700 543.600 301.800 ;
        RECT 550.800 290.700 552.600 297.600 ;
        RECT 556.800 290.700 558.600 297.600 ;
        RECT 565.800 290.700 567.600 297.000 ;
        RECT 571.800 290.700 573.600 297.600 ;
        RECT 575.400 290.700 577.200 297.600 ;
        RECT 587.400 290.700 589.200 297.600 ;
        RECT 594.900 290.700 596.700 303.600 ;
        RECT 603.300 290.700 605.100 303.600 ;
        RECT 610.800 290.700 612.600 297.600 ;
        RECT 628.800 290.700 630.600 301.800 ;
        RECT 643.800 290.700 645.600 297.000 ;
        RECT 649.800 290.700 651.600 297.600 ;
        RECT 658.800 290.700 660.600 297.000 ;
        RECT 664.800 290.700 666.600 297.600 ;
        RECT 676.800 290.700 678.600 301.800 ;
        RECT 691.800 290.700 693.600 297.000 ;
        RECT 697.800 290.700 699.600 297.600 ;
        RECT 701.400 290.700 703.200 297.600 ;
        RECT 707.400 290.700 709.200 297.600 ;
        RECT 718.800 290.700 720.600 297.000 ;
        RECT 724.800 290.700 726.600 297.600 ;
        RECT 731.400 290.700 733.200 301.800 ;
        RECT 749.400 290.700 751.200 301.800 ;
        RECT -9.300 288.300 770.400 290.700 ;
        RECT -9.300 218.700 -0.300 288.300 ;
        RECT 5.400 281.400 7.200 288.300 ;
        RECT 12.900 275.400 14.700 288.300 ;
        RECT 19.800 281.400 21.600 288.300 ;
        RECT 25.800 281.400 27.600 288.300 ;
        RECT 32.400 281.400 34.200 288.300 ;
        RECT 38.400 282.000 40.200 288.300 ;
        RECT 49.800 281.400 51.600 288.300 ;
        RECT 55.800 281.400 57.600 288.300 ;
        RECT 59.400 281.400 61.200 288.300 ;
        RECT 65.400 282.000 67.200 288.300 ;
        RECT 82.800 277.200 84.600 288.300 ;
        RECT 92.400 281.400 94.200 288.300 ;
        RECT 98.400 281.400 100.200 288.300 ;
        RECT 115.800 275.400 117.600 288.300 ;
        RECT 122.400 281.400 124.200 288.300 ;
        RECT 129.900 275.400 131.700 288.300 ;
        RECT 134.400 275.400 136.200 288.300 ;
        RECT 144.900 275.400 146.700 288.300 ;
        RECT 160.800 277.200 162.600 288.300 ;
        RECT 167.400 275.400 169.200 288.300 ;
        RECT 179.400 275.400 181.200 288.300 ;
        RECT 194.400 281.400 196.200 288.300 ;
        RECT 200.400 281.400 202.200 288.300 ;
        RECT 206.400 281.400 208.200 288.300 ;
        RECT 212.400 281.400 214.200 288.300 ;
        RECT 221.400 281.400 223.200 288.300 ;
        RECT 227.400 281.400 229.200 288.300 ;
        RECT 233.400 281.400 235.200 288.300 ;
        RECT 239.400 281.400 241.200 288.300 ;
        RECT 245.400 275.400 247.200 288.300 ;
        RECT 265.800 277.200 267.600 288.300 ;
        RECT 280.500 275.400 282.300 288.300 ;
        RECT 289.800 275.400 291.600 288.300 ;
        RECT 295.800 275.400 297.600 288.300 ;
        RECT 299.400 275.400 301.200 288.300 ;
        RECT 313.800 275.400 315.600 288.300 ;
        RECT 320.700 275.400 322.500 288.300 ;
        RECT 334.800 282.000 336.600 288.300 ;
        RECT 340.800 281.400 342.600 288.300 ;
        RECT 346.800 281.400 348.600 288.300 ;
        RECT 352.800 281.400 354.600 288.300 ;
        RECT 367.800 277.200 369.600 288.300 ;
        RECT 374.400 281.400 376.200 288.300 ;
        RECT 380.400 281.400 382.200 288.300 ;
        RECT 389.700 275.400 391.500 288.300 ;
        RECT 403.200 275.400 405.000 288.300 ;
        RECT 409.800 281.400 411.600 288.300 ;
        RECT 413.400 275.400 415.200 288.300 ;
        RECT 428.700 275.400 430.500 288.300 ;
        RECT 442.200 275.400 444.000 288.300 ;
        RECT 448.800 281.400 450.600 288.300 ;
        RECT 452.400 281.400 454.200 288.300 ;
        RECT 459.000 275.400 460.800 288.300 ;
        RECT 481.800 277.500 483.600 288.300 ;
        RECT 493.200 275.400 495.000 288.300 ;
        RECT 499.800 281.400 501.600 288.300 ;
        RECT 503.400 281.400 505.200 288.300 ;
        RECT 509.400 281.400 511.200 288.300 ;
        RECT 516.300 275.400 518.100 288.300 ;
        RECT 523.800 281.400 525.600 288.300 ;
        RECT 530.400 281.400 532.200 288.300 ;
        RECT 536.400 281.400 538.200 288.300 ;
        RECT 543.300 275.400 545.100 288.300 ;
        RECT 550.800 281.400 552.600 288.300 ;
        RECT 557.400 275.400 559.200 288.300 ;
        RECT 572.700 275.400 574.500 288.300 ;
        RECT 583.800 281.400 585.600 288.300 ;
        RECT 589.800 281.400 591.600 288.300 ;
        RECT 596.400 277.500 598.200 288.300 ;
        RECT 622.800 275.400 624.600 288.300 ;
        RECT 626.400 281.400 628.200 288.300 ;
        RECT 632.400 281.400 634.200 288.300 ;
        RECT 643.800 281.400 645.600 288.300 ;
        RECT 649.800 281.400 651.600 288.300 ;
        RECT 654.300 275.400 656.100 288.300 ;
        RECT 661.800 281.400 663.600 288.300 ;
        RECT 668.400 281.400 670.200 288.300 ;
        RECT 685.800 277.200 687.600 288.300 ;
        RECT 697.800 281.400 699.600 288.300 ;
        RECT 702.300 275.400 704.100 288.300 ;
        RECT 709.800 281.400 711.600 288.300 ;
        RECT 717.300 275.400 719.100 288.300 ;
        RECT 724.800 281.400 726.600 288.300 ;
        RECT 736.800 282.000 738.600 288.300 ;
        RECT 742.800 281.400 744.600 288.300 ;
        RECT 746.400 281.400 748.200 288.300 ;
        RECT 752.400 282.000 754.200 288.300 ;
        RECT 12.300 218.700 14.100 231.450 ;
        RECT 22.800 218.700 24.600 225.600 ;
        RECT 28.800 218.700 30.600 225.600 ;
        RECT 39.300 218.700 41.100 231.450 ;
        RECT 53.400 218.700 55.200 225.600 ;
        RECT 60.900 218.700 62.700 231.600 ;
        RECT 70.800 218.700 72.600 225.600 ;
        RECT 74.400 218.700 76.200 225.600 ;
        RECT 80.400 218.700 82.200 225.000 ;
        RECT 91.800 218.700 93.600 225.600 ;
        RECT 97.800 218.700 99.600 225.600 ;
        RECT 103.800 218.700 105.600 225.600 ;
        RECT 109.800 218.700 111.600 225.600 ;
        RECT 113.400 218.700 115.200 231.600 ;
        RECT 125.400 218.700 127.200 231.600 ;
        RECT 135.900 218.700 137.700 231.600 ;
        RECT 143.400 218.700 145.200 231.600 ;
        RECT 163.800 218.700 165.600 225.600 ;
        RECT 172.800 218.700 174.600 225.600 ;
        RECT 184.800 218.700 186.600 231.600 ;
        RECT 188.400 218.700 190.200 225.600 ;
        RECT 194.400 218.700 196.200 225.600 ;
        RECT 211.800 218.700 213.600 229.500 ;
        RECT 221.400 218.700 223.200 225.600 ;
        RECT 228.000 218.700 229.800 231.600 ;
        RECT 236.400 218.700 238.200 225.600 ;
        RECT 242.400 218.700 244.200 225.600 ;
        RECT 251.400 218.700 253.200 225.600 ;
        RECT 258.900 218.700 260.700 231.600 ;
        RECT 269.400 218.700 271.200 225.600 ;
        RECT 276.900 218.700 278.700 231.600 ;
        RECT 286.200 218.700 288.000 231.600 ;
        RECT 292.800 218.700 294.600 225.600 ;
        RECT 302.400 218.700 304.200 229.500 ;
        RECT 322.500 218.700 324.300 231.600 ;
        RECT 329.400 218.700 331.200 225.600 ;
        RECT 336.000 218.700 337.800 231.600 ;
        RECT 349.500 218.700 351.300 231.600 ;
        RECT 361.800 218.700 363.600 231.600 ;
        RECT 365.400 218.700 367.200 225.600 ;
        RECT 372.000 218.700 373.800 231.600 ;
        RECT 383.400 218.700 385.200 225.600 ;
        RECT 390.000 218.700 391.800 231.600 ;
        RECT 398.400 218.700 400.200 225.600 ;
        RECT 404.400 218.700 406.200 225.600 ;
        RECT 413.400 218.700 415.200 225.600 ;
        RECT 420.900 218.700 422.700 231.600 ;
        RECT 425.400 218.700 427.200 225.600 ;
        RECT 431.400 218.700 433.200 225.600 ;
        RECT 440.400 218.700 442.200 225.600 ;
        RECT 447.900 218.700 449.700 231.600 ;
        RECT 460.800 218.700 462.600 225.000 ;
        RECT 466.800 218.700 468.600 225.600 ;
        RECT 470.400 218.700 472.200 225.600 ;
        RECT 476.400 218.700 478.200 225.600 ;
        RECT 485.400 218.700 487.200 225.600 ;
        RECT 492.900 218.700 494.700 231.600 ;
        RECT 499.800 218.700 501.600 225.600 ;
        RECT 505.800 218.700 507.600 225.600 ;
        RECT 509.400 218.700 511.200 225.600 ;
        RECT 521.400 218.700 523.200 229.500 ;
        RECT 540.300 218.700 542.100 231.600 ;
        RECT 547.800 218.700 549.600 225.600 ;
        RECT 554.400 218.700 556.200 225.600 ;
        RECT 560.400 218.700 562.200 225.000 ;
        RECT 574.800 218.700 576.600 225.600 ;
        RECT 580.800 218.700 582.600 225.600 ;
        RECT 592.800 218.700 594.600 231.600 ;
        RECT 601.800 218.700 603.600 225.600 ;
        RECT 607.800 218.700 609.600 225.600 ;
        RECT 615.900 218.700 617.700 231.450 ;
        RECT 637.800 218.700 639.600 229.800 ;
        RECT 646.800 218.700 648.600 225.600 ;
        RECT 652.800 218.700 654.600 225.600 ;
        RECT 656.400 218.700 658.200 225.600 ;
        RECT 663.000 218.700 664.800 231.600 ;
        RECT 674.400 218.700 676.200 229.500 ;
        RECT 692.400 218.700 694.200 225.600 ;
        RECT 699.900 218.700 701.700 231.600 ;
        RECT 705.300 218.700 707.100 231.600 ;
        RECT 712.800 218.700 714.600 225.600 ;
        RECT 719.400 218.700 721.200 225.600 ;
        RECT 725.400 218.700 727.200 225.000 ;
        RECT 737.400 218.700 739.200 225.600 ;
        RECT 743.400 218.700 745.200 225.000 ;
        RECT 760.800 218.700 762.600 225.000 ;
        RECT 766.800 218.700 768.600 225.600 ;
        RECT -9.300 216.300 770.400 218.700 ;
        RECT -9.300 146.700 -0.300 216.300 ;
        RECT 5.400 209.400 7.200 216.300 ;
        RECT 12.900 203.400 14.700 216.300 ;
        RECT 22.800 209.400 24.600 216.300 ;
        RECT 27.300 203.400 29.100 216.300 ;
        RECT 34.800 209.400 36.600 216.300 ;
        RECT 41.400 209.400 43.200 216.300 ;
        RECT 47.400 210.000 49.200 216.300 ;
        RECT 64.800 209.400 66.600 216.300 ;
        RECT 76.800 205.200 78.600 216.300 ;
        RECT 83.400 209.400 85.200 216.300 ;
        RECT 89.400 209.400 91.200 216.300 ;
        RECT 101.400 209.400 103.200 216.300 ;
        RECT 108.900 203.400 110.700 216.300 ;
        RECT 124.800 203.400 126.600 216.300 ;
        RECT 133.800 209.400 135.600 216.300 ;
        RECT 142.200 203.400 144.000 216.300 ;
        RECT 148.800 209.400 150.600 216.300 ;
        RECT 153.300 203.400 155.100 216.300 ;
        RECT 160.800 209.400 162.600 216.300 ;
        RECT 175.800 203.400 177.600 216.300 ;
        RECT 179.400 203.400 181.200 216.300 ;
        RECT 189.900 203.400 191.700 216.300 ;
        RECT 197.400 209.400 199.200 216.300 ;
        RECT 203.400 209.400 205.200 216.300 ;
        RECT 209.400 209.400 211.200 216.300 ;
        RECT 215.400 209.400 217.200 216.300 ;
        RECT 221.400 209.400 223.200 216.300 ;
        RECT 227.400 209.400 229.200 216.300 ;
        RECT 236.400 205.500 238.200 216.300 ;
        RECT 259.800 205.200 261.600 216.300 ;
        RECT 271.800 210.000 273.600 216.300 ;
        RECT 277.800 209.400 279.600 216.300 ;
        RECT 281.400 209.400 283.200 216.300 ;
        RECT 287.400 209.400 289.200 216.300 ;
        RECT 296.400 209.400 298.200 216.300 ;
        RECT 302.400 209.400 304.200 216.300 ;
        RECT 308.400 209.400 310.200 216.300 ;
        RECT 315.000 203.400 316.800 216.300 ;
        RECT 325.800 209.400 327.600 216.300 ;
        RECT 331.800 209.400 333.600 216.300 ;
        RECT 341.400 209.400 343.200 216.300 ;
        RECT 348.900 203.400 350.700 216.300 ;
        RECT 353.400 209.400 355.200 216.300 ;
        RECT 359.400 210.000 361.200 216.300 ;
        RECT 371.400 209.400 373.200 216.300 ;
        RECT 378.900 203.400 380.700 216.300 ;
        RECT 391.800 203.400 393.600 216.300 ;
        RECT 403.800 205.200 405.600 216.300 ;
        RECT 418.800 203.400 420.600 216.300 ;
        RECT 430.500 203.400 432.300 216.300 ;
        RECT 441.300 203.400 443.100 216.300 ;
        RECT 448.800 209.400 450.600 216.300 ;
        RECT 457.800 209.400 459.600 216.300 ;
        RECT 463.800 209.400 465.600 216.300 ;
        RECT 467.400 209.400 469.200 216.300 ;
        RECT 473.400 210.000 475.200 216.300 ;
        RECT 483.300 203.400 485.100 216.300 ;
        RECT 490.800 209.400 492.600 216.300 ;
        RECT 498.300 203.400 500.100 216.300 ;
        RECT 505.800 209.400 507.600 216.300 ;
        RECT 515.400 209.400 517.200 216.300 ;
        RECT 524.400 209.400 526.200 216.300 ;
        RECT 533.400 209.400 535.200 216.300 ;
        RECT 539.400 210.000 541.200 216.300 ;
        RECT 550.800 209.400 552.600 216.300 ;
        RECT 556.800 209.400 558.600 216.300 ;
        RECT 560.400 209.400 562.200 216.300 ;
        RECT 567.000 203.400 568.800 216.300 ;
        RECT 578.400 205.500 580.200 216.300 ;
        RECT 596.400 209.400 598.200 216.300 ;
        RECT 603.000 203.400 604.800 216.300 ;
        RECT 612.300 203.400 614.100 216.300 ;
        RECT 619.800 209.400 621.600 216.300 ;
        RECT 626.400 209.400 628.200 216.300 ;
        RECT 635.400 209.400 637.200 216.300 ;
        RECT 641.400 209.400 643.200 216.300 ;
        RECT 647.400 209.400 649.200 216.300 ;
        RECT 653.400 210.000 655.200 216.300 ;
        RECT 668.400 205.200 670.200 216.300 ;
        RECT 680.400 209.400 682.200 216.300 ;
        RECT 686.400 210.000 688.200 216.300 ;
        RECT 698.400 205.200 700.200 216.300 ;
        RECT 711.300 203.400 713.100 216.300 ;
        RECT 718.800 209.400 720.600 216.300 ;
        RECT 725.400 209.400 727.200 216.300 ;
        RECT 731.400 210.000 733.200 216.300 ;
        RECT 740.400 209.400 742.200 216.300 ;
        RECT 746.400 210.000 748.200 216.300 ;
        RECT 758.400 209.400 760.200 216.300 ;
        RECT 765.900 203.400 767.700 216.300 ;
        RECT 13.800 146.700 15.600 159.600 ;
        RECT 21.900 146.700 23.700 159.450 ;
        RECT 40.800 146.700 42.600 153.000 ;
        RECT 46.800 146.700 48.600 153.600 ;
        RECT 50.400 146.700 52.200 153.600 ;
        RECT 60.300 146.700 62.100 159.600 ;
        RECT 67.800 146.700 69.600 153.600 ;
        RECT 81.300 146.700 83.100 159.450 ;
        RECT 89.400 146.700 91.200 153.600 ;
        RECT 95.400 146.700 97.200 153.600 ;
        RECT 109.800 146.700 111.600 153.000 ;
        RECT 115.800 146.700 117.600 153.600 ;
        RECT 127.800 146.700 129.600 153.600 ;
        RECT 136.800 146.700 138.600 153.600 ;
        RECT 142.800 146.700 144.600 153.600 ;
        RECT 148.800 146.700 150.600 153.600 ;
        RECT 160.800 146.700 162.600 153.600 ;
        RECT 165.300 146.700 167.100 159.600 ;
        RECT 172.800 146.700 174.600 153.600 ;
        RECT 182.400 146.700 184.200 153.600 ;
        RECT 189.900 146.700 191.700 159.600 ;
        RECT 197.400 146.700 199.200 153.600 ;
        RECT 206.400 146.700 208.200 153.600 ;
        RECT 218.400 146.700 220.200 157.800 ;
        RECT 233.400 146.700 235.200 153.600 ;
        RECT 239.400 146.700 241.200 153.000 ;
        RECT 253.800 146.700 255.600 153.000 ;
        RECT 259.800 146.700 261.600 153.600 ;
        RECT 263.400 146.700 265.200 159.600 ;
        RECT 280.800 146.700 282.600 153.600 ;
        RECT 290.400 146.700 292.200 153.600 ;
        RECT 297.900 146.700 299.700 159.600 ;
        RECT 302.400 146.700 304.200 153.600 ;
        RECT 316.800 146.700 318.600 153.600 ;
        RECT 320.400 146.700 322.200 153.600 ;
        RECT 326.400 146.700 328.200 153.000 ;
        RECT 337.800 146.700 339.600 153.600 ;
        RECT 343.800 146.700 345.600 153.600 ;
        RECT 347.400 146.700 349.200 153.600 ;
        RECT 362.400 146.700 364.200 153.600 ;
        RECT 369.900 146.700 371.700 159.600 ;
        RECT 385.800 146.700 387.600 157.500 ;
        RECT 392.400 146.700 394.200 153.600 ;
        RECT 399.000 146.700 400.800 159.600 ;
        RECT 415.800 146.700 417.600 153.600 ;
        RECT 423.300 146.700 425.100 159.600 ;
        RECT 430.800 146.700 432.600 153.600 ;
        RECT 439.800 146.700 441.600 153.600 ;
        RECT 445.800 146.700 447.600 153.600 ;
        RECT 452.400 146.700 454.200 159.600 ;
        RECT 464.400 146.700 466.200 153.600 ;
        RECT 470.400 146.700 472.200 153.600 ;
        RECT 487.800 146.700 489.600 157.500 ;
        RECT 494.400 146.700 496.200 153.600 ;
        RECT 500.400 146.700 502.200 153.000 ;
        RECT 512.400 146.700 514.200 153.600 ;
        RECT 524.400 146.700 526.200 153.600 ;
        RECT 530.400 146.700 532.200 153.600 ;
        RECT 538.800 146.700 540.600 153.600 ;
        RECT 544.800 146.700 546.600 153.600 ;
        RECT 553.800 146.700 555.600 153.000 ;
        RECT 559.800 146.700 561.600 153.600 ;
        RECT 569.400 146.700 571.200 153.600 ;
        RECT 576.900 146.700 578.700 159.600 ;
        RECT 586.800 146.700 588.600 153.000 ;
        RECT 592.800 146.700 594.600 153.600 ;
        RECT 599.400 146.700 601.200 157.800 ;
        RECT 612.300 146.700 614.100 159.600 ;
        RECT 619.800 146.700 621.600 153.600 ;
        RECT 631.800 146.700 633.600 153.600 ;
        RECT 641.400 146.700 643.200 153.600 ;
        RECT 648.900 146.700 650.700 159.600 ;
        RECT 656.400 146.700 658.200 153.600 ;
        RECT 663.900 146.700 665.700 159.600 ;
        RECT 671.400 146.700 673.200 153.600 ;
        RECT 677.400 146.700 679.200 153.000 ;
        RECT 692.400 146.700 694.200 157.800 ;
        RECT 705.300 146.700 707.100 159.600 ;
        RECT 712.800 146.700 714.600 153.600 ;
        RECT 730.800 146.700 732.600 157.800 ;
        RECT 745.800 146.700 747.600 153.000 ;
        RECT 751.800 146.700 753.600 153.600 ;
        RECT -9.300 144.300 770.400 146.700 ;
        RECT -9.300 74.700 -0.300 144.300 ;
        RECT 7.800 137.400 9.600 144.300 ;
        RECT 16.800 137.400 18.600 144.300 ;
        RECT 25.800 138.000 27.600 144.300 ;
        RECT 31.800 137.400 33.600 144.300 ;
        RECT 41.400 133.200 43.200 144.300 ;
        RECT 55.800 137.400 57.600 144.300 ;
        RECT 61.800 137.400 63.600 144.300 ;
        RECT 68.400 137.400 70.200 144.300 ;
        RECT 75.900 131.400 77.700 144.300 ;
        RECT 80.400 131.400 82.200 144.300 ;
        RECT 97.800 138.000 99.600 144.300 ;
        RECT 103.800 137.400 105.600 144.300 ;
        RECT 109.800 137.400 111.600 144.300 ;
        RECT 115.800 137.400 117.600 144.300 ;
        RECT 121.800 137.400 123.600 144.300 ;
        RECT 127.800 137.400 129.600 144.300 ;
        RECT 136.800 131.400 138.600 144.300 ;
        RECT 142.800 137.400 144.600 144.300 ;
        RECT 148.800 137.400 150.600 144.300 ;
        RECT 157.800 137.400 159.600 144.300 ;
        RECT 163.800 137.400 165.600 144.300 ;
        RECT 172.800 137.400 174.600 144.300 ;
        RECT 178.800 137.400 180.600 144.300 ;
        RECT 185.400 137.400 187.200 144.300 ;
        RECT 192.900 131.400 194.700 144.300 ;
        RECT 205.200 131.400 207.000 144.300 ;
        RECT 211.800 137.400 213.600 144.300 ;
        RECT 217.800 137.400 219.600 144.300 ;
        RECT 223.800 137.400 225.600 144.300 ;
        RECT 232.800 137.400 234.600 144.300 ;
        RECT 240.300 131.400 242.100 144.300 ;
        RECT 250.800 131.400 252.600 144.300 ;
        RECT 256.800 137.400 258.600 144.300 ;
        RECT 262.800 137.400 264.600 144.300 ;
        RECT 272.400 133.200 274.200 144.300 ;
        RECT 287.400 137.400 289.200 144.300 ;
        RECT 294.900 131.400 296.700 144.300 ;
        RECT 299.400 131.400 301.200 144.300 ;
        RECT 313.800 137.400 315.600 144.300 ;
        RECT 319.800 137.400 321.600 144.300 ;
        RECT 323.400 137.400 325.200 144.300 ;
        RECT 329.400 137.400 331.200 144.300 ;
        RECT 346.800 131.400 348.600 144.300 ;
        RECT 350.400 137.400 352.200 144.300 ;
        RECT 356.400 137.400 358.200 144.300 ;
        RECT 364.800 137.400 366.600 144.300 ;
        RECT 370.800 137.400 372.600 144.300 ;
        RECT 374.400 137.400 376.200 144.300 ;
        RECT 380.400 137.400 382.200 144.300 ;
        RECT 394.800 133.200 396.600 144.300 ;
        RECT 401.400 137.400 403.200 144.300 ;
        RECT 407.400 138.000 409.200 144.300 ;
        RECT 424.800 138.000 426.600 144.300 ;
        RECT 430.800 137.400 432.600 144.300 ;
        RECT 440.400 137.400 442.200 144.300 ;
        RECT 447.900 131.400 449.700 144.300 ;
        RECT 460.800 133.200 462.600 144.300 ;
        RECT 478.800 133.200 480.600 144.300 ;
        RECT 487.800 137.400 489.600 144.300 ;
        RECT 493.800 137.400 495.600 144.300 ;
        RECT 497.400 137.400 499.200 144.300 ;
        RECT 509.400 137.400 511.200 144.300 ;
        RECT 516.900 131.400 518.700 144.300 ;
        RECT 524.400 137.400 526.200 144.300 ;
        RECT 531.900 131.400 533.700 144.300 ;
        RECT 537.300 131.400 539.100 144.300 ;
        RECT 544.800 137.400 546.600 144.300 ;
        RECT 551.400 137.400 553.200 144.300 ;
        RECT 557.400 138.000 559.200 144.300 ;
        RECT 569.400 137.400 571.200 144.300 ;
        RECT 575.400 138.000 577.200 144.300 ;
        RECT 595.800 133.500 597.600 144.300 ;
        RECT 602.400 137.400 604.200 144.300 ;
        RECT 608.400 138.000 610.200 144.300 ;
        RECT 617.400 137.400 619.200 144.300 ;
        RECT 623.400 138.000 625.200 144.300 ;
        RECT 635.400 133.200 637.200 144.300 ;
        RECT 658.800 133.200 660.600 144.300 ;
        RECT 665.400 137.400 667.200 144.300 ;
        RECT 671.400 138.000 673.200 144.300 ;
        RECT 685.800 138.000 687.600 144.300 ;
        RECT 691.800 137.400 693.600 144.300 ;
        RECT 696.300 131.400 698.100 144.300 ;
        RECT 703.800 137.400 705.600 144.300 ;
        RECT 718.800 133.200 720.600 144.300 ;
        RECT 725.400 137.400 727.200 144.300 ;
        RECT 731.400 138.000 733.200 144.300 ;
        RECT 751.800 133.200 753.600 144.300 ;
        RECT 10.800 74.700 12.600 81.000 ;
        RECT 16.800 74.700 18.600 81.600 ;
        RECT 21.300 74.700 23.100 87.600 ;
        RECT 28.800 74.700 30.600 81.600 ;
        RECT 35.400 74.700 37.200 81.600 ;
        RECT 41.400 74.700 43.200 81.000 ;
        RECT 51.300 74.700 53.100 87.600 ;
        RECT 58.800 74.700 60.600 81.600 ;
        RECT 68.400 74.700 70.200 81.600 ;
        RECT 77.400 74.700 79.200 81.600 ;
        RECT 83.400 74.700 85.200 81.000 ;
        RECT 98.400 74.700 100.200 81.600 ;
        RECT 105.900 74.700 107.700 87.600 ;
        RECT 110.400 74.700 112.200 81.600 ;
        RECT 130.800 74.700 132.600 85.800 ;
        RECT 144.300 74.700 146.100 87.450 ;
        RECT 160.800 74.700 162.600 85.800 ;
        RECT 175.800 74.700 177.600 81.000 ;
        RECT 181.800 74.700 183.600 81.600 ;
        RECT 189.300 74.700 191.100 87.600 ;
        RECT 196.800 74.700 198.600 81.600 ;
        RECT 203.400 74.700 205.200 81.600 ;
        RECT 212.400 74.700 214.200 81.600 ;
        RECT 218.400 74.700 220.200 81.600 ;
        RECT 224.400 74.700 226.200 81.600 ;
        RECT 230.400 74.700 232.200 81.000 ;
        RECT 247.800 74.700 249.600 87.600 ;
        RECT 258.300 74.700 260.100 87.450 ;
        RECT 271.800 74.700 273.600 81.000 ;
        RECT 277.800 74.700 279.600 81.600 ;
        RECT 292.800 74.700 294.600 85.800 ;
        RECT 299.400 74.700 301.200 81.600 ;
        RECT 305.400 74.700 307.200 81.000 ;
        RECT 317.400 74.700 319.200 81.600 ;
        RECT 324.900 74.700 326.700 87.600 ;
        RECT 337.800 74.700 339.600 85.800 ;
        RECT 352.200 74.700 354.000 87.600 ;
        RECT 358.800 74.700 360.600 81.600 ;
        RECT 365.400 74.700 367.200 85.500 ;
        RECT 380.400 74.700 382.200 81.600 ;
        RECT 386.400 74.700 388.200 81.000 ;
        RECT 400.800 74.700 402.600 81.000 ;
        RECT 406.800 74.700 408.600 81.600 ;
        RECT 413.400 74.700 415.200 85.800 ;
        RECT 436.800 74.700 438.600 85.500 ;
        RECT 446.400 74.700 448.200 81.600 ;
        RECT 452.400 74.700 454.200 81.000 ;
        RECT 469.800 74.700 471.600 85.800 ;
        RECT 481.800 74.700 483.600 81.600 ;
        RECT 490.800 74.700 492.600 81.000 ;
        RECT 496.800 74.700 498.600 81.600 ;
        RECT 506.400 74.700 508.200 81.600 ;
        RECT 513.900 74.700 515.700 87.600 ;
        RECT 523.800 74.700 525.600 81.000 ;
        RECT 529.800 74.700 531.600 81.600 ;
        RECT 541.800 74.700 543.600 85.800 ;
        RECT 556.800 74.700 558.600 85.800 ;
        RECT 563.400 74.700 565.200 81.600 ;
        RECT 569.400 74.700 571.200 81.000 ;
        RECT 578.400 74.700 580.200 81.600 ;
        RECT 590.400 74.700 592.200 81.600 ;
        RECT 604.800 74.700 606.600 81.600 ;
        RECT 610.800 74.700 612.600 81.600 ;
        RECT 614.400 74.700 616.200 81.600 ;
        RECT 621.000 74.700 622.800 87.600 ;
        RECT 637.800 74.700 639.600 85.800 ;
        RECT 647.400 74.700 649.200 81.600 ;
        RECT 654.900 74.700 656.700 87.600 ;
        RECT 663.300 74.700 665.100 87.600 ;
        RECT 670.800 74.700 672.600 81.600 ;
        RECT 678.300 74.700 680.100 87.600 ;
        RECT 685.800 74.700 687.600 81.600 ;
        RECT 692.400 74.700 694.200 81.600 ;
        RECT 698.400 74.700 700.200 81.000 ;
        RECT 710.400 74.700 712.200 81.600 ;
        RECT 716.400 74.700 718.200 81.000 ;
        RECT 733.800 74.700 735.600 85.800 ;
        RECT 740.400 74.700 742.200 81.600 ;
        RECT 746.400 74.700 748.200 81.000 ;
        RECT -9.300 72.300 770.400 74.700 ;
        RECT -9.300 2.700 -0.300 72.300 ;
        RECT 4.800 65.400 6.600 72.300 ;
        RECT 10.800 65.400 12.600 72.300 ;
        RECT 19.800 66.000 21.600 72.300 ;
        RECT 25.800 65.400 27.600 72.300 ;
        RECT 30.300 59.400 32.100 72.300 ;
        RECT 37.800 65.400 39.600 72.300 ;
        RECT 46.800 65.400 48.600 72.300 ;
        RECT 52.800 65.400 54.600 72.300 ;
        RECT 64.800 65.400 66.600 72.300 ;
        RECT 68.400 65.400 70.200 72.300 ;
        RECT 74.400 66.000 76.200 72.300 ;
        RECT 93.300 59.550 95.100 72.300 ;
        RECT 104.400 61.200 106.200 72.300 ;
        RECT 117.300 59.400 119.100 72.300 ;
        RECT 124.800 65.400 126.600 72.300 ;
        RECT 133.800 65.400 135.600 72.300 ;
        RECT 139.800 65.400 141.600 72.300 ;
        RECT 143.400 65.400 145.200 72.300 ;
        RECT 149.400 66.000 151.200 72.300 ;
        RECT 166.800 66.000 168.600 72.300 ;
        RECT 172.800 65.400 174.600 72.300 ;
        RECT 181.800 66.000 183.600 72.300 ;
        RECT 187.800 65.400 189.600 72.300 ;
        RECT 191.400 65.400 193.200 72.300 ;
        RECT 200.400 65.400 202.200 72.300 ;
        RECT 206.400 65.400 208.200 72.300 ;
        RECT 212.400 65.400 214.200 72.300 ;
        RECT 218.400 66.000 220.200 72.300 ;
        RECT 227.400 65.400 229.200 72.300 ;
        RECT 233.400 65.400 235.200 72.300 ;
        RECT 239.400 65.400 241.200 72.300 ;
        RECT 246.000 59.400 247.800 72.300 ;
        RECT 259.800 65.400 261.600 72.300 ;
        RECT 265.800 65.400 267.600 72.300 ;
        RECT 272.400 59.400 274.200 72.300 ;
        RECT 289.800 66.000 291.600 72.300 ;
        RECT 295.800 65.400 297.600 72.300 ;
        RECT 302.400 65.400 304.200 72.300 ;
        RECT 309.900 59.400 311.700 72.300 ;
        RECT 320.400 61.200 322.200 72.300 ;
        RECT 337.800 66.000 339.600 72.300 ;
        RECT 343.800 65.400 345.600 72.300 ;
        RECT 350.400 65.400 352.200 72.300 ;
        RECT 356.400 66.000 358.200 72.300 ;
        RECT 370.800 65.400 372.600 72.300 ;
        RECT 374.400 65.400 376.200 72.300 ;
        RECT 380.400 66.000 382.200 72.300 ;
        RECT 389.400 65.400 391.200 72.300 ;
        RECT 395.400 66.000 397.200 72.300 ;
        RECT 408.300 59.400 410.100 72.300 ;
        RECT 415.800 65.400 417.600 72.300 ;
        RECT 425.400 61.200 427.200 72.300 ;
        RECT 438.300 59.400 440.100 72.300 ;
        RECT 445.800 65.400 447.600 72.300 ;
        RECT 452.400 65.400 454.200 72.300 ;
        RECT 458.400 66.000 460.200 72.300 ;
        RECT 472.800 66.000 474.600 72.300 ;
        RECT 478.800 65.400 480.600 72.300 ;
        RECT 485.400 65.400 487.200 72.300 ;
        RECT 491.400 66.000 493.200 72.300 ;
        RECT 503.400 61.200 505.200 72.300 ;
        RECT 515.400 65.400 517.200 72.300 ;
        RECT 521.400 66.000 523.200 72.300 ;
        RECT 531.300 59.400 533.100 72.300 ;
        RECT 538.800 65.400 540.600 72.300 ;
        RECT 545.400 65.400 547.200 72.300 ;
        RECT 551.400 66.000 553.200 72.300 ;
        RECT 561.300 59.400 563.100 72.300 ;
        RECT 568.800 65.400 570.600 72.300 ;
        RECT 578.400 65.400 580.200 72.300 ;
        RECT 584.400 65.400 586.200 72.300 ;
        RECT 590.400 59.400 592.200 72.300 ;
        RECT 613.800 59.400 615.600 72.300 ;
        RECT 620.400 65.400 622.200 72.300 ;
        RECT 627.900 59.400 629.700 72.300 ;
        RECT 635.400 65.400 637.200 72.300 ;
        RECT 641.400 65.400 643.200 72.300 ;
        RECT 647.400 65.400 649.200 72.300 ;
        RECT 657.300 59.400 659.100 72.300 ;
        RECT 664.800 65.400 666.600 72.300 ;
        RECT 679.800 61.200 681.600 72.300 ;
        RECT 694.800 61.200 696.600 72.300 ;
        RECT 701.400 65.400 703.200 72.300 ;
        RECT 707.400 66.000 709.200 72.300 ;
        RECT 724.800 66.000 726.600 72.300 ;
        RECT 730.800 65.400 732.600 72.300 ;
        RECT 734.400 65.400 736.200 72.300 ;
        RECT 740.400 66.000 742.200 72.300 ;
        RECT 752.400 61.200 754.200 72.300 ;
        RECT 10.800 2.700 12.600 15.600 ;
        RECT 14.400 2.700 16.200 9.600 ;
        RECT 21.000 2.700 22.800 15.600 ;
        RECT 33.300 2.700 35.100 15.600 ;
        RECT 40.800 2.700 42.600 9.600 ;
        RECT 52.200 2.700 54.000 15.600 ;
        RECT 58.800 2.700 60.600 9.600 ;
        RECT 64.800 2.700 66.600 9.600 ;
        RECT 70.800 2.700 72.600 9.600 ;
        RECT 77.400 2.700 79.200 13.500 ;
        RECT 92.400 2.700 94.200 9.600 ;
        RECT 98.400 2.700 100.200 9.000 ;
        RECT 115.800 2.700 117.600 13.800 ;
        RECT 122.400 2.700 124.200 9.600 ;
        RECT 128.400 2.700 130.200 9.000 ;
        RECT 140.400 2.700 142.200 9.600 ;
        RECT 147.900 2.700 149.700 15.600 ;
        RECT 153.300 2.700 155.100 15.600 ;
        RECT 160.800 2.700 162.600 9.600 ;
        RECT 171.300 2.700 173.100 15.600 ;
        RECT 178.800 2.700 180.600 9.600 ;
        RECT 185.400 2.700 187.200 9.600 ;
        RECT 191.400 2.700 193.200 9.000 ;
        RECT 200.400 2.700 202.200 9.600 ;
        RECT 206.400 2.700 208.200 9.000 ;
        RECT 221.400 2.700 223.200 9.600 ;
        RECT 228.900 2.700 230.700 15.600 ;
        RECT 241.800 2.700 243.600 13.800 ;
        RECT 248.400 2.700 250.200 9.600 ;
        RECT 254.400 2.700 256.200 9.000 ;
        RECT 266.400 2.700 268.200 13.800 ;
        RECT 279.300 2.700 281.100 15.600 ;
        RECT 286.800 2.700 288.600 9.600 ;
        RECT 293.400 2.700 295.200 9.600 ;
        RECT 299.400 2.700 301.200 9.000 ;
        RECT 319.800 2.700 321.600 13.800 ;
        RECT 329.400 2.700 331.200 9.600 ;
        RECT 335.400 2.700 337.200 9.000 ;
        RECT 347.400 2.700 349.200 9.600 ;
        RECT 354.900 2.700 356.700 15.600 ;
        RECT 360.300 2.700 362.100 15.600 ;
        RECT 367.800 2.700 369.600 9.600 ;
        RECT 377.400 2.700 379.200 12.600 ;
        RECT 405.300 2.700 407.100 15.600 ;
        RECT 412.800 2.700 414.600 9.600 ;
        RECT 430.800 2.700 432.600 13.800 ;
        RECT 442.200 2.700 444.000 15.600 ;
        RECT 448.800 2.700 450.600 9.600 ;
        RECT 466.800 2.700 468.600 13.500 ;
        RECT 473.400 2.700 475.200 9.600 ;
        RECT 479.400 2.700 481.200 9.600 ;
        RECT 488.400 2.700 490.200 9.600 ;
        RECT 495.900 2.700 497.700 15.600 ;
        RECT 505.200 2.700 507.000 15.600 ;
        RECT 511.800 2.700 513.600 9.600 ;
        RECT 526.800 2.700 528.600 15.600 ;
        RECT 531.300 2.700 533.100 15.600 ;
        RECT 538.800 2.700 540.600 9.600 ;
        RECT 548.400 2.700 550.200 9.600 ;
        RECT 557.400 2.700 559.200 9.600 ;
        RECT 563.400 2.700 565.200 9.000 ;
        RECT 579.300 2.700 581.100 15.450 ;
        RECT 589.800 2.700 591.600 9.600 ;
        RECT 595.800 2.700 597.600 9.600 ;
        RECT 601.800 2.700 603.600 9.600 ;
        RECT 607.800 2.700 609.600 9.600 ;
        RECT 616.800 2.700 618.600 9.000 ;
        RECT 622.800 2.700 624.600 9.600 ;
        RECT 626.400 2.700 628.200 9.600 ;
        RECT 632.400 2.700 634.200 9.000 ;
        RECT 641.400 2.700 643.200 9.600 ;
        RECT 647.400 2.700 649.200 9.600 ;
        RECT 658.800 2.700 660.600 9.000 ;
        RECT 664.800 2.700 666.600 9.600 ;
        RECT 671.400 2.700 673.200 9.600 ;
        RECT 683.400 2.700 685.200 9.600 ;
        RECT 689.400 2.700 691.200 9.000 ;
        RECT 698.400 2.700 700.200 9.600 ;
        RECT 704.400 2.700 706.200 9.600 ;
        RECT 711.300 2.700 713.100 15.600 ;
        RECT 718.800 2.700 720.600 9.600 ;
        RECT 728.400 2.700 730.200 9.600 ;
        RECT 735.900 2.700 737.700 15.600 ;
        RECT 741.300 2.700 743.100 15.600 ;
        RECT 748.800 2.700 750.600 9.600 ;
        RECT -9.300 0.300 770.400 2.700 ;
      LAYER metal2 ;
        RECT 664.500 715.950 666.600 718.050 ;
        RECT 751.500 715.950 753.600 718.050 ;
        RECT 665.400 702.450 666.450 715.950 ;
        RECT 667.950 702.450 670.050 703.050 ;
        RECT 665.400 701.400 670.050 702.450 ;
        RECT 752.400 702.450 753.450 715.950 ;
        RECT 754.950 702.450 757.050 703.050 ;
        RECT 752.400 701.400 757.050 702.450 ;
        RECT 667.950 700.950 670.050 701.400 ;
        RECT 754.950 700.950 757.050 701.400 ;
        RECT 676.950 664.950 679.050 667.050 ;
        RECT 677.400 649.050 678.450 664.950 ;
        RECT 676.950 646.950 679.050 649.050 ;
    END
  END vdd
  PIN ABCmd_i[7]
    PORT
      LAYER metal1 ;
        RECT 205.950 552.450 208.050 553.050 ;
        RECT 211.950 552.450 214.050 553.050 ;
        RECT 205.950 551.550 214.050 552.450 ;
        RECT 205.950 550.950 208.050 551.550 ;
        RECT 211.950 550.950 214.050 551.550 ;
      LAYER metal2 ;
        RECT 482.400 728.400 489.450 729.450 ;
        RECT 488.400 667.050 489.450 728.400 ;
        RECT 478.950 664.950 481.050 667.050 ;
        RECT 487.950 664.950 490.050 667.050 ;
        RECT 479.400 621.450 480.450 664.950 ;
        RECT 479.400 620.400 483.450 621.450 ;
        RECT 482.400 592.050 483.450 620.400 ;
        RECT 466.950 589.950 469.050 592.050 ;
        RECT 481.950 589.950 484.050 592.050 ;
        RECT 313.950 556.950 316.050 559.050 ;
        RECT 205.950 553.950 208.050 556.050 ;
        RECT 206.400 553.050 207.450 553.950 ;
        RECT 205.950 550.950 208.050 553.050 ;
        RECT 211.950 552.450 214.050 553.050 ;
        RECT 211.950 551.400 216.450 552.450 ;
        RECT 211.950 550.950 214.050 551.400 ;
        RECT 215.400 535.050 216.450 551.400 ;
        RECT 232.950 550.950 235.050 553.050 ;
        RECT 331.950 550.950 334.050 553.050 ;
        RECT 233.400 535.050 234.450 550.950 ;
        RECT 214.950 532.950 217.050 535.050 ;
        RECT 232.950 532.950 235.050 535.050 ;
        RECT 233.400 529.050 234.450 532.950 ;
        RECT 232.950 526.950 235.050 529.050 ;
        RECT 332.400 508.050 333.450 550.950 ;
        RECT 331.950 505.950 334.050 508.050 ;
        RECT 385.950 505.950 388.050 508.050 ;
        RECT 332.400 463.050 333.450 505.950 ;
        RECT 386.400 486.450 387.450 505.950 ;
        RECT 467.400 504.450 468.450 589.950 ;
        RECT 467.400 503.400 471.450 504.450 ;
        RECT 388.950 486.450 391.050 487.050 ;
        RECT 386.400 485.400 391.050 486.450 ;
        RECT 388.950 484.950 391.050 485.400 ;
        RECT 265.950 460.950 268.050 463.050 ;
        RECT 304.950 460.950 307.050 463.050 ;
        RECT 331.950 460.950 334.050 463.050 ;
        RECT 266.400 457.050 267.450 460.950 ;
        RECT 265.950 454.950 268.050 457.050 ;
        RECT 305.400 427.050 306.450 460.950 ;
        RECT 389.400 427.050 390.450 484.950 ;
        RECT 470.400 460.050 471.450 503.400 ;
        RECT 493.950 484.950 496.050 487.050 ;
        RECT 494.400 460.050 495.450 484.950 ;
        RECT 451.950 457.950 454.050 460.050 ;
        RECT 469.950 457.950 472.050 460.050 ;
        RECT 493.950 457.950 496.050 460.050 ;
        RECT 452.400 444.450 453.450 457.950 ;
        RECT 452.400 443.400 456.450 444.450 ;
        RECT 455.400 427.050 456.450 443.400 ;
        RECT 280.950 424.950 283.050 427.050 ;
        RECT 304.950 424.950 307.050 427.050 ;
        RECT 388.950 424.950 391.050 427.050 ;
        RECT 397.950 424.950 400.050 427.050 ;
        RECT 454.950 424.950 457.050 427.050 ;
        RECT 148.950 400.950 151.050 403.050 ;
        RECT 163.950 400.950 166.050 403.050 ;
        RECT 214.950 400.950 217.050 403.050 ;
        RECT 149.400 388.050 150.450 400.950 ;
        RECT 148.950 385.950 151.050 388.050 ;
        RECT 164.400 343.050 165.450 400.950 ;
        RECT 215.400 391.050 216.450 400.950 ;
        RECT 281.400 391.050 282.450 424.950 ;
        RECT 305.400 418.050 306.450 424.950 ;
        RECT 304.950 415.950 307.050 418.050 ;
        RECT 398.400 415.050 399.450 424.950 ;
        RECT 331.950 412.950 334.050 415.050 ;
        RECT 397.950 412.950 400.050 415.050 ;
        RECT 214.950 388.950 217.050 391.050 ;
        RECT 229.950 388.950 232.050 391.050 ;
        RECT 280.950 388.950 283.050 391.050 ;
        RECT 298.950 388.950 301.050 391.050 ;
        RECT 215.400 382.050 216.450 388.950 ;
        RECT 230.400 382.050 231.450 388.950 ;
        RECT 214.950 379.950 217.050 382.050 ;
        RECT 229.950 379.950 232.050 382.050 ;
        RECT 299.400 343.050 300.450 388.950 ;
        RECT 455.400 382.050 456.450 424.950 ;
        RECT 454.950 379.950 457.050 382.050 ;
        RECT 157.950 340.950 160.050 343.050 ;
        RECT 163.950 340.950 166.050 343.050 ;
        RECT 298.950 340.950 301.050 343.050 ;
        RECT 307.950 340.950 310.050 343.050 ;
      LAYER metal3 ;
        RECT 478.950 666.600 481.050 667.050 ;
        RECT 487.950 666.600 490.050 667.050 ;
        RECT 478.950 665.400 490.050 666.600 ;
        RECT 478.950 664.950 481.050 665.400 ;
        RECT 487.950 664.950 490.050 665.400 ;
        RECT 466.950 591.600 469.050 592.050 ;
        RECT 481.950 591.600 484.050 592.050 ;
        RECT 466.950 590.400 484.050 591.600 ;
        RECT 466.950 589.950 469.050 590.400 ;
        RECT 481.950 589.950 484.050 590.400 ;
        RECT 313.950 558.600 316.050 559.050 ;
        RECT 308.400 557.400 316.050 558.600 ;
        RECT 232.950 552.600 235.050 553.050 ;
        RECT 308.400 552.600 309.600 557.400 ;
        RECT 313.950 556.950 316.050 557.400 ;
        RECT 331.950 552.600 334.050 553.050 ;
        RECT 232.950 551.400 334.050 552.600 ;
        RECT 232.950 550.950 235.050 551.400 ;
        RECT 331.950 550.950 334.050 551.400 ;
        RECT 214.950 534.600 217.050 535.050 ;
        RECT 232.950 534.600 235.050 535.050 ;
        RECT 214.950 533.400 235.050 534.600 ;
        RECT 214.950 532.950 217.050 533.400 ;
        RECT 232.950 532.950 235.050 533.400 ;
        RECT 331.950 507.600 334.050 508.050 ;
        RECT 385.950 507.600 388.050 508.050 ;
        RECT 331.950 506.400 388.050 507.600 ;
        RECT 331.950 505.950 334.050 506.400 ;
        RECT 385.950 505.950 388.050 506.400 ;
        RECT 265.950 462.600 268.050 463.050 ;
        RECT 304.950 462.600 307.050 463.050 ;
        RECT 331.950 462.600 334.050 463.050 ;
        RECT 265.950 461.400 334.050 462.600 ;
        RECT 265.950 460.950 268.050 461.400 ;
        RECT 304.950 460.950 307.050 461.400 ;
        RECT 331.950 460.950 334.050 461.400 ;
        RECT 451.950 459.600 454.050 460.050 ;
        RECT 469.950 459.600 472.050 460.050 ;
        RECT 493.950 459.600 496.050 460.050 ;
        RECT 451.950 458.400 496.050 459.600 ;
        RECT 451.950 457.950 454.050 458.400 ;
        RECT 469.950 457.950 472.050 458.400 ;
        RECT 493.950 457.950 496.050 458.400 ;
        RECT 280.950 426.600 283.050 427.050 ;
        RECT 304.950 426.600 307.050 427.050 ;
        RECT 280.950 425.400 307.050 426.600 ;
        RECT 280.950 424.950 283.050 425.400 ;
        RECT 304.950 424.950 307.050 425.400 ;
        RECT 388.950 426.600 391.050 427.050 ;
        RECT 397.950 426.600 400.050 427.050 ;
        RECT 454.950 426.600 457.050 427.050 ;
        RECT 388.950 425.400 457.050 426.600 ;
        RECT 388.950 424.950 391.050 425.400 ;
        RECT 397.950 424.950 400.050 425.400 ;
        RECT 454.950 424.950 457.050 425.400 ;
        RECT 304.950 417.600 307.050 418.050 ;
        RECT 304.950 416.400 333.600 417.600 ;
        RECT 304.950 415.950 307.050 416.400 ;
        RECT 332.400 415.050 333.600 416.400 ;
        RECT 331.950 412.950 334.050 415.050 ;
        RECT 148.950 402.600 151.050 403.050 ;
        RECT 163.950 402.600 166.050 403.050 ;
        RECT 214.950 402.600 217.050 403.050 ;
        RECT 148.950 401.400 217.050 402.600 ;
        RECT 148.950 400.950 151.050 401.400 ;
        RECT 163.950 400.950 166.050 401.400 ;
        RECT 214.950 400.950 217.050 401.400 ;
        RECT 214.950 390.600 217.050 391.050 ;
        RECT 229.950 390.600 232.050 391.050 ;
        RECT 280.950 390.600 283.050 391.050 ;
        RECT 298.950 390.600 301.050 391.050 ;
        RECT 214.950 389.400 301.050 390.600 ;
        RECT 214.950 388.950 217.050 389.400 ;
        RECT 229.950 388.950 232.050 389.400 ;
        RECT 280.950 388.950 283.050 389.400 ;
        RECT 298.950 388.950 301.050 389.400 ;
        RECT 157.950 342.600 160.050 343.050 ;
        RECT 163.950 342.600 166.050 343.050 ;
        RECT 157.950 341.400 166.050 342.600 ;
        RECT 157.950 340.950 160.050 341.400 ;
        RECT 163.950 340.950 166.050 341.400 ;
        RECT 298.950 342.600 301.050 343.050 ;
        RECT 307.950 342.600 310.050 343.050 ;
        RECT 298.950 341.400 310.050 342.600 ;
        RECT 298.950 340.950 301.050 341.400 ;
        RECT 307.950 340.950 310.050 341.400 ;
    END
  END ABCmd_i[7]
  PIN ABCmd_i[6]
    PORT
      LAYER metal2 ;
        RECT 476.400 724.050 477.450 729.450 ;
        RECT 445.950 721.950 448.050 724.050 ;
        RECT 475.950 721.950 478.050 724.050 ;
        RECT 446.400 607.050 447.450 721.950 ;
        RECT 397.950 604.950 400.050 607.050 ;
        RECT 445.950 604.950 448.050 607.050 ;
        RECT 475.950 604.950 478.050 607.050 ;
        RECT 100.950 601.950 103.050 604.050 ;
        RECT 112.950 601.950 115.050 604.050 ;
        RECT 103.950 592.950 106.050 595.050 ;
        RECT 104.400 592.050 105.450 592.950 ;
        RECT 113.400 592.050 114.450 601.950 ;
        RECT 103.950 589.950 106.050 592.050 ;
        RECT 112.950 589.950 115.050 592.050 ;
        RECT 136.950 589.950 139.050 592.050 ;
        RECT 137.400 549.450 138.450 589.950 ;
        RECT 134.400 548.400 138.450 549.450 ;
        RECT 134.400 532.050 135.450 548.400 ;
        RECT 398.400 547.050 399.450 604.950 ;
        RECT 476.400 604.050 477.450 604.950 ;
        RECT 475.950 601.950 478.050 604.050 ;
        RECT 196.950 544.950 199.050 547.050 ;
        RECT 397.950 544.950 400.050 547.050 ;
        RECT 133.950 529.950 136.050 532.050 ;
        RECT 148.950 523.950 151.050 526.050 ;
        RECT 149.400 517.050 150.450 523.950 ;
        RECT 197.400 517.050 198.450 544.950 ;
        RECT 148.950 514.950 151.050 517.050 ;
        RECT 196.950 514.950 199.050 517.050 ;
        RECT 149.400 492.450 150.450 514.950 ;
        RECT 146.400 491.400 150.450 492.450 ;
        RECT 146.400 460.050 147.450 491.400 ;
        RECT 145.950 457.950 148.050 460.050 ;
        RECT 154.950 457.950 157.050 460.050 ;
        RECT 163.950 457.950 166.050 460.050 ;
        RECT 155.400 454.050 156.450 457.950 ;
        RECT 164.400 454.050 165.450 457.950 ;
        RECT 154.950 451.950 157.050 454.050 ;
        RECT 163.950 451.950 166.050 454.050 ;
      LAYER metal3 ;
        RECT 445.950 723.600 448.050 724.050 ;
        RECT 475.950 723.600 478.050 724.050 ;
        RECT 445.950 722.400 478.050 723.600 ;
        RECT 445.950 721.950 448.050 722.400 ;
        RECT 475.950 721.950 478.050 722.400 ;
        RECT 397.950 606.600 400.050 607.050 ;
        RECT 445.950 606.600 448.050 607.050 ;
        RECT 475.950 606.600 478.050 607.050 ;
        RECT 397.950 605.400 478.050 606.600 ;
        RECT 397.950 604.950 400.050 605.400 ;
        RECT 445.950 604.950 448.050 605.400 ;
        RECT 475.950 604.950 478.050 605.400 ;
        RECT 100.950 603.600 103.050 604.050 ;
        RECT 112.950 603.600 115.050 604.050 ;
        RECT 100.950 602.400 115.050 603.600 ;
        RECT 100.950 601.950 103.050 602.400 ;
        RECT 112.950 601.950 115.050 602.400 ;
        RECT 103.950 591.600 106.050 592.050 ;
        RECT 112.950 591.600 115.050 592.050 ;
        RECT 136.950 591.600 139.050 592.050 ;
        RECT 103.950 590.400 139.050 591.600 ;
        RECT 103.950 589.950 106.050 590.400 ;
        RECT 112.950 589.950 115.050 590.400 ;
        RECT 136.950 589.950 139.050 590.400 ;
        RECT 196.950 546.600 199.050 547.050 ;
        RECT 397.950 546.600 400.050 547.050 ;
        RECT 196.950 545.400 400.050 546.600 ;
        RECT 196.950 544.950 199.050 545.400 ;
        RECT 397.950 544.950 400.050 545.400 ;
        RECT 133.950 531.600 136.050 532.050 ;
        RECT 133.950 530.400 150.600 531.600 ;
        RECT 133.950 529.950 136.050 530.400 ;
        RECT 149.400 526.050 150.600 530.400 ;
        RECT 148.950 523.950 151.050 526.050 ;
        RECT 148.950 516.600 151.050 517.050 ;
        RECT 196.950 516.600 199.050 517.050 ;
        RECT 148.950 515.400 199.050 516.600 ;
        RECT 148.950 514.950 151.050 515.400 ;
        RECT 196.950 514.950 199.050 515.400 ;
        RECT 145.950 459.600 148.050 460.050 ;
        RECT 154.950 459.600 157.050 460.050 ;
        RECT 163.950 459.600 166.050 460.050 ;
        RECT 145.950 458.400 166.050 459.600 ;
        RECT 145.950 457.950 148.050 458.400 ;
        RECT 154.950 457.950 157.050 458.400 ;
        RECT 163.950 457.950 166.050 458.400 ;
    END
  END ABCmd_i[6]
  PIN ABCmd_i[5]
    PORT
      LAYER metal2 ;
        RECT 395.400 706.050 396.450 729.450 ;
        RECT 394.950 705.450 397.050 706.050 ;
        RECT 392.400 704.400 397.050 705.450 ;
        RECT 250.950 699.450 253.050 700.050 ;
        RECT 253.950 699.450 256.050 700.050 ;
        RECT 250.950 698.400 256.050 699.450 ;
        RECT 250.950 697.950 253.050 698.400 ;
        RECT 253.950 697.950 256.050 698.400 ;
        RECT 251.400 672.450 252.450 697.950 ;
        RECT 392.400 697.050 393.450 704.400 ;
        RECT 394.950 703.950 397.050 704.400 ;
        RECT 391.950 694.950 394.050 697.050 ;
        RECT 412.950 694.950 415.050 697.050 ;
        RECT 248.400 671.400 252.450 672.450 ;
        RECT 413.400 675.450 414.450 694.950 ;
        RECT 415.950 675.450 418.050 676.050 ;
        RECT 413.400 674.400 418.050 675.450 ;
        RECT 248.400 664.050 249.450 671.400 ;
        RECT 265.950 664.950 268.050 667.050 ;
        RECT 266.400 664.050 267.450 664.950 ;
        RECT 247.950 661.950 250.050 664.050 ;
        RECT 265.950 661.950 268.050 664.050 ;
        RECT 248.400 637.050 249.450 661.950 ;
        RECT 413.400 640.050 414.450 674.400 ;
        RECT 415.950 673.950 418.050 674.400 ;
        RECT 277.950 637.950 280.050 640.050 ;
        RECT 412.950 637.950 415.050 640.050 ;
        RECT 226.950 634.950 229.050 637.050 ;
        RECT 241.950 634.950 244.050 637.050 ;
        RECT 247.950 634.950 250.050 637.050 ;
        RECT 160.950 592.950 163.050 595.050 ;
        RECT 184.950 592.950 187.050 595.050 ;
        RECT 161.400 592.050 162.450 592.950 ;
        RECT 185.400 592.050 186.450 592.950 ;
        RECT 160.950 589.950 163.050 592.050 ;
        RECT 184.950 589.950 187.050 592.050 ;
        RECT 185.400 589.050 186.450 589.950 ;
        RECT 227.400 589.050 228.450 634.950 ;
        RECT 242.400 634.050 243.450 634.950 ;
        RECT 278.400 634.050 279.450 637.950 ;
        RECT 241.950 631.950 244.050 634.050 ;
        RECT 277.950 631.950 280.050 634.050 ;
        RECT 184.950 586.950 187.050 589.050 ;
        RECT 226.950 586.950 229.050 589.050 ;
        RECT 227.400 580.050 228.450 586.950 ;
        RECT 226.950 577.950 229.050 580.050 ;
        RECT 307.950 577.950 310.050 580.050 ;
        RECT 227.400 568.050 228.450 577.950 ;
        RECT 220.950 565.950 223.050 568.050 ;
        RECT 226.950 565.950 229.050 568.050 ;
        RECT 221.400 562.050 222.450 565.950 ;
        RECT 220.950 559.950 223.050 562.050 ;
        RECT 308.400 559.050 309.450 577.950 ;
        RECT 307.950 556.950 310.050 559.050 ;
      LAYER metal3 ;
        RECT 391.950 696.600 394.050 697.050 ;
        RECT 412.950 696.600 415.050 697.050 ;
        RECT 391.950 695.400 415.050 696.600 ;
        RECT 391.950 694.950 394.050 695.400 ;
        RECT 412.950 694.950 415.050 695.400 ;
        RECT 247.950 663.600 250.050 664.050 ;
        RECT 265.950 663.600 268.050 664.050 ;
        RECT 247.950 662.400 268.050 663.600 ;
        RECT 247.950 661.950 250.050 662.400 ;
        RECT 265.950 661.950 268.050 662.400 ;
        RECT 277.950 639.600 280.050 640.050 ;
        RECT 412.950 639.600 415.050 640.050 ;
        RECT 277.950 638.400 415.050 639.600 ;
        RECT 277.950 637.950 280.050 638.400 ;
        RECT 412.950 637.950 415.050 638.400 ;
        RECT 226.950 636.600 229.050 637.050 ;
        RECT 241.950 636.600 244.050 637.050 ;
        RECT 247.950 636.600 250.050 637.050 ;
        RECT 226.950 635.400 250.050 636.600 ;
        RECT 226.950 634.950 229.050 635.400 ;
        RECT 241.950 634.950 244.050 635.400 ;
        RECT 247.950 634.950 250.050 635.400 ;
        RECT 241.950 633.600 244.050 634.050 ;
        RECT 277.950 633.600 280.050 634.050 ;
        RECT 241.950 632.400 280.050 633.600 ;
        RECT 241.950 631.950 244.050 632.400 ;
        RECT 277.950 631.950 280.050 632.400 ;
        RECT 160.950 591.600 163.050 592.050 ;
        RECT 184.950 591.600 187.050 592.050 ;
        RECT 160.950 590.400 187.050 591.600 ;
        RECT 160.950 589.950 163.050 590.400 ;
        RECT 184.950 589.950 187.050 590.400 ;
        RECT 184.950 588.600 187.050 589.050 ;
        RECT 226.950 588.600 229.050 589.050 ;
        RECT 184.950 587.400 229.050 588.600 ;
        RECT 184.950 586.950 187.050 587.400 ;
        RECT 226.950 586.950 229.050 587.400 ;
        RECT 226.950 579.600 229.050 580.050 ;
        RECT 307.950 579.600 310.050 580.050 ;
        RECT 226.950 578.400 310.050 579.600 ;
        RECT 226.950 577.950 229.050 578.400 ;
        RECT 307.950 577.950 310.050 578.400 ;
        RECT 220.950 567.600 223.050 568.050 ;
        RECT 226.950 567.600 229.050 568.050 ;
        RECT 220.950 566.400 229.050 567.600 ;
        RECT 220.950 565.950 223.050 566.400 ;
        RECT 226.950 565.950 229.050 566.400 ;
    END
  END ABCmd_i[5]
  PIN ABCmd_i[4]
    PORT
      LAYER metal2 ;
        RECT 365.400 724.050 366.450 729.450 ;
        RECT 286.950 721.950 289.050 724.050 ;
        RECT 364.950 721.950 367.050 724.050 ;
        RECT 283.950 702.450 286.050 703.050 ;
        RECT 287.400 702.450 288.450 721.950 ;
        RECT 283.950 701.400 288.450 702.450 ;
        RECT 283.950 700.950 286.050 701.400 ;
        RECT 287.400 691.050 288.450 701.400 ;
        RECT 286.950 688.950 289.050 691.050 ;
        RECT 313.950 688.950 316.050 691.050 ;
        RECT 314.400 670.050 315.450 688.950 ;
        RECT 313.950 667.950 316.050 670.050 ;
        RECT 310.950 661.950 313.050 664.050 ;
        RECT 367.950 661.950 370.050 664.050 ;
        RECT 311.400 634.050 312.450 661.950 ;
        RECT 283.950 631.950 286.050 634.050 ;
        RECT 310.950 631.950 313.050 634.050 ;
        RECT 368.400 604.050 369.450 661.950 ;
        RECT 367.950 601.950 370.050 604.050 ;
      LAYER metal3 ;
        RECT 286.950 723.600 289.050 724.050 ;
        RECT 364.950 723.600 367.050 724.050 ;
        RECT 286.950 722.400 367.050 723.600 ;
        RECT 286.950 721.950 289.050 722.400 ;
        RECT 364.950 721.950 367.050 722.400 ;
        RECT 286.950 690.600 289.050 691.050 ;
        RECT 313.950 690.600 316.050 691.050 ;
        RECT 286.950 689.400 316.050 690.600 ;
        RECT 286.950 688.950 289.050 689.400 ;
        RECT 313.950 688.950 316.050 689.400 ;
        RECT 313.950 669.600 316.050 670.050 ;
        RECT 313.950 668.400 318.600 669.600 ;
        RECT 313.950 667.950 316.050 668.400 ;
        RECT 310.950 663.600 313.050 664.050 ;
        RECT 317.400 663.600 318.600 668.400 ;
        RECT 367.950 663.600 370.050 664.050 ;
        RECT 310.950 662.400 370.050 663.600 ;
        RECT 310.950 661.950 313.050 662.400 ;
        RECT 367.950 661.950 370.050 662.400 ;
        RECT 283.950 633.600 286.050 634.050 ;
        RECT 310.950 633.600 313.050 634.050 ;
        RECT 283.950 632.400 313.050 633.600 ;
        RECT 283.950 631.950 286.050 632.400 ;
        RECT 310.950 631.950 313.050 632.400 ;
    END
  END ABCmd_i[4]
  PIN ABCmd_i[3]
    PORT
      LAYER metal2 ;
        RECT 341.400 728.400 345.450 729.450 ;
        RECT 344.400 709.050 345.450 728.400 ;
        RECT 343.950 706.950 346.050 709.050 ;
        RECT 406.950 706.950 409.050 709.050 ;
        RECT 344.400 703.050 345.450 706.950 ;
        RECT 343.950 700.950 346.050 703.050 ;
        RECT 407.400 696.450 408.450 706.950 ;
        RECT 409.950 696.450 412.050 697.050 ;
        RECT 407.400 695.400 412.050 696.450 ;
        RECT 409.950 694.950 412.050 695.400 ;
      LAYER metal3 ;
        RECT 343.950 708.600 346.050 709.050 ;
        RECT 406.950 708.600 409.050 709.050 ;
        RECT 343.950 707.400 409.050 708.600 ;
        RECT 343.950 706.950 346.050 707.400 ;
        RECT 406.950 706.950 409.050 707.400 ;
    END
  END ABCmd_i[3]
  PIN ABCmd_i[2]
    PORT
      LAYER metal2 ;
        RECT 769.950 700.950 772.050 703.050 ;
        RECT 154.950 699.450 157.050 700.050 ;
        RECT 154.950 698.400 159.450 699.450 ;
        RECT 154.950 697.950 157.050 698.400 ;
        RECT 158.400 652.050 159.450 698.400 ;
        RECT 430.950 697.950 433.050 700.050 ;
        RECT 431.400 697.050 432.450 697.950 ;
        RECT 424.950 694.950 427.050 697.050 ;
        RECT 430.950 694.950 433.050 697.050 ;
        RECT 425.400 688.050 426.450 694.950 ;
        RECT 770.400 688.050 771.450 700.950 ;
        RECT 424.950 685.950 427.050 688.050 ;
        RECT 769.950 685.950 772.050 688.050 ;
        RECT 425.400 655.050 426.450 685.950 ;
        RECT 424.950 652.950 427.050 655.050 ;
        RECT 130.950 649.950 133.050 652.050 ;
        RECT 157.950 649.950 160.050 652.050 ;
        RECT 131.400 631.050 132.450 649.950 ;
        RECT 130.950 628.950 133.050 631.050 ;
        RECT 139.950 625.950 142.050 628.050 ;
        RECT 140.400 601.050 141.450 625.950 ;
        RECT 133.950 598.950 136.050 601.050 ;
        RECT 139.950 598.950 142.050 601.050 ;
      LAYER metal3 ;
        RECT 769.950 702.600 772.050 703.050 ;
        RECT 769.950 701.400 777.600 702.600 ;
        RECT 769.950 700.950 772.050 701.400 ;
        RECT 424.950 696.600 427.050 697.050 ;
        RECT 430.950 696.600 433.050 697.050 ;
        RECT 424.950 695.400 433.050 696.600 ;
        RECT 424.950 694.950 427.050 695.400 ;
        RECT 430.950 694.950 433.050 695.400 ;
        RECT 424.950 687.600 427.050 688.050 ;
        RECT 769.950 687.600 772.050 688.050 ;
        RECT 424.950 686.400 772.050 687.600 ;
        RECT 424.950 685.950 427.050 686.400 ;
        RECT 769.950 685.950 772.050 686.400 ;
        RECT 424.950 654.600 427.050 655.050 ;
        RECT 377.400 653.400 427.050 654.600 ;
        RECT 130.950 651.600 133.050 652.050 ;
        RECT 157.950 651.600 160.050 652.050 ;
        RECT 377.400 651.600 378.600 653.400 ;
        RECT 424.950 652.950 427.050 653.400 ;
        RECT 130.950 650.400 378.600 651.600 ;
        RECT 130.950 649.950 133.050 650.400 ;
        RECT 157.950 649.950 160.050 650.400 ;
        RECT 130.950 628.950 133.050 631.050 ;
        RECT 131.400 627.600 132.600 628.950 ;
        RECT 139.950 627.600 142.050 628.050 ;
        RECT 131.400 626.400 142.050 627.600 ;
        RECT 139.950 625.950 142.050 626.400 ;
        RECT 133.950 600.600 136.050 601.050 ;
        RECT 139.950 600.600 142.050 601.050 ;
        RECT 133.950 599.400 142.050 600.600 ;
        RECT 133.950 598.950 136.050 599.400 ;
        RECT 139.950 598.950 142.050 599.400 ;
    END
  END ABCmd_i[2]
  PIN ABCmd_i[1]
    PORT
      LAYER metal2 ;
        RECT 403.950 700.950 406.050 703.050 ;
        RECT 427.950 700.950 430.050 703.050 ;
        RECT 404.400 672.450 405.450 700.950 ;
        RECT 619.950 682.950 622.050 685.050 ;
        RECT 401.400 671.400 405.450 672.450 ;
        RECT 401.400 667.050 402.450 671.400 ;
        RECT 400.950 664.950 403.050 667.050 ;
        RECT 409.950 664.950 412.050 667.050 ;
        RECT 401.400 646.050 402.450 664.950 ;
        RECT 620.400 646.050 621.450 682.950 ;
        RECT 400.950 643.950 403.050 646.050 ;
        RECT 619.950 643.950 622.050 646.050 ;
        RECT 349.950 625.950 352.050 628.050 ;
        RECT 350.400 625.050 351.450 625.950 ;
        RECT 401.400 625.050 402.450 643.950 ;
        RECT 349.950 622.950 352.050 625.050 ;
        RECT 400.950 622.950 403.050 625.050 ;
        RECT 620.400 609.450 621.450 643.950 ;
        RECT 617.400 608.400 621.450 609.450 ;
        RECT 617.400 604.050 618.450 608.400 ;
        RECT 616.950 601.950 619.050 604.050 ;
      LAYER metal3 ;
        RECT 403.950 702.600 406.050 703.050 ;
        RECT 427.950 702.600 430.050 703.050 ;
        RECT 403.950 701.400 430.050 702.600 ;
        RECT 403.950 700.950 406.050 701.400 ;
        RECT 427.950 700.950 430.050 701.400 ;
        RECT 619.950 684.600 622.050 685.050 ;
        RECT 619.950 683.400 777.600 684.600 ;
        RECT 619.950 682.950 622.050 683.400 ;
        RECT 776.400 680.400 777.600 683.400 ;
        RECT 400.950 666.600 403.050 667.050 ;
        RECT 409.950 666.600 412.050 667.050 ;
        RECT 400.950 665.400 412.050 666.600 ;
        RECT 400.950 664.950 403.050 665.400 ;
        RECT 409.950 664.950 412.050 665.400 ;
        RECT 400.950 645.600 403.050 646.050 ;
        RECT 619.950 645.600 622.050 646.050 ;
        RECT 400.950 644.400 622.050 645.600 ;
        RECT 400.950 643.950 403.050 644.400 ;
        RECT 619.950 643.950 622.050 644.400 ;
        RECT 349.950 624.600 352.050 625.050 ;
        RECT 400.950 624.600 403.050 625.050 ;
        RECT 349.950 623.400 403.050 624.600 ;
        RECT 349.950 622.950 352.050 623.400 ;
        RECT 400.950 622.950 403.050 623.400 ;
    END
  END ABCmd_i[1]
  PIN ABCmd_i[0]
    PORT
      LAYER metal2 ;
        RECT 340.950 703.950 343.050 706.050 ;
        RECT 346.950 703.950 349.050 706.050 ;
        RECT 341.400 694.050 342.450 703.950 ;
        RECT 340.950 691.950 343.050 694.050 ;
        RECT 379.950 691.950 382.050 694.050 ;
        RECT 526.950 691.950 529.050 694.050 ;
        RECT 766.950 691.950 769.050 694.050 ;
        RECT 380.400 673.050 381.450 691.950 ;
        RECT 527.400 676.050 528.450 691.950 ;
        RECT 767.400 676.050 768.450 691.950 ;
        RECT 526.950 673.950 529.050 676.050 ;
        RECT 766.950 673.950 769.050 676.050 ;
        RECT 379.950 672.450 382.050 673.050 ;
        RECT 377.400 671.400 382.050 672.450 ;
        RECT 377.400 646.050 378.450 671.400 ;
        RECT 379.950 670.950 382.050 671.400 ;
        RECT 295.950 643.950 298.050 646.050 ;
        RECT 313.950 643.950 316.050 646.050 ;
        RECT 337.950 643.950 340.050 646.050 ;
        RECT 376.950 643.950 379.050 646.050 ;
        RECT 296.400 631.050 297.450 643.950 ;
        RECT 295.950 628.950 298.050 631.050 ;
        RECT 310.950 627.450 313.050 628.050 ;
        RECT 314.400 627.450 315.450 643.950 ;
        RECT 338.400 631.050 339.450 643.950 ;
        RECT 337.950 628.950 340.050 631.050 ;
        RECT 310.950 626.400 315.450 627.450 ;
        RECT 310.950 625.950 313.050 626.400 ;
        RECT 311.400 606.450 312.450 625.950 ;
        RECT 308.400 605.400 312.450 606.450 ;
        RECT 308.400 601.050 309.450 605.400 ;
        RECT 307.950 598.950 310.050 601.050 ;
      LAYER metal3 ;
        RECT 340.950 705.600 343.050 706.050 ;
        RECT 346.950 705.600 349.050 706.050 ;
        RECT 340.950 704.400 349.050 705.600 ;
        RECT 340.950 703.950 343.050 704.400 ;
        RECT 346.950 703.950 349.050 704.400 ;
        RECT 340.950 693.600 343.050 694.050 ;
        RECT 379.950 693.600 382.050 694.050 ;
        RECT 340.950 692.400 382.050 693.600 ;
        RECT 340.950 691.950 343.050 692.400 ;
        RECT 379.950 691.950 382.050 692.400 ;
        RECT 526.950 693.600 529.050 694.050 ;
        RECT 766.950 693.600 769.050 694.050 ;
        RECT 526.950 692.400 769.050 693.600 ;
        RECT 526.950 691.950 529.050 692.400 ;
        RECT 766.950 691.950 769.050 692.400 ;
        RECT 526.950 675.600 529.050 676.050 ;
        RECT 485.400 674.400 529.050 675.600 ;
        RECT 379.950 672.600 382.050 673.050 ;
        RECT 485.400 672.600 486.600 674.400 ;
        RECT 526.950 673.950 529.050 674.400 ;
        RECT 766.950 675.600 769.050 676.050 ;
        RECT 766.950 674.400 777.600 675.600 ;
        RECT 766.950 673.950 769.050 674.400 ;
        RECT 379.950 671.400 486.600 672.600 ;
        RECT 379.950 670.950 382.050 671.400 ;
        RECT 295.950 645.600 298.050 646.050 ;
        RECT 313.950 645.600 316.050 646.050 ;
        RECT 337.950 645.600 340.050 646.050 ;
        RECT 376.950 645.600 379.050 646.050 ;
        RECT 295.950 644.400 379.050 645.600 ;
        RECT 295.950 643.950 298.050 644.400 ;
        RECT 313.950 643.950 316.050 644.400 ;
        RECT 337.950 643.950 340.050 644.400 ;
        RECT 376.950 643.950 379.050 644.400 ;
    END
  END ABCmd_i[0]
  PIN ACC_o[7]
    PORT
      LAYER metal2 ;
        RECT 373.950 265.950 376.050 268.050 ;
        RECT 391.950 265.950 394.050 268.050 ;
        RECT 374.400 253.050 375.450 265.950 ;
        RECT 349.950 250.950 352.050 253.050 ;
        RECT 373.950 250.950 376.050 253.050 ;
        RECT 350.400 217.050 351.450 250.950 ;
        RECT 337.950 214.950 340.050 217.050 ;
        RECT 349.950 214.950 352.050 217.050 ;
        RECT 338.400 172.050 339.450 214.950 ;
        RECT 322.950 169.950 325.050 172.050 ;
        RECT 337.950 169.950 340.050 172.050 ;
        RECT 323.400 166.050 324.450 169.950 ;
        RECT 322.950 163.950 325.050 166.050 ;
        RECT 301.950 157.950 304.050 160.050 ;
        RECT 302.400 127.050 303.450 157.950 ;
        RECT 301.950 124.950 304.050 127.050 ;
        RECT 313.950 121.950 316.050 124.050 ;
        RECT 314.400 102.450 315.450 121.950 ;
        RECT 311.400 101.400 315.450 102.450 ;
        RECT 311.400 64.050 312.450 101.400 ;
        RECT 310.950 61.950 313.050 64.050 ;
        RECT 346.950 61.950 349.050 64.050 ;
        RECT 347.400 30.450 348.450 61.950 ;
        RECT 344.400 29.400 348.450 30.450 ;
        RECT 344.400 4.050 345.450 29.400 ;
        RECT 343.950 1.950 346.050 4.050 ;
        RECT 388.950 1.950 391.050 4.050 ;
        RECT 389.400 -3.600 390.450 1.950 ;
      LAYER metal3 ;
        RECT 373.950 267.600 376.050 268.050 ;
        RECT 391.950 267.600 394.050 268.050 ;
        RECT 373.950 266.400 394.050 267.600 ;
        RECT 373.950 265.950 376.050 266.400 ;
        RECT 391.950 265.950 394.050 266.400 ;
        RECT 349.950 252.600 352.050 253.050 ;
        RECT 373.950 252.600 376.050 253.050 ;
        RECT 349.950 251.400 376.050 252.600 ;
        RECT 349.950 250.950 352.050 251.400 ;
        RECT 373.950 250.950 376.050 251.400 ;
        RECT 337.950 216.600 340.050 217.050 ;
        RECT 349.950 216.600 352.050 217.050 ;
        RECT 337.950 215.400 352.050 216.600 ;
        RECT 337.950 214.950 340.050 215.400 ;
        RECT 349.950 214.950 352.050 215.400 ;
        RECT 322.950 171.600 325.050 172.050 ;
        RECT 337.950 171.600 340.050 172.050 ;
        RECT 322.950 170.400 340.050 171.600 ;
        RECT 322.950 169.950 325.050 170.400 ;
        RECT 337.950 169.950 340.050 170.400 ;
        RECT 322.950 165.600 325.050 166.050 ;
        RECT 322.950 164.400 327.600 165.600 ;
        RECT 322.950 163.950 325.050 164.400 ;
        RECT 301.950 159.600 304.050 160.050 ;
        RECT 326.400 159.600 327.600 164.400 ;
        RECT 301.950 158.400 327.600 159.600 ;
        RECT 301.950 157.950 304.050 158.400 ;
        RECT 301.950 126.600 304.050 127.050 ;
        RECT 301.950 125.400 315.600 126.600 ;
        RECT 301.950 124.950 304.050 125.400 ;
        RECT 314.400 124.050 315.600 125.400 ;
        RECT 313.950 121.950 316.050 124.050 ;
        RECT 310.950 63.600 313.050 64.050 ;
        RECT 346.950 63.600 349.050 64.050 ;
        RECT 310.950 62.400 349.050 63.600 ;
        RECT 310.950 61.950 313.050 62.400 ;
        RECT 346.950 61.950 349.050 62.400 ;
        RECT 343.950 3.600 346.050 4.050 ;
        RECT 388.950 3.600 391.050 4.050 ;
        RECT 343.950 2.400 391.050 3.600 ;
        RECT 343.950 1.950 346.050 2.400 ;
        RECT 388.950 1.950 391.050 2.400 ;
    END
  END ACC_o[7]
  PIN ACC_o[6]
    PORT
      LAYER metal2 ;
        RECT 337.950 312.450 340.050 313.050 ;
        RECT 335.400 311.400 340.050 312.450 ;
        RECT 335.400 277.050 336.450 311.400 ;
        RECT 337.950 310.950 340.050 311.400 ;
        RECT 307.950 274.950 310.050 277.050 ;
        RECT 334.950 274.950 337.050 277.050 ;
        RECT 308.400 244.050 309.450 274.950 ;
        RECT 307.950 241.950 310.050 244.050 ;
        RECT 313.950 241.950 316.050 244.050 ;
        RECT 314.400 210.450 315.450 241.950 ;
        RECT 314.400 209.400 318.450 210.450 ;
        RECT 317.400 202.050 318.450 209.400 ;
        RECT 316.950 199.950 319.050 202.050 ;
        RECT 313.950 193.950 316.050 196.050 ;
        RECT 314.400 171.450 315.450 193.950 ;
        RECT 311.400 170.400 315.450 171.450 ;
        RECT 311.400 136.050 312.450 170.400 ;
        RECT 310.950 133.950 313.050 136.050 ;
        RECT 334.950 133.950 337.050 136.050 ;
        RECT 335.400 100.050 336.450 133.950 ;
        RECT 313.950 97.950 316.050 100.050 ;
        RECT 334.950 97.950 337.050 100.050 ;
        RECT 314.400 61.050 315.450 97.950 ;
        RECT 313.950 58.950 316.050 61.050 ;
        RECT 361.950 58.950 364.050 61.050 ;
        RECT 362.400 34.050 363.450 58.950 ;
        RECT 361.950 31.950 364.050 34.050 ;
        RECT 394.950 31.950 397.050 34.050 ;
        RECT 395.400 -3.600 396.450 31.950 ;
      LAYER metal3 ;
        RECT 307.950 276.600 310.050 277.050 ;
        RECT 334.950 276.600 337.050 277.050 ;
        RECT 307.950 275.400 337.050 276.600 ;
        RECT 307.950 274.950 310.050 275.400 ;
        RECT 334.950 274.950 337.050 275.400 ;
        RECT 307.950 243.600 310.050 244.050 ;
        RECT 313.950 243.600 316.050 244.050 ;
        RECT 307.950 242.400 316.050 243.600 ;
        RECT 307.950 241.950 310.050 242.400 ;
        RECT 313.950 241.950 316.050 242.400 ;
        RECT 316.950 201.600 319.050 202.050 ;
        RECT 314.400 200.400 319.050 201.600 ;
        RECT 314.400 196.050 315.600 200.400 ;
        RECT 316.950 199.950 319.050 200.400 ;
        RECT 313.950 193.950 316.050 196.050 ;
        RECT 310.950 135.600 313.050 136.050 ;
        RECT 334.950 135.600 337.050 136.050 ;
        RECT 310.950 134.400 337.050 135.600 ;
        RECT 310.950 133.950 313.050 134.400 ;
        RECT 334.950 133.950 337.050 134.400 ;
        RECT 313.950 99.600 316.050 100.050 ;
        RECT 334.950 99.600 337.050 100.050 ;
        RECT 313.950 98.400 337.050 99.600 ;
        RECT 313.950 97.950 316.050 98.400 ;
        RECT 334.950 97.950 337.050 98.400 ;
        RECT 313.950 60.600 316.050 61.050 ;
        RECT 361.950 60.600 364.050 61.050 ;
        RECT 313.950 59.400 364.050 60.600 ;
        RECT 313.950 58.950 316.050 59.400 ;
        RECT 361.950 58.950 364.050 59.400 ;
        RECT 361.950 33.600 364.050 34.050 ;
        RECT 394.950 33.600 397.050 34.050 ;
        RECT 361.950 32.400 397.050 33.600 ;
        RECT 361.950 31.950 364.050 32.400 ;
        RECT 394.950 31.950 397.050 32.400 ;
    END
  END ACC_o[6]
  PIN ACC_o[5]
    PORT
      LAYER metal2 ;
        RECT 394.950 310.950 397.050 313.050 ;
        RECT 403.950 310.950 406.050 313.050 ;
        RECT 404.400 280.050 405.450 310.950 ;
        RECT 403.950 277.950 406.050 280.050 ;
        RECT 418.950 277.950 421.050 280.050 ;
        RECT 419.400 253.050 420.450 277.950 ;
        RECT 403.950 250.950 406.050 253.050 ;
        RECT 418.950 250.950 421.050 253.050 ;
        RECT 404.400 241.050 405.450 250.950 ;
        RECT 403.950 238.950 406.050 241.050 ;
        RECT 394.950 229.950 397.050 232.050 ;
        RECT 395.400 193.050 396.450 229.950 ;
        RECT 394.950 190.950 397.050 193.050 ;
        RECT 406.950 190.950 409.050 193.050 ;
        RECT 407.400 139.050 408.450 190.950 ;
        RECT 394.950 136.950 397.050 139.050 ;
        RECT 406.950 136.950 409.050 139.050 ;
        RECT 395.400 127.050 396.450 136.950 ;
        RECT 394.950 124.950 397.050 127.050 ;
        RECT 403.950 124.950 406.050 127.050 ;
        RECT 404.400 102.450 405.450 124.950 ;
        RECT 404.400 101.400 408.450 102.450 ;
        RECT 407.400 97.050 408.450 101.400 ;
        RECT 406.950 94.950 409.050 97.050 ;
        RECT 418.950 88.950 421.050 91.050 ;
        RECT 419.400 73.050 420.450 88.950 ;
        RECT 403.950 70.950 406.050 73.050 ;
        RECT 418.950 70.950 421.050 73.050 ;
        RECT 404.400 34.050 405.450 70.950 ;
        RECT 397.950 31.950 400.050 34.050 ;
        RECT 403.950 31.950 406.050 34.050 ;
        RECT 398.400 -2.550 399.450 31.950 ;
        RECT 398.400 -3.600 402.450 -2.550 ;
      LAYER metal3 ;
        RECT 394.950 312.600 397.050 313.050 ;
        RECT 403.950 312.600 406.050 313.050 ;
        RECT 394.950 311.400 406.050 312.600 ;
        RECT 394.950 310.950 397.050 311.400 ;
        RECT 403.950 310.950 406.050 311.400 ;
        RECT 403.950 279.600 406.050 280.050 ;
        RECT 418.950 279.600 421.050 280.050 ;
        RECT 403.950 278.400 421.050 279.600 ;
        RECT 403.950 277.950 406.050 278.400 ;
        RECT 418.950 277.950 421.050 278.400 ;
        RECT 403.950 252.600 406.050 253.050 ;
        RECT 418.950 252.600 421.050 253.050 ;
        RECT 403.950 251.400 421.050 252.600 ;
        RECT 403.950 250.950 406.050 251.400 ;
        RECT 418.950 250.950 421.050 251.400 ;
        RECT 403.950 240.600 406.050 241.050 ;
        RECT 398.400 239.400 406.050 240.600 ;
        RECT 398.400 234.600 399.600 239.400 ;
        RECT 403.950 238.950 406.050 239.400 ;
        RECT 395.400 233.400 399.600 234.600 ;
        RECT 395.400 232.050 396.600 233.400 ;
        RECT 394.950 229.950 397.050 232.050 ;
        RECT 394.950 192.600 397.050 193.050 ;
        RECT 406.950 192.600 409.050 193.050 ;
        RECT 394.950 191.400 409.050 192.600 ;
        RECT 394.950 190.950 397.050 191.400 ;
        RECT 406.950 190.950 409.050 191.400 ;
        RECT 394.950 138.600 397.050 139.050 ;
        RECT 406.950 138.600 409.050 139.050 ;
        RECT 394.950 137.400 409.050 138.600 ;
        RECT 394.950 136.950 397.050 137.400 ;
        RECT 406.950 136.950 409.050 137.400 ;
        RECT 394.950 126.600 397.050 127.050 ;
        RECT 403.950 126.600 406.050 127.050 ;
        RECT 394.950 125.400 406.050 126.600 ;
        RECT 394.950 124.950 397.050 125.400 ;
        RECT 403.950 124.950 406.050 125.400 ;
        RECT 406.950 96.600 409.050 97.050 ;
        RECT 406.950 95.400 420.600 96.600 ;
        RECT 406.950 94.950 409.050 95.400 ;
        RECT 419.400 91.050 420.600 95.400 ;
        RECT 418.950 88.950 421.050 91.050 ;
        RECT 403.950 72.600 406.050 73.050 ;
        RECT 418.950 72.600 421.050 73.050 ;
        RECT 403.950 71.400 421.050 72.600 ;
        RECT 403.950 70.950 406.050 71.400 ;
        RECT 418.950 70.950 421.050 71.400 ;
        RECT 397.950 33.600 400.050 34.050 ;
        RECT 403.950 33.600 406.050 34.050 ;
        RECT 397.950 32.400 406.050 33.600 ;
        RECT 397.950 31.950 400.050 32.400 ;
        RECT 403.950 31.950 406.050 32.400 ;
    END
  END ACC_o[5]
  PIN ACC_o[4]
    PORT
      LAYER metal1 ;
        RECT 148.950 171.450 151.050 172.050 ;
        RECT 148.950 170.550 153.450 171.450 ;
        RECT 148.950 169.950 151.050 170.550 ;
        RECT 152.550 163.050 153.450 170.550 ;
        RECT 151.950 160.950 154.050 163.050 ;
      LAYER metal2 ;
        RECT 373.950 316.950 376.050 319.050 ;
        RECT 406.950 316.950 409.050 319.050 ;
        RECT 374.400 295.050 375.450 316.950 ;
        RECT 407.400 313.050 408.450 316.950 ;
        RECT 406.950 310.950 409.050 313.050 ;
        RECT 358.950 292.950 361.050 295.050 ;
        RECT 373.950 292.950 376.050 295.050 ;
        RECT 359.400 280.050 360.450 292.950 ;
        RECT 253.950 277.950 256.050 280.050 ;
        RECT 358.950 277.950 361.050 280.050 ;
        RECT 254.400 253.050 255.450 277.950 ;
        RECT 196.950 250.950 199.050 253.050 ;
        RECT 253.950 250.950 256.050 253.050 ;
        RECT 197.400 205.050 198.450 250.950 ;
        RECT 163.950 202.950 166.050 205.050 ;
        RECT 196.950 202.950 199.050 205.050 ;
        RECT 164.400 175.050 165.450 202.950 ;
        RECT 148.950 172.950 151.050 175.050 ;
        RECT 163.950 172.950 166.050 175.050 ;
        RECT 149.400 172.050 150.450 172.950 ;
        RECT 148.950 169.950 151.050 172.050 ;
        RECT 151.950 160.950 154.050 163.050 ;
        RECT 152.400 106.050 153.450 160.950 ;
        RECT 136.950 103.950 139.050 106.050 ;
        RECT 151.950 103.950 154.050 106.050 ;
        RECT 137.400 73.050 138.450 103.950 ;
        RECT 136.950 70.950 139.050 73.050 ;
        RECT 283.950 70.950 286.050 73.050 ;
        RECT 284.400 37.050 285.450 70.950 ;
        RECT 283.950 34.950 286.050 37.050 ;
        RECT 310.950 34.950 313.050 37.050 ;
        RECT 311.400 7.050 312.450 34.950 ;
        RECT 310.950 4.950 313.050 7.050 ;
        RECT 406.950 4.950 409.050 7.050 ;
        RECT 407.400 -3.600 408.450 4.950 ;
      LAYER metal3 ;
        RECT 373.950 318.600 376.050 319.050 ;
        RECT 406.950 318.600 409.050 319.050 ;
        RECT 373.950 317.400 409.050 318.600 ;
        RECT 373.950 316.950 376.050 317.400 ;
        RECT 406.950 316.950 409.050 317.400 ;
        RECT 358.950 294.600 361.050 295.050 ;
        RECT 373.950 294.600 376.050 295.050 ;
        RECT 358.950 293.400 376.050 294.600 ;
        RECT 358.950 292.950 361.050 293.400 ;
        RECT 373.950 292.950 376.050 293.400 ;
        RECT 253.950 279.600 256.050 280.050 ;
        RECT 358.950 279.600 361.050 280.050 ;
        RECT 253.950 278.400 361.050 279.600 ;
        RECT 253.950 277.950 256.050 278.400 ;
        RECT 358.950 277.950 361.050 278.400 ;
        RECT 196.950 252.600 199.050 253.050 ;
        RECT 253.950 252.600 256.050 253.050 ;
        RECT 196.950 251.400 256.050 252.600 ;
        RECT 196.950 250.950 199.050 251.400 ;
        RECT 253.950 250.950 256.050 251.400 ;
        RECT 163.950 204.600 166.050 205.050 ;
        RECT 196.950 204.600 199.050 205.050 ;
        RECT 163.950 203.400 199.050 204.600 ;
        RECT 163.950 202.950 166.050 203.400 ;
        RECT 196.950 202.950 199.050 203.400 ;
        RECT 148.950 174.600 151.050 175.050 ;
        RECT 163.950 174.600 166.050 175.050 ;
        RECT 148.950 173.400 166.050 174.600 ;
        RECT 148.950 172.950 151.050 173.400 ;
        RECT 163.950 172.950 166.050 173.400 ;
        RECT 136.950 105.600 139.050 106.050 ;
        RECT 151.950 105.600 154.050 106.050 ;
        RECT 136.950 104.400 154.050 105.600 ;
        RECT 136.950 103.950 139.050 104.400 ;
        RECT 151.950 103.950 154.050 104.400 ;
        RECT 136.950 72.600 139.050 73.050 ;
        RECT 283.950 72.600 286.050 73.050 ;
        RECT 136.950 71.400 286.050 72.600 ;
        RECT 136.950 70.950 139.050 71.400 ;
        RECT 283.950 70.950 286.050 71.400 ;
        RECT 283.950 36.600 286.050 37.050 ;
        RECT 310.950 36.600 313.050 37.050 ;
        RECT 283.950 35.400 313.050 36.600 ;
        RECT 283.950 34.950 286.050 35.400 ;
        RECT 310.950 34.950 313.050 35.400 ;
        RECT 310.950 6.600 313.050 7.050 ;
        RECT 406.950 6.600 409.050 7.050 ;
        RECT 310.950 5.400 409.050 6.600 ;
        RECT 310.950 4.950 313.050 5.400 ;
        RECT 406.950 4.950 409.050 5.400 ;
    END
  END ACC_o[4]
  PIN ACC_o[3]
    PORT
      LAYER metal2 ;
        RECT 262.950 433.950 265.050 436.050 ;
        RECT 424.950 433.950 427.050 436.050 ;
        RECT 263.400 397.050 264.450 433.950 ;
        RECT 425.400 412.050 426.450 433.950 ;
        RECT 424.950 409.950 427.050 412.050 ;
        RECT 433.950 409.950 436.050 412.050 ;
        RECT 124.950 394.950 127.050 397.050 ;
        RECT 262.950 394.950 265.050 397.050 ;
        RECT 125.400 346.050 126.450 394.950 ;
        RECT 109.950 343.950 112.050 346.050 ;
        RECT 124.950 343.950 127.050 346.050 ;
        RECT 110.400 280.050 111.450 343.950 ;
        RECT 70.950 277.950 73.050 280.050 ;
        RECT 109.950 277.950 112.050 280.050 ;
        RECT 71.400 256.050 72.450 277.950 ;
        RECT 46.950 253.950 49.050 256.050 ;
        RECT 70.950 253.950 73.050 256.050 ;
        RECT 47.400 205.050 48.450 253.950 ;
        RECT 46.950 202.950 49.050 205.050 ;
        RECT 55.950 202.950 58.050 205.050 ;
        RECT 56.400 172.050 57.450 202.950 ;
        RECT 55.950 169.950 58.050 172.050 ;
        RECT 130.950 169.950 133.050 172.050 ;
        RECT 131.400 109.050 132.450 169.950 ;
        RECT 130.950 106.950 133.050 109.050 ;
        RECT 208.950 106.950 211.050 109.050 ;
        RECT 209.400 67.050 210.450 106.950 ;
        RECT 208.950 64.950 211.050 67.050 ;
        RECT 400.950 64.950 403.050 67.050 ;
        RECT 401.400 4.050 402.450 64.950 ;
        RECT 400.950 1.950 403.050 4.050 ;
        RECT 430.950 1.950 433.050 4.050 ;
        RECT 431.400 -3.600 432.450 1.950 ;
      LAYER metal3 ;
        RECT 262.950 435.600 265.050 436.050 ;
        RECT 424.950 435.600 427.050 436.050 ;
        RECT 262.950 434.400 427.050 435.600 ;
        RECT 262.950 433.950 265.050 434.400 ;
        RECT 424.950 433.950 427.050 434.400 ;
        RECT 424.950 411.600 427.050 412.050 ;
        RECT 433.950 411.600 436.050 412.050 ;
        RECT 424.950 410.400 436.050 411.600 ;
        RECT 424.950 409.950 427.050 410.400 ;
        RECT 433.950 409.950 436.050 410.400 ;
        RECT 124.950 396.600 127.050 397.050 ;
        RECT 262.950 396.600 265.050 397.050 ;
        RECT 124.950 395.400 265.050 396.600 ;
        RECT 124.950 394.950 127.050 395.400 ;
        RECT 262.950 394.950 265.050 395.400 ;
        RECT 109.950 345.600 112.050 346.050 ;
        RECT 124.950 345.600 127.050 346.050 ;
        RECT 109.950 344.400 127.050 345.600 ;
        RECT 109.950 343.950 112.050 344.400 ;
        RECT 124.950 343.950 127.050 344.400 ;
        RECT 70.950 279.600 73.050 280.050 ;
        RECT 109.950 279.600 112.050 280.050 ;
        RECT 70.950 278.400 112.050 279.600 ;
        RECT 70.950 277.950 73.050 278.400 ;
        RECT 109.950 277.950 112.050 278.400 ;
        RECT 46.950 255.600 49.050 256.050 ;
        RECT 70.950 255.600 73.050 256.050 ;
        RECT 46.950 254.400 73.050 255.600 ;
        RECT 46.950 253.950 49.050 254.400 ;
        RECT 70.950 253.950 73.050 254.400 ;
        RECT 46.950 204.600 49.050 205.050 ;
        RECT 55.950 204.600 58.050 205.050 ;
        RECT 46.950 203.400 58.050 204.600 ;
        RECT 46.950 202.950 49.050 203.400 ;
        RECT 55.950 202.950 58.050 203.400 ;
        RECT 55.950 171.600 58.050 172.050 ;
        RECT 130.950 171.600 133.050 172.050 ;
        RECT 55.950 170.400 133.050 171.600 ;
        RECT 55.950 169.950 58.050 170.400 ;
        RECT 130.950 169.950 133.050 170.400 ;
        RECT 130.950 108.600 133.050 109.050 ;
        RECT 208.950 108.600 211.050 109.050 ;
        RECT 130.950 107.400 211.050 108.600 ;
        RECT 130.950 106.950 133.050 107.400 ;
        RECT 208.950 106.950 211.050 107.400 ;
        RECT 208.950 66.600 211.050 67.050 ;
        RECT 400.950 66.600 403.050 67.050 ;
        RECT 208.950 65.400 403.050 66.600 ;
        RECT 208.950 64.950 211.050 65.400 ;
        RECT 400.950 64.950 403.050 65.400 ;
        RECT 400.950 3.600 403.050 4.050 ;
        RECT 430.950 3.600 433.050 4.050 ;
        RECT 400.950 2.400 433.050 3.600 ;
        RECT 400.950 1.950 403.050 2.400 ;
        RECT 430.950 1.950 433.050 2.400 ;
    END
  END ACC_o[3]
  PIN ACC_o[2]
    PORT
      LAYER metal2 ;
        RECT 112.950 586.950 115.050 589.050 ;
        RECT 113.400 574.050 114.450 586.950 ;
        RECT 526.950 583.950 529.050 586.050 ;
        RECT 1.950 571.950 4.050 574.050 ;
        RECT 112.950 571.950 115.050 574.050 ;
        RECT 2.400 559.050 3.450 571.950 ;
        RECT 1.950 556.950 4.050 559.050 ;
        RECT 523.950 555.450 526.050 556.050 ;
        RECT 527.400 555.450 528.450 583.950 ;
        RECT 523.950 554.400 528.450 555.450 ;
        RECT 523.950 553.950 526.050 554.400 ;
      LAYER metal3 ;
        RECT 112.950 588.600 115.050 589.050 ;
        RECT 112.950 587.400 168.600 588.600 ;
        RECT 112.950 586.950 115.050 587.400 ;
        RECT 167.400 585.600 168.600 587.400 ;
        RECT 251.400 587.400 291.600 588.600 ;
        RECT 251.400 585.600 252.600 587.400 ;
        RECT 167.400 584.400 252.600 585.600 ;
        RECT 290.400 585.600 291.600 587.400 ;
        RECT 526.950 585.600 529.050 586.050 ;
        RECT 290.400 584.400 529.050 585.600 ;
        RECT 526.950 583.950 529.050 584.400 ;
        RECT 1.950 573.600 4.050 574.050 ;
        RECT 112.950 573.600 115.050 574.050 ;
        RECT 1.950 572.400 115.050 573.600 ;
        RECT 1.950 571.950 4.050 572.400 ;
        RECT 112.950 571.950 115.050 572.400 ;
        RECT 1.950 558.600 4.050 559.050 ;
        RECT -3.600 557.400 4.050 558.600 ;
        RECT 1.950 556.950 4.050 557.400 ;
    END
  END ACC_o[2]
  PIN ACC_o[1]
    PORT
      LAYER metal2 ;
        RECT 7.950 562.950 10.050 565.050 ;
        RECT 8.400 529.050 9.450 562.950 ;
        RECT 7.950 526.950 10.050 529.050 ;
      LAYER metal3 ;
        RECT 7.950 564.600 10.050 565.050 ;
        RECT -3.600 563.400 10.050 564.600 ;
        RECT 7.950 562.950 10.050 563.400 ;
    END
  END ACC_o[1]
  PIN ACC_o[0]
    PORT
      LAYER metal2 ;
        RECT 4.950 568.950 7.050 571.050 ;
        RECT 5.400 562.050 6.450 568.950 ;
        RECT 4.950 559.950 7.050 562.050 ;
        RECT 4.950 553.950 7.050 556.050 ;
      LAYER metal3 ;
        RECT 4.950 570.600 7.050 571.050 ;
        RECT -3.600 569.400 7.050 570.600 ;
        RECT 4.950 568.950 7.050 569.400 ;
        RECT 4.950 559.950 7.050 562.050 ;
        RECT 5.400 556.050 6.600 559.950 ;
        RECT 4.950 553.950 7.050 556.050 ;
    END
  END ACC_o[0]
  PIN Done_o
    PORT
      LAYER metal2 ;
        RECT 754.950 526.950 757.050 529.050 ;
        RECT 742.950 523.950 745.050 526.050 ;
        RECT 743.400 489.450 744.450 523.950 ;
        RECT 740.400 488.400 744.450 489.450 ;
        RECT 740.400 438.450 741.450 488.400 ;
        RECT 737.400 437.400 741.450 438.450 ;
        RECT 737.400 406.050 738.450 437.400 ;
        RECT 736.950 403.950 739.050 406.050 ;
        RECT 766.950 403.950 769.050 406.050 ;
        RECT 767.400 292.050 768.450 403.950 ;
        RECT 757.950 289.950 760.050 292.050 ;
        RECT 766.950 289.950 769.050 292.050 ;
        RECT 758.400 259.050 759.450 289.950 ;
        RECT 715.950 256.950 718.050 259.050 ;
        RECT 757.950 256.950 760.050 259.050 ;
        RECT 716.400 235.050 717.450 256.950 ;
        RECT 709.950 232.950 712.050 235.050 ;
        RECT 715.950 232.950 718.050 235.050 ;
        RECT 710.400 205.050 711.450 232.950 ;
        RECT 709.950 202.950 712.050 205.050 ;
        RECT 718.950 190.950 721.050 193.050 ;
        RECT 719.400 142.050 720.450 190.950 ;
        RECT 718.950 139.950 721.050 142.050 ;
        RECT 766.950 139.950 769.050 142.050 ;
        RECT 767.400 4.050 768.450 139.950 ;
        RECT 754.950 1.950 757.050 4.050 ;
        RECT 766.950 1.950 769.050 4.050 ;
        RECT 755.400 -3.600 756.450 1.950 ;
      LAYER metal3 ;
        RECT 754.950 528.600 757.050 529.050 ;
        RECT 743.400 527.400 757.050 528.600 ;
        RECT 743.400 526.050 744.600 527.400 ;
        RECT 754.950 526.950 757.050 527.400 ;
        RECT 742.950 523.950 745.050 526.050 ;
        RECT 736.950 405.600 739.050 406.050 ;
        RECT 766.950 405.600 769.050 406.050 ;
        RECT 736.950 404.400 769.050 405.600 ;
        RECT 736.950 403.950 739.050 404.400 ;
        RECT 766.950 403.950 769.050 404.400 ;
        RECT 757.950 291.600 760.050 292.050 ;
        RECT 766.950 291.600 769.050 292.050 ;
        RECT 757.950 290.400 769.050 291.600 ;
        RECT 757.950 289.950 760.050 290.400 ;
        RECT 766.950 289.950 769.050 290.400 ;
        RECT 715.950 258.600 718.050 259.050 ;
        RECT 757.950 258.600 760.050 259.050 ;
        RECT 715.950 257.400 760.050 258.600 ;
        RECT 715.950 256.950 718.050 257.400 ;
        RECT 757.950 256.950 760.050 257.400 ;
        RECT 709.950 234.600 712.050 235.050 ;
        RECT 715.950 234.600 718.050 235.050 ;
        RECT 709.950 233.400 718.050 234.600 ;
        RECT 709.950 232.950 712.050 233.400 ;
        RECT 715.950 232.950 718.050 233.400 ;
        RECT 709.950 204.600 712.050 205.050 ;
        RECT 709.950 203.400 720.600 204.600 ;
        RECT 709.950 202.950 712.050 203.400 ;
        RECT 719.400 193.050 720.600 203.400 ;
        RECT 718.950 190.950 721.050 193.050 ;
        RECT 718.950 141.600 721.050 142.050 ;
        RECT 766.950 141.600 769.050 142.050 ;
        RECT 718.950 140.400 769.050 141.600 ;
        RECT 718.950 139.950 721.050 140.400 ;
        RECT 766.950 139.950 769.050 140.400 ;
        RECT 754.950 3.600 757.050 4.050 ;
        RECT 766.950 3.600 769.050 4.050 ;
        RECT 754.950 2.400 769.050 3.600 ;
        RECT 754.950 1.950 757.050 2.400 ;
        RECT 766.950 1.950 769.050 2.400 ;
    END
  END Done_o
  PIN LoadA_i
    PORT
      LAYER metal2 ;
        RECT 713.400 637.050 714.450 729.450 ;
        RECT 712.950 634.950 715.050 637.050 ;
        RECT 688.950 625.950 691.050 628.050 ;
        RECT 689.400 610.050 690.450 625.950 ;
        RECT 721.950 622.950 724.050 625.050 ;
        RECT 688.950 607.950 691.050 610.050 ;
        RECT 694.950 607.950 697.050 610.050 ;
        RECT 695.400 604.050 696.450 607.950 ;
        RECT 722.400 604.050 723.450 622.950 ;
        RECT 694.950 601.950 697.050 604.050 ;
        RECT 721.950 601.950 724.050 604.050 ;
        RECT 722.400 601.050 723.450 601.950 ;
        RECT 721.950 598.950 724.050 601.050 ;
      LAYER metal3 ;
        RECT 712.950 636.600 715.050 637.050 ;
        RECT 712.950 635.400 720.600 636.600 ;
        RECT 712.950 634.950 715.050 635.400 ;
        RECT 719.400 624.600 720.600 635.400 ;
        RECT 721.950 624.600 724.050 625.050 ;
        RECT 719.400 623.400 724.050 624.600 ;
        RECT 721.950 622.950 724.050 623.400 ;
        RECT 688.950 609.600 691.050 610.050 ;
        RECT 694.950 609.600 697.050 610.050 ;
        RECT 688.950 608.400 697.050 609.600 ;
        RECT 688.950 607.950 691.050 608.400 ;
        RECT 694.950 607.950 697.050 608.400 ;
        RECT 694.950 603.600 697.050 604.050 ;
        RECT 721.950 603.600 724.050 604.050 ;
        RECT 694.950 602.400 724.050 603.600 ;
        RECT 694.950 601.950 697.050 602.400 ;
        RECT 721.950 601.950 724.050 602.400 ;
    END
  END LoadA_i
  PIN LoadB_i
    PORT
      LAYER metal2 ;
        RECT 719.400 724.050 720.450 729.450 ;
        RECT 700.950 721.950 703.050 724.050 ;
        RECT 718.950 721.950 721.050 724.050 ;
        RECT 701.400 670.050 702.450 721.950 ;
        RECT 700.950 669.450 703.050 670.050 ;
        RECT 698.400 668.400 703.050 669.450 ;
        RECT 698.400 640.050 699.450 668.400 ;
        RECT 700.950 667.950 703.050 668.400 ;
        RECT 685.950 637.950 688.050 640.050 ;
        RECT 697.950 637.950 700.050 640.050 ;
        RECT 686.400 631.050 687.450 637.950 ;
        RECT 685.950 628.950 688.050 631.050 ;
        RECT 697.950 622.950 700.050 625.050 ;
        RECT 698.400 607.050 699.450 622.950 ;
        RECT 697.950 604.950 700.050 607.050 ;
        RECT 709.950 604.950 712.050 607.050 ;
        RECT 698.400 601.050 699.450 604.950 ;
        RECT 710.400 604.050 711.450 604.950 ;
        RECT 709.950 601.950 712.050 604.050 ;
        RECT 697.950 598.950 700.050 601.050 ;
      LAYER metal3 ;
        RECT 700.950 723.600 703.050 724.050 ;
        RECT 718.950 723.600 721.050 724.050 ;
        RECT 700.950 722.400 721.050 723.600 ;
        RECT 700.950 721.950 703.050 722.400 ;
        RECT 718.950 721.950 721.050 722.400 ;
        RECT 685.950 639.600 688.050 640.050 ;
        RECT 697.950 639.600 700.050 640.050 ;
        RECT 685.950 638.400 700.050 639.600 ;
        RECT 685.950 637.950 688.050 638.400 ;
        RECT 697.950 637.950 700.050 638.400 ;
        RECT 685.950 630.600 688.050 631.050 ;
        RECT 685.950 629.400 699.600 630.600 ;
        RECT 685.950 628.950 688.050 629.400 ;
        RECT 698.400 625.050 699.600 629.400 ;
        RECT 697.950 622.950 700.050 625.050 ;
        RECT 697.950 606.600 700.050 607.050 ;
        RECT 709.950 606.600 712.050 607.050 ;
        RECT 697.950 605.400 712.050 606.600 ;
        RECT 697.950 604.950 700.050 605.400 ;
        RECT 709.950 604.950 712.050 605.400 ;
    END
  END LoadB_i
  PIN LoadCmd_i
    PORT
      LAYER metal2 ;
        RECT 740.400 728.400 744.450 729.450 ;
        RECT 740.400 676.050 741.450 728.400 ;
        RECT 724.950 673.950 727.050 676.050 ;
        RECT 739.950 673.950 742.050 676.050 ;
        RECT 745.950 673.950 748.050 676.050 ;
        RECT 725.400 673.050 726.450 673.950 ;
        RECT 724.950 670.950 727.050 673.050 ;
      LAYER metal3 ;
        RECT 724.950 675.600 727.050 676.050 ;
        RECT 739.950 675.600 742.050 676.050 ;
        RECT 745.950 675.600 748.050 676.050 ;
        RECT 724.950 674.400 748.050 675.600 ;
        RECT 724.950 673.950 727.050 674.400 ;
        RECT 739.950 673.950 742.050 674.400 ;
        RECT 745.950 673.950 748.050 674.400 ;
    END
  END LoadCmd_i
  PIN clk
    PORT
      LAYER metal2 ;
        RECT 602.400 709.050 603.450 729.450 ;
        RECT 496.950 706.950 499.050 709.050 ;
        RECT 505.950 706.950 508.050 709.050 ;
        RECT 580.950 706.950 583.050 709.050 ;
        RECT 601.950 706.950 604.050 709.050 ;
        RECT 497.400 594.450 498.450 706.950 ;
        RECT 506.400 703.050 507.450 706.950 ;
        RECT 581.400 703.050 582.450 706.950 ;
        RECT 505.950 700.950 508.050 703.050 ;
        RECT 580.950 700.950 583.050 703.050 ;
        RECT 497.400 593.400 501.450 594.450 ;
        RECT 500.400 520.050 501.450 593.400 ;
        RECT 700.950 523.950 703.050 526.050 ;
        RECT 499.950 517.950 502.050 520.050 ;
        RECT 571.950 517.950 574.050 520.050 ;
        RECT 500.400 514.050 501.450 517.950 ;
        RECT 484.950 511.950 487.050 514.050 ;
        RECT 499.950 511.950 502.050 514.050 ;
        RECT 485.400 487.050 486.450 511.950 ;
        RECT 572.400 508.050 573.450 517.950 ;
        RECT 701.400 508.050 702.450 523.950 ;
        RECT 571.950 505.950 574.050 508.050 ;
        RECT 700.950 505.950 703.050 508.050 ;
        RECT 484.950 486.450 487.050 487.050 ;
        RECT 482.400 485.400 487.050 486.450 ;
        RECT 482.400 469.050 483.450 485.400 ;
        RECT 484.950 484.950 487.050 485.400 ;
        RECT 448.950 466.950 451.050 469.050 ;
        RECT 481.950 466.950 484.050 469.050 ;
        RECT 449.400 454.050 450.450 466.950 ;
        RECT 448.950 451.950 451.050 454.050 ;
        RECT 457.950 451.950 460.050 454.050 ;
      LAYER metal3 ;
        RECT 496.950 708.600 499.050 709.050 ;
        RECT 505.950 708.600 508.050 709.050 ;
        RECT 580.950 708.600 583.050 709.050 ;
        RECT 601.950 708.600 604.050 709.050 ;
        RECT 496.950 707.400 604.050 708.600 ;
        RECT 496.950 706.950 499.050 707.400 ;
        RECT 505.950 706.950 508.050 707.400 ;
        RECT 580.950 706.950 583.050 707.400 ;
        RECT 601.950 706.950 604.050 707.400 ;
        RECT 499.950 519.600 502.050 520.050 ;
        RECT 571.950 519.600 574.050 520.050 ;
        RECT 499.950 518.400 574.050 519.600 ;
        RECT 499.950 517.950 502.050 518.400 ;
        RECT 571.950 517.950 574.050 518.400 ;
        RECT 484.950 513.600 487.050 514.050 ;
        RECT 499.950 513.600 502.050 514.050 ;
        RECT 484.950 512.400 502.050 513.600 ;
        RECT 484.950 511.950 487.050 512.400 ;
        RECT 499.950 511.950 502.050 512.400 ;
        RECT 571.950 507.600 574.050 508.050 ;
        RECT 700.950 507.600 703.050 508.050 ;
        RECT 571.950 506.400 703.050 507.600 ;
        RECT 571.950 505.950 574.050 506.400 ;
        RECT 700.950 505.950 703.050 506.400 ;
        RECT 448.950 468.600 451.050 469.050 ;
        RECT 481.950 468.600 484.050 469.050 ;
        RECT 448.950 467.400 484.050 468.600 ;
        RECT 448.950 466.950 451.050 467.400 ;
        RECT 481.950 466.950 484.050 467.400 ;
        RECT 448.950 453.600 451.050 454.050 ;
        RECT 457.950 453.600 460.050 454.050 ;
        RECT 448.950 452.400 460.050 453.600 ;
        RECT 448.950 451.950 451.050 452.400 ;
        RECT 457.950 451.950 460.050 452.400 ;
    END
  END clk
  PIN reset
    PORT
      LAYER metal2 ;
        RECT 758.400 709.050 759.450 729.450 ;
        RECT 757.950 706.950 760.050 709.050 ;
        RECT 754.950 697.950 757.050 700.050 ;
        RECT 755.400 676.050 756.450 697.950 ;
        RECT 754.950 673.950 757.050 676.050 ;
      LAYER metal3 ;
        RECT 757.950 706.950 760.050 709.050 ;
        RECT 754.950 699.600 757.050 700.050 ;
        RECT 758.400 699.600 759.600 706.950 ;
        RECT 754.950 698.400 759.600 699.600 ;
        RECT 754.950 697.950 757.050 698.400 ;
    END
  END reset
  OBS
      LAYER metal1 ;
        RECT 9.300 708.900 11.100 718.200 ;
        RECT 9.000 708.000 11.100 708.900 ;
        RECT 16.800 712.200 18.600 718.200 ;
        RECT 5.100 702.150 6.900 703.950 ;
        RECT 4.950 700.050 7.050 702.150 ;
        RECT 9.000 700.950 9.900 708.000 ;
        RECT 16.800 707.100 17.700 712.200 ;
        RECT 29.700 707.400 31.500 719.400 ;
        RECT 40.800 713.400 42.600 719.400 ;
        RECT 11.550 706.200 17.700 707.100 ;
        RECT 11.550 703.500 12.750 706.200 ;
        RECT 26.250 705.150 28.050 706.950 ;
        RECT 10.950 701.700 12.750 703.500 ;
        RECT 14.100 702.150 15.900 703.950 ;
        RECT 25.950 703.050 28.050 705.150 ;
        RECT 29.850 702.150 31.050 707.400 ;
        RECT 35.100 702.150 36.900 703.950 ;
        RECT 7.950 698.850 10.050 700.950 ;
        RECT 9.000 694.200 9.900 698.850 ;
        RECT 11.550 696.000 12.750 701.700 ;
        RECT 13.950 700.050 16.050 702.150 ;
        RECT 16.950 698.850 19.050 700.950 ;
        RECT 28.950 700.050 31.050 702.150 ;
        RECT 17.100 697.050 18.900 698.850 ;
        RECT 28.950 696.750 30.150 700.050 ;
        RECT 31.950 698.850 34.050 700.950 ;
        RECT 34.950 700.050 37.050 702.150 ;
        RECT 41.400 700.950 42.600 713.400 ;
        RECT 55.500 707.400 57.300 719.400 ;
        RECT 71.700 707.400 73.500 719.400 ;
        RECT 82.800 707.400 84.600 719.400 ;
        RECT 85.800 708.300 87.600 719.400 ;
        RECT 91.800 708.300 93.600 719.400 ;
        RECT 85.800 707.400 93.600 708.300 ;
        RECT 101.700 707.400 103.500 719.400 ;
        RECT 113.400 713.400 115.200 719.400 ;
        RECT 50.100 702.150 51.900 703.950 ;
        RECT 55.950 702.150 57.150 707.400 ;
        RECT 58.950 705.150 60.750 706.950 ;
        RECT 68.250 705.150 70.050 706.950 ;
        RECT 58.950 703.050 61.050 705.150 ;
        RECT 67.950 703.050 70.050 705.150 ;
        RECT 71.850 702.150 73.050 707.400 ;
        RECT 77.100 702.150 78.900 703.950 ;
        RECT 83.400 702.150 84.300 707.400 ;
        RECT 98.250 705.150 100.050 706.950 ;
        RECT 97.950 703.050 100.050 705.150 ;
        RECT 101.850 702.150 103.050 707.400 ;
        RECT 107.100 702.150 108.900 703.950 ;
        RECT 40.950 698.850 43.050 700.950 ;
        RECT 44.100 699.150 45.900 700.950 ;
        RECT 49.950 700.050 52.050 702.150 ;
        RECT 32.100 697.050 33.900 698.850 ;
        RECT 11.550 695.100 17.850 696.000 ;
        RECT 9.000 693.300 11.100 694.200 ;
        RECT 9.300 688.800 11.100 693.300 ;
        RECT 16.800 691.800 17.850 695.100 ;
        RECT 26.400 695.700 30.150 696.750 ;
        RECT 26.400 693.600 27.600 695.700 ;
        RECT 16.800 688.800 18.600 691.800 ;
        RECT 25.800 687.600 27.600 693.600 ;
        RECT 28.800 692.700 36.600 694.050 ;
        RECT 28.800 687.600 30.600 692.700 ;
        RECT 34.800 687.600 36.600 692.700 ;
        RECT 41.400 690.600 42.600 698.850 ;
        RECT 43.950 697.050 46.050 699.150 ;
        RECT 52.950 698.850 55.050 700.950 ;
        RECT 55.950 700.050 58.050 702.150 ;
        RECT 53.100 697.050 54.900 698.850 ;
        RECT 56.850 696.750 58.050 700.050 ;
        RECT 70.950 700.050 73.050 702.150 ;
        RECT 70.950 696.750 72.150 700.050 ;
        RECT 73.950 698.850 76.050 700.950 ;
        RECT 76.950 700.050 79.050 702.150 ;
        RECT 82.950 700.050 85.050 702.150 ;
        RECT 74.100 697.050 75.900 698.850 ;
        RECT 56.850 695.700 60.600 696.750 ;
        RECT 40.800 687.600 42.600 690.600 ;
        RECT 50.400 692.700 58.200 694.050 ;
        RECT 50.400 687.600 52.200 692.700 ;
        RECT 56.400 687.600 58.200 692.700 ;
        RECT 59.400 693.600 60.600 695.700 ;
        RECT 68.400 695.700 72.150 696.750 ;
        RECT 68.400 693.600 69.600 695.700 ;
        RECT 59.400 687.600 61.200 693.600 ;
        RECT 67.800 687.600 69.600 693.600 ;
        RECT 70.800 692.700 78.600 694.050 ;
        RECT 70.800 687.600 72.600 692.700 ;
        RECT 76.800 687.600 78.600 692.700 ;
        RECT 83.400 693.600 84.300 700.050 ;
        RECT 85.950 698.850 88.050 700.950 ;
        RECT 89.100 699.150 90.900 700.950 ;
        RECT 86.100 697.050 87.900 698.850 ;
        RECT 88.950 697.050 91.050 699.150 ;
        RECT 91.950 698.850 94.050 700.950 ;
        RECT 100.950 700.050 103.050 702.150 ;
        RECT 92.100 697.050 93.900 698.850 ;
        RECT 100.950 696.750 102.150 700.050 ;
        RECT 103.950 698.850 106.050 700.950 ;
        RECT 106.950 700.050 109.050 702.150 ;
        RECT 113.400 700.950 114.600 713.400 ;
        RECT 122.400 712.200 124.200 718.200 ;
        RECT 123.300 707.100 124.200 712.200 ;
        RECT 129.900 708.900 131.700 718.200 ;
        RECT 129.900 708.000 132.000 708.900 ;
        RECT 123.300 706.200 129.450 707.100 ;
        RECT 125.100 702.150 126.900 703.950 ;
        RECT 128.250 703.500 129.450 706.200 ;
        RECT 110.100 699.150 111.900 700.950 ;
        RECT 104.100 697.050 105.900 698.850 ;
        RECT 109.950 697.050 112.050 699.150 ;
        RECT 112.950 698.850 115.050 700.950 ;
        RECT 121.950 698.850 124.050 700.950 ;
        RECT 124.950 700.050 127.050 702.150 ;
        RECT 128.250 701.700 130.050 703.500 ;
        RECT 98.400 695.700 102.150 696.750 ;
        RECT 98.400 693.600 99.600 695.700 ;
        RECT 83.400 691.950 88.800 693.600 ;
        RECT 87.000 687.600 88.800 691.950 ;
        RECT 97.800 687.600 99.600 693.600 ;
        RECT 100.800 692.700 108.600 694.050 ;
        RECT 100.800 687.600 102.600 692.700 ;
        RECT 106.800 687.600 108.600 692.700 ;
        RECT 113.400 690.600 114.600 698.850 ;
        RECT 122.100 697.050 123.900 698.850 ;
        RECT 128.250 696.000 129.450 701.700 ;
        RECT 131.100 700.950 132.000 708.000 ;
        RECT 146.700 707.400 148.500 719.400 ;
        RECT 155.400 713.400 157.200 719.400 ;
        RECT 143.250 705.150 145.050 706.950 ;
        RECT 134.100 702.150 135.900 703.950 ;
        RECT 142.950 703.050 145.050 705.150 ;
        RECT 146.850 702.150 148.050 707.400 ;
        RECT 155.400 706.500 156.600 713.400 ;
        RECT 161.700 707.400 163.500 719.400 ;
        RECT 169.800 707.400 171.600 719.400 ;
        RECT 172.800 708.300 174.600 719.400 ;
        RECT 178.800 708.300 180.600 719.400 ;
        RECT 172.800 707.400 180.600 708.300 ;
        RECT 190.500 707.400 192.300 719.400 ;
        RECT 205.800 713.400 207.600 719.400 ;
        RECT 155.400 705.600 161.100 706.500 ;
        RECT 159.150 704.700 161.100 705.600 ;
        RECT 152.100 702.150 153.900 703.950 ;
        RECT 155.100 702.150 156.900 703.950 ;
        RECT 130.950 698.850 133.050 700.950 ;
        RECT 133.950 700.050 136.050 702.150 ;
        RECT 145.950 700.050 148.050 702.150 ;
        RECT 123.150 695.100 129.450 696.000 ;
        RECT 123.150 691.800 124.200 695.100 ;
        RECT 131.100 694.200 132.000 698.850 ;
        RECT 145.950 696.750 147.150 700.050 ;
        RECT 148.950 698.850 151.050 700.950 ;
        RECT 151.950 700.050 154.050 702.150 ;
        RECT 154.950 700.050 157.050 702.150 ;
        RECT 149.100 697.050 150.900 698.850 ;
        RECT 113.400 687.600 115.200 690.600 ;
        RECT 122.400 688.800 124.200 691.800 ;
        RECT 129.900 693.300 132.000 694.200 ;
        RECT 143.400 695.700 147.150 696.750 ;
        RECT 159.150 696.300 160.050 704.700 ;
        RECT 162.000 702.150 163.200 707.400 ;
        RECT 170.400 702.150 171.300 707.400 ;
        RECT 172.950 705.450 175.050 706.050 ;
        RECT 181.950 705.450 184.050 706.050 ;
        RECT 172.950 704.550 184.050 705.450 ;
        RECT 172.950 703.950 175.050 704.550 ;
        RECT 181.950 703.950 184.050 704.550 ;
        RECT 185.100 702.150 186.900 703.950 ;
        RECT 190.950 702.150 192.150 707.400 ;
        RECT 193.950 705.150 195.750 706.950 ;
        RECT 206.400 705.150 207.600 713.400 ;
        RECT 216.300 708.900 218.100 719.400 ;
        RECT 215.700 707.550 218.100 708.900 ;
        RECT 193.950 703.050 196.050 705.150 ;
        RECT 160.950 700.050 163.200 702.150 ;
        RECT 169.950 700.050 172.050 702.150 ;
        RECT 143.400 693.600 144.600 695.700 ;
        RECT 159.150 695.400 161.100 696.300 ;
        RECT 156.000 694.500 161.100 695.400 ;
        RECT 129.900 688.800 131.700 693.300 ;
        RECT 142.800 687.600 144.600 693.600 ;
        RECT 145.800 692.700 153.600 694.050 ;
        RECT 145.800 687.600 147.600 692.700 ;
        RECT 151.800 687.600 153.600 692.700 ;
        RECT 156.000 690.600 157.200 694.500 ;
        RECT 162.000 693.600 163.200 700.050 ;
        RECT 170.400 693.600 171.300 700.050 ;
        RECT 172.950 698.850 175.050 700.950 ;
        RECT 176.100 699.150 177.900 700.950 ;
        RECT 173.100 697.050 174.900 698.850 ;
        RECT 175.950 697.050 178.050 699.150 ;
        RECT 178.950 698.850 181.050 700.950 ;
        RECT 184.950 700.050 187.050 702.150 ;
        RECT 187.950 698.850 190.050 700.950 ;
        RECT 190.950 700.050 193.050 702.150 ;
        RECT 202.950 701.850 205.050 703.950 ;
        RECT 205.950 703.050 208.050 705.150 ;
        RECT 203.100 700.050 204.900 701.850 ;
        RECT 179.100 697.050 180.900 698.850 ;
        RECT 188.100 697.050 189.900 698.850 ;
        RECT 191.850 696.750 193.050 700.050 ;
        RECT 191.850 695.700 195.600 696.750 ;
        RECT 206.400 695.700 207.600 703.050 ;
        RECT 208.950 701.850 211.050 703.950 ;
        RECT 209.100 700.050 210.900 701.850 ;
        RECT 215.700 700.950 217.050 707.550 ;
        RECT 223.800 707.400 225.600 719.400 ;
        RECT 229.800 713.400 231.600 719.400 ;
        RECT 155.400 687.600 157.200 690.600 ;
        RECT 161.700 687.600 163.500 693.600 ;
        RECT 170.400 691.950 175.800 693.600 ;
        RECT 174.000 687.600 175.800 691.950 ;
        RECT 185.400 692.700 193.200 694.050 ;
        RECT 185.400 687.600 187.200 692.700 ;
        RECT 191.400 687.600 193.200 692.700 ;
        RECT 194.400 693.600 195.600 695.700 ;
        RECT 204.000 694.800 207.600 695.700 ;
        RECT 214.950 698.850 217.050 700.950 ;
        RECT 218.400 706.200 220.200 706.650 ;
        RECT 224.400 706.200 225.600 707.400 ;
        RECT 218.400 705.000 225.600 706.200 ;
        RECT 218.400 704.850 220.200 705.000 ;
        RECT 194.400 687.600 196.200 693.600 ;
        RECT 204.000 687.600 205.800 694.800 ;
        RECT 214.950 693.600 216.000 698.850 ;
        RECT 218.400 696.600 219.300 704.850 ;
        RECT 221.100 702.150 222.900 703.950 ;
        RECT 220.950 700.050 223.050 702.150 ;
        RECT 230.400 700.950 231.600 713.400 ;
        RECT 245.700 707.400 247.500 719.400 ;
        RECT 258.600 707.400 260.400 719.400 ;
        RECT 268.800 713.400 270.600 719.400 ;
        RECT 242.250 705.150 244.050 706.950 ;
        RECT 241.950 703.050 244.050 705.150 ;
        RECT 245.850 702.150 247.050 707.400 ;
        RECT 258.000 706.350 260.400 707.400 ;
        RECT 251.100 702.150 252.900 703.950 ;
        RECT 254.100 702.150 255.900 703.950 ;
        RECT 224.100 699.150 225.900 700.950 ;
        RECT 223.950 697.050 226.050 699.150 ;
        RECT 229.950 698.850 232.050 700.950 ;
        RECT 233.100 699.150 234.900 700.950 ;
        RECT 244.950 700.050 247.050 702.150 ;
        RECT 218.250 695.700 220.050 696.600 ;
        RECT 218.250 694.800 221.700 695.700 ;
        RECT 214.800 687.600 216.600 693.600 ;
        RECT 220.800 690.600 221.700 694.800 ;
        RECT 230.400 690.600 231.600 698.850 ;
        RECT 232.950 697.050 235.050 699.150 ;
        RECT 244.950 696.750 246.150 700.050 ;
        RECT 247.950 698.850 250.050 700.950 ;
        RECT 250.950 700.050 253.050 702.150 ;
        RECT 253.950 700.050 256.050 702.150 ;
        RECT 258.000 699.150 259.050 706.350 ;
        RECT 260.100 702.150 261.900 703.950 ;
        RECT 259.950 700.050 262.050 702.150 ;
        RECT 269.400 700.950 270.600 713.400 ;
        RECT 280.500 707.400 282.300 719.400 ;
        RECT 294.600 707.400 296.400 719.400 ;
        RECT 304.800 707.400 306.600 719.400 ;
        RECT 307.800 708.300 309.600 719.400 ;
        RECT 313.800 708.300 315.600 719.400 ;
        RECT 307.800 707.400 315.600 708.300 ;
        RECT 322.500 707.400 324.300 719.400 ;
        RECT 340.800 707.400 342.600 719.400 ;
        RECT 350.400 713.400 352.200 719.400 ;
        RECT 361.800 718.500 369.600 719.400 ;
        RECT 275.100 702.150 276.900 703.950 ;
        RECT 280.950 702.150 282.150 707.400 ;
        RECT 283.950 705.150 285.750 706.950 ;
        RECT 294.000 706.350 296.400 707.400 ;
        RECT 283.950 703.050 286.050 705.150 ;
        RECT 290.100 702.150 291.900 703.950 ;
        RECT 248.100 697.050 249.900 698.850 ;
        RECT 256.950 697.050 259.050 699.150 ;
        RECT 268.950 698.850 271.050 700.950 ;
        RECT 272.100 699.150 273.900 700.950 ;
        RECT 274.950 700.050 277.050 702.150 ;
        RECT 242.400 695.700 246.150 696.750 ;
        RECT 242.400 693.600 243.600 695.700 ;
        RECT 220.800 687.600 222.600 690.600 ;
        RECT 229.800 687.600 231.600 690.600 ;
        RECT 241.800 687.600 243.600 693.600 ;
        RECT 244.800 692.700 252.600 694.050 ;
        RECT 244.800 687.600 246.600 692.700 ;
        RECT 250.800 687.600 252.600 692.700 ;
        RECT 258.000 690.600 259.050 697.050 ;
        RECT 269.400 690.600 270.600 698.850 ;
        RECT 271.950 697.050 274.050 699.150 ;
        RECT 277.950 698.850 280.050 700.950 ;
        RECT 280.950 700.050 283.050 702.150 ;
        RECT 289.950 700.050 292.050 702.150 ;
        RECT 278.100 697.050 279.900 698.850 ;
        RECT 281.850 696.750 283.050 700.050 ;
        RECT 294.000 699.150 295.050 706.350 ;
        RECT 296.100 702.150 297.900 703.950 ;
        RECT 305.400 702.150 306.300 707.400 ;
        RECT 317.100 702.150 318.900 703.950 ;
        RECT 322.950 702.150 324.150 707.400 ;
        RECT 325.950 705.150 327.750 706.950 ;
        RECT 325.950 703.050 328.050 705.150 ;
        RECT 295.950 700.050 298.050 702.150 ;
        RECT 304.950 700.050 307.050 702.150 ;
        RECT 292.950 697.050 295.050 699.150 ;
        RECT 281.850 695.700 285.600 696.750 ;
        RECT 257.400 687.600 259.200 690.600 ;
        RECT 268.800 687.600 270.600 690.600 ;
        RECT 275.400 692.700 283.200 694.050 ;
        RECT 275.400 687.600 277.200 692.700 ;
        RECT 281.400 687.600 283.200 692.700 ;
        RECT 284.400 693.600 285.600 695.700 ;
        RECT 284.400 687.600 286.200 693.600 ;
        RECT 294.000 690.600 295.050 697.050 ;
        RECT 305.400 693.600 306.300 700.050 ;
        RECT 307.950 698.850 310.050 700.950 ;
        RECT 311.100 699.150 312.900 700.950 ;
        RECT 308.100 697.050 309.900 698.850 ;
        RECT 310.950 697.050 313.050 699.150 ;
        RECT 313.950 698.850 316.050 700.950 ;
        RECT 316.950 700.050 319.050 702.150 ;
        RECT 319.950 698.850 322.050 700.950 ;
        RECT 322.950 700.050 325.050 702.150 ;
        RECT 340.950 700.950 342.300 707.400 ;
        RECT 350.400 705.150 351.600 713.400 ;
        RECT 361.800 707.400 363.600 718.500 ;
        RECT 364.800 706.500 366.600 717.600 ;
        RECT 367.800 708.600 369.600 718.500 ;
        RECT 373.800 708.600 375.600 719.400 ;
        RECT 367.800 707.700 375.600 708.600 ;
        RECT 385.500 707.400 387.300 719.400 ;
        RECT 398.400 713.400 400.200 719.400 ;
        RECT 413.400 713.400 415.200 719.400 ;
        RECT 364.800 705.600 368.850 706.500 ;
        RECT 346.950 701.850 349.050 703.950 ;
        RECT 349.950 703.050 352.050 705.150 ;
        RECT 314.100 697.050 315.900 698.850 ;
        RECT 320.100 697.050 321.900 698.850 ;
        RECT 323.850 696.750 325.050 700.050 ;
        RECT 337.950 698.850 342.300 700.950 ;
        RECT 343.950 698.850 346.050 700.950 ;
        RECT 347.100 700.050 348.900 701.850 ;
        RECT 323.850 695.700 327.600 696.750 ;
        RECT 305.400 691.950 310.800 693.600 ;
        RECT 293.400 687.600 295.200 690.600 ;
        RECT 309.000 687.600 310.800 691.950 ;
        RECT 317.400 692.700 325.200 694.050 ;
        RECT 317.400 687.600 319.200 692.700 ;
        RECT 323.400 687.600 325.200 692.700 ;
        RECT 326.400 693.600 327.600 695.700 ;
        RECT 340.950 693.600 342.300 698.850 ;
        RECT 344.100 697.050 345.900 698.850 ;
        RECT 350.400 695.700 351.600 703.050 ;
        RECT 352.950 701.850 355.050 703.950 ;
        RECT 362.100 702.150 363.900 703.950 ;
        RECT 367.950 702.150 368.850 705.600 ;
        RECT 373.950 702.150 375.750 703.950 ;
        RECT 380.100 702.150 381.900 703.950 ;
        RECT 385.950 702.150 387.150 707.400 ;
        RECT 388.950 705.150 390.750 706.950 ;
        RECT 398.400 705.150 399.600 713.400 ;
        RECT 388.950 703.050 391.050 705.150 ;
        RECT 353.100 700.050 354.900 701.850 ;
        RECT 361.950 700.050 364.050 702.150 ;
        RECT 364.950 698.850 367.050 700.950 ;
        RECT 367.950 700.050 370.050 702.150 ;
        RECT 365.250 697.050 367.050 698.850 ;
        RECT 350.400 694.800 354.000 695.700 ;
        RECT 326.400 687.600 328.200 693.600 ;
        RECT 340.800 687.600 342.600 693.600 ;
        RECT 352.200 687.600 354.000 694.800 ;
        RECT 369.000 693.600 370.050 700.050 ;
        RECT 370.950 698.850 373.050 700.950 ;
        RECT 373.950 700.050 376.050 702.150 ;
        RECT 379.950 700.050 382.050 702.150 ;
        RECT 382.950 698.850 385.050 700.950 ;
        RECT 385.950 700.050 388.050 702.150 ;
        RECT 394.950 701.850 397.050 703.950 ;
        RECT 397.950 703.050 400.050 705.150 ;
        RECT 395.100 700.050 396.900 701.850 ;
        RECT 370.950 697.050 372.750 698.850 ;
        RECT 383.100 697.050 384.900 698.850 ;
        RECT 373.950 696.450 376.050 697.050 ;
        RECT 379.950 696.450 382.050 697.050 ;
        RECT 373.950 695.550 382.050 696.450 ;
        RECT 386.850 696.750 388.050 700.050 ;
        RECT 386.850 695.700 390.600 696.750 ;
        RECT 373.950 694.950 376.050 695.550 ;
        RECT 379.950 694.950 382.050 695.550 ;
        RECT 369.000 687.600 370.800 693.600 ;
        RECT 380.400 692.700 388.200 694.050 ;
        RECT 380.400 687.600 382.200 692.700 ;
        RECT 386.400 687.600 388.200 692.700 ;
        RECT 389.400 693.600 390.600 695.700 ;
        RECT 398.400 695.700 399.600 703.050 ;
        RECT 400.950 701.850 403.050 703.950 ;
        RECT 401.100 700.050 402.900 701.850 ;
        RECT 413.400 700.950 414.600 713.400 ;
        RECT 424.800 707.400 426.600 719.400 ;
        RECT 425.400 702.150 426.600 707.400 ;
        RECT 431.400 713.400 433.200 719.400 ;
        RECT 431.400 706.500 432.600 713.400 ;
        RECT 437.700 707.400 439.500 719.400 ;
        RECT 444.150 707.400 445.950 719.400 ;
        RECT 452.550 713.400 454.350 719.400 ;
        RECT 452.550 712.500 453.750 713.400 ;
        RECT 460.350 712.500 462.150 719.400 ;
        RECT 468.150 713.400 469.950 719.400 ;
        RECT 448.950 710.400 453.750 712.500 ;
        RECT 456.450 711.450 463.050 712.500 ;
        RECT 456.450 710.700 458.250 711.450 ;
        RECT 461.250 710.700 463.050 711.450 ;
        RECT 468.150 711.300 472.050 713.400 ;
        RECT 452.550 709.500 453.750 710.400 ;
        RECT 465.450 709.800 467.250 710.400 ;
        RECT 452.550 708.300 460.050 709.500 ;
        RECT 458.250 707.700 460.050 708.300 ;
        RECT 460.950 708.900 467.250 709.800 ;
        RECT 431.400 705.600 437.100 706.500 ;
        RECT 435.150 704.700 437.100 705.600 ;
        RECT 431.100 702.150 432.900 703.950 ;
        RECT 410.100 699.150 411.900 700.950 ;
        RECT 409.950 697.050 412.050 699.150 ;
        RECT 412.950 698.850 415.050 700.950 ;
        RECT 424.950 700.050 427.050 702.150 ;
        RECT 398.400 694.800 402.000 695.700 ;
        RECT 389.400 687.600 391.200 693.600 ;
        RECT 400.200 687.600 402.000 694.800 ;
        RECT 413.400 690.600 414.600 698.850 ;
        RECT 425.400 693.600 426.600 700.050 ;
        RECT 427.950 698.850 430.050 700.950 ;
        RECT 430.950 700.050 433.050 702.150 ;
        RECT 428.100 697.050 429.900 698.850 ;
        RECT 435.150 696.300 436.050 704.700 ;
        RECT 438.000 702.150 439.200 707.400 ;
        RECT 436.950 700.050 439.200 702.150 ;
        RECT 435.150 695.400 437.100 696.300 ;
        RECT 413.400 687.600 415.200 690.600 ;
        RECT 424.800 687.600 426.600 693.600 ;
        RECT 432.000 694.500 437.100 695.400 ;
        RECT 432.000 690.600 433.200 694.500 ;
        RECT 438.000 693.600 439.200 700.050 ;
        RECT 444.150 706.800 455.250 707.400 ;
        RECT 460.950 706.800 461.850 708.900 ;
        RECT 465.450 708.600 467.250 708.900 ;
        RECT 468.150 708.600 470.850 710.400 ;
        RECT 468.150 707.700 469.050 708.600 ;
        RECT 444.150 706.200 461.850 706.800 ;
        RECT 444.150 693.600 445.050 706.200 ;
        RECT 453.450 705.900 461.850 706.200 ;
        RECT 463.050 706.800 469.050 707.700 ;
        RECT 469.950 706.800 472.050 707.700 ;
        RECT 475.650 707.400 477.450 719.400 ;
        RECT 453.450 705.600 455.250 705.900 ;
        RECT 463.050 702.150 463.950 706.800 ;
        RECT 469.950 705.600 474.150 706.800 ;
        RECT 473.250 703.800 475.050 705.600 ;
        RECT 454.950 701.100 457.050 702.150 ;
        RECT 446.100 699.150 447.900 700.950 ;
        RECT 449.100 700.050 457.050 701.100 ;
        RECT 460.950 700.050 463.950 702.150 ;
        RECT 449.100 699.300 450.900 700.050 ;
        RECT 447.000 698.400 447.900 699.150 ;
        RECT 452.100 698.400 453.900 699.000 ;
        RECT 447.000 697.200 453.900 698.400 ;
        RECT 452.850 696.000 453.900 697.200 ;
        RECT 463.050 696.000 463.950 700.050 ;
        RECT 472.950 699.750 475.050 700.050 ;
        RECT 471.150 697.950 475.050 699.750 ;
        RECT 476.250 697.950 477.450 707.400 ;
        RECT 487.800 706.500 489.600 719.400 ;
        RECT 493.800 706.500 495.600 719.400 ;
        RECT 499.800 706.500 501.600 719.400 ;
        RECT 505.800 706.500 507.600 719.400 ;
        RECT 517.500 707.400 519.300 719.400 ;
        RECT 535.800 713.400 537.600 719.400 ;
        RECT 486.900 705.300 489.600 706.500 ;
        RECT 491.700 705.300 495.600 706.500 ;
        RECT 497.700 705.300 501.600 706.500 ;
        RECT 503.700 705.300 507.600 706.500 ;
        RECT 486.900 700.950 487.800 705.300 ;
        RECT 484.950 698.850 487.800 700.950 ;
        RECT 452.850 695.100 463.950 696.000 ;
        RECT 472.950 695.850 477.450 697.950 ;
        RECT 452.850 694.200 453.900 695.100 ;
        RECT 463.050 694.800 463.950 695.100 ;
        RECT 431.400 687.600 433.200 690.600 ;
        RECT 437.700 687.600 439.500 693.600 ;
        RECT 444.150 687.600 445.950 693.600 ;
        RECT 448.950 691.500 451.050 693.600 ;
        RECT 452.550 692.400 454.350 694.200 ;
        RECT 455.850 693.450 457.650 694.200 ;
        RECT 455.850 692.400 460.800 693.450 ;
        RECT 463.050 693.000 464.850 694.800 ;
        RECT 476.250 693.600 477.450 695.850 ;
        RECT 486.900 695.700 487.800 698.850 ;
        RECT 488.700 697.800 490.500 698.400 ;
        RECT 491.700 697.800 492.900 705.300 ;
        RECT 488.700 696.600 492.900 697.800 ;
        RECT 494.700 697.800 496.500 698.400 ;
        RECT 497.700 697.800 498.900 705.300 ;
        RECT 494.700 696.600 498.900 697.800 ;
        RECT 500.700 697.800 502.500 698.400 ;
        RECT 503.700 697.800 504.900 705.300 ;
        RECT 512.100 702.150 513.900 703.950 ;
        RECT 517.950 702.150 519.150 707.400 ;
        RECT 520.950 705.150 522.750 706.950 ;
        RECT 536.400 705.150 537.600 713.400 ;
        RECT 542.550 707.400 544.350 719.400 ;
        RECT 550.050 713.400 551.850 719.400 ;
        RECT 547.950 711.300 551.850 713.400 ;
        RECT 557.850 712.500 559.650 719.400 ;
        RECT 565.650 713.400 567.450 719.400 ;
        RECT 566.250 712.500 567.450 713.400 ;
        RECT 556.950 711.450 563.550 712.500 ;
        RECT 556.950 710.700 558.750 711.450 ;
        RECT 561.750 710.700 563.550 711.450 ;
        RECT 566.250 710.400 571.050 712.500 ;
        RECT 549.150 708.600 551.850 710.400 ;
        RECT 552.750 709.800 554.550 710.400 ;
        RECT 552.750 708.900 559.050 709.800 ;
        RECT 566.250 709.500 567.450 710.400 ;
        RECT 552.750 708.600 554.550 708.900 ;
        RECT 550.950 707.700 551.850 708.600 ;
        RECT 520.950 703.050 523.050 705.150 ;
        RECT 505.950 698.850 508.050 700.950 ;
        RECT 511.950 700.050 514.050 702.150 ;
        RECT 514.950 698.850 517.050 700.950 ;
        RECT 517.950 700.050 520.050 702.150 ;
        RECT 532.950 701.850 535.050 703.950 ;
        RECT 535.950 703.050 538.050 705.150 ;
        RECT 533.100 700.050 534.900 701.850 ;
        RECT 500.700 696.600 504.900 697.800 ;
        RECT 506.100 697.050 507.900 698.850 ;
        RECT 515.100 697.050 516.900 698.850 ;
        RECT 491.700 695.700 492.900 696.600 ;
        RECT 497.700 695.700 498.900 696.600 ;
        RECT 503.700 695.700 504.900 696.600 ;
        RECT 518.850 696.750 520.050 700.050 ;
        RECT 518.850 695.700 522.600 696.750 ;
        RECT 536.400 695.700 537.600 703.050 ;
        RECT 538.950 701.850 541.050 703.950 ;
        RECT 539.100 700.050 540.900 701.850 ;
        RECT 486.900 694.500 489.600 695.700 ;
        RECT 491.700 694.500 495.600 695.700 ;
        RECT 497.700 694.500 501.600 695.700 ;
        RECT 503.700 694.500 507.600 695.700 ;
        RECT 469.950 692.700 472.050 693.600 ;
        RECT 450.000 690.600 451.050 691.500 ;
        RECT 459.750 690.600 460.800 692.400 ;
        RECT 468.300 691.500 472.050 692.700 ;
        RECT 468.300 690.600 469.350 691.500 ;
        RECT 450.000 689.700 453.750 690.600 ;
        RECT 451.950 687.600 453.750 689.700 ;
        RECT 459.750 687.600 461.550 690.600 ;
        RECT 467.550 687.600 469.350 690.600 ;
        RECT 475.650 687.600 477.450 693.600 ;
        RECT 487.800 687.600 489.600 694.500 ;
        RECT 493.800 687.600 495.600 694.500 ;
        RECT 499.800 687.600 501.600 694.500 ;
        RECT 505.800 687.600 507.600 694.500 ;
        RECT 512.400 692.700 520.200 694.050 ;
        RECT 512.400 687.600 514.200 692.700 ;
        RECT 518.400 687.600 520.200 692.700 ;
        RECT 521.400 693.600 522.600 695.700 ;
        RECT 534.000 694.800 537.600 695.700 ;
        RECT 542.550 697.950 543.750 707.400 ;
        RECT 547.950 706.800 550.050 707.700 ;
        RECT 550.950 706.800 556.950 707.700 ;
        RECT 545.850 705.600 550.050 706.800 ;
        RECT 544.950 703.800 546.750 705.600 ;
        RECT 556.050 702.150 556.950 706.800 ;
        RECT 558.150 706.800 559.050 708.900 ;
        RECT 559.950 708.300 567.450 709.500 ;
        RECT 559.950 707.700 561.750 708.300 ;
        RECT 574.050 707.400 575.850 719.400 ;
        RECT 564.750 706.800 575.850 707.400 ;
        RECT 558.150 706.200 575.850 706.800 ;
        RECT 558.150 705.900 566.550 706.200 ;
        RECT 564.750 705.600 566.550 705.900 ;
        RECT 556.050 700.050 559.050 702.150 ;
        RECT 562.950 701.100 565.050 702.150 ;
        RECT 562.950 700.050 570.900 701.100 ;
        RECT 544.950 699.750 547.050 700.050 ;
        RECT 544.950 697.950 548.850 699.750 ;
        RECT 542.550 695.850 547.050 697.950 ;
        RECT 556.050 696.000 556.950 700.050 ;
        RECT 569.100 699.300 570.900 700.050 ;
        RECT 572.100 699.150 573.900 700.950 ;
        RECT 566.100 698.400 567.900 699.000 ;
        RECT 572.100 698.400 573.000 699.150 ;
        RECT 566.100 697.200 573.000 698.400 ;
        RECT 566.100 696.000 567.150 697.200 ;
        RECT 521.400 687.600 523.200 693.600 ;
        RECT 534.000 687.600 535.800 694.800 ;
        RECT 542.550 693.600 543.750 695.850 ;
        RECT 556.050 695.100 567.150 696.000 ;
        RECT 556.050 694.800 556.950 695.100 ;
        RECT 542.550 687.600 544.350 693.600 ;
        RECT 547.950 692.700 550.050 693.600 ;
        RECT 555.150 693.000 556.950 694.800 ;
        RECT 566.100 694.200 567.150 695.100 ;
        RECT 562.350 693.450 564.150 694.200 ;
        RECT 547.950 691.500 551.700 692.700 ;
        RECT 550.650 690.600 551.700 691.500 ;
        RECT 559.200 692.400 564.150 693.450 ;
        RECT 565.650 692.400 567.450 694.200 ;
        RECT 574.950 693.600 575.850 706.200 ;
        RECT 581.400 706.500 583.200 719.400 ;
        RECT 587.400 706.500 589.200 719.400 ;
        RECT 593.400 706.500 595.200 719.400 ;
        RECT 599.400 706.500 601.200 719.400 ;
        RECT 613.200 713.400 615.000 719.400 ;
        RECT 581.400 705.300 585.300 706.500 ;
        RECT 587.400 705.300 591.300 706.500 ;
        RECT 593.400 705.300 597.300 706.500 ;
        RECT 599.400 705.300 602.100 706.500 ;
        RECT 580.950 698.850 583.050 700.950 ;
        RECT 581.100 697.050 582.900 698.850 ;
        RECT 584.100 697.800 585.300 705.300 ;
        RECT 586.500 697.800 588.300 698.400 ;
        RECT 584.100 696.600 588.300 697.800 ;
        RECT 590.100 697.800 591.300 705.300 ;
        RECT 592.500 697.800 594.300 698.400 ;
        RECT 590.100 696.600 594.300 697.800 ;
        RECT 596.100 697.800 597.300 705.300 ;
        RECT 601.200 700.950 602.100 705.300 ;
        RECT 613.500 700.950 615.000 713.400 ;
        RECT 619.800 713.400 621.600 719.400 ;
        RECT 619.800 709.350 621.000 713.400 ;
        RECT 625.800 712.500 627.600 719.400 ;
        RECT 632.400 716.400 634.200 719.400 ;
        RECT 635.400 716.400 637.200 719.400 ;
        RECT 638.400 716.400 640.200 719.400 ;
        RECT 632.850 715.200 634.050 716.400 ;
        RECT 631.950 713.100 634.050 715.200 ;
        RECT 635.400 712.950 637.050 716.400 ;
        RECT 621.900 711.300 627.600 712.500 ;
        RECT 628.500 712.050 630.300 712.500 ;
        RECT 634.950 712.050 637.050 712.950 ;
        RECT 621.900 710.700 623.700 711.300 ;
        RECT 628.500 710.850 637.050 712.050 ;
        RECT 628.500 710.700 630.300 710.850 ;
        RECT 638.850 709.350 640.050 716.400 ;
        RECT 642.000 712.500 643.800 719.400 ;
        RECT 648.000 713.400 649.800 719.400 ;
        RECT 654.900 716.400 656.850 719.400 ;
        RECT 657.900 716.400 660.000 719.400 ;
        RECT 660.900 716.400 663.150 719.400 ;
        RECT 655.650 715.050 656.850 716.400 ;
        RECT 658.950 715.050 660.000 716.400 ;
        RECT 662.250 715.050 663.150 716.400 ;
        RECT 648.000 712.500 649.050 713.400 ;
        RECT 655.650 712.950 658.050 715.050 ;
        RECT 658.950 712.950 661.050 715.050 ;
        RECT 661.950 712.950 664.050 715.050 ;
        RECT 642.000 712.200 645.000 712.500 ;
        RECT 641.100 710.400 645.000 712.200 ;
        RECT 646.950 710.400 649.050 712.500 ;
        RECT 667.500 710.700 669.300 719.400 ;
        RECT 673.500 713.400 675.300 719.400 ;
        RECT 674.250 712.500 675.300 713.400 ;
        RECT 674.250 711.600 678.300 712.500 ;
        RECT 601.200 698.850 604.050 700.950 ;
        RECT 610.950 698.850 615.000 700.950 ;
        RECT 598.500 697.800 600.300 698.400 ;
        RECT 596.100 696.600 600.300 697.800 ;
        RECT 584.100 695.700 585.300 696.600 ;
        RECT 590.100 695.700 591.300 696.600 ;
        RECT 596.100 695.700 597.300 696.600 ;
        RECT 601.200 695.700 602.100 698.850 ;
        RECT 559.200 690.600 560.250 692.400 ;
        RECT 568.950 691.500 571.050 693.600 ;
        RECT 568.950 690.600 570.000 691.500 ;
        RECT 550.650 687.600 552.450 690.600 ;
        RECT 558.450 687.600 560.250 690.600 ;
        RECT 566.250 689.700 570.000 690.600 ;
        RECT 566.250 687.600 568.050 689.700 ;
        RECT 574.050 687.600 575.850 693.600 ;
        RECT 581.400 694.500 585.300 695.700 ;
        RECT 587.400 694.500 591.300 695.700 ;
        RECT 593.400 694.500 597.300 695.700 ;
        RECT 599.400 694.500 602.100 695.700 ;
        RECT 581.400 687.600 583.200 694.500 ;
        RECT 587.400 687.600 589.200 694.500 ;
        RECT 593.400 687.600 595.200 694.500 ;
        RECT 599.400 687.600 601.200 694.500 ;
        RECT 613.500 690.600 615.000 698.850 ;
        RECT 613.200 687.600 615.000 690.600 ;
        RECT 617.100 708.450 634.050 709.350 ;
        RECT 617.100 693.600 618.000 708.450 ;
        RECT 618.900 706.350 631.050 707.550 ;
        RECT 631.950 707.250 634.050 708.450 ;
        RECT 637.950 708.300 640.050 709.350 ;
        RECT 656.100 709.650 673.800 710.700 ;
        RECT 656.100 708.300 658.050 709.650 ;
        RECT 672.000 708.900 673.800 709.650 ;
        RECT 637.950 707.250 658.050 708.300 ;
        RECT 658.950 708.150 661.050 708.750 ;
        RECT 658.950 706.950 670.500 708.150 ;
        RECT 658.950 706.650 661.050 706.950 ;
        RECT 668.700 706.350 670.500 706.950 ;
        RECT 618.900 705.750 620.700 706.350 ;
        RECT 630.000 705.450 658.050 706.350 ;
        RECT 630.000 705.150 670.050 705.450 ;
        RECT 622.950 701.100 625.050 705.150 ;
        RECT 656.100 704.550 670.050 705.150 ;
        RECT 626.100 702.000 633.150 703.800 ;
        RECT 622.950 700.050 631.200 701.100 ;
        RECT 618.900 698.700 620.700 699.000 ;
        RECT 623.700 698.700 625.500 699.000 ;
        RECT 618.900 697.200 626.700 698.700 ;
        RECT 630.150 698.250 631.200 700.050 ;
        RECT 632.250 700.350 633.150 702.000 ;
        RECT 634.500 703.500 649.050 704.250 ;
        RECT 655.800 703.500 657.600 703.650 ;
        RECT 634.500 703.050 657.600 703.500 ;
        RECT 666.150 703.350 670.050 704.550 ;
        RECT 634.500 701.250 636.300 703.050 ;
        RECT 646.950 702.450 657.600 703.050 ;
        RECT 646.950 702.150 649.050 702.450 ;
        RECT 655.800 701.850 657.600 702.450 ;
        RECT 658.500 702.450 665.250 703.350 ;
        RECT 667.950 703.050 670.050 703.350 ;
        RECT 642.750 701.250 644.850 701.550 ;
        RECT 632.250 699.300 641.850 700.350 ;
        RECT 642.750 699.450 646.650 701.250 ;
        RECT 658.500 700.950 659.550 702.450 ;
        RECT 647.550 700.050 659.550 700.950 ;
        RECT 640.950 698.550 641.850 699.300 ;
        RECT 647.550 698.550 648.600 700.050 ;
        RECT 660.450 699.750 662.250 701.550 ;
        RECT 664.050 700.050 665.250 702.450 ;
        RECT 673.950 701.850 676.050 703.950 ;
        RECT 674.100 700.050 675.900 701.850 ;
        RECT 630.150 697.200 640.050 698.250 ;
        RECT 640.950 697.200 648.600 698.550 ;
        RECT 649.950 697.350 653.850 699.150 ;
        RECT 625.200 693.600 626.700 697.200 ;
        RECT 639.000 696.300 640.050 697.200 ;
        RECT 649.950 697.050 652.050 697.350 ;
        RECT 657.150 696.300 658.950 696.750 ;
        RECT 660.450 696.300 661.500 699.750 ;
        RECT 664.050 699.000 675.900 700.050 ;
        RECT 677.100 698.100 678.300 711.600 ;
        RECT 682.800 707.400 684.600 719.400 ;
        RECT 685.800 708.300 687.600 719.400 ;
        RECT 691.800 708.300 693.600 719.400 ;
        RECT 700.200 713.400 702.000 719.400 ;
        RECT 685.800 707.400 693.600 708.300 ;
        RECT 683.400 702.150 684.300 707.400 ;
        RECT 682.950 700.050 685.050 702.150 ;
        RECT 700.500 700.950 702.000 713.400 ;
        RECT 706.800 713.400 708.600 719.400 ;
        RECT 706.800 709.350 708.000 713.400 ;
        RECT 712.800 712.500 714.600 719.400 ;
        RECT 719.400 716.400 721.200 719.400 ;
        RECT 722.400 716.400 724.200 719.400 ;
        RECT 725.400 716.400 727.200 719.400 ;
        RECT 719.850 715.200 721.050 716.400 ;
        RECT 718.950 713.100 721.050 715.200 ;
        RECT 722.400 712.950 724.050 716.400 ;
        RECT 708.900 711.300 714.600 712.500 ;
        RECT 715.500 712.050 717.300 712.500 ;
        RECT 721.950 712.050 724.050 712.950 ;
        RECT 708.900 710.700 710.700 711.300 ;
        RECT 715.500 710.850 724.050 712.050 ;
        RECT 715.500 710.700 717.300 710.850 ;
        RECT 725.850 709.350 727.050 716.400 ;
        RECT 729.000 712.500 730.800 719.400 ;
        RECT 735.000 713.400 736.800 719.400 ;
        RECT 741.900 716.400 743.850 719.400 ;
        RECT 744.900 716.400 747.000 719.400 ;
        RECT 747.900 716.400 750.150 719.400 ;
        RECT 742.650 715.050 743.850 716.400 ;
        RECT 745.950 715.050 747.000 716.400 ;
        RECT 749.250 715.050 750.150 716.400 ;
        RECT 735.000 712.500 736.050 713.400 ;
        RECT 742.650 712.950 745.050 715.050 ;
        RECT 745.950 712.950 748.050 715.050 ;
        RECT 748.950 712.950 751.050 715.050 ;
        RECT 729.000 712.200 732.000 712.500 ;
        RECT 728.100 710.400 732.000 712.200 ;
        RECT 733.950 710.400 736.050 712.500 ;
        RECT 754.500 710.700 756.300 719.400 ;
        RECT 760.500 713.400 762.300 719.400 ;
        RECT 761.250 712.500 762.300 713.400 ;
        RECT 761.250 711.600 765.300 712.500 ;
        RECT 631.500 694.500 638.100 696.300 ;
        RECT 639.000 694.500 645.900 696.300 ;
        RECT 657.150 695.850 661.500 696.300 ;
        RECT 653.850 695.100 661.500 695.850 ;
        RECT 663.000 697.200 678.300 698.100 ;
        RECT 653.850 694.950 658.950 695.100 ;
        RECT 653.850 693.600 654.750 694.950 ;
        RECT 663.000 694.050 664.050 697.200 ;
        RECT 672.300 695.700 674.100 696.300 ;
        RECT 617.100 687.600 618.900 693.600 ;
        RECT 625.200 692.400 629.400 693.600 ;
        RECT 627.600 687.600 629.400 692.400 ;
        RECT 631.950 691.500 634.050 693.600 ;
        RECT 634.950 691.500 637.050 693.600 ;
        RECT 637.950 691.500 640.050 693.600 ;
        RECT 632.400 690.600 633.750 691.500 ;
        RECT 635.400 690.600 637.050 691.500 ;
        RECT 638.400 690.600 640.050 691.500 ;
        RECT 642.750 691.500 644.850 693.600 ;
        RECT 646.950 691.500 649.050 693.600 ;
        RECT 650.700 692.250 654.750 693.600 ;
        RECT 650.700 691.800 652.500 692.250 ;
        RECT 655.950 691.950 658.050 694.050 ;
        RECT 658.950 691.950 661.050 694.050 ;
        RECT 661.950 691.950 664.050 694.050 ;
        RECT 665.700 694.500 674.100 695.700 ;
        RECT 665.700 693.600 667.200 694.500 ;
        RECT 677.100 693.600 678.300 697.200 ;
        RECT 642.750 690.600 643.800 691.500 ;
        RECT 632.400 687.600 634.200 690.600 ;
        RECT 635.400 687.600 637.200 690.600 ;
        RECT 638.400 687.600 640.200 690.600 ;
        RECT 642.000 687.600 643.800 690.600 ;
        RECT 648.000 690.600 649.050 691.500 ;
        RECT 655.950 690.600 657.300 691.950 ;
        RECT 658.950 690.600 660.300 691.950 ;
        RECT 661.950 690.600 663.300 691.950 ;
        RECT 648.000 687.600 649.800 690.600 ;
        RECT 655.500 687.600 657.300 690.600 ;
        RECT 658.500 687.600 660.300 690.600 ;
        RECT 661.500 687.600 663.300 690.600 ;
        RECT 665.700 687.600 667.500 693.600 ;
        RECT 676.500 687.600 678.300 693.600 ;
        RECT 683.400 693.600 684.300 700.050 ;
        RECT 685.950 698.850 688.050 700.950 ;
        RECT 689.100 699.150 690.900 700.950 ;
        RECT 686.100 697.050 687.900 698.850 ;
        RECT 688.950 697.050 691.050 699.150 ;
        RECT 691.950 698.850 694.050 700.950 ;
        RECT 697.950 698.850 702.000 700.950 ;
        RECT 692.100 697.050 693.900 698.850 ;
        RECT 683.400 691.950 688.800 693.600 ;
        RECT 687.000 687.600 688.800 691.950 ;
        RECT 700.500 690.600 702.000 698.850 ;
        RECT 700.200 687.600 702.000 690.600 ;
        RECT 704.100 708.450 721.050 709.350 ;
        RECT 704.100 693.600 705.000 708.450 ;
        RECT 705.900 706.350 718.050 707.550 ;
        RECT 718.950 707.250 721.050 708.450 ;
        RECT 724.950 708.300 727.050 709.350 ;
        RECT 743.100 709.650 760.800 710.700 ;
        RECT 743.100 708.300 745.050 709.650 ;
        RECT 759.000 708.900 760.800 709.650 ;
        RECT 724.950 707.250 745.050 708.300 ;
        RECT 745.950 708.150 748.050 708.750 ;
        RECT 745.950 706.950 757.500 708.150 ;
        RECT 745.950 706.650 748.050 706.950 ;
        RECT 755.700 706.350 757.500 706.950 ;
        RECT 705.900 705.750 707.700 706.350 ;
        RECT 717.000 705.450 745.050 706.350 ;
        RECT 717.000 705.150 757.050 705.450 ;
        RECT 709.950 701.100 712.050 705.150 ;
        RECT 743.100 704.550 757.050 705.150 ;
        RECT 713.100 702.000 720.150 703.800 ;
        RECT 709.950 700.050 718.200 701.100 ;
        RECT 705.900 698.700 707.700 699.000 ;
        RECT 710.700 698.700 712.500 699.000 ;
        RECT 705.900 697.200 713.700 698.700 ;
        RECT 717.150 698.250 718.200 700.050 ;
        RECT 719.250 700.350 720.150 702.000 ;
        RECT 721.500 703.500 736.050 704.250 ;
        RECT 742.800 703.500 744.600 703.650 ;
        RECT 721.500 703.050 744.600 703.500 ;
        RECT 753.150 703.350 757.050 704.550 ;
        RECT 721.500 701.250 723.300 703.050 ;
        RECT 733.950 702.450 744.600 703.050 ;
        RECT 733.950 702.150 736.050 702.450 ;
        RECT 742.800 701.850 744.600 702.450 ;
        RECT 745.500 702.450 752.250 703.350 ;
        RECT 754.950 703.050 757.050 703.350 ;
        RECT 729.750 701.250 731.850 701.550 ;
        RECT 719.250 699.300 728.850 700.350 ;
        RECT 729.750 699.450 733.650 701.250 ;
        RECT 745.500 700.950 746.550 702.450 ;
        RECT 734.550 700.050 746.550 700.950 ;
        RECT 727.950 698.550 728.850 699.300 ;
        RECT 734.550 698.550 735.600 700.050 ;
        RECT 747.450 699.750 749.250 701.550 ;
        RECT 751.050 700.050 752.250 702.450 ;
        RECT 760.950 701.850 763.050 703.950 ;
        RECT 761.100 700.050 762.900 701.850 ;
        RECT 717.150 697.200 727.050 698.250 ;
        RECT 727.950 697.200 735.600 698.550 ;
        RECT 736.950 697.350 740.850 699.150 ;
        RECT 712.200 693.600 713.700 697.200 ;
        RECT 726.000 696.300 727.050 697.200 ;
        RECT 736.950 697.050 739.050 697.350 ;
        RECT 744.150 696.300 745.950 696.750 ;
        RECT 747.450 696.300 748.500 699.750 ;
        RECT 751.050 699.000 762.900 700.050 ;
        RECT 764.100 698.100 765.300 711.600 ;
        RECT 718.500 694.500 725.100 696.300 ;
        RECT 726.000 694.500 732.900 696.300 ;
        RECT 744.150 695.850 748.500 696.300 ;
        RECT 740.850 695.100 748.500 695.850 ;
        RECT 750.000 697.200 765.300 698.100 ;
        RECT 740.850 694.950 745.950 695.100 ;
        RECT 740.850 693.600 741.750 694.950 ;
        RECT 750.000 694.050 751.050 697.200 ;
        RECT 759.300 695.700 761.100 696.300 ;
        RECT 704.100 687.600 705.900 693.600 ;
        RECT 712.200 692.400 716.400 693.600 ;
        RECT 714.600 687.600 716.400 692.400 ;
        RECT 718.950 691.500 721.050 693.600 ;
        RECT 721.950 691.500 724.050 693.600 ;
        RECT 724.950 691.500 727.050 693.600 ;
        RECT 719.400 690.600 720.750 691.500 ;
        RECT 722.400 690.600 724.050 691.500 ;
        RECT 725.400 690.600 727.050 691.500 ;
        RECT 729.750 691.500 731.850 693.600 ;
        RECT 733.950 691.500 736.050 693.600 ;
        RECT 737.700 692.250 741.750 693.600 ;
        RECT 737.700 691.800 739.500 692.250 ;
        RECT 742.950 691.950 745.050 694.050 ;
        RECT 745.950 691.950 748.050 694.050 ;
        RECT 748.950 691.950 751.050 694.050 ;
        RECT 752.700 694.500 761.100 695.700 ;
        RECT 752.700 693.600 754.200 694.500 ;
        RECT 764.100 693.600 765.300 697.200 ;
        RECT 729.750 690.600 730.800 691.500 ;
        RECT 719.400 687.600 721.200 690.600 ;
        RECT 722.400 687.600 724.200 690.600 ;
        RECT 725.400 687.600 727.200 690.600 ;
        RECT 729.000 687.600 730.800 690.600 ;
        RECT 735.000 690.600 736.050 691.500 ;
        RECT 742.950 690.600 744.300 691.950 ;
        RECT 745.950 690.600 747.300 691.950 ;
        RECT 748.950 690.600 750.300 691.950 ;
        RECT 735.000 687.600 736.800 690.600 ;
        RECT 742.500 687.600 744.300 690.600 ;
        RECT 745.500 687.600 747.300 690.600 ;
        RECT 748.500 687.600 750.300 690.600 ;
        RECT 752.700 687.600 754.500 693.600 ;
        RECT 763.500 687.600 765.300 693.600 ;
        RECT 6.000 676.200 7.800 683.400 ;
        RECT 19.800 677.400 21.600 683.400 ;
        RECT 6.000 675.300 9.600 676.200 ;
        RECT 5.100 669.150 6.900 670.950 ;
        RECT 4.950 667.050 7.050 669.150 ;
        RECT 8.400 667.950 9.600 675.300 ;
        RECT 20.400 675.300 21.600 677.400 ;
        RECT 22.800 678.300 24.600 683.400 ;
        RECT 28.800 678.300 30.600 683.400 ;
        RECT 22.800 676.950 30.600 678.300 ;
        RECT 37.200 676.200 39.000 683.400 ;
        RECT 35.400 675.300 39.000 676.200 ;
        RECT 20.400 674.250 24.150 675.300 ;
        RECT 22.950 670.950 24.150 674.250 ;
        RECT 26.100 672.150 27.900 673.950 ;
        RECT 11.100 669.150 12.900 670.950 ;
        RECT 7.950 665.850 10.050 667.950 ;
        RECT 10.950 667.050 13.050 669.150 ;
        RECT 22.950 668.850 25.050 670.950 ;
        RECT 25.950 670.050 28.050 672.150 ;
        RECT 28.950 668.850 31.050 670.950 ;
        RECT 32.100 669.150 33.900 670.950 ;
        RECT 19.950 665.850 22.050 667.950 ;
        RECT 8.400 657.600 9.600 665.850 ;
        RECT 20.250 664.050 22.050 665.850 ;
        RECT 23.850 663.600 25.050 668.850 ;
        RECT 29.100 667.050 30.900 668.850 ;
        RECT 31.950 667.050 34.050 669.150 ;
        RECT 35.400 667.950 36.600 675.300 ;
        RECT 50.100 675.000 51.900 683.400 ;
        RECT 63.000 676.200 64.800 683.400 ;
        RECT 78.000 676.200 79.800 683.400 ;
        RECT 88.800 677.400 90.600 683.400 ;
        RECT 63.000 675.300 66.600 676.200 ;
        RECT 78.000 675.300 81.600 676.200 ;
        RECT 47.700 673.350 51.900 675.000 ;
        RECT 38.100 669.150 39.900 670.950 ;
        RECT 47.700 669.150 48.600 673.350 ;
        RECT 62.100 669.150 63.900 670.950 ;
        RECT 34.950 665.850 37.050 667.950 ;
        RECT 37.950 667.050 40.050 669.150 ;
        RECT 46.950 667.050 49.050 669.150 ;
        RECT 7.800 651.600 9.600 657.600 ;
        RECT 23.700 651.600 25.500 663.600 ;
        RECT 35.400 657.600 36.600 665.850 ;
        RECT 47.700 658.800 48.600 667.050 ;
        RECT 49.950 665.850 52.050 667.950 ;
        RECT 55.950 665.850 58.050 667.950 ;
        RECT 61.950 667.050 64.050 669.150 ;
        RECT 65.400 667.950 66.600 675.300 ;
        RECT 68.100 669.150 69.900 670.950 ;
        RECT 77.100 669.150 78.900 670.950 ;
        RECT 64.950 665.850 67.050 667.950 ;
        RECT 67.950 667.050 70.050 669.150 ;
        RECT 76.950 667.050 79.050 669.150 ;
        RECT 80.400 667.950 81.600 675.300 ;
        RECT 89.400 675.300 90.600 677.400 ;
        RECT 91.800 678.300 93.600 683.400 ;
        RECT 97.800 678.300 99.600 683.400 ;
        RECT 104.400 680.400 106.200 683.400 ;
        RECT 91.800 676.950 99.600 678.300 ;
        RECT 89.400 674.250 93.150 675.300 ;
        RECT 91.950 670.950 93.150 674.250 ;
        RECT 105.000 673.950 106.050 680.400 ;
        RECT 115.800 677.400 117.600 683.400 ;
        RECT 116.400 675.300 117.600 677.400 ;
        RECT 118.800 678.300 120.600 683.400 ;
        RECT 124.800 678.300 126.600 683.400 ;
        RECT 118.800 676.950 126.600 678.300 ;
        RECT 133.200 676.200 135.000 683.400 ;
        RECT 145.800 677.400 147.600 683.400 ;
        RECT 131.400 675.300 135.000 676.200 ;
        RECT 146.400 675.300 147.600 677.400 ;
        RECT 148.800 678.300 150.600 683.400 ;
        RECT 154.800 678.300 156.600 683.400 ;
        RECT 163.800 680.400 165.600 683.400 ;
        RECT 148.800 676.950 156.600 678.300 ;
        RECT 116.400 674.250 120.150 675.300 ;
        RECT 95.100 672.150 96.900 673.950 ;
        RECT 83.100 669.150 84.900 670.950 ;
        RECT 79.950 665.850 82.050 667.950 ;
        RECT 82.950 667.050 85.050 669.150 ;
        RECT 91.950 668.850 94.050 670.950 ;
        RECT 94.950 670.050 97.050 672.150 ;
        RECT 103.950 671.850 106.050 673.950 ;
        RECT 97.950 668.850 100.050 670.950 ;
        RECT 100.950 668.850 103.050 670.950 ;
        RECT 88.950 665.850 91.050 667.950 ;
        RECT 49.950 664.050 51.750 665.850 ;
        RECT 52.950 662.850 55.050 664.950 ;
        RECT 56.100 664.050 57.900 665.850 ;
        RECT 53.100 661.050 54.900 662.850 ;
        RECT 47.700 657.900 54.300 658.800 ;
        RECT 47.700 657.600 48.600 657.900 ;
        RECT 35.400 651.600 37.200 657.600 ;
        RECT 46.800 651.600 48.600 657.600 ;
        RECT 52.800 657.600 54.300 657.900 ;
        RECT 65.400 657.600 66.600 665.850 ;
        RECT 80.400 657.600 81.600 665.850 ;
        RECT 89.250 664.050 91.050 665.850 ;
        RECT 92.850 663.600 94.050 668.850 ;
        RECT 98.100 667.050 99.900 668.850 ;
        RECT 101.100 667.050 102.900 668.850 ;
        RECT 105.000 664.650 106.050 671.850 ;
        RECT 118.950 670.950 120.150 674.250 ;
        RECT 122.100 672.150 123.900 673.950 ;
        RECT 106.950 668.850 109.050 670.950 ;
        RECT 118.950 668.850 121.050 670.950 ;
        RECT 121.950 670.050 124.050 672.150 ;
        RECT 124.950 668.850 127.050 670.950 ;
        RECT 128.100 669.150 129.900 670.950 ;
        RECT 107.100 667.050 108.900 668.850 ;
        RECT 115.950 665.850 118.050 667.950 ;
        RECT 105.000 663.600 107.400 664.650 ;
        RECT 116.250 664.050 118.050 665.850 ;
        RECT 119.850 663.600 121.050 668.850 ;
        RECT 125.100 667.050 126.900 668.850 ;
        RECT 127.950 667.050 130.050 669.150 ;
        RECT 131.400 667.950 132.600 675.300 ;
        RECT 146.400 674.250 150.150 675.300 ;
        RECT 148.950 670.950 150.150 674.250 ;
        RECT 163.950 673.950 165.000 680.400 ;
        RECT 175.800 677.400 177.600 683.400 ;
        RECT 176.400 675.300 177.600 677.400 ;
        RECT 178.800 678.300 180.600 683.400 ;
        RECT 184.800 678.300 186.600 683.400 ;
        RECT 178.800 676.950 186.600 678.300 ;
        RECT 190.800 677.400 192.600 683.400 ;
        RECT 191.400 675.300 192.600 677.400 ;
        RECT 193.800 678.300 195.600 683.400 ;
        RECT 199.800 678.300 201.600 683.400 ;
        RECT 205.800 680.400 207.600 683.400 ;
        RECT 193.800 676.950 201.600 678.300 ;
        RECT 176.400 674.250 180.150 675.300 ;
        RECT 191.400 674.250 195.150 675.300 ;
        RECT 152.100 672.150 153.900 673.950 ;
        RECT 134.100 669.150 135.900 670.950 ;
        RECT 130.950 665.850 133.050 667.950 ;
        RECT 133.950 667.050 136.050 669.150 ;
        RECT 148.950 668.850 151.050 670.950 ;
        RECT 151.950 670.050 154.050 672.150 ;
        RECT 163.950 671.850 166.050 673.950 ;
        RECT 175.950 672.450 178.050 673.050 ;
        RECT 154.950 668.850 157.050 670.950 ;
        RECT 160.950 668.850 163.050 670.950 ;
        RECT 145.950 665.850 148.050 667.950 ;
        RECT 52.800 651.600 54.600 657.600 ;
        RECT 64.800 651.600 66.600 657.600 ;
        RECT 79.800 651.600 81.600 657.600 ;
        RECT 92.700 651.600 94.500 663.600 ;
        RECT 105.600 651.600 107.400 663.600 ;
        RECT 119.700 651.600 121.500 663.600 ;
        RECT 131.400 657.600 132.600 665.850 ;
        RECT 146.250 664.050 148.050 665.850 ;
        RECT 149.850 663.600 151.050 668.850 ;
        RECT 155.100 667.050 156.900 668.850 ;
        RECT 161.100 667.050 162.900 668.850 ;
        RECT 163.950 664.650 165.000 671.850 ;
        RECT 173.550 671.550 178.050 672.450 ;
        RECT 166.950 668.850 169.050 670.950 ;
        RECT 167.100 667.050 168.900 668.850 ;
        RECT 162.600 663.600 165.000 664.650 ;
        RECT 173.550 664.050 174.450 671.550 ;
        RECT 175.950 670.950 178.050 671.550 ;
        RECT 178.950 670.950 180.150 674.250 ;
        RECT 182.100 672.150 183.900 673.950 ;
        RECT 178.950 668.850 181.050 670.950 ;
        RECT 181.950 670.050 184.050 672.150 ;
        RECT 193.950 670.950 195.150 674.250 ;
        RECT 197.100 672.150 198.900 673.950 ;
        RECT 206.400 672.150 207.600 680.400 ;
        RECT 214.800 677.400 216.600 683.400 ;
        RECT 215.400 675.300 216.600 677.400 ;
        RECT 217.800 678.300 219.600 683.400 ;
        RECT 223.800 678.300 225.600 683.400 ;
        RECT 217.800 676.950 225.600 678.300 ;
        RECT 232.200 677.400 234.000 683.400 ;
        RECT 215.400 674.250 219.150 675.300 ;
        RECT 184.950 668.850 187.050 670.950 ;
        RECT 193.950 668.850 196.050 670.950 ;
        RECT 196.950 670.050 199.050 672.150 ;
        RECT 199.950 668.850 202.050 670.950 ;
        RECT 205.950 670.050 208.050 672.150 ;
        RECT 208.950 671.850 211.050 673.950 ;
        RECT 214.950 672.450 217.050 673.050 ;
        RECT 209.100 670.050 210.900 671.850 ;
        RECT 212.550 671.550 217.050 672.450 ;
        RECT 175.950 665.850 178.050 667.950 ;
        RECT 176.250 664.050 178.050 665.850 ;
        RECT 131.400 651.600 133.200 657.600 ;
        RECT 149.700 651.600 151.500 663.600 ;
        RECT 162.600 651.600 164.400 663.600 ;
        RECT 172.950 661.950 175.050 664.050 ;
        RECT 179.850 663.600 181.050 668.850 ;
        RECT 185.100 667.050 186.900 668.850 ;
        RECT 190.950 665.850 193.050 667.950 ;
        RECT 191.250 664.050 193.050 665.850 ;
        RECT 194.850 663.600 196.050 668.850 ;
        RECT 200.100 667.050 201.900 668.850 ;
        RECT 179.700 651.600 181.500 663.600 ;
        RECT 194.700 651.600 196.500 663.600 ;
        RECT 206.400 657.600 207.600 670.050 ;
        RECT 208.950 666.450 211.050 667.050 ;
        RECT 212.550 666.450 213.450 671.550 ;
        RECT 214.950 670.950 217.050 671.550 ;
        RECT 217.950 670.950 219.150 674.250 ;
        RECT 221.100 672.150 222.900 673.950 ;
        RECT 230.250 672.150 232.050 673.950 ;
        RECT 217.950 668.850 220.050 670.950 ;
        RECT 220.950 670.050 223.050 672.150 ;
        RECT 223.950 668.850 226.050 670.950 ;
        RECT 226.950 668.850 229.050 670.950 ;
        RECT 229.950 670.050 232.050 672.150 ;
        RECT 232.950 670.950 234.000 677.400 ;
        RECT 254.100 675.000 255.900 683.400 ;
        RECT 267.000 676.200 268.800 683.400 ;
        RECT 280.800 677.400 282.600 683.400 ;
        RECT 267.000 675.300 270.600 676.200 ;
        RECT 235.950 672.150 237.750 673.950 ;
        RECT 251.700 673.350 255.900 675.000 ;
        RECT 232.950 668.850 235.050 670.950 ;
        RECT 235.950 670.050 238.050 672.150 ;
        RECT 238.950 668.850 241.050 670.950 ;
        RECT 251.700 669.150 252.600 673.350 ;
        RECT 266.100 669.150 267.900 670.950 ;
        RECT 208.950 665.550 213.450 666.450 ;
        RECT 214.950 665.850 217.050 667.950 ;
        RECT 208.950 664.950 211.050 665.550 ;
        RECT 215.250 664.050 217.050 665.850 ;
        RECT 218.850 663.600 220.050 668.850 ;
        RECT 224.100 667.050 225.900 668.850 ;
        RECT 227.250 667.050 229.050 668.850 ;
        RECT 234.150 665.400 235.050 668.850 ;
        RECT 239.100 667.050 240.900 668.850 ;
        RECT 250.950 667.050 253.050 669.150 ;
        RECT 234.150 664.500 238.200 665.400 ;
        RECT 205.800 651.600 207.600 657.600 ;
        RECT 218.700 651.600 220.500 663.600 ;
        RECT 227.400 662.400 235.200 663.300 ;
        RECT 227.400 651.600 229.200 662.400 ;
        RECT 233.400 652.500 235.200 662.400 ;
        RECT 236.400 653.400 238.200 664.500 ;
        RECT 239.400 652.500 241.200 663.600 ;
        RECT 251.700 658.800 252.600 667.050 ;
        RECT 253.950 665.850 256.050 667.950 ;
        RECT 259.950 665.850 262.050 667.950 ;
        RECT 265.950 667.050 268.050 669.150 ;
        RECT 269.400 667.950 270.600 675.300 ;
        RECT 281.400 675.300 282.600 677.400 ;
        RECT 283.800 678.300 285.600 683.400 ;
        RECT 289.800 678.300 291.600 683.400 ;
        RECT 283.800 676.950 291.600 678.300 ;
        RECT 298.200 676.200 300.000 683.400 ;
        RECT 296.400 675.300 300.000 676.200 ;
        RECT 281.400 674.250 285.150 675.300 ;
        RECT 283.950 670.950 285.150 674.250 ;
        RECT 287.100 672.150 288.900 673.950 ;
        RECT 272.100 669.150 273.900 670.950 ;
        RECT 268.950 665.850 271.050 667.950 ;
        RECT 271.950 667.050 274.050 669.150 ;
        RECT 283.950 668.850 286.050 670.950 ;
        RECT 286.950 670.050 289.050 672.150 ;
        RECT 289.950 668.850 292.050 670.950 ;
        RECT 293.100 669.150 294.900 670.950 ;
        RECT 280.950 665.850 283.050 667.950 ;
        RECT 253.950 664.050 255.750 665.850 ;
        RECT 256.950 662.850 259.050 664.950 ;
        RECT 260.100 664.050 261.900 665.850 ;
        RECT 257.100 661.050 258.900 662.850 ;
        RECT 251.700 657.900 258.300 658.800 ;
        RECT 251.700 657.600 252.600 657.900 ;
        RECT 233.400 651.600 241.200 652.500 ;
        RECT 250.800 651.600 252.600 657.600 ;
        RECT 256.800 657.600 258.300 657.900 ;
        RECT 269.400 657.600 270.600 665.850 ;
        RECT 281.250 664.050 283.050 665.850 ;
        RECT 284.850 663.600 286.050 668.850 ;
        RECT 290.100 667.050 291.900 668.850 ;
        RECT 292.950 667.050 295.050 669.150 ;
        RECT 296.400 667.950 297.600 675.300 ;
        RECT 311.100 675.000 312.900 683.400 ;
        RECT 324.000 676.200 325.800 683.400 ;
        RECT 342.000 677.400 343.800 683.400 ;
        RECT 352.800 677.400 354.600 683.400 ;
        RECT 324.000 675.300 327.600 676.200 ;
        RECT 308.700 673.350 312.900 675.000 ;
        RECT 299.100 669.150 300.900 670.950 ;
        RECT 308.700 669.150 309.600 673.350 ;
        RECT 323.100 669.150 324.900 670.950 ;
        RECT 295.950 665.850 298.050 667.950 ;
        RECT 298.950 667.050 301.050 669.150 ;
        RECT 307.950 667.050 310.050 669.150 ;
        RECT 256.800 651.600 258.600 657.600 ;
        RECT 268.800 651.600 270.600 657.600 ;
        RECT 284.700 651.600 286.500 663.600 ;
        RECT 296.400 657.600 297.600 665.850 ;
        RECT 308.700 658.800 309.600 667.050 ;
        RECT 310.950 665.850 313.050 667.950 ;
        RECT 316.950 665.850 319.050 667.950 ;
        RECT 322.950 667.050 325.050 669.150 ;
        RECT 326.400 667.950 327.600 675.300 ;
        RECT 338.250 672.150 340.050 673.950 ;
        RECT 329.100 669.150 330.900 670.950 ;
        RECT 325.950 665.850 328.050 667.950 ;
        RECT 328.950 667.050 331.050 669.150 ;
        RECT 334.950 668.850 337.050 670.950 ;
        RECT 337.950 670.050 340.050 672.150 ;
        RECT 342.000 670.950 343.050 677.400 ;
        RECT 353.400 675.300 354.600 677.400 ;
        RECT 355.800 678.300 357.600 683.400 ;
        RECT 361.800 678.300 363.600 683.400 ;
        RECT 355.800 676.950 363.600 678.300 ;
        RECT 370.200 676.200 372.000 683.400 ;
        RECT 383.400 680.400 385.200 683.400 ;
        RECT 395.400 680.400 397.200 683.400 ;
        RECT 368.400 675.300 372.000 676.200 ;
        RECT 353.400 674.250 357.150 675.300 ;
        RECT 340.950 668.850 343.050 670.950 ;
        RECT 343.950 672.150 345.750 673.950 ;
        RECT 343.950 670.050 346.050 672.150 ;
        RECT 355.950 670.950 357.150 674.250 ;
        RECT 359.100 672.150 360.900 673.950 ;
        RECT 346.950 668.850 349.050 670.950 ;
        RECT 355.950 668.850 358.050 670.950 ;
        RECT 358.950 670.050 361.050 672.150 ;
        RECT 361.950 668.850 364.050 670.950 ;
        RECT 365.100 669.150 366.900 670.950 ;
        RECT 335.100 667.050 336.900 668.850 ;
        RECT 310.950 664.050 312.750 665.850 ;
        RECT 313.950 662.850 316.050 664.950 ;
        RECT 317.100 664.050 318.900 665.850 ;
        RECT 314.100 661.050 315.900 662.850 ;
        RECT 308.700 657.900 315.300 658.800 ;
        RECT 308.700 657.600 309.600 657.900 ;
        RECT 296.400 651.600 298.200 657.600 ;
        RECT 307.800 651.600 309.600 657.600 ;
        RECT 313.800 657.600 315.300 657.900 ;
        RECT 326.400 657.600 327.600 665.850 ;
        RECT 340.950 665.400 341.850 668.850 ;
        RECT 346.950 667.050 348.750 668.850 ;
        RECT 352.950 665.850 355.050 667.950 ;
        RECT 337.800 664.500 341.850 665.400 ;
        RECT 313.800 651.600 315.600 657.600 ;
        RECT 325.800 651.600 327.600 657.600 ;
        RECT 334.800 652.500 336.600 663.600 ;
        RECT 337.800 653.400 339.600 664.500 ;
        RECT 353.250 664.050 355.050 665.850 ;
        RECT 356.850 663.600 358.050 668.850 ;
        RECT 362.100 667.050 363.900 668.850 ;
        RECT 364.950 667.050 367.050 669.150 ;
        RECT 368.400 667.950 369.600 675.300 ;
        RECT 384.000 673.950 385.050 680.400 ;
        RECT 382.950 671.850 385.050 673.950 ;
        RECT 391.950 671.850 394.050 673.950 ;
        RECT 395.400 672.150 396.600 680.400 ;
        RECT 409.200 676.200 411.000 683.400 ;
        RECT 407.400 675.300 411.000 676.200 ;
        RECT 419.400 680.400 421.200 683.400 ;
        RECT 371.100 669.150 372.900 670.950 ;
        RECT 367.950 665.850 370.050 667.950 ;
        RECT 370.950 667.050 373.050 669.150 ;
        RECT 379.950 668.850 382.050 670.950 ;
        RECT 380.100 667.050 381.900 668.850 ;
        RECT 340.800 662.400 348.600 663.300 ;
        RECT 340.800 652.500 342.600 662.400 ;
        RECT 334.800 651.600 342.600 652.500 ;
        RECT 346.800 651.600 348.600 662.400 ;
        RECT 356.700 651.600 358.500 663.600 ;
        RECT 368.400 657.600 369.600 665.850 ;
        RECT 384.000 664.650 385.050 671.850 ;
        RECT 385.950 668.850 388.050 670.950 ;
        RECT 392.100 670.050 393.900 671.850 ;
        RECT 394.950 670.050 397.050 672.150 ;
        RECT 386.100 667.050 387.900 668.850 ;
        RECT 384.000 663.600 386.400 664.650 ;
        RECT 368.400 651.600 370.200 657.600 ;
        RECT 384.600 651.600 386.400 663.600 ;
        RECT 395.400 657.600 396.600 670.050 ;
        RECT 404.100 669.150 405.900 670.950 ;
        RECT 403.950 667.050 406.050 669.150 ;
        RECT 407.400 667.950 408.600 675.300 ;
        RECT 415.950 671.850 418.050 673.950 ;
        RECT 419.400 672.150 420.600 680.400 ;
        RECT 429.000 676.200 430.800 683.400 ;
        RECT 440.400 680.400 442.200 683.400 ;
        RECT 429.000 675.300 432.600 676.200 ;
        RECT 410.100 669.150 411.900 670.950 ;
        RECT 416.100 670.050 417.900 671.850 ;
        RECT 418.950 670.050 421.050 672.150 ;
        RECT 406.950 665.850 409.050 667.950 ;
        RECT 409.950 667.050 412.050 669.150 ;
        RECT 407.400 657.600 408.600 665.850 ;
        RECT 419.400 657.600 420.600 670.050 ;
        RECT 428.100 669.150 429.900 670.950 ;
        RECT 427.950 667.050 430.050 669.150 ;
        RECT 431.400 667.950 432.600 675.300 ;
        RECT 436.950 671.850 439.050 673.950 ;
        RECT 440.400 672.150 441.600 680.400 ;
        RECT 451.800 677.400 453.600 683.400 ;
        RECT 452.400 675.300 453.600 677.400 ;
        RECT 454.800 678.300 456.600 683.400 ;
        RECT 460.800 678.300 462.600 683.400 ;
        RECT 454.800 676.950 462.600 678.300 ;
        RECT 464.550 677.400 466.350 683.400 ;
        RECT 472.650 680.400 474.450 683.400 ;
        RECT 480.450 680.400 482.250 683.400 ;
        RECT 488.250 681.300 490.050 683.400 ;
        RECT 488.250 680.400 492.000 681.300 ;
        RECT 472.650 679.500 473.700 680.400 ;
        RECT 469.950 678.300 473.700 679.500 ;
        RECT 481.200 678.600 482.250 680.400 ;
        RECT 490.950 679.500 492.000 680.400 ;
        RECT 469.950 677.400 472.050 678.300 ;
        RECT 452.400 674.250 456.150 675.300 ;
        RECT 434.100 669.150 435.900 670.950 ;
        RECT 437.100 670.050 438.900 671.850 ;
        RECT 439.950 670.050 442.050 672.150 ;
        RECT 454.950 670.950 456.150 674.250 ;
        RECT 464.550 675.150 465.750 677.400 ;
        RECT 477.150 676.200 478.950 678.000 ;
        RECT 481.200 677.550 486.150 678.600 ;
        RECT 484.350 676.800 486.150 677.550 ;
        RECT 487.650 676.800 489.450 678.600 ;
        RECT 490.950 677.400 493.050 679.500 ;
        RECT 496.050 677.400 497.850 683.400 ;
        RECT 478.050 675.900 478.950 676.200 ;
        RECT 488.100 675.900 489.150 676.800 ;
        RECT 458.100 672.150 459.900 673.950 ;
        RECT 464.550 673.050 469.050 675.150 ;
        RECT 478.050 675.000 489.150 675.900 ;
        RECT 430.950 665.850 433.050 667.950 ;
        RECT 433.950 667.050 436.050 669.150 ;
        RECT 431.400 657.600 432.600 665.850 ;
        RECT 395.400 651.600 397.200 657.600 ;
        RECT 407.400 651.600 409.200 657.600 ;
        RECT 419.400 651.600 421.200 657.600 ;
        RECT 430.800 651.600 432.600 657.600 ;
        RECT 440.400 657.600 441.600 670.050 ;
        RECT 454.950 668.850 457.050 670.950 ;
        RECT 457.950 670.050 460.050 672.150 ;
        RECT 460.950 668.850 463.050 670.950 ;
        RECT 451.950 665.850 454.050 667.950 ;
        RECT 452.250 664.050 454.050 665.850 ;
        RECT 455.850 663.600 457.050 668.850 ;
        RECT 461.100 667.050 462.900 668.850 ;
        RECT 464.550 663.600 465.750 673.050 ;
        RECT 466.950 671.250 470.850 673.050 ;
        RECT 466.950 670.950 469.050 671.250 ;
        RECT 478.050 670.950 478.950 675.000 ;
        RECT 488.100 673.800 489.150 675.000 ;
        RECT 488.100 672.600 495.000 673.800 ;
        RECT 488.100 672.000 489.900 672.600 ;
        RECT 494.100 671.850 495.000 672.600 ;
        RECT 491.100 670.950 492.900 671.700 ;
        RECT 478.050 668.850 481.050 670.950 ;
        RECT 484.950 669.900 492.900 670.950 ;
        RECT 494.100 670.050 495.900 671.850 ;
        RECT 484.950 668.850 487.050 669.900 ;
        RECT 466.950 665.400 468.750 667.200 ;
        RECT 467.850 664.200 472.050 665.400 ;
        RECT 478.050 664.200 478.950 668.850 ;
        RECT 486.750 665.100 488.550 665.400 ;
        RECT 440.400 651.600 442.200 657.600 ;
        RECT 455.700 651.600 457.500 663.600 ;
        RECT 464.550 651.600 466.350 663.600 ;
        RECT 469.950 663.300 472.050 664.200 ;
        RECT 472.950 663.300 478.950 664.200 ;
        RECT 480.150 664.800 488.550 665.100 ;
        RECT 496.950 664.800 497.850 677.400 ;
        RECT 500.400 678.300 502.200 683.400 ;
        RECT 506.400 678.300 508.200 683.400 ;
        RECT 500.400 676.950 508.200 678.300 ;
        RECT 509.400 677.400 511.200 683.400 ;
        RECT 509.400 675.300 510.600 677.400 ;
        RECT 520.200 676.200 522.000 683.400 ;
        RECT 506.850 674.250 510.600 675.300 ;
        RECT 518.400 675.300 522.000 676.200 ;
        RECT 530.400 680.400 532.200 683.400 ;
        RECT 503.100 672.150 504.900 673.950 ;
        RECT 499.950 668.850 502.050 670.950 ;
        RECT 502.950 670.050 505.050 672.150 ;
        RECT 506.850 670.950 508.050 674.250 ;
        RECT 505.950 668.850 508.050 670.950 ;
        RECT 515.100 669.150 516.900 670.950 ;
        RECT 500.100 667.050 501.900 668.850 ;
        RECT 480.150 664.200 497.850 664.800 ;
        RECT 472.950 662.400 473.850 663.300 ;
        RECT 471.150 660.600 473.850 662.400 ;
        RECT 474.750 662.100 476.550 662.400 ;
        RECT 480.150 662.100 481.050 664.200 ;
        RECT 486.750 663.600 497.850 664.200 ;
        RECT 505.950 663.600 507.150 668.850 ;
        RECT 508.950 665.850 511.050 667.950 ;
        RECT 514.950 667.050 517.050 669.150 ;
        RECT 518.400 667.950 519.600 675.300 ;
        RECT 526.950 671.850 529.050 673.950 ;
        RECT 530.400 672.150 531.600 680.400 ;
        RECT 536.400 678.300 538.200 683.400 ;
        RECT 542.400 678.300 544.200 683.400 ;
        RECT 536.400 676.950 544.200 678.300 ;
        RECT 545.400 677.400 547.200 683.400 ;
        RECT 545.400 675.300 546.600 677.400 ;
        RECT 555.000 676.200 556.800 683.400 ;
        RECT 564.150 677.400 565.950 683.400 ;
        RECT 571.950 681.300 573.750 683.400 ;
        RECT 570.000 680.400 573.750 681.300 ;
        RECT 579.750 680.400 581.550 683.400 ;
        RECT 587.550 680.400 589.350 683.400 ;
        RECT 570.000 679.500 571.050 680.400 ;
        RECT 568.950 677.400 571.050 679.500 ;
        RECT 579.750 678.600 580.800 680.400 ;
        RECT 555.000 675.300 558.600 676.200 ;
        RECT 542.850 674.250 546.600 675.300 ;
        RECT 539.100 672.150 540.900 673.950 ;
        RECT 521.100 669.150 522.900 670.950 ;
        RECT 527.100 670.050 528.900 671.850 ;
        RECT 529.950 670.050 532.050 672.150 ;
        RECT 517.950 665.850 520.050 667.950 ;
        RECT 520.950 667.050 523.050 669.150 ;
        RECT 508.950 664.050 510.750 665.850 ;
        RECT 474.750 661.200 481.050 662.100 ;
        RECT 481.950 662.700 483.750 663.300 ;
        RECT 481.950 661.500 489.450 662.700 ;
        RECT 474.750 660.600 476.550 661.200 ;
        RECT 488.250 660.600 489.450 661.500 ;
        RECT 469.950 657.600 473.850 659.700 ;
        RECT 478.950 659.550 480.750 660.300 ;
        RECT 483.750 659.550 485.550 660.300 ;
        RECT 478.950 658.500 485.550 659.550 ;
        RECT 488.250 658.500 493.050 660.600 ;
        RECT 472.050 651.600 473.850 657.600 ;
        RECT 479.850 651.600 481.650 658.500 ;
        RECT 488.250 657.600 489.450 658.500 ;
        RECT 487.650 651.600 489.450 657.600 ;
        RECT 496.050 651.600 497.850 663.600 ;
        RECT 505.500 651.600 507.300 663.600 ;
        RECT 518.400 657.600 519.600 665.850 ;
        RECT 530.400 657.600 531.600 670.050 ;
        RECT 535.950 668.850 538.050 670.950 ;
        RECT 538.950 670.050 541.050 672.150 ;
        RECT 542.850 670.950 544.050 674.250 ;
        RECT 541.950 668.850 544.050 670.950 ;
        RECT 554.100 669.150 555.900 670.950 ;
        RECT 536.100 667.050 537.900 668.850 ;
        RECT 541.950 663.600 543.150 668.850 ;
        RECT 544.950 665.850 547.050 667.950 ;
        RECT 553.950 667.050 556.050 669.150 ;
        RECT 557.400 667.950 558.600 675.300 ;
        RECT 560.100 669.150 561.900 670.950 ;
        RECT 556.950 665.850 559.050 667.950 ;
        RECT 559.950 667.050 562.050 669.150 ;
        RECT 544.950 664.050 546.750 665.850 ;
        RECT 518.400 651.600 520.200 657.600 ;
        RECT 530.400 651.600 532.200 657.600 ;
        RECT 541.500 651.600 543.300 663.600 ;
        RECT 557.400 657.600 558.600 665.850 ;
        RECT 556.800 651.600 558.600 657.600 ;
        RECT 564.150 664.800 565.050 677.400 ;
        RECT 572.550 676.800 574.350 678.600 ;
        RECT 575.850 677.550 580.800 678.600 ;
        RECT 588.300 679.500 589.350 680.400 ;
        RECT 588.300 678.300 592.050 679.500 ;
        RECT 575.850 676.800 577.650 677.550 ;
        RECT 572.850 675.900 573.900 676.800 ;
        RECT 583.050 676.200 584.850 678.000 ;
        RECT 589.950 677.400 592.050 678.300 ;
        RECT 595.650 677.400 597.450 683.400 ;
        RECT 583.050 675.900 583.950 676.200 ;
        RECT 572.850 675.000 583.950 675.900 ;
        RECT 596.250 675.150 597.450 677.400 ;
        RECT 603.000 676.200 604.800 683.400 ;
        RECT 616.200 680.400 618.000 683.400 ;
        RECT 603.000 675.300 606.600 676.200 ;
        RECT 572.850 673.800 573.900 675.000 ;
        RECT 567.000 672.600 573.900 673.800 ;
        RECT 567.000 671.850 567.900 672.600 ;
        RECT 572.100 672.000 573.900 672.600 ;
        RECT 566.100 670.050 567.900 671.850 ;
        RECT 569.100 670.950 570.900 671.700 ;
        RECT 583.050 670.950 583.950 675.000 ;
        RECT 592.950 673.050 597.450 675.150 ;
        RECT 591.150 671.250 595.050 673.050 ;
        RECT 592.950 670.950 595.050 671.250 ;
        RECT 569.100 669.900 577.050 670.950 ;
        RECT 574.950 668.850 577.050 669.900 ;
        RECT 580.950 668.850 583.950 670.950 ;
        RECT 573.450 665.100 575.250 665.400 ;
        RECT 573.450 664.800 581.850 665.100 ;
        RECT 564.150 664.200 581.850 664.800 ;
        RECT 564.150 663.600 575.250 664.200 ;
        RECT 564.150 651.600 565.950 663.600 ;
        RECT 578.250 662.700 580.050 663.300 ;
        RECT 572.550 661.500 580.050 662.700 ;
        RECT 580.950 662.100 581.850 664.200 ;
        RECT 583.050 664.200 583.950 668.850 ;
        RECT 593.250 665.400 595.050 667.200 ;
        RECT 589.950 664.200 594.150 665.400 ;
        RECT 583.050 663.300 589.050 664.200 ;
        RECT 589.950 663.300 592.050 664.200 ;
        RECT 596.250 663.600 597.450 673.050 ;
        RECT 602.100 669.150 603.900 670.950 ;
        RECT 601.950 667.050 604.050 669.150 ;
        RECT 605.400 667.950 606.600 675.300 ;
        RECT 616.500 672.150 618.000 680.400 ;
        RECT 608.100 669.150 609.900 670.950 ;
        RECT 613.950 670.050 618.000 672.150 ;
        RECT 604.950 665.850 607.050 667.950 ;
        RECT 607.950 667.050 610.050 669.150 ;
        RECT 588.150 662.400 589.050 663.300 ;
        RECT 585.450 662.100 587.250 662.400 ;
        RECT 572.550 660.600 573.750 661.500 ;
        RECT 580.950 661.200 587.250 662.100 ;
        RECT 585.450 660.600 587.250 661.200 ;
        RECT 588.150 660.600 590.850 662.400 ;
        RECT 568.950 658.500 573.750 660.600 ;
        RECT 576.450 659.550 578.250 660.300 ;
        RECT 581.250 659.550 583.050 660.300 ;
        RECT 576.450 658.500 583.050 659.550 ;
        RECT 572.550 657.600 573.750 658.500 ;
        RECT 572.550 651.600 574.350 657.600 ;
        RECT 580.350 651.600 582.150 658.500 ;
        RECT 588.150 657.600 592.050 659.700 ;
        RECT 588.150 651.600 589.950 657.600 ;
        RECT 595.650 651.600 597.450 663.600 ;
        RECT 605.400 657.600 606.600 665.850 ;
        RECT 616.500 657.600 618.000 670.050 ;
        RECT 620.100 677.400 621.900 683.400 ;
        RECT 630.600 678.600 632.400 683.400 ;
        RECT 635.400 680.400 637.200 683.400 ;
        RECT 638.400 680.400 640.200 683.400 ;
        RECT 641.400 680.400 643.200 683.400 ;
        RECT 645.000 680.400 646.800 683.400 ;
        RECT 635.400 679.500 636.750 680.400 ;
        RECT 638.400 679.500 640.050 680.400 ;
        RECT 641.400 679.500 643.050 680.400 ;
        RECT 628.200 677.400 632.400 678.600 ;
        RECT 634.950 677.400 637.050 679.500 ;
        RECT 637.950 677.400 640.050 679.500 ;
        RECT 640.950 677.400 643.050 679.500 ;
        RECT 645.750 679.500 646.800 680.400 ;
        RECT 651.000 680.400 652.800 683.400 ;
        RECT 658.500 680.400 660.300 683.400 ;
        RECT 661.500 680.400 663.300 683.400 ;
        RECT 664.500 680.400 666.300 683.400 ;
        RECT 651.000 679.500 652.050 680.400 ;
        RECT 645.750 677.400 647.850 679.500 ;
        RECT 649.950 677.400 652.050 679.500 ;
        RECT 653.700 678.750 655.500 679.200 ;
        RECT 658.950 679.050 660.300 680.400 ;
        RECT 661.950 679.050 663.300 680.400 ;
        RECT 664.950 679.050 666.300 680.400 ;
        RECT 653.700 677.400 657.750 678.750 ;
        RECT 620.100 662.550 621.000 677.400 ;
        RECT 628.200 673.800 629.700 677.400 ;
        RECT 634.500 674.700 641.100 676.500 ;
        RECT 642.000 674.700 648.900 676.500 ;
        RECT 656.850 676.050 657.750 677.400 ;
        RECT 658.950 676.950 661.050 679.050 ;
        RECT 661.950 676.950 664.050 679.050 ;
        RECT 664.950 676.950 667.050 679.050 ;
        RECT 656.850 675.900 661.950 676.050 ;
        RECT 656.850 675.150 664.500 675.900 ;
        RECT 660.150 674.700 664.500 675.150 ;
        RECT 642.000 673.800 643.050 674.700 ;
        RECT 660.150 674.250 661.950 674.700 ;
        RECT 621.900 672.300 629.700 673.800 ;
        RECT 633.150 672.750 643.050 673.800 ;
        RECT 621.900 672.000 623.700 672.300 ;
        RECT 626.700 672.000 628.500 672.300 ;
        RECT 633.150 670.950 634.200 672.750 ;
        RECT 643.950 672.450 651.600 673.800 ;
        RECT 643.950 671.700 644.850 672.450 ;
        RECT 625.950 669.900 634.200 670.950 ;
        RECT 635.250 670.650 644.850 671.700 ;
        RECT 625.950 665.850 628.050 669.900 ;
        RECT 635.250 669.000 636.150 670.650 ;
        RECT 645.750 669.750 649.650 671.550 ;
        RECT 650.550 670.950 651.600 672.450 ;
        RECT 652.950 673.650 655.050 673.950 ;
        RECT 652.950 671.850 656.850 673.650 ;
        RECT 663.450 671.250 664.500 674.700 ;
        RECT 666.000 673.800 667.050 676.950 ;
        RECT 668.700 677.400 670.500 683.400 ;
        RECT 679.500 677.400 681.300 683.400 ;
        RECT 668.700 676.500 670.200 677.400 ;
        RECT 668.700 675.300 677.100 676.500 ;
        RECT 675.300 674.700 677.100 675.300 ;
        RECT 680.100 673.800 681.300 677.400 ;
        RECT 691.200 676.200 693.000 683.400 ;
        RECT 700.800 677.400 702.600 683.400 ;
        RECT 666.000 672.900 681.300 673.800 ;
        RECT 650.550 670.050 662.550 670.950 ;
        RECT 629.100 667.200 636.150 669.000 ;
        RECT 637.500 667.950 639.300 669.750 ;
        RECT 645.750 669.450 647.850 669.750 ;
        RECT 649.950 668.550 652.050 668.850 ;
        RECT 658.800 668.550 660.600 669.150 ;
        RECT 649.950 667.950 660.600 668.550 ;
        RECT 637.500 667.500 660.600 667.950 ;
        RECT 661.500 668.550 662.550 670.050 ;
        RECT 663.450 669.450 665.250 671.250 ;
        RECT 667.050 670.950 678.900 672.000 ;
        RECT 667.050 668.550 668.250 670.950 ;
        RECT 677.100 669.150 678.900 670.950 ;
        RECT 661.500 667.650 668.250 668.550 ;
        RECT 670.950 667.650 673.050 667.950 ;
        RECT 637.500 666.750 652.050 667.500 ;
        RECT 658.800 667.350 660.600 667.500 ;
        RECT 669.150 666.450 673.050 667.650 ;
        RECT 676.950 667.050 679.050 669.150 ;
        RECT 659.100 665.850 673.050 666.450 ;
        RECT 633.000 665.550 673.050 665.850 ;
        RECT 621.900 664.650 623.700 665.250 ;
        RECT 633.000 664.650 661.050 665.550 ;
        RECT 621.900 663.450 634.050 664.650 ;
        RECT 661.950 664.050 664.050 664.350 ;
        RECT 671.700 664.050 673.500 664.650 ;
        RECT 634.950 662.550 637.050 663.750 ;
        RECT 620.100 661.650 637.050 662.550 ;
        RECT 640.950 662.700 661.050 663.750 ;
        RECT 640.950 661.650 643.050 662.700 ;
        RECT 604.800 651.600 606.600 657.600 ;
        RECT 616.200 651.600 618.000 657.600 ;
        RECT 622.800 657.600 624.000 661.650 ;
        RECT 624.900 659.700 626.700 660.300 ;
        RECT 631.500 660.150 633.300 660.300 ;
        RECT 624.900 658.500 630.600 659.700 ;
        RECT 631.500 658.950 640.050 660.150 ;
        RECT 631.500 658.500 633.300 658.950 ;
        RECT 622.800 651.600 624.600 657.600 ;
        RECT 628.800 651.600 630.600 658.500 ;
        RECT 637.950 658.050 640.050 658.950 ;
        RECT 634.950 655.800 637.050 657.900 ;
        RECT 635.850 654.600 637.050 655.800 ;
        RECT 638.400 654.600 640.050 658.050 ;
        RECT 641.850 654.600 643.050 661.650 ;
        RECT 659.100 661.350 661.050 662.700 ;
        RECT 661.950 662.850 673.500 664.050 ;
        RECT 661.950 662.250 664.050 662.850 ;
        RECT 675.000 661.350 676.800 662.100 ;
        RECT 644.100 658.800 648.000 660.600 ;
        RECT 645.000 658.500 648.000 658.800 ;
        RECT 649.950 658.500 652.050 660.600 ;
        RECT 659.100 660.300 676.800 661.350 ;
        RECT 635.400 651.600 637.200 654.600 ;
        RECT 638.400 651.600 640.200 654.600 ;
        RECT 641.400 651.600 643.200 654.600 ;
        RECT 645.000 651.600 646.800 658.500 ;
        RECT 651.000 657.600 652.050 658.500 ;
        RECT 651.000 651.600 652.800 657.600 ;
        RECT 658.650 655.950 661.050 658.050 ;
        RECT 661.950 655.950 664.050 658.050 ;
        RECT 664.950 655.950 667.050 658.050 ;
        RECT 658.650 654.600 659.850 655.950 ;
        RECT 661.950 654.600 663.000 655.950 ;
        RECT 665.250 654.600 666.150 655.950 ;
        RECT 657.900 651.600 659.850 654.600 ;
        RECT 660.900 651.600 663.000 654.600 ;
        RECT 663.900 651.600 666.150 654.600 ;
        RECT 670.500 651.600 672.300 660.300 ;
        RECT 680.100 659.400 681.300 672.900 ;
        RECT 689.400 675.300 693.000 676.200 ;
        RECT 701.400 675.300 702.600 677.400 ;
        RECT 703.800 678.300 705.600 683.400 ;
        RECT 709.800 678.300 711.600 683.400 ;
        RECT 721.800 680.400 723.600 683.400 ;
        RECT 703.800 676.950 711.600 678.300 ;
        RECT 686.100 669.150 687.900 670.950 ;
        RECT 685.950 667.050 688.050 669.150 ;
        RECT 689.400 667.950 690.600 675.300 ;
        RECT 701.400 674.250 705.150 675.300 ;
        RECT 703.950 670.950 705.150 674.250 ;
        RECT 721.950 673.950 723.000 680.400 ;
        RECT 734.100 675.000 735.900 683.400 ;
        RECT 707.100 672.150 708.900 673.950 ;
        RECT 692.100 669.150 693.900 670.950 ;
        RECT 688.950 665.850 691.050 667.950 ;
        RECT 691.950 667.050 694.050 669.150 ;
        RECT 703.950 668.850 706.050 670.950 ;
        RECT 706.950 670.050 709.050 672.150 ;
        RECT 721.950 671.850 724.050 673.950 ;
        RECT 731.700 673.350 735.900 675.000 ;
        RECT 749.400 680.400 751.200 683.400 ;
        RECT 758.400 680.400 760.200 683.400 ;
        RECT 709.950 668.850 712.050 670.950 ;
        RECT 718.950 668.850 721.050 670.950 ;
        RECT 700.950 665.850 703.050 667.950 ;
        RECT 677.250 658.500 681.300 659.400 ;
        RECT 677.250 657.600 678.300 658.500 ;
        RECT 676.500 651.600 678.300 657.600 ;
        RECT 689.400 657.600 690.600 665.850 ;
        RECT 701.250 664.050 703.050 665.850 ;
        RECT 704.850 663.600 706.050 668.850 ;
        RECT 710.100 667.050 711.900 668.850 ;
        RECT 719.100 667.050 720.900 668.850 ;
        RECT 721.950 664.650 723.000 671.850 ;
        RECT 724.950 668.850 727.050 670.950 ;
        RECT 731.700 669.150 732.600 673.350 ;
        RECT 745.950 671.850 748.050 673.950 ;
        RECT 749.400 672.150 750.600 680.400 ;
        RECT 746.100 670.050 747.900 671.850 ;
        RECT 748.950 670.050 751.050 672.150 ;
        RECT 754.950 671.850 757.050 673.950 ;
        RECT 758.400 672.150 759.600 680.400 ;
        RECT 755.100 670.050 756.900 671.850 ;
        RECT 757.950 670.050 760.050 672.150 ;
        RECT 725.100 667.050 726.900 668.850 ;
        RECT 730.950 667.050 733.050 669.150 ;
        RECT 720.600 663.600 723.000 664.650 ;
        RECT 689.400 651.600 691.200 657.600 ;
        RECT 704.700 651.600 706.500 663.600 ;
        RECT 720.600 651.600 722.400 663.600 ;
        RECT 731.700 658.800 732.600 667.050 ;
        RECT 733.950 665.850 736.050 667.950 ;
        RECT 739.950 665.850 742.050 667.950 ;
        RECT 733.950 664.050 735.750 665.850 ;
        RECT 736.950 662.850 739.050 664.950 ;
        RECT 740.100 664.050 741.900 665.850 ;
        RECT 737.100 661.050 738.900 662.850 ;
        RECT 731.700 657.900 738.300 658.800 ;
        RECT 731.700 657.600 732.600 657.900 ;
        RECT 730.800 651.600 732.600 657.600 ;
        RECT 736.800 657.600 738.300 657.900 ;
        RECT 749.400 657.600 750.600 670.050 ;
        RECT 758.400 657.600 759.600 670.050 ;
        RECT 736.800 651.600 738.600 657.600 ;
        RECT 749.400 651.600 751.200 657.600 ;
        RECT 758.400 651.600 760.200 657.600 ;
        RECT 6.600 635.400 8.400 647.400 ;
        RECT 17.400 641.400 19.200 647.400 ;
        RECT 6.600 634.350 9.000 635.400 ;
        RECT 5.100 630.150 6.900 631.950 ;
        RECT 4.950 628.050 7.050 630.150 ;
        RECT 7.950 627.150 9.000 634.350 ;
        RECT 11.100 630.150 12.900 631.950 ;
        RECT 14.100 630.150 15.900 631.950 ;
        RECT 10.950 628.050 13.050 630.150 ;
        RECT 13.950 628.050 16.050 630.150 ;
        RECT 7.950 625.050 10.050 627.150 ;
        RECT 7.950 618.600 9.000 625.050 ;
        RECT 17.550 624.300 18.600 641.400 ;
        RECT 24.000 635.400 25.800 647.400 ;
        RECT 34.800 641.400 36.600 647.400 ;
        RECT 44.400 641.400 46.200 647.400 ;
        RECT 19.950 629.850 22.050 631.950 ;
        RECT 24.000 630.150 25.050 635.400 ;
        RECT 35.400 633.150 36.600 641.400 ;
        RECT 44.700 641.100 46.200 641.400 ;
        RECT 50.400 641.400 52.200 647.400 ;
        RECT 62.400 641.400 64.200 647.400 ;
        RECT 50.400 641.100 51.300 641.400 ;
        RECT 44.700 640.200 51.300 641.100 ;
        RECT 44.100 636.150 45.900 637.950 ;
        RECT 41.100 633.150 42.900 634.950 ;
        RECT 43.950 634.050 46.050 636.150 ;
        RECT 47.250 633.150 49.050 634.950 ;
        RECT 20.100 628.050 21.900 629.850 ;
        RECT 22.950 628.050 25.050 630.150 ;
        RECT 31.950 629.850 34.050 631.950 ;
        RECT 34.950 631.050 37.050 633.150 ;
        RECT 32.100 628.050 33.900 629.850 ;
        RECT 14.400 623.100 21.900 624.300 ;
        RECT 7.800 615.600 9.600 618.600 ;
        RECT 14.400 615.600 16.200 623.100 ;
        RECT 20.100 622.500 21.900 623.100 ;
        RECT 24.000 621.600 25.050 628.050 ;
        RECT 35.400 623.700 36.600 631.050 ;
        RECT 37.950 629.850 40.050 631.950 ;
        RECT 40.950 631.050 43.050 633.150 ;
        RECT 46.950 631.050 49.050 633.150 ;
        RECT 50.400 631.950 51.300 640.200 ;
        RECT 49.950 629.850 52.050 631.950 ;
        RECT 38.100 628.050 39.900 629.850 ;
        RECT 50.400 625.650 51.300 629.850 ;
        RECT 62.400 628.950 63.600 641.400 ;
        RECT 68.400 636.300 70.200 647.400 ;
        RECT 74.400 636.300 76.200 647.400 ;
        RECT 68.400 635.400 76.200 636.300 ;
        RECT 77.400 635.400 79.200 647.400 ;
        RECT 85.800 641.400 87.600 647.400 ;
        RECT 77.700 630.150 78.600 635.400 ;
        RECT 59.100 627.150 60.900 628.950 ;
        RECT 21.900 620.100 25.050 621.600 ;
        RECT 33.000 622.800 36.600 623.700 ;
        RECT 47.100 624.000 51.300 625.650 ;
        RECT 58.950 625.050 61.050 627.150 ;
        RECT 61.950 626.850 64.050 628.950 ;
        RECT 67.950 626.850 70.050 628.950 ;
        RECT 71.100 627.150 72.900 628.950 ;
        RECT 21.900 615.600 23.700 620.100 ;
        RECT 33.000 615.600 34.800 622.800 ;
        RECT 47.100 615.600 48.900 624.000 ;
        RECT 62.400 618.600 63.600 626.850 ;
        RECT 68.100 625.050 69.900 626.850 ;
        RECT 70.950 625.050 73.050 627.150 ;
        RECT 73.950 626.850 76.050 628.950 ;
        RECT 76.950 628.050 79.050 630.150 ;
        RECT 86.400 628.950 87.600 641.400 ;
        RECT 98.700 635.400 100.500 647.400 ;
        RECT 113.700 635.400 115.500 647.400 ;
        RECT 124.800 635.400 126.600 647.400 ;
        RECT 127.800 636.300 129.600 647.400 ;
        RECT 133.800 636.300 135.600 647.400 ;
        RECT 127.800 635.400 135.600 636.300 ;
        RECT 146.700 635.400 148.500 647.400 ;
        RECT 161.700 635.400 163.500 647.400 ;
        RECT 176.700 635.400 178.500 647.400 ;
        RECT 191.400 641.400 193.200 647.400 ;
        RECT 202.800 646.500 210.600 647.400 ;
        RECT 95.250 633.150 97.050 634.950 ;
        RECT 94.950 631.050 97.050 633.150 ;
        RECT 98.850 630.150 100.050 635.400 ;
        RECT 110.250 633.150 112.050 634.950 ;
        RECT 104.100 630.150 105.900 631.950 ;
        RECT 109.950 631.050 112.050 633.150 ;
        RECT 113.850 630.150 115.050 635.400 ;
        RECT 119.100 630.150 120.900 631.950 ;
        RECT 125.400 630.150 126.300 635.400 ;
        RECT 127.950 633.450 130.050 634.050 ;
        RECT 127.950 632.550 138.450 633.450 ;
        RECT 143.250 633.150 145.050 634.950 ;
        RECT 127.950 631.950 130.050 632.550 ;
        RECT 74.100 625.050 75.900 626.850 ;
        RECT 77.700 621.600 78.600 628.050 ;
        RECT 85.950 626.850 88.050 628.950 ;
        RECT 89.100 627.150 90.900 628.950 ;
        RECT 97.950 628.050 100.050 630.150 ;
        RECT 73.200 619.950 78.600 621.600 ;
        RECT 62.400 615.600 64.200 618.600 ;
        RECT 73.200 615.600 75.000 619.950 ;
        RECT 86.400 618.600 87.600 626.850 ;
        RECT 88.950 625.050 91.050 627.150 ;
        RECT 97.950 624.750 99.150 628.050 ;
        RECT 100.950 626.850 103.050 628.950 ;
        RECT 103.950 628.050 106.050 630.150 ;
        RECT 112.950 628.050 115.050 630.150 ;
        RECT 101.100 625.050 102.900 626.850 ;
        RECT 112.950 624.750 114.150 628.050 ;
        RECT 115.950 626.850 118.050 628.950 ;
        RECT 118.950 628.050 121.050 630.150 ;
        RECT 124.950 628.050 127.050 630.150 ;
        RECT 116.100 625.050 117.900 626.850 ;
        RECT 95.400 623.700 99.150 624.750 ;
        RECT 110.400 623.700 114.150 624.750 ;
        RECT 95.400 621.600 96.600 623.700 ;
        RECT 85.800 615.600 87.600 618.600 ;
        RECT 94.800 615.600 96.600 621.600 ;
        RECT 97.800 620.700 105.600 622.050 ;
        RECT 110.400 621.600 111.600 623.700 ;
        RECT 97.800 615.600 99.600 620.700 ;
        RECT 103.800 615.600 105.600 620.700 ;
        RECT 109.800 615.600 111.600 621.600 ;
        RECT 112.800 620.700 120.600 622.050 ;
        RECT 112.800 615.600 114.600 620.700 ;
        RECT 118.800 615.600 120.600 620.700 ;
        RECT 125.400 621.600 126.300 628.050 ;
        RECT 127.950 626.850 130.050 628.950 ;
        RECT 131.100 627.150 132.900 628.950 ;
        RECT 128.100 625.050 129.900 626.850 ;
        RECT 130.950 625.050 133.050 627.150 ;
        RECT 133.950 626.850 136.050 628.950 ;
        RECT 137.550 627.450 138.450 632.550 ;
        RECT 142.950 631.050 145.050 633.150 ;
        RECT 146.850 630.150 148.050 635.400 ;
        RECT 158.250 633.150 160.050 634.950 ;
        RECT 152.100 630.150 153.900 631.950 ;
        RECT 157.950 631.050 160.050 633.150 ;
        RECT 161.850 630.150 163.050 635.400 ;
        RECT 173.250 633.150 175.050 634.950 ;
        RECT 167.100 630.150 168.900 631.950 ;
        RECT 172.950 631.050 175.050 633.150 ;
        RECT 176.850 630.150 178.050 635.400 ;
        RECT 184.950 634.950 187.050 637.050 ;
        RECT 182.100 630.150 183.900 631.950 ;
        RECT 145.950 628.050 148.050 630.150 ;
        RECT 142.950 627.450 145.050 628.050 ;
        RECT 134.100 625.050 135.900 626.850 ;
        RECT 137.550 626.550 145.050 627.450 ;
        RECT 142.950 625.950 145.050 626.550 ;
        RECT 145.950 624.750 147.150 628.050 ;
        RECT 148.950 626.850 151.050 628.950 ;
        RECT 151.950 628.050 154.050 630.150 ;
        RECT 160.950 628.050 163.050 630.150 ;
        RECT 149.100 625.050 150.900 626.850 ;
        RECT 160.950 624.750 162.150 628.050 ;
        RECT 163.950 626.850 166.050 628.950 ;
        RECT 166.950 628.050 169.050 630.150 ;
        RECT 175.950 628.050 178.050 630.150 ;
        RECT 164.100 625.050 165.900 626.850 ;
        RECT 175.950 624.750 177.150 628.050 ;
        RECT 178.950 626.850 181.050 628.950 ;
        RECT 181.950 628.050 184.050 630.150 ;
        RECT 179.100 625.050 180.900 626.850 ;
        RECT 143.400 623.700 147.150 624.750 ;
        RECT 158.400 623.700 162.150 624.750 ;
        RECT 173.400 623.700 177.150 624.750 ;
        RECT 185.550 624.450 186.450 634.950 ;
        RECT 191.400 633.150 192.600 641.400 ;
        RECT 202.800 635.400 204.600 646.500 ;
        RECT 205.800 634.500 207.600 645.600 ;
        RECT 208.800 636.600 210.600 646.500 ;
        RECT 214.800 636.600 216.600 647.400 ;
        RECT 208.800 635.700 216.600 636.600 ;
        RECT 220.200 635.400 222.000 647.400 ;
        RECT 226.800 641.400 228.600 647.400 ;
        RECT 238.800 641.400 240.600 647.400 ;
        RECT 205.800 633.600 209.850 634.500 ;
        RECT 187.950 629.850 190.050 631.950 ;
        RECT 190.950 631.050 193.050 633.150 ;
        RECT 188.100 628.050 189.900 629.850 ;
        RECT 187.950 624.450 190.050 625.050 ;
        RECT 143.400 621.600 144.600 623.700 ;
        RECT 125.400 619.950 130.800 621.600 ;
        RECT 129.000 615.600 130.800 619.950 ;
        RECT 142.800 615.600 144.600 621.600 ;
        RECT 145.800 620.700 153.600 622.050 ;
        RECT 158.400 621.600 159.600 623.700 ;
        RECT 145.800 615.600 147.600 620.700 ;
        RECT 151.800 615.600 153.600 620.700 ;
        RECT 157.800 615.600 159.600 621.600 ;
        RECT 160.800 620.700 168.600 622.050 ;
        RECT 173.400 621.600 174.600 623.700 ;
        RECT 185.550 623.550 190.050 624.450 ;
        RECT 187.950 622.950 190.050 623.550 ;
        RECT 191.400 623.700 192.600 631.050 ;
        RECT 193.950 629.850 196.050 631.950 ;
        RECT 203.100 630.150 204.900 631.950 ;
        RECT 208.950 630.150 209.850 633.600 ;
        RECT 214.950 630.150 216.750 631.950 ;
        RECT 220.950 630.150 222.000 635.400 ;
        RECT 194.100 628.050 195.900 629.850 ;
        RECT 202.950 628.050 205.050 630.150 ;
        RECT 205.950 626.850 208.050 628.950 ;
        RECT 208.950 628.050 211.050 630.150 ;
        RECT 206.250 625.050 208.050 626.850 ;
        RECT 191.400 622.800 195.000 623.700 ;
        RECT 160.800 615.600 162.600 620.700 ;
        RECT 166.800 615.600 168.600 620.700 ;
        RECT 172.800 615.600 174.600 621.600 ;
        RECT 175.800 620.700 183.600 622.050 ;
        RECT 175.800 615.600 177.600 620.700 ;
        RECT 181.800 615.600 183.600 620.700 ;
        RECT 193.200 615.600 195.000 622.800 ;
        RECT 210.000 621.600 211.050 628.050 ;
        RECT 211.950 626.850 214.050 628.950 ;
        RECT 214.950 628.050 217.050 630.150 ;
        RECT 220.950 628.050 223.050 630.150 ;
        RECT 223.950 629.850 226.050 631.950 ;
        RECT 224.100 628.050 225.900 629.850 ;
        RECT 211.950 625.050 213.750 626.850 ;
        RECT 220.950 621.600 222.000 628.050 ;
        RECT 227.400 624.300 228.450 641.400 ;
        RECT 239.400 633.150 240.600 641.400 ;
        RECT 251.700 635.400 253.500 647.400 ;
        RECT 260.400 636.600 262.200 647.400 ;
        RECT 266.400 646.500 274.200 647.400 ;
        RECT 266.400 636.600 268.200 646.500 ;
        RECT 260.400 635.700 268.200 636.600 ;
        RECT 248.250 633.150 250.050 634.950 ;
        RECT 230.100 630.150 231.900 631.950 ;
        RECT 229.950 628.050 232.050 630.150 ;
        RECT 235.950 629.850 238.050 631.950 ;
        RECT 238.950 631.050 241.050 633.150 ;
        RECT 236.100 628.050 237.900 629.850 ;
        RECT 224.100 623.100 231.600 624.300 ;
        RECT 239.400 623.700 240.600 631.050 ;
        RECT 241.950 629.850 244.050 631.950 ;
        RECT 247.950 631.050 250.050 633.150 ;
        RECT 251.850 630.150 253.050 635.400 ;
        RECT 269.400 634.500 271.200 645.600 ;
        RECT 272.400 635.400 274.200 646.500 ;
        RECT 281.400 641.400 283.200 647.400 ;
        RECT 267.150 633.600 271.200 634.500 ;
        RECT 257.100 630.150 258.900 631.950 ;
        RECT 260.250 630.150 262.050 631.950 ;
        RECT 267.150 630.150 268.050 633.600 ;
        RECT 281.400 633.150 282.600 641.400 ;
        RECT 292.800 635.400 294.600 647.400 ;
        RECT 305.700 635.400 307.500 647.400 ;
        RECT 316.800 641.400 318.600 647.400 ;
        RECT 328.800 641.400 330.600 647.400 ;
        RECT 272.100 630.150 273.900 631.950 ;
        RECT 242.100 628.050 243.900 629.850 ;
        RECT 250.950 628.050 253.050 630.150 ;
        RECT 250.950 624.750 252.150 628.050 ;
        RECT 253.950 626.850 256.050 628.950 ;
        RECT 256.950 628.050 259.050 630.150 ;
        RECT 259.950 628.050 262.050 630.150 ;
        RECT 262.950 626.850 265.050 628.950 ;
        RECT 254.100 625.050 255.900 626.850 ;
        RECT 263.250 625.050 265.050 626.850 ;
        RECT 265.950 628.050 268.050 630.150 ;
        RECT 224.100 622.500 225.900 623.100 ;
        RECT 210.000 615.600 211.800 621.600 ;
        RECT 220.950 620.100 224.100 621.600 ;
        RECT 222.300 615.600 224.100 620.100 ;
        RECT 229.800 615.600 231.600 623.100 ;
        RECT 237.000 622.800 240.600 623.700 ;
        RECT 248.400 623.700 252.150 624.750 ;
        RECT 237.000 615.600 238.800 622.800 ;
        RECT 248.400 621.600 249.600 623.700 ;
        RECT 247.800 615.600 249.600 621.600 ;
        RECT 250.800 620.700 258.600 622.050 ;
        RECT 265.950 621.600 267.000 628.050 ;
        RECT 268.950 626.850 271.050 628.950 ;
        RECT 271.950 628.050 274.050 630.150 ;
        RECT 277.950 629.850 280.050 631.950 ;
        RECT 280.950 631.050 283.050 633.150 ;
        RECT 278.100 628.050 279.900 629.850 ;
        RECT 268.950 625.050 270.750 626.850 ;
        RECT 281.400 623.700 282.600 631.050 ;
        RECT 283.950 629.850 286.050 631.950 ;
        RECT 286.950 630.450 289.050 631.050 ;
        RECT 284.100 628.050 285.900 629.850 ;
        RECT 286.950 629.550 291.450 630.450 ;
        RECT 293.400 630.150 294.600 635.400 ;
        RECT 302.250 633.150 304.050 634.950 ;
        RECT 301.950 631.050 304.050 633.150 ;
        RECT 305.850 630.150 307.050 635.400 ;
        RECT 311.100 630.150 312.900 631.950 ;
        RECT 286.950 628.950 289.050 629.550 ;
        RECT 290.550 625.050 291.450 629.550 ;
        RECT 292.950 628.050 295.050 630.150 ;
        RECT 281.400 622.800 285.000 623.700 ;
        RECT 289.950 622.950 292.050 625.050 ;
        RECT 250.800 615.600 252.600 620.700 ;
        RECT 256.800 615.600 258.600 620.700 ;
        RECT 265.200 615.600 267.000 621.600 ;
        RECT 283.200 615.600 285.000 622.800 ;
        RECT 293.400 621.600 294.600 628.050 ;
        RECT 295.950 626.850 298.050 628.950 ;
        RECT 304.950 628.050 307.050 630.150 ;
        RECT 296.100 625.050 297.900 626.850 ;
        RECT 304.950 624.750 306.150 628.050 ;
        RECT 307.950 626.850 310.050 628.950 ;
        RECT 310.950 628.050 313.050 630.150 ;
        RECT 317.400 628.950 318.600 641.400 ;
        RECT 329.400 633.150 330.600 641.400 ;
        RECT 338.400 640.200 340.200 646.200 ;
        RECT 339.300 635.100 340.200 640.200 ;
        RECT 345.900 636.900 347.700 646.200 ;
        RECT 359.400 641.400 361.200 647.400 ;
        RECT 345.900 636.000 348.000 636.900 ;
        RECT 339.300 634.200 345.450 635.100 ;
        RECT 325.950 629.850 328.050 631.950 ;
        RECT 328.950 631.050 331.050 633.150 ;
        RECT 316.950 626.850 319.050 628.950 ;
        RECT 320.100 627.150 321.900 628.950 ;
        RECT 326.100 628.050 327.900 629.850 ;
        RECT 308.100 625.050 309.900 626.850 ;
        RECT 302.400 623.700 306.150 624.750 ;
        RECT 302.400 621.600 303.600 623.700 ;
        RECT 292.800 615.600 294.600 621.600 ;
        RECT 301.800 615.600 303.600 621.600 ;
        RECT 304.800 620.700 312.600 622.050 ;
        RECT 304.800 615.600 306.600 620.700 ;
        RECT 310.800 615.600 312.600 620.700 ;
        RECT 317.400 618.600 318.600 626.850 ;
        RECT 319.950 625.050 322.050 627.150 ;
        RECT 329.400 623.700 330.600 631.050 ;
        RECT 331.950 629.850 334.050 631.950 ;
        RECT 341.100 630.150 342.900 631.950 ;
        RECT 344.250 631.500 345.450 634.200 ;
        RECT 332.100 628.050 333.900 629.850 ;
        RECT 337.950 626.850 340.050 628.950 ;
        RECT 340.950 628.050 343.050 630.150 ;
        RECT 344.250 629.700 346.050 631.500 ;
        RECT 338.100 625.050 339.900 626.850 ;
        RECT 344.250 624.000 345.450 629.700 ;
        RECT 347.100 628.950 348.000 636.000 ;
        RECT 359.400 634.500 360.600 641.400 ;
        RECT 365.700 635.400 367.500 647.400 ;
        RECT 374.400 641.400 376.200 647.400 ;
        RECT 359.400 633.600 365.100 634.500 ;
        RECT 363.150 632.700 365.100 633.600 ;
        RECT 350.100 630.150 351.900 631.950 ;
        RECT 359.100 630.150 360.900 631.950 ;
        RECT 346.950 626.850 349.050 628.950 ;
        RECT 349.950 628.050 352.050 630.150 ;
        RECT 358.950 628.050 361.050 630.150 ;
        RECT 316.800 615.600 318.600 618.600 ;
        RECT 327.000 622.800 330.600 623.700 ;
        RECT 339.150 623.100 345.450 624.000 ;
        RECT 327.000 615.600 328.800 622.800 ;
        RECT 339.150 619.800 340.200 623.100 ;
        RECT 347.100 622.200 348.000 626.850 ;
        RECT 363.150 624.300 364.050 632.700 ;
        RECT 366.000 630.150 367.200 635.400 ;
        RECT 374.400 633.150 375.600 641.400 ;
        RECT 389.700 635.400 391.500 647.400 ;
        RECT 403.500 635.400 405.300 647.400 ;
        RECT 409.800 641.400 411.600 647.400 ;
        RECT 386.250 633.150 388.050 634.950 ;
        RECT 364.950 628.050 367.200 630.150 ;
        RECT 370.950 629.850 373.050 631.950 ;
        RECT 373.950 631.050 376.050 633.150 ;
        RECT 371.100 628.050 372.900 629.850 ;
        RECT 363.150 623.400 365.100 624.300 ;
        RECT 338.400 616.800 340.200 619.800 ;
        RECT 345.900 621.300 348.000 622.200 ;
        RECT 360.000 622.500 365.100 623.400 ;
        RECT 345.900 616.800 347.700 621.300 ;
        RECT 360.000 618.600 361.200 622.500 ;
        RECT 366.000 621.600 367.200 628.050 ;
        RECT 374.400 623.700 375.600 631.050 ;
        RECT 376.950 629.850 379.050 631.950 ;
        RECT 385.950 631.050 388.050 633.150 ;
        RECT 389.850 630.150 391.050 635.400 ;
        RECT 395.100 630.150 396.900 631.950 ;
        RECT 403.800 630.150 405.000 635.400 ;
        RECT 410.400 634.500 411.600 641.400 ;
        RECT 405.900 633.600 411.600 634.500 ;
        RECT 413.550 635.400 415.350 647.400 ;
        RECT 421.050 641.400 422.850 647.400 ;
        RECT 418.950 639.300 422.850 641.400 ;
        RECT 428.850 640.500 430.650 647.400 ;
        RECT 436.650 641.400 438.450 647.400 ;
        RECT 437.250 640.500 438.450 641.400 ;
        RECT 427.950 639.450 434.550 640.500 ;
        RECT 427.950 638.700 429.750 639.450 ;
        RECT 432.750 638.700 434.550 639.450 ;
        RECT 437.250 638.400 442.050 640.500 ;
        RECT 420.150 636.600 422.850 638.400 ;
        RECT 423.750 637.800 425.550 638.400 ;
        RECT 423.750 636.900 430.050 637.800 ;
        RECT 437.250 637.500 438.450 638.400 ;
        RECT 423.750 636.600 425.550 636.900 ;
        RECT 421.950 635.700 422.850 636.600 ;
        RECT 405.900 632.700 407.850 633.600 ;
        RECT 377.100 628.050 378.900 629.850 ;
        RECT 388.950 628.050 391.050 630.150 ;
        RECT 388.950 624.750 390.150 628.050 ;
        RECT 391.950 626.850 394.050 628.950 ;
        RECT 394.950 628.050 397.050 630.150 ;
        RECT 403.800 628.050 406.050 630.150 ;
        RECT 392.100 625.050 393.900 626.850 ;
        RECT 386.400 623.700 390.150 624.750 ;
        RECT 374.400 622.800 378.000 623.700 ;
        RECT 359.400 615.600 361.200 618.600 ;
        RECT 365.700 615.600 367.500 621.600 ;
        RECT 376.200 615.600 378.000 622.800 ;
        RECT 386.400 621.600 387.600 623.700 ;
        RECT 385.800 615.600 387.600 621.600 ;
        RECT 388.800 620.700 396.600 622.050 ;
        RECT 403.800 621.600 405.000 628.050 ;
        RECT 406.950 624.300 407.850 632.700 ;
        RECT 410.100 630.150 411.900 631.950 ;
        RECT 409.950 628.050 412.050 630.150 ;
        RECT 405.900 623.400 407.850 624.300 ;
        RECT 413.550 625.950 414.750 635.400 ;
        RECT 418.950 634.800 421.050 635.700 ;
        RECT 421.950 634.800 427.950 635.700 ;
        RECT 416.850 633.600 421.050 634.800 ;
        RECT 415.950 631.800 417.750 633.600 ;
        RECT 427.050 630.150 427.950 634.800 ;
        RECT 429.150 634.800 430.050 636.900 ;
        RECT 430.950 636.300 438.450 637.500 ;
        RECT 430.950 635.700 432.750 636.300 ;
        RECT 445.050 635.400 446.850 647.400 ;
        RECT 458.700 635.400 460.500 647.400 ;
        RECT 470.400 641.400 472.200 647.400 ;
        RECT 435.750 634.800 446.850 635.400 ;
        RECT 429.150 634.200 446.850 634.800 ;
        RECT 429.150 633.900 437.550 634.200 ;
        RECT 435.750 633.600 437.550 633.900 ;
        RECT 427.050 628.050 430.050 630.150 ;
        RECT 433.950 629.100 436.050 630.150 ;
        RECT 433.950 628.050 441.900 629.100 ;
        RECT 415.950 627.750 418.050 628.050 ;
        RECT 415.950 625.950 419.850 627.750 ;
        RECT 413.550 623.850 418.050 625.950 ;
        RECT 427.050 624.000 427.950 628.050 ;
        RECT 440.100 627.300 441.900 628.050 ;
        RECT 443.100 627.150 444.900 628.950 ;
        RECT 437.100 626.400 438.900 627.000 ;
        RECT 443.100 626.400 444.000 627.150 ;
        RECT 437.100 625.200 444.000 626.400 ;
        RECT 437.100 624.000 438.150 625.200 ;
        RECT 405.900 622.500 411.000 623.400 ;
        RECT 388.800 615.600 390.600 620.700 ;
        RECT 394.800 615.600 396.600 620.700 ;
        RECT 403.500 615.600 405.300 621.600 ;
        RECT 409.800 618.600 411.000 622.500 ;
        RECT 413.550 621.600 414.750 623.850 ;
        RECT 427.050 623.100 438.150 624.000 ;
        RECT 427.050 622.800 427.950 623.100 ;
        RECT 409.800 615.600 411.600 618.600 ;
        RECT 413.550 615.600 415.350 621.600 ;
        RECT 418.950 620.700 421.050 621.600 ;
        RECT 426.150 621.000 427.950 622.800 ;
        RECT 437.100 622.200 438.150 623.100 ;
        RECT 433.350 621.450 435.150 622.200 ;
        RECT 418.950 619.500 422.700 620.700 ;
        RECT 421.650 618.600 422.700 619.500 ;
        RECT 430.200 620.400 435.150 621.450 ;
        RECT 436.650 620.400 438.450 622.200 ;
        RECT 445.950 621.600 446.850 634.200 ;
        RECT 455.250 633.150 457.050 634.950 ;
        RECT 454.950 631.050 457.050 633.150 ;
        RECT 458.850 630.150 460.050 635.400 ;
        RECT 470.400 633.150 471.600 641.400 ;
        RECT 479.550 635.400 481.350 647.400 ;
        RECT 487.050 641.400 488.850 647.400 ;
        RECT 484.950 639.300 488.850 641.400 ;
        RECT 494.850 640.500 496.650 647.400 ;
        RECT 502.650 641.400 504.450 647.400 ;
        RECT 503.250 640.500 504.450 641.400 ;
        RECT 493.950 639.450 500.550 640.500 ;
        RECT 493.950 638.700 495.750 639.450 ;
        RECT 498.750 638.700 500.550 639.450 ;
        RECT 503.250 638.400 508.050 640.500 ;
        RECT 486.150 636.600 488.850 638.400 ;
        RECT 489.750 637.800 491.550 638.400 ;
        RECT 489.750 636.900 496.050 637.800 ;
        RECT 503.250 637.500 504.450 638.400 ;
        RECT 489.750 636.600 491.550 636.900 ;
        RECT 487.950 635.700 488.850 636.600 ;
        RECT 464.100 630.150 465.900 631.950 ;
        RECT 457.950 628.050 460.050 630.150 ;
        RECT 457.950 624.750 459.150 628.050 ;
        RECT 460.950 626.850 463.050 628.950 ;
        RECT 463.950 628.050 466.050 630.150 ;
        RECT 466.950 629.850 469.050 631.950 ;
        RECT 469.950 631.050 472.050 633.150 ;
        RECT 467.100 628.050 468.900 629.850 ;
        RECT 461.100 625.050 462.900 626.850 ;
        RECT 455.400 623.700 459.150 624.750 ;
        RECT 470.400 623.700 471.600 631.050 ;
        RECT 472.950 629.850 475.050 631.950 ;
        RECT 473.100 628.050 474.900 629.850 ;
        RECT 479.550 625.950 480.750 635.400 ;
        RECT 484.950 634.800 487.050 635.700 ;
        RECT 487.950 634.800 493.950 635.700 ;
        RECT 482.850 633.600 487.050 634.800 ;
        RECT 481.950 631.800 483.750 633.600 ;
        RECT 493.050 630.150 493.950 634.800 ;
        RECT 495.150 634.800 496.050 636.900 ;
        RECT 496.950 636.300 504.450 637.500 ;
        RECT 496.950 635.700 498.750 636.300 ;
        RECT 511.050 635.400 512.850 647.400 ;
        RECT 501.750 634.800 512.850 635.400 ;
        RECT 495.150 634.200 512.850 634.800 ;
        RECT 495.150 633.900 503.550 634.200 ;
        RECT 501.750 633.600 503.550 633.900 ;
        RECT 493.050 628.050 496.050 630.150 ;
        RECT 499.950 629.100 502.050 630.150 ;
        RECT 499.950 628.050 507.900 629.100 ;
        RECT 481.950 627.750 484.050 628.050 ;
        RECT 481.950 625.950 485.850 627.750 ;
        RECT 479.550 623.850 484.050 625.950 ;
        RECT 493.050 624.000 493.950 628.050 ;
        RECT 506.100 627.300 507.900 628.050 ;
        RECT 509.100 627.150 510.900 628.950 ;
        RECT 503.100 626.400 504.900 627.000 ;
        RECT 509.100 626.400 510.000 627.150 ;
        RECT 503.100 625.200 510.000 626.400 ;
        RECT 503.100 624.000 504.150 625.200 ;
        RECT 455.400 621.600 456.600 623.700 ;
        RECT 470.400 622.800 474.000 623.700 ;
        RECT 430.200 618.600 431.250 620.400 ;
        RECT 439.950 619.500 442.050 621.600 ;
        RECT 439.950 618.600 441.000 619.500 ;
        RECT 421.650 615.600 423.450 618.600 ;
        RECT 429.450 615.600 431.250 618.600 ;
        RECT 437.250 617.700 441.000 618.600 ;
        RECT 437.250 615.600 439.050 617.700 ;
        RECT 445.050 615.600 446.850 621.600 ;
        RECT 454.800 615.600 456.600 621.600 ;
        RECT 457.800 620.700 465.600 622.050 ;
        RECT 457.800 615.600 459.600 620.700 ;
        RECT 463.800 615.600 465.600 620.700 ;
        RECT 472.200 615.600 474.000 622.800 ;
        RECT 479.550 621.600 480.750 623.850 ;
        RECT 493.050 623.100 504.150 624.000 ;
        RECT 493.050 622.800 493.950 623.100 ;
        RECT 479.550 615.600 481.350 621.600 ;
        RECT 484.950 620.700 487.050 621.600 ;
        RECT 492.150 621.000 493.950 622.800 ;
        RECT 503.100 622.200 504.150 623.100 ;
        RECT 499.350 621.450 501.150 622.200 ;
        RECT 484.950 619.500 488.700 620.700 ;
        RECT 487.650 618.600 488.700 619.500 ;
        RECT 496.200 620.400 501.150 621.450 ;
        RECT 502.650 620.400 504.450 622.200 ;
        RECT 511.950 621.600 512.850 634.200 ;
        RECT 515.400 641.400 517.200 647.400 ;
        RECT 515.400 634.500 516.600 641.400 ;
        RECT 521.700 635.400 523.500 647.400 ;
        RECT 535.800 641.400 537.600 647.400 ;
        RECT 515.400 633.600 521.100 634.500 ;
        RECT 519.150 632.700 521.100 633.600 ;
        RECT 515.100 630.150 516.900 631.950 ;
        RECT 514.950 628.050 517.050 630.150 ;
        RECT 519.150 624.300 520.050 632.700 ;
        RECT 522.000 630.150 523.200 635.400 ;
        RECT 536.400 633.150 537.600 641.400 ;
        RECT 548.700 635.400 550.500 647.400 ;
        RECT 562.800 641.400 564.600 647.400 ;
        RECT 545.250 633.150 547.050 634.950 ;
        RECT 520.950 628.050 523.200 630.150 ;
        RECT 532.950 629.850 535.050 631.950 ;
        RECT 535.950 631.050 538.050 633.150 ;
        RECT 533.100 628.050 534.900 629.850 ;
        RECT 519.150 623.400 521.100 624.300 ;
        RECT 496.200 618.600 497.250 620.400 ;
        RECT 505.950 619.500 508.050 621.600 ;
        RECT 505.950 618.600 507.000 619.500 ;
        RECT 487.650 615.600 489.450 618.600 ;
        RECT 495.450 615.600 497.250 618.600 ;
        RECT 503.250 617.700 507.000 618.600 ;
        RECT 503.250 615.600 505.050 617.700 ;
        RECT 511.050 615.600 512.850 621.600 ;
        RECT 516.000 622.500 521.100 623.400 ;
        RECT 516.000 618.600 517.200 622.500 ;
        RECT 522.000 621.600 523.200 628.050 ;
        RECT 536.400 623.700 537.600 631.050 ;
        RECT 538.950 629.850 541.050 631.950 ;
        RECT 544.950 631.050 547.050 633.150 ;
        RECT 548.850 630.150 550.050 635.400 ;
        RECT 563.400 633.150 564.600 641.400 ;
        RECT 575.700 635.400 577.500 647.400 ;
        RECT 584.400 641.400 586.200 647.400 ;
        RECT 572.250 633.150 574.050 634.950 ;
        RECT 554.100 630.150 555.900 631.950 ;
        RECT 539.100 628.050 540.900 629.850 ;
        RECT 547.950 628.050 550.050 630.150 ;
        RECT 547.950 624.750 549.150 628.050 ;
        RECT 550.950 626.850 553.050 628.950 ;
        RECT 553.950 628.050 556.050 630.150 ;
        RECT 559.950 629.850 562.050 631.950 ;
        RECT 562.950 631.050 565.050 633.150 ;
        RECT 560.100 628.050 561.900 629.850 ;
        RECT 551.100 625.050 552.900 626.850 ;
        RECT 534.000 622.800 537.600 623.700 ;
        RECT 545.400 623.700 549.150 624.750 ;
        RECT 563.400 623.700 564.600 631.050 ;
        RECT 565.950 629.850 568.050 631.950 ;
        RECT 571.950 631.050 574.050 633.150 ;
        RECT 575.850 630.150 577.050 635.400 ;
        RECT 584.400 634.500 585.600 641.400 ;
        RECT 590.700 635.400 592.500 647.400 ;
        RECT 601.500 635.400 603.300 647.400 ;
        RECT 612.150 635.400 613.950 647.400 ;
        RECT 620.550 641.400 622.350 647.400 ;
        RECT 620.550 640.500 621.750 641.400 ;
        RECT 628.350 640.500 630.150 647.400 ;
        RECT 636.150 641.400 637.950 647.400 ;
        RECT 616.950 638.400 621.750 640.500 ;
        RECT 624.450 639.450 631.050 640.500 ;
        RECT 624.450 638.700 626.250 639.450 ;
        RECT 629.250 638.700 631.050 639.450 ;
        RECT 636.150 639.300 640.050 641.400 ;
        RECT 620.550 637.500 621.750 638.400 ;
        RECT 633.450 637.800 635.250 638.400 ;
        RECT 620.550 636.300 628.050 637.500 ;
        RECT 626.250 635.700 628.050 636.300 ;
        RECT 628.950 636.900 635.250 637.800 ;
        RECT 584.400 633.600 590.100 634.500 ;
        RECT 588.150 632.700 590.100 633.600 ;
        RECT 581.100 630.150 582.900 631.950 ;
        RECT 584.100 630.150 585.900 631.950 ;
        RECT 566.100 628.050 567.900 629.850 ;
        RECT 574.950 628.050 577.050 630.150 ;
        RECT 574.950 624.750 576.150 628.050 ;
        RECT 577.950 626.850 580.050 628.950 ;
        RECT 580.950 628.050 583.050 630.150 ;
        RECT 583.950 628.050 586.050 630.150 ;
        RECT 578.100 625.050 579.900 626.850 ;
        RECT 515.400 615.600 517.200 618.600 ;
        RECT 521.700 615.600 523.500 621.600 ;
        RECT 534.000 615.600 535.800 622.800 ;
        RECT 545.400 621.600 546.600 623.700 ;
        RECT 561.000 622.800 564.600 623.700 ;
        RECT 572.400 623.700 576.150 624.750 ;
        RECT 588.150 624.300 589.050 632.700 ;
        RECT 591.000 630.150 592.200 635.400 ;
        RECT 596.100 630.150 597.900 631.950 ;
        RECT 601.950 630.150 603.150 635.400 ;
        RECT 604.950 633.150 606.750 634.950 ;
        RECT 612.150 634.800 623.250 635.400 ;
        RECT 628.950 634.800 629.850 636.900 ;
        RECT 633.450 636.600 635.250 636.900 ;
        RECT 636.150 636.600 638.850 638.400 ;
        RECT 636.150 635.700 637.050 636.600 ;
        RECT 612.150 634.200 629.850 634.800 ;
        RECT 604.950 631.050 607.050 633.150 ;
        RECT 589.950 628.050 592.200 630.150 ;
        RECT 595.950 628.050 598.050 630.150 ;
        RECT 544.800 615.600 546.600 621.600 ;
        RECT 547.800 620.700 555.600 622.050 ;
        RECT 547.800 615.600 549.600 620.700 ;
        RECT 553.800 615.600 555.600 620.700 ;
        RECT 561.000 615.600 562.800 622.800 ;
        RECT 572.400 621.600 573.600 623.700 ;
        RECT 588.150 623.400 590.100 624.300 ;
        RECT 585.000 622.500 590.100 623.400 ;
        RECT 571.800 615.600 573.600 621.600 ;
        RECT 574.800 620.700 582.600 622.050 ;
        RECT 574.800 615.600 576.600 620.700 ;
        RECT 580.800 615.600 582.600 620.700 ;
        RECT 585.000 618.600 586.200 622.500 ;
        RECT 591.000 621.600 592.200 628.050 ;
        RECT 598.950 626.850 601.050 628.950 ;
        RECT 601.950 628.050 604.050 630.150 ;
        RECT 599.100 625.050 600.900 626.850 ;
        RECT 602.850 624.750 604.050 628.050 ;
        RECT 602.850 623.700 606.600 624.750 ;
        RECT 584.400 615.600 586.200 618.600 ;
        RECT 590.700 615.600 592.500 621.600 ;
        RECT 596.400 620.700 604.200 622.050 ;
        RECT 596.400 615.600 598.200 620.700 ;
        RECT 602.400 615.600 604.200 620.700 ;
        RECT 605.400 621.600 606.600 623.700 ;
        RECT 612.150 621.600 613.050 634.200 ;
        RECT 621.450 633.900 629.850 634.200 ;
        RECT 631.050 634.800 637.050 635.700 ;
        RECT 637.950 634.800 640.050 635.700 ;
        RECT 643.650 635.400 645.450 647.400 ;
        RECT 651.300 636.900 653.100 647.400 ;
        RECT 621.450 633.600 623.250 633.900 ;
        RECT 631.050 630.150 631.950 634.800 ;
        RECT 637.950 633.600 642.150 634.800 ;
        RECT 641.250 631.800 643.050 633.600 ;
        RECT 622.950 629.100 625.050 630.150 ;
        RECT 614.100 627.150 615.900 628.950 ;
        RECT 617.100 628.050 625.050 629.100 ;
        RECT 628.950 628.050 631.950 630.150 ;
        RECT 617.100 627.300 618.900 628.050 ;
        RECT 615.000 626.400 615.900 627.150 ;
        RECT 620.100 626.400 621.900 627.000 ;
        RECT 615.000 625.200 621.900 626.400 ;
        RECT 620.850 624.000 621.900 625.200 ;
        RECT 631.050 624.000 631.950 628.050 ;
        RECT 640.950 627.750 643.050 628.050 ;
        RECT 639.150 625.950 643.050 627.750 ;
        RECT 644.250 625.950 645.450 635.400 ;
        RECT 650.700 635.550 653.100 636.900 ;
        RECT 650.700 628.950 652.050 635.550 ;
        RECT 658.800 635.400 660.600 647.400 ;
        RECT 668.700 635.400 670.500 647.400 ;
        RECT 683.700 635.400 685.500 647.400 ;
        RECT 700.800 635.400 704.100 647.400 ;
        RECT 713.400 641.400 715.200 647.400 ;
        RECT 721.800 646.500 729.600 647.400 ;
        RECT 620.850 623.100 631.950 624.000 ;
        RECT 640.950 623.850 645.450 625.950 ;
        RECT 620.850 622.200 621.900 623.100 ;
        RECT 631.050 622.800 631.950 623.100 ;
        RECT 605.400 615.600 607.200 621.600 ;
        RECT 612.150 615.600 613.950 621.600 ;
        RECT 616.950 619.500 619.050 621.600 ;
        RECT 620.550 620.400 622.350 622.200 ;
        RECT 623.850 621.450 625.650 622.200 ;
        RECT 623.850 620.400 628.800 621.450 ;
        RECT 631.050 621.000 632.850 622.800 ;
        RECT 644.250 621.600 645.450 623.850 ;
        RECT 649.950 626.850 652.050 628.950 ;
        RECT 653.400 634.200 655.200 634.650 ;
        RECT 659.400 634.200 660.600 635.400 ;
        RECT 653.400 633.000 660.600 634.200 ;
        RECT 665.250 633.150 667.050 634.950 ;
        RECT 653.400 632.850 655.200 633.000 ;
        RECT 649.950 621.600 651.000 626.850 ;
        RECT 653.400 624.600 654.300 632.850 ;
        RECT 656.100 630.150 657.900 631.950 ;
        RECT 664.950 631.050 667.050 633.150 ;
        RECT 668.850 630.150 670.050 635.400 ;
        RECT 676.950 631.950 679.050 634.050 ;
        RECT 680.250 633.150 682.050 634.950 ;
        RECT 674.100 630.150 675.900 631.950 ;
        RECT 655.950 628.050 658.050 630.150 ;
        RECT 659.100 627.150 660.900 628.950 ;
        RECT 667.950 628.050 670.050 630.150 ;
        RECT 658.950 625.050 661.050 627.150 ;
        RECT 667.950 624.750 669.150 628.050 ;
        RECT 670.950 626.850 673.050 628.950 ;
        RECT 673.950 628.050 676.050 630.150 ;
        RECT 677.550 627.450 678.450 631.950 ;
        RECT 679.950 631.050 682.050 633.150 ;
        RECT 683.850 630.150 685.050 635.400 ;
        RECT 689.100 630.150 690.900 631.950 ;
        RECT 695.250 630.150 697.050 631.950 ;
        RECT 701.400 630.150 702.600 635.400 ;
        RECT 707.100 630.150 708.900 631.950 ;
        RECT 682.950 628.050 685.050 630.150 ;
        RECT 679.950 627.450 682.050 628.050 ;
        RECT 671.100 625.050 672.900 626.850 ;
        RECT 677.550 626.550 682.050 627.450 ;
        RECT 679.950 625.950 682.050 626.550 ;
        RECT 682.950 624.750 684.150 628.050 ;
        RECT 685.950 626.850 688.050 628.950 ;
        RECT 688.950 628.050 691.050 630.150 ;
        RECT 694.950 628.050 697.050 630.150 ;
        RECT 697.950 626.850 700.050 628.950 ;
        RECT 700.950 628.050 703.050 630.150 ;
        RECT 686.100 625.050 687.900 626.850 ;
        RECT 698.700 625.050 700.500 626.850 ;
        RECT 653.250 623.700 655.050 624.600 ;
        RECT 665.400 623.700 669.150 624.750 ;
        RECT 680.400 623.700 684.150 624.750 ;
        RECT 701.400 624.150 702.600 628.050 ;
        RECT 703.950 626.850 706.050 628.950 ;
        RECT 706.950 628.050 709.050 630.150 ;
        RECT 713.400 628.950 714.600 641.400 ;
        RECT 721.800 635.400 723.600 646.500 ;
        RECT 724.800 634.500 726.600 645.600 ;
        RECT 727.800 636.600 729.600 646.500 ;
        RECT 733.800 636.600 735.600 647.400 ;
        RECT 727.800 635.700 735.600 636.600 ;
        RECT 743.400 641.400 745.200 647.400 ;
        RECT 724.800 633.600 728.850 634.500 ;
        RECT 722.100 630.150 723.900 631.950 ;
        RECT 727.950 630.150 728.850 633.600 ;
        RECT 733.950 630.150 735.750 631.950 ;
        RECT 710.100 627.150 711.900 628.950 ;
        RECT 704.100 625.050 705.900 626.850 ;
        RECT 709.950 625.050 712.050 627.150 ;
        RECT 712.950 626.850 715.050 628.950 ;
        RECT 721.950 628.050 724.050 630.150 ;
        RECT 724.950 626.850 727.050 628.950 ;
        RECT 727.950 628.050 730.050 630.150 ;
        RECT 653.250 622.800 656.700 623.700 ;
        RECT 637.950 620.700 640.050 621.600 ;
        RECT 618.000 618.600 619.050 619.500 ;
        RECT 627.750 618.600 628.800 620.400 ;
        RECT 636.300 619.500 640.050 620.700 ;
        RECT 636.300 618.600 637.350 619.500 ;
        RECT 618.000 617.700 621.750 618.600 ;
        RECT 619.950 615.600 621.750 617.700 ;
        RECT 627.750 615.600 629.550 618.600 ;
        RECT 635.550 615.600 637.350 618.600 ;
        RECT 643.650 615.600 645.450 621.600 ;
        RECT 649.800 615.600 651.600 621.600 ;
        RECT 655.800 618.600 656.700 622.800 ;
        RECT 665.400 621.600 666.600 623.700 ;
        RECT 655.800 615.600 657.600 618.600 ;
        RECT 664.800 615.600 666.600 621.600 ;
        RECT 667.800 620.700 675.600 622.050 ;
        RECT 680.400 621.600 681.600 623.700 ;
        RECT 698.400 623.100 702.600 624.150 ;
        RECT 667.800 615.600 669.600 620.700 ;
        RECT 673.800 615.600 675.600 620.700 ;
        RECT 679.800 615.600 681.600 621.600 ;
        RECT 682.800 620.700 690.600 622.050 ;
        RECT 698.400 621.600 699.300 623.100 ;
        RECT 682.800 615.600 684.600 620.700 ;
        RECT 688.800 615.600 690.600 620.700 ;
        RECT 694.800 616.500 696.600 621.600 ;
        RECT 697.800 617.400 699.600 621.600 ;
        RECT 700.800 621.000 708.600 621.900 ;
        RECT 700.800 616.500 702.600 621.000 ;
        RECT 694.800 615.600 702.600 616.500 ;
        RECT 706.800 615.600 708.600 621.000 ;
        RECT 713.400 618.600 714.600 626.850 ;
        RECT 725.250 625.050 727.050 626.850 ;
        RECT 729.000 621.600 730.050 628.050 ;
        RECT 730.950 626.850 733.050 628.950 ;
        RECT 733.950 628.050 736.050 630.150 ;
        RECT 743.400 628.950 744.600 641.400 ;
        RECT 755.700 635.400 757.500 647.400 ;
        RECT 752.250 633.150 754.050 634.950 ;
        RECT 751.950 631.050 754.050 633.150 ;
        RECT 755.850 630.150 757.050 635.400 ;
        RECT 761.100 630.150 762.900 631.950 ;
        RECT 740.100 627.150 741.900 628.950 ;
        RECT 730.950 625.050 732.750 626.850 ;
        RECT 739.950 625.050 742.050 627.150 ;
        RECT 742.950 626.850 745.050 628.950 ;
        RECT 754.950 628.050 757.050 630.150 ;
        RECT 713.400 615.600 715.200 618.600 ;
        RECT 729.000 615.600 730.800 621.600 ;
        RECT 743.400 618.600 744.600 626.850 ;
        RECT 754.950 624.750 756.150 628.050 ;
        RECT 757.950 626.850 760.050 628.950 ;
        RECT 760.950 628.050 763.050 630.150 ;
        RECT 758.100 625.050 759.900 626.850 ;
        RECT 752.400 623.700 756.150 624.750 ;
        RECT 752.400 621.600 753.600 623.700 ;
        RECT 743.400 615.600 745.200 618.600 ;
        RECT 751.800 615.600 753.600 621.600 ;
        RECT 754.800 620.700 762.600 622.050 ;
        RECT 754.800 615.600 756.600 620.700 ;
        RECT 760.800 615.600 762.600 620.700 ;
        RECT 5.400 606.300 7.200 611.400 ;
        RECT 11.400 606.300 13.200 611.400 ;
        RECT 5.400 604.950 13.200 606.300 ;
        RECT 14.400 605.400 16.200 611.400 ;
        RECT 25.800 608.400 27.600 611.400 ;
        RECT 14.400 603.300 15.600 605.400 ;
        RECT 11.850 602.250 15.600 603.300 ;
        RECT 8.100 600.150 9.900 601.950 ;
        RECT 4.950 596.850 7.050 598.950 ;
        RECT 7.950 598.050 10.050 600.150 ;
        RECT 11.850 598.950 13.050 602.250 ;
        RECT 26.400 600.150 27.600 608.400 ;
        RECT 32.400 606.300 34.200 611.400 ;
        RECT 38.400 606.300 40.200 611.400 ;
        RECT 32.400 604.950 40.200 606.300 ;
        RECT 41.400 605.400 43.200 611.400 ;
        RECT 41.400 603.300 42.600 605.400 ;
        RECT 54.000 604.200 55.800 611.400 ;
        RECT 54.000 603.300 57.600 604.200 ;
        RECT 38.850 602.250 42.600 603.300 ;
        RECT 10.950 596.850 13.050 598.950 ;
        RECT 25.950 598.050 28.050 600.150 ;
        RECT 28.950 599.850 31.050 601.950 ;
        RECT 35.100 600.150 36.900 601.950 ;
        RECT 29.100 598.050 30.900 599.850 ;
        RECT 5.100 595.050 6.900 596.850 ;
        RECT 10.950 591.600 12.150 596.850 ;
        RECT 13.950 593.850 16.050 595.950 ;
        RECT 13.950 592.050 15.750 593.850 ;
        RECT 10.500 579.600 12.300 591.600 ;
        RECT 26.400 585.600 27.600 598.050 ;
        RECT 31.950 596.850 34.050 598.950 ;
        RECT 34.950 598.050 37.050 600.150 ;
        RECT 38.850 598.950 40.050 602.250 ;
        RECT 37.950 596.850 40.050 598.950 ;
        RECT 53.100 597.150 54.900 598.950 ;
        RECT 32.100 595.050 33.900 596.850 ;
        RECT 37.950 591.600 39.150 596.850 ;
        RECT 40.950 593.850 43.050 595.950 ;
        RECT 52.950 595.050 55.050 597.150 ;
        RECT 56.400 595.950 57.600 603.300 ;
        RECT 71.100 603.000 72.900 611.400 ;
        RECT 87.000 607.050 88.800 611.400 ;
        RECT 97.800 608.400 99.600 611.400 ;
        RECT 83.400 605.400 88.800 607.050 ;
        RECT 71.100 601.350 75.300 603.000 ;
        RECT 59.100 597.150 60.900 598.950 ;
        RECT 74.400 597.150 75.300 601.350 ;
        RECT 83.400 598.950 84.300 605.400 ;
        RECT 86.100 600.150 87.900 601.950 ;
        RECT 55.950 593.850 58.050 595.950 ;
        RECT 58.950 595.050 61.050 597.150 ;
        RECT 64.950 593.850 67.050 595.950 ;
        RECT 70.950 593.850 73.050 595.950 ;
        RECT 73.950 595.050 76.050 597.150 ;
        RECT 82.950 596.850 85.050 598.950 ;
        RECT 85.950 598.050 88.050 600.150 ;
        RECT 88.950 599.850 91.050 601.950 ;
        RECT 92.100 600.150 93.900 601.950 ;
        RECT 98.400 600.150 99.600 608.400 ;
        RECT 109.200 604.200 111.000 611.400 ;
        RECT 107.400 603.300 111.000 604.200 ;
        RECT 119.400 608.400 121.200 611.400 ;
        RECT 89.100 598.050 90.900 599.850 ;
        RECT 91.950 598.050 94.050 600.150 ;
        RECT 97.950 598.050 100.050 600.150 ;
        RECT 100.950 599.850 103.050 601.950 ;
        RECT 101.100 598.050 102.900 599.850 ;
        RECT 40.950 592.050 42.750 593.850 ;
        RECT 25.800 579.600 27.600 585.600 ;
        RECT 37.500 579.600 39.300 591.600 ;
        RECT 56.400 585.600 57.600 593.850 ;
        RECT 65.100 592.050 66.900 593.850 ;
        RECT 67.950 590.850 70.050 592.950 ;
        RECT 71.250 592.050 73.050 593.850 ;
        RECT 68.100 589.050 69.900 590.850 ;
        RECT 74.400 586.800 75.300 595.050 ;
        RECT 83.400 591.600 84.300 596.850 ;
        RECT 68.700 585.900 75.300 586.800 ;
        RECT 68.700 585.600 70.200 585.900 ;
        RECT 55.800 579.600 57.600 585.600 ;
        RECT 68.400 579.600 70.200 585.600 ;
        RECT 74.400 585.600 75.300 585.900 ;
        RECT 74.400 579.600 76.200 585.600 ;
        RECT 82.800 579.600 84.600 591.600 ;
        RECT 85.800 590.700 93.600 591.600 ;
        RECT 85.800 579.600 87.600 590.700 ;
        RECT 91.800 579.600 93.600 590.700 ;
        RECT 98.400 585.600 99.600 598.050 ;
        RECT 104.100 597.150 105.900 598.950 ;
        RECT 103.950 595.050 106.050 597.150 ;
        RECT 107.400 595.950 108.600 603.300 ;
        RECT 115.950 599.850 118.050 601.950 ;
        RECT 119.400 600.150 120.600 608.400 ;
        RECT 127.500 605.400 129.300 611.400 ;
        RECT 133.800 608.400 135.600 611.400 ;
        RECT 140.400 608.400 142.200 611.400 ;
        RECT 110.100 597.150 111.900 598.950 ;
        RECT 116.100 598.050 117.900 599.850 ;
        RECT 118.950 598.050 121.050 600.150 ;
        RECT 127.800 598.950 129.000 605.400 ;
        RECT 133.800 604.500 135.000 608.400 ;
        RECT 129.900 603.600 135.000 604.500 ;
        RECT 141.000 604.500 142.200 608.400 ;
        RECT 146.700 605.400 148.500 611.400 ;
        RECT 141.000 603.600 146.100 604.500 ;
        RECT 129.900 602.700 131.850 603.600 ;
        RECT 106.950 593.850 109.050 595.950 ;
        RECT 109.950 595.050 112.050 597.150 ;
        RECT 97.800 579.600 99.600 585.600 ;
        RECT 107.400 585.600 108.600 593.850 ;
        RECT 119.400 585.600 120.600 598.050 ;
        RECT 127.800 596.850 130.050 598.950 ;
        RECT 127.800 591.600 129.000 596.850 ;
        RECT 130.950 594.300 131.850 602.700 ;
        RECT 144.150 602.700 146.100 603.600 ;
        RECT 133.950 596.850 136.050 598.950 ;
        RECT 139.950 596.850 142.050 598.950 ;
        RECT 134.100 595.050 135.900 596.850 ;
        RECT 140.100 595.050 141.900 596.850 ;
        RECT 129.900 593.400 131.850 594.300 ;
        RECT 144.150 594.300 145.050 602.700 ;
        RECT 147.000 598.950 148.200 605.400 ;
        RECT 156.000 604.200 157.800 611.400 ;
        RECT 169.800 608.400 171.600 611.400 ;
        RECT 178.800 608.400 180.600 611.400 ;
        RECT 156.000 603.300 159.600 604.200 ;
        RECT 145.950 596.850 148.200 598.950 ;
        RECT 155.100 597.150 156.900 598.950 ;
        RECT 144.150 593.400 146.100 594.300 ;
        RECT 129.900 592.500 135.600 593.400 ;
        RECT 107.400 579.600 109.200 585.600 ;
        RECT 119.400 579.600 121.200 585.600 ;
        RECT 127.500 579.600 129.300 591.600 ;
        RECT 134.400 585.600 135.600 592.500 ;
        RECT 133.800 579.600 135.600 585.600 ;
        RECT 140.400 592.500 146.100 593.400 ;
        RECT 140.400 585.600 141.600 592.500 ;
        RECT 147.000 591.600 148.200 596.850 ;
        RECT 154.950 595.050 157.050 597.150 ;
        RECT 158.400 595.950 159.600 603.300 ;
        RECT 169.950 601.950 171.000 608.400 ;
        RECT 169.950 599.850 172.050 601.950 ;
        RECT 179.400 600.150 180.600 608.400 ;
        RECT 190.200 604.200 192.000 611.400 ;
        RECT 199.800 605.400 201.600 611.400 ;
        RECT 188.400 603.300 192.000 604.200 ;
        RECT 200.400 603.300 201.600 605.400 ;
        RECT 202.800 606.300 204.600 611.400 ;
        RECT 208.800 606.300 210.600 611.400 ;
        RECT 202.800 604.950 210.600 606.300 ;
        RECT 217.200 605.400 219.000 611.400 ;
        RECT 161.100 597.150 162.900 598.950 ;
        RECT 157.950 593.850 160.050 595.950 ;
        RECT 160.950 595.050 163.050 597.150 ;
        RECT 166.950 596.850 169.050 598.950 ;
        RECT 167.100 595.050 168.900 596.850 ;
        RECT 140.400 579.600 142.200 585.600 ;
        RECT 146.700 579.600 148.500 591.600 ;
        RECT 158.400 585.600 159.600 593.850 ;
        RECT 169.950 592.650 171.000 599.850 ;
        RECT 172.950 596.850 175.050 598.950 ;
        RECT 178.950 598.050 181.050 600.150 ;
        RECT 181.950 599.850 184.050 601.950 ;
        RECT 182.100 598.050 183.900 599.850 ;
        RECT 173.100 595.050 174.900 596.850 ;
        RECT 157.800 579.600 159.600 585.600 ;
        RECT 168.600 591.600 171.000 592.650 ;
        RECT 168.600 579.600 170.400 591.600 ;
        RECT 179.400 585.600 180.600 598.050 ;
        RECT 185.100 597.150 186.900 598.950 ;
        RECT 184.950 595.050 187.050 597.150 ;
        RECT 188.400 595.950 189.600 603.300 ;
        RECT 200.400 602.250 204.150 603.300 ;
        RECT 202.950 598.950 204.150 602.250 ;
        RECT 206.100 600.150 207.900 601.950 ;
        RECT 215.250 600.150 217.050 601.950 ;
        RECT 191.100 597.150 192.900 598.950 ;
        RECT 187.950 593.850 190.050 595.950 ;
        RECT 190.950 595.050 193.050 597.150 ;
        RECT 202.950 596.850 205.050 598.950 ;
        RECT 205.950 598.050 208.050 600.150 ;
        RECT 208.950 596.850 211.050 598.950 ;
        RECT 211.950 596.850 214.050 598.950 ;
        RECT 214.950 598.050 217.050 600.150 ;
        RECT 217.950 598.950 219.000 605.400 ;
        RECT 235.200 604.200 237.000 611.400 ;
        RECT 245.400 606.300 247.200 611.400 ;
        RECT 251.400 606.300 253.200 611.400 ;
        RECT 245.400 604.950 253.200 606.300 ;
        RECT 254.400 605.400 256.200 611.400 ;
        RECT 267.300 606.900 269.100 611.400 ;
        RECT 265.950 605.400 269.100 606.900 ;
        RECT 233.400 603.300 237.000 604.200 ;
        RECT 254.400 603.300 255.600 605.400 ;
        RECT 220.950 600.150 222.750 601.950 ;
        RECT 217.950 596.850 220.050 598.950 ;
        RECT 220.950 598.050 223.050 600.150 ;
        RECT 223.950 596.850 226.050 598.950 ;
        RECT 230.100 597.150 231.900 598.950 ;
        RECT 199.950 593.850 202.050 595.950 ;
        RECT 178.800 579.600 180.600 585.600 ;
        RECT 188.400 585.600 189.600 593.850 ;
        RECT 200.250 592.050 202.050 593.850 ;
        RECT 203.850 591.600 205.050 596.850 ;
        RECT 209.100 595.050 210.900 596.850 ;
        RECT 212.250 595.050 214.050 596.850 ;
        RECT 219.150 593.400 220.050 596.850 ;
        RECT 224.100 595.050 225.900 596.850 ;
        RECT 229.950 595.050 232.050 597.150 ;
        RECT 233.400 595.950 234.600 603.300 ;
        RECT 251.850 602.250 255.600 603.300 ;
        RECT 248.100 600.150 249.900 601.950 ;
        RECT 236.100 597.150 237.900 598.950 ;
        RECT 232.950 593.850 235.050 595.950 ;
        RECT 235.950 595.050 238.050 597.150 ;
        RECT 244.950 596.850 247.050 598.950 ;
        RECT 247.950 598.050 250.050 600.150 ;
        RECT 251.850 598.950 253.050 602.250 ;
        RECT 250.950 596.850 253.050 598.950 ;
        RECT 265.950 598.950 267.000 605.400 ;
        RECT 269.100 603.900 270.900 604.500 ;
        RECT 274.800 603.900 276.600 611.400 ;
        RECT 269.100 602.700 276.600 603.900 ;
        RECT 284.100 603.000 285.900 611.400 ;
        RECT 295.800 605.400 297.600 611.400 ;
        RECT 265.950 596.850 268.050 598.950 ;
        RECT 269.100 597.150 270.900 598.950 ;
        RECT 245.100 595.050 246.900 596.850 ;
        RECT 219.150 592.500 223.200 593.400 ;
        RECT 188.400 579.600 190.200 585.600 ;
        RECT 203.700 579.600 205.500 591.600 ;
        RECT 212.400 590.400 220.200 591.300 ;
        RECT 212.400 579.600 214.200 590.400 ;
        RECT 218.400 580.500 220.200 590.400 ;
        RECT 221.400 581.400 223.200 592.500 ;
        RECT 224.400 580.500 226.200 591.600 ;
        RECT 218.400 579.600 226.200 580.500 ;
        RECT 233.400 585.600 234.600 593.850 ;
        RECT 250.950 591.600 252.150 596.850 ;
        RECT 253.950 593.850 256.050 595.950 ;
        RECT 253.950 592.050 255.750 593.850 ;
        RECT 265.950 591.600 267.000 596.850 ;
        RECT 268.950 595.050 271.050 597.150 ;
        RECT 233.400 579.600 235.200 585.600 ;
        RECT 250.500 579.600 252.300 591.600 ;
        RECT 265.200 579.600 267.000 591.600 ;
        RECT 272.400 585.600 273.450 602.700 ;
        RECT 281.700 601.350 285.900 603.000 ;
        RECT 296.400 603.300 297.600 605.400 ;
        RECT 298.800 606.300 300.600 611.400 ;
        RECT 304.800 606.300 306.600 611.400 ;
        RECT 311.400 608.400 313.200 611.400 ;
        RECT 325.800 608.400 327.600 611.400 ;
        RECT 298.800 604.950 306.600 606.300 ;
        RECT 296.400 602.250 300.150 603.300 ;
        RECT 274.950 596.850 277.050 598.950 ;
        RECT 281.700 597.150 282.600 601.350 ;
        RECT 298.950 598.950 300.150 602.250 ;
        RECT 312.000 601.950 313.050 608.400 ;
        RECT 302.100 600.150 303.900 601.950 ;
        RECT 275.100 595.050 276.900 596.850 ;
        RECT 280.950 595.050 283.050 597.150 ;
        RECT 298.950 596.850 301.050 598.950 ;
        RECT 301.950 598.050 304.050 600.150 ;
        RECT 310.950 599.850 313.050 601.950 ;
        RECT 326.400 600.150 327.600 608.400 ;
        RECT 332.400 606.300 334.200 611.400 ;
        RECT 338.400 606.300 340.200 611.400 ;
        RECT 332.400 604.950 340.200 606.300 ;
        RECT 341.400 605.400 343.200 611.400 ;
        RECT 350.400 608.400 352.200 611.400 ;
        RECT 361.800 608.400 363.600 611.400 ;
        RECT 341.400 603.300 342.600 605.400 ;
        RECT 338.850 602.250 342.600 603.300 ;
        RECT 304.950 596.850 307.050 598.950 ;
        RECT 307.950 596.850 310.050 598.950 ;
        RECT 281.700 586.800 282.600 595.050 ;
        RECT 283.950 593.850 286.050 595.950 ;
        RECT 289.950 593.850 292.050 595.950 ;
        RECT 295.950 593.850 298.050 595.950 ;
        RECT 283.950 592.050 285.750 593.850 ;
        RECT 286.950 590.850 289.050 592.950 ;
        RECT 290.100 592.050 291.900 593.850 ;
        RECT 296.250 592.050 298.050 593.850 ;
        RECT 299.850 591.600 301.050 596.850 ;
        RECT 305.100 595.050 306.900 596.850 ;
        RECT 308.100 595.050 309.900 596.850 ;
        RECT 312.000 592.650 313.050 599.850 ;
        RECT 313.950 596.850 316.050 598.950 ;
        RECT 325.950 598.050 328.050 600.150 ;
        RECT 328.950 599.850 331.050 601.950 ;
        RECT 335.100 600.150 336.900 601.950 ;
        RECT 329.100 598.050 330.900 599.850 ;
        RECT 314.100 595.050 315.900 596.850 ;
        RECT 312.000 591.600 314.400 592.650 ;
        RECT 287.100 589.050 288.900 590.850 ;
        RECT 281.700 585.900 288.300 586.800 ;
        RECT 281.700 585.600 282.600 585.900 ;
        RECT 271.800 579.600 273.600 585.600 ;
        RECT 280.800 579.600 282.600 585.600 ;
        RECT 286.800 585.600 288.300 585.900 ;
        RECT 286.800 579.600 288.600 585.600 ;
        RECT 299.700 579.600 301.500 591.600 ;
        RECT 312.600 579.600 314.400 591.600 ;
        RECT 326.400 585.600 327.600 598.050 ;
        RECT 331.950 596.850 334.050 598.950 ;
        RECT 334.950 598.050 337.050 600.150 ;
        RECT 338.850 598.950 340.050 602.250 ;
        RECT 340.950 600.450 343.050 601.050 ;
        RECT 340.950 599.550 345.450 600.450 ;
        RECT 346.950 599.850 349.050 601.950 ;
        RECT 350.400 600.150 351.600 608.400 ;
        RECT 362.400 600.150 363.600 608.400 ;
        RECT 371.400 608.400 373.200 611.400 ;
        RECT 340.950 598.950 343.050 599.550 ;
        RECT 337.950 596.850 340.050 598.950 ;
        RECT 332.100 595.050 333.900 596.850 ;
        RECT 337.950 591.600 339.150 596.850 ;
        RECT 340.950 593.850 343.050 595.950 ;
        RECT 344.550 594.450 345.450 599.550 ;
        RECT 347.100 598.050 348.900 599.850 ;
        RECT 349.950 598.050 352.050 600.150 ;
        RECT 361.950 598.050 364.050 600.150 ;
        RECT 364.950 599.850 367.050 601.950 ;
        RECT 367.950 599.850 370.050 601.950 ;
        RECT 371.400 600.150 372.600 608.400 ;
        RECT 378.150 605.400 379.950 611.400 ;
        RECT 385.950 609.300 387.750 611.400 ;
        RECT 384.000 608.400 387.750 609.300 ;
        RECT 393.750 608.400 395.550 611.400 ;
        RECT 401.550 608.400 403.350 611.400 ;
        RECT 384.000 607.500 385.050 608.400 ;
        RECT 382.950 605.400 385.050 607.500 ;
        RECT 393.750 606.600 394.800 608.400 ;
        RECT 365.100 598.050 366.900 599.850 ;
        RECT 368.100 598.050 369.900 599.850 ;
        RECT 370.950 598.050 373.050 600.150 ;
        RECT 346.950 594.450 349.050 595.050 ;
        RECT 340.950 592.050 342.750 593.850 ;
        RECT 344.550 593.550 349.050 594.450 ;
        RECT 346.950 592.950 349.050 593.550 ;
        RECT 325.800 579.600 327.600 585.600 ;
        RECT 337.500 579.600 339.300 591.600 ;
        RECT 350.400 585.600 351.600 598.050 ;
        RECT 362.400 585.600 363.600 598.050 ;
        RECT 350.400 579.600 352.200 585.600 ;
        RECT 361.800 579.600 363.600 585.600 ;
        RECT 371.400 585.600 372.600 598.050 ;
        RECT 378.150 592.800 379.050 605.400 ;
        RECT 386.550 604.800 388.350 606.600 ;
        RECT 389.850 605.550 394.800 606.600 ;
        RECT 402.300 607.500 403.350 608.400 ;
        RECT 402.300 606.300 406.050 607.500 ;
        RECT 389.850 604.800 391.650 605.550 ;
        RECT 386.850 603.900 387.900 604.800 ;
        RECT 397.050 604.200 398.850 606.000 ;
        RECT 403.950 605.400 406.050 606.300 ;
        RECT 409.650 605.400 411.450 611.400 ;
        RECT 397.050 603.900 397.950 604.200 ;
        RECT 386.850 603.000 397.950 603.900 ;
        RECT 410.250 603.150 411.450 605.400 ;
        RECT 386.850 601.800 387.900 603.000 ;
        RECT 381.000 600.600 387.900 601.800 ;
        RECT 381.000 599.850 381.900 600.600 ;
        RECT 386.100 600.000 387.900 600.600 ;
        RECT 380.100 598.050 381.900 599.850 ;
        RECT 383.100 598.950 384.900 599.700 ;
        RECT 397.050 598.950 397.950 603.000 ;
        RECT 406.950 601.050 411.450 603.150 ;
        RECT 405.150 599.250 409.050 601.050 ;
        RECT 406.950 598.950 409.050 599.250 ;
        RECT 383.100 597.900 391.050 598.950 ;
        RECT 388.950 596.850 391.050 597.900 ;
        RECT 394.950 596.850 397.950 598.950 ;
        RECT 387.450 593.100 389.250 593.400 ;
        RECT 387.450 592.800 395.850 593.100 ;
        RECT 378.150 592.200 395.850 592.800 ;
        RECT 378.150 591.600 389.250 592.200 ;
        RECT 371.400 579.600 373.200 585.600 ;
        RECT 378.150 579.600 379.950 591.600 ;
        RECT 392.250 590.700 394.050 591.300 ;
        RECT 386.550 589.500 394.050 590.700 ;
        RECT 394.950 590.100 395.850 592.200 ;
        RECT 397.050 592.200 397.950 596.850 ;
        RECT 407.250 593.400 409.050 595.200 ;
        RECT 403.950 592.200 408.150 593.400 ;
        RECT 397.050 591.300 403.050 592.200 ;
        RECT 403.950 591.300 406.050 592.200 ;
        RECT 410.250 591.600 411.450 601.050 ;
        RECT 402.150 590.400 403.050 591.300 ;
        RECT 399.450 590.100 401.250 590.400 ;
        RECT 386.550 588.600 387.750 589.500 ;
        RECT 394.950 589.200 401.250 590.100 ;
        RECT 399.450 588.600 401.250 589.200 ;
        RECT 402.150 588.600 404.850 590.400 ;
        RECT 382.950 586.500 387.750 588.600 ;
        RECT 390.450 587.550 392.250 588.300 ;
        RECT 395.250 587.550 397.050 588.300 ;
        RECT 390.450 586.500 397.050 587.550 ;
        RECT 386.550 585.600 387.750 586.500 ;
        RECT 386.550 579.600 388.350 585.600 ;
        RECT 394.350 579.600 396.150 586.500 ;
        RECT 402.150 585.600 406.050 587.700 ;
        RECT 402.150 579.600 403.950 585.600 ;
        RECT 409.650 579.600 411.450 591.600 ;
        RECT 413.550 605.400 415.350 611.400 ;
        RECT 421.650 608.400 423.450 611.400 ;
        RECT 429.450 608.400 431.250 611.400 ;
        RECT 437.250 609.300 439.050 611.400 ;
        RECT 437.250 608.400 441.000 609.300 ;
        RECT 421.650 607.500 422.700 608.400 ;
        RECT 418.950 606.300 422.700 607.500 ;
        RECT 430.200 606.600 431.250 608.400 ;
        RECT 439.950 607.500 441.000 608.400 ;
        RECT 418.950 605.400 421.050 606.300 ;
        RECT 413.550 603.150 414.750 605.400 ;
        RECT 426.150 604.200 427.950 606.000 ;
        RECT 430.200 605.550 435.150 606.600 ;
        RECT 433.350 604.800 435.150 605.550 ;
        RECT 436.650 604.800 438.450 606.600 ;
        RECT 439.950 605.400 442.050 607.500 ;
        RECT 445.050 605.400 446.850 611.400 ;
        RECT 427.050 603.900 427.950 604.200 ;
        RECT 437.100 603.900 438.150 604.800 ;
        RECT 413.550 601.050 418.050 603.150 ;
        RECT 427.050 603.000 438.150 603.900 ;
        RECT 413.550 591.600 414.750 601.050 ;
        RECT 415.950 599.250 419.850 601.050 ;
        RECT 415.950 598.950 418.050 599.250 ;
        RECT 427.050 598.950 427.950 603.000 ;
        RECT 437.100 601.800 438.150 603.000 ;
        RECT 437.100 600.600 444.000 601.800 ;
        RECT 437.100 600.000 438.900 600.600 ;
        RECT 443.100 599.850 444.000 600.600 ;
        RECT 440.100 598.950 441.900 599.700 ;
        RECT 427.050 596.850 430.050 598.950 ;
        RECT 433.950 597.900 441.900 598.950 ;
        RECT 443.100 598.050 444.900 599.850 ;
        RECT 433.950 596.850 436.050 597.900 ;
        RECT 415.950 593.400 417.750 595.200 ;
        RECT 416.850 592.200 421.050 593.400 ;
        RECT 427.050 592.200 427.950 596.850 ;
        RECT 435.750 593.100 437.550 593.400 ;
        RECT 413.550 579.600 415.350 591.600 ;
        RECT 418.950 591.300 421.050 592.200 ;
        RECT 421.950 591.300 427.950 592.200 ;
        RECT 429.150 592.800 437.550 593.100 ;
        RECT 445.950 592.800 446.850 605.400 ;
        RECT 454.200 604.200 456.000 611.400 ;
        RECT 463.800 605.400 465.600 611.400 ;
        RECT 452.400 603.300 456.000 604.200 ;
        RECT 464.400 603.300 465.600 605.400 ;
        RECT 466.800 606.300 468.600 611.400 ;
        RECT 472.800 606.300 474.600 611.400 ;
        RECT 466.800 604.950 474.600 606.300 ;
        RECT 479.400 608.400 481.200 611.400 ;
        RECT 449.100 597.150 450.900 598.950 ;
        RECT 448.950 595.050 451.050 597.150 ;
        RECT 452.400 595.950 453.600 603.300 ;
        RECT 464.400 602.250 468.150 603.300 ;
        RECT 466.950 598.950 468.150 602.250 ;
        RECT 470.100 600.150 471.900 601.950 ;
        RECT 455.100 597.150 456.900 598.950 ;
        RECT 451.950 593.850 454.050 595.950 ;
        RECT 454.950 595.050 457.050 597.150 ;
        RECT 466.950 596.850 469.050 598.950 ;
        RECT 469.950 598.050 472.050 600.150 ;
        RECT 475.950 599.850 478.050 601.950 ;
        RECT 479.400 600.150 480.600 608.400 ;
        RECT 487.500 605.400 489.300 611.400 ;
        RECT 493.800 608.400 495.600 611.400 ;
        RECT 472.950 596.850 475.050 598.950 ;
        RECT 476.100 598.050 477.900 599.850 ;
        RECT 478.950 598.050 481.050 600.150 ;
        RECT 487.800 598.950 489.000 605.400 ;
        RECT 493.800 604.500 495.000 608.400 ;
        RECT 499.500 605.400 501.300 611.400 ;
        RECT 505.800 608.400 507.600 611.400 ;
        RECT 489.900 603.600 495.000 604.500 ;
        RECT 489.900 602.700 491.850 603.600 ;
        RECT 463.950 593.850 466.050 595.950 ;
        RECT 429.150 592.200 446.850 592.800 ;
        RECT 421.950 590.400 422.850 591.300 ;
        RECT 420.150 588.600 422.850 590.400 ;
        RECT 423.750 590.100 425.550 590.400 ;
        RECT 429.150 590.100 430.050 592.200 ;
        RECT 435.750 591.600 446.850 592.200 ;
        RECT 423.750 589.200 430.050 590.100 ;
        RECT 430.950 590.700 432.750 591.300 ;
        RECT 430.950 589.500 438.450 590.700 ;
        RECT 423.750 588.600 425.550 589.200 ;
        RECT 437.250 588.600 438.450 589.500 ;
        RECT 418.950 585.600 422.850 587.700 ;
        RECT 427.950 587.550 429.750 588.300 ;
        RECT 432.750 587.550 434.550 588.300 ;
        RECT 427.950 586.500 434.550 587.550 ;
        RECT 437.250 586.500 442.050 588.600 ;
        RECT 421.050 579.600 422.850 585.600 ;
        RECT 428.850 579.600 430.650 586.500 ;
        RECT 437.250 585.600 438.450 586.500 ;
        RECT 436.650 579.600 438.450 585.600 ;
        RECT 445.050 579.600 446.850 591.600 ;
        RECT 452.400 585.600 453.600 593.850 ;
        RECT 464.250 592.050 466.050 593.850 ;
        RECT 467.850 591.600 469.050 596.850 ;
        RECT 473.100 595.050 474.900 596.850 ;
        RECT 452.400 579.600 454.200 585.600 ;
        RECT 467.700 579.600 469.500 591.600 ;
        RECT 479.400 585.600 480.600 598.050 ;
        RECT 487.800 596.850 490.050 598.950 ;
        RECT 487.800 591.600 489.000 596.850 ;
        RECT 490.950 594.300 491.850 602.700 ;
        RECT 499.800 598.950 501.000 605.400 ;
        RECT 505.800 604.500 507.000 608.400 ;
        RECT 501.900 603.600 507.000 604.500 ;
        RECT 516.000 604.200 517.800 611.400 ;
        RECT 526.800 605.400 528.600 611.400 ;
        RECT 501.900 602.700 503.850 603.600 ;
        RECT 516.000 603.300 519.600 604.200 ;
        RECT 493.950 596.850 496.050 598.950 ;
        RECT 499.800 596.850 502.050 598.950 ;
        RECT 494.100 595.050 495.900 596.850 ;
        RECT 489.900 593.400 491.850 594.300 ;
        RECT 489.900 592.500 495.600 593.400 ;
        RECT 479.400 579.600 481.200 585.600 ;
        RECT 487.500 579.600 489.300 591.600 ;
        RECT 494.400 585.600 495.600 592.500 ;
        RECT 499.800 591.600 501.000 596.850 ;
        RECT 502.950 594.300 503.850 602.700 ;
        RECT 505.950 596.850 508.050 598.950 ;
        RECT 515.100 597.150 516.900 598.950 ;
        RECT 506.100 595.050 507.900 596.850 ;
        RECT 514.950 595.050 517.050 597.150 ;
        RECT 518.400 595.950 519.600 603.300 ;
        RECT 527.400 603.300 528.600 605.400 ;
        RECT 529.800 606.300 531.600 611.400 ;
        RECT 535.800 606.300 537.600 611.400 ;
        RECT 529.800 604.950 537.600 606.300 ;
        RECT 539.550 605.400 541.350 611.400 ;
        RECT 547.650 608.400 549.450 611.400 ;
        RECT 555.450 608.400 557.250 611.400 ;
        RECT 563.250 609.300 565.050 611.400 ;
        RECT 563.250 608.400 567.000 609.300 ;
        RECT 547.650 607.500 548.700 608.400 ;
        RECT 544.950 606.300 548.700 607.500 ;
        RECT 556.200 606.600 557.250 608.400 ;
        RECT 565.950 607.500 567.000 608.400 ;
        RECT 544.950 605.400 547.050 606.300 ;
        RECT 527.400 602.250 531.150 603.300 ;
        RECT 529.950 598.950 531.150 602.250 ;
        RECT 539.550 603.150 540.750 605.400 ;
        RECT 552.150 604.200 553.950 606.000 ;
        RECT 556.200 605.550 561.150 606.600 ;
        RECT 559.350 604.800 561.150 605.550 ;
        RECT 562.650 604.800 564.450 606.600 ;
        RECT 565.950 605.400 568.050 607.500 ;
        RECT 571.050 605.400 572.850 611.400 ;
        RECT 553.050 603.900 553.950 604.200 ;
        RECT 563.100 603.900 564.150 604.800 ;
        RECT 533.100 600.150 534.900 601.950 ;
        RECT 539.550 601.050 544.050 603.150 ;
        RECT 553.050 603.000 564.150 603.900 ;
        RECT 521.100 597.150 522.900 598.950 ;
        RECT 501.900 593.400 503.850 594.300 ;
        RECT 517.950 593.850 520.050 595.950 ;
        RECT 520.950 595.050 523.050 597.150 ;
        RECT 529.950 596.850 532.050 598.950 ;
        RECT 532.950 598.050 535.050 600.150 ;
        RECT 535.950 596.850 538.050 598.950 ;
        RECT 526.950 593.850 529.050 595.950 ;
        RECT 501.900 592.500 507.600 593.400 ;
        RECT 493.800 579.600 495.600 585.600 ;
        RECT 499.500 579.600 501.300 591.600 ;
        RECT 506.400 585.600 507.600 592.500 ;
        RECT 518.400 585.600 519.600 593.850 ;
        RECT 527.250 592.050 529.050 593.850 ;
        RECT 530.850 591.600 532.050 596.850 ;
        RECT 536.100 595.050 537.900 596.850 ;
        RECT 539.550 591.600 540.750 601.050 ;
        RECT 541.950 599.250 545.850 601.050 ;
        RECT 541.950 598.950 544.050 599.250 ;
        RECT 553.050 598.950 553.950 603.000 ;
        RECT 563.100 601.800 564.150 603.000 ;
        RECT 563.100 600.600 570.000 601.800 ;
        RECT 563.100 600.000 564.900 600.600 ;
        RECT 569.100 599.850 570.000 600.600 ;
        RECT 566.100 598.950 567.900 599.700 ;
        RECT 553.050 596.850 556.050 598.950 ;
        RECT 559.950 597.900 567.900 598.950 ;
        RECT 569.100 598.050 570.900 599.850 ;
        RECT 559.950 596.850 562.050 597.900 ;
        RECT 541.950 593.400 543.750 595.200 ;
        RECT 542.850 592.200 547.050 593.400 ;
        RECT 553.050 592.200 553.950 596.850 ;
        RECT 561.750 593.100 563.550 593.400 ;
        RECT 505.800 579.600 507.600 585.600 ;
        RECT 517.800 579.600 519.600 585.600 ;
        RECT 530.700 579.600 532.500 591.600 ;
        RECT 539.550 579.600 541.350 591.600 ;
        RECT 544.950 591.300 547.050 592.200 ;
        RECT 547.950 591.300 553.950 592.200 ;
        RECT 555.150 592.800 563.550 593.100 ;
        RECT 571.950 592.800 572.850 605.400 ;
        RECT 555.150 592.200 572.850 592.800 ;
        RECT 547.950 590.400 548.850 591.300 ;
        RECT 546.150 588.600 548.850 590.400 ;
        RECT 549.750 590.100 551.550 590.400 ;
        RECT 555.150 590.100 556.050 592.200 ;
        RECT 561.750 591.600 572.850 592.200 ;
        RECT 549.750 589.200 556.050 590.100 ;
        RECT 556.950 590.700 558.750 591.300 ;
        RECT 556.950 589.500 564.450 590.700 ;
        RECT 549.750 588.600 551.550 589.200 ;
        RECT 563.250 588.600 564.450 589.500 ;
        RECT 544.950 585.600 548.850 587.700 ;
        RECT 553.950 587.550 555.750 588.300 ;
        RECT 558.750 587.550 560.550 588.300 ;
        RECT 553.950 586.500 560.550 587.550 ;
        RECT 563.250 586.500 568.050 588.600 ;
        RECT 547.050 579.600 548.850 585.600 ;
        RECT 554.850 579.600 556.650 586.500 ;
        RECT 563.250 585.600 564.450 586.500 ;
        RECT 562.650 579.600 564.450 585.600 ;
        RECT 571.050 579.600 572.850 591.600 ;
        RECT 576.150 605.400 577.950 611.400 ;
        RECT 583.950 609.300 585.750 611.400 ;
        RECT 582.000 608.400 585.750 609.300 ;
        RECT 591.750 608.400 593.550 611.400 ;
        RECT 599.550 608.400 601.350 611.400 ;
        RECT 582.000 607.500 583.050 608.400 ;
        RECT 580.950 605.400 583.050 607.500 ;
        RECT 591.750 606.600 592.800 608.400 ;
        RECT 576.150 592.800 577.050 605.400 ;
        RECT 584.550 604.800 586.350 606.600 ;
        RECT 587.850 605.550 592.800 606.600 ;
        RECT 600.300 607.500 601.350 608.400 ;
        RECT 600.300 606.300 604.050 607.500 ;
        RECT 587.850 604.800 589.650 605.550 ;
        RECT 584.850 603.900 585.900 604.800 ;
        RECT 595.050 604.200 596.850 606.000 ;
        RECT 601.950 605.400 604.050 606.300 ;
        RECT 607.650 605.400 609.450 611.400 ;
        RECT 613.800 608.400 615.600 611.400 ;
        RECT 595.050 603.900 595.950 604.200 ;
        RECT 584.850 603.000 595.950 603.900 ;
        RECT 608.250 603.150 609.450 605.400 ;
        RECT 584.850 601.800 585.900 603.000 ;
        RECT 579.000 600.600 585.900 601.800 ;
        RECT 579.000 599.850 579.900 600.600 ;
        RECT 584.100 600.000 585.900 600.600 ;
        RECT 578.100 598.050 579.900 599.850 ;
        RECT 581.100 598.950 582.900 599.700 ;
        RECT 595.050 598.950 595.950 603.000 ;
        RECT 604.950 601.050 609.450 603.150 ;
        RECT 603.150 599.250 607.050 601.050 ;
        RECT 604.950 598.950 607.050 599.250 ;
        RECT 581.100 597.900 589.050 598.950 ;
        RECT 586.950 596.850 589.050 597.900 ;
        RECT 592.950 596.850 595.950 598.950 ;
        RECT 585.450 593.100 587.250 593.400 ;
        RECT 585.450 592.800 593.850 593.100 ;
        RECT 576.150 592.200 593.850 592.800 ;
        RECT 576.150 591.600 587.250 592.200 ;
        RECT 576.150 579.600 577.950 591.600 ;
        RECT 590.250 590.700 592.050 591.300 ;
        RECT 584.550 589.500 592.050 590.700 ;
        RECT 592.950 590.100 593.850 592.200 ;
        RECT 595.050 592.200 595.950 596.850 ;
        RECT 605.250 593.400 607.050 595.200 ;
        RECT 601.950 592.200 606.150 593.400 ;
        RECT 595.050 591.300 601.050 592.200 ;
        RECT 601.950 591.300 604.050 592.200 ;
        RECT 608.250 591.600 609.450 601.050 ;
        RECT 614.400 600.150 615.600 608.400 ;
        RECT 625.500 605.400 627.300 611.400 ;
        RECT 631.800 608.400 633.600 611.400 ;
        RECT 613.950 598.050 616.050 600.150 ;
        RECT 616.950 599.850 619.050 601.950 ;
        RECT 617.100 598.050 618.900 599.850 ;
        RECT 625.800 598.950 627.000 605.400 ;
        RECT 631.800 604.500 633.000 608.400 ;
        RECT 627.900 603.600 633.000 604.500 ;
        RECT 640.200 604.200 642.000 611.400 ;
        RECT 652.800 608.400 654.600 611.400 ;
        RECT 627.900 602.700 629.850 603.600 ;
        RECT 600.150 590.400 601.050 591.300 ;
        RECT 597.450 590.100 599.250 590.400 ;
        RECT 584.550 588.600 585.750 589.500 ;
        RECT 592.950 589.200 599.250 590.100 ;
        RECT 597.450 588.600 599.250 589.200 ;
        RECT 600.150 588.600 602.850 590.400 ;
        RECT 580.950 586.500 585.750 588.600 ;
        RECT 588.450 587.550 590.250 588.300 ;
        RECT 593.250 587.550 595.050 588.300 ;
        RECT 588.450 586.500 595.050 587.550 ;
        RECT 584.550 585.600 585.750 586.500 ;
        RECT 584.550 579.600 586.350 585.600 ;
        RECT 592.350 579.600 594.150 586.500 ;
        RECT 600.150 585.600 604.050 587.700 ;
        RECT 600.150 579.600 601.950 585.600 ;
        RECT 607.650 579.600 609.450 591.600 ;
        RECT 614.400 585.600 615.600 598.050 ;
        RECT 625.800 596.850 628.050 598.950 ;
        RECT 625.800 591.600 627.000 596.850 ;
        RECT 628.950 594.300 629.850 602.700 ;
        RECT 638.400 603.300 642.000 604.200 ;
        RECT 631.950 596.850 634.050 598.950 ;
        RECT 635.100 597.150 636.900 598.950 ;
        RECT 632.100 595.050 633.900 596.850 ;
        RECT 634.950 595.050 637.050 597.150 ;
        RECT 638.400 595.950 639.600 603.300 ;
        RECT 652.950 601.950 654.000 608.400 ;
        RECT 664.200 607.050 666.000 611.400 ;
        RECT 664.200 605.400 669.600 607.050 ;
        RECT 652.950 599.850 655.050 601.950 ;
        RECT 659.100 600.150 660.900 601.950 ;
        RECT 641.100 597.150 642.900 598.950 ;
        RECT 627.900 593.400 629.850 594.300 ;
        RECT 637.950 593.850 640.050 595.950 ;
        RECT 640.950 595.050 643.050 597.150 ;
        RECT 649.950 596.850 652.050 598.950 ;
        RECT 650.100 595.050 651.900 596.850 ;
        RECT 627.900 592.500 633.600 593.400 ;
        RECT 613.800 579.600 615.600 585.600 ;
        RECT 625.500 579.600 627.300 591.600 ;
        RECT 632.400 585.600 633.600 592.500 ;
        RECT 631.800 579.600 633.600 585.600 ;
        RECT 638.400 585.600 639.600 593.850 ;
        RECT 652.950 592.650 654.000 599.850 ;
        RECT 655.950 596.850 658.050 598.950 ;
        RECT 658.950 598.050 661.050 600.150 ;
        RECT 661.950 599.850 664.050 601.950 ;
        RECT 665.100 600.150 666.900 601.950 ;
        RECT 662.100 598.050 663.900 599.850 ;
        RECT 664.950 598.050 667.050 600.150 ;
        RECT 668.700 598.950 669.600 605.400 ;
        RECT 674.400 606.300 676.200 611.400 ;
        RECT 680.400 606.300 682.200 611.400 ;
        RECT 674.400 604.950 682.200 606.300 ;
        RECT 683.400 605.400 685.200 611.400 ;
        RECT 691.800 608.400 693.600 611.400 ;
        RECT 701.400 608.400 703.200 611.400 ;
        RECT 713.400 608.400 715.200 611.400 ;
        RECT 725.400 608.400 727.200 611.400 ;
        RECT 683.400 603.300 684.600 605.400 ;
        RECT 680.850 602.250 684.600 603.300 ;
        RECT 677.100 600.150 678.900 601.950 ;
        RECT 667.950 596.850 670.050 598.950 ;
        RECT 673.950 596.850 676.050 598.950 ;
        RECT 676.950 598.050 679.050 600.150 ;
        RECT 680.850 598.950 682.050 602.250 ;
        RECT 692.400 600.150 693.600 608.400 ;
        RECT 702.000 601.950 703.050 608.400 ;
        RECT 679.950 596.850 682.050 598.950 ;
        RECT 691.950 598.050 694.050 600.150 ;
        RECT 694.950 599.850 697.050 601.950 ;
        RECT 700.950 599.850 703.050 601.950 ;
        RECT 709.950 599.850 712.050 601.950 ;
        RECT 713.400 600.150 714.600 608.400 ;
        RECT 726.000 601.950 727.050 608.400 ;
        RECT 734.400 606.300 736.200 611.400 ;
        RECT 740.400 606.300 742.200 611.400 ;
        RECT 734.400 604.950 742.200 606.300 ;
        RECT 743.400 605.400 745.200 611.400 ;
        RECT 754.200 607.050 756.000 611.400 ;
        RECT 754.200 605.400 759.600 607.050 ;
        RECT 743.400 603.300 744.600 605.400 ;
        RECT 740.850 602.250 744.600 603.300 ;
        RECT 695.100 598.050 696.900 599.850 ;
        RECT 656.100 595.050 657.900 596.850 ;
        RECT 651.600 591.600 654.000 592.650 ;
        RECT 668.700 591.600 669.600 596.850 ;
        RECT 674.100 595.050 675.900 596.850 ;
        RECT 679.950 591.600 681.150 596.850 ;
        RECT 682.950 593.850 685.050 595.950 ;
        RECT 682.950 592.050 684.750 593.850 ;
        RECT 638.400 579.600 640.200 585.600 ;
        RECT 651.600 579.600 653.400 591.600 ;
        RECT 659.400 590.700 667.200 591.600 ;
        RECT 659.400 579.600 661.200 590.700 ;
        RECT 665.400 579.600 667.200 590.700 ;
        RECT 668.400 579.600 670.200 591.600 ;
        RECT 679.500 579.600 681.300 591.600 ;
        RECT 692.400 585.600 693.600 598.050 ;
        RECT 697.950 596.850 700.050 598.950 ;
        RECT 698.100 595.050 699.900 596.850 ;
        RECT 702.000 592.650 703.050 599.850 ;
        RECT 703.950 596.850 706.050 598.950 ;
        RECT 710.100 598.050 711.900 599.850 ;
        RECT 712.950 598.050 715.050 600.150 ;
        RECT 724.950 599.850 727.050 601.950 ;
        RECT 737.100 600.150 738.900 601.950 ;
        RECT 704.100 595.050 705.900 596.850 ;
        RECT 702.000 591.600 704.400 592.650 ;
        RECT 691.800 579.600 693.600 585.600 ;
        RECT 702.600 579.600 704.400 591.600 ;
        RECT 713.400 585.600 714.600 598.050 ;
        RECT 721.950 596.850 724.050 598.950 ;
        RECT 722.100 595.050 723.900 596.850 ;
        RECT 726.000 592.650 727.050 599.850 ;
        RECT 727.950 596.850 730.050 598.950 ;
        RECT 733.950 596.850 736.050 598.950 ;
        RECT 736.950 598.050 739.050 600.150 ;
        RECT 740.850 598.950 742.050 602.250 ;
        RECT 749.100 600.150 750.900 601.950 ;
        RECT 739.950 596.850 742.050 598.950 ;
        RECT 748.950 598.050 751.050 600.150 ;
        RECT 751.950 599.850 754.050 601.950 ;
        RECT 755.100 600.150 756.900 601.950 ;
        RECT 752.100 598.050 753.900 599.850 ;
        RECT 754.950 598.050 757.050 600.150 ;
        RECT 758.700 598.950 759.600 605.400 ;
        RECT 757.950 596.850 760.050 598.950 ;
        RECT 728.100 595.050 729.900 596.850 ;
        RECT 734.100 595.050 735.900 596.850 ;
        RECT 726.000 591.600 728.400 592.650 ;
        RECT 739.950 591.600 741.150 596.850 ;
        RECT 742.950 593.850 745.050 595.950 ;
        RECT 742.950 592.050 744.750 593.850 ;
        RECT 758.700 591.600 759.600 596.850 ;
        RECT 713.400 579.600 715.200 585.600 ;
        RECT 726.600 579.600 728.400 591.600 ;
        RECT 739.500 579.600 741.300 591.600 ;
        RECT 749.400 590.700 757.200 591.600 ;
        RECT 749.400 579.600 751.200 590.700 ;
        RECT 755.400 579.600 757.200 590.700 ;
        RECT 758.400 579.600 760.200 591.600 ;
        RECT 4.500 563.400 6.300 575.400 ;
        RECT 10.800 569.400 12.600 575.400 ;
        RECT 4.800 558.150 6.000 563.400 ;
        RECT 11.400 562.500 12.600 569.400 ;
        RECT 23.700 563.400 25.500 575.400 ;
        RECT 37.500 563.400 39.300 575.400 ;
        RECT 49.800 563.400 51.600 575.400 ;
        RECT 52.800 564.300 54.600 575.400 ;
        RECT 58.800 564.300 60.600 575.400 ;
        RECT 52.800 563.400 60.600 564.300 ;
        RECT 67.500 563.400 69.300 575.400 ;
        RECT 77.400 564.300 79.200 575.400 ;
        RECT 83.400 564.300 85.200 575.400 ;
        RECT 77.400 563.400 85.200 564.300 ;
        RECT 86.400 563.400 88.200 575.400 ;
        RECT 98.700 563.400 100.500 575.400 ;
        RECT 113.700 563.400 115.500 575.400 ;
        RECT 130.500 563.400 132.300 575.400 ;
        RECT 146.700 563.400 148.500 575.400 ;
        RECT 157.800 563.400 159.600 575.400 ;
        RECT 160.800 564.300 162.600 575.400 ;
        RECT 166.800 564.300 168.600 575.400 ;
        RECT 160.800 563.400 168.600 564.300 ;
        RECT 175.500 563.400 177.300 575.400 ;
        RECT 190.800 569.400 192.600 575.400 ;
        RECT 6.900 561.600 12.600 562.500 ;
        RECT 6.900 560.700 8.850 561.600 ;
        RECT 20.250 561.150 22.050 562.950 ;
        RECT 4.800 556.050 7.050 558.150 ;
        RECT 4.800 549.600 6.000 556.050 ;
        RECT 7.950 552.300 8.850 560.700 ;
        RECT 11.100 558.150 12.900 559.950 ;
        RECT 19.950 559.050 22.050 561.150 ;
        RECT 23.850 558.150 25.050 563.400 ;
        RECT 29.100 558.150 30.900 559.950 ;
        RECT 32.100 558.150 33.900 559.950 ;
        RECT 37.950 558.150 39.150 563.400 ;
        RECT 40.950 561.150 42.750 562.950 ;
        RECT 40.950 559.050 43.050 561.150 ;
        RECT 50.400 558.150 51.300 563.400 ;
        RECT 62.100 558.150 63.900 559.950 ;
        RECT 67.950 558.150 69.150 563.400 ;
        RECT 70.950 561.150 72.750 562.950 ;
        RECT 70.950 559.050 73.050 561.150 ;
        RECT 86.700 558.150 87.600 563.400 ;
        RECT 95.250 561.150 97.050 562.950 ;
        RECT 94.950 559.050 97.050 561.150 ;
        RECT 98.850 558.150 100.050 563.400 ;
        RECT 110.250 561.150 112.050 562.950 ;
        RECT 104.100 558.150 105.900 559.950 ;
        RECT 109.950 559.050 112.050 561.150 ;
        RECT 113.850 558.150 115.050 563.400 ;
        RECT 121.950 559.950 124.050 562.050 ;
        RECT 119.100 558.150 120.900 559.950 ;
        RECT 10.950 556.050 13.050 558.150 ;
        RECT 22.950 556.050 25.050 558.150 ;
        RECT 22.950 552.750 24.150 556.050 ;
        RECT 25.950 554.850 28.050 556.950 ;
        RECT 28.950 556.050 31.050 558.150 ;
        RECT 31.950 556.050 34.050 558.150 ;
        RECT 34.950 554.850 37.050 556.950 ;
        RECT 37.950 556.050 40.050 558.150 ;
        RECT 49.950 556.050 52.050 558.150 ;
        RECT 26.100 553.050 27.900 554.850 ;
        RECT 35.100 553.050 36.900 554.850 ;
        RECT 6.900 551.400 8.850 552.300 ;
        RECT 20.400 551.700 24.150 552.750 ;
        RECT 38.850 552.750 40.050 556.050 ;
        RECT 38.850 551.700 42.600 552.750 ;
        RECT 6.900 550.500 12.000 551.400 ;
        RECT 4.500 543.600 6.300 549.600 ;
        RECT 10.800 546.600 12.000 550.500 ;
        RECT 20.400 549.600 21.600 551.700 ;
        RECT 10.800 543.600 12.600 546.600 ;
        RECT 19.800 543.600 21.600 549.600 ;
        RECT 22.800 548.700 30.600 550.050 ;
        RECT 22.800 543.600 24.600 548.700 ;
        RECT 28.800 543.600 30.600 548.700 ;
        RECT 32.400 548.700 40.200 550.050 ;
        RECT 32.400 543.600 34.200 548.700 ;
        RECT 38.400 543.600 40.200 548.700 ;
        RECT 41.400 549.600 42.600 551.700 ;
        RECT 50.400 549.600 51.300 556.050 ;
        RECT 52.950 554.850 55.050 556.950 ;
        RECT 56.100 555.150 57.900 556.950 ;
        RECT 53.100 553.050 54.900 554.850 ;
        RECT 55.950 553.050 58.050 555.150 ;
        RECT 58.950 554.850 61.050 556.950 ;
        RECT 61.950 556.050 64.050 558.150 ;
        RECT 64.950 554.850 67.050 556.950 ;
        RECT 67.950 556.050 70.050 558.150 ;
        RECT 59.100 553.050 60.900 554.850 ;
        RECT 65.100 553.050 66.900 554.850 ;
        RECT 68.850 552.750 70.050 556.050 ;
        RECT 76.950 554.850 79.050 556.950 ;
        RECT 80.100 555.150 81.900 556.950 ;
        RECT 77.100 553.050 78.900 554.850 ;
        RECT 79.950 553.050 82.050 555.150 ;
        RECT 82.950 554.850 85.050 556.950 ;
        RECT 85.950 556.050 88.050 558.150 ;
        RECT 97.950 556.050 100.050 558.150 ;
        RECT 83.100 553.050 84.900 554.850 ;
        RECT 68.850 551.700 72.600 552.750 ;
        RECT 41.400 543.600 43.200 549.600 ;
        RECT 50.400 547.950 55.800 549.600 ;
        RECT 54.000 543.600 55.800 547.950 ;
        RECT 62.400 548.700 70.200 550.050 ;
        RECT 62.400 543.600 64.200 548.700 ;
        RECT 68.400 543.600 70.200 548.700 ;
        RECT 71.400 549.600 72.600 551.700 ;
        RECT 86.700 549.600 87.600 556.050 ;
        RECT 97.950 552.750 99.150 556.050 ;
        RECT 100.950 554.850 103.050 556.950 ;
        RECT 103.950 556.050 106.050 558.150 ;
        RECT 112.950 556.050 115.050 558.150 ;
        RECT 101.100 553.050 102.900 554.850 ;
        RECT 112.950 552.750 114.150 556.050 ;
        RECT 115.950 554.850 118.050 556.950 ;
        RECT 118.950 556.050 121.050 558.150 ;
        RECT 116.100 553.050 117.900 554.850 ;
        RECT 95.400 551.700 99.150 552.750 ;
        RECT 110.400 551.700 114.150 552.750 ;
        RECT 122.550 552.450 123.450 559.950 ;
        RECT 125.100 558.150 126.900 559.950 ;
        RECT 130.950 558.150 132.150 563.400 ;
        RECT 133.950 561.150 135.750 562.950 ;
        RECT 143.250 561.150 145.050 562.950 ;
        RECT 133.950 559.050 136.050 561.150 ;
        RECT 142.950 559.050 145.050 561.150 ;
        RECT 146.850 558.150 148.050 563.400 ;
        RECT 152.100 558.150 153.900 559.950 ;
        RECT 158.400 558.150 159.300 563.400 ;
        RECT 170.100 558.150 171.900 559.950 ;
        RECT 175.950 558.150 177.150 563.400 ;
        RECT 178.950 561.150 180.750 562.950 ;
        RECT 191.400 561.150 192.600 569.400 ;
        RECT 201.600 563.400 203.400 575.400 ;
        RECT 217.800 569.400 219.600 575.400 ;
        RECT 201.600 562.350 204.000 563.400 ;
        RECT 178.950 559.050 181.050 561.150 ;
        RECT 124.950 556.050 127.050 558.150 ;
        RECT 127.950 554.850 130.050 556.950 ;
        RECT 130.950 556.050 133.050 558.150 ;
        RECT 128.100 553.050 129.900 554.850 ;
        RECT 124.950 552.450 127.050 553.050 ;
        RECT 95.400 549.600 96.600 551.700 ;
        RECT 71.400 543.600 73.200 549.600 ;
        RECT 82.200 547.950 87.600 549.600 ;
        RECT 82.200 543.600 84.000 547.950 ;
        RECT 94.800 543.600 96.600 549.600 ;
        RECT 97.800 548.700 105.600 550.050 ;
        RECT 110.400 549.600 111.600 551.700 ;
        RECT 122.550 551.550 127.050 552.450 ;
        RECT 131.850 552.750 133.050 556.050 ;
        RECT 145.950 556.050 148.050 558.150 ;
        RECT 145.950 552.750 147.150 556.050 ;
        RECT 148.950 554.850 151.050 556.950 ;
        RECT 151.950 556.050 154.050 558.150 ;
        RECT 157.950 556.050 160.050 558.150 ;
        RECT 149.100 553.050 150.900 554.850 ;
        RECT 131.850 551.700 135.600 552.750 ;
        RECT 124.950 550.950 127.050 551.550 ;
        RECT 97.800 543.600 99.600 548.700 ;
        RECT 103.800 543.600 105.600 548.700 ;
        RECT 109.800 543.600 111.600 549.600 ;
        RECT 112.800 548.700 120.600 550.050 ;
        RECT 112.800 543.600 114.600 548.700 ;
        RECT 118.800 543.600 120.600 548.700 ;
        RECT 125.400 548.700 133.200 550.050 ;
        RECT 125.400 543.600 127.200 548.700 ;
        RECT 131.400 543.600 133.200 548.700 ;
        RECT 134.400 549.600 135.600 551.700 ;
        RECT 143.400 551.700 147.150 552.750 ;
        RECT 143.400 549.600 144.600 551.700 ;
        RECT 134.400 543.600 136.200 549.600 ;
        RECT 142.800 543.600 144.600 549.600 ;
        RECT 145.800 548.700 153.600 550.050 ;
        RECT 145.800 543.600 147.600 548.700 ;
        RECT 151.800 543.600 153.600 548.700 ;
        RECT 158.400 549.600 159.300 556.050 ;
        RECT 160.950 554.850 163.050 556.950 ;
        RECT 164.100 555.150 165.900 556.950 ;
        RECT 161.100 553.050 162.900 554.850 ;
        RECT 163.950 553.050 166.050 555.150 ;
        RECT 166.950 554.850 169.050 556.950 ;
        RECT 169.950 556.050 172.050 558.150 ;
        RECT 172.950 554.850 175.050 556.950 ;
        RECT 175.950 556.050 178.050 558.150 ;
        RECT 187.950 557.850 190.050 559.950 ;
        RECT 190.950 559.050 193.050 561.150 ;
        RECT 188.100 556.050 189.900 557.850 ;
        RECT 167.100 553.050 168.900 554.850 ;
        RECT 173.100 553.050 174.900 554.850 ;
        RECT 176.850 552.750 178.050 556.050 ;
        RECT 176.850 551.700 180.600 552.750 ;
        RECT 191.400 551.700 192.600 559.050 ;
        RECT 193.950 557.850 196.050 559.950 ;
        RECT 200.100 558.150 201.900 559.950 ;
        RECT 194.100 556.050 195.900 557.850 ;
        RECT 199.950 556.050 202.050 558.150 ;
        RECT 158.400 547.950 163.800 549.600 ;
        RECT 162.000 543.600 163.800 547.950 ;
        RECT 170.400 548.700 178.200 550.050 ;
        RECT 170.400 543.600 172.200 548.700 ;
        RECT 176.400 543.600 178.200 548.700 ;
        RECT 179.400 549.600 180.600 551.700 ;
        RECT 189.000 550.800 192.600 551.700 ;
        RECT 202.950 555.150 204.000 562.350 ;
        RECT 218.400 561.150 219.600 569.400 ;
        RECT 230.700 563.400 232.500 575.400 ;
        RECT 239.400 564.600 241.200 575.400 ;
        RECT 245.400 574.500 253.200 575.400 ;
        RECT 245.400 564.600 247.200 574.500 ;
        RECT 239.400 563.700 247.200 564.600 ;
        RECT 227.250 561.150 229.050 562.950 ;
        RECT 206.100 558.150 207.900 559.950 ;
        RECT 205.950 556.050 208.050 558.150 ;
        RECT 214.950 557.850 217.050 559.950 ;
        RECT 217.950 559.050 220.050 561.150 ;
        RECT 215.100 556.050 216.900 557.850 ;
        RECT 202.950 553.050 205.050 555.150 ;
        RECT 179.400 543.600 181.200 549.600 ;
        RECT 189.000 543.600 190.800 550.800 ;
        RECT 202.950 546.600 204.000 553.050 ;
        RECT 218.400 551.700 219.600 559.050 ;
        RECT 220.950 557.850 223.050 559.950 ;
        RECT 226.950 559.050 229.050 561.150 ;
        RECT 230.850 558.150 232.050 563.400 ;
        RECT 248.400 562.500 250.200 573.600 ;
        RECT 251.400 563.400 253.200 574.500 ;
        RECT 260.400 569.400 262.200 575.400 ;
        RECT 246.150 561.600 250.200 562.500 ;
        RECT 236.100 558.150 237.900 559.950 ;
        RECT 239.250 558.150 241.050 559.950 ;
        RECT 246.150 558.150 247.050 561.600 ;
        RECT 260.400 561.150 261.600 569.400 ;
        RECT 277.500 563.400 279.300 575.400 ;
        RECT 289.200 563.400 291.000 575.400 ;
        RECT 295.800 569.400 297.600 575.400 ;
        RECT 251.100 558.150 252.900 559.950 ;
        RECT 221.100 556.050 222.900 557.850 ;
        RECT 229.950 556.050 232.050 558.150 ;
        RECT 229.950 552.750 231.150 556.050 ;
        RECT 232.950 554.850 235.050 556.950 ;
        RECT 235.950 556.050 238.050 558.150 ;
        RECT 238.950 556.050 241.050 558.150 ;
        RECT 241.950 554.850 244.050 556.950 ;
        RECT 233.100 553.050 234.900 554.850 ;
        RECT 242.250 553.050 244.050 554.850 ;
        RECT 244.950 556.050 247.050 558.150 ;
        RECT 216.000 550.800 219.600 551.700 ;
        RECT 227.400 551.700 231.150 552.750 ;
        RECT 202.800 543.600 204.600 546.600 ;
        RECT 216.000 543.600 217.800 550.800 ;
        RECT 227.400 549.600 228.600 551.700 ;
        RECT 226.800 543.600 228.600 549.600 ;
        RECT 229.800 548.700 237.600 550.050 ;
        RECT 244.950 549.600 246.000 556.050 ;
        RECT 247.950 554.850 250.050 556.950 ;
        RECT 250.950 556.050 253.050 558.150 ;
        RECT 256.950 557.850 259.050 559.950 ;
        RECT 259.950 559.050 262.050 561.150 ;
        RECT 257.100 556.050 258.900 557.850 ;
        RECT 247.950 553.050 249.750 554.850 ;
        RECT 250.950 552.450 253.050 553.050 ;
        RECT 256.950 552.450 259.050 553.050 ;
        RECT 250.950 551.550 259.050 552.450 ;
        RECT 250.950 550.950 253.050 551.550 ;
        RECT 256.950 550.950 259.050 551.550 ;
        RECT 260.400 551.700 261.600 559.050 ;
        RECT 262.950 557.850 265.050 559.950 ;
        RECT 272.100 558.150 273.900 559.950 ;
        RECT 277.950 558.150 279.150 563.400 ;
        RECT 280.950 561.150 282.750 562.950 ;
        RECT 280.950 559.050 283.050 561.150 ;
        RECT 289.950 558.150 291.000 563.400 ;
        RECT 263.100 556.050 264.900 557.850 ;
        RECT 271.950 556.050 274.050 558.150 ;
        RECT 274.950 554.850 277.050 556.950 ;
        RECT 277.950 556.050 280.050 558.150 ;
        RECT 275.100 553.050 276.900 554.850 ;
        RECT 278.850 552.750 280.050 556.050 ;
        RECT 289.950 556.050 292.050 558.150 ;
        RECT 292.950 557.850 295.050 559.950 ;
        RECT 293.100 556.050 294.900 557.850 ;
        RECT 278.850 551.700 282.600 552.750 ;
        RECT 260.400 550.800 264.000 551.700 ;
        RECT 229.800 543.600 231.600 548.700 ;
        RECT 235.800 543.600 237.600 548.700 ;
        RECT 244.200 543.600 246.000 549.600 ;
        RECT 262.200 543.600 264.000 550.800 ;
        RECT 272.400 548.700 280.200 550.050 ;
        RECT 272.400 543.600 274.200 548.700 ;
        RECT 278.400 543.600 280.200 548.700 ;
        RECT 281.400 549.600 282.600 551.700 ;
        RECT 289.950 549.600 291.000 556.050 ;
        RECT 296.400 552.300 297.450 569.400 ;
        RECT 304.800 563.400 306.600 575.400 ;
        RECT 316.500 563.400 318.300 575.400 ;
        RECT 328.500 563.400 330.300 575.400 ;
        RECT 334.800 569.400 336.600 575.400 ;
        RECT 299.100 558.150 300.900 559.950 ;
        RECT 305.400 558.150 306.600 563.400 ;
        RECT 311.100 558.150 312.900 559.950 ;
        RECT 316.950 558.150 318.150 563.400 ;
        RECT 319.950 561.150 321.750 562.950 ;
        RECT 319.950 559.050 322.050 561.150 ;
        RECT 328.800 558.150 330.000 563.400 ;
        RECT 335.400 562.500 336.600 569.400 ;
        RECT 330.900 561.600 336.600 562.500 ;
        RECT 338.550 563.400 340.350 575.400 ;
        RECT 346.050 569.400 347.850 575.400 ;
        RECT 343.950 567.300 347.850 569.400 ;
        RECT 353.850 568.500 355.650 575.400 ;
        RECT 361.650 569.400 363.450 575.400 ;
        RECT 362.250 568.500 363.450 569.400 ;
        RECT 352.950 567.450 359.550 568.500 ;
        RECT 352.950 566.700 354.750 567.450 ;
        RECT 357.750 566.700 359.550 567.450 ;
        RECT 362.250 566.400 367.050 568.500 ;
        RECT 345.150 564.600 347.850 566.400 ;
        RECT 348.750 565.800 350.550 566.400 ;
        RECT 348.750 564.900 355.050 565.800 ;
        RECT 362.250 565.500 363.450 566.400 ;
        RECT 348.750 564.600 350.550 564.900 ;
        RECT 346.950 563.700 347.850 564.600 ;
        RECT 330.900 560.700 332.850 561.600 ;
        RECT 298.950 556.050 301.050 558.150 ;
        RECT 304.950 556.050 307.050 558.150 ;
        RECT 293.100 551.100 300.600 552.300 ;
        RECT 293.100 550.500 294.900 551.100 ;
        RECT 281.400 543.600 283.200 549.600 ;
        RECT 289.950 548.100 293.100 549.600 ;
        RECT 291.300 543.600 293.100 548.100 ;
        RECT 298.800 543.600 300.600 551.100 ;
        RECT 305.400 549.600 306.600 556.050 ;
        RECT 307.950 554.850 310.050 556.950 ;
        RECT 310.950 556.050 313.050 558.150 ;
        RECT 313.950 554.850 316.050 556.950 ;
        RECT 316.950 556.050 319.050 558.150 ;
        RECT 308.100 553.050 309.900 554.850 ;
        RECT 314.100 553.050 315.900 554.850 ;
        RECT 317.850 552.750 319.050 556.050 ;
        RECT 328.800 556.050 331.050 558.150 ;
        RECT 317.850 551.700 321.600 552.750 ;
        RECT 304.800 543.600 306.600 549.600 ;
        RECT 311.400 548.700 319.200 550.050 ;
        RECT 311.400 543.600 313.200 548.700 ;
        RECT 317.400 543.600 319.200 548.700 ;
        RECT 320.400 549.600 321.600 551.700 ;
        RECT 328.800 549.600 330.000 556.050 ;
        RECT 331.950 552.300 332.850 560.700 ;
        RECT 335.100 558.150 336.900 559.950 ;
        RECT 334.950 556.050 337.050 558.150 ;
        RECT 330.900 551.400 332.850 552.300 ;
        RECT 338.550 553.950 339.750 563.400 ;
        RECT 343.950 562.800 346.050 563.700 ;
        RECT 346.950 562.800 352.950 563.700 ;
        RECT 341.850 561.600 346.050 562.800 ;
        RECT 340.950 559.800 342.750 561.600 ;
        RECT 352.050 558.150 352.950 562.800 ;
        RECT 354.150 562.800 355.050 564.900 ;
        RECT 355.950 564.300 363.450 565.500 ;
        RECT 355.950 563.700 357.750 564.300 ;
        RECT 370.050 563.400 371.850 575.400 ;
        RECT 360.750 562.800 371.850 563.400 ;
        RECT 354.150 562.200 371.850 562.800 ;
        RECT 354.150 561.900 362.550 562.200 ;
        RECT 360.750 561.600 362.550 561.900 ;
        RECT 352.050 556.050 355.050 558.150 ;
        RECT 358.950 557.100 361.050 558.150 ;
        RECT 358.950 556.050 366.900 557.100 ;
        RECT 340.950 555.750 343.050 556.050 ;
        RECT 340.950 553.950 344.850 555.750 ;
        RECT 338.550 551.850 343.050 553.950 ;
        RECT 352.050 552.000 352.950 556.050 ;
        RECT 365.100 555.300 366.900 556.050 ;
        RECT 368.100 555.150 369.900 556.950 ;
        RECT 362.100 554.400 363.900 555.000 ;
        RECT 368.100 554.400 369.000 555.150 ;
        RECT 362.100 553.200 369.000 554.400 ;
        RECT 362.100 552.000 363.150 553.200 ;
        RECT 330.900 550.500 336.000 551.400 ;
        RECT 320.400 543.600 322.200 549.600 ;
        RECT 328.500 543.600 330.300 549.600 ;
        RECT 334.800 546.600 336.000 550.500 ;
        RECT 338.550 549.600 339.750 551.850 ;
        RECT 352.050 551.100 363.150 552.000 ;
        RECT 352.050 550.800 352.950 551.100 ;
        RECT 334.800 543.600 336.600 546.600 ;
        RECT 338.550 543.600 340.350 549.600 ;
        RECT 343.950 548.700 346.050 549.600 ;
        RECT 351.150 549.000 352.950 550.800 ;
        RECT 362.100 550.200 363.150 551.100 ;
        RECT 358.350 549.450 360.150 550.200 ;
        RECT 343.950 547.500 347.700 548.700 ;
        RECT 346.650 546.600 347.700 547.500 ;
        RECT 355.200 548.400 360.150 549.450 ;
        RECT 361.650 548.400 363.450 550.200 ;
        RECT 370.950 549.600 371.850 562.200 ;
        RECT 377.400 569.400 379.200 575.400 ;
        RECT 377.400 556.950 378.600 569.400 ;
        RECT 388.500 563.400 390.300 575.400 ;
        RECT 404.400 569.400 406.200 575.400 ;
        RECT 383.100 558.150 384.900 559.950 ;
        RECT 388.950 558.150 390.150 563.400 ;
        RECT 391.950 561.150 393.750 562.950 ;
        RECT 404.400 561.150 405.600 569.400 ;
        RECT 419.700 563.400 421.500 575.400 ;
        RECT 436.500 563.400 438.300 575.400 ;
        RECT 451.800 569.400 453.600 575.400 ;
        RECT 391.950 559.050 394.050 561.150 ;
        RECT 374.100 555.150 375.900 556.950 ;
        RECT 373.950 553.050 376.050 555.150 ;
        RECT 376.950 554.850 379.050 556.950 ;
        RECT 382.950 556.050 385.050 558.150 ;
        RECT 385.950 554.850 388.050 556.950 ;
        RECT 388.950 556.050 391.050 558.150 ;
        RECT 400.950 557.850 403.050 559.950 ;
        RECT 403.950 559.050 406.050 561.150 ;
        RECT 412.950 559.950 415.050 562.050 ;
        RECT 416.250 561.150 418.050 562.950 ;
        RECT 401.100 556.050 402.900 557.850 ;
        RECT 355.200 546.600 356.250 548.400 ;
        RECT 364.950 547.500 367.050 549.600 ;
        RECT 364.950 546.600 366.000 547.500 ;
        RECT 346.650 543.600 348.450 546.600 ;
        RECT 354.450 543.600 356.250 546.600 ;
        RECT 362.250 545.700 366.000 546.600 ;
        RECT 362.250 543.600 364.050 545.700 ;
        RECT 370.050 543.600 371.850 549.600 ;
        RECT 377.400 546.600 378.600 554.850 ;
        RECT 386.100 553.050 387.900 554.850 ;
        RECT 389.850 552.750 391.050 556.050 ;
        RECT 389.850 551.700 393.600 552.750 ;
        RECT 383.400 548.700 391.200 550.050 ;
        RECT 377.400 543.600 379.200 546.600 ;
        RECT 383.400 543.600 385.200 548.700 ;
        RECT 389.400 543.600 391.200 548.700 ;
        RECT 392.400 549.600 393.600 551.700 ;
        RECT 404.400 551.700 405.600 559.050 ;
        RECT 406.950 557.850 409.050 559.950 ;
        RECT 407.100 556.050 408.900 557.850 ;
        RECT 413.550 556.050 414.450 559.950 ;
        RECT 415.950 559.050 418.050 561.150 ;
        RECT 419.850 558.150 421.050 563.400 ;
        RECT 425.100 558.150 426.900 559.950 ;
        RECT 431.100 558.150 432.900 559.950 ;
        RECT 436.950 558.150 438.150 563.400 ;
        RECT 439.950 561.150 441.750 562.950 ;
        RECT 452.400 561.150 453.600 569.400 ;
        RECT 459.150 563.400 460.950 575.400 ;
        RECT 467.550 569.400 469.350 575.400 ;
        RECT 467.550 568.500 468.750 569.400 ;
        RECT 475.350 568.500 477.150 575.400 ;
        RECT 483.150 569.400 484.950 575.400 ;
        RECT 463.950 566.400 468.750 568.500 ;
        RECT 471.450 567.450 478.050 568.500 ;
        RECT 471.450 566.700 473.250 567.450 ;
        RECT 476.250 566.700 478.050 567.450 ;
        RECT 483.150 567.300 487.050 569.400 ;
        RECT 467.550 565.500 468.750 566.400 ;
        RECT 480.450 565.800 482.250 566.400 ;
        RECT 467.550 564.300 475.050 565.500 ;
        RECT 473.250 563.700 475.050 564.300 ;
        RECT 475.950 564.900 482.250 565.800 ;
        RECT 459.150 562.800 470.250 563.400 ;
        RECT 475.950 562.800 476.850 564.900 ;
        RECT 480.450 564.600 482.250 564.900 ;
        RECT 483.150 564.600 485.850 566.400 ;
        RECT 483.150 563.700 484.050 564.600 ;
        RECT 459.150 562.200 476.850 562.800 ;
        RECT 439.950 559.050 442.050 561.150 ;
        RECT 418.950 556.050 421.050 558.150 ;
        RECT 412.950 553.950 415.050 556.050 ;
        RECT 418.950 552.750 420.150 556.050 ;
        RECT 421.950 554.850 424.050 556.950 ;
        RECT 424.950 556.050 427.050 558.150 ;
        RECT 430.950 556.050 433.050 558.150 ;
        RECT 433.950 554.850 436.050 556.950 ;
        RECT 436.950 556.050 439.050 558.150 ;
        RECT 448.950 557.850 451.050 559.950 ;
        RECT 451.950 559.050 454.050 561.150 ;
        RECT 449.100 556.050 450.900 557.850 ;
        RECT 422.100 553.050 423.900 554.850 ;
        RECT 434.100 553.050 435.900 554.850 ;
        RECT 416.400 551.700 420.150 552.750 ;
        RECT 437.850 552.750 439.050 556.050 ;
        RECT 437.850 551.700 441.600 552.750 ;
        RECT 452.400 551.700 453.600 559.050 ;
        RECT 454.950 557.850 457.050 559.950 ;
        RECT 455.100 556.050 456.900 557.850 ;
        RECT 404.400 550.800 408.000 551.700 ;
        RECT 392.400 543.600 394.200 549.600 ;
        RECT 406.200 543.600 408.000 550.800 ;
        RECT 416.400 549.600 417.600 551.700 ;
        RECT 415.800 543.600 417.600 549.600 ;
        RECT 418.800 548.700 426.600 550.050 ;
        RECT 418.800 543.600 420.600 548.700 ;
        RECT 424.800 543.600 426.600 548.700 ;
        RECT 431.400 548.700 439.200 550.050 ;
        RECT 431.400 543.600 433.200 548.700 ;
        RECT 437.400 543.600 439.200 548.700 ;
        RECT 440.400 549.600 441.600 551.700 ;
        RECT 450.000 550.800 453.600 551.700 ;
        RECT 440.400 543.600 442.200 549.600 ;
        RECT 450.000 543.600 451.800 550.800 ;
        RECT 459.150 549.600 460.050 562.200 ;
        RECT 468.450 561.900 476.850 562.200 ;
        RECT 478.050 562.800 484.050 563.700 ;
        RECT 484.950 562.800 487.050 563.700 ;
        RECT 490.650 563.400 492.450 575.400 ;
        RECT 468.450 561.600 470.250 561.900 ;
        RECT 478.050 558.150 478.950 562.800 ;
        RECT 484.950 561.600 489.150 562.800 ;
        RECT 488.250 559.800 490.050 561.600 ;
        RECT 469.950 557.100 472.050 558.150 ;
        RECT 461.100 555.150 462.900 556.950 ;
        RECT 464.100 556.050 472.050 557.100 ;
        RECT 475.950 556.050 478.950 558.150 ;
        RECT 464.100 555.300 465.900 556.050 ;
        RECT 462.000 554.400 462.900 555.150 ;
        RECT 467.100 554.400 468.900 555.000 ;
        RECT 462.000 553.200 468.900 554.400 ;
        RECT 467.850 552.000 468.900 553.200 ;
        RECT 478.050 552.000 478.950 556.050 ;
        RECT 487.950 555.750 490.050 556.050 ;
        RECT 486.150 553.950 490.050 555.750 ;
        RECT 491.250 553.950 492.450 563.400 ;
        RECT 497.400 569.400 499.200 575.400 ;
        RECT 497.400 562.500 498.600 569.400 ;
        RECT 503.700 563.400 505.500 575.400 ;
        RECT 511.500 563.400 513.300 575.400 ;
        RECT 517.800 569.400 519.600 575.400 ;
        RECT 497.400 561.600 503.100 562.500 ;
        RECT 501.150 560.700 503.100 561.600 ;
        RECT 497.100 558.150 498.900 559.950 ;
        RECT 496.950 556.050 499.050 558.150 ;
        RECT 467.850 551.100 478.950 552.000 ;
        RECT 487.950 551.850 492.450 553.950 ;
        RECT 467.850 550.200 468.900 551.100 ;
        RECT 478.050 550.800 478.950 551.100 ;
        RECT 459.150 543.600 460.950 549.600 ;
        RECT 463.950 547.500 466.050 549.600 ;
        RECT 467.550 548.400 469.350 550.200 ;
        RECT 470.850 549.450 472.650 550.200 ;
        RECT 470.850 548.400 475.800 549.450 ;
        RECT 478.050 549.000 479.850 550.800 ;
        RECT 491.250 549.600 492.450 551.850 ;
        RECT 501.150 552.300 502.050 560.700 ;
        RECT 504.000 558.150 505.200 563.400 ;
        RECT 502.950 556.050 505.200 558.150 ;
        RECT 501.150 551.400 503.100 552.300 ;
        RECT 484.950 548.700 487.050 549.600 ;
        RECT 465.000 546.600 466.050 547.500 ;
        RECT 474.750 546.600 475.800 548.400 ;
        RECT 483.300 547.500 487.050 548.700 ;
        RECT 483.300 546.600 484.350 547.500 ;
        RECT 465.000 545.700 468.750 546.600 ;
        RECT 466.950 543.600 468.750 545.700 ;
        RECT 474.750 543.600 476.550 546.600 ;
        RECT 482.550 543.600 484.350 546.600 ;
        RECT 490.650 543.600 492.450 549.600 ;
        RECT 498.000 550.500 503.100 551.400 ;
        RECT 498.000 546.600 499.200 550.500 ;
        RECT 504.000 549.600 505.200 556.050 ;
        RECT 511.800 558.150 513.000 563.400 ;
        RECT 518.400 562.500 519.600 569.400 ;
        RECT 523.500 563.400 525.300 575.400 ;
        RECT 529.800 569.400 531.600 575.400 ;
        RECT 513.900 561.600 519.600 562.500 ;
        RECT 513.900 560.700 515.850 561.600 ;
        RECT 511.800 556.050 514.050 558.150 ;
        RECT 511.800 549.600 513.000 556.050 ;
        RECT 514.950 552.300 515.850 560.700 ;
        RECT 518.100 558.150 519.900 559.950 ;
        RECT 523.800 558.150 525.000 563.400 ;
        RECT 530.400 562.500 531.600 569.400 ;
        RECT 525.900 561.600 531.600 562.500 ;
        RECT 533.550 563.400 535.350 575.400 ;
        RECT 541.050 569.400 542.850 575.400 ;
        RECT 538.950 567.300 542.850 569.400 ;
        RECT 548.850 568.500 550.650 575.400 ;
        RECT 556.650 569.400 558.450 575.400 ;
        RECT 557.250 568.500 558.450 569.400 ;
        RECT 547.950 567.450 554.550 568.500 ;
        RECT 547.950 566.700 549.750 567.450 ;
        RECT 552.750 566.700 554.550 567.450 ;
        RECT 557.250 566.400 562.050 568.500 ;
        RECT 540.150 564.600 542.850 566.400 ;
        RECT 543.750 565.800 545.550 566.400 ;
        RECT 543.750 564.900 550.050 565.800 ;
        RECT 557.250 565.500 558.450 566.400 ;
        RECT 543.750 564.600 545.550 564.900 ;
        RECT 541.950 563.700 542.850 564.600 ;
        RECT 525.900 560.700 527.850 561.600 ;
        RECT 517.950 556.050 520.050 558.150 ;
        RECT 523.800 556.050 526.050 558.150 ;
        RECT 513.900 551.400 515.850 552.300 ;
        RECT 513.900 550.500 519.000 551.400 ;
        RECT 497.400 543.600 499.200 546.600 ;
        RECT 503.700 543.600 505.500 549.600 ;
        RECT 511.500 543.600 513.300 549.600 ;
        RECT 517.800 546.600 519.000 550.500 ;
        RECT 523.800 549.600 525.000 556.050 ;
        RECT 526.950 552.300 527.850 560.700 ;
        RECT 530.100 558.150 531.900 559.950 ;
        RECT 529.950 556.050 532.050 558.150 ;
        RECT 525.900 551.400 527.850 552.300 ;
        RECT 533.550 553.950 534.750 563.400 ;
        RECT 538.950 562.800 541.050 563.700 ;
        RECT 541.950 562.800 547.950 563.700 ;
        RECT 536.850 561.600 541.050 562.800 ;
        RECT 535.950 559.800 537.750 561.600 ;
        RECT 547.050 558.150 547.950 562.800 ;
        RECT 549.150 562.800 550.050 564.900 ;
        RECT 550.950 564.300 558.450 565.500 ;
        RECT 550.950 563.700 552.750 564.300 ;
        RECT 565.050 563.400 566.850 575.400 ;
        RECT 555.750 562.800 566.850 563.400 ;
        RECT 549.150 562.200 566.850 562.800 ;
        RECT 549.150 561.900 557.550 562.200 ;
        RECT 555.750 561.600 557.550 561.900 ;
        RECT 547.050 556.050 550.050 558.150 ;
        RECT 553.950 557.100 556.050 558.150 ;
        RECT 553.950 556.050 561.900 557.100 ;
        RECT 535.950 555.750 538.050 556.050 ;
        RECT 535.950 553.950 539.850 555.750 ;
        RECT 533.550 551.850 538.050 553.950 ;
        RECT 547.050 552.000 547.950 556.050 ;
        RECT 560.100 555.300 561.900 556.050 ;
        RECT 563.100 555.150 564.900 556.950 ;
        RECT 557.100 554.400 558.900 555.000 ;
        RECT 563.100 554.400 564.000 555.150 ;
        RECT 557.100 553.200 564.000 554.400 ;
        RECT 557.100 552.000 558.150 553.200 ;
        RECT 525.900 550.500 531.000 551.400 ;
        RECT 517.800 543.600 519.600 546.600 ;
        RECT 523.500 543.600 525.300 549.600 ;
        RECT 529.800 546.600 531.000 550.500 ;
        RECT 533.550 549.600 534.750 551.850 ;
        RECT 547.050 551.100 558.150 552.000 ;
        RECT 547.050 550.800 547.950 551.100 ;
        RECT 529.800 543.600 531.600 546.600 ;
        RECT 533.550 543.600 535.350 549.600 ;
        RECT 538.950 548.700 541.050 549.600 ;
        RECT 546.150 549.000 547.950 550.800 ;
        RECT 557.100 550.200 558.150 551.100 ;
        RECT 553.350 549.450 555.150 550.200 ;
        RECT 538.950 547.500 542.700 548.700 ;
        RECT 541.650 546.600 542.700 547.500 ;
        RECT 550.200 548.400 555.150 549.450 ;
        RECT 556.650 548.400 558.450 550.200 ;
        RECT 565.950 549.600 566.850 562.200 ;
        RECT 569.400 569.400 571.200 575.400 ;
        RECT 569.400 562.500 570.600 569.400 ;
        RECT 575.700 563.400 577.500 575.400 ;
        RECT 590.700 563.400 592.500 575.400 ;
        RECT 603.600 563.400 605.400 575.400 ;
        RECT 607.950 567.450 610.050 568.050 ;
        RECT 607.950 566.550 612.450 567.450 ;
        RECT 607.950 565.950 610.050 566.550 ;
        RECT 569.400 561.600 575.100 562.500 ;
        RECT 573.150 560.700 575.100 561.600 ;
        RECT 569.100 558.150 570.900 559.950 ;
        RECT 568.950 556.050 571.050 558.150 ;
        RECT 573.150 552.300 574.050 560.700 ;
        RECT 576.000 558.150 577.200 563.400 ;
        RECT 587.250 561.150 589.050 562.950 ;
        RECT 586.950 559.050 589.050 561.150 ;
        RECT 590.850 558.150 592.050 563.400 ;
        RECT 603.000 562.350 605.400 563.400 ;
        RECT 596.100 558.150 597.900 559.950 ;
        RECT 599.100 558.150 600.900 559.950 ;
        RECT 574.950 556.050 577.200 558.150 ;
        RECT 573.150 551.400 575.100 552.300 ;
        RECT 550.200 546.600 551.250 548.400 ;
        RECT 559.950 547.500 562.050 549.600 ;
        RECT 559.950 546.600 561.000 547.500 ;
        RECT 541.650 543.600 543.450 546.600 ;
        RECT 549.450 543.600 551.250 546.600 ;
        RECT 557.250 545.700 561.000 546.600 ;
        RECT 557.250 543.600 559.050 545.700 ;
        RECT 565.050 543.600 566.850 549.600 ;
        RECT 570.000 550.500 575.100 551.400 ;
        RECT 570.000 546.600 571.200 550.500 ;
        RECT 576.000 549.600 577.200 556.050 ;
        RECT 589.950 556.050 592.050 558.150 ;
        RECT 589.950 552.750 591.150 556.050 ;
        RECT 592.950 554.850 595.050 556.950 ;
        RECT 595.950 556.050 598.050 558.150 ;
        RECT 598.950 556.050 601.050 558.150 ;
        RECT 603.000 555.150 604.050 562.350 ;
        RECT 605.100 558.150 606.900 559.950 ;
        RECT 604.950 556.050 607.050 558.150 ;
        RECT 593.100 553.050 594.900 554.850 ;
        RECT 601.950 553.050 604.050 555.150 ;
        RECT 587.400 551.700 591.150 552.750 ;
        RECT 587.400 549.600 588.600 551.700 ;
        RECT 569.400 543.600 571.200 546.600 ;
        RECT 575.700 543.600 577.500 549.600 ;
        RECT 586.800 543.600 588.600 549.600 ;
        RECT 589.800 548.700 597.600 550.050 ;
        RECT 589.800 543.600 591.600 548.700 ;
        RECT 595.800 543.600 597.600 548.700 ;
        RECT 603.000 546.600 604.050 553.050 ;
        RECT 611.550 550.050 612.450 566.550 ;
        RECT 619.500 563.400 621.300 575.400 ;
        RECT 632.400 569.400 634.200 575.400 ;
        RECT 643.800 569.400 645.600 575.400 ;
        RECT 614.100 558.150 615.900 559.950 ;
        RECT 619.950 558.150 621.150 563.400 ;
        RECT 622.950 561.150 624.750 562.950 ;
        RECT 622.950 559.050 625.050 561.150 ;
        RECT 613.950 556.050 616.050 558.150 ;
        RECT 616.950 554.850 619.050 556.950 ;
        RECT 619.950 556.050 622.050 558.150 ;
        RECT 632.400 556.950 633.600 569.400 ;
        RECT 644.400 556.950 645.600 569.400 ;
        RECT 656.400 569.400 658.200 575.400 ;
        RECT 656.400 561.150 657.600 569.400 ;
        RECT 658.950 564.450 661.050 565.050 ;
        RECT 658.950 563.550 663.450 564.450 ;
        RECT 658.950 562.950 661.050 563.550 ;
        RECT 649.950 556.950 652.050 559.050 ;
        RECT 652.950 557.850 655.050 559.950 ;
        RECT 655.950 559.050 658.050 561.150 ;
        RECT 617.100 553.050 618.900 554.850 ;
        RECT 620.850 552.750 622.050 556.050 ;
        RECT 629.100 555.150 630.900 556.950 ;
        RECT 628.950 553.050 631.050 555.150 ;
        RECT 631.950 554.850 634.050 556.950 ;
        RECT 643.950 554.850 646.050 556.950 ;
        RECT 647.100 555.150 648.900 556.950 ;
        RECT 620.850 551.700 624.600 552.750 ;
        RECT 610.950 547.950 613.050 550.050 ;
        RECT 614.400 548.700 622.200 550.050 ;
        RECT 602.400 543.600 604.200 546.600 ;
        RECT 614.400 543.600 616.200 548.700 ;
        RECT 620.400 543.600 622.200 548.700 ;
        RECT 623.400 549.600 624.600 551.700 ;
        RECT 623.400 543.600 625.200 549.600 ;
        RECT 632.400 546.600 633.600 554.850 ;
        RECT 644.400 546.600 645.600 554.850 ;
        RECT 646.950 553.050 649.050 555.150 ;
        RECT 650.550 552.450 651.450 556.950 ;
        RECT 653.100 556.050 654.900 557.850 ;
        RECT 652.950 552.450 655.050 553.050 ;
        RECT 650.550 551.550 655.050 552.450 ;
        RECT 652.950 550.950 655.050 551.550 ;
        RECT 656.400 551.700 657.600 559.050 ;
        RECT 658.950 557.850 661.050 559.950 ;
        RECT 659.100 556.050 660.900 557.850 ;
        RECT 662.550 552.450 663.450 563.550 ;
        RECT 669.600 563.400 671.400 575.400 ;
        RECT 677.400 564.600 679.200 575.400 ;
        RECT 683.400 574.500 691.200 575.400 ;
        RECT 683.400 564.600 685.200 574.500 ;
        RECT 677.400 563.700 685.200 564.600 ;
        RECT 669.000 562.350 671.400 563.400 ;
        RECT 686.400 562.500 688.200 573.600 ;
        RECT 689.400 563.400 691.200 574.500 ;
        RECT 700.500 563.400 702.300 575.400 ;
        RECT 713.400 569.400 715.200 575.400 ;
        RECT 713.700 569.100 715.200 569.400 ;
        RECT 719.400 569.400 721.200 575.400 ;
        RECT 719.400 569.100 720.300 569.400 ;
        RECT 713.700 568.200 720.300 569.100 ;
        RECT 706.950 565.950 709.050 568.050 ;
        RECT 665.100 558.150 666.900 559.950 ;
        RECT 664.950 556.050 667.050 558.150 ;
        RECT 669.000 555.150 670.050 562.350 ;
        RECT 684.150 561.600 688.200 562.500 ;
        RECT 671.100 558.150 672.900 559.950 ;
        RECT 677.250 558.150 679.050 559.950 ;
        RECT 684.150 558.150 685.050 561.600 ;
        RECT 689.100 558.150 690.900 559.950 ;
        RECT 695.100 558.150 696.900 559.950 ;
        RECT 700.950 558.150 702.150 563.400 ;
        RECT 703.950 561.150 705.750 562.950 ;
        RECT 703.950 559.050 706.050 561.150 ;
        RECT 670.950 556.050 673.050 558.150 ;
        RECT 676.950 556.050 679.050 558.150 ;
        RECT 667.950 553.050 670.050 555.150 ;
        RECT 679.950 554.850 682.050 556.950 ;
        RECT 680.250 553.050 682.050 554.850 ;
        RECT 682.950 556.050 685.050 558.150 ;
        RECT 664.950 552.450 667.050 553.050 ;
        RECT 656.400 550.800 660.000 551.700 ;
        RECT 662.550 551.550 667.050 552.450 ;
        RECT 664.950 550.950 667.050 551.550 ;
        RECT 632.400 543.600 634.200 546.600 ;
        RECT 643.800 543.600 645.600 546.600 ;
        RECT 658.200 543.600 660.000 550.800 ;
        RECT 669.000 546.600 670.050 553.050 ;
        RECT 682.950 549.600 684.000 556.050 ;
        RECT 685.950 554.850 688.050 556.950 ;
        RECT 688.950 556.050 691.050 558.150 ;
        RECT 694.950 556.050 697.050 558.150 ;
        RECT 697.950 554.850 700.050 556.950 ;
        RECT 700.950 556.050 703.050 558.150 ;
        RECT 685.950 553.050 687.750 554.850 ;
        RECT 698.100 553.050 699.900 554.850 ;
        RECT 701.850 552.750 703.050 556.050 ;
        RECT 703.950 555.450 706.050 556.050 ;
        RECT 707.550 555.450 708.450 565.950 ;
        RECT 713.100 564.150 714.900 565.950 ;
        RECT 710.100 561.150 711.900 562.950 ;
        RECT 712.950 562.050 715.050 564.150 ;
        RECT 716.250 561.150 718.050 562.950 ;
        RECT 709.950 559.050 712.050 561.150 ;
        RECT 715.950 559.050 718.050 561.150 ;
        RECT 719.400 559.950 720.300 568.200 ;
        RECT 730.800 563.400 732.600 575.400 ;
        RECT 743.400 569.400 745.200 575.400 ;
        RECT 718.950 557.850 721.050 559.950 ;
        RECT 703.950 554.550 708.450 555.450 ;
        RECT 703.950 553.950 706.050 554.550 ;
        RECT 719.400 553.650 720.300 557.850 ;
        RECT 730.950 556.950 732.300 563.400 ;
        RECT 740.100 558.150 741.900 559.950 ;
        RECT 727.950 554.850 732.300 556.950 ;
        RECT 733.950 554.850 736.050 556.950 ;
        RECT 739.950 556.050 742.050 558.150 ;
        RECT 701.850 551.700 705.600 552.750 ;
        RECT 668.400 543.600 670.200 546.600 ;
        RECT 682.200 543.600 684.000 549.600 ;
        RECT 695.400 548.700 703.200 550.050 ;
        RECT 695.400 543.600 697.200 548.700 ;
        RECT 701.400 543.600 703.200 548.700 ;
        RECT 704.400 549.600 705.600 551.700 ;
        RECT 716.100 552.000 720.300 553.650 ;
        RECT 704.400 543.600 706.200 549.600 ;
        RECT 716.100 543.600 717.900 552.000 ;
        RECT 730.950 549.600 732.300 554.850 ;
        RECT 734.100 553.050 735.900 554.850 ;
        RECT 743.550 552.300 744.600 569.400 ;
        RECT 750.000 563.400 751.800 575.400 ;
        RECT 745.950 557.850 748.050 559.950 ;
        RECT 750.000 558.150 751.050 563.400 ;
        RECT 746.100 556.050 747.900 557.850 ;
        RECT 748.950 556.050 751.050 558.150 ;
        RECT 740.400 551.100 747.900 552.300 ;
        RECT 730.800 543.600 732.600 549.600 ;
        RECT 740.400 543.600 742.200 551.100 ;
        RECT 746.100 550.500 747.900 551.100 ;
        RECT 750.000 549.600 751.050 556.050 ;
        RECT 747.900 548.100 751.050 549.600 ;
        RECT 747.900 543.600 749.700 548.100 ;
        RECT 7.500 533.400 9.300 539.400 ;
        RECT 13.800 536.400 15.600 539.400 ;
        RECT 7.800 526.950 9.000 533.400 ;
        RECT 13.800 532.500 15.000 536.400 ;
        RECT 27.000 535.050 28.800 539.400 ;
        RECT 40.800 536.400 42.600 539.400 ;
        RECT 9.900 531.600 15.000 532.500 ;
        RECT 23.400 533.400 28.800 535.050 ;
        RECT 9.900 530.700 11.850 531.600 ;
        RECT 7.800 524.850 10.050 526.950 ;
        RECT 7.800 519.600 9.000 524.850 ;
        RECT 10.950 522.300 11.850 530.700 ;
        RECT 23.400 526.950 24.300 533.400 ;
        RECT 26.100 528.150 27.900 529.950 ;
        RECT 13.950 524.850 16.050 526.950 ;
        RECT 22.950 524.850 25.050 526.950 ;
        RECT 25.950 526.050 28.050 528.150 ;
        RECT 28.950 527.850 31.050 529.950 ;
        RECT 32.100 528.150 33.900 529.950 ;
        RECT 41.400 528.150 42.600 536.400 ;
        RECT 49.800 533.400 51.600 539.400 ;
        RECT 50.400 531.300 51.600 533.400 ;
        RECT 52.800 534.300 54.600 539.400 ;
        RECT 58.800 534.300 60.600 539.400 ;
        RECT 52.800 532.950 60.600 534.300 ;
        RECT 66.000 532.200 67.800 539.400 ;
        RECT 76.800 533.400 78.600 539.400 ;
        RECT 66.000 531.300 69.600 532.200 ;
        RECT 50.400 530.250 54.150 531.300 ;
        RECT 29.100 526.050 30.900 527.850 ;
        RECT 31.950 526.050 34.050 528.150 ;
        RECT 40.950 526.050 43.050 528.150 ;
        RECT 43.950 527.850 46.050 529.950 ;
        RECT 44.100 526.050 45.900 527.850 ;
        RECT 52.950 526.950 54.150 530.250 ;
        RECT 56.100 528.150 57.900 529.950 ;
        RECT 14.100 523.050 15.900 524.850 ;
        RECT 9.900 521.400 11.850 522.300 ;
        RECT 9.900 520.500 15.600 521.400 ;
        RECT 7.500 507.600 9.300 519.600 ;
        RECT 14.400 513.600 15.600 520.500 ;
        RECT 23.400 519.600 24.300 524.850 ;
        RECT 13.800 507.600 15.600 513.600 ;
        RECT 22.800 507.600 24.600 519.600 ;
        RECT 25.800 518.700 33.600 519.600 ;
        RECT 25.800 507.600 27.600 518.700 ;
        RECT 31.800 507.600 33.600 518.700 ;
        RECT 41.400 513.600 42.600 526.050 ;
        RECT 52.950 524.850 55.050 526.950 ;
        RECT 55.950 526.050 58.050 528.150 ;
        RECT 61.950 526.950 64.050 529.050 ;
        RECT 58.950 524.850 61.050 526.950 ;
        RECT 49.950 521.850 52.050 523.950 ;
        RECT 50.250 520.050 52.050 521.850 ;
        RECT 53.850 519.600 55.050 524.850 ;
        RECT 59.100 523.050 60.900 524.850 ;
        RECT 62.550 520.050 63.450 526.950 ;
        RECT 65.100 525.150 66.900 526.950 ;
        RECT 64.950 523.050 67.050 525.150 ;
        RECT 68.400 523.950 69.600 531.300 ;
        RECT 77.400 531.300 78.600 533.400 ;
        RECT 79.800 534.300 81.600 539.400 ;
        RECT 85.800 534.300 87.600 539.400 ;
        RECT 79.800 532.950 87.600 534.300 ;
        RECT 91.800 533.400 93.600 539.400 ;
        RECT 92.400 531.300 93.600 533.400 ;
        RECT 94.800 534.300 96.600 539.400 ;
        RECT 100.800 534.300 102.600 539.400 ;
        RECT 94.800 532.950 102.600 534.300 ;
        RECT 109.200 532.200 111.000 539.400 ;
        RECT 121.200 535.050 123.000 539.400 ;
        RECT 133.800 536.400 135.600 539.400 ;
        RECT 121.200 533.400 126.600 535.050 ;
        RECT 107.400 531.300 111.000 532.200 ;
        RECT 77.400 530.250 81.150 531.300 ;
        RECT 92.400 530.250 96.150 531.300 ;
        RECT 79.950 526.950 81.150 530.250 ;
        RECT 83.100 528.150 84.900 529.950 ;
        RECT 71.100 525.150 72.900 526.950 ;
        RECT 67.950 521.850 70.050 523.950 ;
        RECT 70.950 523.050 73.050 525.150 ;
        RECT 79.950 524.850 82.050 526.950 ;
        RECT 82.950 526.050 85.050 528.150 ;
        RECT 94.950 526.950 96.150 530.250 ;
        RECT 98.100 528.150 99.900 529.950 ;
        RECT 85.950 524.850 88.050 526.950 ;
        RECT 94.950 524.850 97.050 526.950 ;
        RECT 97.950 526.050 100.050 528.150 ;
        RECT 100.950 524.850 103.050 526.950 ;
        RECT 104.100 525.150 105.900 526.950 ;
        RECT 76.950 521.850 79.050 523.950 ;
        RECT 40.800 507.600 42.600 513.600 ;
        RECT 53.700 507.600 55.500 519.600 ;
        RECT 61.950 517.950 64.050 520.050 ;
        RECT 68.400 513.600 69.600 521.850 ;
        RECT 77.250 520.050 79.050 521.850 ;
        RECT 80.850 519.600 82.050 524.850 ;
        RECT 86.100 523.050 87.900 524.850 ;
        RECT 91.950 521.850 94.050 523.950 ;
        RECT 92.250 520.050 94.050 521.850 ;
        RECT 95.850 519.600 97.050 524.850 ;
        RECT 101.100 523.050 102.900 524.850 ;
        RECT 103.950 523.050 106.050 525.150 ;
        RECT 107.400 523.950 108.600 531.300 ;
        RECT 116.100 528.150 117.900 529.950 ;
        RECT 110.100 525.150 111.900 526.950 ;
        RECT 115.950 526.050 118.050 528.150 ;
        RECT 118.950 527.850 121.050 529.950 ;
        RECT 122.100 528.150 123.900 529.950 ;
        RECT 119.100 526.050 120.900 527.850 ;
        RECT 121.950 526.050 124.050 528.150 ;
        RECT 125.700 526.950 126.600 533.400 ;
        RECT 127.950 529.950 130.050 532.050 ;
        RECT 106.950 521.850 109.050 523.950 ;
        RECT 109.950 523.050 112.050 525.150 ;
        RECT 124.950 524.850 127.050 526.950 ;
        RECT 67.800 507.600 69.600 513.600 ;
        RECT 80.700 507.600 82.500 519.600 ;
        RECT 95.700 507.600 97.500 519.600 ;
        RECT 107.400 513.600 108.600 521.850 ;
        RECT 125.700 519.600 126.600 524.850 ;
        RECT 128.550 522.450 129.450 529.950 ;
        RECT 134.400 528.150 135.600 536.400 ;
        RECT 147.000 535.050 148.800 539.400 ;
        RECT 143.400 533.400 148.800 535.050 ;
        RECT 158.400 536.400 160.200 539.400 ;
        RECT 133.950 526.050 136.050 528.150 ;
        RECT 136.950 527.850 139.050 529.950 ;
        RECT 137.100 526.050 138.900 527.850 ;
        RECT 143.400 526.950 144.300 533.400 ;
        RECT 146.100 528.150 147.900 529.950 ;
        RECT 130.950 522.450 133.050 523.050 ;
        RECT 128.550 521.550 133.050 522.450 ;
        RECT 130.950 520.950 133.050 521.550 ;
        RECT 116.400 518.700 124.200 519.600 ;
        RECT 107.400 507.600 109.200 513.600 ;
        RECT 116.400 507.600 118.200 518.700 ;
        RECT 122.400 507.600 124.200 518.700 ;
        RECT 125.400 507.600 127.200 519.600 ;
        RECT 134.400 513.600 135.600 526.050 ;
        RECT 142.950 524.850 145.050 526.950 ;
        RECT 145.950 526.050 148.050 528.150 ;
        RECT 148.950 527.850 151.050 529.950 ;
        RECT 152.100 528.150 153.900 529.950 ;
        RECT 149.100 526.050 150.900 527.850 ;
        RECT 151.950 526.050 154.050 528.150 ;
        RECT 154.950 527.850 157.050 529.950 ;
        RECT 158.400 528.150 159.600 536.400 ;
        RECT 169.200 535.050 171.000 539.400 ;
        RECT 169.200 533.400 174.600 535.050 ;
        RECT 164.100 528.150 165.900 529.950 ;
        RECT 155.100 526.050 156.900 527.850 ;
        RECT 157.950 526.050 160.050 528.150 ;
        RECT 163.950 526.050 166.050 528.150 ;
        RECT 166.950 527.850 169.050 529.950 ;
        RECT 170.100 528.150 171.900 529.950 ;
        RECT 167.100 526.050 168.900 527.850 ;
        RECT 169.950 526.050 172.050 528.150 ;
        RECT 173.700 526.950 174.600 533.400 ;
        RECT 182.400 534.300 184.200 539.400 ;
        RECT 188.400 534.300 190.200 539.400 ;
        RECT 182.400 532.950 190.200 534.300 ;
        RECT 191.400 533.400 193.200 539.400 ;
        RECT 203.400 536.400 205.200 539.400 ;
        RECT 215.400 536.400 217.200 539.400 ;
        RECT 229.800 536.400 231.600 539.400 ;
        RECT 191.400 531.300 192.600 533.400 ;
        RECT 188.850 530.250 192.600 531.300 ;
        RECT 185.100 528.150 186.900 529.950 ;
        RECT 143.400 519.600 144.300 524.850 ;
        RECT 133.800 507.600 135.600 513.600 ;
        RECT 142.800 507.600 144.600 519.600 ;
        RECT 145.800 518.700 153.600 519.600 ;
        RECT 145.800 507.600 147.600 518.700 ;
        RECT 151.800 507.600 153.600 518.700 ;
        RECT 158.400 513.600 159.600 526.050 ;
        RECT 172.950 524.850 175.050 526.950 ;
        RECT 181.950 524.850 184.050 526.950 ;
        RECT 184.950 526.050 187.050 528.150 ;
        RECT 188.850 526.950 190.050 530.250 ;
        RECT 204.000 529.950 205.050 536.400 ;
        RECT 216.000 529.950 217.050 536.400 ;
        RECT 202.950 527.850 205.050 529.950 ;
        RECT 214.950 527.850 217.050 529.950 ;
        RECT 187.950 524.850 190.050 526.950 ;
        RECT 199.950 524.850 202.050 526.950 ;
        RECT 173.700 519.600 174.600 524.850 ;
        RECT 182.100 523.050 183.900 524.850 ;
        RECT 187.950 519.600 189.150 524.850 ;
        RECT 190.950 521.850 193.050 523.950 ;
        RECT 200.100 523.050 201.900 524.850 ;
        RECT 190.950 520.050 192.750 521.850 ;
        RECT 204.000 520.650 205.050 527.850 ;
        RECT 205.950 524.850 208.050 526.950 ;
        RECT 211.950 524.850 214.050 526.950 ;
        RECT 206.100 523.050 207.900 524.850 ;
        RECT 212.100 523.050 213.900 524.850 ;
        RECT 216.000 520.650 217.050 527.850 ;
        RECT 229.950 529.950 231.000 536.400 ;
        RECT 241.200 533.400 243.000 539.400 ;
        RECT 229.950 527.850 232.050 529.950 ;
        RECT 239.250 528.150 241.050 529.950 ;
        RECT 217.950 524.850 220.050 526.950 ;
        RECT 226.950 524.850 229.050 526.950 ;
        RECT 218.100 523.050 219.900 524.850 ;
        RECT 227.100 523.050 228.900 524.850 ;
        RECT 229.950 520.650 231.000 527.850 ;
        RECT 232.950 524.850 235.050 526.950 ;
        RECT 235.950 524.850 238.050 526.950 ;
        RECT 238.950 526.050 241.050 528.150 ;
        RECT 241.950 526.950 243.000 533.400 ;
        RECT 259.200 532.200 261.000 539.400 ;
        RECT 270.300 534.900 272.100 539.400 ;
        RECT 257.400 531.300 261.000 532.200 ;
        RECT 268.950 533.400 272.100 534.900 ;
        RECT 244.950 528.150 246.750 529.950 ;
        RECT 241.950 524.850 244.050 526.950 ;
        RECT 244.950 526.050 247.050 528.150 ;
        RECT 247.950 524.850 250.050 526.950 ;
        RECT 254.100 525.150 255.900 526.950 ;
        RECT 233.100 523.050 234.900 524.850 ;
        RECT 236.250 523.050 238.050 524.850 ;
        RECT 204.000 519.600 206.400 520.650 ;
        RECT 216.000 519.600 218.400 520.650 ;
        RECT 164.400 518.700 172.200 519.600 ;
        RECT 158.400 507.600 160.200 513.600 ;
        RECT 164.400 507.600 166.200 518.700 ;
        RECT 170.400 507.600 172.200 518.700 ;
        RECT 173.400 507.600 175.200 519.600 ;
        RECT 187.500 507.600 189.300 519.600 ;
        RECT 204.600 507.600 206.400 519.600 ;
        RECT 216.600 507.600 218.400 519.600 ;
        RECT 228.600 519.600 231.000 520.650 ;
        RECT 243.150 521.400 244.050 524.850 ;
        RECT 248.100 523.050 249.900 524.850 ;
        RECT 253.950 523.050 256.050 525.150 ;
        RECT 257.400 523.950 258.600 531.300 ;
        RECT 268.950 526.950 270.000 533.400 ;
        RECT 272.100 531.900 273.900 532.500 ;
        RECT 277.800 531.900 279.600 539.400 ;
        RECT 283.800 533.400 285.600 539.400 ;
        RECT 272.100 530.700 279.600 531.900 ;
        RECT 284.400 531.300 285.600 533.400 ;
        RECT 286.800 534.300 288.600 539.400 ;
        RECT 292.800 534.300 294.600 539.400 ;
        RECT 286.800 532.950 294.600 534.300 ;
        RECT 301.200 533.400 303.000 539.400 ;
        RECT 260.100 525.150 261.900 526.950 ;
        RECT 256.950 521.850 259.050 523.950 ;
        RECT 259.950 523.050 262.050 525.150 ;
        RECT 268.950 524.850 271.050 526.950 ;
        RECT 272.100 525.150 273.900 526.950 ;
        RECT 243.150 520.500 247.200 521.400 ;
        RECT 228.600 507.600 230.400 519.600 ;
        RECT 236.400 518.400 244.200 519.300 ;
        RECT 236.400 507.600 238.200 518.400 ;
        RECT 242.400 508.500 244.200 518.400 ;
        RECT 245.400 509.400 247.200 520.500 ;
        RECT 248.400 508.500 250.200 519.600 ;
        RECT 242.400 507.600 250.200 508.500 ;
        RECT 257.400 513.600 258.600 521.850 ;
        RECT 268.950 519.600 270.000 524.850 ;
        RECT 271.950 523.050 274.050 525.150 ;
        RECT 257.400 507.600 259.200 513.600 ;
        RECT 268.200 507.600 270.000 519.600 ;
        RECT 275.400 513.600 276.450 530.700 ;
        RECT 284.400 530.250 288.150 531.300 ;
        RECT 286.950 526.950 288.150 530.250 ;
        RECT 290.100 528.150 291.900 529.950 ;
        RECT 299.250 528.150 301.050 529.950 ;
        RECT 277.950 524.850 280.050 526.950 ;
        RECT 286.950 524.850 289.050 526.950 ;
        RECT 289.950 526.050 292.050 528.150 ;
        RECT 292.950 524.850 295.050 526.950 ;
        RECT 295.950 524.850 298.050 526.950 ;
        RECT 298.950 526.050 301.050 528.150 ;
        RECT 301.950 526.950 303.000 533.400 ;
        RECT 322.200 532.200 324.000 539.400 ;
        RECT 325.950 532.950 328.050 535.050 ;
        RECT 320.400 531.300 324.000 532.200 ;
        RECT 304.950 528.150 306.750 529.950 ;
        RECT 301.950 524.850 304.050 526.950 ;
        RECT 304.950 526.050 307.050 528.150 ;
        RECT 307.950 524.850 310.050 526.950 ;
        RECT 317.100 525.150 318.900 526.950 ;
        RECT 278.100 523.050 279.900 524.850 ;
        RECT 283.950 521.850 286.050 523.950 ;
        RECT 284.250 520.050 286.050 521.850 ;
        RECT 287.850 519.600 289.050 524.850 ;
        RECT 293.100 523.050 294.900 524.850 ;
        RECT 296.250 523.050 298.050 524.850 ;
        RECT 303.150 521.400 304.050 524.850 ;
        RECT 308.100 523.050 309.900 524.850 ;
        RECT 316.950 523.050 319.050 525.150 ;
        RECT 320.400 523.950 321.600 531.300 ;
        RECT 323.100 525.150 324.900 526.950 ;
        RECT 319.950 521.850 322.050 523.950 ;
        RECT 322.950 523.050 325.050 525.150 ;
        RECT 303.150 520.500 307.200 521.400 ;
        RECT 274.800 507.600 276.600 513.600 ;
        RECT 287.700 507.600 289.500 519.600 ;
        RECT 296.400 518.400 304.200 519.300 ;
        RECT 296.400 507.600 298.200 518.400 ;
        RECT 302.400 508.500 304.200 518.400 ;
        RECT 305.400 509.400 307.200 520.500 ;
        RECT 308.400 508.500 310.200 519.600 ;
        RECT 302.400 507.600 310.200 508.500 ;
        RECT 320.400 513.600 321.600 521.850 ;
        RECT 326.550 519.450 327.450 532.950 ;
        RECT 329.400 531.900 331.200 539.400 ;
        RECT 336.900 534.900 338.700 539.400 ;
        RECT 336.900 533.400 340.050 534.900 ;
        RECT 335.100 531.900 336.900 532.500 ;
        RECT 329.400 530.700 336.900 531.900 ;
        RECT 328.950 524.850 331.050 526.950 ;
        RECT 329.100 523.050 330.900 524.850 ;
        RECT 328.950 519.450 331.050 520.050 ;
        RECT 326.550 518.550 331.050 519.450 ;
        RECT 328.950 517.950 331.050 518.550 ;
        RECT 332.550 513.600 333.600 530.700 ;
        RECT 339.000 526.950 340.050 533.400 ;
        RECT 344.400 534.300 346.200 539.400 ;
        RECT 350.400 534.300 352.200 539.400 ;
        RECT 344.400 532.950 352.200 534.300 ;
        RECT 353.400 533.400 355.200 539.400 ;
        RECT 365.400 536.400 367.200 539.400 ;
        RECT 353.400 531.300 354.600 533.400 ;
        RECT 350.850 530.250 354.600 531.300 ;
        RECT 347.100 528.150 348.900 529.950 ;
        RECT 335.100 525.150 336.900 526.950 ;
        RECT 334.950 523.050 337.050 525.150 ;
        RECT 337.950 524.850 340.050 526.950 ;
        RECT 343.950 524.850 346.050 526.950 ;
        RECT 346.950 526.050 349.050 528.150 ;
        RECT 350.850 526.950 352.050 530.250 ;
        RECT 366.000 529.950 367.050 536.400 ;
        RECT 376.800 533.400 378.600 539.400 ;
        RECT 377.400 531.300 378.600 533.400 ;
        RECT 379.800 534.300 381.600 539.400 ;
        RECT 385.800 534.300 387.600 539.400 ;
        RECT 379.800 532.950 387.600 534.300 ;
        RECT 394.200 532.200 396.000 539.400 ;
        RECT 406.800 533.400 408.600 539.400 ;
        RECT 392.400 531.300 396.000 532.200 ;
        RECT 407.400 531.300 408.600 533.400 ;
        RECT 409.800 534.300 411.600 539.400 ;
        RECT 415.800 534.300 417.600 539.400 ;
        RECT 409.800 532.950 417.600 534.300 ;
        RECT 422.400 536.400 424.200 539.400 ;
        RECT 377.400 530.250 381.150 531.300 ;
        RECT 364.950 527.850 367.050 529.950 ;
        RECT 349.950 524.850 352.050 526.950 ;
        RECT 361.950 524.850 364.050 526.950 ;
        RECT 339.000 519.600 340.050 524.850 ;
        RECT 344.100 523.050 345.900 524.850 ;
        RECT 349.950 519.600 351.150 524.850 ;
        RECT 352.950 521.850 355.050 523.950 ;
        RECT 362.100 523.050 363.900 524.850 ;
        RECT 352.950 520.050 354.750 521.850 ;
        RECT 366.000 520.650 367.050 527.850 ;
        RECT 379.950 526.950 381.150 530.250 ;
        RECT 383.100 528.150 384.900 529.950 ;
        RECT 367.950 524.850 370.050 526.950 ;
        RECT 379.950 524.850 382.050 526.950 ;
        RECT 382.950 526.050 385.050 528.150 ;
        RECT 385.950 524.850 388.050 526.950 ;
        RECT 389.100 525.150 390.900 526.950 ;
        RECT 368.100 523.050 369.900 524.850 ;
        RECT 376.950 521.850 379.050 523.950 ;
        RECT 366.000 519.600 368.400 520.650 ;
        RECT 377.250 520.050 379.050 521.850 ;
        RECT 380.850 519.600 382.050 524.850 ;
        RECT 386.100 523.050 387.900 524.850 ;
        RECT 388.950 523.050 391.050 525.150 ;
        RECT 392.400 523.950 393.600 531.300 ;
        RECT 407.400 530.250 411.150 531.300 ;
        RECT 409.950 526.950 411.150 530.250 ;
        RECT 413.100 528.150 414.900 529.950 ;
        RECT 395.100 525.150 396.900 526.950 ;
        RECT 391.950 521.850 394.050 523.950 ;
        RECT 394.950 523.050 397.050 525.150 ;
        RECT 409.950 524.850 412.050 526.950 ;
        RECT 412.950 526.050 415.050 528.150 ;
        RECT 418.950 527.850 421.050 529.950 ;
        RECT 422.400 528.150 423.600 536.400 ;
        RECT 433.200 532.200 435.000 539.400 ;
        RECT 447.000 535.050 448.800 539.400 ;
        RECT 427.950 531.450 430.050 532.050 ;
        RECT 425.550 530.550 430.050 531.450 ;
        RECT 415.950 524.850 418.050 526.950 ;
        RECT 419.100 526.050 420.900 527.850 ;
        RECT 421.950 526.050 424.050 528.150 ;
        RECT 406.950 521.850 409.050 523.950 ;
        RECT 320.400 507.600 322.200 513.600 ;
        RECT 332.400 507.600 334.200 513.600 ;
        RECT 339.000 507.600 340.800 519.600 ;
        RECT 349.500 507.600 351.300 519.600 ;
        RECT 366.600 507.600 368.400 519.600 ;
        RECT 380.700 507.600 382.500 519.600 ;
        RECT 392.400 513.600 393.600 521.850 ;
        RECT 407.250 520.050 409.050 521.850 ;
        RECT 410.850 519.600 412.050 524.850 ;
        RECT 416.100 523.050 417.900 524.850 ;
        RECT 392.400 507.600 394.200 513.600 ;
        RECT 410.700 507.600 412.500 519.600 ;
        RECT 422.400 513.600 423.600 526.050 ;
        RECT 425.550 520.050 426.450 530.550 ;
        RECT 427.950 529.950 430.050 530.550 ;
        RECT 431.400 531.300 435.000 532.200 ;
        RECT 443.400 533.400 448.800 535.050 ;
        RECT 455.400 534.300 457.200 539.400 ;
        RECT 461.400 534.300 463.200 539.400 ;
        RECT 428.100 525.150 429.900 526.950 ;
        RECT 427.950 523.050 430.050 525.150 ;
        RECT 431.400 523.950 432.600 531.300 ;
        RECT 443.400 526.950 444.300 533.400 ;
        RECT 455.400 532.950 463.200 534.300 ;
        RECT 464.400 533.400 466.200 539.400 ;
        RECT 464.400 531.300 465.600 533.400 ;
        RECT 475.200 532.200 477.000 539.400 ;
        RECT 461.850 530.250 465.600 531.300 ;
        RECT 473.400 531.300 477.000 532.200 ;
        RECT 482.550 533.400 484.350 539.400 ;
        RECT 490.650 536.400 492.450 539.400 ;
        RECT 498.450 536.400 500.250 539.400 ;
        RECT 506.250 537.300 508.050 539.400 ;
        RECT 506.250 536.400 510.000 537.300 ;
        RECT 490.650 535.500 491.700 536.400 ;
        RECT 487.950 534.300 491.700 535.500 ;
        RECT 499.200 534.600 500.250 536.400 ;
        RECT 508.950 535.500 510.000 536.400 ;
        RECT 487.950 533.400 490.050 534.300 ;
        RECT 446.100 528.150 447.900 529.950 ;
        RECT 434.100 525.150 435.900 526.950 ;
        RECT 430.950 521.850 433.050 523.950 ;
        RECT 433.950 523.050 436.050 525.150 ;
        RECT 442.950 524.850 445.050 526.950 ;
        RECT 445.950 526.050 448.050 528.150 ;
        RECT 448.950 527.850 451.050 529.950 ;
        RECT 452.100 528.150 453.900 529.950 ;
        RECT 458.100 528.150 459.900 529.950 ;
        RECT 449.100 526.050 450.900 527.850 ;
        RECT 451.950 526.050 454.050 528.150 ;
        RECT 454.950 524.850 457.050 526.950 ;
        RECT 457.950 526.050 460.050 528.150 ;
        RECT 461.850 526.950 463.050 530.250 ;
        RECT 460.950 524.850 463.050 526.950 ;
        RECT 470.100 525.150 471.900 526.950 ;
        RECT 424.950 517.950 427.050 520.050 ;
        RECT 431.400 513.600 432.600 521.850 ;
        RECT 443.400 519.600 444.300 524.850 ;
        RECT 455.100 523.050 456.900 524.850 ;
        RECT 460.950 519.600 462.150 524.850 ;
        RECT 463.950 521.850 466.050 523.950 ;
        RECT 469.950 523.050 472.050 525.150 ;
        RECT 473.400 523.950 474.600 531.300 ;
        RECT 482.550 531.150 483.750 533.400 ;
        RECT 495.150 532.200 496.950 534.000 ;
        RECT 499.200 533.550 504.150 534.600 ;
        RECT 502.350 532.800 504.150 533.550 ;
        RECT 505.650 532.800 507.450 534.600 ;
        RECT 508.950 533.400 511.050 535.500 ;
        RECT 514.050 533.400 515.850 539.400 ;
        RECT 496.050 531.900 496.950 532.200 ;
        RECT 506.100 531.900 507.150 532.800 ;
        RECT 482.550 529.050 487.050 531.150 ;
        RECT 496.050 531.000 507.150 531.900 ;
        RECT 476.100 525.150 477.900 526.950 ;
        RECT 472.950 521.850 475.050 523.950 ;
        RECT 475.950 523.050 478.050 525.150 ;
        RECT 463.950 520.050 465.750 521.850 ;
        RECT 422.400 507.600 424.200 513.600 ;
        RECT 431.400 507.600 433.200 513.600 ;
        RECT 442.800 507.600 444.600 519.600 ;
        RECT 445.800 518.700 453.600 519.600 ;
        RECT 445.800 507.600 447.600 518.700 ;
        RECT 451.800 507.600 453.600 518.700 ;
        RECT 460.500 507.600 462.300 519.600 ;
        RECT 473.400 513.600 474.600 521.850 ;
        RECT 482.550 519.600 483.750 529.050 ;
        RECT 484.950 527.250 488.850 529.050 ;
        RECT 484.950 526.950 487.050 527.250 ;
        RECT 496.050 526.950 496.950 531.000 ;
        RECT 506.100 529.800 507.150 531.000 ;
        RECT 506.100 528.600 513.000 529.800 ;
        RECT 506.100 528.000 507.900 528.600 ;
        RECT 512.100 527.850 513.000 528.600 ;
        RECT 509.100 526.950 510.900 527.700 ;
        RECT 496.050 524.850 499.050 526.950 ;
        RECT 502.950 525.900 510.900 526.950 ;
        RECT 512.100 526.050 513.900 527.850 ;
        RECT 502.950 524.850 505.050 525.900 ;
        RECT 484.950 521.400 486.750 523.200 ;
        RECT 485.850 520.200 490.050 521.400 ;
        RECT 496.050 520.200 496.950 524.850 ;
        RECT 504.750 521.100 506.550 521.400 ;
        RECT 473.400 507.600 475.200 513.600 ;
        RECT 482.550 507.600 484.350 519.600 ;
        RECT 487.950 519.300 490.050 520.200 ;
        RECT 490.950 519.300 496.950 520.200 ;
        RECT 498.150 520.800 506.550 521.100 ;
        RECT 514.950 520.800 515.850 533.400 ;
        RECT 518.400 534.300 520.200 539.400 ;
        RECT 524.400 534.300 526.200 539.400 ;
        RECT 518.400 532.950 526.200 534.300 ;
        RECT 527.400 533.400 529.200 539.400 ;
        RECT 527.400 531.300 528.600 533.400 ;
        RECT 538.200 532.200 540.000 539.400 ;
        RECT 545.400 536.400 547.200 539.400 ;
        RECT 532.950 531.450 535.050 532.050 ;
        RECT 524.850 530.250 528.600 531.300 ;
        RECT 530.550 530.550 535.050 531.450 ;
        RECT 521.100 528.150 522.900 529.950 ;
        RECT 517.950 524.850 520.050 526.950 ;
        RECT 520.950 526.050 523.050 528.150 ;
        RECT 524.850 526.950 526.050 530.250 ;
        RECT 523.950 524.850 526.050 526.950 ;
        RECT 518.100 523.050 519.900 524.850 ;
        RECT 498.150 520.200 515.850 520.800 ;
        RECT 490.950 518.400 491.850 519.300 ;
        RECT 489.150 516.600 491.850 518.400 ;
        RECT 492.750 518.100 494.550 518.400 ;
        RECT 498.150 518.100 499.050 520.200 ;
        RECT 504.750 519.600 515.850 520.200 ;
        RECT 523.950 519.600 525.150 524.850 ;
        RECT 526.950 521.850 529.050 523.950 ;
        RECT 526.950 520.050 528.750 521.850 ;
        RECT 492.750 517.200 499.050 518.100 ;
        RECT 499.950 518.700 501.750 519.300 ;
        RECT 499.950 517.500 507.450 518.700 ;
        RECT 492.750 516.600 494.550 517.200 ;
        RECT 506.250 516.600 507.450 517.500 ;
        RECT 487.950 513.600 491.850 515.700 ;
        RECT 496.950 515.550 498.750 516.300 ;
        RECT 501.750 515.550 503.550 516.300 ;
        RECT 496.950 514.500 503.550 515.550 ;
        RECT 506.250 514.500 511.050 516.600 ;
        RECT 490.050 507.600 491.850 513.600 ;
        RECT 497.850 507.600 499.650 514.500 ;
        RECT 506.250 513.600 507.450 514.500 ;
        RECT 505.650 507.600 507.450 513.600 ;
        RECT 514.050 507.600 515.850 519.600 ;
        RECT 523.500 507.600 525.300 519.600 ;
        RECT 526.950 516.450 529.050 517.050 ;
        RECT 530.550 516.450 531.450 530.550 ;
        RECT 532.950 529.950 535.050 530.550 ;
        RECT 536.400 531.300 540.000 532.200 ;
        RECT 546.000 532.500 547.200 536.400 ;
        RECT 551.700 533.400 553.500 539.400 ;
        RECT 557.400 534.300 559.200 539.400 ;
        RECT 563.400 534.300 565.200 539.400 ;
        RECT 546.000 531.600 551.100 532.500 ;
        RECT 533.100 525.150 534.900 526.950 ;
        RECT 532.950 523.050 535.050 525.150 ;
        RECT 536.400 523.950 537.600 531.300 ;
        RECT 549.150 530.700 551.100 531.600 ;
        RECT 539.100 525.150 540.900 526.950 ;
        RECT 535.950 521.850 538.050 523.950 ;
        RECT 538.950 523.050 541.050 525.150 ;
        RECT 544.950 524.850 547.050 526.950 ;
        RECT 545.100 523.050 546.900 524.850 ;
        RECT 549.150 522.300 550.050 530.700 ;
        RECT 552.000 526.950 553.200 533.400 ;
        RECT 557.400 532.950 565.200 534.300 ;
        RECT 566.400 533.400 568.200 539.400 ;
        RECT 572.550 533.400 574.350 539.400 ;
        RECT 580.650 536.400 582.450 539.400 ;
        RECT 588.450 536.400 590.250 539.400 ;
        RECT 596.250 537.300 598.050 539.400 ;
        RECT 596.250 536.400 600.000 537.300 ;
        RECT 580.650 535.500 581.700 536.400 ;
        RECT 577.950 534.300 581.700 535.500 ;
        RECT 589.200 534.600 590.250 536.400 ;
        RECT 598.950 535.500 600.000 536.400 ;
        RECT 577.950 533.400 580.050 534.300 ;
        RECT 566.400 531.300 567.600 533.400 ;
        RECT 563.850 530.250 567.600 531.300 ;
        RECT 572.550 531.150 573.750 533.400 ;
        RECT 585.150 532.200 586.950 534.000 ;
        RECT 589.200 533.550 594.150 534.600 ;
        RECT 592.350 532.800 594.150 533.550 ;
        RECT 595.650 532.800 597.450 534.600 ;
        RECT 598.950 533.400 601.050 535.500 ;
        RECT 604.050 533.400 605.850 539.400 ;
        RECT 586.050 531.900 586.950 532.200 ;
        RECT 596.100 531.900 597.150 532.800 ;
        RECT 560.100 528.150 561.900 529.950 ;
        RECT 550.950 524.850 553.200 526.950 ;
        RECT 556.950 524.850 559.050 526.950 ;
        RECT 559.950 526.050 562.050 528.150 ;
        RECT 563.850 526.950 565.050 530.250 ;
        RECT 562.950 524.850 565.050 526.950 ;
        RECT 572.550 529.050 577.050 531.150 ;
        RECT 586.050 531.000 597.150 531.900 ;
        RECT 526.950 515.550 531.450 516.450 ;
        RECT 526.950 514.950 529.050 515.550 ;
        RECT 536.400 513.600 537.600 521.850 ;
        RECT 549.150 521.400 551.100 522.300 ;
        RECT 545.400 520.500 551.100 521.400 ;
        RECT 545.400 513.600 546.600 520.500 ;
        RECT 552.000 519.600 553.200 524.850 ;
        RECT 557.100 523.050 558.900 524.850 ;
        RECT 562.950 519.600 564.150 524.850 ;
        RECT 565.950 521.850 568.050 523.950 ;
        RECT 565.950 520.050 567.750 521.850 ;
        RECT 572.550 519.600 573.750 529.050 ;
        RECT 574.950 527.250 578.850 529.050 ;
        RECT 574.950 526.950 577.050 527.250 ;
        RECT 586.050 526.950 586.950 531.000 ;
        RECT 596.100 529.800 597.150 531.000 ;
        RECT 596.100 528.600 603.000 529.800 ;
        RECT 596.100 528.000 597.900 528.600 ;
        RECT 602.100 527.850 603.000 528.600 ;
        RECT 599.100 526.950 600.900 527.700 ;
        RECT 586.050 524.850 589.050 526.950 ;
        RECT 592.950 525.900 600.900 526.950 ;
        RECT 602.100 526.050 603.900 527.850 ;
        RECT 592.950 524.850 595.050 525.900 ;
        RECT 574.950 521.400 576.750 523.200 ;
        RECT 575.850 520.200 580.050 521.400 ;
        RECT 586.050 520.200 586.950 524.850 ;
        RECT 594.750 521.100 596.550 521.400 ;
        RECT 536.400 507.600 538.200 513.600 ;
        RECT 545.400 507.600 547.200 513.600 ;
        RECT 551.700 507.600 553.500 519.600 ;
        RECT 562.500 507.600 564.300 519.600 ;
        RECT 572.550 507.600 574.350 519.600 ;
        RECT 577.950 519.300 580.050 520.200 ;
        RECT 580.950 519.300 586.950 520.200 ;
        RECT 588.150 520.800 596.550 521.100 ;
        RECT 604.950 520.800 605.850 533.400 ;
        RECT 611.400 534.300 613.200 539.400 ;
        RECT 617.400 534.300 619.200 539.400 ;
        RECT 611.400 532.950 619.200 534.300 ;
        RECT 620.400 533.400 622.200 539.400 ;
        RECT 620.400 531.300 621.600 533.400 ;
        RECT 631.200 532.200 633.000 539.400 ;
        RECT 638.400 536.400 640.200 539.400 ;
        RECT 617.850 530.250 621.600 531.300 ;
        RECT 629.400 531.300 633.000 532.200 ;
        RECT 639.000 532.500 640.200 536.400 ;
        RECT 644.700 533.400 646.500 539.400 ;
        RECT 639.000 531.600 644.100 532.500 ;
        RECT 614.100 528.150 615.900 529.950 ;
        RECT 610.950 524.850 613.050 526.950 ;
        RECT 613.950 526.050 616.050 528.150 ;
        RECT 617.850 526.950 619.050 530.250 ;
        RECT 616.950 524.850 619.050 526.950 ;
        RECT 626.100 525.150 627.900 526.950 ;
        RECT 611.100 523.050 612.900 524.850 ;
        RECT 588.150 520.200 605.850 520.800 ;
        RECT 580.950 518.400 581.850 519.300 ;
        RECT 579.150 516.600 581.850 518.400 ;
        RECT 582.750 518.100 584.550 518.400 ;
        RECT 588.150 518.100 589.050 520.200 ;
        RECT 594.750 519.600 605.850 520.200 ;
        RECT 616.950 519.600 618.150 524.850 ;
        RECT 619.950 521.850 622.050 523.950 ;
        RECT 625.950 523.050 628.050 525.150 ;
        RECT 629.400 523.950 630.600 531.300 ;
        RECT 642.150 530.700 644.100 531.600 ;
        RECT 632.100 525.150 633.900 526.950 ;
        RECT 628.950 521.850 631.050 523.950 ;
        RECT 631.950 523.050 634.050 525.150 ;
        RECT 637.950 524.850 640.050 526.950 ;
        RECT 638.100 523.050 639.900 524.850 ;
        RECT 642.150 522.300 643.050 530.700 ;
        RECT 645.000 526.950 646.200 533.400 ;
        RECT 658.200 532.200 660.000 539.400 ;
        RECT 670.200 532.200 672.000 539.400 ;
        RECT 682.800 532.500 684.600 539.400 ;
        RECT 688.800 532.500 690.600 539.400 ;
        RECT 694.800 532.500 696.600 539.400 ;
        RECT 700.800 532.500 702.600 539.400 ;
        RECT 709.800 536.400 711.600 539.400 ;
        RECT 719.400 536.400 721.200 539.400 ;
        RECT 656.400 531.300 660.000 532.200 ;
        RECT 668.400 531.300 672.000 532.200 ;
        RECT 681.900 531.300 684.600 532.500 ;
        RECT 686.700 531.300 690.600 532.500 ;
        RECT 692.700 531.300 696.600 532.500 ;
        RECT 698.700 531.300 702.600 532.500 ;
        RECT 643.950 524.850 646.200 526.950 ;
        RECT 653.100 525.150 654.900 526.950 ;
        RECT 619.950 520.050 621.750 521.850 ;
        RECT 582.750 517.200 589.050 518.100 ;
        RECT 589.950 518.700 591.750 519.300 ;
        RECT 589.950 517.500 597.450 518.700 ;
        RECT 582.750 516.600 584.550 517.200 ;
        RECT 596.250 516.600 597.450 517.500 ;
        RECT 577.950 513.600 581.850 515.700 ;
        RECT 586.950 515.550 588.750 516.300 ;
        RECT 591.750 515.550 593.550 516.300 ;
        RECT 586.950 514.500 593.550 515.550 ;
        RECT 596.250 514.500 601.050 516.600 ;
        RECT 580.050 507.600 581.850 513.600 ;
        RECT 587.850 507.600 589.650 514.500 ;
        RECT 596.250 513.600 597.450 514.500 ;
        RECT 595.650 507.600 597.450 513.600 ;
        RECT 604.050 507.600 605.850 519.600 ;
        RECT 616.500 507.600 618.300 519.600 ;
        RECT 629.400 513.600 630.600 521.850 ;
        RECT 642.150 521.400 644.100 522.300 ;
        RECT 638.400 520.500 644.100 521.400 ;
        RECT 638.400 513.600 639.600 520.500 ;
        RECT 645.000 519.600 646.200 524.850 ;
        RECT 652.950 523.050 655.050 525.150 ;
        RECT 656.400 523.950 657.600 531.300 ;
        RECT 659.100 525.150 660.900 526.950 ;
        RECT 665.100 525.150 666.900 526.950 ;
        RECT 655.950 521.850 658.050 523.950 ;
        RECT 658.950 523.050 661.050 525.150 ;
        RECT 664.950 523.050 667.050 525.150 ;
        RECT 668.400 523.950 669.600 531.300 ;
        RECT 681.900 528.150 682.800 531.300 ;
        RECT 686.700 530.400 687.900 531.300 ;
        RECT 692.700 530.400 693.900 531.300 ;
        RECT 698.700 530.400 699.900 531.300 ;
        RECT 683.700 529.200 687.900 530.400 ;
        RECT 683.700 528.600 685.500 529.200 ;
        RECT 671.100 525.150 672.900 526.950 ;
        RECT 679.950 526.050 682.800 528.150 ;
        RECT 667.950 521.850 670.050 523.950 ;
        RECT 670.950 523.050 673.050 525.150 ;
        RECT 629.400 507.600 631.200 513.600 ;
        RECT 638.400 507.600 640.200 513.600 ;
        RECT 644.700 507.600 646.500 519.600 ;
        RECT 656.400 513.600 657.600 521.850 ;
        RECT 668.400 513.600 669.600 521.850 ;
        RECT 681.900 521.700 682.800 526.050 ;
        RECT 686.700 521.700 687.900 529.200 ;
        RECT 689.700 529.200 693.900 530.400 ;
        RECT 689.700 528.600 691.500 529.200 ;
        RECT 692.700 521.700 693.900 529.200 ;
        RECT 695.700 529.200 699.900 530.400 ;
        RECT 695.700 528.600 697.500 529.200 ;
        RECT 698.700 521.700 699.900 529.200 ;
        RECT 701.100 528.150 702.900 529.950 ;
        RECT 710.400 528.150 711.600 536.400 ;
        RECT 720.000 529.950 721.050 536.400 ;
        RECT 733.200 532.200 735.000 539.400 ;
        RECT 700.950 526.050 703.050 528.150 ;
        RECT 709.950 526.050 712.050 528.150 ;
        RECT 712.950 527.850 715.050 529.950 ;
        RECT 718.950 527.850 721.050 529.950 ;
        RECT 713.100 526.050 714.900 527.850 ;
        RECT 681.900 520.500 684.600 521.700 ;
        RECT 686.700 520.500 690.600 521.700 ;
        RECT 692.700 520.500 696.600 521.700 ;
        RECT 698.700 520.500 702.600 521.700 ;
        RECT 656.400 507.600 658.200 513.600 ;
        RECT 668.400 507.600 670.200 513.600 ;
        RECT 682.800 507.600 684.600 520.500 ;
        RECT 688.800 507.600 690.600 520.500 ;
        RECT 694.800 507.600 696.600 520.500 ;
        RECT 700.800 507.600 702.600 520.500 ;
        RECT 710.400 513.600 711.600 526.050 ;
        RECT 715.950 524.850 718.050 526.950 ;
        RECT 716.100 523.050 717.900 524.850 ;
        RECT 720.000 520.650 721.050 527.850 ;
        RECT 731.400 531.300 735.000 532.200 ;
        RECT 746.400 536.400 748.200 539.400 ;
        RECT 721.950 524.850 724.050 526.950 ;
        RECT 728.100 525.150 729.900 526.950 ;
        RECT 722.100 523.050 723.900 524.850 ;
        RECT 727.950 523.050 730.050 525.150 ;
        RECT 731.400 523.950 732.600 531.300 ;
        RECT 742.950 527.850 745.050 529.950 ;
        RECT 746.400 528.150 747.600 536.400 ;
        RECT 754.500 533.400 756.300 539.400 ;
        RECT 760.800 536.400 762.600 539.400 ;
        RECT 734.100 525.150 735.900 526.950 ;
        RECT 743.100 526.050 744.900 527.850 ;
        RECT 745.950 526.050 748.050 528.150 ;
        RECT 754.800 526.950 756.000 533.400 ;
        RECT 760.800 532.500 762.000 536.400 ;
        RECT 756.900 531.600 762.000 532.500 ;
        RECT 756.900 530.700 758.850 531.600 ;
        RECT 730.950 521.850 733.050 523.950 ;
        RECT 733.950 523.050 736.050 525.150 ;
        RECT 720.000 519.600 722.400 520.650 ;
        RECT 709.800 507.600 711.600 513.600 ;
        RECT 720.600 507.600 722.400 519.600 ;
        RECT 731.400 513.600 732.600 521.850 ;
        RECT 746.400 513.600 747.600 526.050 ;
        RECT 754.800 524.850 757.050 526.950 ;
        RECT 754.800 519.600 756.000 524.850 ;
        RECT 757.950 522.300 758.850 530.700 ;
        RECT 760.950 524.850 763.050 526.950 ;
        RECT 761.100 523.050 762.900 524.850 ;
        RECT 756.900 521.400 758.850 522.300 ;
        RECT 756.900 520.500 762.600 521.400 ;
        RECT 731.400 507.600 733.200 513.600 ;
        RECT 746.400 507.600 748.200 513.600 ;
        RECT 754.500 507.600 756.300 519.600 ;
        RECT 761.400 513.600 762.600 520.500 ;
        RECT 760.800 507.600 762.600 513.600 ;
        RECT 7.800 497.400 9.600 503.400 ;
        RECT 19.800 497.400 21.600 503.400 ;
        RECT 8.400 484.950 9.600 497.400 ;
        RECT 20.400 489.150 21.600 497.400 ;
        RECT 31.800 491.400 33.600 503.400 ;
        RECT 34.800 492.300 36.600 503.400 ;
        RECT 40.800 492.300 42.600 503.400 ;
        RECT 46.800 497.400 48.600 503.400 ;
        RECT 34.800 491.400 42.600 492.300 ;
        RECT 47.700 497.100 48.600 497.400 ;
        RECT 52.800 497.400 54.600 503.400 ;
        RECT 64.800 497.400 66.600 503.400 ;
        RECT 74.400 497.400 76.200 503.400 ;
        RECT 52.800 497.100 54.300 497.400 ;
        RECT 47.700 496.200 54.300 497.100 ;
        RECT 16.950 485.850 19.050 487.950 ;
        RECT 19.950 487.050 22.050 489.150 ;
        RECT 7.950 482.850 10.050 484.950 ;
        RECT 11.100 483.150 12.900 484.950 ;
        RECT 17.100 484.050 18.900 485.850 ;
        RECT 8.400 474.600 9.600 482.850 ;
        RECT 10.950 481.050 13.050 483.150 ;
        RECT 20.400 479.700 21.600 487.050 ;
        RECT 22.950 485.850 25.050 487.950 ;
        RECT 32.400 486.150 33.300 491.400 ;
        RECT 47.700 487.950 48.600 496.200 ;
        RECT 58.950 493.950 61.050 496.050 ;
        RECT 53.100 492.150 54.900 493.950 ;
        RECT 49.950 489.150 51.750 490.950 ;
        RECT 52.950 490.050 55.050 492.150 ;
        RECT 56.100 489.150 57.900 490.950 ;
        RECT 23.100 484.050 24.900 485.850 ;
        RECT 31.950 484.050 34.050 486.150 ;
        RECT 46.950 485.850 49.050 487.950 ;
        RECT 49.950 487.050 52.050 489.150 ;
        RECT 55.950 487.050 58.050 489.150 ;
        RECT 7.800 471.600 9.600 474.600 ;
        RECT 18.000 478.800 21.600 479.700 ;
        RECT 18.000 471.600 19.800 478.800 ;
        RECT 32.400 477.600 33.300 484.050 ;
        RECT 34.950 482.850 37.050 484.950 ;
        RECT 38.100 483.150 39.900 484.950 ;
        RECT 35.100 481.050 36.900 482.850 ;
        RECT 37.950 481.050 40.050 483.150 ;
        RECT 40.950 482.850 43.050 484.950 ;
        RECT 41.100 481.050 42.900 482.850 ;
        RECT 47.700 481.650 48.600 485.850 ;
        RECT 52.950 483.450 55.050 484.050 ;
        RECT 59.550 483.450 60.450 493.950 ;
        RECT 65.400 489.150 66.600 497.400 ;
        RECT 74.700 497.100 76.200 497.400 ;
        RECT 80.400 497.400 82.200 503.400 ;
        RECT 80.400 497.100 81.300 497.400 ;
        RECT 74.700 496.200 81.300 497.100 ;
        RECT 74.100 492.150 75.900 493.950 ;
        RECT 71.100 489.150 72.900 490.950 ;
        RECT 73.950 490.050 76.050 492.150 ;
        RECT 77.250 489.150 79.050 490.950 ;
        RECT 61.950 485.850 64.050 487.950 ;
        RECT 64.950 487.050 67.050 489.150 ;
        RECT 62.100 484.050 63.900 485.850 ;
        RECT 52.950 482.550 60.450 483.450 ;
        RECT 52.950 481.950 55.050 482.550 ;
        RECT 47.700 480.000 51.900 481.650 ;
        RECT 32.400 475.950 37.800 477.600 ;
        RECT 36.000 471.600 37.800 475.950 ;
        RECT 50.100 471.600 51.900 480.000 ;
        RECT 65.400 479.700 66.600 487.050 ;
        RECT 67.950 485.850 70.050 487.950 ;
        RECT 70.950 487.050 73.050 489.150 ;
        RECT 76.950 487.050 79.050 489.150 ;
        RECT 80.400 487.950 81.300 496.200 ;
        RECT 91.500 491.400 93.300 503.400 ;
        RECT 106.800 497.400 108.600 503.400 ;
        RECT 79.950 485.850 82.050 487.950 ;
        RECT 86.100 486.150 87.900 487.950 ;
        RECT 91.950 486.150 93.150 491.400 ;
        RECT 94.950 489.150 96.750 490.950 ;
        RECT 107.400 489.150 108.600 497.400 ;
        RECT 119.700 491.400 121.500 503.400 ;
        RECT 136.500 491.400 138.300 503.400 ;
        RECT 152.700 491.400 154.500 503.400 ;
        RECT 167.700 491.400 169.500 503.400 ;
        RECT 179.400 497.400 181.200 503.400 ;
        RECT 116.250 489.150 118.050 490.950 ;
        RECT 94.950 487.050 97.050 489.150 ;
        RECT 68.100 484.050 69.900 485.850 ;
        RECT 80.400 481.650 81.300 485.850 ;
        RECT 85.950 484.050 88.050 486.150 ;
        RECT 88.950 482.850 91.050 484.950 ;
        RECT 91.950 484.050 94.050 486.150 ;
        RECT 103.950 485.850 106.050 487.950 ;
        RECT 106.950 487.050 109.050 489.150 ;
        RECT 104.100 484.050 105.900 485.850 ;
        RECT 63.000 478.800 66.600 479.700 ;
        RECT 77.100 480.000 81.300 481.650 ;
        RECT 89.100 481.050 90.900 482.850 ;
        RECT 92.850 480.750 94.050 484.050 ;
        RECT 63.000 471.600 64.800 478.800 ;
        RECT 77.100 471.600 78.900 480.000 ;
        RECT 92.850 479.700 96.600 480.750 ;
        RECT 107.400 479.700 108.600 487.050 ;
        RECT 109.950 485.850 112.050 487.950 ;
        RECT 115.950 487.050 118.050 489.150 ;
        RECT 119.850 486.150 121.050 491.400 ;
        RECT 125.100 486.150 126.900 487.950 ;
        RECT 131.100 486.150 132.900 487.950 ;
        RECT 136.950 486.150 138.150 491.400 ;
        RECT 139.950 489.150 141.750 490.950 ;
        RECT 149.250 489.150 151.050 490.950 ;
        RECT 139.950 487.050 142.050 489.150 ;
        RECT 148.950 487.050 151.050 489.150 ;
        RECT 152.850 486.150 154.050 491.400 ;
        RECT 164.250 489.150 166.050 490.950 ;
        RECT 158.100 486.150 159.900 487.950 ;
        RECT 163.950 487.050 166.050 489.150 ;
        RECT 167.850 486.150 169.050 491.400 ;
        RECT 173.100 486.150 174.900 487.950 ;
        RECT 110.100 484.050 111.900 485.850 ;
        RECT 118.950 484.050 121.050 486.150 ;
        RECT 118.950 480.750 120.150 484.050 ;
        RECT 121.950 482.850 124.050 484.950 ;
        RECT 124.950 484.050 127.050 486.150 ;
        RECT 130.950 484.050 133.050 486.150 ;
        RECT 133.950 482.850 136.050 484.950 ;
        RECT 136.950 484.050 139.050 486.150 ;
        RECT 122.100 481.050 123.900 482.850 ;
        RECT 134.100 481.050 135.900 482.850 ;
        RECT 86.400 476.700 94.200 478.050 ;
        RECT 86.400 471.600 88.200 476.700 ;
        RECT 92.400 471.600 94.200 476.700 ;
        RECT 95.400 477.600 96.600 479.700 ;
        RECT 105.000 478.800 108.600 479.700 ;
        RECT 116.400 479.700 120.150 480.750 ;
        RECT 137.850 480.750 139.050 484.050 ;
        RECT 151.950 484.050 154.050 486.150 ;
        RECT 151.950 480.750 153.150 484.050 ;
        RECT 154.950 482.850 157.050 484.950 ;
        RECT 157.950 484.050 160.050 486.150 ;
        RECT 166.950 484.050 169.050 486.150 ;
        RECT 155.100 481.050 156.900 482.850 ;
        RECT 166.950 480.750 168.150 484.050 ;
        RECT 169.950 482.850 172.050 484.950 ;
        RECT 172.950 484.050 175.050 486.150 ;
        RECT 179.400 484.950 180.600 497.400 ;
        RECT 187.800 491.400 189.600 503.400 ;
        RECT 190.800 492.300 192.600 503.400 ;
        RECT 196.800 492.300 198.600 503.400 ;
        RECT 190.800 491.400 198.600 492.300 ;
        RECT 203.400 497.400 205.200 503.400 ;
        RECT 218.400 497.400 220.200 503.400 ;
        RECT 188.400 486.150 189.300 491.400 ;
        RECT 203.400 489.150 204.600 497.400 ;
        RECT 176.100 483.150 177.900 484.950 ;
        RECT 170.100 481.050 171.900 482.850 ;
        RECT 175.950 481.050 178.050 483.150 ;
        RECT 178.950 482.850 181.050 484.950 ;
        RECT 187.950 484.050 190.050 486.150 ;
        RECT 199.950 485.850 202.050 487.950 ;
        RECT 202.950 487.050 205.050 489.150 ;
        RECT 137.850 479.700 141.600 480.750 ;
        RECT 95.400 471.600 97.200 477.600 ;
        RECT 105.000 471.600 106.800 478.800 ;
        RECT 116.400 477.600 117.600 479.700 ;
        RECT 115.800 471.600 117.600 477.600 ;
        RECT 118.800 476.700 126.600 478.050 ;
        RECT 118.800 471.600 120.600 476.700 ;
        RECT 124.800 471.600 126.600 476.700 ;
        RECT 131.400 476.700 139.200 478.050 ;
        RECT 131.400 471.600 133.200 476.700 ;
        RECT 137.400 471.600 139.200 476.700 ;
        RECT 140.400 477.600 141.600 479.700 ;
        RECT 149.400 479.700 153.150 480.750 ;
        RECT 164.400 479.700 168.150 480.750 ;
        RECT 149.400 477.600 150.600 479.700 ;
        RECT 140.400 471.600 142.200 477.600 ;
        RECT 148.800 471.600 150.600 477.600 ;
        RECT 151.800 476.700 159.600 478.050 ;
        RECT 164.400 477.600 165.600 479.700 ;
        RECT 151.800 471.600 153.600 476.700 ;
        RECT 157.800 471.600 159.600 476.700 ;
        RECT 163.800 471.600 165.600 477.600 ;
        RECT 166.800 476.700 174.600 478.050 ;
        RECT 166.800 471.600 168.600 476.700 ;
        RECT 172.800 471.600 174.600 476.700 ;
        RECT 179.400 474.600 180.600 482.850 ;
        RECT 188.400 477.600 189.300 484.050 ;
        RECT 190.950 482.850 193.050 484.950 ;
        RECT 194.100 483.150 195.900 484.950 ;
        RECT 191.100 481.050 192.900 482.850 ;
        RECT 193.950 481.050 196.050 483.150 ;
        RECT 196.950 482.850 199.050 484.950 ;
        RECT 200.100 484.050 201.900 485.850 ;
        RECT 197.100 481.050 198.900 482.850 ;
        RECT 203.400 479.700 204.600 487.050 ;
        RECT 205.950 485.850 208.050 487.950 ;
        RECT 206.100 484.050 207.900 485.850 ;
        RECT 218.400 484.950 219.600 497.400 ;
        RECT 228.900 491.400 232.200 503.400 ;
        RECT 251.700 491.400 253.500 503.400 ;
        RECT 267.600 491.400 269.400 503.400 ;
        RECT 274.950 493.950 277.050 496.050 ;
        RECT 224.100 486.150 225.900 487.950 ;
        RECT 230.400 486.150 231.600 491.400 ;
        RECT 248.250 489.150 250.050 490.950 ;
        RECT 235.950 486.150 237.750 487.950 ;
        RECT 247.950 487.050 250.050 489.150 ;
        RECT 251.850 486.150 253.050 491.400 ;
        RECT 267.600 490.350 270.000 491.400 ;
        RECT 257.100 486.150 258.900 487.950 ;
        RECT 266.100 486.150 267.900 487.950 ;
        RECT 215.100 483.150 216.900 484.950 ;
        RECT 214.950 481.050 217.050 483.150 ;
        RECT 217.950 482.850 220.050 484.950 ;
        RECT 223.950 484.050 226.050 486.150 ;
        RECT 226.950 482.850 229.050 484.950 ;
        RECT 229.950 484.050 232.050 486.150 ;
        RECT 203.400 478.800 207.000 479.700 ;
        RECT 188.400 475.950 193.800 477.600 ;
        RECT 179.400 471.600 181.200 474.600 ;
        RECT 192.000 471.600 193.800 475.950 ;
        RECT 205.200 471.600 207.000 478.800 ;
        RECT 218.400 474.600 219.600 482.850 ;
        RECT 227.100 481.050 228.900 482.850 ;
        RECT 230.400 480.150 231.600 484.050 ;
        RECT 232.950 482.850 235.050 484.950 ;
        RECT 235.950 484.050 238.050 486.150 ;
        RECT 250.950 484.050 253.050 486.150 ;
        RECT 232.500 481.050 234.300 482.850 ;
        RECT 250.950 480.750 252.150 484.050 ;
        RECT 253.950 482.850 256.050 484.950 ;
        RECT 256.950 484.050 259.050 486.150 ;
        RECT 265.950 484.050 268.050 486.150 ;
        RECT 268.950 483.150 270.000 490.350 ;
        RECT 272.100 486.150 273.900 487.950 ;
        RECT 271.950 484.050 274.050 486.150 ;
        RECT 254.100 481.050 255.900 482.850 ;
        RECT 268.950 481.050 271.050 483.150 ;
        RECT 230.400 479.100 234.600 480.150 ;
        RECT 224.400 477.000 232.200 477.900 ;
        RECT 233.700 477.600 234.600 479.100 ;
        RECT 248.400 479.700 252.150 480.750 ;
        RECT 248.400 477.600 249.600 479.700 ;
        RECT 218.400 471.600 220.200 474.600 ;
        RECT 224.400 471.600 226.200 477.000 ;
        RECT 230.400 472.500 232.200 477.000 ;
        RECT 233.400 473.400 235.200 477.600 ;
        RECT 236.400 472.500 238.200 477.600 ;
        RECT 230.400 471.600 238.200 472.500 ;
        RECT 247.800 471.600 249.600 477.600 ;
        RECT 250.800 476.700 258.600 478.050 ;
        RECT 250.800 471.600 252.600 476.700 ;
        RECT 256.800 471.600 258.600 476.700 ;
        RECT 268.950 474.600 270.000 481.050 ;
        RECT 275.550 480.450 276.450 493.950 ;
        RECT 282.600 491.400 284.400 503.400 ;
        RECT 292.800 502.500 300.600 503.400 ;
        RECT 292.800 491.400 294.600 502.500 ;
        RECT 282.600 490.350 285.000 491.400 ;
        RECT 281.100 486.150 282.900 487.950 ;
        RECT 280.950 484.050 283.050 486.150 ;
        RECT 283.950 483.150 285.000 490.350 ;
        RECT 295.800 490.500 297.600 501.600 ;
        RECT 298.800 492.600 300.600 502.500 ;
        RECT 304.800 492.600 306.600 503.400 ;
        RECT 298.800 491.700 306.600 492.600 ;
        RECT 308.550 491.400 310.350 503.400 ;
        RECT 316.050 497.400 317.850 503.400 ;
        RECT 313.950 495.300 317.850 497.400 ;
        RECT 323.850 496.500 325.650 503.400 ;
        RECT 331.650 497.400 333.450 503.400 ;
        RECT 332.250 496.500 333.450 497.400 ;
        RECT 322.950 495.450 329.550 496.500 ;
        RECT 322.950 494.700 324.750 495.450 ;
        RECT 327.750 494.700 329.550 495.450 ;
        RECT 332.250 494.400 337.050 496.500 ;
        RECT 315.150 492.600 317.850 494.400 ;
        RECT 318.750 493.800 320.550 494.400 ;
        RECT 318.750 492.900 325.050 493.800 ;
        RECT 332.250 493.500 333.450 494.400 ;
        RECT 318.750 492.600 320.550 492.900 ;
        RECT 316.950 491.700 317.850 492.600 ;
        RECT 295.800 489.600 299.850 490.500 ;
        RECT 287.100 486.150 288.900 487.950 ;
        RECT 293.100 486.150 294.900 487.950 ;
        RECT 298.950 486.150 299.850 489.600 ;
        RECT 304.950 486.150 306.750 487.950 ;
        RECT 286.950 484.050 289.050 486.150 ;
        RECT 292.950 484.050 295.050 486.150 ;
        RECT 283.950 481.050 286.050 483.150 ;
        RECT 295.950 482.850 298.050 484.950 ;
        RECT 298.950 484.050 301.050 486.150 ;
        RECT 296.250 481.050 298.050 482.850 ;
        RECT 280.950 480.450 283.050 481.050 ;
        RECT 275.550 479.550 283.050 480.450 ;
        RECT 280.950 478.950 283.050 479.550 ;
        RECT 283.950 474.600 285.000 481.050 ;
        RECT 300.000 477.600 301.050 484.050 ;
        RECT 301.950 482.850 304.050 484.950 ;
        RECT 304.950 484.050 307.050 486.150 ;
        RECT 301.950 481.050 303.750 482.850 ;
        RECT 308.550 481.950 309.750 491.400 ;
        RECT 313.950 490.800 316.050 491.700 ;
        RECT 316.950 490.800 322.950 491.700 ;
        RECT 311.850 489.600 316.050 490.800 ;
        RECT 310.950 487.800 312.750 489.600 ;
        RECT 322.050 486.150 322.950 490.800 ;
        RECT 324.150 490.800 325.050 492.900 ;
        RECT 325.950 492.300 333.450 493.500 ;
        RECT 325.950 491.700 327.750 492.300 ;
        RECT 340.050 491.400 341.850 503.400 ;
        RECT 330.750 490.800 341.850 491.400 ;
        RECT 324.150 490.200 341.850 490.800 ;
        RECT 324.150 489.900 332.550 490.200 ;
        RECT 330.750 489.600 332.550 489.900 ;
        RECT 322.050 484.050 325.050 486.150 ;
        RECT 328.950 485.100 331.050 486.150 ;
        RECT 328.950 484.050 336.900 485.100 ;
        RECT 310.950 483.750 313.050 484.050 ;
        RECT 310.950 481.950 314.850 483.750 ;
        RECT 308.550 479.850 313.050 481.950 ;
        RECT 322.050 480.000 322.950 484.050 ;
        RECT 335.100 483.300 336.900 484.050 ;
        RECT 338.100 483.150 339.900 484.950 ;
        RECT 332.100 482.400 333.900 483.000 ;
        RECT 338.100 482.400 339.000 483.150 ;
        RECT 332.100 481.200 339.000 482.400 ;
        RECT 332.100 480.000 333.150 481.200 ;
        RECT 308.550 477.600 309.750 479.850 ;
        RECT 322.050 479.100 333.150 480.000 ;
        RECT 322.050 478.800 322.950 479.100 ;
        RECT 268.800 471.600 270.600 474.600 ;
        RECT 283.800 471.600 285.600 474.600 ;
        RECT 300.000 471.600 301.800 477.600 ;
        RECT 308.550 471.600 310.350 477.600 ;
        RECT 313.950 476.700 316.050 477.600 ;
        RECT 321.150 477.000 322.950 478.800 ;
        RECT 332.100 478.200 333.150 479.100 ;
        RECT 328.350 477.450 330.150 478.200 ;
        RECT 313.950 475.500 317.700 476.700 ;
        RECT 316.650 474.600 317.700 475.500 ;
        RECT 325.200 476.400 330.150 477.450 ;
        RECT 331.650 476.400 333.450 478.200 ;
        RECT 340.950 477.600 341.850 490.200 ;
        RECT 344.400 497.400 346.200 503.400 ;
        RECT 344.400 490.500 345.600 497.400 ;
        RECT 350.700 491.400 352.500 503.400 ;
        RECT 359.400 497.400 361.200 503.400 ;
        RECT 344.400 489.600 350.100 490.500 ;
        RECT 348.150 488.700 350.100 489.600 ;
        RECT 344.100 486.150 345.900 487.950 ;
        RECT 343.950 484.050 346.050 486.150 ;
        RECT 348.150 480.300 349.050 488.700 ;
        RECT 351.000 486.150 352.200 491.400 ;
        RECT 359.400 489.150 360.600 497.400 ;
        RECT 374.700 491.400 376.500 503.400 ;
        RECT 392.700 491.400 394.500 503.400 ;
        RECT 403.200 491.400 405.000 503.400 ;
        RECT 409.800 497.400 411.600 503.400 ;
        RECT 371.250 489.150 373.050 490.950 ;
        RECT 349.950 484.050 352.200 486.150 ;
        RECT 355.950 485.850 358.050 487.950 ;
        RECT 358.950 487.050 361.050 489.150 ;
        RECT 356.100 484.050 357.900 485.850 ;
        RECT 348.150 479.400 350.100 480.300 ;
        RECT 325.200 474.600 326.250 476.400 ;
        RECT 334.950 475.500 337.050 477.600 ;
        RECT 334.950 474.600 336.000 475.500 ;
        RECT 316.650 471.600 318.450 474.600 ;
        RECT 324.450 471.600 326.250 474.600 ;
        RECT 332.250 473.700 336.000 474.600 ;
        RECT 332.250 471.600 334.050 473.700 ;
        RECT 340.050 471.600 341.850 477.600 ;
        RECT 345.000 478.500 350.100 479.400 ;
        RECT 345.000 474.600 346.200 478.500 ;
        RECT 351.000 477.600 352.200 484.050 ;
        RECT 359.400 479.700 360.600 487.050 ;
        RECT 361.950 485.850 364.050 487.950 ;
        RECT 370.950 487.050 373.050 489.150 ;
        RECT 374.850 486.150 376.050 491.400 ;
        RECT 389.250 489.150 391.050 490.950 ;
        RECT 380.100 486.150 381.900 487.950 ;
        RECT 388.950 487.050 391.050 489.150 ;
        RECT 392.850 486.150 394.050 491.400 ;
        RECT 398.100 486.150 399.900 487.950 ;
        RECT 403.950 486.150 405.000 491.400 ;
        RECT 362.100 484.050 363.900 485.850 ;
        RECT 373.950 484.050 376.050 486.150 ;
        RECT 373.950 480.750 375.150 484.050 ;
        RECT 376.950 482.850 379.050 484.950 ;
        RECT 379.950 484.050 382.050 486.150 ;
        RECT 391.950 484.050 394.050 486.150 ;
        RECT 377.100 481.050 378.900 482.850 ;
        RECT 391.950 480.750 393.150 484.050 ;
        RECT 394.950 482.850 397.050 484.950 ;
        RECT 397.950 484.050 400.050 486.150 ;
        RECT 403.950 484.050 406.050 486.150 ;
        RECT 406.950 485.850 409.050 487.950 ;
        RECT 407.100 484.050 408.900 485.850 ;
        RECT 395.100 481.050 396.900 482.850 ;
        RECT 371.400 479.700 375.150 480.750 ;
        RECT 389.400 479.700 393.150 480.750 ;
        RECT 359.400 478.800 363.000 479.700 ;
        RECT 344.400 471.600 346.200 474.600 ;
        RECT 350.700 471.600 352.500 477.600 ;
        RECT 361.200 471.600 363.000 478.800 ;
        RECT 371.400 477.600 372.600 479.700 ;
        RECT 370.800 471.600 372.600 477.600 ;
        RECT 373.800 476.700 381.600 478.050 ;
        RECT 389.400 477.600 390.600 479.700 ;
        RECT 373.800 471.600 375.600 476.700 ;
        RECT 379.800 471.600 381.600 476.700 ;
        RECT 388.800 471.600 390.600 477.600 ;
        RECT 391.800 476.700 399.600 478.050 ;
        RECT 391.800 471.600 393.600 476.700 ;
        RECT 397.800 471.600 399.600 476.700 ;
        RECT 403.950 477.600 405.000 484.050 ;
        RECT 410.400 480.300 411.450 497.400 ;
        RECT 418.800 491.400 420.600 503.400 ;
        RECT 413.100 486.150 414.900 487.950 ;
        RECT 419.400 486.150 420.600 491.400 ;
        RECT 425.550 491.400 427.350 503.400 ;
        RECT 433.050 497.400 434.850 503.400 ;
        RECT 430.950 495.300 434.850 497.400 ;
        RECT 440.850 496.500 442.650 503.400 ;
        RECT 448.650 497.400 450.450 503.400 ;
        RECT 449.250 496.500 450.450 497.400 ;
        RECT 439.950 495.450 446.550 496.500 ;
        RECT 439.950 494.700 441.750 495.450 ;
        RECT 444.750 494.700 446.550 495.450 ;
        RECT 449.250 494.400 454.050 496.500 ;
        RECT 432.150 492.600 434.850 494.400 ;
        RECT 435.750 493.800 437.550 494.400 ;
        RECT 435.750 492.900 442.050 493.800 ;
        RECT 449.250 493.500 450.450 494.400 ;
        RECT 435.750 492.600 437.550 492.900 ;
        RECT 433.950 491.700 434.850 492.600 ;
        RECT 412.950 484.050 415.050 486.150 ;
        RECT 418.950 484.050 421.050 486.150 ;
        RECT 407.100 479.100 414.600 480.300 ;
        RECT 407.100 478.500 408.900 479.100 ;
        RECT 403.950 476.100 407.100 477.600 ;
        RECT 405.300 471.600 407.100 476.100 ;
        RECT 412.800 471.600 414.600 479.100 ;
        RECT 419.400 477.600 420.600 484.050 ;
        RECT 421.950 482.850 424.050 484.950 ;
        RECT 422.100 481.050 423.900 482.850 ;
        RECT 425.550 481.950 426.750 491.400 ;
        RECT 430.950 490.800 433.050 491.700 ;
        RECT 433.950 490.800 439.950 491.700 ;
        RECT 428.850 489.600 433.050 490.800 ;
        RECT 427.950 487.800 429.750 489.600 ;
        RECT 439.050 486.150 439.950 490.800 ;
        RECT 441.150 490.800 442.050 492.900 ;
        RECT 442.950 492.300 450.450 493.500 ;
        RECT 442.950 491.700 444.750 492.300 ;
        RECT 457.050 491.400 458.850 503.400 ;
        RECT 447.750 490.800 458.850 491.400 ;
        RECT 441.150 490.200 458.850 490.800 ;
        RECT 466.800 490.500 468.600 503.400 ;
        RECT 472.800 490.500 474.600 503.400 ;
        RECT 478.800 490.500 480.600 503.400 ;
        RECT 484.800 490.500 486.600 503.400 ;
        RECT 497.700 491.400 499.500 503.400 ;
        RECT 508.800 497.400 510.600 503.400 ;
        RECT 441.150 489.900 449.550 490.200 ;
        RECT 447.750 489.600 449.550 489.900 ;
        RECT 439.050 484.050 442.050 486.150 ;
        RECT 445.950 485.100 448.050 486.150 ;
        RECT 445.950 484.050 453.900 485.100 ;
        RECT 427.950 483.750 430.050 484.050 ;
        RECT 427.950 481.950 431.850 483.750 ;
        RECT 418.800 471.600 420.600 477.600 ;
        RECT 425.550 479.850 430.050 481.950 ;
        RECT 439.050 480.000 439.950 484.050 ;
        RECT 452.100 483.300 453.900 484.050 ;
        RECT 455.100 483.150 456.900 484.950 ;
        RECT 449.100 482.400 450.900 483.000 ;
        RECT 455.100 482.400 456.000 483.150 ;
        RECT 449.100 481.200 456.000 482.400 ;
        RECT 449.100 480.000 450.150 481.200 ;
        RECT 425.550 477.600 426.750 479.850 ;
        RECT 439.050 479.100 450.150 480.000 ;
        RECT 439.050 478.800 439.950 479.100 ;
        RECT 425.550 471.600 427.350 477.600 ;
        RECT 430.950 476.700 433.050 477.600 ;
        RECT 438.150 477.000 439.950 478.800 ;
        RECT 449.100 478.200 450.150 479.100 ;
        RECT 445.350 477.450 447.150 478.200 ;
        RECT 430.950 475.500 434.700 476.700 ;
        RECT 433.650 474.600 434.700 475.500 ;
        RECT 442.200 476.400 447.150 477.450 ;
        RECT 448.650 476.400 450.450 478.200 ;
        RECT 457.950 477.600 458.850 490.200 ;
        RECT 465.900 489.300 468.600 490.500 ;
        RECT 470.700 489.300 474.600 490.500 ;
        RECT 476.700 489.300 480.600 490.500 ;
        RECT 482.700 489.300 486.600 490.500 ;
        RECT 465.900 484.950 466.800 489.300 ;
        RECT 463.950 482.850 466.800 484.950 ;
        RECT 465.900 479.700 466.800 482.850 ;
        RECT 467.700 481.800 469.500 482.400 ;
        RECT 470.700 481.800 471.900 489.300 ;
        RECT 467.700 480.600 471.900 481.800 ;
        RECT 473.700 481.800 475.500 482.400 ;
        RECT 476.700 481.800 477.900 489.300 ;
        RECT 473.700 480.600 477.900 481.800 ;
        RECT 479.700 481.800 481.500 482.400 ;
        RECT 482.700 481.800 483.900 489.300 ;
        RECT 494.250 489.150 496.050 490.950 ;
        RECT 493.950 487.050 496.050 489.150 ;
        RECT 497.850 486.150 499.050 491.400 ;
        RECT 503.100 486.150 504.900 487.950 ;
        RECT 484.950 482.850 487.050 484.950 ;
        RECT 496.950 484.050 499.050 486.150 ;
        RECT 479.700 480.600 483.900 481.800 ;
        RECT 485.100 481.050 486.900 482.850 ;
        RECT 496.950 480.750 498.150 484.050 ;
        RECT 499.950 482.850 502.050 484.950 ;
        RECT 502.950 484.050 505.050 486.150 ;
        RECT 509.400 484.950 510.600 497.400 ;
        RECT 518.400 497.400 520.200 503.400 ;
        RECT 518.400 489.150 519.600 497.400 ;
        RECT 529.800 491.400 531.600 503.400 ;
        RECT 532.800 492.300 534.600 503.400 ;
        RECT 538.800 492.300 540.600 503.400 ;
        RECT 544.800 497.400 546.600 503.400 ;
        RECT 532.800 491.400 540.600 492.300 ;
        RECT 545.700 497.100 546.600 497.400 ;
        RECT 550.800 497.400 552.600 503.400 ;
        RECT 550.800 497.100 552.300 497.400 ;
        RECT 545.700 496.200 552.300 497.100 ;
        RECT 514.950 485.850 517.050 487.950 ;
        RECT 517.950 487.050 520.050 489.150 ;
        RECT 508.950 482.850 511.050 484.950 ;
        RECT 512.100 483.150 513.900 484.950 ;
        RECT 515.100 484.050 516.900 485.850 ;
        RECT 500.100 481.050 501.900 482.850 ;
        RECT 470.700 479.700 471.900 480.600 ;
        RECT 476.700 479.700 477.900 480.600 ;
        RECT 482.700 479.700 483.900 480.600 ;
        RECT 494.400 479.700 498.150 480.750 ;
        RECT 465.900 478.500 468.600 479.700 ;
        RECT 470.700 478.500 474.600 479.700 ;
        RECT 476.700 478.500 480.600 479.700 ;
        RECT 482.700 478.500 486.600 479.700 ;
        RECT 442.200 474.600 443.250 476.400 ;
        RECT 451.950 475.500 454.050 477.600 ;
        RECT 451.950 474.600 453.000 475.500 ;
        RECT 433.650 471.600 435.450 474.600 ;
        RECT 441.450 471.600 443.250 474.600 ;
        RECT 449.250 473.700 453.000 474.600 ;
        RECT 449.250 471.600 451.050 473.700 ;
        RECT 457.050 471.600 458.850 477.600 ;
        RECT 466.800 471.600 468.600 478.500 ;
        RECT 472.800 471.600 474.600 478.500 ;
        RECT 478.800 471.600 480.600 478.500 ;
        RECT 484.800 471.600 486.600 478.500 ;
        RECT 494.400 477.600 495.600 479.700 ;
        RECT 493.800 471.600 495.600 477.600 ;
        RECT 496.800 476.700 504.600 478.050 ;
        RECT 496.800 471.600 498.600 476.700 ;
        RECT 502.800 471.600 504.600 476.700 ;
        RECT 509.400 474.600 510.600 482.850 ;
        RECT 511.950 481.050 514.050 483.150 ;
        RECT 518.400 479.700 519.600 487.050 ;
        RECT 520.950 485.850 523.050 487.950 ;
        RECT 530.400 486.150 531.300 491.400 ;
        RECT 545.700 487.950 546.600 496.200 ;
        RECT 551.100 492.150 552.900 493.950 ;
        RECT 547.950 489.150 549.750 490.950 ;
        RECT 550.950 490.050 553.050 492.150 ;
        RECT 561.600 491.400 563.400 503.400 ;
        RECT 554.100 489.150 555.900 490.950 ;
        RECT 561.000 490.350 563.400 491.400 ;
        RECT 572.400 497.400 574.200 503.400 ;
        RECT 521.100 484.050 522.900 485.850 ;
        RECT 529.950 484.050 532.050 486.150 ;
        RECT 544.950 485.850 547.050 487.950 ;
        RECT 547.950 487.050 550.050 489.150 ;
        RECT 553.950 487.050 556.050 489.150 ;
        RECT 557.100 486.150 558.900 487.950 ;
        RECT 518.400 478.800 522.000 479.700 ;
        RECT 508.800 471.600 510.600 474.600 ;
        RECT 520.200 471.600 522.000 478.800 ;
        RECT 530.400 477.600 531.300 484.050 ;
        RECT 532.950 482.850 535.050 484.950 ;
        RECT 536.100 483.150 537.900 484.950 ;
        RECT 533.100 481.050 534.900 482.850 ;
        RECT 535.950 481.050 538.050 483.150 ;
        RECT 538.950 482.850 541.050 484.950 ;
        RECT 539.100 481.050 540.900 482.850 ;
        RECT 545.700 481.650 546.600 485.850 ;
        RECT 556.950 484.050 559.050 486.150 ;
        RECT 561.000 483.150 562.050 490.350 ;
        RECT 572.400 489.150 573.600 497.400 ;
        RECT 574.950 492.450 577.050 493.050 ;
        RECT 581.400 492.600 583.200 503.400 ;
        RECT 587.400 502.500 595.200 503.400 ;
        RECT 587.400 492.600 589.200 502.500 ;
        RECT 574.950 491.550 579.450 492.450 ;
        RECT 581.400 491.700 589.200 492.600 ;
        RECT 574.950 490.950 577.050 491.550 ;
        RECT 563.100 486.150 564.900 487.950 ;
        RECT 562.950 484.050 565.050 486.150 ;
        RECT 568.950 485.850 571.050 487.950 ;
        RECT 571.950 487.050 574.050 489.150 ;
        RECT 569.100 484.050 570.900 485.850 ;
        RECT 545.700 480.000 549.900 481.650 ;
        RECT 559.950 481.050 562.050 483.150 ;
        RECT 530.400 475.950 535.800 477.600 ;
        RECT 534.000 471.600 535.800 475.950 ;
        RECT 548.100 471.600 549.900 480.000 ;
        RECT 561.000 474.600 562.050 481.050 ;
        RECT 572.400 479.700 573.600 487.050 ;
        RECT 574.950 485.850 577.050 487.950 ;
        RECT 575.100 484.050 576.900 485.850 ;
        RECT 578.550 480.450 579.450 491.550 ;
        RECT 590.400 490.500 592.200 501.600 ;
        RECT 593.400 491.400 595.200 502.500 ;
        RECT 604.800 497.400 606.600 503.400 ;
        RECT 601.950 492.450 604.050 493.050 ;
        RECT 599.550 491.550 604.050 492.450 ;
        RECT 588.150 489.600 592.200 490.500 ;
        RECT 581.250 486.150 583.050 487.950 ;
        RECT 588.150 486.150 589.050 489.600 ;
        RECT 593.100 486.150 594.900 487.950 ;
        RECT 580.950 484.050 583.050 486.150 ;
        RECT 583.950 482.850 586.050 484.950 ;
        RECT 584.250 481.050 586.050 482.850 ;
        RECT 586.950 484.050 589.050 486.150 ;
        RECT 580.950 480.450 583.050 481.050 ;
        RECT 572.400 478.800 576.000 479.700 ;
        RECT 578.550 479.550 583.050 480.450 ;
        RECT 580.950 478.950 583.050 479.550 ;
        RECT 560.400 471.600 562.200 474.600 ;
        RECT 574.200 471.600 576.000 478.800 ;
        RECT 586.950 477.600 588.000 484.050 ;
        RECT 589.950 482.850 592.050 484.950 ;
        RECT 592.950 484.050 595.050 486.150 ;
        RECT 589.950 481.050 591.750 482.850 ;
        RECT 595.950 480.450 598.050 481.050 ;
        RECT 599.550 480.450 600.450 491.550 ;
        RECT 601.950 490.950 604.050 491.550 ;
        RECT 605.400 489.150 606.600 497.400 ;
        RECT 607.950 492.450 610.050 493.050 ;
        RECT 607.950 491.550 612.450 492.450 ;
        RECT 607.950 490.950 610.050 491.550 ;
        RECT 601.950 485.850 604.050 487.950 ;
        RECT 604.950 487.050 607.050 489.150 ;
        RECT 602.100 484.050 603.900 485.850 ;
        RECT 595.950 479.550 600.450 480.450 ;
        RECT 605.400 479.700 606.600 487.050 ;
        RECT 607.950 485.850 610.050 487.950 ;
        RECT 608.100 484.050 609.900 485.850 ;
        RECT 595.950 478.950 598.050 479.550 ;
        RECT 586.200 471.600 588.000 477.600 ;
        RECT 603.000 478.800 606.600 479.700 ;
        RECT 607.950 480.450 610.050 481.050 ;
        RECT 611.550 480.450 612.450 491.550 ;
        RECT 618.600 491.400 620.400 503.400 ;
        RECT 628.800 497.400 630.600 503.400 ;
        RECT 618.000 490.350 620.400 491.400 ;
        RECT 614.100 486.150 615.900 487.950 ;
        RECT 613.950 484.050 616.050 486.150 ;
        RECT 618.000 483.150 619.050 490.350 ;
        RECT 620.100 486.150 621.900 487.950 ;
        RECT 619.950 484.050 622.050 486.150 ;
        RECT 629.400 484.950 630.600 497.400 ;
        RECT 643.500 491.400 645.300 503.400 ;
        RECT 661.800 491.400 665.100 503.400 ;
        RECT 675.600 491.400 677.400 503.400 ;
        RECT 686.400 497.400 688.200 503.400 ;
        RECT 682.950 492.450 685.050 493.050 ;
        RECT 638.100 486.150 639.900 487.950 ;
        RECT 643.950 486.150 645.150 491.400 ;
        RECT 646.950 489.150 648.750 490.950 ;
        RECT 646.950 487.050 649.050 489.150 ;
        RECT 656.250 486.150 658.050 487.950 ;
        RECT 662.400 486.150 663.600 491.400 ;
        RECT 675.000 490.350 677.400 491.400 ;
        RECT 680.550 491.550 685.050 492.450 ;
        RECT 668.100 486.150 669.900 487.950 ;
        RECT 671.100 486.150 672.900 487.950 ;
        RECT 616.950 481.050 619.050 483.150 ;
        RECT 628.950 482.850 631.050 484.950 ;
        RECT 632.100 483.150 633.900 484.950 ;
        RECT 637.950 484.050 640.050 486.150 ;
        RECT 607.950 479.550 612.450 480.450 ;
        RECT 607.950 478.950 610.050 479.550 ;
        RECT 603.000 471.600 604.800 478.800 ;
        RECT 618.000 474.600 619.050 481.050 ;
        RECT 629.400 474.600 630.600 482.850 ;
        RECT 631.950 481.050 634.050 483.150 ;
        RECT 640.950 482.850 643.050 484.950 ;
        RECT 643.950 484.050 646.050 486.150 ;
        RECT 655.950 484.050 658.050 486.150 ;
        RECT 641.100 481.050 642.900 482.850 ;
        RECT 644.850 480.750 646.050 484.050 ;
        RECT 658.950 482.850 661.050 484.950 ;
        RECT 661.950 484.050 664.050 486.150 ;
        RECT 659.700 481.050 661.500 482.850 ;
        RECT 644.850 479.700 648.600 480.750 ;
        RECT 662.400 480.150 663.600 484.050 ;
        RECT 664.950 482.850 667.050 484.950 ;
        RECT 667.950 484.050 670.050 486.150 ;
        RECT 670.950 484.050 673.050 486.150 ;
        RECT 675.000 483.150 676.050 490.350 ;
        RECT 677.100 486.150 678.900 487.950 ;
        RECT 676.950 484.050 679.050 486.150 ;
        RECT 665.100 481.050 666.900 482.850 ;
        RECT 673.950 481.050 676.050 483.150 ;
        RECT 617.400 471.600 619.200 474.600 ;
        RECT 628.800 471.600 630.600 474.600 ;
        RECT 638.400 476.700 646.200 478.050 ;
        RECT 638.400 471.600 640.200 476.700 ;
        RECT 644.400 471.600 646.200 476.700 ;
        RECT 647.400 477.600 648.600 479.700 ;
        RECT 659.400 479.100 663.600 480.150 ;
        RECT 659.400 477.600 660.300 479.100 ;
        RECT 647.400 471.600 649.200 477.600 ;
        RECT 655.800 472.500 657.600 477.600 ;
        RECT 658.800 473.400 660.600 477.600 ;
        RECT 661.800 477.000 669.600 477.900 ;
        RECT 661.800 472.500 663.600 477.000 ;
        RECT 655.800 471.600 663.600 472.500 ;
        RECT 667.800 471.600 669.600 477.000 ;
        RECT 675.000 474.600 676.050 481.050 ;
        RECT 676.950 480.450 679.050 481.050 ;
        RECT 680.550 480.450 681.450 491.550 ;
        RECT 682.950 490.950 685.050 491.550 ;
        RECT 686.400 489.150 687.600 497.400 ;
        RECT 701.700 491.400 703.500 503.400 ;
        RECT 715.500 491.400 717.300 503.400 ;
        RECT 698.250 489.150 700.050 490.950 ;
        RECT 682.950 485.850 685.050 487.950 ;
        RECT 685.950 487.050 688.050 489.150 ;
        RECT 683.100 484.050 684.900 485.850 ;
        RECT 676.950 479.550 681.450 480.450 ;
        RECT 686.400 479.700 687.600 487.050 ;
        RECT 688.950 485.850 691.050 487.950 ;
        RECT 697.950 487.050 700.050 489.150 ;
        RECT 694.950 486.450 697.050 487.050 ;
        RECT 689.100 484.050 690.900 485.850 ;
        RECT 692.550 485.550 697.050 486.450 ;
        RECT 701.850 486.150 703.050 491.400 ;
        RECT 707.100 486.150 708.900 487.950 ;
        RECT 710.100 486.150 711.900 487.950 ;
        RECT 715.950 486.150 717.150 491.400 ;
        RECT 721.950 490.950 724.050 493.050 ;
        RECT 729.600 491.400 731.400 503.400 ;
        RECT 744.300 492.900 746.100 503.400 ;
        RECT 718.950 489.150 720.750 490.950 ;
        RECT 718.950 487.050 721.050 489.150 ;
        RECT 692.550 481.050 693.450 485.550 ;
        RECT 694.950 484.950 697.050 485.550 ;
        RECT 700.950 484.050 703.050 486.150 ;
        RECT 676.950 478.950 679.050 479.550 ;
        RECT 686.400 478.800 690.000 479.700 ;
        RECT 691.950 478.950 694.050 481.050 ;
        RECT 700.950 480.750 702.150 484.050 ;
        RECT 703.950 482.850 706.050 484.950 ;
        RECT 706.950 484.050 709.050 486.150 ;
        RECT 709.950 484.050 712.050 486.150 ;
        RECT 712.950 482.850 715.050 484.950 ;
        RECT 715.950 484.050 718.050 486.150 ;
        RECT 704.100 481.050 705.900 482.850 ;
        RECT 713.100 481.050 714.900 482.850 ;
        RECT 698.400 479.700 702.150 480.750 ;
        RECT 716.850 480.750 718.050 484.050 ;
        RECT 716.850 479.700 720.600 480.750 ;
        RECT 674.400 471.600 676.200 474.600 ;
        RECT 688.200 471.600 690.000 478.800 ;
        RECT 698.400 477.600 699.600 479.700 ;
        RECT 697.800 471.600 699.600 477.600 ;
        RECT 700.800 476.700 708.600 478.050 ;
        RECT 700.800 471.600 702.600 476.700 ;
        RECT 706.800 471.600 708.600 476.700 ;
        RECT 710.400 476.700 718.200 478.050 ;
        RECT 710.400 471.600 712.200 476.700 ;
        RECT 716.400 471.600 718.200 476.700 ;
        RECT 719.400 477.600 720.600 479.700 ;
        RECT 722.550 480.450 723.450 490.950 ;
        RECT 729.000 490.350 731.400 491.400 ;
        RECT 743.700 491.550 746.100 492.900 ;
        RECT 725.100 486.150 726.900 487.950 ;
        RECT 724.950 484.050 727.050 486.150 ;
        RECT 729.000 483.150 730.050 490.350 ;
        RECT 731.100 486.150 732.900 487.950 ;
        RECT 730.950 484.050 733.050 486.150 ;
        RECT 733.950 484.950 736.050 487.050 ;
        RECT 743.700 484.950 745.050 491.550 ;
        RECT 751.800 491.400 753.600 503.400 ;
        RECT 758.400 497.400 760.200 503.400 ;
        RECT 727.950 481.050 730.050 483.150 ;
        RECT 724.950 480.450 727.050 481.050 ;
        RECT 722.550 479.550 727.050 480.450 ;
        RECT 724.950 478.950 727.050 479.550 ;
        RECT 719.400 471.600 721.200 477.600 ;
        RECT 729.000 474.600 730.050 481.050 ;
        RECT 730.950 480.450 733.050 481.050 ;
        RECT 734.550 480.450 735.450 484.950 ;
        RECT 730.950 479.550 735.450 480.450 ;
        RECT 742.950 482.850 745.050 484.950 ;
        RECT 746.400 490.200 748.200 490.650 ;
        RECT 752.400 490.200 753.600 491.400 ;
        RECT 746.400 489.000 753.600 490.200 ;
        RECT 746.400 488.850 748.200 489.000 ;
        RECT 730.950 478.950 733.050 479.550 ;
        RECT 742.950 477.600 744.000 482.850 ;
        RECT 746.400 480.600 747.300 488.850 ;
        RECT 749.100 486.150 750.900 487.950 ;
        RECT 755.100 486.150 756.900 487.950 ;
        RECT 748.950 484.050 751.050 486.150 ;
        RECT 752.100 483.150 753.900 484.950 ;
        RECT 754.950 484.050 757.050 486.150 ;
        RECT 751.950 481.050 754.050 483.150 ;
        RECT 746.250 479.700 748.050 480.600 ;
        RECT 758.550 480.300 759.600 497.400 ;
        RECT 765.000 491.400 766.800 503.400 ;
        RECT 760.950 485.850 763.050 487.950 ;
        RECT 765.000 486.150 766.050 491.400 ;
        RECT 761.100 484.050 762.900 485.850 ;
        RECT 763.950 484.050 766.050 486.150 ;
        RECT 746.250 478.800 749.700 479.700 ;
        RECT 728.400 471.600 730.200 474.600 ;
        RECT 742.800 471.600 744.600 477.600 ;
        RECT 748.800 474.600 749.700 478.800 ;
        RECT 755.400 479.100 762.900 480.300 ;
        RECT 748.800 471.600 750.600 474.600 ;
        RECT 755.400 471.600 757.200 479.100 ;
        RECT 761.100 478.500 762.900 479.100 ;
        RECT 765.000 477.600 766.050 484.050 ;
        RECT 762.900 476.100 766.050 477.600 ;
        RECT 762.900 471.600 764.700 476.100 ;
        RECT 4.800 464.400 6.600 467.400 ;
        RECT 5.400 456.150 6.600 464.400 ;
        RECT 13.800 461.400 15.600 467.400 ;
        RECT 14.400 459.300 15.600 461.400 ;
        RECT 16.800 462.300 18.600 467.400 ;
        RECT 22.800 462.300 24.600 467.400 ;
        RECT 16.800 460.950 24.600 462.300 ;
        RECT 26.400 459.900 28.200 467.400 ;
        RECT 33.900 462.900 35.700 467.400 ;
        RECT 33.900 461.400 37.050 462.900 ;
        RECT 32.100 459.900 33.900 460.500 ;
        RECT 14.400 458.250 18.150 459.300 ;
        RECT 26.400 458.700 33.900 459.900 ;
        RECT 4.950 454.050 7.050 456.150 ;
        RECT 7.950 455.850 10.050 457.950 ;
        RECT 8.100 454.050 9.900 455.850 ;
        RECT 16.950 454.950 18.150 458.250 ;
        RECT 20.100 456.150 21.900 457.950 ;
        RECT 5.400 441.600 6.600 454.050 ;
        RECT 16.950 452.850 19.050 454.950 ;
        RECT 19.950 454.050 22.050 456.150 ;
        RECT 22.950 452.850 25.050 454.950 ;
        RECT 25.950 452.850 28.050 454.950 ;
        RECT 13.950 449.850 16.050 451.950 ;
        RECT 14.250 448.050 16.050 449.850 ;
        RECT 17.850 447.600 19.050 452.850 ;
        RECT 23.100 451.050 24.900 452.850 ;
        RECT 26.100 451.050 27.900 452.850 ;
        RECT 4.800 435.600 6.600 441.600 ;
        RECT 17.700 435.600 19.500 447.600 ;
        RECT 29.550 441.600 30.600 458.700 ;
        RECT 36.000 454.950 37.050 461.400 ;
        RECT 50.100 459.000 51.900 467.400 ;
        RECT 32.100 453.150 33.900 454.950 ;
        RECT 31.950 451.050 34.050 453.150 ;
        RECT 34.950 452.850 37.050 454.950 ;
        RECT 47.700 457.350 51.900 459.000 ;
        RECT 62.400 464.400 64.200 467.400 ;
        RECT 70.800 464.400 72.600 467.400 ;
        RECT 47.700 453.150 48.600 457.350 ;
        RECT 58.950 455.850 61.050 457.950 ;
        RECT 62.400 456.150 63.600 464.400 ;
        RECT 71.400 456.150 72.600 464.400 ;
        RECT 86.100 459.000 87.900 467.400 ;
        RECT 101.400 464.400 103.200 467.400 ;
        RECT 59.100 454.050 60.900 455.850 ;
        RECT 61.950 454.050 64.050 456.150 ;
        RECT 70.950 454.050 73.050 456.150 ;
        RECT 73.950 455.850 76.050 457.950 ;
        RECT 86.100 457.350 90.300 459.000 ;
        RECT 74.100 454.050 75.900 455.850 ;
        RECT 36.000 447.600 37.050 452.850 ;
        RECT 46.950 451.050 49.050 453.150 ;
        RECT 29.400 435.600 31.200 441.600 ;
        RECT 36.000 435.600 37.800 447.600 ;
        RECT 47.700 442.800 48.600 451.050 ;
        RECT 49.950 449.850 52.050 451.950 ;
        RECT 55.950 449.850 58.050 451.950 ;
        RECT 49.950 448.050 51.750 449.850 ;
        RECT 52.950 446.850 55.050 448.950 ;
        RECT 56.100 448.050 57.900 449.850 ;
        RECT 53.100 445.050 54.900 446.850 ;
        RECT 47.700 441.900 54.300 442.800 ;
        RECT 47.700 441.600 48.600 441.900 ;
        RECT 46.800 435.600 48.600 441.600 ;
        RECT 52.800 441.600 54.300 441.900 ;
        RECT 62.400 441.600 63.600 454.050 ;
        RECT 71.400 441.600 72.600 454.050 ;
        RECT 89.400 453.150 90.300 457.350 ;
        RECT 97.950 455.850 100.050 457.950 ;
        RECT 101.400 456.150 102.600 464.400 ;
        RECT 111.000 460.200 112.800 467.400 ;
        RECT 111.000 459.300 114.600 460.200 ;
        RECT 98.100 454.050 99.900 455.850 ;
        RECT 100.950 454.050 103.050 456.150 ;
        RECT 79.950 449.850 82.050 451.950 ;
        RECT 85.950 449.850 88.050 451.950 ;
        RECT 88.950 451.050 91.050 453.150 ;
        RECT 80.100 448.050 81.900 449.850 ;
        RECT 82.950 446.850 85.050 448.950 ;
        RECT 86.250 448.050 88.050 449.850 ;
        RECT 83.100 445.050 84.900 446.850 ;
        RECT 89.400 442.800 90.300 451.050 ;
        RECT 83.700 441.900 90.300 442.800 ;
        RECT 83.700 441.600 85.200 441.900 ;
        RECT 52.800 435.600 54.600 441.600 ;
        RECT 62.400 435.600 64.200 441.600 ;
        RECT 70.800 435.600 72.600 441.600 ;
        RECT 83.400 435.600 85.200 441.600 ;
        RECT 89.400 441.600 90.300 441.900 ;
        RECT 101.400 441.600 102.600 454.050 ;
        RECT 110.100 453.150 111.900 454.950 ;
        RECT 109.950 451.050 112.050 453.150 ;
        RECT 113.400 451.950 114.600 459.300 ;
        RECT 125.100 459.000 126.900 467.400 ;
        RECT 140.400 464.400 142.200 467.400 ;
        RECT 125.100 457.350 129.300 459.000 ;
        RECT 116.100 453.150 117.900 454.950 ;
        RECT 128.400 453.150 129.300 457.350 ;
        RECT 136.950 455.850 139.050 457.950 ;
        RECT 140.400 456.150 141.600 464.400 ;
        RECT 146.400 462.300 148.200 467.400 ;
        RECT 152.400 462.300 154.200 467.400 ;
        RECT 146.400 460.950 154.200 462.300 ;
        RECT 155.400 461.400 157.200 467.400 ;
        RECT 155.400 459.300 156.600 461.400 ;
        RECT 152.850 458.250 156.600 459.300 ;
        RECT 170.100 459.000 171.900 467.400 ;
        RECT 184.800 464.400 186.600 467.400 ;
        RECT 194.400 464.400 196.200 467.400 ;
        RECT 149.100 456.150 150.900 457.950 ;
        RECT 137.100 454.050 138.900 455.850 ;
        RECT 139.950 454.050 142.050 456.150 ;
        RECT 112.950 449.850 115.050 451.950 ;
        RECT 115.950 451.050 118.050 453.150 ;
        RECT 118.950 449.850 121.050 451.950 ;
        RECT 124.950 449.850 127.050 451.950 ;
        RECT 127.950 451.050 130.050 453.150 ;
        RECT 113.400 441.600 114.600 449.850 ;
        RECT 119.100 448.050 120.900 449.850 ;
        RECT 121.950 446.850 124.050 448.950 ;
        RECT 125.250 448.050 127.050 449.850 ;
        RECT 122.100 445.050 123.900 446.850 ;
        RECT 128.400 442.800 129.300 451.050 ;
        RECT 122.700 441.900 129.300 442.800 ;
        RECT 122.700 441.600 124.200 441.900 ;
        RECT 89.400 435.600 91.200 441.600 ;
        RECT 101.400 435.600 103.200 441.600 ;
        RECT 112.800 435.600 114.600 441.600 ;
        RECT 122.400 435.600 124.200 441.600 ;
        RECT 128.400 441.600 129.300 441.900 ;
        RECT 140.400 441.600 141.600 454.050 ;
        RECT 145.950 452.850 148.050 454.950 ;
        RECT 148.950 454.050 151.050 456.150 ;
        RECT 152.850 454.950 154.050 458.250 ;
        RECT 170.100 457.350 174.300 459.000 ;
        RECT 151.950 452.850 154.050 454.950 ;
        RECT 173.400 453.150 174.300 457.350 ;
        RECT 184.950 457.950 186.000 464.400 ;
        RECT 195.000 457.950 196.050 464.400 ;
        RECT 211.200 460.200 213.000 467.400 ;
        RECT 221.400 464.400 223.200 467.400 ;
        RECT 233.400 464.400 235.200 467.400 ;
        RECT 184.950 455.850 187.050 457.950 ;
        RECT 193.950 455.850 196.050 457.950 ;
        RECT 146.100 451.050 147.900 452.850 ;
        RECT 151.950 447.600 153.150 452.850 ;
        RECT 154.950 449.850 157.050 451.950 ;
        RECT 163.950 449.850 166.050 451.950 ;
        RECT 169.950 449.850 172.050 451.950 ;
        RECT 172.950 451.050 175.050 453.150 ;
        RECT 181.950 452.850 184.050 454.950 ;
        RECT 182.100 451.050 183.900 452.850 ;
        RECT 154.950 448.050 156.750 449.850 ;
        RECT 164.100 448.050 165.900 449.850 ;
        RECT 128.400 435.600 130.200 441.600 ;
        RECT 140.400 435.600 142.200 441.600 ;
        RECT 151.500 435.600 153.300 447.600 ;
        RECT 166.950 446.850 169.050 448.950 ;
        RECT 170.250 448.050 172.050 449.850 ;
        RECT 167.100 445.050 168.900 446.850 ;
        RECT 173.400 442.800 174.300 451.050 ;
        RECT 184.950 448.650 186.000 455.850 ;
        RECT 187.950 452.850 190.050 454.950 ;
        RECT 190.950 452.850 193.050 454.950 ;
        RECT 188.100 451.050 189.900 452.850 ;
        RECT 191.100 451.050 192.900 452.850 ;
        RECT 167.700 441.900 174.300 442.800 ;
        RECT 167.700 441.600 169.200 441.900 ;
        RECT 167.400 435.600 169.200 441.600 ;
        RECT 173.400 441.600 174.300 441.900 ;
        RECT 183.600 447.600 186.000 448.650 ;
        RECT 195.000 448.650 196.050 455.850 ;
        RECT 209.400 459.300 213.000 460.200 ;
        RECT 196.950 452.850 199.050 454.950 ;
        RECT 206.100 453.150 207.900 454.950 ;
        RECT 197.100 451.050 198.900 452.850 ;
        RECT 205.950 451.050 208.050 453.150 ;
        RECT 209.400 451.950 210.600 459.300 ;
        RECT 222.000 457.950 223.050 464.400 ;
        RECT 234.000 457.950 235.050 464.400 ;
        RECT 242.400 459.900 244.200 467.400 ;
        RECT 249.900 462.900 251.700 467.400 ;
        RECT 262.800 464.400 264.600 467.400 ;
        RECT 275.400 464.400 277.200 467.400 ;
        RECT 290.400 464.400 292.200 467.400 ;
        RECT 249.900 461.400 253.050 462.900 ;
        RECT 248.100 459.900 249.900 460.500 ;
        RECT 242.400 458.700 249.900 459.900 ;
        RECT 220.950 455.850 223.050 457.950 ;
        RECT 232.950 455.850 235.050 457.950 ;
        RECT 212.100 453.150 213.900 454.950 ;
        RECT 208.950 449.850 211.050 451.950 ;
        RECT 211.950 451.050 214.050 453.150 ;
        RECT 217.950 452.850 220.050 454.950 ;
        RECT 218.100 451.050 219.900 452.850 ;
        RECT 195.000 447.600 197.400 448.650 ;
        RECT 173.400 435.600 175.200 441.600 ;
        RECT 183.600 435.600 185.400 447.600 ;
        RECT 195.600 435.600 197.400 447.600 ;
        RECT 209.400 441.600 210.600 449.850 ;
        RECT 222.000 448.650 223.050 455.850 ;
        RECT 223.950 452.850 226.050 454.950 ;
        RECT 229.950 452.850 232.050 454.950 ;
        RECT 224.100 451.050 225.900 452.850 ;
        RECT 230.100 451.050 231.900 452.850 ;
        RECT 234.000 448.650 235.050 455.850 ;
        RECT 235.950 452.850 238.050 454.950 ;
        RECT 241.950 452.850 244.050 454.950 ;
        RECT 236.100 451.050 237.900 452.850 ;
        RECT 242.100 451.050 243.900 452.850 ;
        RECT 222.000 447.600 224.400 448.650 ;
        RECT 234.000 447.600 236.400 448.650 ;
        RECT 209.400 435.600 211.200 441.600 ;
        RECT 222.600 435.600 224.400 447.600 ;
        RECT 234.600 435.600 236.400 447.600 ;
        RECT 245.550 441.600 246.600 458.700 ;
        RECT 252.000 454.950 253.050 461.400 ;
        RECT 262.950 457.950 264.000 464.400 ;
        RECT 276.000 457.950 277.050 464.400 ;
        RECT 262.950 455.850 265.050 457.950 ;
        RECT 274.950 455.850 277.050 457.950 ;
        RECT 286.950 455.850 289.050 457.950 ;
        RECT 290.400 456.150 291.600 464.400 ;
        RECT 301.200 460.200 303.000 467.400 ;
        RECT 299.400 459.300 303.000 460.200 ;
        RECT 311.400 464.400 313.200 467.400 ;
        RECT 248.100 453.150 249.900 454.950 ;
        RECT 247.950 451.050 250.050 453.150 ;
        RECT 250.950 452.850 253.050 454.950 ;
        RECT 259.950 452.850 262.050 454.950 ;
        RECT 252.000 447.600 253.050 452.850 ;
        RECT 260.100 451.050 261.900 452.850 ;
        RECT 262.950 448.650 264.000 455.850 ;
        RECT 265.950 452.850 268.050 454.950 ;
        RECT 271.950 452.850 274.050 454.950 ;
        RECT 266.100 451.050 267.900 452.850 ;
        RECT 272.100 451.050 273.900 452.850 ;
        RECT 261.600 447.600 264.000 448.650 ;
        RECT 276.000 448.650 277.050 455.850 ;
        RECT 277.950 452.850 280.050 454.950 ;
        RECT 287.100 454.050 288.900 455.850 ;
        RECT 289.950 454.050 292.050 456.150 ;
        RECT 278.100 451.050 279.900 452.850 ;
        RECT 276.000 447.600 278.400 448.650 ;
        RECT 245.400 435.600 247.200 441.600 ;
        RECT 252.000 435.600 253.800 447.600 ;
        RECT 261.600 435.600 263.400 447.600 ;
        RECT 276.600 435.600 278.400 447.600 ;
        RECT 290.400 441.600 291.600 454.050 ;
        RECT 296.100 453.150 297.900 454.950 ;
        RECT 295.950 451.050 298.050 453.150 ;
        RECT 299.400 451.950 300.600 459.300 ;
        RECT 307.950 455.850 310.050 457.950 ;
        RECT 311.400 456.150 312.600 464.400 ;
        RECT 322.200 461.400 324.000 467.400 ;
        RECT 340.200 463.050 342.000 467.400 ;
        RECT 357.000 463.050 358.800 467.400 ;
        RECT 340.200 461.400 345.600 463.050 ;
        RECT 320.250 456.150 322.050 457.950 ;
        RECT 302.100 453.150 303.900 454.950 ;
        RECT 308.100 454.050 309.900 455.850 ;
        RECT 310.950 454.050 313.050 456.150 ;
        RECT 298.950 449.850 301.050 451.950 ;
        RECT 301.950 451.050 304.050 453.150 ;
        RECT 299.400 441.600 300.600 449.850 ;
        RECT 311.400 441.600 312.600 454.050 ;
        RECT 316.950 452.850 319.050 454.950 ;
        RECT 319.950 454.050 322.050 456.150 ;
        RECT 322.950 454.950 324.000 461.400 ;
        RECT 325.950 456.150 327.750 457.950 ;
        RECT 335.100 456.150 336.900 457.950 ;
        RECT 322.950 452.850 325.050 454.950 ;
        RECT 325.950 454.050 328.050 456.150 ;
        RECT 328.950 452.850 331.050 454.950 ;
        RECT 334.950 454.050 337.050 456.150 ;
        RECT 337.950 455.850 340.050 457.950 ;
        RECT 341.100 456.150 342.900 457.950 ;
        RECT 338.100 454.050 339.900 455.850 ;
        RECT 340.950 454.050 343.050 456.150 ;
        RECT 344.700 454.950 345.600 461.400 ;
        RECT 353.400 461.400 358.800 463.050 ;
        RECT 365.550 461.400 367.350 467.400 ;
        RECT 373.650 464.400 375.450 467.400 ;
        RECT 381.450 464.400 383.250 467.400 ;
        RECT 389.250 465.300 391.050 467.400 ;
        RECT 389.250 464.400 393.000 465.300 ;
        RECT 373.650 463.500 374.700 464.400 ;
        RECT 370.950 462.300 374.700 463.500 ;
        RECT 382.200 462.600 383.250 464.400 ;
        RECT 391.950 463.500 393.000 464.400 ;
        RECT 370.950 461.400 373.050 462.300 ;
        RECT 353.400 454.950 354.300 461.400 ;
        RECT 365.550 459.150 366.750 461.400 ;
        RECT 378.150 460.200 379.950 462.000 ;
        RECT 382.200 461.550 387.150 462.600 ;
        RECT 385.350 460.800 387.150 461.550 ;
        RECT 388.650 460.800 390.450 462.600 ;
        RECT 391.950 461.400 394.050 463.500 ;
        RECT 397.050 461.400 398.850 467.400 ;
        RECT 411.000 463.050 412.800 467.400 ;
        RECT 379.050 459.900 379.950 460.200 ;
        RECT 389.100 459.900 390.150 460.800 ;
        RECT 356.100 456.150 357.900 457.950 ;
        RECT 343.950 452.850 346.050 454.950 ;
        RECT 352.950 452.850 355.050 454.950 ;
        RECT 355.950 454.050 358.050 456.150 ;
        RECT 358.950 455.850 361.050 457.950 ;
        RECT 362.100 456.150 363.900 457.950 ;
        RECT 365.550 457.050 370.050 459.150 ;
        RECT 379.050 459.000 390.150 459.900 ;
        RECT 359.100 454.050 360.900 455.850 ;
        RECT 361.950 454.050 364.050 456.150 ;
        RECT 317.250 451.050 319.050 452.850 ;
        RECT 324.150 449.400 325.050 452.850 ;
        RECT 329.100 451.050 330.900 452.850 ;
        RECT 324.150 448.500 328.200 449.400 ;
        RECT 317.400 446.400 325.200 447.300 ;
        RECT 290.400 435.600 292.200 441.600 ;
        RECT 299.400 435.600 301.200 441.600 ;
        RECT 311.400 435.600 313.200 441.600 ;
        RECT 317.400 435.600 319.200 446.400 ;
        RECT 323.400 436.500 325.200 446.400 ;
        RECT 326.400 437.400 328.200 448.500 ;
        RECT 344.700 447.600 345.600 452.850 ;
        RECT 353.400 447.600 354.300 452.850 ;
        RECT 365.550 447.600 366.750 457.050 ;
        RECT 367.950 455.250 371.850 457.050 ;
        RECT 367.950 454.950 370.050 455.250 ;
        RECT 379.050 454.950 379.950 459.000 ;
        RECT 389.100 457.800 390.150 459.000 ;
        RECT 389.100 456.600 396.000 457.800 ;
        RECT 389.100 456.000 390.900 456.600 ;
        RECT 395.100 455.850 396.000 456.600 ;
        RECT 392.100 454.950 393.900 455.700 ;
        RECT 379.050 452.850 382.050 454.950 ;
        RECT 385.950 453.900 393.900 454.950 ;
        RECT 395.100 454.050 396.900 455.850 ;
        RECT 385.950 452.850 388.050 453.900 ;
        RECT 367.950 449.400 369.750 451.200 ;
        RECT 368.850 448.200 373.050 449.400 ;
        RECT 379.050 448.200 379.950 452.850 ;
        RECT 387.750 449.100 389.550 449.400 ;
        RECT 329.400 436.500 331.200 447.600 ;
        RECT 323.400 435.600 331.200 436.500 ;
        RECT 335.400 446.700 343.200 447.600 ;
        RECT 335.400 435.600 337.200 446.700 ;
        RECT 341.400 435.600 343.200 446.700 ;
        RECT 344.400 435.600 346.200 447.600 ;
        RECT 352.800 435.600 354.600 447.600 ;
        RECT 355.800 446.700 363.600 447.600 ;
        RECT 355.800 435.600 357.600 446.700 ;
        RECT 361.800 435.600 363.600 446.700 ;
        RECT 365.550 435.600 367.350 447.600 ;
        RECT 370.950 447.300 373.050 448.200 ;
        RECT 373.950 447.300 379.950 448.200 ;
        RECT 381.150 448.800 389.550 449.100 ;
        RECT 397.950 448.800 398.850 461.400 ;
        RECT 407.400 461.400 412.800 463.050 ;
        RECT 419.400 462.300 421.200 467.400 ;
        RECT 425.400 462.300 427.200 467.400 ;
        RECT 407.400 454.950 408.300 461.400 ;
        RECT 419.400 460.950 427.200 462.300 ;
        RECT 428.400 461.400 430.200 467.400 ;
        RECT 428.400 459.300 429.600 461.400 ;
        RECT 439.800 460.500 441.600 467.400 ;
        RECT 445.800 460.500 447.600 467.400 ;
        RECT 451.800 460.500 453.600 467.400 ;
        RECT 457.800 460.500 459.600 467.400 ;
        RECT 425.850 458.250 429.600 459.300 ;
        RECT 438.900 459.300 441.600 460.500 ;
        RECT 443.700 459.300 447.600 460.500 ;
        RECT 449.700 459.300 453.600 460.500 ;
        RECT 455.700 459.300 459.600 460.500 ;
        RECT 471.000 460.200 472.800 467.400 ;
        RECT 483.000 460.200 484.800 467.400 ;
        RECT 495.000 460.200 496.800 467.400 ;
        RECT 471.000 459.300 474.600 460.200 ;
        RECT 483.000 459.300 486.600 460.200 ;
        RECT 495.000 459.300 498.600 460.200 ;
        RECT 410.100 456.150 411.900 457.950 ;
        RECT 406.950 452.850 409.050 454.950 ;
        RECT 409.950 454.050 412.050 456.150 ;
        RECT 412.950 455.850 415.050 457.950 ;
        RECT 416.100 456.150 417.900 457.950 ;
        RECT 422.100 456.150 423.900 457.950 ;
        RECT 413.100 454.050 414.900 455.850 ;
        RECT 415.950 454.050 418.050 456.150 ;
        RECT 418.950 452.850 421.050 454.950 ;
        RECT 421.950 454.050 424.050 456.150 ;
        RECT 425.850 454.950 427.050 458.250 ;
        RECT 438.900 456.150 439.800 459.300 ;
        RECT 443.700 458.400 444.900 459.300 ;
        RECT 449.700 458.400 450.900 459.300 ;
        RECT 455.700 458.400 456.900 459.300 ;
        RECT 440.700 457.200 444.900 458.400 ;
        RECT 440.700 456.600 442.500 457.200 ;
        RECT 424.950 452.850 427.050 454.950 ;
        RECT 436.950 454.050 439.800 456.150 ;
        RECT 381.150 448.200 398.850 448.800 ;
        RECT 373.950 446.400 374.850 447.300 ;
        RECT 372.150 444.600 374.850 446.400 ;
        RECT 375.750 446.100 377.550 446.400 ;
        RECT 381.150 446.100 382.050 448.200 ;
        RECT 387.750 447.600 398.850 448.200 ;
        RECT 407.400 447.600 408.300 452.850 ;
        RECT 419.100 451.050 420.900 452.850 ;
        RECT 424.950 447.600 426.150 452.850 ;
        RECT 427.950 449.850 430.050 451.950 ;
        RECT 427.950 448.050 429.750 449.850 ;
        RECT 438.900 449.700 439.800 454.050 ;
        RECT 443.700 449.700 444.900 457.200 ;
        RECT 446.700 457.200 450.900 458.400 ;
        RECT 446.700 456.600 448.500 457.200 ;
        RECT 449.700 449.700 450.900 457.200 ;
        RECT 452.700 457.200 456.900 458.400 ;
        RECT 452.700 456.600 454.500 457.200 ;
        RECT 455.700 449.700 456.900 457.200 ;
        RECT 458.100 456.150 459.900 457.950 ;
        RECT 457.950 454.050 460.050 456.150 ;
        RECT 470.100 453.150 471.900 454.950 ;
        RECT 469.950 451.050 472.050 453.150 ;
        RECT 473.400 451.950 474.600 459.300 ;
        RECT 476.100 453.150 477.900 454.950 ;
        RECT 482.100 453.150 483.900 454.950 ;
        RECT 472.950 449.850 475.050 451.950 ;
        RECT 475.950 451.050 478.050 453.150 ;
        RECT 481.950 451.050 484.050 453.150 ;
        RECT 485.400 451.950 486.600 459.300 ;
        RECT 488.100 453.150 489.900 454.950 ;
        RECT 494.100 453.150 495.900 454.950 ;
        RECT 484.950 449.850 487.050 451.950 ;
        RECT 487.950 451.050 490.050 453.150 ;
        RECT 493.950 451.050 496.050 453.150 ;
        RECT 497.400 451.950 498.600 459.300 ;
        RECT 509.100 459.000 510.900 467.400 ;
        RECT 524.100 459.000 525.900 467.400 ;
        RECT 538.800 464.400 540.600 467.400 ;
        RECT 509.100 457.350 513.300 459.000 ;
        RECT 500.100 453.150 501.900 454.950 ;
        RECT 512.400 453.150 513.300 457.350 ;
        RECT 521.700 457.350 525.900 459.000 ;
        RECT 521.700 453.150 522.600 457.350 ;
        RECT 539.400 456.150 540.600 464.400 ;
        RECT 550.800 461.400 552.600 467.400 ;
        RECT 551.400 459.300 552.600 461.400 ;
        RECT 553.800 462.300 555.600 467.400 ;
        RECT 559.800 462.300 561.600 467.400 ;
        RECT 553.800 460.950 561.600 462.300 ;
        RECT 566.400 464.400 568.200 467.400 ;
        RECT 551.400 458.250 555.150 459.300 ;
        RECT 538.950 454.050 541.050 456.150 ;
        RECT 541.950 455.850 544.050 457.950 ;
        RECT 544.950 456.450 547.050 457.050 ;
        RECT 550.950 456.450 553.050 457.050 ;
        RECT 542.100 454.050 543.900 455.850 ;
        RECT 544.950 455.550 553.050 456.450 ;
        RECT 544.950 454.950 547.050 455.550 ;
        RECT 550.950 454.950 553.050 455.550 ;
        RECT 553.950 454.950 555.150 458.250 ;
        RECT 557.100 456.150 558.900 457.950 ;
        RECT 496.950 449.850 499.050 451.950 ;
        RECT 499.950 451.050 502.050 453.150 ;
        RECT 502.950 449.850 505.050 451.950 ;
        RECT 508.950 449.850 511.050 451.950 ;
        RECT 511.950 451.050 514.050 453.150 ;
        RECT 520.950 451.050 523.050 453.150 ;
        RECT 438.900 448.500 441.600 449.700 ;
        RECT 443.700 448.500 447.600 449.700 ;
        RECT 449.700 448.500 453.600 449.700 ;
        RECT 455.700 448.500 459.600 449.700 ;
        RECT 375.750 445.200 382.050 446.100 ;
        RECT 382.950 446.700 384.750 447.300 ;
        RECT 382.950 445.500 390.450 446.700 ;
        RECT 375.750 444.600 377.550 445.200 ;
        RECT 389.250 444.600 390.450 445.500 ;
        RECT 370.950 441.600 374.850 443.700 ;
        RECT 379.950 443.550 381.750 444.300 ;
        RECT 384.750 443.550 386.550 444.300 ;
        RECT 379.950 442.500 386.550 443.550 ;
        RECT 389.250 442.500 394.050 444.600 ;
        RECT 373.050 435.600 374.850 441.600 ;
        RECT 380.850 435.600 382.650 442.500 ;
        RECT 389.250 441.600 390.450 442.500 ;
        RECT 388.650 435.600 390.450 441.600 ;
        RECT 397.050 435.600 398.850 447.600 ;
        RECT 406.800 435.600 408.600 447.600 ;
        RECT 409.800 446.700 417.600 447.600 ;
        RECT 409.800 435.600 411.600 446.700 ;
        RECT 415.800 435.600 417.600 446.700 ;
        RECT 424.500 435.600 426.300 447.600 ;
        RECT 439.800 435.600 441.600 448.500 ;
        RECT 445.800 435.600 447.600 448.500 ;
        RECT 451.800 435.600 453.600 448.500 ;
        RECT 457.800 435.600 459.600 448.500 ;
        RECT 473.400 441.600 474.600 449.850 ;
        RECT 485.400 441.600 486.600 449.850 ;
        RECT 497.400 441.600 498.600 449.850 ;
        RECT 503.100 448.050 504.900 449.850 ;
        RECT 505.950 446.850 508.050 448.950 ;
        RECT 509.250 448.050 511.050 449.850 ;
        RECT 506.100 445.050 507.900 446.850 ;
        RECT 512.400 442.800 513.300 451.050 ;
        RECT 506.700 441.900 513.300 442.800 ;
        RECT 506.700 441.600 508.200 441.900 ;
        RECT 472.800 435.600 474.600 441.600 ;
        RECT 484.800 435.600 486.600 441.600 ;
        RECT 496.800 435.600 498.600 441.600 ;
        RECT 506.400 435.600 508.200 441.600 ;
        RECT 512.400 441.600 513.300 441.900 ;
        RECT 521.700 442.800 522.600 451.050 ;
        RECT 523.950 449.850 526.050 451.950 ;
        RECT 529.950 449.850 532.050 451.950 ;
        RECT 523.950 448.050 525.750 449.850 ;
        RECT 526.950 446.850 529.050 448.950 ;
        RECT 530.100 448.050 531.900 449.850 ;
        RECT 527.100 445.050 528.900 446.850 ;
        RECT 521.700 441.900 528.300 442.800 ;
        RECT 521.700 441.600 522.600 441.900 ;
        RECT 512.400 435.600 514.200 441.600 ;
        RECT 520.800 435.600 522.600 441.600 ;
        RECT 526.800 441.600 528.300 441.900 ;
        RECT 539.400 441.600 540.600 454.050 ;
        RECT 553.950 452.850 556.050 454.950 ;
        RECT 556.950 454.050 559.050 456.150 ;
        RECT 562.950 455.850 565.050 457.950 ;
        RECT 566.400 456.150 567.600 464.400 ;
        RECT 572.400 462.300 574.200 467.400 ;
        RECT 578.400 462.300 580.200 467.400 ;
        RECT 572.400 460.950 580.200 462.300 ;
        RECT 581.400 461.400 583.200 467.400 ;
        RECT 581.400 459.300 582.600 461.400 ;
        RECT 578.850 458.250 582.600 459.300 ;
        RECT 596.100 459.000 597.900 467.400 ;
        RECT 612.000 463.050 613.800 467.400 ;
        RECT 575.100 456.150 576.900 457.950 ;
        RECT 559.950 452.850 562.050 454.950 ;
        RECT 563.100 454.050 564.900 455.850 ;
        RECT 565.950 454.050 568.050 456.150 ;
        RECT 550.950 449.850 553.050 451.950 ;
        RECT 551.250 448.050 553.050 449.850 ;
        RECT 554.850 447.600 556.050 452.850 ;
        RECT 560.100 451.050 561.900 452.850 ;
        RECT 526.800 435.600 528.600 441.600 ;
        RECT 538.800 435.600 540.600 441.600 ;
        RECT 554.700 435.600 556.500 447.600 ;
        RECT 566.400 441.600 567.600 454.050 ;
        RECT 571.950 452.850 574.050 454.950 ;
        RECT 574.950 454.050 577.050 456.150 ;
        RECT 578.850 454.950 580.050 458.250 ;
        RECT 577.950 452.850 580.050 454.950 ;
        RECT 593.700 457.350 597.900 459.000 ;
        RECT 608.400 461.400 613.800 463.050 ;
        RECT 630.000 461.400 631.800 467.400 ;
        RECT 593.700 453.150 594.600 457.350 ;
        RECT 608.400 454.950 609.300 461.400 ;
        RECT 611.100 456.150 612.900 457.950 ;
        RECT 572.100 451.050 573.900 452.850 ;
        RECT 577.950 447.600 579.150 452.850 ;
        RECT 580.950 449.850 583.050 451.950 ;
        RECT 592.950 451.050 595.050 453.150 ;
        RECT 607.950 452.850 610.050 454.950 ;
        RECT 610.950 454.050 613.050 456.150 ;
        RECT 613.950 455.850 616.050 457.950 ;
        RECT 617.100 456.150 618.900 457.950 ;
        RECT 626.250 456.150 628.050 457.950 ;
        RECT 614.100 454.050 615.900 455.850 ;
        RECT 616.950 454.050 619.050 456.150 ;
        RECT 622.950 452.850 625.050 454.950 ;
        RECT 625.950 454.050 628.050 456.150 ;
        RECT 630.000 454.950 631.050 461.400 ;
        RECT 642.000 460.200 643.800 467.400 ;
        RECT 653.400 464.400 655.200 467.400 ;
        RECT 642.000 459.300 645.600 460.200 ;
        RECT 628.950 452.850 631.050 454.950 ;
        RECT 631.950 456.150 633.750 457.950 ;
        RECT 631.950 454.050 634.050 456.150 ;
        RECT 634.950 452.850 637.050 454.950 ;
        RECT 641.100 453.150 642.900 454.950 ;
        RECT 580.950 448.050 582.750 449.850 ;
        RECT 566.400 435.600 568.200 441.600 ;
        RECT 577.500 435.600 579.300 447.600 ;
        RECT 593.700 442.800 594.600 451.050 ;
        RECT 595.950 449.850 598.050 451.950 ;
        RECT 601.950 449.850 604.050 451.950 ;
        RECT 595.950 448.050 597.750 449.850 ;
        RECT 598.950 446.850 601.050 448.950 ;
        RECT 602.100 448.050 603.900 449.850 ;
        RECT 608.400 447.600 609.300 452.850 ;
        RECT 623.100 451.050 624.900 452.850 ;
        RECT 628.950 449.400 629.850 452.850 ;
        RECT 634.950 451.050 636.750 452.850 ;
        RECT 640.950 451.050 643.050 453.150 ;
        RECT 644.400 451.950 645.600 459.300 ;
        RECT 649.950 455.850 652.050 457.950 ;
        RECT 653.400 456.150 654.600 464.400 ;
        RECT 659.400 462.300 661.200 467.400 ;
        RECT 665.400 462.300 667.200 467.400 ;
        RECT 659.400 460.950 667.200 462.300 ;
        RECT 668.400 461.400 670.200 467.400 ;
        RECT 676.950 462.450 679.050 463.050 ;
        RECT 674.550 461.550 679.050 462.450 ;
        RECT 668.400 459.300 669.600 461.400 ;
        RECT 665.850 458.250 669.600 459.300 ;
        RECT 662.100 456.150 663.900 457.950 ;
        RECT 647.100 453.150 648.900 454.950 ;
        RECT 650.100 454.050 651.900 455.850 ;
        RECT 652.950 454.050 655.050 456.150 ;
        RECT 643.950 449.850 646.050 451.950 ;
        RECT 646.950 451.050 649.050 453.150 ;
        RECT 625.800 448.500 629.850 449.400 ;
        RECT 599.100 445.050 600.900 446.850 ;
        RECT 593.700 441.900 600.300 442.800 ;
        RECT 593.700 441.600 594.600 441.900 ;
        RECT 592.800 435.600 594.600 441.600 ;
        RECT 598.800 441.600 600.300 441.900 ;
        RECT 598.800 435.600 600.600 441.600 ;
        RECT 607.800 435.600 609.600 447.600 ;
        RECT 610.800 446.700 618.600 447.600 ;
        RECT 610.800 435.600 612.600 446.700 ;
        RECT 616.800 435.600 618.600 446.700 ;
        RECT 622.800 436.500 624.600 447.600 ;
        RECT 625.800 437.400 627.600 448.500 ;
        RECT 628.800 446.400 636.600 447.300 ;
        RECT 628.800 436.500 630.600 446.400 ;
        RECT 622.800 435.600 630.600 436.500 ;
        RECT 634.800 435.600 636.600 446.400 ;
        RECT 644.400 441.600 645.600 449.850 ;
        RECT 643.800 435.600 645.600 441.600 ;
        RECT 653.400 441.600 654.600 454.050 ;
        RECT 658.950 452.850 661.050 454.950 ;
        RECT 661.950 454.050 664.050 456.150 ;
        RECT 665.850 454.950 667.050 458.250 ;
        RECT 664.950 452.850 667.050 454.950 ;
        RECT 659.100 451.050 660.900 452.850 ;
        RECT 664.950 447.600 666.150 452.850 ;
        RECT 667.950 449.850 670.050 451.950 ;
        RECT 667.950 448.050 669.750 449.850 ;
        RECT 674.550 448.050 675.450 461.550 ;
        RECT 676.950 460.950 679.050 461.550 ;
        RECT 680.100 459.000 681.900 467.400 ;
        RECT 694.800 464.400 696.600 467.400 ;
        RECT 677.700 457.350 681.900 459.000 ;
        RECT 677.700 453.150 678.600 457.350 ;
        RECT 695.400 456.150 696.600 464.400 ;
        RECT 706.200 463.050 708.000 467.400 ;
        RECT 722.400 464.400 724.200 467.400 ;
        RECT 737.400 464.400 739.200 467.400 ;
        RECT 706.200 461.400 711.600 463.050 ;
        RECT 694.950 454.050 697.050 456.150 ;
        RECT 697.950 455.850 700.050 457.950 ;
        RECT 701.100 456.150 702.900 457.950 ;
        RECT 698.100 454.050 699.900 455.850 ;
        RECT 700.950 454.050 703.050 456.150 ;
        RECT 703.950 455.850 706.050 457.950 ;
        RECT 707.100 456.150 708.900 457.950 ;
        RECT 704.100 454.050 705.900 455.850 ;
        RECT 706.950 454.050 709.050 456.150 ;
        RECT 710.700 454.950 711.600 461.400 ;
        RECT 723.000 457.950 724.050 464.400 ;
        RECT 738.300 460.200 739.200 464.400 ;
        RECT 743.400 461.400 745.200 467.400 ;
        RECT 749.400 462.300 751.200 467.400 ;
        RECT 755.400 462.300 757.200 467.400 ;
        RECT 730.950 457.950 733.050 460.050 ;
        RECT 738.300 459.300 741.750 460.200 ;
        RECT 739.950 458.400 741.750 459.300 ;
        RECT 721.950 455.850 724.050 457.950 ;
        RECT 691.950 453.450 694.050 454.050 ;
        RECT 676.950 451.050 679.050 453.150 ;
        RECT 689.550 452.550 694.050 453.450 ;
        RECT 653.400 435.600 655.200 441.600 ;
        RECT 664.500 435.600 666.300 447.600 ;
        RECT 673.950 445.950 676.050 448.050 ;
        RECT 677.700 442.800 678.600 451.050 ;
        RECT 679.950 449.850 682.050 451.950 ;
        RECT 685.950 449.850 688.050 451.950 ;
        RECT 679.950 448.050 681.750 449.850 ;
        RECT 682.950 446.850 685.050 448.950 ;
        RECT 686.100 448.050 687.900 449.850 ;
        RECT 683.100 445.050 684.900 446.850 ;
        RECT 685.950 444.450 688.050 445.050 ;
        RECT 689.550 444.450 690.450 452.550 ;
        RECT 691.950 451.950 694.050 452.550 ;
        RECT 685.950 443.550 690.450 444.450 ;
        RECT 685.950 442.950 688.050 443.550 ;
        RECT 677.700 441.900 684.300 442.800 ;
        RECT 677.700 441.600 678.600 441.900 ;
        RECT 676.800 435.600 678.600 441.600 ;
        RECT 682.800 441.600 684.300 441.900 ;
        RECT 695.400 441.600 696.600 454.050 ;
        RECT 709.950 452.850 712.050 454.950 ;
        RECT 718.950 452.850 721.050 454.950 ;
        RECT 710.700 447.600 711.600 452.850 ;
        RECT 719.100 451.050 720.900 452.850 ;
        RECT 723.000 448.650 724.050 455.850 ;
        RECT 724.950 452.850 727.050 454.950 ;
        RECT 725.100 451.050 726.900 452.850 ;
        RECT 723.000 447.600 725.400 448.650 ;
        RECT 682.800 435.600 684.600 441.600 ;
        RECT 694.800 435.600 696.600 441.600 ;
        RECT 701.400 446.700 709.200 447.600 ;
        RECT 701.400 435.600 703.200 446.700 ;
        RECT 707.400 435.600 709.200 446.700 ;
        RECT 710.400 435.600 712.200 447.600 ;
        RECT 723.600 435.600 725.400 447.600 ;
        RECT 727.950 447.450 730.050 448.050 ;
        RECT 731.550 447.450 732.450 457.950 ;
        RECT 733.950 455.850 736.050 457.950 ;
        RECT 734.100 454.050 735.900 455.850 ;
        RECT 736.950 452.850 739.050 454.950 ;
        RECT 737.100 451.050 738.900 452.850 ;
        RECT 740.700 450.150 741.600 458.400 ;
        RECT 744.000 456.150 745.050 461.400 ;
        RECT 749.400 460.950 757.200 462.300 ;
        RECT 758.400 461.400 760.200 467.400 ;
        RECT 758.400 459.300 759.600 461.400 ;
        RECT 755.850 458.250 759.600 459.300 ;
        RECT 752.100 456.150 753.900 457.950 ;
        RECT 739.800 450.000 741.600 450.150 ;
        RECT 727.950 446.550 732.450 447.450 ;
        RECT 734.400 448.800 741.600 450.000 ;
        RECT 734.400 447.600 735.600 448.800 ;
        RECT 739.800 448.350 741.600 448.800 ;
        RECT 742.950 454.050 745.050 456.150 ;
        RECT 727.950 445.950 730.050 446.550 ;
        RECT 734.400 435.600 736.200 447.600 ;
        RECT 742.950 447.450 744.300 454.050 ;
        RECT 748.950 452.850 751.050 454.950 ;
        RECT 751.950 454.050 754.050 456.150 ;
        RECT 755.850 454.950 757.050 458.250 ;
        RECT 754.950 452.850 757.050 454.950 ;
        RECT 749.100 451.050 750.900 452.850 ;
        RECT 754.950 447.600 756.150 452.850 ;
        RECT 757.950 449.850 760.050 451.950 ;
        RECT 757.950 448.050 759.750 449.850 ;
        RECT 741.900 446.100 744.300 447.450 ;
        RECT 741.900 435.600 743.700 446.100 ;
        RECT 754.500 435.600 756.300 447.600 ;
        RECT 4.800 425.400 6.600 431.400 ;
        RECT 5.400 412.950 6.600 425.400 ;
        RECT 17.700 419.400 19.500 431.400 ;
        RECT 34.500 419.400 36.300 431.400 ;
        RECT 52.800 425.400 54.600 431.400 ;
        RECT 61.800 425.400 63.600 431.400 ;
        RECT 14.250 417.150 16.050 418.950 ;
        RECT 13.950 415.050 16.050 417.150 ;
        RECT 17.850 414.150 19.050 419.400 ;
        RECT 23.100 414.150 24.900 415.950 ;
        RECT 29.100 414.150 30.900 415.950 ;
        RECT 34.950 414.150 36.150 419.400 ;
        RECT 37.950 417.150 39.750 418.950 ;
        RECT 53.400 417.150 54.600 425.400 ;
        RECT 62.700 425.100 63.600 425.400 ;
        RECT 67.800 425.400 69.600 431.400 ;
        RECT 77.400 425.400 79.200 431.400 ;
        RECT 67.800 425.100 69.300 425.400 ;
        RECT 62.700 424.200 69.300 425.100 ;
        RECT 77.700 425.100 79.200 425.400 ;
        RECT 83.400 425.400 85.200 431.400 ;
        RECT 94.800 425.400 96.600 431.400 ;
        RECT 104.400 425.400 106.200 431.400 ;
        RECT 83.400 425.100 84.300 425.400 ;
        RECT 77.700 424.200 84.300 425.100 ;
        RECT 37.950 415.050 40.050 417.150 ;
        RECT 4.950 410.850 7.050 412.950 ;
        RECT 8.100 411.150 9.900 412.950 ;
        RECT 16.950 412.050 19.050 414.150 ;
        RECT 5.400 402.600 6.600 410.850 ;
        RECT 7.950 409.050 10.050 411.150 ;
        RECT 16.950 408.750 18.150 412.050 ;
        RECT 19.950 410.850 22.050 412.950 ;
        RECT 22.950 412.050 25.050 414.150 ;
        RECT 28.950 412.050 31.050 414.150 ;
        RECT 31.950 410.850 34.050 412.950 ;
        RECT 34.950 412.050 37.050 414.150 ;
        RECT 49.950 413.850 52.050 415.950 ;
        RECT 52.950 415.050 55.050 417.150 ;
        RECT 62.700 415.950 63.600 424.200 ;
        RECT 68.100 420.150 69.900 421.950 ;
        RECT 77.100 420.150 78.900 421.950 ;
        RECT 64.950 417.150 66.750 418.950 ;
        RECT 67.950 418.050 70.050 420.150 ;
        RECT 71.100 417.150 72.900 418.950 ;
        RECT 74.100 417.150 75.900 418.950 ;
        RECT 76.950 418.050 79.050 420.150 ;
        RECT 80.250 417.150 82.050 418.950 ;
        RECT 50.100 412.050 51.900 413.850 ;
        RECT 20.100 409.050 21.900 410.850 ;
        RECT 32.100 409.050 33.900 410.850 ;
        RECT 14.400 407.700 18.150 408.750 ;
        RECT 35.850 408.750 37.050 412.050 ;
        RECT 35.850 407.700 39.600 408.750 ;
        RECT 53.400 407.700 54.600 415.050 ;
        RECT 55.950 413.850 58.050 415.950 ;
        RECT 61.950 413.850 64.050 415.950 ;
        RECT 64.950 415.050 67.050 417.150 ;
        RECT 70.950 415.050 73.050 417.150 ;
        RECT 73.950 415.050 76.050 417.150 ;
        RECT 79.950 415.050 82.050 417.150 ;
        RECT 83.400 415.950 84.300 424.200 ;
        RECT 95.400 417.150 96.600 425.400 ;
        RECT 104.700 425.100 106.200 425.400 ;
        RECT 110.400 425.400 112.200 431.400 ;
        RECT 121.800 425.400 123.600 431.400 ;
        RECT 134.400 425.400 136.200 431.400 ;
        RECT 110.400 425.100 111.300 425.400 ;
        RECT 104.700 424.200 111.300 425.100 ;
        RECT 104.100 420.150 105.900 421.950 ;
        RECT 101.100 417.150 102.900 418.950 ;
        RECT 103.950 418.050 106.050 420.150 ;
        RECT 107.250 417.150 109.050 418.950 ;
        RECT 82.950 413.850 85.050 415.950 ;
        RECT 91.950 413.850 94.050 415.950 ;
        RECT 94.950 415.050 97.050 417.150 ;
        RECT 56.100 412.050 57.900 413.850 ;
        RECT 62.700 409.650 63.600 413.850 ;
        RECT 83.400 409.650 84.300 413.850 ;
        RECT 92.100 412.050 93.900 413.850 ;
        RECT 62.700 408.000 66.900 409.650 ;
        RECT 14.400 405.600 15.600 407.700 ;
        RECT 4.800 399.600 6.600 402.600 ;
        RECT 13.800 399.600 15.600 405.600 ;
        RECT 16.800 404.700 24.600 406.050 ;
        RECT 16.800 399.600 18.600 404.700 ;
        RECT 22.800 399.600 24.600 404.700 ;
        RECT 29.400 404.700 37.200 406.050 ;
        RECT 29.400 399.600 31.200 404.700 ;
        RECT 35.400 399.600 37.200 404.700 ;
        RECT 38.400 405.600 39.600 407.700 ;
        RECT 51.000 406.800 54.600 407.700 ;
        RECT 38.400 399.600 40.200 405.600 ;
        RECT 51.000 399.600 52.800 406.800 ;
        RECT 65.100 399.600 66.900 408.000 ;
        RECT 80.100 408.000 84.300 409.650 ;
        RECT 80.100 399.600 81.900 408.000 ;
        RECT 95.400 407.700 96.600 415.050 ;
        RECT 97.950 413.850 100.050 415.950 ;
        RECT 100.950 415.050 103.050 417.150 ;
        RECT 106.950 415.050 109.050 417.150 ;
        RECT 110.400 415.950 111.300 424.200 ;
        RECT 122.400 417.150 123.600 425.400 ;
        RECT 109.950 413.850 112.050 415.950 ;
        RECT 118.950 413.850 121.050 415.950 ;
        RECT 121.950 415.050 124.050 417.150 ;
        RECT 98.100 412.050 99.900 413.850 ;
        RECT 110.400 409.650 111.300 413.850 ;
        RECT 119.100 412.050 120.900 413.850 ;
        RECT 93.000 406.800 96.600 407.700 ;
        RECT 107.100 408.000 111.300 409.650 ;
        RECT 93.000 399.600 94.800 406.800 ;
        RECT 107.100 399.600 108.900 408.000 ;
        RECT 122.400 407.700 123.600 415.050 ;
        RECT 124.950 413.850 127.050 415.950 ;
        RECT 131.100 414.150 132.900 415.950 ;
        RECT 125.100 412.050 126.900 413.850 ;
        RECT 130.950 412.050 133.050 414.150 ;
        RECT 134.550 408.300 135.600 425.400 ;
        RECT 141.000 419.400 142.800 431.400 ;
        RECT 151.500 419.400 153.300 431.400 ;
        RECT 164.400 425.400 166.200 431.400 ;
        RECT 176.400 425.400 178.200 431.400 ;
        RECT 136.950 413.850 139.050 415.950 ;
        RECT 141.000 414.150 142.050 419.400 ;
        RECT 146.100 414.150 147.900 415.950 ;
        RECT 151.950 414.150 153.150 419.400 ;
        RECT 154.950 417.150 156.750 418.950 ;
        RECT 164.400 417.150 165.600 425.400 ;
        RECT 176.700 425.100 178.200 425.400 ;
        RECT 182.400 425.400 184.200 431.400 ;
        RECT 191.400 425.400 193.200 431.400 ;
        RECT 206.400 425.400 208.200 431.400 ;
        RECT 182.400 425.100 183.300 425.400 ;
        RECT 176.700 424.200 183.300 425.100 ;
        RECT 176.100 420.150 177.900 421.950 ;
        RECT 173.100 417.150 174.900 418.950 ;
        RECT 175.950 418.050 178.050 420.150 ;
        RECT 179.250 417.150 181.050 418.950 ;
        RECT 154.950 415.050 157.050 417.150 ;
        RECT 137.100 412.050 138.900 413.850 ;
        RECT 139.950 412.050 142.050 414.150 ;
        RECT 145.950 412.050 148.050 414.150 ;
        RECT 120.000 406.800 123.600 407.700 ;
        RECT 131.400 407.100 138.900 408.300 ;
        RECT 120.000 399.600 121.800 406.800 ;
        RECT 131.400 399.600 133.200 407.100 ;
        RECT 137.100 406.500 138.900 407.100 ;
        RECT 141.000 405.600 142.050 412.050 ;
        RECT 148.950 410.850 151.050 412.950 ;
        RECT 151.950 412.050 154.050 414.150 ;
        RECT 160.950 413.850 163.050 415.950 ;
        RECT 163.950 415.050 166.050 417.150 ;
        RECT 161.100 412.050 162.900 413.850 ;
        RECT 149.100 409.050 150.900 410.850 ;
        RECT 152.850 408.750 154.050 412.050 ;
        RECT 152.850 407.700 156.600 408.750 ;
        RECT 138.900 404.100 142.050 405.600 ;
        RECT 146.400 404.700 154.200 406.050 ;
        RECT 138.900 399.600 140.700 404.100 ;
        RECT 146.400 399.600 148.200 404.700 ;
        RECT 152.400 399.600 154.200 404.700 ;
        RECT 155.400 405.600 156.600 407.700 ;
        RECT 164.400 407.700 165.600 415.050 ;
        RECT 166.950 413.850 169.050 415.950 ;
        RECT 172.950 415.050 175.050 417.150 ;
        RECT 178.950 415.050 181.050 417.150 ;
        RECT 182.400 415.950 183.300 424.200 ;
        RECT 191.400 417.150 192.600 425.400 ;
        RECT 181.950 413.850 184.050 415.950 ;
        RECT 187.950 413.850 190.050 415.950 ;
        RECT 190.950 415.050 193.050 417.150 ;
        RECT 167.100 412.050 168.900 413.850 ;
        RECT 182.400 409.650 183.300 413.850 ;
        RECT 188.100 412.050 189.900 413.850 ;
        RECT 179.100 408.000 183.300 409.650 ;
        RECT 164.400 406.800 168.000 407.700 ;
        RECT 155.400 399.600 157.200 405.600 ;
        RECT 166.200 399.600 168.000 406.800 ;
        RECT 179.100 399.600 180.900 408.000 ;
        RECT 191.400 407.700 192.600 415.050 ;
        RECT 193.950 413.850 196.050 415.950 ;
        RECT 194.100 412.050 195.900 413.850 ;
        RECT 206.400 412.950 207.600 425.400 ;
        RECT 217.500 419.400 219.300 431.400 ;
        RECT 232.500 419.400 234.300 431.400 ;
        RECT 248.400 425.400 250.200 431.400 ;
        RECT 257.400 425.400 259.200 431.400 ;
        RECT 212.100 414.150 213.900 415.950 ;
        RECT 217.950 414.150 219.150 419.400 ;
        RECT 220.950 417.150 222.750 418.950 ;
        RECT 220.950 415.050 223.050 417.150 ;
        RECT 227.100 414.150 228.900 415.950 ;
        RECT 232.950 414.150 234.150 419.400 ;
        RECT 235.950 417.150 237.750 418.950 ;
        RECT 235.950 415.050 238.050 417.150 ;
        RECT 203.100 411.150 204.900 412.950 ;
        RECT 202.950 409.050 205.050 411.150 ;
        RECT 205.950 410.850 208.050 412.950 ;
        RECT 211.950 412.050 214.050 414.150 ;
        RECT 214.950 410.850 217.050 412.950 ;
        RECT 217.950 412.050 220.050 414.150 ;
        RECT 226.950 412.050 229.050 414.150 ;
        RECT 191.400 406.800 195.000 407.700 ;
        RECT 193.200 399.600 195.000 406.800 ;
        RECT 206.400 402.600 207.600 410.850 ;
        RECT 215.100 409.050 216.900 410.850 ;
        RECT 218.850 408.750 220.050 412.050 ;
        RECT 229.950 410.850 232.050 412.950 ;
        RECT 232.950 412.050 235.050 414.150 ;
        RECT 248.400 412.950 249.600 425.400 ;
        RECT 257.400 417.150 258.600 425.400 ;
        RECT 271.500 419.400 273.300 431.400 ;
        RECT 283.800 419.400 285.600 431.400 ;
        RECT 286.800 420.300 288.600 431.400 ;
        RECT 292.800 420.300 294.600 431.400 ;
        RECT 286.800 419.400 294.600 420.300 ;
        RECT 305.700 419.400 307.500 431.400 ;
        RECT 320.700 419.400 322.500 431.400 ;
        RECT 335.700 419.400 337.500 431.400 ;
        RECT 347.400 425.400 349.200 431.400 ;
        RECT 253.950 413.850 256.050 415.950 ;
        RECT 256.950 415.050 259.050 417.150 ;
        RECT 230.100 409.050 231.900 410.850 ;
        RECT 233.850 408.750 235.050 412.050 ;
        RECT 245.100 411.150 246.900 412.950 ;
        RECT 244.950 409.050 247.050 411.150 ;
        RECT 247.950 410.850 250.050 412.950 ;
        RECT 254.100 412.050 255.900 413.850 ;
        RECT 218.850 407.700 222.600 408.750 ;
        RECT 233.850 407.700 237.600 408.750 ;
        RECT 212.400 404.700 220.200 406.050 ;
        RECT 206.400 399.600 208.200 402.600 ;
        RECT 212.400 399.600 214.200 404.700 ;
        RECT 218.400 399.600 220.200 404.700 ;
        RECT 221.400 405.600 222.600 407.700 ;
        RECT 221.400 399.600 223.200 405.600 ;
        RECT 227.400 404.700 235.200 406.050 ;
        RECT 227.400 399.600 229.200 404.700 ;
        RECT 233.400 399.600 235.200 404.700 ;
        RECT 236.400 405.600 237.600 407.700 ;
        RECT 236.400 399.600 238.200 405.600 ;
        RECT 248.400 402.600 249.600 410.850 ;
        RECT 257.400 407.700 258.600 415.050 ;
        RECT 259.950 413.850 262.050 415.950 ;
        RECT 266.100 414.150 267.900 415.950 ;
        RECT 271.950 414.150 273.150 419.400 ;
        RECT 274.950 417.150 276.750 418.950 ;
        RECT 274.950 415.050 277.050 417.150 ;
        RECT 284.400 414.150 285.300 419.400 ;
        RECT 302.250 417.150 304.050 418.950 ;
        RECT 301.950 415.050 304.050 417.150 ;
        RECT 305.850 414.150 307.050 419.400 ;
        RECT 317.250 417.150 319.050 418.950 ;
        RECT 311.100 414.150 312.900 415.950 ;
        RECT 316.950 415.050 319.050 417.150 ;
        RECT 320.850 414.150 322.050 419.400 ;
        RECT 332.250 417.150 334.050 418.950 ;
        RECT 326.100 414.150 327.900 415.950 ;
        RECT 331.950 415.050 334.050 417.150 ;
        RECT 335.850 414.150 337.050 419.400 ;
        RECT 347.400 417.150 348.600 425.400 ;
        RECT 358.800 419.400 360.600 431.400 ;
        RECT 361.800 420.300 363.600 431.400 ;
        RECT 367.800 420.300 369.600 431.400 ;
        RECT 361.800 419.400 369.600 420.300 ;
        RECT 377.700 419.400 379.500 431.400 ;
        RECT 385.950 421.950 388.050 424.050 ;
        RECT 341.100 414.150 342.900 415.950 ;
        RECT 260.100 412.050 261.900 413.850 ;
        RECT 265.950 412.050 268.050 414.150 ;
        RECT 268.950 410.850 271.050 412.950 ;
        RECT 271.950 412.050 274.050 414.150 ;
        RECT 283.950 412.050 286.050 414.150 ;
        RECT 269.100 409.050 270.900 410.850 ;
        RECT 272.850 408.750 274.050 412.050 ;
        RECT 272.850 407.700 276.600 408.750 ;
        RECT 257.400 406.800 261.000 407.700 ;
        RECT 248.400 399.600 250.200 402.600 ;
        RECT 259.200 399.600 261.000 406.800 ;
        RECT 266.400 404.700 274.200 406.050 ;
        RECT 266.400 399.600 268.200 404.700 ;
        RECT 272.400 399.600 274.200 404.700 ;
        RECT 275.400 405.600 276.600 407.700 ;
        RECT 284.400 405.600 285.300 412.050 ;
        RECT 286.950 410.850 289.050 412.950 ;
        RECT 290.100 411.150 291.900 412.950 ;
        RECT 287.100 409.050 288.900 410.850 ;
        RECT 289.950 409.050 292.050 411.150 ;
        RECT 292.950 410.850 295.050 412.950 ;
        RECT 304.950 412.050 307.050 414.150 ;
        RECT 293.100 409.050 294.900 410.850 ;
        RECT 304.950 408.750 306.150 412.050 ;
        RECT 307.950 410.850 310.050 412.950 ;
        RECT 310.950 412.050 313.050 414.150 ;
        RECT 319.950 412.050 322.050 414.150 ;
        RECT 308.100 409.050 309.900 410.850 ;
        RECT 319.950 408.750 321.150 412.050 ;
        RECT 322.950 410.850 325.050 412.950 ;
        RECT 325.950 412.050 328.050 414.150 ;
        RECT 334.950 412.050 337.050 414.150 ;
        RECT 323.100 409.050 324.900 410.850 ;
        RECT 334.950 408.750 336.150 412.050 ;
        RECT 337.950 410.850 340.050 412.950 ;
        RECT 340.950 412.050 343.050 414.150 ;
        RECT 343.950 413.850 346.050 415.950 ;
        RECT 346.950 415.050 349.050 417.150 ;
        RECT 344.100 412.050 345.900 413.850 ;
        RECT 338.100 409.050 339.900 410.850 ;
        RECT 302.400 407.700 306.150 408.750 ;
        RECT 317.400 407.700 321.150 408.750 ;
        RECT 332.400 407.700 336.150 408.750 ;
        RECT 347.400 407.700 348.600 415.050 ;
        RECT 349.950 413.850 352.050 415.950 ;
        RECT 359.400 414.150 360.300 419.400 ;
        RECT 374.250 417.150 376.050 418.950 ;
        RECT 373.950 415.050 376.050 417.150 ;
        RECT 377.850 414.150 379.050 419.400 ;
        RECT 383.100 414.150 384.900 415.950 ;
        RECT 350.100 412.050 351.900 413.850 ;
        RECT 358.950 412.050 361.050 414.150 ;
        RECT 302.400 405.600 303.600 407.700 ;
        RECT 275.400 399.600 277.200 405.600 ;
        RECT 284.400 403.950 289.800 405.600 ;
        RECT 288.000 399.600 289.800 403.950 ;
        RECT 301.800 399.600 303.600 405.600 ;
        RECT 304.800 404.700 312.600 406.050 ;
        RECT 317.400 405.600 318.600 407.700 ;
        RECT 304.800 399.600 306.600 404.700 ;
        RECT 310.800 399.600 312.600 404.700 ;
        RECT 316.800 399.600 318.600 405.600 ;
        RECT 319.800 404.700 327.600 406.050 ;
        RECT 332.400 405.600 333.600 407.700 ;
        RECT 347.400 406.800 351.000 407.700 ;
        RECT 319.800 399.600 321.600 404.700 ;
        RECT 325.800 399.600 327.600 404.700 ;
        RECT 331.800 399.600 333.600 405.600 ;
        RECT 334.800 404.700 342.600 406.050 ;
        RECT 334.800 399.600 336.600 404.700 ;
        RECT 340.800 399.600 342.600 404.700 ;
        RECT 349.200 399.600 351.000 406.800 ;
        RECT 359.400 405.600 360.300 412.050 ;
        RECT 361.950 410.850 364.050 412.950 ;
        RECT 365.100 411.150 366.900 412.950 ;
        RECT 362.100 409.050 363.900 410.850 ;
        RECT 364.950 409.050 367.050 411.150 ;
        RECT 367.950 410.850 370.050 412.950 ;
        RECT 376.950 412.050 379.050 414.150 ;
        RECT 368.100 409.050 369.900 410.850 ;
        RECT 376.950 408.750 378.150 412.050 ;
        RECT 379.950 410.850 382.050 412.950 ;
        RECT 382.950 412.050 385.050 414.150 ;
        RECT 380.100 409.050 381.900 410.850 ;
        RECT 374.400 407.700 378.150 408.750 ;
        RECT 386.550 408.450 387.450 421.950 ;
        RECT 394.800 419.400 396.600 431.400 ;
        RECT 403.800 430.500 411.600 431.400 ;
        RECT 403.800 419.400 405.600 430.500 ;
        RECT 394.950 412.950 396.300 419.400 ;
        RECT 406.800 418.500 408.600 429.600 ;
        RECT 409.800 420.600 411.600 430.500 ;
        RECT 415.800 420.600 417.600 431.400 ;
        RECT 409.800 419.700 417.600 420.600 ;
        RECT 422.400 425.400 424.200 431.400 ;
        RECT 428.400 425.400 430.200 431.400 ;
        RECT 406.800 417.600 410.850 418.500 ;
        RECT 404.100 414.150 405.900 415.950 ;
        RECT 409.950 414.150 410.850 417.600 ;
        RECT 415.950 414.150 417.750 415.950 ;
        RECT 391.950 410.850 396.300 412.950 ;
        RECT 397.950 410.850 400.050 412.950 ;
        RECT 403.950 412.050 406.050 414.150 ;
        RECT 406.950 410.850 409.050 412.950 ;
        RECT 409.950 412.050 412.050 414.150 ;
        RECT 391.950 408.450 394.050 409.050 ;
        RECT 374.400 405.600 375.600 407.700 ;
        RECT 386.550 407.550 394.050 408.450 ;
        RECT 391.950 406.950 394.050 407.550 ;
        RECT 359.400 403.950 364.800 405.600 ;
        RECT 363.000 399.600 364.800 403.950 ;
        RECT 373.800 399.600 375.600 405.600 ;
        RECT 376.800 404.700 384.600 406.050 ;
        RECT 394.950 405.600 396.300 410.850 ;
        RECT 398.100 409.050 399.900 410.850 ;
        RECT 407.250 409.050 409.050 410.850 ;
        RECT 411.000 405.600 412.050 412.050 ;
        RECT 412.950 410.850 415.050 412.950 ;
        RECT 415.950 412.050 418.050 414.150 ;
        RECT 422.400 412.950 423.600 425.400 ;
        RECT 428.400 418.500 429.600 425.400 ;
        RECT 434.700 419.400 436.500 431.400 ;
        RECT 442.500 419.400 444.300 431.400 ;
        RECT 448.800 425.400 450.600 431.400 ;
        RECT 460.800 425.400 462.600 431.400 ;
        RECT 469.800 425.400 471.600 431.400 ;
        RECT 428.400 417.600 434.100 418.500 ;
        RECT 432.150 416.700 434.100 417.600 ;
        RECT 428.100 414.150 429.900 415.950 ;
        RECT 419.100 411.150 420.900 412.950 ;
        RECT 412.950 409.050 414.750 410.850 ;
        RECT 418.950 409.050 421.050 411.150 ;
        RECT 421.950 410.850 424.050 412.950 ;
        RECT 427.950 412.050 430.050 414.150 ;
        RECT 376.800 399.600 378.600 404.700 ;
        RECT 382.800 399.600 384.600 404.700 ;
        RECT 394.800 399.600 396.600 405.600 ;
        RECT 411.000 399.600 412.800 405.600 ;
        RECT 422.400 402.600 423.600 410.850 ;
        RECT 432.150 408.300 433.050 416.700 ;
        RECT 435.000 414.150 436.200 419.400 ;
        RECT 433.950 412.050 436.200 414.150 ;
        RECT 432.150 407.400 434.100 408.300 ;
        RECT 429.000 406.500 434.100 407.400 ;
        RECT 429.000 402.600 430.200 406.500 ;
        RECT 435.000 405.600 436.200 412.050 ;
        RECT 442.800 414.150 444.000 419.400 ;
        RECT 449.400 418.500 450.600 425.400 ;
        RECT 444.900 417.600 450.600 418.500 ;
        RECT 444.900 416.700 446.850 417.600 ;
        RECT 461.400 417.150 462.600 425.400 ;
        RECT 442.800 412.050 445.050 414.150 ;
        RECT 442.800 405.600 444.000 412.050 ;
        RECT 445.950 408.300 446.850 416.700 ;
        RECT 449.100 414.150 450.900 415.950 ;
        RECT 448.950 412.050 451.050 414.150 ;
        RECT 457.950 413.850 460.050 415.950 ;
        RECT 460.950 415.050 463.050 417.150 ;
        RECT 458.100 412.050 459.900 413.850 ;
        RECT 444.900 407.400 446.850 408.300 ;
        RECT 461.400 407.700 462.600 415.050 ;
        RECT 463.950 413.850 466.050 415.950 ;
        RECT 464.100 412.050 465.900 413.850 ;
        RECT 470.400 412.950 471.600 425.400 ;
        RECT 482.700 419.400 484.500 431.400 ;
        RECT 493.200 430.500 501.000 431.400 ;
        RECT 493.200 421.200 495.000 430.500 ;
        RECT 496.200 421.800 498.000 429.600 ;
        RECT 496.800 419.400 498.000 421.800 ;
        RECT 499.200 421.800 501.000 430.500 ;
        RECT 502.800 430.500 510.600 431.400 ;
        RECT 502.800 422.700 504.600 430.500 ;
        RECT 505.800 421.800 507.600 429.600 ;
        RECT 499.200 420.900 507.600 421.800 ;
        RECT 508.800 421.500 510.600 430.500 ;
        RECT 514.800 421.500 516.600 431.400 ;
        RECT 508.800 420.600 516.600 421.500 ;
        RECT 527.700 419.400 529.500 431.400 ;
        RECT 539.400 425.400 541.200 431.400 ;
        RECT 545.400 425.400 547.200 431.400 ;
        RECT 479.250 417.150 481.050 418.950 ;
        RECT 478.950 415.050 481.050 417.150 ;
        RECT 482.850 414.150 484.050 419.400 ;
        RECT 496.800 418.200 500.250 419.400 ;
        RECT 488.100 414.150 489.900 415.950 ;
        RECT 469.950 410.850 472.050 412.950 ;
        RECT 473.100 411.150 474.900 412.950 ;
        RECT 481.950 412.050 484.050 414.150 ;
        RECT 444.900 406.500 450.000 407.400 ;
        RECT 422.400 399.600 424.200 402.600 ;
        RECT 428.400 399.600 430.200 402.600 ;
        RECT 434.700 399.600 436.500 405.600 ;
        RECT 442.500 399.600 444.300 405.600 ;
        RECT 448.800 402.600 450.000 406.500 ;
        RECT 459.000 406.800 462.600 407.700 ;
        RECT 448.800 399.600 450.600 402.600 ;
        RECT 459.000 399.600 460.800 406.800 ;
        RECT 470.400 402.600 471.600 410.850 ;
        RECT 472.950 409.050 475.050 411.150 ;
        RECT 481.950 408.750 483.150 412.050 ;
        RECT 484.950 410.850 487.050 412.950 ;
        RECT 487.950 412.050 490.050 414.150 ;
        RECT 499.050 412.800 500.250 418.200 ;
        RECT 524.250 417.150 526.050 418.950 ;
        RECT 503.100 414.000 504.900 415.800 ;
        RECT 512.100 414.000 513.900 415.800 ;
        RECT 523.950 415.050 526.050 417.150 ;
        RECT 527.850 414.150 529.050 419.400 ;
        RECT 533.100 414.150 534.900 415.950 ;
        RECT 485.100 409.050 486.900 410.850 ;
        RECT 496.950 410.700 500.250 412.800 ;
        RECT 502.950 411.900 505.050 414.000 ;
        RECT 505.950 410.700 508.050 412.800 ;
        RECT 511.950 411.900 514.050 414.000 ;
        RECT 526.950 412.050 529.050 414.150 ;
        RECT 479.400 407.700 483.150 408.750 ;
        RECT 479.400 405.600 480.600 407.700 ;
        RECT 469.800 399.600 471.600 402.600 ;
        RECT 478.800 399.600 480.600 405.600 ;
        RECT 481.800 404.700 489.600 406.050 ;
        RECT 481.800 399.600 483.600 404.700 ;
        RECT 487.800 399.600 489.600 404.700 ;
        RECT 499.050 404.400 500.250 410.700 ;
        RECT 506.100 408.900 507.900 410.700 ;
        RECT 526.950 408.750 528.150 412.050 ;
        RECT 529.950 410.850 532.050 412.950 ;
        RECT 532.950 412.050 535.050 414.150 ;
        RECT 539.400 412.950 540.600 425.400 ;
        RECT 545.400 418.500 546.600 425.400 ;
        RECT 551.700 419.400 553.500 431.400 ;
        RECT 562.800 425.400 564.600 431.400 ;
        RECT 563.700 425.100 564.600 425.400 ;
        RECT 568.800 425.400 570.600 431.400 ;
        RECT 568.800 425.100 570.300 425.400 ;
        RECT 563.700 424.200 570.300 425.100 ;
        RECT 545.400 417.600 551.100 418.500 ;
        RECT 549.150 416.700 551.100 417.600 ;
        RECT 545.100 414.150 546.900 415.950 ;
        RECT 536.100 411.150 537.900 412.950 ;
        RECT 530.100 409.050 531.900 410.850 ;
        RECT 535.950 409.050 538.050 411.150 ;
        RECT 538.950 410.850 541.050 412.950 ;
        RECT 544.950 412.050 547.050 414.150 ;
        RECT 524.400 407.700 528.150 408.750 ;
        RECT 524.400 405.600 525.600 407.700 ;
        RECT 499.050 403.500 509.850 404.400 ;
        RECT 502.800 402.600 503.850 403.500 ;
        RECT 508.800 402.600 509.850 403.500 ;
        RECT 502.800 399.600 504.600 402.600 ;
        RECT 508.800 399.600 510.600 402.600 ;
        RECT 523.800 399.600 525.600 405.600 ;
        RECT 526.800 404.700 534.600 406.050 ;
        RECT 526.800 399.600 528.600 404.700 ;
        RECT 532.800 399.600 534.600 404.700 ;
        RECT 539.400 402.600 540.600 410.850 ;
        RECT 549.150 408.300 550.050 416.700 ;
        RECT 552.000 414.150 553.200 419.400 ;
        RECT 563.700 415.950 564.600 424.200 ;
        RECT 569.100 420.150 570.900 421.950 ;
        RECT 565.950 417.150 567.750 418.950 ;
        RECT 568.950 418.050 571.050 420.150 ;
        RECT 577.800 419.400 579.600 431.400 ;
        RECT 580.800 420.300 582.600 431.400 ;
        RECT 586.800 420.300 588.600 431.400 ;
        RECT 580.800 419.400 588.600 420.300 ;
        RECT 596.700 419.400 598.500 431.400 ;
        RECT 610.500 419.400 612.300 431.400 ;
        RECT 622.800 425.400 624.600 431.400 ;
        RECT 623.700 425.100 624.600 425.400 ;
        RECT 628.800 425.400 630.600 431.400 ;
        RECT 628.800 425.100 630.300 425.400 ;
        RECT 623.700 424.200 630.300 425.100 ;
        RECT 613.950 423.450 616.050 424.050 ;
        RECT 613.950 422.550 618.450 423.450 ;
        RECT 613.950 421.950 616.050 422.550 ;
        RECT 572.100 417.150 573.900 418.950 ;
        RECT 550.950 412.050 553.200 414.150 ;
        RECT 562.950 413.850 565.050 415.950 ;
        RECT 565.950 415.050 568.050 417.150 ;
        RECT 571.950 415.050 574.050 417.150 ;
        RECT 578.400 414.150 579.300 419.400 ;
        RECT 593.250 417.150 595.050 418.950 ;
        RECT 592.950 415.050 595.050 417.150 ;
        RECT 596.850 414.150 598.050 419.400 ;
        RECT 602.100 414.150 603.900 415.950 ;
        RECT 605.100 414.150 606.900 415.950 ;
        RECT 610.950 414.150 612.150 419.400 ;
        RECT 613.950 417.150 615.750 418.950 ;
        RECT 613.950 415.050 616.050 417.150 ;
        RECT 549.150 407.400 551.100 408.300 ;
        RECT 546.000 406.500 551.100 407.400 ;
        RECT 546.000 402.600 547.200 406.500 ;
        RECT 552.000 405.600 553.200 412.050 ;
        RECT 563.700 409.650 564.600 413.850 ;
        RECT 577.950 412.050 580.050 414.150 ;
        RECT 563.700 408.000 567.900 409.650 ;
        RECT 539.400 399.600 541.200 402.600 ;
        RECT 545.400 399.600 547.200 402.600 ;
        RECT 551.700 399.600 553.500 405.600 ;
        RECT 566.100 399.600 567.900 408.000 ;
        RECT 578.400 405.600 579.300 412.050 ;
        RECT 580.950 410.850 583.050 412.950 ;
        RECT 584.100 411.150 585.900 412.950 ;
        RECT 581.100 409.050 582.900 410.850 ;
        RECT 583.950 409.050 586.050 411.150 ;
        RECT 586.950 410.850 589.050 412.950 ;
        RECT 595.950 412.050 598.050 414.150 ;
        RECT 587.100 409.050 588.900 410.850 ;
        RECT 595.950 408.750 597.150 412.050 ;
        RECT 598.950 410.850 601.050 412.950 ;
        RECT 601.950 412.050 604.050 414.150 ;
        RECT 604.950 412.050 607.050 414.150 ;
        RECT 607.950 410.850 610.050 412.950 ;
        RECT 610.950 412.050 613.050 414.150 ;
        RECT 617.550 412.050 618.450 422.550 ;
        RECT 623.700 415.950 624.600 424.200 ;
        RECT 629.100 420.150 630.900 421.950 ;
        RECT 635.400 420.300 637.200 431.400 ;
        RECT 641.400 420.300 643.200 431.400 ;
        RECT 625.950 417.150 627.750 418.950 ;
        RECT 628.950 418.050 631.050 420.150 ;
        RECT 635.400 419.400 643.200 420.300 ;
        RECT 644.400 419.400 646.200 431.400 ;
        RECT 650.400 420.600 652.200 431.400 ;
        RECT 656.400 430.500 664.200 431.400 ;
        RECT 656.400 420.600 658.200 430.500 ;
        RECT 650.400 419.700 658.200 420.600 ;
        RECT 632.100 417.150 633.900 418.950 ;
        RECT 622.950 413.850 625.050 415.950 ;
        RECT 625.950 415.050 628.050 417.150 ;
        RECT 631.950 415.050 634.050 417.150 ;
        RECT 644.700 414.150 645.600 419.400 ;
        RECT 659.400 418.500 661.200 429.600 ;
        RECT 662.400 419.400 664.200 430.500 ;
        RECT 673.800 425.400 675.600 431.400 ;
        RECT 646.950 415.950 649.050 418.050 ;
        RECT 657.150 417.600 661.200 418.500 ;
        RECT 599.100 409.050 600.900 410.850 ;
        RECT 608.100 409.050 609.900 410.850 ;
        RECT 593.400 407.700 597.150 408.750 ;
        RECT 611.850 408.750 613.050 412.050 ;
        RECT 616.950 409.950 619.050 412.050 ;
        RECT 623.700 409.650 624.600 413.850 ;
        RECT 634.950 410.850 637.050 412.950 ;
        RECT 638.100 411.150 639.900 412.950 ;
        RECT 611.850 407.700 615.600 408.750 ;
        RECT 623.700 408.000 627.900 409.650 ;
        RECT 635.100 409.050 636.900 410.850 ;
        RECT 637.950 409.050 640.050 411.150 ;
        RECT 640.950 410.850 643.050 412.950 ;
        RECT 643.950 412.050 646.050 414.150 ;
        RECT 641.100 409.050 642.900 410.850 ;
        RECT 593.400 405.600 594.600 407.700 ;
        RECT 578.400 403.950 583.800 405.600 ;
        RECT 582.000 399.600 583.800 403.950 ;
        RECT 592.800 399.600 594.600 405.600 ;
        RECT 595.800 404.700 603.600 406.050 ;
        RECT 595.800 399.600 597.600 404.700 ;
        RECT 601.800 399.600 603.600 404.700 ;
        RECT 605.400 404.700 613.200 406.050 ;
        RECT 605.400 399.600 607.200 404.700 ;
        RECT 611.400 399.600 613.200 404.700 ;
        RECT 614.400 405.600 615.600 407.700 ;
        RECT 614.400 399.600 616.200 405.600 ;
        RECT 626.100 399.600 627.900 408.000 ;
        RECT 644.700 405.600 645.600 412.050 ;
        RECT 647.550 408.450 648.450 415.950 ;
        RECT 650.250 414.150 652.050 415.950 ;
        RECT 657.150 414.150 658.050 417.600 ;
        RECT 674.400 417.150 675.600 425.400 ;
        RECT 682.800 419.400 684.600 431.400 ;
        RECT 685.800 420.300 687.600 431.400 ;
        RECT 691.800 420.300 693.600 431.400 ;
        RECT 698.400 425.400 700.200 431.400 ;
        RECT 698.700 425.100 700.200 425.400 ;
        RECT 704.400 425.400 706.200 431.400 ;
        RECT 704.400 425.100 705.300 425.400 ;
        RECT 698.700 424.200 705.300 425.100 ;
        RECT 685.800 419.400 693.600 420.300 ;
        RECT 698.100 420.150 699.900 421.950 ;
        RECT 662.100 414.150 663.900 415.950 ;
        RECT 649.950 412.050 652.050 414.150 ;
        RECT 652.950 410.850 655.050 412.950 ;
        RECT 653.250 409.050 655.050 410.850 ;
        RECT 655.950 412.050 658.050 414.150 ;
        RECT 649.950 408.450 652.050 409.050 ;
        RECT 647.550 407.550 652.050 408.450 ;
        RECT 649.950 406.950 652.050 407.550 ;
        RECT 655.950 405.600 657.000 412.050 ;
        RECT 658.950 410.850 661.050 412.950 ;
        RECT 661.950 412.050 664.050 414.150 ;
        RECT 670.950 413.850 673.050 415.950 ;
        RECT 673.950 415.050 676.050 417.150 ;
        RECT 671.100 412.050 672.900 413.850 ;
        RECT 658.950 409.050 660.750 410.850 ;
        RECT 674.400 407.700 675.600 415.050 ;
        RECT 676.950 413.850 679.050 415.950 ;
        RECT 683.400 414.150 684.300 419.400 ;
        RECT 695.100 417.150 696.900 418.950 ;
        RECT 697.950 418.050 700.050 420.150 ;
        RECT 701.250 417.150 703.050 418.950 ;
        RECT 694.950 415.050 697.050 417.150 ;
        RECT 700.950 415.050 703.050 417.150 ;
        RECT 704.400 415.950 705.300 424.200 ;
        RECT 712.800 419.400 714.600 431.400 ;
        RECT 715.800 420.300 717.600 431.400 ;
        RECT 721.800 420.300 723.600 431.400 ;
        RECT 728.400 425.400 730.200 431.400 ;
        RECT 728.700 425.100 730.200 425.400 ;
        RECT 734.400 425.400 736.200 431.400 ;
        RECT 743.400 425.400 745.200 431.400 ;
        RECT 734.400 425.100 735.300 425.400 ;
        RECT 728.700 424.200 735.300 425.100 ;
        RECT 743.700 425.100 745.200 425.400 ;
        RECT 749.400 425.400 751.200 431.400 ;
        RECT 749.400 425.100 750.300 425.400 ;
        RECT 743.700 424.200 750.300 425.100 ;
        RECT 715.800 419.400 723.600 420.300 ;
        RECT 728.100 420.150 729.900 421.950 ;
        RECT 677.100 412.050 678.900 413.850 ;
        RECT 682.950 412.050 685.050 414.150 ;
        RECT 703.950 413.850 706.050 415.950 ;
        RECT 713.400 414.150 714.300 419.400 ;
        RECT 725.100 417.150 726.900 418.950 ;
        RECT 727.950 418.050 730.050 420.150 ;
        RECT 731.250 417.150 733.050 418.950 ;
        RECT 724.950 415.050 727.050 417.150 ;
        RECT 730.950 415.050 733.050 417.150 ;
        RECT 734.400 415.950 735.300 424.200 ;
        RECT 743.100 420.150 744.900 421.950 ;
        RECT 740.100 417.150 741.900 418.950 ;
        RECT 742.950 418.050 745.050 420.150 ;
        RECT 746.250 417.150 748.050 418.950 ;
        RECT 640.200 403.950 645.600 405.600 ;
        RECT 640.200 399.600 642.000 403.950 ;
        RECT 655.200 399.600 657.000 405.600 ;
        RECT 672.000 406.800 675.600 407.700 ;
        RECT 672.000 399.600 673.800 406.800 ;
        RECT 683.400 405.600 684.300 412.050 ;
        RECT 685.950 410.850 688.050 412.950 ;
        RECT 689.100 411.150 690.900 412.950 ;
        RECT 686.100 409.050 687.900 410.850 ;
        RECT 688.950 409.050 691.050 411.150 ;
        RECT 691.950 410.850 694.050 412.950 ;
        RECT 692.100 409.050 693.900 410.850 ;
        RECT 704.400 409.650 705.300 413.850 ;
        RECT 712.950 412.050 715.050 414.150 ;
        RECT 733.950 413.850 736.050 415.950 ;
        RECT 739.950 415.050 742.050 417.150 ;
        RECT 745.950 415.050 748.050 417.150 ;
        RECT 749.400 415.950 750.300 424.200 ;
        RECT 748.950 413.850 751.050 415.950 ;
        RECT 701.100 408.000 705.300 409.650 ;
        RECT 683.400 403.950 688.800 405.600 ;
        RECT 687.000 399.600 688.800 403.950 ;
        RECT 701.100 399.600 702.900 408.000 ;
        RECT 713.400 405.600 714.300 412.050 ;
        RECT 715.950 410.850 718.050 412.950 ;
        RECT 719.100 411.150 720.900 412.950 ;
        RECT 716.100 409.050 717.900 410.850 ;
        RECT 718.950 409.050 721.050 411.150 ;
        RECT 721.950 410.850 724.050 412.950 ;
        RECT 722.100 409.050 723.900 410.850 ;
        RECT 734.400 409.650 735.300 413.850 ;
        RECT 749.400 409.650 750.300 413.850 ;
        RECT 731.100 408.000 735.300 409.650 ;
        RECT 746.100 408.000 750.300 409.650 ;
        RECT 713.400 403.950 718.800 405.600 ;
        RECT 717.000 399.600 718.800 403.950 ;
        RECT 731.100 399.600 732.900 408.000 ;
        RECT 746.100 399.600 747.900 408.000 ;
        RECT 4.800 389.400 6.600 395.400 ;
        RECT 10.800 392.400 12.600 395.400 ;
        RECT 4.950 384.150 6.000 389.400 ;
        RECT 10.800 388.200 11.700 392.400 ;
        RECT 8.250 387.300 11.700 388.200 ;
        RECT 21.000 388.200 22.800 395.400 ;
        RECT 37.200 388.200 39.000 395.400 ;
        RECT 21.000 387.300 24.600 388.200 ;
        RECT 8.250 386.400 10.050 387.300 ;
        RECT 4.950 382.050 7.050 384.150 ;
        RECT 5.700 375.450 7.050 382.050 ;
        RECT 8.400 378.150 9.300 386.400 ;
        RECT 13.950 383.850 16.050 385.950 ;
        RECT 10.950 380.850 13.050 382.950 ;
        RECT 14.100 382.050 15.900 383.850 ;
        RECT 20.100 381.150 21.900 382.950 ;
        RECT 11.100 379.050 12.900 380.850 ;
        RECT 19.950 379.050 22.050 381.150 ;
        RECT 23.400 379.950 24.600 387.300 ;
        RECT 25.950 387.450 28.050 388.050 ;
        RECT 25.950 386.550 30.450 387.450 ;
        RECT 25.950 385.950 28.050 386.550 ;
        RECT 26.100 381.150 27.900 382.950 ;
        RECT 8.400 378.000 10.200 378.150 ;
        RECT 8.400 376.800 15.600 378.000 ;
        RECT 22.950 377.850 25.050 379.950 ;
        RECT 25.950 379.050 28.050 381.150 ;
        RECT 8.400 376.350 10.200 376.800 ;
        RECT 14.400 375.600 15.600 376.800 ;
        RECT 5.700 374.100 8.100 375.450 ;
        RECT 6.300 363.600 8.100 374.100 ;
        RECT 13.800 363.600 15.600 375.600 ;
        RECT 23.400 369.600 24.600 377.850 ;
        RECT 29.550 375.450 30.450 386.550 ;
        RECT 35.400 387.300 39.000 388.200 ;
        RECT 47.400 392.400 49.200 395.400 ;
        RECT 32.100 381.150 33.900 382.950 ;
        RECT 31.950 379.050 34.050 381.150 ;
        RECT 35.400 379.950 36.600 387.300 ;
        RECT 43.950 383.850 46.050 385.950 ;
        RECT 47.400 384.150 48.600 392.400 ;
        RECT 55.800 389.400 57.600 395.400 ;
        RECT 56.400 387.300 57.600 389.400 ;
        RECT 58.800 390.300 60.600 395.400 ;
        RECT 64.800 390.300 66.600 395.400 ;
        RECT 70.800 392.400 72.600 395.400 ;
        RECT 58.800 388.950 66.600 390.300 ;
        RECT 56.400 386.250 60.150 387.300 ;
        RECT 38.100 381.150 39.900 382.950 ;
        RECT 44.100 382.050 45.900 383.850 ;
        RECT 46.950 382.050 49.050 384.150 ;
        RECT 58.950 382.950 60.150 386.250 ;
        RECT 62.100 384.150 63.900 385.950 ;
        RECT 71.400 384.150 72.600 392.400 ;
        RECT 85.200 391.050 87.000 395.400 ;
        RECT 85.200 389.400 90.600 391.050 ;
        RECT 34.950 377.850 37.050 379.950 ;
        RECT 37.950 379.050 40.050 381.150 ;
        RECT 31.950 375.450 34.050 376.050 ;
        RECT 29.550 374.550 34.050 375.450 ;
        RECT 31.950 373.950 34.050 374.550 ;
        RECT 22.800 363.600 24.600 369.600 ;
        RECT 35.400 369.600 36.600 377.850 ;
        RECT 47.400 369.600 48.600 382.050 ;
        RECT 58.950 380.850 61.050 382.950 ;
        RECT 61.950 382.050 64.050 384.150 ;
        RECT 64.950 380.850 67.050 382.950 ;
        RECT 70.950 382.050 73.050 384.150 ;
        RECT 73.950 383.850 76.050 385.950 ;
        RECT 80.100 384.150 81.900 385.950 ;
        RECT 74.100 382.050 75.900 383.850 ;
        RECT 79.950 382.050 82.050 384.150 ;
        RECT 82.950 383.850 85.050 385.950 ;
        RECT 86.100 384.150 87.900 385.950 ;
        RECT 83.100 382.050 84.900 383.850 ;
        RECT 85.950 382.050 88.050 384.150 ;
        RECT 89.700 382.950 90.600 389.400 ;
        RECT 101.100 387.000 102.900 395.400 ;
        RECT 116.100 387.000 117.900 395.400 ;
        RECT 127.800 392.400 129.600 395.400 ;
        RECT 101.100 385.350 105.300 387.000 ;
        RECT 116.100 385.350 120.300 387.000 ;
        RECT 55.950 377.850 58.050 379.950 ;
        RECT 56.250 376.050 58.050 377.850 ;
        RECT 59.850 375.600 61.050 380.850 ;
        RECT 65.100 379.050 66.900 380.850 ;
        RECT 35.400 363.600 37.200 369.600 ;
        RECT 47.400 363.600 49.200 369.600 ;
        RECT 59.700 363.600 61.500 375.600 ;
        RECT 71.400 369.600 72.600 382.050 ;
        RECT 88.950 380.850 91.050 382.950 ;
        RECT 104.400 381.150 105.300 385.350 ;
        RECT 119.400 381.150 120.300 385.350 ;
        RECT 128.400 384.150 129.600 392.400 ;
        RECT 139.800 389.400 141.600 395.400 ;
        RECT 145.800 392.400 147.600 395.400 ;
        RECT 127.950 382.050 130.050 384.150 ;
        RECT 130.950 383.850 133.050 385.950 ;
        RECT 139.950 384.150 141.000 389.400 ;
        RECT 145.800 388.200 146.700 392.400 ;
        RECT 143.250 387.300 146.700 388.200 ;
        RECT 143.250 386.400 145.050 387.300 ;
        RECT 158.100 387.000 159.900 395.400 ;
        RECT 178.800 392.400 180.600 395.400 ;
        RECT 184.800 392.400 186.600 395.400 ;
        RECT 197.400 392.400 199.200 395.400 ;
        RECT 178.800 391.500 179.850 392.400 ;
        RECT 184.800 391.500 185.850 392.400 ;
        RECT 175.050 390.600 185.850 391.500 ;
        RECT 131.100 382.050 132.900 383.850 ;
        RECT 139.950 382.050 142.050 384.150 ;
        RECT 89.700 375.600 90.600 380.850 ;
        RECT 94.950 377.850 97.050 379.950 ;
        RECT 100.950 377.850 103.050 379.950 ;
        RECT 103.950 379.050 106.050 381.150 ;
        RECT 95.100 376.050 96.900 377.850 ;
        RECT 70.800 363.600 72.600 369.600 ;
        RECT 80.400 374.700 88.200 375.600 ;
        RECT 80.400 363.600 82.200 374.700 ;
        RECT 86.400 363.600 88.200 374.700 ;
        RECT 89.400 363.600 91.200 375.600 ;
        RECT 97.950 374.850 100.050 376.950 ;
        RECT 101.250 376.050 103.050 377.850 ;
        RECT 98.100 373.050 99.900 374.850 ;
        RECT 104.400 370.800 105.300 379.050 ;
        RECT 109.950 377.850 112.050 379.950 ;
        RECT 115.950 377.850 118.050 379.950 ;
        RECT 118.950 379.050 121.050 381.150 ;
        RECT 110.100 376.050 111.900 377.850 ;
        RECT 112.950 374.850 115.050 376.950 ;
        RECT 116.250 376.050 118.050 377.850 ;
        RECT 113.100 373.050 114.900 374.850 ;
        RECT 119.400 370.800 120.300 379.050 ;
        RECT 98.700 369.900 105.300 370.800 ;
        RECT 98.700 369.600 100.200 369.900 ;
        RECT 98.400 363.600 100.200 369.600 ;
        RECT 104.400 369.600 105.300 369.900 ;
        RECT 113.700 369.900 120.300 370.800 ;
        RECT 113.700 369.600 115.200 369.900 ;
        RECT 104.400 363.600 106.200 369.600 ;
        RECT 113.400 363.600 115.200 369.600 ;
        RECT 119.400 369.600 120.300 369.900 ;
        RECT 128.400 369.600 129.600 382.050 ;
        RECT 140.700 375.450 142.050 382.050 ;
        RECT 143.400 378.150 144.300 386.400 ;
        RECT 148.950 383.850 151.050 385.950 ;
        RECT 158.100 385.350 162.300 387.000 ;
        RECT 145.950 380.850 148.050 382.950 ;
        RECT 149.100 382.050 150.900 383.850 ;
        RECT 161.400 381.150 162.300 385.350 ;
        RECT 175.050 384.300 176.250 390.600 ;
        RECT 182.100 384.300 183.900 386.100 ;
        RECT 172.950 382.200 176.250 384.300 ;
        RECT 146.100 379.050 147.900 380.850 ;
        RECT 143.400 378.000 145.200 378.150 ;
        RECT 143.400 376.800 150.600 378.000 ;
        RECT 151.950 377.850 154.050 379.950 ;
        RECT 157.950 377.850 160.050 379.950 ;
        RECT 160.950 379.050 163.050 381.150 ;
        RECT 143.400 376.350 145.200 376.800 ;
        RECT 149.400 375.600 150.600 376.800 ;
        RECT 152.100 376.050 153.900 377.850 ;
        RECT 140.700 374.100 143.100 375.450 ;
        RECT 119.400 363.600 121.200 369.600 ;
        RECT 127.800 363.600 129.600 369.600 ;
        RECT 141.300 363.600 143.100 374.100 ;
        RECT 148.800 363.600 150.600 375.600 ;
        RECT 154.950 374.850 157.050 376.950 ;
        RECT 158.250 376.050 160.050 377.850 ;
        RECT 155.100 373.050 156.900 374.850 ;
        RECT 161.400 370.800 162.300 379.050 ;
        RECT 175.050 376.800 176.250 382.200 ;
        RECT 178.950 381.000 181.050 383.100 ;
        RECT 181.950 382.200 184.050 384.300 ;
        RECT 193.950 383.850 196.050 385.950 ;
        RECT 197.400 384.150 198.600 392.400 ;
        RECT 206.400 390.300 208.200 395.400 ;
        RECT 212.400 390.300 214.200 395.400 ;
        RECT 206.400 388.950 214.200 390.300 ;
        RECT 215.400 389.400 217.200 395.400 ;
        RECT 221.400 390.300 223.200 395.400 ;
        RECT 227.400 390.300 229.200 395.400 ;
        RECT 215.400 387.300 216.600 389.400 ;
        RECT 221.400 388.950 229.200 390.300 ;
        RECT 230.400 389.400 232.200 395.400 ;
        RECT 246.000 391.050 247.800 395.400 ;
        RECT 242.400 389.400 247.800 391.050 ;
        RECT 256.800 389.400 258.600 395.400 ;
        RECT 230.400 387.300 231.600 389.400 ;
        RECT 212.850 386.250 216.600 387.300 ;
        RECT 227.850 386.250 231.600 387.300 ;
        RECT 209.100 384.150 210.900 385.950 ;
        RECT 187.950 381.000 190.050 383.100 ;
        RECT 194.100 382.050 195.900 383.850 ;
        RECT 196.950 382.050 199.050 384.150 ;
        RECT 179.100 379.200 180.900 381.000 ;
        RECT 188.100 379.200 189.900 381.000 ;
        RECT 172.800 375.600 176.250 376.800 ;
        RECT 155.700 369.900 162.300 370.800 ;
        RECT 155.700 369.600 157.200 369.900 ;
        RECT 155.400 363.600 157.200 369.600 ;
        RECT 161.400 369.600 162.300 369.900 ;
        RECT 161.400 363.600 163.200 369.600 ;
        RECT 169.200 364.500 171.000 373.800 ;
        RECT 172.800 373.200 174.000 375.600 ;
        RECT 172.200 365.400 174.000 373.200 ;
        RECT 175.200 373.200 183.600 374.100 ;
        RECT 175.200 364.500 177.000 373.200 ;
        RECT 169.200 363.600 177.000 364.500 ;
        RECT 178.800 364.500 180.600 372.300 ;
        RECT 181.800 365.400 183.600 373.200 ;
        RECT 184.800 373.500 192.600 374.400 ;
        RECT 184.800 364.500 186.600 373.500 ;
        RECT 178.800 363.600 186.600 364.500 ;
        RECT 190.800 363.600 192.600 373.500 ;
        RECT 197.400 369.600 198.600 382.050 ;
        RECT 205.950 380.850 208.050 382.950 ;
        RECT 208.950 382.050 211.050 384.150 ;
        RECT 212.850 382.950 214.050 386.250 ;
        RECT 224.100 384.150 225.900 385.950 ;
        RECT 211.950 380.850 214.050 382.950 ;
        RECT 220.950 380.850 223.050 382.950 ;
        RECT 223.950 382.050 226.050 384.150 ;
        RECT 227.850 382.950 229.050 386.250 ;
        RECT 242.400 382.950 243.300 389.400 ;
        RECT 257.400 387.300 258.600 389.400 ;
        RECT 259.800 390.300 261.600 395.400 ;
        RECT 265.800 390.300 267.600 395.400 ;
        RECT 259.800 388.950 267.600 390.300 ;
        RECT 279.000 389.400 280.800 395.400 ;
        RECT 292.800 392.400 294.600 395.400 ;
        RECT 257.400 386.250 261.150 387.300 ;
        RECT 245.100 384.150 246.900 385.950 ;
        RECT 226.950 380.850 229.050 382.950 ;
        RECT 241.950 380.850 244.050 382.950 ;
        RECT 244.950 382.050 247.050 384.150 ;
        RECT 247.950 383.850 250.050 385.950 ;
        RECT 251.100 384.150 252.900 385.950 ;
        RECT 248.100 382.050 249.900 383.850 ;
        RECT 250.950 382.050 253.050 384.150 ;
        RECT 259.950 382.950 261.150 386.250 ;
        RECT 263.100 384.150 264.900 385.950 ;
        RECT 275.250 384.150 277.050 385.950 ;
        RECT 259.950 380.850 262.050 382.950 ;
        RECT 262.950 382.050 265.050 384.150 ;
        RECT 265.950 380.850 268.050 382.950 ;
        RECT 271.950 380.850 274.050 382.950 ;
        RECT 274.950 382.050 277.050 384.150 ;
        RECT 279.000 382.950 280.050 389.400 ;
        RECT 277.950 380.850 280.050 382.950 ;
        RECT 280.950 384.150 282.750 385.950 ;
        RECT 293.400 384.150 294.600 392.400 ;
        RECT 300.150 389.400 301.950 395.400 ;
        RECT 307.950 393.300 309.750 395.400 ;
        RECT 306.000 392.400 309.750 393.300 ;
        RECT 315.750 392.400 317.550 395.400 ;
        RECT 323.550 392.400 325.350 395.400 ;
        RECT 306.000 391.500 307.050 392.400 ;
        RECT 304.950 389.400 307.050 391.500 ;
        RECT 315.750 390.600 316.800 392.400 ;
        RECT 280.950 382.050 283.050 384.150 ;
        RECT 283.950 380.850 286.050 382.950 ;
        RECT 292.950 382.050 295.050 384.150 ;
        RECT 295.950 383.850 298.050 385.950 ;
        RECT 296.100 382.050 297.900 383.850 ;
        RECT 206.100 379.050 207.900 380.850 ;
        RECT 211.950 375.600 213.150 380.850 ;
        RECT 214.950 377.850 217.050 379.950 ;
        RECT 221.100 379.050 222.900 380.850 ;
        RECT 214.950 376.050 216.750 377.850 ;
        RECT 226.950 375.600 228.150 380.850 ;
        RECT 229.950 377.850 232.050 379.950 ;
        RECT 229.950 376.050 231.750 377.850 ;
        RECT 242.400 375.600 243.300 380.850 ;
        RECT 256.950 377.850 259.050 379.950 ;
        RECT 257.250 376.050 259.050 377.850 ;
        RECT 260.850 375.600 262.050 380.850 ;
        RECT 266.100 379.050 267.900 380.850 ;
        RECT 272.100 379.050 273.900 380.850 ;
        RECT 277.950 377.400 278.850 380.850 ;
        RECT 283.950 379.050 285.750 380.850 ;
        RECT 274.800 376.500 278.850 377.400 ;
        RECT 197.400 363.600 199.200 369.600 ;
        RECT 211.500 363.600 213.300 375.600 ;
        RECT 226.500 363.600 228.300 375.600 ;
        RECT 241.800 363.600 243.600 375.600 ;
        RECT 244.800 374.700 252.600 375.600 ;
        RECT 244.800 363.600 246.600 374.700 ;
        RECT 250.800 363.600 252.600 374.700 ;
        RECT 260.700 363.600 262.500 375.600 ;
        RECT 271.800 364.500 273.600 375.600 ;
        RECT 274.800 365.400 276.600 376.500 ;
        RECT 277.800 374.400 285.600 375.300 ;
        RECT 277.800 364.500 279.600 374.400 ;
        RECT 271.800 363.600 279.600 364.500 ;
        RECT 283.800 363.600 285.600 374.400 ;
        RECT 293.400 369.600 294.600 382.050 ;
        RECT 292.800 363.600 294.600 369.600 ;
        RECT 300.150 376.800 301.050 389.400 ;
        RECT 308.550 388.800 310.350 390.600 ;
        RECT 311.850 389.550 316.800 390.600 ;
        RECT 324.300 391.500 325.350 392.400 ;
        RECT 324.300 390.300 328.050 391.500 ;
        RECT 311.850 388.800 313.650 389.550 ;
        RECT 308.850 387.900 309.900 388.800 ;
        RECT 319.050 388.200 320.850 390.000 ;
        RECT 325.950 389.400 328.050 390.300 ;
        RECT 331.650 389.400 333.450 395.400 ;
        RECT 342.000 391.050 343.800 395.400 ;
        RECT 319.050 387.900 319.950 388.200 ;
        RECT 308.850 387.000 319.950 387.900 ;
        RECT 332.250 387.150 333.450 389.400 ;
        RECT 308.850 385.800 309.900 387.000 ;
        RECT 303.000 384.600 309.900 385.800 ;
        RECT 303.000 383.850 303.900 384.600 ;
        RECT 308.100 384.000 309.900 384.600 ;
        RECT 302.100 382.050 303.900 383.850 ;
        RECT 305.100 382.950 306.900 383.700 ;
        RECT 319.050 382.950 319.950 387.000 ;
        RECT 328.950 385.050 333.450 387.150 ;
        RECT 327.150 383.250 331.050 385.050 ;
        RECT 328.950 382.950 331.050 383.250 ;
        RECT 305.100 381.900 313.050 382.950 ;
        RECT 310.950 380.850 313.050 381.900 ;
        RECT 316.950 380.850 319.950 382.950 ;
        RECT 309.450 377.100 311.250 377.400 ;
        RECT 309.450 376.800 317.850 377.100 ;
        RECT 300.150 376.200 317.850 376.800 ;
        RECT 300.150 375.600 311.250 376.200 ;
        RECT 300.150 363.600 301.950 375.600 ;
        RECT 314.250 374.700 316.050 375.300 ;
        RECT 308.550 373.500 316.050 374.700 ;
        RECT 316.950 374.100 317.850 376.200 ;
        RECT 319.050 376.200 319.950 380.850 ;
        RECT 329.250 377.400 331.050 379.200 ;
        RECT 325.950 376.200 330.150 377.400 ;
        RECT 319.050 375.300 325.050 376.200 ;
        RECT 325.950 375.300 328.050 376.200 ;
        RECT 332.250 375.600 333.450 385.050 ;
        RECT 338.400 389.400 343.800 391.050 ;
        RECT 363.000 389.400 364.800 395.400 ;
        RECT 373.800 392.400 375.600 395.400 ;
        RECT 338.400 382.950 339.300 389.400 ;
        RECT 341.100 384.150 342.900 385.950 ;
        RECT 337.950 380.850 340.050 382.950 ;
        RECT 340.950 382.050 343.050 384.150 ;
        RECT 343.950 383.850 346.050 385.950 ;
        RECT 347.100 384.150 348.900 385.950 ;
        RECT 359.250 384.150 361.050 385.950 ;
        RECT 344.100 382.050 345.900 383.850 ;
        RECT 346.950 382.050 349.050 384.150 ;
        RECT 355.950 380.850 358.050 382.950 ;
        RECT 358.950 382.050 361.050 384.150 ;
        RECT 363.000 382.950 364.050 389.400 ;
        RECT 361.950 380.850 364.050 382.950 ;
        RECT 364.950 384.150 366.750 385.950 ;
        RECT 374.400 384.150 375.600 392.400 ;
        RECT 380.550 389.400 382.350 395.400 ;
        RECT 388.650 392.400 390.450 395.400 ;
        RECT 396.450 392.400 398.250 395.400 ;
        RECT 404.250 393.300 406.050 395.400 ;
        RECT 404.250 392.400 408.000 393.300 ;
        RECT 388.650 391.500 389.700 392.400 ;
        RECT 385.950 390.300 389.700 391.500 ;
        RECT 397.200 390.600 398.250 392.400 ;
        RECT 406.950 391.500 408.000 392.400 ;
        RECT 385.950 389.400 388.050 390.300 ;
        RECT 380.550 387.150 381.750 389.400 ;
        RECT 393.150 388.200 394.950 390.000 ;
        RECT 397.200 389.550 402.150 390.600 ;
        RECT 400.350 388.800 402.150 389.550 ;
        RECT 403.650 388.800 405.450 390.600 ;
        RECT 406.950 389.400 409.050 391.500 ;
        RECT 412.050 389.400 413.850 395.400 ;
        RECT 394.050 387.900 394.950 388.200 ;
        RECT 404.100 387.900 405.150 388.800 ;
        RECT 364.950 382.050 367.050 384.150 ;
        RECT 367.950 380.850 370.050 382.950 ;
        RECT 373.950 382.050 376.050 384.150 ;
        RECT 376.950 383.850 379.050 385.950 ;
        RECT 380.550 385.050 385.050 387.150 ;
        RECT 394.050 387.000 405.150 387.900 ;
        RECT 377.100 382.050 378.900 383.850 ;
        RECT 338.400 375.600 339.300 380.850 ;
        RECT 356.100 379.050 357.900 380.850 ;
        RECT 361.950 377.400 362.850 380.850 ;
        RECT 367.950 379.050 369.750 380.850 ;
        RECT 358.800 376.500 362.850 377.400 ;
        RECT 324.150 374.400 325.050 375.300 ;
        RECT 321.450 374.100 323.250 374.400 ;
        RECT 308.550 372.600 309.750 373.500 ;
        RECT 316.950 373.200 323.250 374.100 ;
        RECT 321.450 372.600 323.250 373.200 ;
        RECT 324.150 372.600 326.850 374.400 ;
        RECT 304.950 370.500 309.750 372.600 ;
        RECT 312.450 371.550 314.250 372.300 ;
        RECT 317.250 371.550 319.050 372.300 ;
        RECT 312.450 370.500 319.050 371.550 ;
        RECT 308.550 369.600 309.750 370.500 ;
        RECT 308.550 363.600 310.350 369.600 ;
        RECT 316.350 363.600 318.150 370.500 ;
        RECT 324.150 369.600 328.050 371.700 ;
        RECT 324.150 363.600 325.950 369.600 ;
        RECT 331.650 363.600 333.450 375.600 ;
        RECT 337.800 363.600 339.600 375.600 ;
        RECT 340.800 374.700 348.600 375.600 ;
        RECT 340.800 363.600 342.600 374.700 ;
        RECT 346.800 363.600 348.600 374.700 ;
        RECT 355.800 364.500 357.600 375.600 ;
        RECT 358.800 365.400 360.600 376.500 ;
        RECT 361.800 374.400 369.600 375.300 ;
        RECT 361.800 364.500 363.600 374.400 ;
        RECT 355.800 363.600 363.600 364.500 ;
        RECT 367.800 363.600 369.600 374.400 ;
        RECT 374.400 369.600 375.600 382.050 ;
        RECT 373.800 363.600 375.600 369.600 ;
        RECT 380.550 375.600 381.750 385.050 ;
        RECT 382.950 383.250 386.850 385.050 ;
        RECT 382.950 382.950 385.050 383.250 ;
        RECT 394.050 382.950 394.950 387.000 ;
        RECT 404.100 385.800 405.150 387.000 ;
        RECT 404.100 384.600 411.000 385.800 ;
        RECT 404.100 384.000 405.900 384.600 ;
        RECT 410.100 383.850 411.000 384.600 ;
        RECT 407.100 382.950 408.900 383.700 ;
        RECT 394.050 380.850 397.050 382.950 ;
        RECT 400.950 381.900 408.900 382.950 ;
        RECT 410.100 382.050 411.900 383.850 ;
        RECT 400.950 380.850 403.050 381.900 ;
        RECT 382.950 377.400 384.750 379.200 ;
        RECT 383.850 376.200 388.050 377.400 ;
        RECT 394.050 376.200 394.950 380.850 ;
        RECT 402.750 377.100 404.550 377.400 ;
        RECT 380.550 363.600 382.350 375.600 ;
        RECT 385.950 375.300 388.050 376.200 ;
        RECT 388.950 375.300 394.950 376.200 ;
        RECT 396.150 376.800 404.550 377.100 ;
        RECT 412.950 376.800 413.850 389.400 ;
        RECT 396.150 376.200 413.850 376.800 ;
        RECT 388.950 374.400 389.850 375.300 ;
        RECT 387.150 372.600 389.850 374.400 ;
        RECT 390.750 374.100 392.550 374.400 ;
        RECT 396.150 374.100 397.050 376.200 ;
        RECT 402.750 375.600 413.850 376.200 ;
        RECT 390.750 373.200 397.050 374.100 ;
        RECT 397.950 374.700 399.750 375.300 ;
        RECT 397.950 373.500 405.450 374.700 ;
        RECT 390.750 372.600 392.550 373.200 ;
        RECT 404.250 372.600 405.450 373.500 ;
        RECT 385.950 369.600 389.850 371.700 ;
        RECT 394.950 371.550 396.750 372.300 ;
        RECT 399.750 371.550 401.550 372.300 ;
        RECT 394.950 370.500 401.550 371.550 ;
        RECT 404.250 370.500 409.050 372.600 ;
        RECT 388.050 363.600 389.850 369.600 ;
        RECT 395.850 363.600 397.650 370.500 ;
        RECT 404.250 369.600 405.450 370.500 ;
        RECT 403.650 363.600 405.450 369.600 ;
        RECT 412.050 363.600 413.850 375.600 ;
        RECT 416.550 389.400 418.350 395.400 ;
        RECT 424.650 392.400 426.450 395.400 ;
        RECT 432.450 392.400 434.250 395.400 ;
        RECT 440.250 393.300 442.050 395.400 ;
        RECT 440.250 392.400 444.000 393.300 ;
        RECT 424.650 391.500 425.700 392.400 ;
        RECT 421.950 390.300 425.700 391.500 ;
        RECT 433.200 390.600 434.250 392.400 ;
        RECT 442.950 391.500 444.000 392.400 ;
        RECT 421.950 389.400 424.050 390.300 ;
        RECT 416.550 387.150 417.750 389.400 ;
        RECT 429.150 388.200 430.950 390.000 ;
        RECT 433.200 389.550 438.150 390.600 ;
        RECT 436.350 388.800 438.150 389.550 ;
        RECT 439.650 388.800 441.450 390.600 ;
        RECT 442.950 389.400 445.050 391.500 ;
        RECT 448.050 389.400 449.850 395.400 ;
        RECT 454.800 389.400 456.600 395.400 ;
        RECT 430.050 387.900 430.950 388.200 ;
        RECT 440.100 387.900 441.150 388.800 ;
        RECT 416.550 385.050 421.050 387.150 ;
        RECT 430.050 387.000 441.150 387.900 ;
        RECT 416.550 375.600 417.750 385.050 ;
        RECT 418.950 383.250 422.850 385.050 ;
        RECT 418.950 382.950 421.050 383.250 ;
        RECT 430.050 382.950 430.950 387.000 ;
        RECT 440.100 385.800 441.150 387.000 ;
        RECT 440.100 384.600 447.000 385.800 ;
        RECT 440.100 384.000 441.900 384.600 ;
        RECT 446.100 383.850 447.000 384.600 ;
        RECT 443.100 382.950 444.900 383.700 ;
        RECT 430.050 380.850 433.050 382.950 ;
        RECT 436.950 381.900 444.900 382.950 ;
        RECT 446.100 382.050 447.900 383.850 ;
        RECT 436.950 380.850 439.050 381.900 ;
        RECT 418.950 377.400 420.750 379.200 ;
        RECT 419.850 376.200 424.050 377.400 ;
        RECT 430.050 376.200 430.950 380.850 ;
        RECT 438.750 377.100 440.550 377.400 ;
        RECT 416.550 363.600 418.350 375.600 ;
        RECT 421.950 375.300 424.050 376.200 ;
        RECT 424.950 375.300 430.950 376.200 ;
        RECT 432.150 376.800 440.550 377.100 ;
        RECT 448.950 376.800 449.850 389.400 ;
        RECT 455.400 387.300 456.600 389.400 ;
        RECT 457.800 390.300 459.600 395.400 ;
        RECT 463.800 390.300 465.600 395.400 ;
        RECT 474.000 391.050 475.800 395.400 ;
        RECT 457.800 388.950 465.600 390.300 ;
        RECT 470.400 389.400 475.800 391.050 ;
        RECT 455.400 386.250 459.150 387.300 ;
        RECT 457.950 382.950 459.150 386.250 ;
        RECT 461.100 384.150 462.900 385.950 ;
        RECT 457.950 380.850 460.050 382.950 ;
        RECT 460.950 382.050 463.050 384.150 ;
        RECT 470.400 382.950 471.300 389.400 ;
        RECT 488.100 387.000 489.900 395.400 ;
        RECT 503.400 392.400 505.200 395.400 ;
        RECT 473.100 384.150 474.900 385.950 ;
        RECT 463.950 380.850 466.050 382.950 ;
        RECT 469.950 380.850 472.050 382.950 ;
        RECT 472.950 382.050 475.050 384.150 ;
        RECT 475.950 383.850 478.050 385.950 ;
        RECT 479.100 384.150 480.900 385.950 ;
        RECT 488.100 385.350 492.300 387.000 ;
        RECT 476.100 382.050 477.900 383.850 ;
        RECT 478.950 382.050 481.050 384.150 ;
        RECT 491.400 381.150 492.300 385.350 ;
        RECT 499.950 383.850 502.050 385.950 ;
        RECT 503.400 384.150 504.600 392.400 ;
        RECT 512.400 387.900 514.200 395.400 ;
        RECT 519.900 390.900 521.700 395.400 ;
        RECT 529.800 392.400 531.600 395.400 ;
        RECT 519.900 389.400 523.050 390.900 ;
        RECT 518.100 387.900 519.900 388.500 ;
        RECT 512.400 386.700 519.900 387.900 ;
        RECT 500.100 382.050 501.900 383.850 ;
        RECT 502.950 382.050 505.050 384.150 ;
        RECT 454.950 377.850 457.050 379.950 ;
        RECT 432.150 376.200 449.850 376.800 ;
        RECT 424.950 374.400 425.850 375.300 ;
        RECT 423.150 372.600 425.850 374.400 ;
        RECT 426.750 374.100 428.550 374.400 ;
        RECT 432.150 374.100 433.050 376.200 ;
        RECT 438.750 375.600 449.850 376.200 ;
        RECT 455.250 376.050 457.050 377.850 ;
        RECT 458.850 375.600 460.050 380.850 ;
        RECT 464.100 379.050 465.900 380.850 ;
        RECT 470.400 375.600 471.300 380.850 ;
        RECT 481.950 377.850 484.050 379.950 ;
        RECT 487.950 377.850 490.050 379.950 ;
        RECT 490.950 379.050 493.050 381.150 ;
        RECT 482.100 376.050 483.900 377.850 ;
        RECT 426.750 373.200 433.050 374.100 ;
        RECT 433.950 374.700 435.750 375.300 ;
        RECT 433.950 373.500 441.450 374.700 ;
        RECT 426.750 372.600 428.550 373.200 ;
        RECT 440.250 372.600 441.450 373.500 ;
        RECT 421.950 369.600 425.850 371.700 ;
        RECT 430.950 371.550 432.750 372.300 ;
        RECT 435.750 371.550 437.550 372.300 ;
        RECT 430.950 370.500 437.550 371.550 ;
        RECT 440.250 370.500 445.050 372.600 ;
        RECT 424.050 363.600 425.850 369.600 ;
        RECT 431.850 363.600 433.650 370.500 ;
        RECT 440.250 369.600 441.450 370.500 ;
        RECT 439.650 363.600 441.450 369.600 ;
        RECT 448.050 363.600 449.850 375.600 ;
        RECT 458.700 363.600 460.500 375.600 ;
        RECT 469.800 363.600 471.600 375.600 ;
        RECT 472.800 374.700 480.600 375.600 ;
        RECT 484.950 374.850 487.050 376.950 ;
        RECT 488.250 376.050 490.050 377.850 ;
        RECT 472.800 363.600 474.600 374.700 ;
        RECT 478.800 363.600 480.600 374.700 ;
        RECT 485.100 373.050 486.900 374.850 ;
        RECT 491.400 370.800 492.300 379.050 ;
        RECT 485.700 369.900 492.300 370.800 ;
        RECT 485.700 369.600 487.200 369.900 ;
        RECT 485.400 363.600 487.200 369.600 ;
        RECT 491.400 369.600 492.300 369.900 ;
        RECT 503.400 369.600 504.600 382.050 ;
        RECT 511.950 380.850 514.050 382.950 ;
        RECT 512.100 379.050 513.900 380.850 ;
        RECT 515.550 369.600 516.600 386.700 ;
        RECT 522.000 382.950 523.050 389.400 ;
        RECT 530.400 384.150 531.600 392.400 ;
        RECT 542.100 387.000 543.900 395.400 ;
        RECT 560.100 387.000 561.900 395.400 ;
        RECT 571.800 389.400 573.600 395.400 ;
        RECT 518.100 381.150 519.900 382.950 ;
        RECT 517.950 379.050 520.050 381.150 ;
        RECT 520.950 380.850 523.050 382.950 ;
        RECT 529.950 382.050 532.050 384.150 ;
        RECT 532.950 383.850 535.050 385.950 ;
        RECT 539.700 385.350 543.900 387.000 ;
        RECT 557.700 385.350 561.900 387.000 ;
        RECT 572.400 387.300 573.600 389.400 ;
        RECT 574.800 390.300 576.600 395.400 ;
        RECT 580.800 390.300 582.600 395.400 ;
        RECT 574.800 388.950 582.600 390.300 ;
        RECT 587.400 390.300 589.200 395.400 ;
        RECT 593.400 390.300 595.200 395.400 ;
        RECT 587.400 388.950 595.200 390.300 ;
        RECT 596.400 389.400 598.200 395.400 ;
        RECT 605.400 392.400 607.200 395.400 ;
        RECT 596.400 387.300 597.600 389.400 ;
        RECT 572.400 386.250 576.150 387.300 ;
        RECT 533.100 382.050 534.900 383.850 ;
        RECT 522.000 375.600 523.050 380.850 ;
        RECT 491.400 363.600 493.200 369.600 ;
        RECT 503.400 363.600 505.200 369.600 ;
        RECT 515.400 363.600 517.200 369.600 ;
        RECT 522.000 363.600 523.800 375.600 ;
        RECT 530.400 369.600 531.600 382.050 ;
        RECT 539.700 381.150 540.600 385.350 ;
        RECT 557.700 381.150 558.600 385.350 ;
        RECT 574.950 382.950 576.150 386.250 ;
        RECT 593.850 386.250 597.600 387.300 ;
        RECT 578.100 384.150 579.900 385.950 ;
        RECT 590.100 384.150 591.900 385.950 ;
        RECT 538.950 379.050 541.050 381.150 ;
        RECT 539.700 370.800 540.600 379.050 ;
        RECT 541.950 377.850 544.050 379.950 ;
        RECT 547.950 377.850 550.050 379.950 ;
        RECT 556.950 379.050 559.050 381.150 ;
        RECT 574.950 380.850 577.050 382.950 ;
        RECT 577.950 382.050 580.050 384.150 ;
        RECT 580.950 380.850 583.050 382.950 ;
        RECT 586.950 380.850 589.050 382.950 ;
        RECT 589.950 382.050 592.050 384.150 ;
        RECT 593.850 382.950 595.050 386.250 ;
        RECT 601.950 383.850 604.050 385.950 ;
        RECT 605.400 384.150 606.600 392.400 ;
        RECT 617.100 387.000 618.900 395.400 ;
        RECT 614.700 385.350 618.900 387.000 ;
        RECT 632.100 387.000 633.900 395.400 ;
        RECT 647.100 387.000 648.900 395.400 ;
        RECT 658.800 392.400 660.600 395.400 ;
        RECT 632.100 385.350 636.300 387.000 ;
        RECT 592.950 380.850 595.050 382.950 ;
        RECT 602.100 382.050 603.900 383.850 ;
        RECT 604.950 382.050 607.050 384.150 ;
        RECT 541.950 376.050 543.750 377.850 ;
        RECT 544.950 374.850 547.050 376.950 ;
        RECT 548.100 376.050 549.900 377.850 ;
        RECT 545.100 373.050 546.900 374.850 ;
        RECT 557.700 370.800 558.600 379.050 ;
        RECT 559.950 377.850 562.050 379.950 ;
        RECT 565.950 377.850 568.050 379.950 ;
        RECT 571.950 377.850 574.050 379.950 ;
        RECT 559.950 376.050 561.750 377.850 ;
        RECT 562.950 374.850 565.050 376.950 ;
        RECT 566.100 376.050 567.900 377.850 ;
        RECT 572.250 376.050 574.050 377.850 ;
        RECT 575.850 375.600 577.050 380.850 ;
        RECT 581.100 379.050 582.900 380.850 ;
        RECT 587.100 379.050 588.900 380.850 ;
        RECT 592.950 375.600 594.150 380.850 ;
        RECT 595.950 377.850 598.050 379.950 ;
        RECT 595.950 376.050 597.750 377.850 ;
        RECT 563.100 373.050 564.900 374.850 ;
        RECT 539.700 369.900 546.300 370.800 ;
        RECT 539.700 369.600 540.600 369.900 ;
        RECT 529.800 363.600 531.600 369.600 ;
        RECT 538.800 363.600 540.600 369.600 ;
        RECT 544.800 369.600 546.300 369.900 ;
        RECT 557.700 369.900 564.300 370.800 ;
        RECT 557.700 369.600 558.600 369.900 ;
        RECT 544.800 363.600 546.600 369.600 ;
        RECT 556.800 363.600 558.600 369.600 ;
        RECT 562.800 369.600 564.300 369.900 ;
        RECT 562.800 363.600 564.600 369.600 ;
        RECT 575.700 363.600 577.500 375.600 ;
        RECT 592.500 363.600 594.300 375.600 ;
        RECT 605.400 369.600 606.600 382.050 ;
        RECT 614.700 381.150 615.600 385.350 ;
        RECT 635.400 381.150 636.300 385.350 ;
        RECT 644.700 385.350 648.900 387.000 ;
        RECT 644.700 381.150 645.600 385.350 ;
        RECT 652.950 384.450 655.050 385.050 ;
        RECT 650.550 383.550 655.050 384.450 ;
        RECT 659.400 384.150 660.600 392.400 ;
        RECT 667.800 389.400 669.600 395.400 ;
        RECT 668.400 387.300 669.600 389.400 ;
        RECT 670.800 390.300 672.600 395.400 ;
        RECT 676.800 390.300 678.600 395.400 ;
        RECT 690.000 391.050 691.800 395.400 ;
        RECT 670.800 388.950 678.600 390.300 ;
        RECT 686.400 389.400 691.800 391.050 ;
        RECT 700.950 390.450 703.050 391.050 ;
        RECT 698.550 389.550 703.050 390.450 ;
        RECT 668.400 386.250 672.150 387.300 ;
        RECT 650.550 382.050 651.450 383.550 ;
        RECT 652.950 382.950 655.050 383.550 ;
        RECT 658.950 382.050 661.050 384.150 ;
        RECT 661.950 383.850 664.050 385.950 ;
        RECT 662.100 382.050 663.900 383.850 ;
        RECT 670.950 382.950 672.150 386.250 ;
        RECT 674.100 384.150 675.900 385.950 ;
        RECT 613.950 379.050 616.050 381.150 ;
        RECT 614.700 370.800 615.600 379.050 ;
        RECT 616.950 377.850 619.050 379.950 ;
        RECT 622.950 377.850 625.050 379.950 ;
        RECT 625.950 377.850 628.050 379.950 ;
        RECT 631.950 377.850 634.050 379.950 ;
        RECT 634.950 379.050 637.050 381.150 ;
        RECT 643.950 379.050 646.050 381.150 ;
        RECT 649.950 379.950 652.050 382.050 ;
        RECT 616.950 376.050 618.750 377.850 ;
        RECT 619.950 374.850 622.050 376.950 ;
        RECT 623.100 376.050 624.900 377.850 ;
        RECT 626.100 376.050 627.900 377.850 ;
        RECT 628.950 374.850 631.050 376.950 ;
        RECT 632.250 376.050 634.050 377.850 ;
        RECT 620.100 373.050 621.900 374.850 ;
        RECT 629.100 373.050 630.900 374.850 ;
        RECT 635.400 370.800 636.300 379.050 ;
        RECT 614.700 369.900 621.300 370.800 ;
        RECT 614.700 369.600 615.600 369.900 ;
        RECT 605.400 363.600 607.200 369.600 ;
        RECT 613.800 363.600 615.600 369.600 ;
        RECT 619.800 369.600 621.300 369.900 ;
        RECT 629.700 369.900 636.300 370.800 ;
        RECT 629.700 369.600 631.200 369.900 ;
        RECT 619.800 363.600 621.600 369.600 ;
        RECT 629.400 363.600 631.200 369.600 ;
        RECT 635.400 369.600 636.300 369.900 ;
        RECT 644.700 370.800 645.600 379.050 ;
        RECT 646.950 377.850 649.050 379.950 ;
        RECT 652.950 377.850 655.050 379.950 ;
        RECT 646.950 376.050 648.750 377.850 ;
        RECT 649.950 374.850 652.050 376.950 ;
        RECT 653.100 376.050 654.900 377.850 ;
        RECT 650.100 373.050 651.900 374.850 ;
        RECT 644.700 369.900 651.300 370.800 ;
        RECT 644.700 369.600 645.600 369.900 ;
        RECT 635.400 363.600 637.200 369.600 ;
        RECT 643.800 363.600 645.600 369.600 ;
        RECT 649.800 369.600 651.300 369.900 ;
        RECT 659.400 369.600 660.600 382.050 ;
        RECT 670.950 380.850 673.050 382.950 ;
        RECT 673.950 382.050 676.050 384.150 ;
        RECT 686.400 382.950 687.300 389.400 ;
        RECT 689.100 384.150 690.900 385.950 ;
        RECT 676.950 380.850 679.050 382.950 ;
        RECT 685.950 380.850 688.050 382.950 ;
        RECT 688.950 382.050 691.050 384.150 ;
        RECT 691.950 383.850 694.050 385.950 ;
        RECT 695.100 384.150 696.900 385.950 ;
        RECT 692.100 382.050 693.900 383.850 ;
        RECT 694.950 382.050 697.050 384.150 ;
        RECT 667.950 377.850 670.050 379.950 ;
        RECT 668.250 376.050 670.050 377.850 ;
        RECT 671.850 375.600 673.050 380.850 ;
        RECT 677.100 379.050 678.900 380.850 ;
        RECT 686.400 375.600 687.300 380.850 ;
        RECT 691.950 378.450 694.050 379.050 ;
        RECT 698.550 378.450 699.450 389.550 ;
        RECT 700.950 388.950 703.050 389.550 ;
        RECT 704.100 387.000 705.900 395.400 ;
        RECT 716.400 390.300 718.200 395.400 ;
        RECT 722.400 390.300 724.200 395.400 ;
        RECT 716.400 388.950 724.200 390.300 ;
        RECT 725.400 389.400 727.200 395.400 ;
        RECT 733.800 392.400 735.600 395.400 ;
        RECT 725.400 387.300 726.600 389.400 ;
        RECT 701.700 385.350 705.900 387.000 ;
        RECT 722.850 386.250 726.600 387.300 ;
        RECT 701.700 381.150 702.600 385.350 ;
        RECT 706.950 384.450 709.050 385.050 ;
        RECT 706.950 383.550 714.450 384.450 ;
        RECT 719.100 384.150 720.900 385.950 ;
        RECT 706.950 382.950 709.050 383.550 ;
        RECT 700.950 379.050 703.050 381.150 ;
        RECT 691.950 377.550 699.450 378.450 ;
        RECT 691.950 376.950 694.050 377.550 ;
        RECT 649.800 363.600 651.600 369.600 ;
        RECT 658.800 363.600 660.600 369.600 ;
        RECT 671.700 363.600 673.500 375.600 ;
        RECT 685.800 363.600 687.600 375.600 ;
        RECT 688.800 374.700 696.600 375.600 ;
        RECT 688.800 363.600 690.600 374.700 ;
        RECT 694.800 363.600 696.600 374.700 ;
        RECT 701.700 370.800 702.600 379.050 ;
        RECT 703.950 377.850 706.050 379.950 ;
        RECT 709.950 377.850 712.050 379.950 ;
        RECT 703.950 376.050 705.750 377.850 ;
        RECT 706.950 374.850 709.050 376.950 ;
        RECT 710.100 376.050 711.900 377.850 ;
        RECT 707.100 373.050 708.900 374.850 ;
        RECT 709.950 372.450 712.050 373.050 ;
        RECT 713.550 372.450 714.450 383.550 ;
        RECT 715.950 380.850 718.050 382.950 ;
        RECT 718.950 382.050 721.050 384.150 ;
        RECT 722.850 382.950 724.050 386.250 ;
        RECT 734.400 384.150 735.600 392.400 ;
        RECT 740.400 390.300 742.200 395.400 ;
        RECT 746.400 390.300 748.200 395.400 ;
        RECT 740.400 388.950 748.200 390.300 ;
        RECT 749.400 389.400 751.200 395.400 ;
        RECT 749.400 387.300 750.600 389.400 ;
        RECT 746.850 386.250 750.600 387.300 ;
        RECT 721.950 380.850 724.050 382.950 ;
        RECT 733.950 382.050 736.050 384.150 ;
        RECT 736.950 383.850 739.050 385.950 ;
        RECT 743.100 384.150 744.900 385.950 ;
        RECT 737.100 382.050 738.900 383.850 ;
        RECT 716.100 379.050 717.900 380.850 ;
        RECT 721.950 375.600 723.150 380.850 ;
        RECT 724.950 377.850 727.050 379.950 ;
        RECT 724.950 376.050 726.750 377.850 ;
        RECT 709.950 371.550 714.450 372.450 ;
        RECT 709.950 370.950 712.050 371.550 ;
        RECT 701.700 369.900 708.300 370.800 ;
        RECT 701.700 369.600 702.600 369.900 ;
        RECT 700.800 363.600 702.600 369.600 ;
        RECT 706.800 369.600 708.300 369.900 ;
        RECT 706.800 363.600 708.600 369.600 ;
        RECT 721.500 363.600 723.300 375.600 ;
        RECT 734.400 369.600 735.600 382.050 ;
        RECT 739.950 380.850 742.050 382.950 ;
        RECT 742.950 382.050 745.050 384.150 ;
        RECT 746.850 382.950 748.050 386.250 ;
        RECT 748.950 384.450 751.050 385.050 ;
        RECT 757.950 384.450 760.050 385.050 ;
        RECT 748.950 383.550 760.050 384.450 ;
        RECT 748.950 382.950 751.050 383.550 ;
        RECT 757.950 382.950 760.050 383.550 ;
        RECT 745.950 380.850 748.050 382.950 ;
        RECT 740.100 379.050 741.900 380.850 ;
        RECT 745.950 375.600 747.150 380.850 ;
        RECT 748.950 377.850 751.050 379.950 ;
        RECT 748.950 376.050 750.750 377.850 ;
        RECT 733.800 363.600 735.600 369.600 ;
        RECT 745.500 363.600 747.300 375.600 ;
        RECT 7.800 353.400 9.600 359.400 ;
        RECT 8.400 340.950 9.600 353.400 ;
        RECT 19.500 347.400 21.300 359.400 ;
        RECT 33.300 348.900 35.100 359.400 ;
        RECT 32.700 347.550 35.100 348.900 ;
        RECT 14.100 342.150 15.900 343.950 ;
        RECT 19.950 342.150 21.150 347.400 ;
        RECT 22.950 345.150 24.750 346.950 ;
        RECT 22.950 343.050 25.050 345.150 ;
        RECT 7.950 338.850 10.050 340.950 ;
        RECT 11.100 339.150 12.900 340.950 ;
        RECT 13.950 340.050 16.050 342.150 ;
        RECT 8.400 330.600 9.600 338.850 ;
        RECT 10.950 337.050 13.050 339.150 ;
        RECT 16.950 338.850 19.050 340.950 ;
        RECT 19.950 340.050 22.050 342.150 ;
        RECT 32.700 340.950 34.050 347.550 ;
        RECT 40.800 347.400 42.600 359.400 ;
        RECT 50.400 353.400 52.200 359.400 ;
        RECT 17.100 337.050 18.900 338.850 ;
        RECT 20.850 336.750 22.050 340.050 ;
        RECT 31.950 338.850 34.050 340.950 ;
        RECT 35.400 346.200 37.200 346.650 ;
        RECT 41.400 346.200 42.600 347.400 ;
        RECT 35.400 345.000 42.600 346.200 ;
        RECT 35.400 344.850 37.200 345.000 ;
        RECT 20.850 335.700 24.600 336.750 ;
        RECT 7.800 327.600 9.600 330.600 ;
        RECT 14.400 332.700 22.200 334.050 ;
        RECT 14.400 327.600 16.200 332.700 ;
        RECT 20.400 327.600 22.200 332.700 ;
        RECT 23.400 333.600 24.600 335.700 ;
        RECT 31.950 333.600 33.000 338.850 ;
        RECT 35.400 336.600 36.300 344.850 ;
        RECT 38.100 342.150 39.900 343.950 ;
        RECT 47.100 342.150 48.900 343.950 ;
        RECT 37.950 340.050 40.050 342.150 ;
        RECT 41.100 339.150 42.900 340.950 ;
        RECT 46.950 340.050 49.050 342.150 ;
        RECT 40.950 337.050 43.050 339.150 ;
        RECT 35.250 335.700 37.050 336.600 ;
        RECT 50.550 336.300 51.600 353.400 ;
        RECT 57.000 347.400 58.800 359.400 ;
        RECT 65.400 353.400 67.200 359.400 ;
        RECT 65.700 353.100 67.200 353.400 ;
        RECT 71.400 353.400 73.200 359.400 ;
        RECT 80.400 353.400 82.200 359.400 ;
        RECT 71.400 353.100 72.300 353.400 ;
        RECT 65.700 352.200 72.300 353.100 ;
        RECT 80.700 353.100 82.200 353.400 ;
        RECT 86.400 353.400 88.200 359.400 ;
        RECT 86.400 353.100 87.300 353.400 ;
        RECT 80.700 352.200 87.300 353.100 ;
        RECT 65.100 348.150 66.900 349.950 ;
        RECT 52.950 341.850 55.050 343.950 ;
        RECT 57.000 342.150 58.050 347.400 ;
        RECT 62.100 345.150 63.900 346.950 ;
        RECT 64.950 346.050 67.050 348.150 ;
        RECT 68.250 345.150 70.050 346.950 ;
        RECT 61.950 343.050 64.050 345.150 ;
        RECT 67.950 343.050 70.050 345.150 ;
        RECT 71.400 343.950 72.300 352.200 ;
        RECT 80.100 348.150 81.900 349.950 ;
        RECT 77.100 345.150 78.900 346.950 ;
        RECT 79.950 346.050 82.050 348.150 ;
        RECT 83.250 345.150 85.050 346.950 ;
        RECT 53.100 340.050 54.900 341.850 ;
        RECT 55.950 340.050 58.050 342.150 ;
        RECT 70.950 341.850 73.050 343.950 ;
        RECT 76.950 343.050 79.050 345.150 ;
        RECT 82.950 343.050 85.050 345.150 ;
        RECT 86.400 343.950 87.300 352.200 ;
        RECT 97.500 347.400 99.300 359.400 ;
        RECT 112.800 353.400 114.600 359.400 ;
        RECT 113.700 353.100 114.600 353.400 ;
        RECT 118.800 353.400 120.600 359.400 ;
        RECT 128.400 353.400 130.200 359.400 ;
        RECT 118.800 353.100 120.300 353.400 ;
        RECT 113.700 352.200 120.300 353.100 ;
        RECT 85.950 341.850 88.050 343.950 ;
        RECT 92.100 342.150 93.900 343.950 ;
        RECT 97.950 342.150 99.150 347.400 ;
        RECT 100.950 345.150 102.750 346.950 ;
        RECT 100.950 343.050 103.050 345.150 ;
        RECT 113.700 343.950 114.600 352.200 ;
        RECT 119.100 348.150 120.900 349.950 ;
        RECT 115.950 345.150 117.750 346.950 ;
        RECT 118.950 346.050 121.050 348.150 ;
        RECT 122.100 345.150 123.900 346.950 ;
        RECT 35.250 334.800 38.700 335.700 ;
        RECT 23.400 327.600 25.200 333.600 ;
        RECT 31.800 327.600 33.600 333.600 ;
        RECT 37.800 330.600 38.700 334.800 ;
        RECT 47.400 335.100 54.900 336.300 ;
        RECT 37.800 327.600 39.600 330.600 ;
        RECT 47.400 327.600 49.200 335.100 ;
        RECT 53.100 334.500 54.900 335.100 ;
        RECT 57.000 333.600 58.050 340.050 ;
        RECT 71.400 337.650 72.300 341.850 ;
        RECT 86.400 337.650 87.300 341.850 ;
        RECT 91.950 340.050 94.050 342.150 ;
        RECT 94.950 338.850 97.050 340.950 ;
        RECT 97.950 340.050 100.050 342.150 ;
        RECT 112.950 341.850 115.050 343.950 ;
        RECT 115.950 343.050 118.050 345.150 ;
        RECT 121.950 343.050 124.050 345.150 ;
        RECT 54.900 332.100 58.050 333.600 ;
        RECT 68.100 336.000 72.300 337.650 ;
        RECT 83.100 336.000 87.300 337.650 ;
        RECT 95.100 337.050 96.900 338.850 ;
        RECT 98.850 336.750 100.050 340.050 ;
        RECT 113.700 337.650 114.600 341.850 ;
        RECT 128.400 340.950 129.600 353.400 ;
        RECT 134.400 348.300 136.200 359.400 ;
        RECT 140.400 348.300 142.200 359.400 ;
        RECT 134.400 347.400 142.200 348.300 ;
        RECT 143.400 347.400 145.200 359.400 ;
        RECT 154.500 347.400 156.300 359.400 ;
        RECT 169.800 353.400 171.600 359.400 ;
        RECT 143.700 342.150 144.600 347.400 ;
        RECT 149.100 342.150 150.900 343.950 ;
        RECT 154.950 342.150 156.150 347.400 ;
        RECT 157.950 345.150 159.750 346.950 ;
        RECT 157.950 343.050 160.050 345.150 ;
        RECT 125.100 339.150 126.900 340.950 ;
        RECT 54.900 327.600 56.700 332.100 ;
        RECT 68.100 327.600 69.900 336.000 ;
        RECT 83.100 327.600 84.900 336.000 ;
        RECT 98.850 335.700 102.600 336.750 ;
        RECT 113.700 336.000 117.900 337.650 ;
        RECT 124.950 337.050 127.050 339.150 ;
        RECT 127.950 338.850 130.050 340.950 ;
        RECT 133.950 338.850 136.050 340.950 ;
        RECT 137.100 339.150 138.900 340.950 ;
        RECT 92.400 332.700 100.200 334.050 ;
        RECT 92.400 327.600 94.200 332.700 ;
        RECT 98.400 327.600 100.200 332.700 ;
        RECT 101.400 333.600 102.600 335.700 ;
        RECT 101.400 327.600 103.200 333.600 ;
        RECT 116.100 327.600 117.900 336.000 ;
        RECT 128.400 330.600 129.600 338.850 ;
        RECT 134.100 337.050 135.900 338.850 ;
        RECT 136.950 337.050 139.050 339.150 ;
        RECT 139.950 338.850 142.050 340.950 ;
        RECT 142.950 340.050 145.050 342.150 ;
        RECT 148.950 340.050 151.050 342.150 ;
        RECT 140.100 337.050 141.900 338.850 ;
        RECT 143.700 333.600 144.600 340.050 ;
        RECT 151.950 338.850 154.050 340.950 ;
        RECT 154.950 340.050 157.050 342.150 ;
        RECT 170.400 340.950 171.600 353.400 ;
        RECT 183.600 347.400 185.400 359.400 ;
        RECT 193.800 353.400 195.600 359.400 ;
        RECT 183.600 346.350 186.000 347.400 ;
        RECT 182.100 342.150 183.900 343.950 ;
        RECT 152.100 337.050 153.900 338.850 ;
        RECT 155.850 336.750 157.050 340.050 ;
        RECT 169.950 338.850 172.050 340.950 ;
        RECT 173.100 339.150 174.900 340.950 ;
        RECT 181.950 340.050 184.050 342.150 ;
        RECT 184.950 339.150 186.000 346.350 ;
        RECT 188.100 342.150 189.900 343.950 ;
        RECT 187.950 340.050 190.050 342.150 ;
        RECT 194.400 340.950 195.600 353.400 ;
        RECT 202.800 347.400 204.600 359.400 ;
        RECT 205.800 348.300 207.600 359.400 ;
        RECT 211.800 348.300 213.600 359.400 ;
        RECT 205.800 347.400 213.600 348.300 ;
        RECT 219.600 347.400 221.400 359.400 ;
        RECT 229.800 358.500 237.600 359.400 ;
        RECT 229.800 347.400 231.600 358.500 ;
        RECT 203.400 342.150 204.300 347.400 ;
        RECT 219.000 346.350 221.400 347.400 ;
        RECT 232.800 346.500 234.600 357.600 ;
        RECT 235.800 348.600 237.600 358.500 ;
        RECT 241.800 348.600 243.600 359.400 ;
        RECT 247.800 353.400 249.600 359.400 ;
        RECT 235.800 347.700 243.600 348.600 ;
        RECT 215.100 342.150 216.900 343.950 ;
        RECT 155.850 335.700 159.600 336.750 ;
        RECT 139.200 331.950 144.600 333.600 ;
        RECT 149.400 332.700 157.200 334.050 ;
        RECT 128.400 327.600 130.200 330.600 ;
        RECT 139.200 327.600 141.000 331.950 ;
        RECT 149.400 327.600 151.200 332.700 ;
        RECT 155.400 327.600 157.200 332.700 ;
        RECT 158.400 333.600 159.600 335.700 ;
        RECT 158.400 327.600 160.200 333.600 ;
        RECT 170.400 330.600 171.600 338.850 ;
        RECT 172.950 337.050 175.050 339.150 ;
        RECT 184.950 337.050 187.050 339.150 ;
        RECT 193.950 338.850 196.050 340.950 ;
        RECT 197.100 339.150 198.900 340.950 ;
        RECT 202.950 340.050 205.050 342.150 ;
        RECT 184.950 330.600 186.000 337.050 ;
        RECT 194.400 330.600 195.600 338.850 ;
        RECT 196.950 337.050 199.050 339.150 ;
        RECT 203.400 333.600 204.300 340.050 ;
        RECT 205.950 338.850 208.050 340.950 ;
        RECT 209.100 339.150 210.900 340.950 ;
        RECT 206.100 337.050 207.900 338.850 ;
        RECT 208.950 337.050 211.050 339.150 ;
        RECT 211.950 338.850 214.050 340.950 ;
        RECT 214.950 340.050 217.050 342.150 ;
        RECT 219.000 339.150 220.050 346.350 ;
        RECT 232.800 345.600 236.850 346.500 ;
        RECT 221.100 342.150 222.900 343.950 ;
        RECT 230.100 342.150 231.900 343.950 ;
        RECT 235.950 342.150 236.850 345.600 ;
        RECT 241.950 342.150 243.750 343.950 ;
        RECT 220.950 340.050 223.050 342.150 ;
        RECT 229.950 340.050 232.050 342.150 ;
        RECT 212.100 337.050 213.900 338.850 ;
        RECT 217.950 337.050 220.050 339.150 ;
        RECT 232.950 338.850 235.050 340.950 ;
        RECT 235.950 340.050 238.050 342.150 ;
        RECT 233.250 337.050 235.050 338.850 ;
        RECT 203.400 331.950 208.800 333.600 ;
        RECT 169.800 327.600 171.600 330.600 ;
        RECT 184.800 327.600 186.600 330.600 ;
        RECT 193.800 327.600 195.600 330.600 ;
        RECT 207.000 327.600 208.800 331.950 ;
        RECT 219.000 330.600 220.050 337.050 ;
        RECT 237.000 333.600 238.050 340.050 ;
        RECT 238.950 338.850 241.050 340.950 ;
        RECT 241.950 340.050 244.050 342.150 ;
        RECT 248.400 340.950 249.600 353.400 ;
        RECT 255.150 347.400 256.950 359.400 ;
        RECT 263.550 353.400 265.350 359.400 ;
        RECT 263.550 352.500 264.750 353.400 ;
        RECT 271.350 352.500 273.150 359.400 ;
        RECT 279.150 353.400 280.950 359.400 ;
        RECT 259.950 350.400 264.750 352.500 ;
        RECT 267.450 351.450 274.050 352.500 ;
        RECT 267.450 350.700 269.250 351.450 ;
        RECT 272.250 350.700 274.050 351.450 ;
        RECT 279.150 351.300 283.050 353.400 ;
        RECT 263.550 349.500 264.750 350.400 ;
        RECT 276.450 349.800 278.250 350.400 ;
        RECT 263.550 348.300 271.050 349.500 ;
        RECT 269.250 347.700 271.050 348.300 ;
        RECT 271.950 348.900 278.250 349.800 ;
        RECT 255.150 346.800 266.250 347.400 ;
        RECT 271.950 346.800 272.850 348.900 ;
        RECT 276.450 348.600 278.250 348.900 ;
        RECT 279.150 348.600 281.850 350.400 ;
        RECT 279.150 347.700 280.050 348.600 ;
        RECT 255.150 346.200 272.850 346.800 ;
        RECT 247.950 338.850 250.050 340.950 ;
        RECT 251.100 339.150 252.900 340.950 ;
        RECT 238.950 337.050 240.750 338.850 ;
        RECT 218.400 327.600 220.200 330.600 ;
        RECT 237.000 327.600 238.800 333.600 ;
        RECT 248.400 330.600 249.600 338.850 ;
        RECT 250.950 337.050 253.050 339.150 ;
        RECT 247.800 327.600 249.600 330.600 ;
        RECT 255.150 333.600 256.050 346.200 ;
        RECT 264.450 345.900 272.850 346.200 ;
        RECT 274.050 346.800 280.050 347.700 ;
        RECT 280.950 346.800 283.050 347.700 ;
        RECT 286.650 347.400 288.450 359.400 ;
        RECT 264.450 345.600 266.250 345.900 ;
        RECT 274.050 342.150 274.950 346.800 ;
        RECT 280.950 345.600 285.150 346.800 ;
        RECT 284.250 343.800 286.050 345.600 ;
        RECT 265.950 341.100 268.050 342.150 ;
        RECT 257.100 339.150 258.900 340.950 ;
        RECT 260.100 340.050 268.050 341.100 ;
        RECT 271.950 340.050 274.950 342.150 ;
        RECT 260.100 339.300 261.900 340.050 ;
        RECT 258.000 338.400 258.900 339.150 ;
        RECT 263.100 338.400 264.900 339.000 ;
        RECT 258.000 337.200 264.900 338.400 ;
        RECT 263.850 336.000 264.900 337.200 ;
        RECT 274.050 336.000 274.950 340.050 ;
        RECT 283.950 339.750 286.050 340.050 ;
        RECT 282.150 337.950 286.050 339.750 ;
        RECT 287.250 337.950 288.450 347.400 ;
        RECT 290.400 353.400 292.200 359.400 ;
        RECT 290.400 346.500 291.600 353.400 ;
        RECT 296.700 347.400 298.500 359.400 ;
        RECT 311.700 347.400 313.500 359.400 ;
        RECT 322.800 358.500 330.600 359.400 ;
        RECT 322.800 347.400 324.600 358.500 ;
        RECT 290.400 345.600 296.100 346.500 ;
        RECT 294.150 344.700 296.100 345.600 ;
        RECT 290.100 342.150 291.900 343.950 ;
        RECT 289.950 340.050 292.050 342.150 ;
        RECT 263.850 335.100 274.950 336.000 ;
        RECT 283.950 335.850 288.450 337.950 ;
        RECT 263.850 334.200 264.900 335.100 ;
        RECT 274.050 334.800 274.950 335.100 ;
        RECT 255.150 327.600 256.950 333.600 ;
        RECT 259.950 331.500 262.050 333.600 ;
        RECT 263.550 332.400 265.350 334.200 ;
        RECT 266.850 333.450 268.650 334.200 ;
        RECT 266.850 332.400 271.800 333.450 ;
        RECT 274.050 333.000 275.850 334.800 ;
        RECT 287.250 333.600 288.450 335.850 ;
        RECT 294.150 336.300 295.050 344.700 ;
        RECT 297.000 342.150 298.200 347.400 ;
        RECT 308.250 345.150 310.050 346.950 ;
        RECT 307.950 343.050 310.050 345.150 ;
        RECT 311.850 342.150 313.050 347.400 ;
        RECT 325.800 346.500 327.600 357.600 ;
        RECT 328.800 348.600 330.600 358.500 ;
        RECT 334.800 348.600 336.600 359.400 ;
        RECT 340.800 353.400 342.600 359.400 ;
        RECT 328.800 347.700 336.600 348.600 ;
        RECT 325.800 345.600 329.850 346.500 ;
        RECT 317.100 342.150 318.900 343.950 ;
        RECT 323.100 342.150 324.900 343.950 ;
        RECT 328.950 342.150 329.850 345.600 ;
        RECT 334.950 342.150 336.750 343.950 ;
        RECT 295.950 340.050 298.200 342.150 ;
        RECT 294.150 335.400 296.100 336.300 ;
        RECT 280.950 332.700 283.050 333.600 ;
        RECT 261.000 330.600 262.050 331.500 ;
        RECT 270.750 330.600 271.800 332.400 ;
        RECT 279.300 331.500 283.050 332.700 ;
        RECT 279.300 330.600 280.350 331.500 ;
        RECT 261.000 329.700 264.750 330.600 ;
        RECT 262.950 327.600 264.750 329.700 ;
        RECT 270.750 327.600 272.550 330.600 ;
        RECT 278.550 327.600 280.350 330.600 ;
        RECT 286.650 327.600 288.450 333.600 ;
        RECT 291.000 334.500 296.100 335.400 ;
        RECT 291.000 330.600 292.200 334.500 ;
        RECT 297.000 333.600 298.200 340.050 ;
        RECT 310.950 340.050 313.050 342.150 ;
        RECT 310.950 336.750 312.150 340.050 ;
        RECT 313.950 338.850 316.050 340.950 ;
        RECT 316.950 340.050 319.050 342.150 ;
        RECT 322.950 340.050 325.050 342.150 ;
        RECT 325.950 338.850 328.050 340.950 ;
        RECT 328.950 340.050 331.050 342.150 ;
        RECT 314.100 337.050 315.900 338.850 ;
        RECT 326.250 337.050 328.050 338.850 ;
        RECT 308.400 335.700 312.150 336.750 ;
        RECT 308.400 333.600 309.600 335.700 ;
        RECT 290.400 327.600 292.200 330.600 ;
        RECT 296.700 327.600 298.500 333.600 ;
        RECT 307.800 327.600 309.600 333.600 ;
        RECT 310.800 332.700 318.600 334.050 ;
        RECT 310.800 327.600 312.600 332.700 ;
        RECT 316.800 327.600 318.600 332.700 ;
        RECT 330.000 333.600 331.050 340.050 ;
        RECT 331.950 338.850 334.050 340.950 ;
        RECT 334.950 340.050 337.050 342.150 ;
        RECT 341.400 340.950 342.600 353.400 ;
        RECT 348.150 347.400 349.950 359.400 ;
        RECT 356.550 353.400 358.350 359.400 ;
        RECT 356.550 352.500 357.750 353.400 ;
        RECT 364.350 352.500 366.150 359.400 ;
        RECT 372.150 353.400 373.950 359.400 ;
        RECT 352.950 350.400 357.750 352.500 ;
        RECT 360.450 351.450 367.050 352.500 ;
        RECT 360.450 350.700 362.250 351.450 ;
        RECT 365.250 350.700 367.050 351.450 ;
        RECT 372.150 351.300 376.050 353.400 ;
        RECT 356.550 349.500 357.750 350.400 ;
        RECT 369.450 349.800 371.250 350.400 ;
        RECT 356.550 348.300 364.050 349.500 ;
        RECT 362.250 347.700 364.050 348.300 ;
        RECT 364.950 348.900 371.250 349.800 ;
        RECT 348.150 346.800 359.250 347.400 ;
        RECT 364.950 346.800 365.850 348.900 ;
        RECT 369.450 348.600 371.250 348.900 ;
        RECT 372.150 348.600 374.850 350.400 ;
        RECT 372.150 347.700 373.050 348.600 ;
        RECT 348.150 346.200 365.850 346.800 ;
        RECT 340.950 338.850 343.050 340.950 ;
        RECT 344.100 339.150 345.900 340.950 ;
        RECT 331.950 337.050 333.750 338.850 ;
        RECT 330.000 327.600 331.800 333.600 ;
        RECT 341.400 330.600 342.600 338.850 ;
        RECT 343.950 337.050 346.050 339.150 ;
        RECT 340.800 327.600 342.600 330.600 ;
        RECT 348.150 333.600 349.050 346.200 ;
        RECT 357.450 345.900 365.850 346.200 ;
        RECT 367.050 346.800 373.050 347.700 ;
        RECT 373.950 346.800 376.050 347.700 ;
        RECT 379.650 347.400 381.450 359.400 ;
        RECT 389.400 353.400 391.200 359.400 ;
        RECT 357.450 345.600 359.250 345.900 ;
        RECT 367.050 342.150 367.950 346.800 ;
        RECT 373.950 345.600 378.150 346.800 ;
        RECT 377.250 343.800 379.050 345.600 ;
        RECT 358.950 341.100 361.050 342.150 ;
        RECT 350.100 339.150 351.900 340.950 ;
        RECT 353.100 340.050 361.050 341.100 ;
        RECT 364.950 340.050 367.950 342.150 ;
        RECT 353.100 339.300 354.900 340.050 ;
        RECT 351.000 338.400 351.900 339.150 ;
        RECT 356.100 338.400 357.900 339.000 ;
        RECT 351.000 337.200 357.900 338.400 ;
        RECT 356.850 336.000 357.900 337.200 ;
        RECT 367.050 336.000 367.950 340.050 ;
        RECT 376.950 339.750 379.050 340.050 ;
        RECT 375.150 337.950 379.050 339.750 ;
        RECT 380.250 337.950 381.450 347.400 ;
        RECT 386.100 342.150 387.900 343.950 ;
        RECT 385.950 340.050 388.050 342.150 ;
        RECT 356.850 335.100 367.950 336.000 ;
        RECT 376.950 335.850 381.450 337.950 ;
        RECT 389.550 336.300 390.600 353.400 ;
        RECT 396.000 347.400 397.800 359.400 ;
        RECT 409.800 353.400 411.600 359.400 ;
        RECT 421.800 353.400 423.600 359.400 ;
        RECT 391.950 341.850 394.050 343.950 ;
        RECT 396.000 342.150 397.050 347.400 ;
        RECT 410.400 345.150 411.600 353.400 ;
        RECT 392.100 340.050 393.900 341.850 ;
        RECT 394.950 340.050 397.050 342.150 ;
        RECT 406.950 341.850 409.050 343.950 ;
        RECT 409.950 343.050 412.050 345.150 ;
        RECT 407.100 340.050 408.900 341.850 ;
        RECT 356.850 334.200 357.900 335.100 ;
        RECT 367.050 334.800 367.950 335.100 ;
        RECT 348.150 327.600 349.950 333.600 ;
        RECT 352.950 331.500 355.050 333.600 ;
        RECT 356.550 332.400 358.350 334.200 ;
        RECT 359.850 333.450 361.650 334.200 ;
        RECT 359.850 332.400 364.800 333.450 ;
        RECT 367.050 333.000 368.850 334.800 ;
        RECT 380.250 333.600 381.450 335.850 ;
        RECT 373.950 332.700 376.050 333.600 ;
        RECT 354.000 330.600 355.050 331.500 ;
        RECT 363.750 330.600 364.800 332.400 ;
        RECT 372.300 331.500 376.050 332.700 ;
        RECT 372.300 330.600 373.350 331.500 ;
        RECT 354.000 329.700 357.750 330.600 ;
        RECT 355.950 327.600 357.750 329.700 ;
        RECT 363.750 327.600 365.550 330.600 ;
        RECT 371.550 327.600 373.350 330.600 ;
        RECT 379.650 327.600 381.450 333.600 ;
        RECT 386.400 335.100 393.900 336.300 ;
        RECT 386.400 327.600 388.200 335.100 ;
        RECT 392.100 334.500 393.900 335.100 ;
        RECT 396.000 333.600 397.050 340.050 ;
        RECT 410.400 335.700 411.600 343.050 ;
        RECT 412.950 341.850 415.050 343.950 ;
        RECT 413.100 340.050 414.900 341.850 ;
        RECT 422.400 340.950 423.600 353.400 ;
        RECT 433.500 347.400 435.300 359.400 ;
        RECT 448.800 353.400 450.600 359.400 ;
        RECT 460.800 353.400 462.600 359.400 ;
        RECT 428.100 342.150 429.900 343.950 ;
        RECT 433.950 342.150 435.150 347.400 ;
        RECT 436.950 345.150 438.750 346.950 ;
        RECT 449.400 345.150 450.600 353.400 ;
        RECT 457.950 345.450 460.050 346.050 ;
        RECT 436.950 343.050 439.050 345.150 ;
        RECT 421.950 338.850 424.050 340.950 ;
        RECT 425.100 339.150 426.900 340.950 ;
        RECT 427.950 340.050 430.050 342.150 ;
        RECT 393.900 332.100 397.050 333.600 ;
        RECT 408.000 334.800 411.600 335.700 ;
        RECT 393.900 327.600 395.700 332.100 ;
        RECT 408.000 327.600 409.800 334.800 ;
        RECT 422.400 330.600 423.600 338.850 ;
        RECT 424.950 337.050 427.050 339.150 ;
        RECT 430.950 338.850 433.050 340.950 ;
        RECT 433.950 340.050 436.050 342.150 ;
        RECT 445.950 341.850 448.050 343.950 ;
        RECT 448.950 343.050 451.050 345.150 ;
        RECT 455.550 344.550 460.050 345.450 ;
        RECT 446.100 340.050 447.900 341.850 ;
        RECT 431.100 337.050 432.900 338.850 ;
        RECT 434.850 336.750 436.050 340.050 ;
        RECT 434.850 335.700 438.600 336.750 ;
        RECT 449.400 335.700 450.600 343.050 ;
        RECT 451.950 341.850 454.050 343.950 ;
        RECT 452.100 340.050 453.900 341.850 ;
        RECT 421.800 327.600 423.600 330.600 ;
        RECT 428.400 332.700 436.200 334.050 ;
        RECT 428.400 327.600 430.200 332.700 ;
        RECT 434.400 327.600 436.200 332.700 ;
        RECT 437.400 333.600 438.600 335.700 ;
        RECT 447.000 334.800 450.600 335.700 ;
        RECT 451.950 336.450 454.050 337.050 ;
        RECT 455.550 336.450 456.450 344.550 ;
        RECT 457.950 343.950 460.050 344.550 ;
        RECT 461.400 340.950 462.600 353.400 ;
        RECT 470.400 353.400 472.200 359.400 ;
        RECT 470.400 345.150 471.600 353.400 ;
        RECT 472.950 348.450 475.050 349.050 ;
        RECT 472.950 347.550 477.450 348.450 ;
        RECT 472.950 346.950 475.050 347.550 ;
        RECT 466.950 341.850 469.050 343.950 ;
        RECT 469.950 343.050 472.050 345.150 ;
        RECT 460.950 338.850 463.050 340.950 ;
        RECT 464.100 339.150 465.900 340.950 ;
        RECT 467.100 340.050 468.900 341.850 ;
        RECT 451.950 335.550 456.450 336.450 ;
        RECT 451.950 334.950 454.050 335.550 ;
        RECT 437.400 327.600 439.200 333.600 ;
        RECT 447.000 327.600 448.800 334.800 ;
        RECT 461.400 330.600 462.600 338.850 ;
        RECT 463.950 337.050 466.050 339.150 ;
        RECT 470.400 335.700 471.600 343.050 ;
        RECT 472.950 341.850 475.050 343.950 ;
        RECT 473.100 340.050 474.900 341.850 ;
        RECT 476.550 340.050 477.450 347.550 ;
        RECT 483.600 347.400 485.400 359.400 ;
        RECT 496.800 353.400 498.600 359.400 ;
        RECT 483.000 346.350 485.400 347.400 ;
        RECT 497.700 353.100 498.600 353.400 ;
        RECT 502.800 353.400 504.600 359.400 ;
        RECT 502.800 353.100 504.300 353.400 ;
        RECT 497.700 352.200 504.300 353.100 ;
        RECT 479.100 342.150 480.900 343.950 ;
        RECT 478.950 340.050 481.050 342.150 ;
        RECT 475.950 337.950 478.050 340.050 ;
        RECT 483.000 339.150 484.050 346.350 ;
        RECT 497.700 343.950 498.600 352.200 ;
        RECT 503.100 348.150 504.900 349.950 ;
        RECT 499.950 345.150 501.750 346.950 ;
        RECT 502.950 346.050 505.050 348.150 ;
        RECT 515.700 347.400 517.500 359.400 ;
        RECT 529.500 347.400 531.300 359.400 ;
        RECT 539.400 348.300 541.200 359.400 ;
        RECT 545.400 348.300 547.200 359.400 ;
        RECT 539.400 347.400 547.200 348.300 ;
        RECT 548.400 347.400 550.200 359.400 ;
        RECT 553.950 349.950 556.050 352.050 ;
        RECT 506.100 345.150 507.900 346.950 ;
        RECT 512.250 345.150 514.050 346.950 ;
        RECT 485.100 342.150 486.900 343.950 ;
        RECT 484.950 340.050 487.050 342.150 ;
        RECT 496.950 341.850 499.050 343.950 ;
        RECT 499.950 343.050 502.050 345.150 ;
        RECT 505.950 343.050 508.050 345.150 ;
        RECT 511.950 343.050 514.050 345.150 ;
        RECT 515.850 342.150 517.050 347.400 ;
        RECT 521.100 342.150 522.900 343.950 ;
        RECT 524.100 342.150 525.900 343.950 ;
        RECT 529.950 342.150 531.150 347.400 ;
        RECT 532.950 345.150 534.750 346.950 ;
        RECT 532.950 343.050 535.050 345.150 ;
        RECT 548.700 342.150 549.600 347.400 ;
        RECT 481.950 337.050 484.050 339.150 ;
        RECT 470.400 334.800 474.000 335.700 ;
        RECT 460.800 327.600 462.600 330.600 ;
        RECT 472.200 327.600 474.000 334.800 ;
        RECT 483.000 330.600 484.050 337.050 ;
        RECT 497.700 337.650 498.600 341.850 ;
        RECT 514.950 340.050 517.050 342.150 ;
        RECT 497.700 336.000 501.900 337.650 ;
        RECT 514.950 336.750 516.150 340.050 ;
        RECT 517.950 338.850 520.050 340.950 ;
        RECT 520.950 340.050 523.050 342.150 ;
        RECT 523.950 340.050 526.050 342.150 ;
        RECT 526.950 338.850 529.050 340.950 ;
        RECT 529.950 340.050 532.050 342.150 ;
        RECT 518.100 337.050 519.900 338.850 ;
        RECT 527.100 337.050 528.900 338.850 ;
        RECT 482.400 327.600 484.200 330.600 ;
        RECT 500.100 327.600 501.900 336.000 ;
        RECT 512.400 335.700 516.150 336.750 ;
        RECT 530.850 336.750 532.050 340.050 ;
        RECT 538.950 338.850 541.050 340.950 ;
        RECT 542.100 339.150 543.900 340.950 ;
        RECT 539.100 337.050 540.900 338.850 ;
        RECT 541.950 337.050 544.050 339.150 ;
        RECT 544.950 338.850 547.050 340.950 ;
        RECT 547.950 340.050 550.050 342.150 ;
        RECT 554.550 340.050 555.450 349.950 ;
        RECT 560.700 347.400 562.500 359.400 ;
        RECT 571.200 358.500 579.000 359.400 ;
        RECT 571.200 349.200 573.000 358.500 ;
        RECT 574.200 349.800 576.000 357.600 ;
        RECT 574.800 347.400 576.000 349.800 ;
        RECT 577.200 349.800 579.000 358.500 ;
        RECT 580.800 358.500 588.600 359.400 ;
        RECT 580.800 350.700 582.600 358.500 ;
        RECT 583.800 349.800 585.600 357.600 ;
        RECT 577.200 348.900 585.600 349.800 ;
        RECT 586.800 349.500 588.600 358.500 ;
        RECT 592.800 349.500 594.600 359.400 ;
        RECT 586.800 348.600 594.600 349.500 ;
        RECT 599.400 353.400 601.200 359.400 ;
        RECT 557.250 345.150 559.050 346.950 ;
        RECT 556.950 343.050 559.050 345.150 ;
        RECT 560.850 342.150 562.050 347.400 ;
        RECT 574.800 346.200 578.250 347.400 ;
        RECT 566.100 342.150 567.900 343.950 ;
        RECT 559.950 340.050 562.050 342.150 ;
        RECT 545.100 337.050 546.900 338.850 ;
        RECT 530.850 335.700 534.600 336.750 ;
        RECT 512.400 333.600 513.600 335.700 ;
        RECT 511.800 327.600 513.600 333.600 ;
        RECT 514.800 332.700 522.600 334.050 ;
        RECT 514.800 327.600 516.600 332.700 ;
        RECT 520.800 327.600 522.600 332.700 ;
        RECT 524.400 332.700 532.200 334.050 ;
        RECT 524.400 327.600 526.200 332.700 ;
        RECT 530.400 327.600 532.200 332.700 ;
        RECT 533.400 333.600 534.600 335.700 ;
        RECT 548.700 333.600 549.600 340.050 ;
        RECT 553.950 337.950 556.050 340.050 ;
        RECT 559.950 336.750 561.150 340.050 ;
        RECT 562.950 338.850 565.050 340.950 ;
        RECT 565.950 340.050 568.050 342.150 ;
        RECT 577.050 340.800 578.250 346.200 ;
        RECT 583.950 345.450 586.050 346.050 ;
        RECT 583.950 344.550 588.450 345.450 ;
        RECT 583.950 343.950 586.050 344.550 ;
        RECT 581.100 342.000 582.900 343.800 ;
        RECT 563.100 337.050 564.900 338.850 ;
        RECT 574.950 338.700 578.250 340.800 ;
        RECT 580.950 339.900 583.050 342.000 ;
        RECT 583.950 338.700 586.050 340.800 ;
        RECT 557.400 335.700 561.150 336.750 ;
        RECT 557.400 333.600 558.600 335.700 ;
        RECT 533.400 327.600 535.200 333.600 ;
        RECT 544.200 331.950 549.600 333.600 ;
        RECT 544.200 327.600 546.000 331.950 ;
        RECT 556.800 327.600 558.600 333.600 ;
        RECT 559.800 332.700 567.600 334.050 ;
        RECT 559.800 327.600 561.600 332.700 ;
        RECT 565.800 327.600 567.600 332.700 ;
        RECT 577.050 332.400 578.250 338.700 ;
        RECT 584.100 336.900 585.900 338.700 ;
        RECT 587.550 336.450 588.450 344.550 ;
        RECT 590.100 342.000 591.900 343.800 ;
        RECT 589.950 339.900 592.050 342.000 ;
        RECT 599.400 340.950 600.600 353.400 ;
        RECT 607.800 347.400 609.600 359.400 ;
        RECT 610.800 348.300 612.600 359.400 ;
        RECT 616.800 348.300 618.600 359.400 ;
        RECT 626.400 353.400 628.200 359.400 ;
        RECT 626.700 353.100 628.200 353.400 ;
        RECT 632.400 353.400 634.200 359.400 ;
        RECT 632.400 353.100 633.300 353.400 ;
        RECT 626.700 352.200 633.300 353.100 ;
        RECT 610.800 347.400 618.600 348.300 ;
        RECT 626.100 348.150 627.900 349.950 ;
        RECT 608.400 342.150 609.300 347.400 ;
        RECT 623.100 345.150 624.900 346.950 ;
        RECT 625.950 346.050 628.050 348.150 ;
        RECT 629.250 345.150 631.050 346.950 ;
        RECT 622.950 343.050 625.050 345.150 ;
        RECT 628.950 343.050 631.050 345.150 ;
        RECT 632.400 343.950 633.300 352.200 ;
        RECT 643.500 347.400 645.300 359.400 ;
        RECT 655.800 347.400 657.600 359.400 ;
        RECT 658.800 348.300 660.600 359.400 ;
        RECT 664.800 348.300 666.600 359.400 ;
        RECT 670.800 353.400 672.600 359.400 ;
        RECT 658.800 347.400 666.600 348.300 ;
        RECT 671.700 353.100 672.600 353.400 ;
        RECT 676.800 353.400 678.600 359.400 ;
        RECT 688.800 353.400 690.600 359.400 ;
        RECT 676.800 353.100 678.300 353.400 ;
        RECT 671.700 352.200 678.300 353.100 ;
        RECT 689.700 353.100 690.600 353.400 ;
        RECT 694.800 353.400 696.600 359.400 ;
        RECT 706.800 353.400 708.600 359.400 ;
        RECT 694.800 353.100 696.300 353.400 ;
        RECT 689.700 352.200 696.300 353.100 ;
        RECT 707.700 353.100 708.600 353.400 ;
        RECT 712.800 353.400 714.600 359.400 ;
        RECT 712.800 353.100 714.300 353.400 ;
        RECT 707.700 352.200 714.300 353.100 ;
        RECT 596.100 339.150 597.900 340.950 ;
        RECT 595.950 337.050 598.050 339.150 ;
        RECT 598.950 338.850 601.050 340.950 ;
        RECT 607.950 340.050 610.050 342.150 ;
        RECT 631.950 341.850 634.050 343.950 ;
        RECT 638.100 342.150 639.900 343.950 ;
        RECT 643.950 342.150 645.150 347.400 ;
        RECT 646.950 345.150 648.750 346.950 ;
        RECT 646.950 343.050 649.050 345.150 ;
        RECT 656.400 342.150 657.300 347.400 ;
        RECT 661.950 345.450 664.050 346.050 ;
        RECT 661.950 344.550 669.450 345.450 ;
        RECT 661.950 343.950 664.050 344.550 ;
        RECT 587.550 335.550 594.450 336.450 ;
        RECT 593.550 333.450 594.450 335.550 ;
        RECT 595.950 333.450 598.050 334.050 ;
        RECT 593.550 332.550 598.050 333.450 ;
        RECT 577.050 331.500 587.850 332.400 ;
        RECT 595.950 331.950 598.050 332.550 ;
        RECT 580.800 330.600 581.850 331.500 ;
        RECT 586.800 330.600 587.850 331.500 ;
        RECT 599.400 330.600 600.600 338.850 ;
        RECT 608.400 333.600 609.300 340.050 ;
        RECT 610.950 338.850 613.050 340.950 ;
        RECT 614.100 339.150 615.900 340.950 ;
        RECT 611.100 337.050 612.900 338.850 ;
        RECT 613.950 337.050 616.050 339.150 ;
        RECT 616.950 338.850 619.050 340.950 ;
        RECT 617.100 337.050 618.900 338.850 ;
        RECT 632.400 337.650 633.300 341.850 ;
        RECT 637.950 340.050 640.050 342.150 ;
        RECT 640.950 338.850 643.050 340.950 ;
        RECT 643.950 340.050 646.050 342.150 ;
        RECT 655.950 340.050 658.050 342.150 ;
        RECT 629.100 336.000 633.300 337.650 ;
        RECT 641.100 337.050 642.900 338.850 ;
        RECT 644.850 336.750 646.050 340.050 ;
        RECT 608.400 331.950 613.800 333.600 ;
        RECT 580.800 327.600 582.600 330.600 ;
        RECT 586.800 327.600 588.600 330.600 ;
        RECT 599.400 327.600 601.200 330.600 ;
        RECT 612.000 327.600 613.800 331.950 ;
        RECT 629.100 327.600 630.900 336.000 ;
        RECT 644.850 335.700 648.600 336.750 ;
        RECT 638.400 332.700 646.200 334.050 ;
        RECT 638.400 327.600 640.200 332.700 ;
        RECT 644.400 327.600 646.200 332.700 ;
        RECT 647.400 333.600 648.600 335.700 ;
        RECT 656.400 333.600 657.300 340.050 ;
        RECT 658.950 338.850 661.050 340.950 ;
        RECT 662.100 339.150 663.900 340.950 ;
        RECT 659.100 337.050 660.900 338.850 ;
        RECT 661.950 337.050 664.050 339.150 ;
        RECT 664.950 338.850 667.050 340.950 ;
        RECT 665.100 337.050 666.900 338.850 ;
        RECT 668.550 337.050 669.450 344.550 ;
        RECT 671.700 343.950 672.600 352.200 ;
        RECT 677.100 348.150 678.900 349.950 ;
        RECT 673.950 345.150 675.750 346.950 ;
        RECT 676.950 346.050 679.050 348.150 ;
        RECT 680.100 345.150 681.900 346.950 ;
        RECT 670.950 341.850 673.050 343.950 ;
        RECT 673.950 343.050 676.050 345.150 ;
        RECT 679.950 343.050 682.050 345.150 ;
        RECT 689.700 343.950 690.600 352.200 ;
        RECT 695.100 348.150 696.900 349.950 ;
        RECT 691.950 345.150 693.750 346.950 ;
        RECT 694.950 346.050 697.050 348.150 ;
        RECT 698.100 345.150 699.900 346.950 ;
        RECT 688.950 341.850 691.050 343.950 ;
        RECT 691.950 343.050 694.050 345.150 ;
        RECT 697.950 343.050 700.050 345.150 ;
        RECT 707.700 343.950 708.600 352.200 ;
        RECT 713.100 348.150 714.900 349.950 ;
        RECT 709.950 345.150 711.750 346.950 ;
        RECT 712.950 346.050 715.050 348.150 ;
        RECT 728.700 347.400 730.500 359.400 ;
        RECT 742.500 347.400 744.300 359.400 ;
        RECT 755.400 353.400 757.200 359.400 ;
        RECT 755.700 353.100 757.200 353.400 ;
        RECT 761.400 353.400 763.200 359.400 ;
        RECT 761.400 353.100 762.300 353.400 ;
        RECT 755.700 352.200 762.300 353.100 ;
        RECT 755.100 348.150 756.900 349.950 ;
        RECT 716.100 345.150 717.900 346.950 ;
        RECT 725.250 345.150 727.050 346.950 ;
        RECT 706.950 341.850 709.050 343.950 ;
        RECT 709.950 343.050 712.050 345.150 ;
        RECT 715.950 343.050 718.050 345.150 ;
        RECT 724.950 343.050 727.050 345.150 ;
        RECT 728.850 342.150 730.050 347.400 ;
        RECT 734.100 342.150 735.900 343.950 ;
        RECT 737.100 342.150 738.900 343.950 ;
        RECT 742.950 342.150 744.150 347.400 ;
        RECT 745.950 345.150 747.750 346.950 ;
        RECT 752.100 345.150 753.900 346.950 ;
        RECT 754.950 346.050 757.050 348.150 ;
        RECT 758.250 345.150 760.050 346.950 ;
        RECT 745.950 343.050 748.050 345.150 ;
        RECT 751.950 343.050 754.050 345.150 ;
        RECT 757.950 343.050 760.050 345.150 ;
        RECT 761.400 343.950 762.300 352.200 ;
        RECT 671.700 337.650 672.600 341.850 ;
        RECT 689.700 337.650 690.600 341.850 ;
        RECT 707.700 337.650 708.600 341.850 ;
        RECT 727.950 340.050 730.050 342.150 ;
        RECT 667.950 334.950 670.050 337.050 ;
        RECT 671.700 336.000 675.900 337.650 ;
        RECT 689.700 336.000 693.900 337.650 ;
        RECT 707.700 336.000 711.900 337.650 ;
        RECT 727.950 336.750 729.150 340.050 ;
        RECT 730.950 338.850 733.050 340.950 ;
        RECT 733.950 340.050 736.050 342.150 ;
        RECT 736.950 340.050 739.050 342.150 ;
        RECT 739.950 338.850 742.050 340.950 ;
        RECT 742.950 340.050 745.050 342.150 ;
        RECT 760.950 341.850 763.050 343.950 ;
        RECT 731.100 337.050 732.900 338.850 ;
        RECT 740.100 337.050 741.900 338.850 ;
        RECT 647.400 327.600 649.200 333.600 ;
        RECT 656.400 331.950 661.800 333.600 ;
        RECT 660.000 327.600 661.800 331.950 ;
        RECT 674.100 327.600 675.900 336.000 ;
        RECT 692.100 327.600 693.900 336.000 ;
        RECT 700.950 333.450 703.050 334.050 ;
        RECT 706.950 333.450 709.050 334.050 ;
        RECT 700.950 332.550 709.050 333.450 ;
        RECT 700.950 331.950 703.050 332.550 ;
        RECT 706.950 331.950 709.050 332.550 ;
        RECT 710.100 327.600 711.900 336.000 ;
        RECT 725.400 335.700 729.150 336.750 ;
        RECT 743.850 336.750 745.050 340.050 ;
        RECT 761.400 337.650 762.300 341.850 ;
        RECT 743.850 335.700 747.600 336.750 ;
        RECT 725.400 333.600 726.600 335.700 ;
        RECT 724.800 327.600 726.600 333.600 ;
        RECT 727.800 332.700 735.600 334.050 ;
        RECT 727.800 327.600 729.600 332.700 ;
        RECT 733.800 327.600 735.600 332.700 ;
        RECT 737.400 332.700 745.200 334.050 ;
        RECT 737.400 327.600 739.200 332.700 ;
        RECT 743.400 327.600 745.200 332.700 ;
        RECT 746.400 333.600 747.600 335.700 ;
        RECT 758.100 336.000 762.300 337.650 ;
        RECT 746.400 327.600 748.200 333.600 ;
        RECT 758.100 327.600 759.900 336.000 ;
        RECT 7.800 320.400 9.600 323.400 ;
        RECT 8.400 312.150 9.600 320.400 ;
        RECT 18.000 316.200 19.800 323.400 ;
        RECT 31.200 316.200 33.000 323.400 ;
        RECT 18.000 315.300 21.600 316.200 ;
        RECT 7.950 310.050 10.050 312.150 ;
        RECT 10.950 311.850 13.050 313.950 ;
        RECT 11.100 310.050 12.900 311.850 ;
        RECT 8.400 297.600 9.600 310.050 ;
        RECT 17.100 309.150 18.900 310.950 ;
        RECT 16.950 307.050 19.050 309.150 ;
        RECT 20.400 307.950 21.600 315.300 ;
        RECT 29.400 315.300 33.000 316.200 ;
        RECT 23.100 309.150 24.900 310.950 ;
        RECT 26.100 309.150 27.900 310.950 ;
        RECT 19.950 305.850 22.050 307.950 ;
        RECT 22.950 307.050 25.050 309.150 ;
        RECT 25.950 307.050 28.050 309.150 ;
        RECT 29.400 307.950 30.600 315.300 ;
        RECT 47.100 315.000 48.900 323.400 ;
        RECT 61.200 316.200 63.000 323.400 ;
        RECT 70.800 317.400 72.600 323.400 ;
        RECT 59.400 315.300 63.000 316.200 ;
        RECT 71.400 315.300 72.600 317.400 ;
        RECT 73.800 318.300 75.600 323.400 ;
        RECT 79.800 318.300 81.600 323.400 ;
        RECT 73.800 316.950 81.600 318.300 ;
        RECT 88.200 316.200 90.000 323.400 ;
        RECT 98.400 320.400 100.200 323.400 ;
        RECT 86.400 315.300 90.000 316.200 ;
        RECT 99.300 316.200 100.200 320.400 ;
        RECT 104.400 317.400 106.200 323.400 ;
        RECT 99.300 315.300 102.750 316.200 ;
        RECT 47.100 313.350 51.300 315.000 ;
        RECT 32.100 309.150 33.900 310.950 ;
        RECT 50.400 309.150 51.300 313.350 ;
        RECT 56.100 309.150 57.900 310.950 ;
        RECT 28.950 305.850 31.050 307.950 ;
        RECT 31.950 307.050 34.050 309.150 ;
        RECT 40.950 305.850 43.050 307.950 ;
        RECT 46.950 305.850 49.050 307.950 ;
        RECT 49.950 307.050 52.050 309.150 ;
        RECT 55.950 307.050 58.050 309.150 ;
        RECT 59.400 307.950 60.600 315.300 ;
        RECT 71.400 314.250 75.150 315.300 ;
        RECT 73.950 310.950 75.150 314.250 ;
        RECT 77.100 312.150 78.900 313.950 ;
        RECT 62.100 309.150 63.900 310.950 ;
        RECT 20.400 297.600 21.600 305.850 ;
        RECT 7.800 291.600 9.600 297.600 ;
        RECT 19.800 291.600 21.600 297.600 ;
        RECT 29.400 297.600 30.600 305.850 ;
        RECT 41.100 304.050 42.900 305.850 ;
        RECT 43.950 302.850 46.050 304.950 ;
        RECT 47.250 304.050 49.050 305.850 ;
        RECT 44.100 301.050 45.900 302.850 ;
        RECT 50.400 298.800 51.300 307.050 ;
        RECT 58.950 305.850 61.050 307.950 ;
        RECT 61.950 307.050 64.050 309.150 ;
        RECT 73.950 308.850 76.050 310.950 ;
        RECT 76.950 310.050 79.050 312.150 ;
        RECT 79.950 308.850 82.050 310.950 ;
        RECT 83.100 309.150 84.900 310.950 ;
        RECT 70.950 305.850 73.050 307.950 ;
        RECT 44.700 297.900 51.300 298.800 ;
        RECT 44.700 297.600 46.200 297.900 ;
        RECT 29.400 291.600 31.200 297.600 ;
        RECT 44.400 291.600 46.200 297.600 ;
        RECT 50.400 297.600 51.300 297.900 ;
        RECT 59.400 297.600 60.600 305.850 ;
        RECT 71.250 304.050 73.050 305.850 ;
        RECT 74.850 303.600 76.050 308.850 ;
        RECT 80.100 307.050 81.900 308.850 ;
        RECT 82.950 307.050 85.050 309.150 ;
        RECT 86.400 307.950 87.600 315.300 ;
        RECT 100.950 314.400 102.750 315.300 ;
        RECT 94.950 311.850 97.050 313.950 ;
        RECT 89.100 309.150 90.900 310.950 ;
        RECT 95.100 310.050 96.900 311.850 ;
        RECT 85.950 305.850 88.050 307.950 ;
        RECT 88.950 307.050 91.050 309.150 ;
        RECT 97.950 308.850 100.050 310.950 ;
        RECT 98.100 307.050 99.900 308.850 ;
        RECT 101.700 306.150 102.600 314.400 ;
        RECT 105.000 312.150 106.050 317.400 ;
        RECT 117.000 316.200 118.800 323.400 ;
        RECT 117.000 315.300 120.600 316.200 ;
        RECT 100.800 306.000 102.600 306.150 ;
        RECT 50.400 291.600 52.200 297.600 ;
        RECT 59.400 291.600 61.200 297.600 ;
        RECT 74.700 291.600 76.500 303.600 ;
        RECT 86.400 297.600 87.600 305.850 ;
        RECT 95.400 304.800 102.600 306.000 ;
        RECT 95.400 303.600 96.600 304.800 ;
        RECT 100.800 304.350 102.600 304.800 ;
        RECT 103.950 310.050 106.050 312.150 ;
        RECT 86.400 291.600 88.200 297.600 ;
        RECT 95.400 291.600 97.200 303.600 ;
        RECT 103.950 303.450 105.300 310.050 ;
        RECT 116.100 309.150 117.900 310.950 ;
        RECT 115.950 307.050 118.050 309.150 ;
        RECT 119.400 307.950 120.600 315.300 ;
        RECT 131.100 315.000 132.900 323.400 ;
        RECT 143.400 320.400 145.200 323.400 ;
        RECT 128.700 313.350 132.900 315.000 ;
        RECT 144.000 313.950 145.050 320.400 ;
        RECT 162.000 319.050 163.800 323.400 ;
        RECT 180.000 319.050 181.800 323.400 ;
        RECT 122.100 309.150 123.900 310.950 ;
        RECT 128.700 309.150 129.600 313.350 ;
        RECT 142.950 311.850 145.050 313.950 ;
        RECT 118.950 305.850 121.050 307.950 ;
        RECT 121.950 307.050 124.050 309.150 ;
        RECT 127.950 307.050 130.050 309.150 ;
        RECT 139.950 308.850 142.050 310.950 ;
        RECT 102.900 302.100 105.300 303.450 ;
        RECT 102.900 291.600 104.700 302.100 ;
        RECT 119.400 297.600 120.600 305.850 ;
        RECT 128.700 298.800 129.600 307.050 ;
        RECT 130.950 305.850 133.050 307.950 ;
        RECT 136.950 305.850 139.050 307.950 ;
        RECT 140.100 307.050 141.900 308.850 ;
        RECT 130.950 304.050 132.750 305.850 ;
        RECT 133.950 302.850 136.050 304.950 ;
        RECT 137.100 304.050 138.900 305.850 ;
        RECT 144.000 304.650 145.050 311.850 ;
        RECT 158.400 317.400 163.800 319.050 ;
        RECT 176.400 317.400 181.800 319.050 ;
        RECT 188.400 318.300 190.200 323.400 ;
        RECT 194.400 318.300 196.200 323.400 ;
        RECT 158.400 310.950 159.300 317.400 ;
        RECT 161.100 312.150 162.900 313.950 ;
        RECT 145.950 308.850 148.050 310.950 ;
        RECT 157.950 308.850 160.050 310.950 ;
        RECT 160.950 310.050 163.050 312.150 ;
        RECT 163.950 311.850 166.050 313.950 ;
        RECT 167.100 312.150 168.900 313.950 ;
        RECT 164.100 310.050 165.900 311.850 ;
        RECT 166.950 310.050 169.050 312.150 ;
        RECT 176.400 310.950 177.300 317.400 ;
        RECT 188.400 316.950 196.200 318.300 ;
        RECT 197.400 317.400 199.200 323.400 ;
        RECT 197.400 315.300 198.600 317.400 ;
        RECT 208.200 316.200 210.000 323.400 ;
        RECT 220.200 317.400 222.000 323.400 ;
        RECT 241.200 319.050 243.000 323.400 ;
        RECT 241.200 317.400 246.600 319.050 ;
        RECT 253.800 317.400 255.600 323.400 ;
        RECT 194.850 314.250 198.600 315.300 ;
        RECT 206.400 315.300 210.000 316.200 ;
        RECT 179.100 312.150 180.900 313.950 ;
        RECT 175.950 308.850 178.050 310.950 ;
        RECT 178.950 310.050 181.050 312.150 ;
        RECT 181.950 311.850 184.050 313.950 ;
        RECT 185.100 312.150 186.900 313.950 ;
        RECT 191.100 312.150 192.900 313.950 ;
        RECT 182.100 310.050 183.900 311.850 ;
        RECT 184.950 310.050 187.050 312.150 ;
        RECT 187.950 308.850 190.050 310.950 ;
        RECT 190.950 310.050 193.050 312.150 ;
        RECT 194.850 310.950 196.050 314.250 ;
        RECT 193.950 308.850 196.050 310.950 ;
        RECT 203.100 309.150 204.900 310.950 ;
        RECT 146.100 307.050 147.900 308.850 ;
        RECT 144.000 303.600 146.400 304.650 ;
        RECT 158.400 303.600 159.300 308.850 ;
        RECT 176.400 303.600 177.300 308.850 ;
        RECT 188.100 307.050 189.900 308.850 ;
        RECT 193.950 303.600 195.150 308.850 ;
        RECT 196.950 305.850 199.050 307.950 ;
        RECT 202.950 307.050 205.050 309.150 ;
        RECT 206.400 307.950 207.600 315.300 ;
        RECT 218.250 312.150 220.050 313.950 ;
        RECT 209.100 309.150 210.900 310.950 ;
        RECT 205.950 305.850 208.050 307.950 ;
        RECT 208.950 307.050 211.050 309.150 ;
        RECT 214.950 308.850 217.050 310.950 ;
        RECT 217.950 310.050 220.050 312.150 ;
        RECT 220.950 310.950 222.000 317.400 ;
        RECT 223.950 312.150 225.750 313.950 ;
        RECT 236.100 312.150 237.900 313.950 ;
        RECT 220.950 308.850 223.050 310.950 ;
        RECT 223.950 310.050 226.050 312.150 ;
        RECT 226.950 308.850 229.050 310.950 ;
        RECT 235.950 310.050 238.050 312.150 ;
        RECT 238.950 311.850 241.050 313.950 ;
        RECT 242.100 312.150 243.900 313.950 ;
        RECT 239.100 310.050 240.900 311.850 ;
        RECT 241.950 310.050 244.050 312.150 ;
        RECT 245.700 310.950 246.600 317.400 ;
        RECT 254.400 315.300 255.600 317.400 ;
        RECT 256.800 318.300 258.600 323.400 ;
        RECT 262.800 318.300 264.600 323.400 ;
        RECT 256.800 316.950 264.600 318.300 ;
        RECT 266.400 318.300 268.200 323.400 ;
        RECT 272.400 318.300 274.200 323.400 ;
        RECT 266.400 316.950 274.200 318.300 ;
        RECT 275.400 317.400 277.200 323.400 ;
        RECT 284.400 320.400 286.200 323.400 ;
        RECT 275.400 315.300 276.600 317.400 ;
        RECT 254.400 314.250 258.150 315.300 ;
        RECT 256.950 310.950 258.150 314.250 ;
        RECT 272.850 314.250 276.600 315.300 ;
        RECT 260.100 312.150 261.900 313.950 ;
        RECT 269.100 312.150 270.900 313.950 ;
        RECT 244.950 308.850 247.050 310.950 ;
        RECT 256.950 308.850 259.050 310.950 ;
        RECT 259.950 310.050 262.050 312.150 ;
        RECT 262.950 308.850 265.050 310.950 ;
        RECT 265.950 308.850 268.050 310.950 ;
        RECT 268.950 310.050 271.050 312.150 ;
        RECT 272.850 310.950 274.050 314.250 ;
        RECT 280.950 311.850 283.050 313.950 ;
        RECT 284.400 312.150 285.600 320.400 ;
        RECT 296.100 315.000 297.900 323.400 ;
        RECT 310.800 320.400 312.600 323.400 ;
        RECT 293.700 313.350 297.900 315.000 ;
        RECT 310.950 313.950 312.000 320.400 ;
        RECT 317.400 318.300 319.200 323.400 ;
        RECT 323.400 318.300 325.200 323.400 ;
        RECT 317.400 316.950 325.200 318.300 ;
        RECT 326.400 317.400 328.200 323.400 ;
        RECT 332.400 320.400 334.200 323.400 ;
        RECT 326.400 315.300 327.600 317.400 ;
        RECT 333.000 316.500 334.200 320.400 ;
        RECT 338.700 317.400 340.500 323.400 ;
        RECT 333.000 315.600 338.100 316.500 ;
        RECT 323.850 314.250 327.600 315.300 ;
        RECT 336.150 314.700 338.100 315.600 ;
        RECT 271.950 308.850 274.050 310.950 ;
        RECT 281.100 310.050 282.900 311.850 ;
        RECT 283.950 310.050 286.050 312.150 ;
        RECT 215.250 307.050 217.050 308.850 ;
        RECT 196.950 304.050 198.750 305.850 ;
        RECT 134.100 301.050 135.900 302.850 ;
        RECT 128.700 297.900 135.300 298.800 ;
        RECT 128.700 297.600 129.600 297.900 ;
        RECT 118.800 291.600 120.600 297.600 ;
        RECT 127.800 291.600 129.600 297.600 ;
        RECT 133.800 297.600 135.300 297.900 ;
        RECT 133.800 291.600 135.600 297.600 ;
        RECT 144.600 291.600 146.400 303.600 ;
        RECT 157.800 291.600 159.600 303.600 ;
        RECT 160.800 302.700 168.600 303.600 ;
        RECT 160.800 291.600 162.600 302.700 ;
        RECT 166.800 291.600 168.600 302.700 ;
        RECT 175.800 291.600 177.600 303.600 ;
        RECT 178.800 302.700 186.600 303.600 ;
        RECT 178.800 291.600 180.600 302.700 ;
        RECT 184.800 291.600 186.600 302.700 ;
        RECT 193.500 291.600 195.300 303.600 ;
        RECT 206.400 297.600 207.600 305.850 ;
        RECT 222.150 305.400 223.050 308.850 ;
        RECT 227.100 307.050 228.900 308.850 ;
        RECT 222.150 304.500 226.200 305.400 ;
        RECT 215.400 302.400 223.200 303.300 ;
        RECT 206.400 291.600 208.200 297.600 ;
        RECT 215.400 291.600 217.200 302.400 ;
        RECT 221.400 292.500 223.200 302.400 ;
        RECT 224.400 293.400 226.200 304.500 ;
        RECT 245.700 303.600 246.600 308.850 ;
        RECT 253.950 305.850 256.050 307.950 ;
        RECT 254.250 304.050 256.050 305.850 ;
        RECT 257.850 303.600 259.050 308.850 ;
        RECT 263.100 307.050 264.900 308.850 ;
        RECT 266.100 307.050 267.900 308.850 ;
        RECT 271.950 303.600 273.150 308.850 ;
        RECT 274.950 305.850 277.050 307.950 ;
        RECT 274.950 304.050 276.750 305.850 ;
        RECT 227.400 292.500 229.200 303.600 ;
        RECT 221.400 291.600 229.200 292.500 ;
        RECT 236.400 302.700 244.200 303.600 ;
        RECT 236.400 291.600 238.200 302.700 ;
        RECT 242.400 291.600 244.200 302.700 ;
        RECT 245.400 291.600 247.200 303.600 ;
        RECT 257.700 291.600 259.500 303.600 ;
        RECT 271.500 291.600 273.300 303.600 ;
        RECT 284.400 297.600 285.600 310.050 ;
        RECT 293.700 309.150 294.600 313.350 ;
        RECT 310.950 311.850 313.050 313.950 ;
        RECT 320.100 312.150 321.900 313.950 ;
        RECT 292.950 307.050 295.050 309.150 ;
        RECT 307.950 308.850 310.050 310.950 ;
        RECT 293.700 298.800 294.600 307.050 ;
        RECT 295.950 305.850 298.050 307.950 ;
        RECT 301.950 305.850 304.050 307.950 ;
        RECT 308.100 307.050 309.900 308.850 ;
        RECT 295.950 304.050 297.750 305.850 ;
        RECT 298.950 302.850 301.050 304.950 ;
        RECT 302.100 304.050 303.900 305.850 ;
        RECT 310.950 304.650 312.000 311.850 ;
        RECT 313.950 308.850 316.050 310.950 ;
        RECT 316.950 308.850 319.050 310.950 ;
        RECT 319.950 310.050 322.050 312.150 ;
        RECT 323.850 310.950 325.050 314.250 ;
        RECT 322.950 308.850 325.050 310.950 ;
        RECT 331.950 308.850 334.050 310.950 ;
        RECT 314.100 307.050 315.900 308.850 ;
        RECT 317.100 307.050 318.900 308.850 ;
        RECT 309.600 303.600 312.000 304.650 ;
        RECT 322.950 303.600 324.150 308.850 ;
        RECT 325.950 305.850 328.050 307.950 ;
        RECT 332.100 307.050 333.900 308.850 ;
        RECT 336.150 306.300 337.050 314.700 ;
        RECT 339.000 310.950 340.200 317.400 ;
        RECT 352.200 316.200 354.000 323.400 ;
        RECT 364.200 316.200 366.000 323.400 ;
        RECT 350.400 315.300 354.000 316.200 ;
        RECT 362.400 315.300 366.000 316.200 ;
        RECT 371.400 315.900 373.200 323.400 ;
        RECT 378.900 318.900 380.700 323.400 ;
        RECT 389.400 320.400 391.200 323.400 ;
        RECT 378.900 317.400 382.050 318.900 ;
        RECT 377.100 315.900 378.900 316.500 ;
        RECT 337.950 308.850 340.200 310.950 ;
        RECT 347.100 309.150 348.900 310.950 ;
        RECT 325.950 304.050 327.750 305.850 ;
        RECT 336.150 305.400 338.100 306.300 ;
        RECT 332.400 304.500 338.100 305.400 ;
        RECT 299.100 301.050 300.900 302.850 ;
        RECT 293.700 297.900 300.300 298.800 ;
        RECT 293.700 297.600 294.600 297.900 ;
        RECT 284.400 291.600 286.200 297.600 ;
        RECT 292.800 291.600 294.600 297.600 ;
        RECT 298.800 297.600 300.300 297.900 ;
        RECT 298.800 291.600 300.600 297.600 ;
        RECT 309.600 291.600 311.400 303.600 ;
        RECT 322.500 291.600 324.300 303.600 ;
        RECT 332.400 297.600 333.600 304.500 ;
        RECT 339.000 303.600 340.200 308.850 ;
        RECT 346.950 307.050 349.050 309.150 ;
        RECT 350.400 307.950 351.600 315.300 ;
        RECT 353.100 309.150 354.900 310.950 ;
        RECT 359.100 309.150 360.900 310.950 ;
        RECT 349.950 305.850 352.050 307.950 ;
        RECT 352.950 307.050 355.050 309.150 ;
        RECT 358.950 307.050 361.050 309.150 ;
        RECT 362.400 307.950 363.600 315.300 ;
        RECT 371.400 314.700 378.900 315.900 ;
        RECT 365.100 309.150 366.900 310.950 ;
        RECT 361.950 305.850 364.050 307.950 ;
        RECT 364.950 307.050 367.050 309.150 ;
        RECT 370.950 308.850 373.050 310.950 ;
        RECT 371.100 307.050 372.900 308.850 ;
        RECT 332.400 291.600 334.200 297.600 ;
        RECT 338.700 291.600 340.500 303.600 ;
        RECT 350.400 297.600 351.600 305.850 ;
        RECT 362.400 297.600 363.600 305.850 ;
        RECT 374.550 297.600 375.600 314.700 ;
        RECT 381.000 310.950 382.050 317.400 ;
        RECT 390.000 316.500 391.200 320.400 ;
        RECT 395.700 317.400 397.500 323.400 ;
        RECT 401.400 320.400 403.200 323.400 ;
        RECT 390.000 315.600 395.100 316.500 ;
        RECT 393.150 314.700 395.100 315.600 ;
        RECT 377.100 309.150 378.900 310.950 ;
        RECT 376.950 307.050 379.050 309.150 ;
        RECT 379.950 308.850 382.050 310.950 ;
        RECT 388.950 308.850 391.050 310.950 ;
        RECT 381.000 303.600 382.050 308.850 ;
        RECT 389.100 307.050 390.900 308.850 ;
        RECT 393.150 306.300 394.050 314.700 ;
        RECT 396.000 310.950 397.200 317.400 ;
        RECT 402.000 316.500 403.200 320.400 ;
        RECT 407.700 317.400 409.500 323.400 ;
        RECT 415.800 317.400 417.600 323.400 ;
        RECT 402.000 315.600 407.100 316.500 ;
        RECT 405.150 314.700 407.100 315.600 ;
        RECT 394.950 308.850 397.200 310.950 ;
        RECT 400.950 308.850 403.050 310.950 ;
        RECT 393.150 305.400 395.100 306.300 ;
        RECT 389.400 304.500 395.100 305.400 ;
        RECT 350.400 291.600 352.200 297.600 ;
        RECT 362.400 291.600 364.200 297.600 ;
        RECT 374.400 291.600 376.200 297.600 ;
        RECT 381.000 291.600 382.800 303.600 ;
        RECT 389.400 297.600 390.600 304.500 ;
        RECT 396.000 303.600 397.200 308.850 ;
        RECT 401.100 307.050 402.900 308.850 ;
        RECT 405.150 306.300 406.050 314.700 ;
        RECT 408.000 310.950 409.200 317.400 ;
        RECT 416.400 315.300 417.600 317.400 ;
        RECT 418.800 318.300 420.600 323.400 ;
        RECT 424.800 318.300 426.600 323.400 ;
        RECT 418.800 316.950 426.600 318.300 ;
        RECT 435.000 316.200 436.800 323.400 ;
        RECT 446.400 320.400 448.200 323.400 ;
        RECT 435.000 315.300 438.600 316.200 ;
        RECT 416.400 314.250 420.150 315.300 ;
        RECT 406.950 308.850 409.200 310.950 ;
        RECT 418.950 310.950 420.150 314.250 ;
        RECT 422.100 312.150 423.900 313.950 ;
        RECT 418.950 308.850 421.050 310.950 ;
        RECT 421.950 310.050 424.050 312.150 ;
        RECT 424.950 308.850 427.050 310.950 ;
        RECT 434.100 309.150 435.900 310.950 ;
        RECT 405.150 305.400 407.100 306.300 ;
        RECT 401.400 304.500 407.100 305.400 ;
        RECT 389.400 291.600 391.200 297.600 ;
        RECT 395.700 291.600 397.500 303.600 ;
        RECT 401.400 297.600 402.600 304.500 ;
        RECT 408.000 303.600 409.200 308.850 ;
        RECT 415.950 305.850 418.050 307.950 ;
        RECT 416.250 304.050 418.050 305.850 ;
        RECT 419.850 303.600 421.050 308.850 ;
        RECT 425.100 307.050 426.900 308.850 ;
        RECT 433.950 307.050 436.050 309.150 ;
        RECT 437.400 307.950 438.600 315.300 ;
        RECT 442.950 311.850 445.050 313.950 ;
        RECT 446.400 312.150 447.600 320.400 ;
        RECT 458.100 315.000 459.900 323.400 ;
        RECT 472.200 316.200 474.000 323.400 ;
        RECT 466.950 315.450 469.050 316.050 ;
        RECT 458.100 313.350 462.300 315.000 ;
        RECT 440.100 309.150 441.900 310.950 ;
        RECT 443.100 310.050 444.900 311.850 ;
        RECT 445.950 310.050 448.050 312.150 ;
        RECT 436.950 305.850 439.050 307.950 ;
        RECT 439.950 307.050 442.050 309.150 ;
        RECT 401.400 291.600 403.200 297.600 ;
        RECT 407.700 291.600 409.500 303.600 ;
        RECT 419.700 291.600 421.500 303.600 ;
        RECT 437.400 297.600 438.600 305.850 ;
        RECT 436.800 291.600 438.600 297.600 ;
        RECT 446.400 297.600 447.600 310.050 ;
        RECT 461.400 309.150 462.300 313.350 ;
        RECT 464.550 314.550 469.050 315.450 ;
        RECT 451.950 305.850 454.050 307.950 ;
        RECT 457.950 305.850 460.050 307.950 ;
        RECT 460.950 307.050 463.050 309.150 ;
        RECT 452.100 304.050 453.900 305.850 ;
        RECT 454.950 302.850 457.050 304.950 ;
        RECT 458.250 304.050 460.050 305.850 ;
        RECT 455.100 301.050 456.900 302.850 ;
        RECT 461.400 298.800 462.300 307.050 ;
        RECT 464.550 303.450 465.450 314.550 ;
        RECT 466.950 313.950 469.050 314.550 ;
        RECT 470.400 315.300 474.000 316.200 ;
        RECT 467.100 309.150 468.900 310.950 ;
        RECT 466.950 307.050 469.050 309.150 ;
        RECT 470.400 307.950 471.600 315.300 ;
        RECT 485.100 315.000 486.900 323.400 ;
        RECT 498.000 316.200 499.800 323.400 ;
        RECT 498.000 315.300 501.600 316.200 ;
        RECT 485.100 313.350 489.300 315.000 ;
        RECT 473.100 309.150 474.900 310.950 ;
        RECT 488.400 309.150 489.300 313.350 ;
        RECT 497.100 309.150 498.900 310.950 ;
        RECT 469.950 305.850 472.050 307.950 ;
        RECT 472.950 307.050 475.050 309.150 ;
        RECT 478.950 305.850 481.050 307.950 ;
        RECT 484.950 305.850 487.050 307.950 ;
        RECT 487.950 307.050 490.050 309.150 ;
        RECT 496.950 307.050 499.050 309.150 ;
        RECT 500.400 307.950 501.600 315.300 ;
        RECT 506.400 315.900 508.200 323.400 ;
        RECT 513.900 318.900 515.700 323.400 ;
        RECT 513.900 317.400 517.050 318.900 ;
        RECT 512.100 315.900 513.900 316.500 ;
        RECT 506.400 314.700 513.900 315.900 ;
        RECT 503.100 309.150 504.900 310.950 ;
        RECT 466.950 303.450 469.050 304.050 ;
        RECT 464.550 302.550 469.050 303.450 ;
        RECT 466.950 301.950 469.050 302.550 ;
        RECT 455.700 297.900 462.300 298.800 ;
        RECT 455.700 297.600 457.200 297.900 ;
        RECT 446.400 291.600 448.200 297.600 ;
        RECT 455.400 291.600 457.200 297.600 ;
        RECT 461.400 297.600 462.300 297.900 ;
        RECT 470.400 297.600 471.600 305.850 ;
        RECT 479.100 304.050 480.900 305.850 ;
        RECT 481.950 302.850 484.050 304.950 ;
        RECT 485.250 304.050 487.050 305.850 ;
        RECT 482.100 301.050 483.900 302.850 ;
        RECT 488.400 298.800 489.300 307.050 ;
        RECT 499.950 305.850 502.050 307.950 ;
        RECT 502.950 307.050 505.050 309.150 ;
        RECT 505.950 308.850 508.050 310.950 ;
        RECT 506.100 307.050 507.900 308.850 ;
        RECT 482.700 297.900 489.300 298.800 ;
        RECT 482.700 297.600 484.200 297.900 ;
        RECT 461.400 291.600 463.200 297.600 ;
        RECT 470.400 291.600 472.200 297.600 ;
        RECT 482.400 291.600 484.200 297.600 ;
        RECT 488.400 297.600 489.300 297.900 ;
        RECT 500.400 297.600 501.600 305.850 ;
        RECT 509.550 297.600 510.600 314.700 ;
        RECT 516.000 310.950 517.050 317.400 ;
        RECT 525.000 316.200 526.800 323.400 ;
        RECT 540.000 319.050 541.800 323.400 ;
        RECT 536.400 317.400 541.800 319.050 ;
        RECT 525.000 315.300 528.600 316.200 ;
        RECT 512.100 309.150 513.900 310.950 ;
        RECT 511.950 307.050 514.050 309.150 ;
        RECT 514.950 308.850 517.050 310.950 ;
        RECT 524.100 309.150 525.900 310.950 ;
        RECT 516.000 303.600 517.050 308.850 ;
        RECT 523.950 307.050 526.050 309.150 ;
        RECT 527.400 307.950 528.600 315.300 ;
        RECT 536.400 310.950 537.300 317.400 ;
        RECT 552.000 316.200 553.800 323.400 ;
        RECT 552.000 315.300 555.600 316.200 ;
        RECT 539.100 312.150 540.900 313.950 ;
        RECT 530.100 309.150 531.900 310.950 ;
        RECT 526.950 305.850 529.050 307.950 ;
        RECT 529.950 307.050 532.050 309.150 ;
        RECT 535.950 308.850 538.050 310.950 ;
        RECT 538.950 310.050 541.050 312.150 ;
        RECT 541.950 311.850 544.050 313.950 ;
        RECT 545.100 312.150 546.900 313.950 ;
        RECT 542.100 310.050 543.900 311.850 ;
        RECT 544.950 310.050 547.050 312.150 ;
        RECT 551.100 309.150 552.900 310.950 ;
        RECT 488.400 291.600 490.200 297.600 ;
        RECT 499.800 291.600 501.600 297.600 ;
        RECT 509.400 291.600 511.200 297.600 ;
        RECT 516.000 291.600 517.800 303.600 ;
        RECT 527.400 297.600 528.600 305.850 ;
        RECT 536.400 303.600 537.300 308.850 ;
        RECT 550.950 307.050 553.050 309.150 ;
        RECT 554.400 307.950 555.600 315.300 ;
        RECT 566.100 315.000 567.900 323.400 ;
        RECT 563.700 313.350 567.900 315.000 ;
        RECT 578.400 320.400 580.200 323.400 ;
        RECT 557.100 309.150 558.900 310.950 ;
        RECT 563.700 309.150 564.600 313.350 ;
        RECT 574.950 311.850 577.050 313.950 ;
        RECT 578.400 312.150 579.600 320.400 ;
        RECT 586.800 317.400 588.600 323.400 ;
        RECT 583.950 315.450 586.050 316.050 ;
        RECT 581.550 314.550 586.050 315.450 ;
        RECT 575.100 310.050 576.900 311.850 ;
        RECT 577.950 310.050 580.050 312.150 ;
        RECT 553.950 305.850 556.050 307.950 ;
        RECT 556.950 307.050 559.050 309.150 ;
        RECT 562.950 307.050 565.050 309.150 ;
        RECT 526.800 291.600 528.600 297.600 ;
        RECT 535.800 291.600 537.600 303.600 ;
        RECT 538.800 302.700 546.600 303.600 ;
        RECT 538.800 291.600 540.600 302.700 ;
        RECT 544.800 291.600 546.600 302.700 ;
        RECT 554.400 297.600 555.600 305.850 ;
        RECT 563.700 298.800 564.600 307.050 ;
        RECT 565.950 305.850 568.050 307.950 ;
        RECT 571.950 305.850 574.050 307.950 ;
        RECT 565.950 304.050 567.750 305.850 ;
        RECT 568.950 302.850 571.050 304.950 ;
        RECT 572.100 304.050 573.900 305.850 ;
        RECT 569.100 301.050 570.900 302.850 ;
        RECT 563.700 297.900 570.300 298.800 ;
        RECT 563.700 297.600 564.600 297.900 ;
        RECT 553.800 291.600 555.600 297.600 ;
        RECT 562.800 291.600 564.600 297.600 ;
        RECT 568.800 297.600 570.300 297.900 ;
        RECT 578.400 297.600 579.600 310.050 ;
        RECT 581.550 304.050 582.450 314.550 ;
        RECT 583.950 313.950 586.050 314.550 ;
        RECT 587.400 315.300 588.600 317.400 ;
        RECT 589.800 318.300 591.600 323.400 ;
        RECT 595.800 318.300 597.600 323.400 ;
        RECT 589.800 316.950 597.600 318.300 ;
        RECT 602.400 318.300 604.200 323.400 ;
        RECT 608.400 318.300 610.200 323.400 ;
        RECT 602.400 316.950 610.200 318.300 ;
        RECT 611.400 317.400 613.200 323.400 ;
        RECT 627.000 319.050 628.800 323.400 ;
        RECT 623.400 317.400 628.800 319.050 ;
        RECT 611.400 315.300 612.600 317.400 ;
        RECT 587.400 314.250 591.150 315.300 ;
        RECT 589.950 310.950 591.150 314.250 ;
        RECT 608.850 314.250 612.600 315.300 ;
        RECT 593.100 312.150 594.900 313.950 ;
        RECT 605.100 312.150 606.900 313.950 ;
        RECT 589.950 308.850 592.050 310.950 ;
        RECT 592.950 310.050 595.050 312.150 ;
        RECT 595.950 308.850 598.050 310.950 ;
        RECT 601.950 308.850 604.050 310.950 ;
        RECT 604.950 310.050 607.050 312.150 ;
        RECT 608.850 310.950 610.050 314.250 ;
        RECT 610.950 312.450 613.050 313.050 ;
        RECT 610.950 311.550 618.450 312.450 ;
        RECT 610.950 310.950 613.050 311.550 ;
        RECT 607.950 308.850 610.050 310.950 ;
        RECT 586.950 305.850 589.050 307.950 ;
        RECT 587.250 304.050 589.050 305.850 ;
        RECT 580.950 301.950 583.050 304.050 ;
        RECT 590.850 303.600 592.050 308.850 ;
        RECT 596.100 307.050 597.900 308.850 ;
        RECT 602.100 307.050 603.900 308.850 ;
        RECT 607.950 303.600 609.150 308.850 ;
        RECT 610.950 305.850 613.050 307.950 ;
        RECT 617.550 307.050 618.450 311.550 ;
        RECT 623.400 310.950 624.300 317.400 ;
        RECT 644.100 315.000 645.900 323.400 ;
        RECT 659.100 315.000 660.900 323.400 ;
        RECT 675.000 319.050 676.800 323.400 ;
        RECT 626.100 312.150 627.900 313.950 ;
        RECT 622.950 308.850 625.050 310.950 ;
        RECT 625.950 310.050 628.050 312.150 ;
        RECT 628.950 311.850 631.050 313.950 ;
        RECT 632.100 312.150 633.900 313.950 ;
        RECT 641.700 313.350 645.900 315.000 ;
        RECT 656.700 313.350 660.900 315.000 ;
        RECT 671.400 317.400 676.800 319.050 ;
        RECT 629.100 310.050 630.900 311.850 ;
        RECT 631.950 310.050 634.050 312.150 ;
        RECT 641.700 309.150 642.600 313.350 ;
        RECT 656.700 309.150 657.600 313.350 ;
        RECT 671.400 310.950 672.300 317.400 ;
        RECT 692.100 315.000 693.900 323.400 ;
        RECT 706.200 316.200 708.000 323.400 ;
        RECT 674.100 312.150 675.900 313.950 ;
        RECT 610.950 304.050 612.750 305.850 ;
        RECT 616.950 304.950 619.050 307.050 ;
        RECT 623.400 303.600 624.300 308.850 ;
        RECT 640.950 307.050 643.050 309.150 ;
        RECT 568.800 291.600 570.600 297.600 ;
        RECT 578.400 291.600 580.200 297.600 ;
        RECT 590.700 291.600 592.500 303.600 ;
        RECT 607.500 291.600 609.300 303.600 ;
        RECT 622.800 291.600 624.600 303.600 ;
        RECT 625.800 302.700 633.600 303.600 ;
        RECT 625.800 291.600 627.600 302.700 ;
        RECT 631.800 291.600 633.600 302.700 ;
        RECT 641.700 298.800 642.600 307.050 ;
        RECT 643.950 305.850 646.050 307.950 ;
        RECT 649.950 305.850 652.050 307.950 ;
        RECT 655.950 307.050 658.050 309.150 ;
        RECT 670.950 308.850 673.050 310.950 ;
        RECT 673.950 310.050 676.050 312.150 ;
        RECT 676.950 311.850 679.050 313.950 ;
        RECT 680.100 312.150 681.900 313.950 ;
        RECT 689.700 313.350 693.900 315.000 ;
        RECT 704.400 315.300 708.000 316.200 ;
        RECT 677.100 310.050 678.900 311.850 ;
        RECT 679.950 310.050 682.050 312.150 ;
        RECT 689.700 309.150 690.600 313.350 ;
        RECT 701.100 309.150 702.900 310.950 ;
        RECT 643.950 304.050 645.750 305.850 ;
        RECT 646.950 302.850 649.050 304.950 ;
        RECT 650.100 304.050 651.900 305.850 ;
        RECT 647.100 301.050 648.900 302.850 ;
        RECT 656.700 298.800 657.600 307.050 ;
        RECT 658.950 305.850 661.050 307.950 ;
        RECT 664.950 305.850 667.050 307.950 ;
        RECT 658.950 304.050 660.750 305.850 ;
        RECT 661.950 302.850 664.050 304.950 ;
        RECT 665.100 304.050 666.900 305.850 ;
        RECT 671.400 303.600 672.300 308.850 ;
        RECT 688.950 307.050 691.050 309.150 ;
        RECT 662.100 301.050 663.900 302.850 ;
        RECT 641.700 297.900 648.300 298.800 ;
        RECT 641.700 297.600 642.600 297.900 ;
        RECT 640.800 291.600 642.600 297.600 ;
        RECT 646.800 297.600 648.300 297.900 ;
        RECT 656.700 297.900 663.300 298.800 ;
        RECT 656.700 297.600 657.600 297.900 ;
        RECT 646.800 291.600 648.600 297.600 ;
        RECT 655.800 291.600 657.600 297.600 ;
        RECT 661.800 297.600 663.300 297.900 ;
        RECT 661.800 291.600 663.600 297.600 ;
        RECT 670.800 291.600 672.600 303.600 ;
        RECT 673.800 302.700 681.600 303.600 ;
        RECT 673.800 291.600 675.600 302.700 ;
        RECT 679.800 291.600 681.600 302.700 ;
        RECT 689.700 298.800 690.600 307.050 ;
        RECT 691.950 305.850 694.050 307.950 ;
        RECT 697.950 305.850 700.050 307.950 ;
        RECT 700.950 307.050 703.050 309.150 ;
        RECT 704.400 307.950 705.600 315.300 ;
        RECT 719.100 315.000 720.900 323.400 ;
        RECT 733.200 319.050 735.000 323.400 ;
        RECT 751.200 319.050 753.000 323.400 ;
        RECT 733.200 317.400 738.600 319.050 ;
        RECT 751.200 317.400 756.600 319.050 ;
        RECT 716.700 313.350 720.900 315.000 ;
        RECT 707.100 309.150 708.900 310.950 ;
        RECT 716.700 309.150 717.600 313.350 ;
        RECT 728.100 312.150 729.900 313.950 ;
        RECT 727.950 310.050 730.050 312.150 ;
        RECT 730.950 311.850 733.050 313.950 ;
        RECT 734.100 312.150 735.900 313.950 ;
        RECT 731.100 310.050 732.900 311.850 ;
        RECT 733.950 310.050 736.050 312.150 ;
        RECT 737.700 310.950 738.600 317.400 ;
        RECT 746.100 312.150 747.900 313.950 ;
        RECT 703.950 305.850 706.050 307.950 ;
        RECT 706.950 307.050 709.050 309.150 ;
        RECT 715.950 307.050 718.050 309.150 ;
        RECT 736.950 308.850 739.050 310.950 ;
        RECT 745.950 310.050 748.050 312.150 ;
        RECT 748.950 311.850 751.050 313.950 ;
        RECT 752.100 312.150 753.900 313.950 ;
        RECT 749.100 310.050 750.900 311.850 ;
        RECT 751.950 310.050 754.050 312.150 ;
        RECT 755.700 310.950 756.600 317.400 ;
        RECT 754.950 308.850 757.050 310.950 ;
        RECT 691.950 304.050 693.750 305.850 ;
        RECT 694.950 302.850 697.050 304.950 ;
        RECT 698.100 304.050 699.900 305.850 ;
        RECT 695.100 301.050 696.900 302.850 ;
        RECT 689.700 297.900 696.300 298.800 ;
        RECT 689.700 297.600 690.600 297.900 ;
        RECT 688.800 291.600 690.600 297.600 ;
        RECT 694.800 297.600 696.300 297.900 ;
        RECT 704.400 297.600 705.600 305.850 ;
        RECT 716.700 298.800 717.600 307.050 ;
        RECT 718.950 305.850 721.050 307.950 ;
        RECT 724.950 305.850 727.050 307.950 ;
        RECT 718.950 304.050 720.750 305.850 ;
        RECT 721.950 302.850 724.050 304.950 ;
        RECT 725.100 304.050 726.900 305.850 ;
        RECT 737.700 303.600 738.600 308.850 ;
        RECT 755.700 303.600 756.600 308.850 ;
        RECT 722.100 301.050 723.900 302.850 ;
        RECT 728.400 302.700 736.200 303.600 ;
        RECT 716.700 297.900 723.300 298.800 ;
        RECT 716.700 297.600 717.600 297.900 ;
        RECT 694.800 291.600 696.600 297.600 ;
        RECT 704.400 291.600 706.200 297.600 ;
        RECT 715.800 291.600 717.600 297.600 ;
        RECT 721.800 297.600 723.300 297.900 ;
        RECT 721.800 291.600 723.600 297.600 ;
        RECT 728.400 291.600 730.200 302.700 ;
        RECT 734.400 291.600 736.200 302.700 ;
        RECT 737.400 291.600 739.200 303.600 ;
        RECT 746.400 302.700 754.200 303.600 ;
        RECT 746.400 291.600 748.200 302.700 ;
        RECT 752.400 291.600 754.200 302.700 ;
        RECT 755.400 291.600 757.200 303.600 ;
        RECT 8.700 275.400 10.500 287.400 ;
        RECT 22.800 281.400 24.600 287.400 ;
        RECT 35.400 281.400 37.200 287.400 ;
        RECT 5.250 273.150 7.050 274.950 ;
        RECT 4.950 271.050 7.050 273.150 ;
        RECT 8.850 270.150 10.050 275.400 ;
        RECT 23.400 273.150 24.600 281.400 ;
        RECT 35.700 281.100 37.200 281.400 ;
        RECT 41.400 281.400 43.200 287.400 ;
        RECT 52.800 281.400 54.600 287.400 ;
        RECT 62.400 281.400 64.200 287.400 ;
        RECT 41.400 281.100 42.300 281.400 ;
        RECT 35.700 280.200 42.300 281.100 ;
        RECT 35.100 276.150 36.900 277.950 ;
        RECT 32.100 273.150 33.900 274.950 ;
        RECT 34.950 274.050 37.050 276.150 ;
        RECT 38.250 273.150 40.050 274.950 ;
        RECT 14.100 270.150 15.900 271.950 ;
        RECT 7.950 268.050 10.050 270.150 ;
        RECT 7.950 264.750 9.150 268.050 ;
        RECT 10.950 266.850 13.050 268.950 ;
        RECT 13.950 268.050 16.050 270.150 ;
        RECT 19.950 269.850 22.050 271.950 ;
        RECT 22.950 271.050 25.050 273.150 ;
        RECT 20.100 268.050 21.900 269.850 ;
        RECT 11.100 265.050 12.900 266.850 ;
        RECT 5.400 263.700 9.150 264.750 ;
        RECT 23.400 263.700 24.600 271.050 ;
        RECT 25.950 269.850 28.050 271.950 ;
        RECT 31.950 271.050 34.050 273.150 ;
        RECT 37.950 271.050 40.050 273.150 ;
        RECT 41.400 271.950 42.300 280.200 ;
        RECT 53.400 273.150 54.600 281.400 ;
        RECT 62.700 281.100 64.200 281.400 ;
        RECT 68.400 281.400 70.200 287.400 ;
        RECT 68.400 281.100 69.300 281.400 ;
        RECT 62.700 280.200 69.300 281.100 ;
        RECT 62.100 276.150 63.900 277.950 ;
        RECT 59.100 273.150 60.900 274.950 ;
        RECT 61.950 274.050 64.050 276.150 ;
        RECT 65.250 273.150 67.050 274.950 ;
        RECT 40.950 269.850 43.050 271.950 ;
        RECT 49.950 269.850 52.050 271.950 ;
        RECT 52.950 271.050 55.050 273.150 ;
        RECT 26.100 268.050 27.900 269.850 ;
        RECT 41.400 265.650 42.300 269.850 ;
        RECT 50.100 268.050 51.900 269.850 ;
        RECT 5.400 261.600 6.600 263.700 ;
        RECT 21.000 262.800 24.600 263.700 ;
        RECT 38.100 264.000 42.300 265.650 ;
        RECT 4.800 255.600 6.600 261.600 ;
        RECT 7.800 260.700 15.600 262.050 ;
        RECT 7.800 255.600 9.600 260.700 ;
        RECT 13.800 255.600 15.600 260.700 ;
        RECT 21.000 255.600 22.800 262.800 ;
        RECT 38.100 255.600 39.900 264.000 ;
        RECT 53.400 263.700 54.600 271.050 ;
        RECT 55.950 269.850 58.050 271.950 ;
        RECT 58.950 271.050 61.050 273.150 ;
        RECT 64.950 271.050 67.050 273.150 ;
        RECT 68.400 271.950 69.300 280.200 ;
        RECT 76.800 275.400 78.600 287.400 ;
        RECT 79.800 276.300 81.600 287.400 ;
        RECT 85.800 276.300 87.600 287.400 ;
        RECT 79.800 275.400 87.600 276.300 ;
        RECT 95.400 281.400 97.200 287.400 ;
        RECT 67.950 269.850 70.050 271.950 ;
        RECT 77.400 270.150 78.300 275.400 ;
        RECT 95.400 273.150 96.600 281.400 ;
        RECT 111.600 275.400 113.400 287.400 ;
        RECT 125.700 275.400 127.500 287.400 ;
        RECT 138.900 275.400 142.200 287.400 ;
        RECT 154.800 275.400 156.600 287.400 ;
        RECT 157.800 276.300 159.600 287.400 ;
        RECT 163.800 276.300 165.600 287.400 ;
        RECT 157.800 275.400 165.600 276.300 ;
        RECT 171.600 275.400 173.400 287.400 ;
        RECT 183.600 275.400 185.400 287.400 ;
        RECT 111.600 274.350 114.000 275.400 ;
        RECT 56.100 268.050 57.900 269.850 ;
        RECT 68.400 265.650 69.300 269.850 ;
        RECT 76.950 268.050 79.050 270.150 ;
        RECT 91.950 269.850 94.050 271.950 ;
        RECT 94.950 271.050 97.050 273.150 ;
        RECT 51.000 262.800 54.600 263.700 ;
        RECT 65.100 264.000 69.300 265.650 ;
        RECT 51.000 255.600 52.800 262.800 ;
        RECT 65.100 255.600 66.900 264.000 ;
        RECT 77.400 261.600 78.300 268.050 ;
        RECT 79.950 266.850 82.050 268.950 ;
        RECT 83.100 267.150 84.900 268.950 ;
        RECT 80.100 265.050 81.900 266.850 ;
        RECT 82.950 265.050 85.050 267.150 ;
        RECT 85.950 266.850 88.050 268.950 ;
        RECT 92.100 268.050 93.900 269.850 ;
        RECT 86.100 265.050 87.900 266.850 ;
        RECT 95.400 263.700 96.600 271.050 ;
        RECT 97.950 269.850 100.050 271.950 ;
        RECT 110.100 270.150 111.900 271.950 ;
        RECT 98.100 268.050 99.900 269.850 ;
        RECT 109.950 268.050 112.050 270.150 ;
        RECT 112.950 267.150 114.000 274.350 ;
        RECT 122.250 273.150 124.050 274.950 ;
        RECT 116.100 270.150 117.900 271.950 ;
        RECT 121.950 271.050 124.050 273.150 ;
        RECT 125.850 270.150 127.050 275.400 ;
        RECT 131.100 270.150 132.900 271.950 ;
        RECT 134.100 270.150 135.900 271.950 ;
        RECT 140.400 270.150 141.600 275.400 ;
        RECT 145.950 270.150 147.750 271.950 ;
        RECT 155.400 270.150 156.300 275.400 ;
        RECT 171.000 274.350 173.400 275.400 ;
        RECT 183.000 274.350 185.400 275.400 ;
        RECT 197.400 281.400 199.200 287.400 ;
        RECT 209.400 281.400 211.200 287.400 ;
        RECT 224.400 281.400 226.200 287.400 ;
        RECT 236.400 281.400 238.200 287.400 ;
        RECT 167.100 270.150 168.900 271.950 ;
        RECT 115.950 268.050 118.050 270.150 ;
        RECT 124.950 268.050 127.050 270.150 ;
        RECT 112.950 265.050 115.050 267.150 ;
        RECT 95.400 262.800 99.000 263.700 ;
        RECT 77.400 259.950 82.800 261.600 ;
        RECT 81.000 255.600 82.800 259.950 ;
        RECT 97.200 255.600 99.000 262.800 ;
        RECT 112.950 258.600 114.000 265.050 ;
        RECT 124.950 264.750 126.150 268.050 ;
        RECT 127.950 266.850 130.050 268.950 ;
        RECT 130.950 268.050 133.050 270.150 ;
        RECT 133.950 268.050 136.050 270.150 ;
        RECT 136.950 266.850 139.050 268.950 ;
        RECT 139.950 268.050 142.050 270.150 ;
        RECT 128.100 265.050 129.900 266.850 ;
        RECT 137.100 265.050 138.900 266.850 ;
        RECT 122.400 263.700 126.150 264.750 ;
        RECT 140.400 264.150 141.600 268.050 ;
        RECT 142.950 266.850 145.050 268.950 ;
        RECT 145.950 268.050 148.050 270.150 ;
        RECT 154.950 268.050 157.050 270.150 ;
        RECT 142.500 265.050 144.300 266.850 ;
        RECT 122.400 261.600 123.600 263.700 ;
        RECT 140.400 263.100 144.600 264.150 ;
        RECT 112.800 255.600 114.600 258.600 ;
        RECT 121.800 255.600 123.600 261.600 ;
        RECT 124.800 260.700 132.600 262.050 ;
        RECT 124.800 255.600 126.600 260.700 ;
        RECT 130.800 255.600 132.600 260.700 ;
        RECT 134.400 261.000 142.200 261.900 ;
        RECT 143.700 261.600 144.600 263.100 ;
        RECT 155.400 261.600 156.300 268.050 ;
        RECT 157.950 266.850 160.050 268.950 ;
        RECT 161.100 267.150 162.900 268.950 ;
        RECT 158.100 265.050 159.900 266.850 ;
        RECT 160.950 265.050 163.050 267.150 ;
        RECT 163.950 266.850 166.050 268.950 ;
        RECT 166.950 268.050 169.050 270.150 ;
        RECT 171.000 267.150 172.050 274.350 ;
        RECT 173.100 270.150 174.900 271.950 ;
        RECT 179.100 270.150 180.900 271.950 ;
        RECT 172.950 268.050 175.050 270.150 ;
        RECT 178.950 268.050 181.050 270.150 ;
        RECT 183.000 267.150 184.050 274.350 ;
        RECT 197.400 273.150 198.600 281.400 ;
        RECT 209.400 273.150 210.600 281.400 ;
        RECT 224.400 273.150 225.600 281.400 ;
        RECT 236.400 273.150 237.600 281.400 ;
        RECT 248.400 275.400 250.200 287.400 ;
        RECT 259.800 275.400 261.600 287.400 ;
        RECT 262.800 276.300 264.600 287.400 ;
        RECT 268.800 276.300 270.600 287.400 ;
        RECT 262.800 275.400 270.600 276.300 ;
        RECT 277.500 275.400 279.300 287.400 ;
        RECT 283.800 281.400 285.600 287.400 ;
        RECT 185.100 270.150 186.900 271.950 ;
        RECT 184.950 268.050 187.050 270.150 ;
        RECT 193.950 269.850 196.050 271.950 ;
        RECT 196.950 271.050 199.050 273.150 ;
        RECT 194.100 268.050 195.900 269.850 ;
        RECT 164.100 265.050 165.900 266.850 ;
        RECT 169.950 265.050 172.050 267.150 ;
        RECT 181.950 265.050 184.050 267.150 ;
        RECT 134.400 255.600 136.200 261.000 ;
        RECT 140.400 256.500 142.200 261.000 ;
        RECT 143.400 257.400 145.200 261.600 ;
        RECT 146.400 256.500 148.200 261.600 ;
        RECT 155.400 259.950 160.800 261.600 ;
        RECT 140.400 255.600 148.200 256.500 ;
        RECT 159.000 255.600 160.800 259.950 ;
        RECT 171.000 258.600 172.050 265.050 ;
        RECT 183.000 258.600 184.050 265.050 ;
        RECT 197.400 263.700 198.600 271.050 ;
        RECT 199.950 269.850 202.050 271.950 ;
        RECT 205.950 269.850 208.050 271.950 ;
        RECT 208.950 271.050 211.050 273.150 ;
        RECT 200.100 268.050 201.900 269.850 ;
        RECT 206.100 268.050 207.900 269.850 ;
        RECT 209.400 263.700 210.600 271.050 ;
        RECT 211.950 269.850 214.050 271.950 ;
        RECT 220.950 269.850 223.050 271.950 ;
        RECT 223.950 271.050 226.050 273.150 ;
        RECT 212.100 268.050 213.900 269.850 ;
        RECT 221.100 268.050 222.900 269.850 ;
        RECT 224.400 263.700 225.600 271.050 ;
        RECT 226.950 269.850 229.050 271.950 ;
        RECT 232.950 269.850 235.050 271.950 ;
        RECT 235.950 271.050 238.050 273.150 ;
        RECT 227.100 268.050 228.900 269.850 ;
        RECT 233.100 268.050 234.900 269.850 ;
        RECT 236.400 263.700 237.600 271.050 ;
        RECT 238.950 269.850 241.050 271.950 ;
        RECT 248.400 270.150 249.600 275.400 ;
        RECT 260.400 270.150 261.300 275.400 ;
        RECT 277.800 270.150 279.000 275.400 ;
        RECT 284.400 274.500 285.600 281.400 ;
        RECT 292.800 275.400 294.600 287.400 ;
        RECT 302.400 275.400 304.200 287.400 ;
        RECT 310.800 275.400 312.600 287.400 ;
        RECT 279.900 273.600 285.600 274.500 ;
        RECT 279.900 272.700 281.850 273.600 ;
        RECT 239.100 268.050 240.900 269.850 ;
        RECT 244.950 266.850 247.050 268.950 ;
        RECT 247.950 268.050 250.050 270.150 ;
        RECT 259.950 268.050 262.050 270.150 ;
        RECT 245.100 265.050 246.900 266.850 ;
        RECT 197.400 262.800 201.000 263.700 ;
        RECT 209.400 262.800 213.000 263.700 ;
        RECT 224.400 262.800 228.000 263.700 ;
        RECT 236.400 262.800 240.000 263.700 ;
        RECT 170.400 255.600 172.200 258.600 ;
        RECT 182.400 255.600 184.200 258.600 ;
        RECT 199.200 255.600 201.000 262.800 ;
        RECT 211.200 255.600 213.000 262.800 ;
        RECT 226.200 255.600 228.000 262.800 ;
        RECT 238.200 255.600 240.000 262.800 ;
        RECT 248.400 261.600 249.600 268.050 ;
        RECT 260.400 261.600 261.300 268.050 ;
        RECT 262.950 266.850 265.050 268.950 ;
        RECT 266.100 267.150 267.900 268.950 ;
        RECT 263.100 265.050 264.900 266.850 ;
        RECT 265.950 265.050 268.050 267.150 ;
        RECT 268.950 266.850 271.050 268.950 ;
        RECT 277.800 268.050 280.050 270.150 ;
        RECT 269.100 265.050 270.900 266.850 ;
        RECT 277.800 261.600 279.000 268.050 ;
        RECT 280.950 264.300 281.850 272.700 ;
        RECT 284.100 270.150 285.900 271.950 ;
        RECT 283.950 268.050 286.050 270.150 ;
        RECT 292.950 268.950 294.300 275.400 ;
        RECT 302.400 270.150 303.600 275.400 ;
        RECT 311.400 270.150 312.600 275.400 ;
        RECT 317.400 281.400 319.200 287.400 ;
        RECT 317.400 274.500 318.600 281.400 ;
        RECT 323.700 275.400 325.500 287.400 ;
        RECT 331.800 281.400 333.600 287.400 ;
        RECT 332.700 281.100 333.600 281.400 ;
        RECT 337.800 281.400 339.600 287.400 ;
        RECT 349.800 281.400 351.600 287.400 ;
        RECT 337.800 281.100 339.300 281.400 ;
        RECT 332.700 280.200 339.300 281.100 ;
        RECT 317.400 273.600 323.100 274.500 ;
        RECT 321.150 272.700 323.100 273.600 ;
        RECT 317.100 270.150 318.900 271.950 ;
        RECT 289.950 266.850 294.300 268.950 ;
        RECT 295.950 266.850 298.050 268.950 ;
        RECT 298.950 266.850 301.050 268.950 ;
        RECT 301.950 268.050 304.050 270.150 ;
        RECT 310.950 268.050 313.050 270.150 ;
        RECT 279.900 263.400 281.850 264.300 ;
        RECT 279.900 262.500 285.000 263.400 ;
        RECT 248.400 255.600 250.200 261.600 ;
        RECT 260.400 259.950 265.800 261.600 ;
        RECT 264.000 255.600 265.800 259.950 ;
        RECT 277.500 255.600 279.300 261.600 ;
        RECT 283.800 258.600 285.000 262.500 ;
        RECT 292.950 261.600 294.300 266.850 ;
        RECT 296.100 265.050 297.900 266.850 ;
        RECT 299.100 265.050 300.900 266.850 ;
        RECT 302.400 261.600 303.600 268.050 ;
        RECT 311.400 261.600 312.600 268.050 ;
        RECT 313.950 266.850 316.050 268.950 ;
        RECT 316.950 268.050 319.050 270.150 ;
        RECT 314.100 265.050 315.900 266.850 ;
        RECT 321.150 264.300 322.050 272.700 ;
        RECT 324.000 270.150 325.200 275.400 ;
        RECT 332.700 271.950 333.600 280.200 ;
        RECT 340.950 279.450 343.050 280.050 ;
        RECT 340.950 278.550 345.450 279.450 ;
        RECT 340.950 277.950 343.050 278.550 ;
        RECT 338.100 276.150 339.900 277.950 ;
        RECT 334.950 273.150 336.750 274.950 ;
        RECT 337.950 274.050 340.050 276.150 ;
        RECT 341.100 273.150 342.900 274.950 ;
        RECT 322.950 268.050 325.200 270.150 ;
        RECT 331.950 269.850 334.050 271.950 ;
        RECT 334.950 271.050 337.050 273.150 ;
        RECT 340.950 271.050 343.050 273.150 ;
        RECT 321.150 263.400 323.100 264.300 ;
        RECT 283.800 255.600 285.600 258.600 ;
        RECT 292.800 255.600 294.600 261.600 ;
        RECT 302.400 255.600 304.200 261.600 ;
        RECT 310.800 255.600 312.600 261.600 ;
        RECT 318.000 262.500 323.100 263.400 ;
        RECT 318.000 258.600 319.200 262.500 ;
        RECT 324.000 261.600 325.200 268.050 ;
        RECT 332.700 265.650 333.600 269.850 ;
        RECT 337.950 267.450 340.050 268.050 ;
        RECT 344.550 267.450 345.450 278.550 ;
        RECT 350.400 273.150 351.600 281.400 ;
        RECT 352.950 276.450 355.050 277.050 ;
        RECT 352.950 275.550 357.450 276.450 ;
        RECT 352.950 274.950 355.050 275.550 ;
        RECT 346.950 269.850 349.050 271.950 ;
        RECT 349.950 271.050 352.050 273.150 ;
        RECT 347.100 268.050 348.900 269.850 ;
        RECT 337.950 266.550 345.450 267.450 ;
        RECT 337.950 265.950 340.050 266.550 ;
        RECT 332.700 264.000 336.900 265.650 ;
        RECT 317.400 255.600 319.200 258.600 ;
        RECT 323.700 255.600 325.500 261.600 ;
        RECT 335.100 255.600 336.900 264.000 ;
        RECT 350.400 263.700 351.600 271.050 ;
        RECT 352.950 269.850 355.050 271.950 ;
        RECT 353.100 268.050 354.900 269.850 ;
        RECT 348.000 262.800 351.600 263.700 ;
        RECT 352.950 264.450 355.050 265.050 ;
        RECT 356.550 264.450 357.450 275.550 ;
        RECT 361.800 275.400 363.600 287.400 ;
        RECT 364.800 276.300 366.600 287.400 ;
        RECT 370.800 276.300 372.600 287.400 ;
        RECT 364.800 275.400 372.600 276.300 ;
        RECT 377.400 281.400 379.200 287.400 ;
        RECT 386.400 281.400 388.200 287.400 ;
        RECT 362.400 270.150 363.300 275.400 ;
        RECT 377.400 273.150 378.600 281.400 ;
        RECT 386.400 274.500 387.600 281.400 ;
        RECT 392.700 275.400 394.500 287.400 ;
        RECT 400.200 275.400 402.000 287.400 ;
        RECT 406.800 281.400 408.600 287.400 ;
        RECT 386.400 273.600 392.100 274.500 ;
        RECT 361.950 268.050 364.050 270.150 ;
        RECT 373.950 269.850 376.050 271.950 ;
        RECT 376.950 271.050 379.050 273.150 ;
        RECT 390.150 272.700 392.100 273.600 ;
        RECT 352.950 263.550 357.450 264.450 ;
        RECT 352.950 262.950 355.050 263.550 ;
        RECT 348.000 255.600 349.800 262.800 ;
        RECT 362.400 261.600 363.300 268.050 ;
        RECT 364.950 266.850 367.050 268.950 ;
        RECT 368.100 267.150 369.900 268.950 ;
        RECT 365.100 265.050 366.900 266.850 ;
        RECT 367.950 265.050 370.050 267.150 ;
        RECT 370.950 266.850 373.050 268.950 ;
        RECT 374.100 268.050 375.900 269.850 ;
        RECT 371.100 265.050 372.900 266.850 ;
        RECT 377.400 263.700 378.600 271.050 ;
        RECT 379.950 269.850 382.050 271.950 ;
        RECT 386.100 270.150 387.900 271.950 ;
        RECT 380.100 268.050 381.900 269.850 ;
        RECT 385.950 268.050 388.050 270.150 ;
        RECT 390.150 264.300 391.050 272.700 ;
        RECT 393.000 270.150 394.200 275.400 ;
        RECT 391.950 268.050 394.200 270.150 ;
        RECT 377.400 262.800 381.000 263.700 ;
        RECT 390.150 263.400 392.100 264.300 ;
        RECT 362.400 259.950 367.800 261.600 ;
        RECT 366.000 255.600 367.800 259.950 ;
        RECT 379.200 255.600 381.000 262.800 ;
        RECT 387.000 262.500 392.100 263.400 ;
        RECT 387.000 258.600 388.200 262.500 ;
        RECT 393.000 261.600 394.200 268.050 ;
        RECT 400.950 270.150 402.000 275.400 ;
        RECT 400.950 268.050 403.050 270.150 ;
        RECT 403.950 269.850 406.050 271.950 ;
        RECT 404.100 268.050 405.900 269.850 ;
        RECT 400.950 261.600 402.000 268.050 ;
        RECT 407.400 264.300 408.450 281.400 ;
        RECT 416.400 275.400 418.200 287.400 ;
        RECT 425.400 281.400 427.200 287.400 ;
        RECT 410.100 270.150 411.900 271.950 ;
        RECT 416.400 270.150 417.600 275.400 ;
        RECT 425.400 274.500 426.600 281.400 ;
        RECT 431.700 275.400 433.500 287.400 ;
        RECT 439.200 275.400 441.000 287.400 ;
        RECT 445.800 281.400 447.600 287.400 ;
        RECT 455.400 281.400 457.200 287.400 ;
        RECT 425.400 273.600 431.100 274.500 ;
        RECT 429.150 272.700 431.100 273.600 ;
        RECT 425.100 270.150 426.900 271.950 ;
        RECT 409.950 268.050 412.050 270.150 ;
        RECT 412.950 266.850 415.050 268.950 ;
        RECT 415.950 268.050 418.050 270.150 ;
        RECT 424.950 268.050 427.050 270.150 ;
        RECT 413.100 265.050 414.900 266.850 ;
        RECT 404.100 263.100 411.600 264.300 ;
        RECT 404.100 262.500 405.900 263.100 ;
        RECT 386.400 255.600 388.200 258.600 ;
        RECT 392.700 255.600 394.500 261.600 ;
        RECT 400.950 260.100 404.100 261.600 ;
        RECT 402.300 255.600 404.100 260.100 ;
        RECT 409.800 255.600 411.600 263.100 ;
        RECT 416.400 261.600 417.600 268.050 ;
        RECT 429.150 264.300 430.050 272.700 ;
        RECT 432.000 270.150 433.200 275.400 ;
        RECT 430.950 268.050 433.200 270.150 ;
        RECT 429.150 263.400 431.100 264.300 ;
        RECT 426.000 262.500 431.100 263.400 ;
        RECT 416.400 255.600 418.200 261.600 ;
        RECT 426.000 258.600 427.200 262.500 ;
        RECT 432.000 261.600 433.200 268.050 ;
        RECT 439.950 270.150 441.000 275.400 ;
        RECT 439.950 268.050 442.050 270.150 ;
        RECT 442.950 269.850 445.050 271.950 ;
        RECT 443.100 268.050 444.900 269.850 ;
        RECT 439.950 261.600 441.000 268.050 ;
        RECT 446.400 264.300 447.450 281.400 ;
        RECT 449.100 270.150 450.900 271.950 ;
        RECT 452.100 270.150 453.900 271.950 ;
        RECT 448.950 268.050 451.050 270.150 ;
        RECT 451.950 268.050 454.050 270.150 ;
        RECT 455.550 264.300 456.600 281.400 ;
        RECT 462.000 275.400 463.800 287.400 ;
        RECT 472.800 286.500 480.600 287.400 ;
        RECT 472.800 275.400 474.600 286.500 ;
        RECT 457.950 269.850 460.050 271.950 ;
        RECT 462.000 270.150 463.050 275.400 ;
        RECT 475.800 274.500 477.600 285.600 ;
        RECT 478.800 276.600 480.600 286.500 ;
        RECT 484.800 276.600 486.600 287.400 ;
        RECT 478.800 275.700 486.600 276.600 ;
        RECT 490.200 275.400 492.000 287.400 ;
        RECT 496.800 281.400 498.600 287.400 ;
        RECT 506.400 281.400 508.200 287.400 ;
        RECT 475.800 273.600 479.850 274.500 ;
        RECT 473.100 270.150 474.900 271.950 ;
        RECT 478.950 270.150 479.850 273.600 ;
        RECT 484.950 270.150 486.750 271.950 ;
        RECT 490.950 270.150 492.000 275.400 ;
        RECT 458.100 268.050 459.900 269.850 ;
        RECT 460.950 268.050 463.050 270.150 ;
        RECT 472.950 268.050 475.050 270.150 ;
        RECT 443.100 263.100 450.600 264.300 ;
        RECT 443.100 262.500 444.900 263.100 ;
        RECT 425.400 255.600 427.200 258.600 ;
        RECT 431.700 255.600 433.500 261.600 ;
        RECT 439.950 260.100 443.100 261.600 ;
        RECT 441.300 255.600 443.100 260.100 ;
        RECT 448.800 255.600 450.600 263.100 ;
        RECT 452.400 263.100 459.900 264.300 ;
        RECT 452.400 255.600 454.200 263.100 ;
        RECT 458.100 262.500 459.900 263.100 ;
        RECT 462.000 261.600 463.050 268.050 ;
        RECT 475.950 266.850 478.050 268.950 ;
        RECT 478.950 268.050 481.050 270.150 ;
        RECT 476.250 265.050 478.050 266.850 ;
        RECT 463.950 264.450 466.050 265.050 ;
        RECT 472.950 264.450 475.050 265.050 ;
        RECT 463.950 263.550 475.050 264.450 ;
        RECT 463.950 262.950 466.050 263.550 ;
        RECT 472.950 262.950 475.050 263.550 ;
        RECT 459.900 260.100 463.050 261.600 ;
        RECT 480.000 261.600 481.050 268.050 ;
        RECT 481.950 266.850 484.050 268.950 ;
        RECT 484.950 268.050 487.050 270.150 ;
        RECT 490.950 268.050 493.050 270.150 ;
        RECT 493.950 269.850 496.050 271.950 ;
        RECT 494.100 268.050 495.900 269.850 ;
        RECT 481.950 265.050 483.750 266.850 ;
        RECT 490.950 261.600 492.000 268.050 ;
        RECT 497.400 264.300 498.450 281.400 ;
        RECT 506.400 273.150 507.600 281.400 ;
        RECT 520.500 275.400 522.300 287.400 ;
        RECT 533.400 281.400 535.200 287.400 ;
        RECT 500.100 270.150 501.900 271.950 ;
        RECT 499.950 268.050 502.050 270.150 ;
        RECT 502.950 269.850 505.050 271.950 ;
        RECT 505.950 271.050 508.050 273.150 ;
        RECT 503.100 268.050 504.900 269.850 ;
        RECT 494.100 263.100 501.600 264.300 ;
        RECT 494.100 262.500 495.900 263.100 ;
        RECT 459.900 255.600 461.700 260.100 ;
        RECT 480.000 255.600 481.800 261.600 ;
        RECT 490.950 260.100 494.100 261.600 ;
        RECT 492.300 255.600 494.100 260.100 ;
        RECT 499.800 255.600 501.600 263.100 ;
        RECT 506.400 263.700 507.600 271.050 ;
        RECT 508.950 269.850 511.050 271.950 ;
        RECT 515.100 270.150 516.900 271.950 ;
        RECT 520.950 270.150 522.150 275.400 ;
        RECT 526.950 274.950 529.050 277.050 ;
        RECT 523.950 273.150 525.750 274.950 ;
        RECT 523.950 271.050 526.050 273.150 ;
        RECT 509.100 268.050 510.900 269.850 ;
        RECT 514.950 268.050 517.050 270.150 ;
        RECT 517.950 266.850 520.050 268.950 ;
        RECT 520.950 268.050 523.050 270.150 ;
        RECT 518.100 265.050 519.900 266.850 ;
        RECT 521.850 264.750 523.050 268.050 ;
        RECT 523.950 267.450 526.050 268.050 ;
        RECT 527.550 267.450 528.450 274.950 ;
        RECT 533.400 273.150 534.600 281.400 ;
        RECT 547.500 275.400 549.300 287.400 ;
        RECT 561.600 275.400 563.400 287.400 ;
        RECT 529.950 269.850 532.050 271.950 ;
        RECT 532.950 271.050 535.050 273.150 ;
        RECT 530.100 268.050 531.900 269.850 ;
        RECT 523.950 266.550 528.450 267.450 ;
        RECT 523.950 265.950 526.050 266.550 ;
        RECT 521.850 263.700 525.600 264.750 ;
        RECT 506.400 262.800 510.000 263.700 ;
        RECT 508.200 255.600 510.000 262.800 ;
        RECT 515.400 260.700 523.200 262.050 ;
        RECT 515.400 255.600 517.200 260.700 ;
        RECT 521.400 255.600 523.200 260.700 ;
        RECT 524.400 261.600 525.600 263.700 ;
        RECT 533.400 263.700 534.600 271.050 ;
        RECT 535.950 269.850 538.050 271.950 ;
        RECT 542.100 270.150 543.900 271.950 ;
        RECT 547.950 270.150 549.150 275.400 ;
        RECT 550.950 273.150 552.750 274.950 ;
        RECT 561.000 274.350 563.400 275.400 ;
        RECT 569.400 281.400 571.200 287.400 ;
        RECT 569.400 274.500 570.600 281.400 ;
        RECT 575.700 275.400 577.500 287.400 ;
        RECT 586.800 281.400 588.600 287.400 ;
        RECT 550.950 271.050 553.050 273.150 ;
        RECT 557.100 270.150 558.900 271.950 ;
        RECT 536.100 268.050 537.900 269.850 ;
        RECT 541.950 268.050 544.050 270.150 ;
        RECT 544.950 266.850 547.050 268.950 ;
        RECT 547.950 268.050 550.050 270.150 ;
        RECT 556.950 268.050 559.050 270.150 ;
        RECT 545.100 265.050 546.900 266.850 ;
        RECT 548.850 264.750 550.050 268.050 ;
        RECT 561.000 267.150 562.050 274.350 ;
        RECT 569.400 273.600 575.100 274.500 ;
        RECT 573.150 272.700 575.100 273.600 ;
        RECT 563.100 270.150 564.900 271.950 ;
        RECT 569.100 270.150 570.900 271.950 ;
        RECT 562.950 268.050 565.050 270.150 ;
        RECT 568.950 268.050 571.050 270.150 ;
        RECT 559.950 265.050 562.050 267.150 ;
        RECT 548.850 263.700 552.600 264.750 ;
        RECT 533.400 262.800 537.000 263.700 ;
        RECT 524.400 255.600 526.200 261.600 ;
        RECT 535.200 255.600 537.000 262.800 ;
        RECT 542.400 260.700 550.200 262.050 ;
        RECT 542.400 255.600 544.200 260.700 ;
        RECT 548.400 255.600 550.200 260.700 ;
        RECT 551.400 261.600 552.600 263.700 ;
        RECT 551.400 255.600 553.200 261.600 ;
        RECT 561.000 258.600 562.050 265.050 ;
        RECT 573.150 264.300 574.050 272.700 ;
        RECT 576.000 270.150 577.200 275.400 ;
        RECT 587.400 273.150 588.600 281.400 ;
        RECT 593.400 276.600 595.200 287.400 ;
        RECT 599.400 286.500 607.200 287.400 ;
        RECT 599.400 276.600 601.200 286.500 ;
        RECT 593.400 275.700 601.200 276.600 ;
        RECT 602.400 274.500 604.200 285.600 ;
        RECT 605.400 275.400 607.200 286.500 ;
        RECT 618.600 275.400 620.400 287.400 ;
        RECT 629.400 281.400 631.200 287.400 ;
        RECT 646.800 281.400 648.600 287.400 ;
        RECT 600.150 273.600 604.200 274.500 ;
        RECT 618.600 274.350 621.000 275.400 ;
        RECT 574.950 268.050 577.200 270.150 ;
        RECT 583.950 269.850 586.050 271.950 ;
        RECT 586.950 271.050 589.050 273.150 ;
        RECT 584.100 268.050 585.900 269.850 ;
        RECT 573.150 263.400 575.100 264.300 ;
        RECT 570.000 262.500 575.100 263.400 ;
        RECT 570.000 258.600 571.200 262.500 ;
        RECT 576.000 261.600 577.200 268.050 ;
        RECT 587.400 263.700 588.600 271.050 ;
        RECT 589.950 269.850 592.050 271.950 ;
        RECT 593.250 270.150 595.050 271.950 ;
        RECT 600.150 270.150 601.050 273.600 ;
        RECT 605.100 270.150 606.900 271.950 ;
        RECT 617.100 270.150 618.900 271.950 ;
        RECT 590.100 268.050 591.900 269.850 ;
        RECT 592.950 268.050 595.050 270.150 ;
        RECT 595.950 266.850 598.050 268.950 ;
        RECT 596.250 265.050 598.050 266.850 ;
        RECT 598.950 268.050 601.050 270.150 ;
        RECT 585.000 262.800 588.600 263.700 ;
        RECT 560.400 255.600 562.200 258.600 ;
        RECT 569.400 255.600 571.200 258.600 ;
        RECT 575.700 255.600 577.500 261.600 ;
        RECT 585.000 255.600 586.800 262.800 ;
        RECT 598.950 261.600 600.000 268.050 ;
        RECT 601.950 266.850 604.050 268.950 ;
        RECT 604.950 268.050 607.050 270.150 ;
        RECT 616.950 268.050 619.050 270.150 ;
        RECT 619.950 267.150 621.000 274.350 ;
        RECT 629.400 273.150 630.600 281.400 ;
        RECT 647.400 273.150 648.600 281.400 ;
        RECT 658.500 275.400 660.300 287.400 ;
        RECT 671.400 281.400 673.200 287.400 ;
        RECT 623.100 270.150 624.900 271.950 ;
        RECT 622.950 268.050 625.050 270.150 ;
        RECT 625.950 269.850 628.050 271.950 ;
        RECT 628.950 271.050 631.050 273.150 ;
        RECT 626.100 268.050 627.900 269.850 ;
        RECT 601.950 265.050 603.750 266.850 ;
        RECT 619.950 265.050 622.050 267.150 ;
        RECT 598.200 255.600 600.000 261.600 ;
        RECT 619.950 258.600 621.000 265.050 ;
        RECT 629.400 263.700 630.600 271.050 ;
        RECT 631.950 269.850 634.050 271.950 ;
        RECT 643.950 269.850 646.050 271.950 ;
        RECT 646.950 271.050 649.050 273.150 ;
        RECT 632.100 268.050 633.900 269.850 ;
        RECT 644.100 268.050 645.900 269.850 ;
        RECT 647.400 263.700 648.600 271.050 ;
        RECT 649.950 269.850 652.050 271.950 ;
        RECT 653.100 270.150 654.900 271.950 ;
        RECT 658.950 270.150 660.150 275.400 ;
        RECT 661.950 273.150 663.750 274.950 ;
        RECT 667.950 273.450 670.050 274.050 ;
        RECT 661.950 271.050 664.050 273.150 ;
        RECT 665.550 272.550 670.050 273.450 ;
        RECT 650.100 268.050 651.900 269.850 ;
        RECT 652.950 268.050 655.050 270.150 ;
        RECT 655.950 266.850 658.050 268.950 ;
        RECT 658.950 268.050 661.050 270.150 ;
        RECT 656.100 265.050 657.900 266.850 ;
        RECT 659.850 264.750 661.050 268.050 ;
        RECT 661.950 267.450 664.050 268.050 ;
        RECT 665.550 267.450 666.450 272.550 ;
        RECT 667.950 271.950 670.050 272.550 ;
        RECT 671.400 268.950 672.600 281.400 ;
        RECT 679.800 275.400 681.600 287.400 ;
        RECT 682.800 276.300 684.600 287.400 ;
        RECT 688.800 276.300 690.600 287.400 ;
        RECT 694.800 281.400 696.600 287.400 ;
        RECT 682.800 275.400 690.600 276.300 ;
        RECT 680.400 270.150 681.300 275.400 ;
        RECT 691.950 274.950 694.050 277.050 ;
        RECT 661.950 266.550 666.450 267.450 ;
        RECT 668.100 267.150 669.900 268.950 ;
        RECT 661.950 265.950 664.050 266.550 ;
        RECT 667.950 265.050 670.050 267.150 ;
        RECT 670.950 266.850 673.050 268.950 ;
        RECT 679.950 268.050 682.050 270.150 ;
        RECT 659.850 263.700 663.600 264.750 ;
        RECT 629.400 262.800 633.000 263.700 ;
        RECT 619.800 255.600 621.600 258.600 ;
        RECT 631.200 255.600 633.000 262.800 ;
        RECT 645.000 262.800 648.600 263.700 ;
        RECT 645.000 255.600 646.800 262.800 ;
        RECT 653.400 260.700 661.200 262.050 ;
        RECT 653.400 255.600 655.200 260.700 ;
        RECT 659.400 255.600 661.200 260.700 ;
        RECT 662.400 261.600 663.600 263.700 ;
        RECT 662.400 255.600 664.200 261.600 ;
        RECT 671.400 258.600 672.600 266.850 ;
        RECT 680.400 261.600 681.300 268.050 ;
        RECT 682.950 266.850 685.050 268.950 ;
        RECT 686.100 267.150 687.900 268.950 ;
        RECT 683.100 265.050 684.900 266.850 ;
        RECT 685.950 265.050 688.050 267.150 ;
        RECT 688.950 266.850 691.050 268.950 ;
        RECT 689.100 265.050 690.900 266.850 ;
        RECT 692.550 262.050 693.450 274.950 ;
        RECT 695.400 268.950 696.600 281.400 ;
        RECT 706.500 275.400 708.300 287.400 ;
        RECT 721.500 275.400 723.300 287.400 ;
        RECT 733.800 281.400 735.600 287.400 ;
        RECT 734.700 281.100 735.600 281.400 ;
        RECT 739.800 281.400 741.600 287.400 ;
        RECT 749.400 281.400 751.200 287.400 ;
        RECT 739.800 281.100 741.300 281.400 ;
        RECT 734.700 280.200 741.300 281.100 ;
        RECT 749.700 281.100 751.200 281.400 ;
        RECT 755.400 281.400 757.200 287.400 ;
        RECT 755.400 281.100 756.300 281.400 ;
        RECT 749.700 280.200 756.300 281.100 ;
        RECT 727.950 279.450 730.050 280.050 ;
        RECT 727.950 278.550 732.450 279.450 ;
        RECT 727.950 277.950 730.050 278.550 ;
        RECT 701.100 270.150 702.900 271.950 ;
        RECT 706.950 270.150 708.150 275.400 ;
        RECT 709.950 273.150 711.750 274.950 ;
        RECT 709.950 271.050 712.050 273.150 ;
        RECT 716.100 270.150 717.900 271.950 ;
        RECT 721.950 270.150 723.150 275.400 ;
        RECT 724.950 273.150 726.750 274.950 ;
        RECT 724.950 271.050 727.050 273.150 ;
        RECT 694.950 266.850 697.050 268.950 ;
        RECT 698.100 267.150 699.900 268.950 ;
        RECT 700.950 268.050 703.050 270.150 ;
        RECT 680.400 259.950 685.800 261.600 ;
        RECT 691.950 259.950 694.050 262.050 ;
        RECT 671.400 255.600 673.200 258.600 ;
        RECT 684.000 255.600 685.800 259.950 ;
        RECT 695.400 258.600 696.600 266.850 ;
        RECT 697.950 265.050 700.050 267.150 ;
        RECT 703.950 266.850 706.050 268.950 ;
        RECT 706.950 268.050 709.050 270.150 ;
        RECT 715.950 268.050 718.050 270.150 ;
        RECT 704.100 265.050 705.900 266.850 ;
        RECT 707.850 264.750 709.050 268.050 ;
        RECT 718.950 266.850 721.050 268.950 ;
        RECT 721.950 268.050 724.050 270.150 ;
        RECT 719.100 265.050 720.900 266.850 ;
        RECT 722.850 264.750 724.050 268.050 ;
        RECT 707.850 263.700 711.600 264.750 ;
        RECT 722.850 263.700 726.600 264.750 ;
        RECT 694.800 255.600 696.600 258.600 ;
        RECT 701.400 260.700 709.200 262.050 ;
        RECT 701.400 255.600 703.200 260.700 ;
        RECT 707.400 255.600 709.200 260.700 ;
        RECT 710.400 261.600 711.600 263.700 ;
        RECT 710.400 255.600 712.200 261.600 ;
        RECT 716.400 260.700 724.200 262.050 ;
        RECT 716.400 255.600 718.200 260.700 ;
        RECT 722.400 255.600 724.200 260.700 ;
        RECT 725.400 261.600 726.600 263.700 ;
        RECT 725.400 255.600 727.200 261.600 ;
        RECT 731.550 261.450 732.450 278.550 ;
        RECT 734.700 271.950 735.600 280.200 ;
        RECT 740.100 276.150 741.900 277.950 ;
        RECT 749.100 276.150 750.900 277.950 ;
        RECT 736.950 273.150 738.750 274.950 ;
        RECT 739.950 274.050 742.050 276.150 ;
        RECT 743.100 273.150 744.900 274.950 ;
        RECT 746.100 273.150 747.900 274.950 ;
        RECT 748.950 274.050 751.050 276.150 ;
        RECT 752.250 273.150 754.050 274.950 ;
        RECT 733.950 269.850 736.050 271.950 ;
        RECT 736.950 271.050 739.050 273.150 ;
        RECT 742.950 271.050 745.050 273.150 ;
        RECT 745.950 271.050 748.050 273.150 ;
        RECT 751.950 271.050 754.050 273.150 ;
        RECT 755.400 271.950 756.300 280.200 ;
        RECT 754.950 269.850 757.050 271.950 ;
        RECT 734.700 265.650 735.600 269.850 ;
        RECT 755.400 265.650 756.300 269.850 ;
        RECT 734.700 264.000 738.900 265.650 ;
        RECT 733.950 261.450 736.050 262.050 ;
        RECT 731.550 260.550 736.050 261.450 ;
        RECT 733.950 259.950 736.050 260.550 ;
        RECT 737.100 255.600 738.900 264.000 ;
        RECT 752.100 264.000 756.300 265.650 ;
        RECT 752.100 255.600 753.900 264.000 ;
        RECT 7.800 245.400 9.600 251.400 ;
        RECT 13.800 248.400 15.600 251.400 ;
        RECT 7.950 240.150 9.000 245.400 ;
        RECT 13.800 244.200 14.700 248.400 ;
        RECT 11.250 243.300 14.700 244.200 ;
        RECT 24.000 244.200 25.800 251.400 ;
        RECT 34.800 245.400 36.600 251.400 ;
        RECT 40.800 248.400 42.600 251.400 ;
        RECT 24.000 243.300 27.600 244.200 ;
        RECT 11.250 242.400 13.050 243.300 ;
        RECT 7.950 238.050 10.050 240.150 ;
        RECT 8.700 231.450 10.050 238.050 ;
        RECT 11.400 234.150 12.300 242.400 ;
        RECT 16.950 239.850 19.050 241.950 ;
        RECT 13.950 236.850 16.050 238.950 ;
        RECT 17.100 238.050 18.900 239.850 ;
        RECT 23.100 237.150 24.900 238.950 ;
        RECT 14.100 235.050 15.900 236.850 ;
        RECT 22.950 235.050 25.050 237.150 ;
        RECT 26.400 235.950 27.600 243.300 ;
        RECT 31.950 238.950 34.050 241.050 ;
        RECT 34.950 240.150 36.000 245.400 ;
        RECT 40.800 244.200 41.700 248.400 ;
        RECT 52.800 245.400 54.600 251.400 ;
        RECT 38.250 243.300 41.700 244.200 ;
        RECT 53.400 243.300 54.600 245.400 ;
        RECT 55.800 246.300 57.600 251.400 ;
        RECT 61.800 246.300 63.600 251.400 ;
        RECT 67.800 248.400 69.600 251.400 ;
        RECT 55.800 244.950 63.600 246.300 ;
        RECT 38.250 242.400 40.050 243.300 ;
        RECT 29.100 237.150 30.900 238.950 ;
        RECT 11.400 234.000 13.200 234.150 ;
        RECT 11.400 232.800 18.600 234.000 ;
        RECT 25.950 233.850 28.050 235.950 ;
        RECT 28.950 235.050 31.050 237.150 ;
        RECT 11.400 232.350 13.200 232.800 ;
        RECT 17.400 231.600 18.600 232.800 ;
        RECT 8.700 230.100 11.100 231.450 ;
        RECT 9.300 219.600 11.100 230.100 ;
        RECT 16.800 219.600 18.600 231.600 ;
        RECT 26.400 225.600 27.600 233.850 ;
        RECT 32.550 232.050 33.450 238.950 ;
        RECT 34.950 238.050 37.050 240.150 ;
        RECT 31.950 229.950 34.050 232.050 ;
        RECT 35.700 231.450 37.050 238.050 ;
        RECT 38.400 234.150 39.300 242.400 ;
        RECT 53.400 242.250 57.150 243.300 ;
        RECT 43.950 239.850 46.050 241.950 ;
        RECT 40.950 236.850 43.050 238.950 ;
        RECT 44.100 238.050 45.900 239.850 ;
        RECT 55.950 238.950 57.150 242.250 ;
        RECT 59.100 240.150 60.900 241.950 ;
        RECT 68.400 240.150 69.600 248.400 ;
        RECT 80.100 243.000 81.900 251.400 ;
        RECT 93.000 244.200 94.800 251.400 ;
        RECT 105.000 244.200 106.800 251.400 ;
        RECT 116.400 248.400 118.200 251.400 ;
        RECT 93.000 243.300 96.600 244.200 ;
        RECT 105.000 243.300 108.600 244.200 ;
        RECT 55.950 236.850 58.050 238.950 ;
        RECT 58.950 238.050 61.050 240.150 ;
        RECT 61.950 236.850 64.050 238.950 ;
        RECT 67.950 238.050 70.050 240.150 ;
        RECT 70.950 239.850 73.050 241.950 ;
        RECT 80.100 241.350 84.300 243.000 ;
        RECT 71.100 238.050 72.900 239.850 ;
        RECT 41.100 235.050 42.900 236.850 ;
        RECT 38.400 234.000 40.200 234.150 ;
        RECT 38.400 232.800 45.600 234.000 ;
        RECT 52.950 233.850 55.050 235.950 ;
        RECT 38.400 232.350 40.200 232.800 ;
        RECT 44.400 231.600 45.600 232.800 ;
        RECT 53.250 232.050 55.050 233.850 ;
        RECT 56.850 231.600 58.050 236.850 ;
        RECT 62.100 235.050 63.900 236.850 ;
        RECT 35.700 230.100 38.100 231.450 ;
        RECT 25.800 219.600 27.600 225.600 ;
        RECT 36.300 219.600 38.100 230.100 ;
        RECT 43.800 219.600 45.600 231.600 ;
        RECT 56.700 219.600 58.500 231.600 ;
        RECT 68.400 225.600 69.600 238.050 ;
        RECT 83.400 237.150 84.300 241.350 ;
        RECT 92.100 237.150 93.900 238.950 ;
        RECT 73.950 233.850 76.050 235.950 ;
        RECT 79.950 233.850 82.050 235.950 ;
        RECT 82.950 235.050 85.050 237.150 ;
        RECT 91.950 235.050 94.050 237.150 ;
        RECT 95.400 235.950 96.600 243.300 ;
        RECT 98.100 237.150 99.900 238.950 ;
        RECT 104.100 237.150 105.900 238.950 ;
        RECT 74.100 232.050 75.900 233.850 ;
        RECT 76.950 230.850 79.050 232.950 ;
        RECT 80.250 232.050 82.050 233.850 ;
        RECT 77.100 229.050 78.900 230.850 ;
        RECT 83.400 226.800 84.300 235.050 ;
        RECT 94.950 233.850 97.050 235.950 ;
        RECT 97.950 235.050 100.050 237.150 ;
        RECT 103.950 235.050 106.050 237.150 ;
        RECT 107.400 235.950 108.600 243.300 ;
        RECT 117.000 241.950 118.050 248.400 ;
        RECT 125.400 246.000 127.200 251.400 ;
        RECT 131.400 250.500 139.200 251.400 ;
        RECT 131.400 246.000 133.200 250.500 ;
        RECT 125.400 245.100 133.200 246.000 ;
        RECT 134.400 245.400 136.200 249.600 ;
        RECT 137.400 245.400 139.200 250.500 ;
        RECT 146.400 248.400 148.200 251.400 ;
        RECT 160.800 248.400 162.600 251.400 ;
        RECT 169.800 248.400 171.600 251.400 ;
        RECT 181.800 248.400 183.600 251.400 ;
        RECT 134.700 243.900 135.600 245.400 ;
        RECT 131.400 242.850 135.600 243.900 ;
        RECT 115.950 239.850 118.050 241.950 ;
        RECT 128.100 240.150 129.900 241.950 ;
        RECT 110.100 237.150 111.900 238.950 ;
        RECT 106.950 233.850 109.050 235.950 ;
        RECT 109.950 235.050 112.050 237.150 ;
        RECT 112.950 236.850 115.050 238.950 ;
        RECT 113.100 235.050 114.900 236.850 ;
        RECT 77.700 225.900 84.300 226.800 ;
        RECT 77.700 225.600 79.200 225.900 ;
        RECT 67.800 219.600 69.600 225.600 ;
        RECT 77.400 219.600 79.200 225.600 ;
        RECT 83.400 225.600 84.300 225.900 ;
        RECT 95.400 225.600 96.600 233.850 ;
        RECT 107.400 225.600 108.600 233.850 ;
        RECT 117.000 232.650 118.050 239.850 ;
        RECT 118.950 236.850 121.050 238.950 ;
        RECT 124.950 236.850 127.050 238.950 ;
        RECT 127.950 238.050 130.050 240.150 ;
        RECT 131.400 238.950 132.600 242.850 ;
        RECT 147.000 241.950 148.050 248.400 ;
        RECT 133.500 240.150 135.300 241.950 ;
        RECT 130.950 236.850 133.050 238.950 ;
        RECT 133.950 238.050 136.050 240.150 ;
        RECT 145.950 239.850 148.050 241.950 ;
        RECT 161.400 240.150 162.600 248.400 ;
        RECT 136.950 236.850 139.050 238.950 ;
        RECT 142.950 236.850 145.050 238.950 ;
        RECT 119.100 235.050 120.900 236.850 ;
        RECT 125.100 235.050 126.900 236.850 ;
        RECT 117.000 231.600 119.400 232.650 ;
        RECT 131.400 231.600 132.600 236.850 ;
        RECT 136.950 235.050 138.750 236.850 ;
        RECT 143.100 235.050 144.900 236.850 ;
        RECT 147.000 232.650 148.050 239.850 ;
        RECT 148.950 236.850 151.050 238.950 ;
        RECT 160.950 238.050 163.050 240.150 ;
        RECT 163.950 239.850 166.050 241.950 ;
        RECT 170.400 240.150 171.600 248.400 ;
        RECT 175.950 244.950 178.050 247.050 ;
        RECT 164.100 238.050 165.900 239.850 ;
        RECT 169.950 238.050 172.050 240.150 ;
        RECT 172.950 239.850 175.050 241.950 ;
        RECT 173.100 238.050 174.900 239.850 ;
        RECT 149.100 235.050 150.900 236.850 ;
        RECT 147.000 231.600 149.400 232.650 ;
        RECT 83.400 219.600 85.200 225.600 ;
        RECT 94.800 219.600 96.600 225.600 ;
        RECT 106.800 219.600 108.600 225.600 ;
        RECT 117.600 219.600 119.400 231.600 ;
        RECT 129.900 219.600 133.200 231.600 ;
        RECT 147.600 219.600 149.400 231.600 ;
        RECT 161.400 225.600 162.600 238.050 ;
        RECT 170.400 225.600 171.600 238.050 ;
        RECT 172.950 234.450 175.050 235.050 ;
        RECT 176.550 234.450 177.450 244.950 ;
        RECT 181.950 241.950 183.000 248.400 ;
        RECT 193.200 244.200 195.000 251.400 ;
        RECT 191.400 243.300 195.000 244.200 ;
        RECT 210.000 245.400 211.800 251.400 ;
        RECT 181.950 239.850 184.050 241.950 ;
        RECT 178.950 236.850 181.050 238.950 ;
        RECT 179.100 235.050 180.900 236.850 ;
        RECT 172.950 233.550 177.450 234.450 ;
        RECT 172.950 232.950 175.050 233.550 ;
        RECT 181.950 232.650 183.000 239.850 ;
        RECT 184.950 236.850 187.050 238.950 ;
        RECT 188.100 237.150 189.900 238.950 ;
        RECT 185.100 235.050 186.900 236.850 ;
        RECT 187.950 235.050 190.050 237.150 ;
        RECT 191.400 235.950 192.600 243.300 ;
        RECT 206.250 240.150 208.050 241.950 ;
        RECT 194.100 237.150 195.900 238.950 ;
        RECT 190.950 233.850 193.050 235.950 ;
        RECT 193.950 235.050 196.050 237.150 ;
        RECT 202.950 236.850 205.050 238.950 ;
        RECT 205.950 238.050 208.050 240.150 ;
        RECT 210.000 238.950 211.050 245.400 ;
        RECT 221.400 243.900 223.200 251.400 ;
        RECT 228.900 246.900 230.700 251.400 ;
        RECT 228.900 245.400 232.050 246.900 ;
        RECT 227.100 243.900 228.900 244.500 ;
        RECT 221.400 242.700 228.900 243.900 ;
        RECT 208.950 236.850 211.050 238.950 ;
        RECT 211.950 240.150 213.750 241.950 ;
        RECT 211.950 238.050 214.050 240.150 ;
        RECT 214.950 236.850 217.050 238.950 ;
        RECT 220.950 236.850 223.050 238.950 ;
        RECT 203.100 235.050 204.900 236.850 ;
        RECT 160.800 219.600 162.600 225.600 ;
        RECT 169.800 219.600 171.600 225.600 ;
        RECT 180.600 231.600 183.000 232.650 ;
        RECT 180.600 219.600 182.400 231.600 ;
        RECT 191.400 225.600 192.600 233.850 ;
        RECT 208.950 233.400 209.850 236.850 ;
        RECT 214.950 235.050 216.750 236.850 ;
        RECT 221.100 235.050 222.900 236.850 ;
        RECT 205.800 232.500 209.850 233.400 ;
        RECT 191.400 219.600 193.200 225.600 ;
        RECT 202.800 220.500 204.600 231.600 ;
        RECT 205.800 221.400 207.600 232.500 ;
        RECT 208.800 230.400 216.600 231.300 ;
        RECT 208.800 220.500 210.600 230.400 ;
        RECT 202.800 219.600 210.600 220.500 ;
        RECT 214.800 219.600 216.600 230.400 ;
        RECT 224.550 225.600 225.600 242.700 ;
        RECT 231.000 238.950 232.050 245.400 ;
        RECT 241.200 244.200 243.000 251.400 ;
        RECT 250.800 245.400 252.600 251.400 ;
        RECT 239.400 243.300 243.000 244.200 ;
        RECT 251.400 243.300 252.600 245.400 ;
        RECT 253.800 246.300 255.600 251.400 ;
        RECT 259.800 246.300 261.600 251.400 ;
        RECT 253.800 244.950 261.600 246.300 ;
        RECT 268.800 245.400 270.600 251.400 ;
        RECT 269.400 243.300 270.600 245.400 ;
        RECT 271.800 246.300 273.600 251.400 ;
        RECT 277.800 246.300 279.600 251.400 ;
        RECT 285.300 246.900 287.100 251.400 ;
        RECT 271.800 244.950 279.600 246.300 ;
        RECT 283.950 245.400 287.100 246.900 ;
        RECT 227.100 237.150 228.900 238.950 ;
        RECT 226.950 235.050 229.050 237.150 ;
        RECT 229.950 236.850 232.050 238.950 ;
        RECT 236.100 237.150 237.900 238.950 ;
        RECT 231.000 231.600 232.050 236.850 ;
        RECT 235.950 235.050 238.050 237.150 ;
        RECT 239.400 235.950 240.600 243.300 ;
        RECT 251.400 242.250 255.150 243.300 ;
        RECT 269.400 242.250 273.150 243.300 ;
        RECT 253.950 238.950 255.150 242.250 ;
        RECT 257.100 240.150 258.900 241.950 ;
        RECT 242.100 237.150 243.900 238.950 ;
        RECT 238.950 233.850 241.050 235.950 ;
        RECT 241.950 235.050 244.050 237.150 ;
        RECT 253.950 236.850 256.050 238.950 ;
        RECT 256.950 238.050 259.050 240.150 ;
        RECT 271.950 238.950 273.150 242.250 ;
        RECT 275.100 240.150 276.900 241.950 ;
        RECT 259.950 236.850 262.050 238.950 ;
        RECT 271.950 236.850 274.050 238.950 ;
        RECT 274.950 238.050 277.050 240.150 ;
        RECT 283.950 238.950 285.000 245.400 ;
        RECT 287.100 243.900 288.900 244.500 ;
        RECT 292.800 243.900 294.600 251.400 ;
        RECT 304.200 245.400 306.000 251.400 ;
        RECT 319.500 245.400 321.300 251.400 ;
        RECT 325.800 248.400 327.600 251.400 ;
        RECT 287.100 242.700 294.600 243.900 ;
        RECT 277.950 236.850 280.050 238.950 ;
        RECT 283.950 236.850 286.050 238.950 ;
        RECT 287.100 237.150 288.900 238.950 ;
        RECT 250.950 233.850 253.050 235.950 ;
        RECT 224.400 219.600 226.200 225.600 ;
        RECT 231.000 219.600 232.800 231.600 ;
        RECT 239.400 225.600 240.600 233.850 ;
        RECT 251.250 232.050 253.050 233.850 ;
        RECT 254.850 231.600 256.050 236.850 ;
        RECT 260.100 235.050 261.900 236.850 ;
        RECT 268.950 233.850 271.050 235.950 ;
        RECT 269.250 232.050 271.050 233.850 ;
        RECT 272.850 231.600 274.050 236.850 ;
        RECT 278.100 235.050 279.900 236.850 ;
        RECT 283.950 231.600 285.000 236.850 ;
        RECT 286.950 235.050 289.050 237.150 ;
        RECT 239.400 219.600 241.200 225.600 ;
        RECT 254.700 219.600 256.500 231.600 ;
        RECT 272.700 219.600 274.500 231.600 ;
        RECT 283.200 219.600 285.000 231.600 ;
        RECT 290.400 225.600 291.450 242.700 ;
        RECT 302.250 240.150 304.050 241.950 ;
        RECT 292.950 236.850 295.050 238.950 ;
        RECT 298.950 236.850 301.050 238.950 ;
        RECT 301.950 238.050 304.050 240.150 ;
        RECT 304.950 238.950 306.000 245.400 ;
        RECT 307.950 240.150 309.750 241.950 ;
        RECT 304.950 236.850 307.050 238.950 ;
        RECT 307.950 238.050 310.050 240.150 ;
        RECT 319.800 238.950 321.000 245.400 ;
        RECT 325.800 244.500 327.000 248.400 ;
        RECT 321.900 243.600 327.000 244.500 ;
        RECT 329.400 243.900 331.200 251.400 ;
        RECT 336.900 246.900 338.700 251.400 ;
        RECT 336.900 245.400 340.050 246.900 ;
        RECT 346.500 245.400 348.300 251.400 ;
        RECT 352.800 248.400 354.600 251.400 ;
        RECT 335.100 243.900 336.900 244.500 ;
        RECT 321.900 242.700 323.850 243.600 ;
        RECT 329.400 242.700 336.900 243.900 ;
        RECT 310.950 236.850 313.050 238.950 ;
        RECT 319.800 236.850 322.050 238.950 ;
        RECT 293.100 235.050 294.900 236.850 ;
        RECT 299.250 235.050 301.050 236.850 ;
        RECT 306.150 233.400 307.050 236.850 ;
        RECT 311.100 235.050 312.900 236.850 ;
        RECT 306.150 232.500 310.200 233.400 ;
        RECT 299.400 230.400 307.200 231.300 ;
        RECT 289.800 219.600 291.600 225.600 ;
        RECT 299.400 219.600 301.200 230.400 ;
        RECT 305.400 220.500 307.200 230.400 ;
        RECT 308.400 221.400 310.200 232.500 ;
        RECT 319.800 231.600 321.000 236.850 ;
        RECT 322.950 234.300 323.850 242.700 ;
        RECT 325.950 236.850 328.050 238.950 ;
        RECT 328.950 236.850 331.050 238.950 ;
        RECT 326.100 235.050 327.900 236.850 ;
        RECT 329.100 235.050 330.900 236.850 ;
        RECT 321.900 233.400 323.850 234.300 ;
        RECT 321.900 232.500 327.600 233.400 ;
        RECT 311.400 220.500 313.200 231.600 ;
        RECT 305.400 219.600 313.200 220.500 ;
        RECT 319.500 219.600 321.300 231.600 ;
        RECT 326.400 225.600 327.600 232.500 ;
        RECT 332.550 225.600 333.600 242.700 ;
        RECT 339.000 238.950 340.050 245.400 ;
        RECT 335.100 237.150 336.900 238.950 ;
        RECT 334.950 235.050 337.050 237.150 ;
        RECT 337.950 236.850 340.050 238.950 ;
        RECT 339.000 231.600 340.050 236.850 ;
        RECT 346.800 238.950 348.000 245.400 ;
        RECT 352.800 244.500 354.000 248.400 ;
        RECT 358.800 245.400 360.600 251.400 ;
        RECT 348.900 243.600 354.000 244.500 ;
        RECT 348.900 242.700 350.850 243.600 ;
        RECT 346.800 236.850 349.050 238.950 ;
        RECT 346.800 231.600 348.000 236.850 ;
        RECT 349.950 234.300 350.850 242.700 ;
        RECT 359.400 238.950 360.600 245.400 ;
        RECT 365.400 243.900 367.200 251.400 ;
        RECT 372.900 246.900 374.700 251.400 ;
        RECT 372.900 245.400 376.050 246.900 ;
        RECT 371.100 243.900 372.900 244.500 ;
        RECT 365.400 242.700 372.900 243.900 ;
        RECT 362.100 240.150 363.900 241.950 ;
        RECT 352.950 236.850 355.050 238.950 ;
        RECT 358.950 236.850 361.050 238.950 ;
        RECT 361.950 238.050 364.050 240.150 ;
        RECT 364.950 236.850 367.050 238.950 ;
        RECT 353.100 235.050 354.900 236.850 ;
        RECT 348.900 233.400 350.850 234.300 ;
        RECT 348.900 232.500 354.600 233.400 ;
        RECT 325.800 219.600 327.600 225.600 ;
        RECT 332.400 219.600 334.200 225.600 ;
        RECT 339.000 219.600 340.800 231.600 ;
        RECT 346.500 219.600 348.300 231.600 ;
        RECT 353.400 225.600 354.600 232.500 ;
        RECT 359.400 231.600 360.600 236.850 ;
        RECT 365.100 235.050 366.900 236.850 ;
        RECT 352.800 219.600 354.600 225.600 ;
        RECT 358.800 219.600 360.600 231.600 ;
        RECT 368.550 225.600 369.600 242.700 ;
        RECT 375.000 238.950 376.050 245.400 ;
        RECT 383.400 243.900 385.200 251.400 ;
        RECT 390.900 246.900 392.700 251.400 ;
        RECT 390.900 245.400 394.050 246.900 ;
        RECT 389.100 243.900 390.900 244.500 ;
        RECT 383.400 242.700 390.900 243.900 ;
        RECT 371.100 237.150 372.900 238.950 ;
        RECT 370.950 235.050 373.050 237.150 ;
        RECT 373.950 236.850 376.050 238.950 ;
        RECT 382.950 236.850 385.050 238.950 ;
        RECT 375.000 231.600 376.050 236.850 ;
        RECT 383.100 235.050 384.900 236.850 ;
        RECT 368.400 219.600 370.200 225.600 ;
        RECT 375.000 219.600 376.800 231.600 ;
        RECT 386.550 225.600 387.600 242.700 ;
        RECT 393.000 238.950 394.050 245.400 ;
        RECT 403.200 244.200 405.000 251.400 ;
        RECT 412.800 245.400 414.600 251.400 ;
        RECT 401.400 243.300 405.000 244.200 ;
        RECT 413.400 243.300 414.600 245.400 ;
        RECT 415.800 246.300 417.600 251.400 ;
        RECT 421.800 246.300 423.600 251.400 ;
        RECT 415.800 244.950 423.600 246.300 ;
        RECT 430.200 244.200 432.000 251.400 ;
        RECT 439.800 245.400 441.600 251.400 ;
        RECT 428.400 243.300 432.000 244.200 ;
        RECT 440.400 243.300 441.600 245.400 ;
        RECT 442.800 246.300 444.600 251.400 ;
        RECT 448.800 246.300 450.600 251.400 ;
        RECT 442.800 244.950 450.600 246.300 ;
        RECT 389.100 237.150 390.900 238.950 ;
        RECT 388.950 235.050 391.050 237.150 ;
        RECT 391.950 236.850 394.050 238.950 ;
        RECT 398.100 237.150 399.900 238.950 ;
        RECT 393.000 231.600 394.050 236.850 ;
        RECT 397.950 235.050 400.050 237.150 ;
        RECT 401.400 235.950 402.600 243.300 ;
        RECT 413.400 242.250 417.150 243.300 ;
        RECT 415.950 238.950 417.150 242.250 ;
        RECT 419.100 240.150 420.900 241.950 ;
        RECT 404.100 237.150 405.900 238.950 ;
        RECT 400.950 233.850 403.050 235.950 ;
        RECT 403.950 235.050 406.050 237.150 ;
        RECT 415.950 236.850 418.050 238.950 ;
        RECT 418.950 238.050 421.050 240.150 ;
        RECT 421.950 236.850 424.050 238.950 ;
        RECT 425.100 237.150 426.900 238.950 ;
        RECT 412.950 233.850 415.050 235.950 ;
        RECT 386.400 219.600 388.200 225.600 ;
        RECT 393.000 219.600 394.800 231.600 ;
        RECT 401.400 225.600 402.600 233.850 ;
        RECT 413.250 232.050 415.050 233.850 ;
        RECT 416.850 231.600 418.050 236.850 ;
        RECT 422.100 235.050 423.900 236.850 ;
        RECT 424.950 235.050 427.050 237.150 ;
        RECT 428.400 235.950 429.600 243.300 ;
        RECT 440.400 242.250 444.150 243.300 ;
        RECT 461.100 243.000 462.900 251.400 ;
        RECT 475.200 244.200 477.000 251.400 ;
        RECT 484.800 245.400 486.600 251.400 ;
        RECT 442.950 238.950 444.150 242.250 ;
        RECT 446.100 240.150 447.900 241.950 ;
        RECT 458.700 241.350 462.900 243.000 ;
        RECT 473.400 243.300 477.000 244.200 ;
        RECT 485.400 243.300 486.600 245.400 ;
        RECT 487.800 246.300 489.600 251.400 ;
        RECT 493.800 246.300 495.600 251.400 ;
        RECT 487.800 244.950 495.600 246.300 ;
        RECT 501.000 244.200 502.800 251.400 ;
        RECT 512.400 248.400 514.200 251.400 ;
        RECT 493.950 243.450 496.050 244.050 ;
        RECT 431.100 237.150 432.900 238.950 ;
        RECT 427.950 233.850 430.050 235.950 ;
        RECT 430.950 235.050 433.050 237.150 ;
        RECT 442.950 236.850 445.050 238.950 ;
        RECT 445.950 238.050 448.050 240.150 ;
        RECT 448.950 236.850 451.050 238.950 ;
        RECT 458.700 237.150 459.600 241.350 ;
        RECT 470.100 237.150 471.900 238.950 ;
        RECT 439.950 233.850 442.050 235.950 ;
        RECT 401.400 219.600 403.200 225.600 ;
        RECT 416.700 219.600 418.500 231.600 ;
        RECT 428.400 225.600 429.600 233.850 ;
        RECT 440.250 232.050 442.050 233.850 ;
        RECT 443.850 231.600 445.050 236.850 ;
        RECT 449.100 235.050 450.900 236.850 ;
        RECT 457.950 235.050 460.050 237.150 ;
        RECT 428.400 219.600 430.200 225.600 ;
        RECT 443.700 219.600 445.500 231.600 ;
        RECT 458.700 226.800 459.600 235.050 ;
        RECT 460.950 233.850 463.050 235.950 ;
        RECT 466.950 233.850 469.050 235.950 ;
        RECT 469.950 235.050 472.050 237.150 ;
        RECT 473.400 235.950 474.600 243.300 ;
        RECT 485.400 242.250 489.150 243.300 ;
        RECT 487.950 238.950 489.150 242.250 ;
        RECT 493.950 242.550 498.450 243.450 ;
        RECT 501.000 243.300 504.600 244.200 ;
        RECT 493.950 241.950 496.050 242.550 ;
        RECT 491.100 240.150 492.900 241.950 ;
        RECT 476.100 237.150 477.900 238.950 ;
        RECT 472.950 233.850 475.050 235.950 ;
        RECT 475.950 235.050 478.050 237.150 ;
        RECT 487.950 236.850 490.050 238.950 ;
        RECT 490.950 238.050 493.050 240.150 ;
        RECT 493.950 236.850 496.050 238.950 ;
        RECT 484.950 233.850 487.050 235.950 ;
        RECT 460.950 232.050 462.750 233.850 ;
        RECT 463.950 230.850 466.050 232.950 ;
        RECT 467.100 232.050 468.900 233.850 ;
        RECT 464.100 229.050 465.900 230.850 ;
        RECT 458.700 225.900 465.300 226.800 ;
        RECT 458.700 225.600 459.600 225.900 ;
        RECT 457.800 219.600 459.600 225.600 ;
        RECT 463.800 225.600 465.300 225.900 ;
        RECT 473.400 225.600 474.600 233.850 ;
        RECT 485.250 232.050 487.050 233.850 ;
        RECT 488.850 231.600 490.050 236.850 ;
        RECT 494.100 235.050 495.900 236.850 ;
        RECT 463.800 219.600 465.600 225.600 ;
        RECT 473.400 219.600 475.200 225.600 ;
        RECT 488.700 219.600 490.500 231.600 ;
        RECT 497.550 231.450 498.450 242.550 ;
        RECT 500.100 237.150 501.900 238.950 ;
        RECT 499.950 235.050 502.050 237.150 ;
        RECT 503.400 235.950 504.600 243.300 ;
        RECT 508.950 239.850 511.050 241.950 ;
        RECT 512.400 240.150 513.600 248.400 ;
        RECT 523.200 245.400 525.000 251.400 ;
        RECT 521.250 240.150 523.050 241.950 ;
        RECT 506.100 237.150 507.900 238.950 ;
        RECT 509.100 238.050 510.900 239.850 ;
        RECT 511.950 238.050 514.050 240.150 ;
        RECT 502.950 233.850 505.050 235.950 ;
        RECT 505.950 235.050 508.050 237.150 ;
        RECT 499.950 231.450 502.050 232.050 ;
        RECT 497.550 230.550 502.050 231.450 ;
        RECT 499.950 229.950 502.050 230.550 ;
        RECT 503.400 225.600 504.600 233.850 ;
        RECT 502.800 219.600 504.600 225.600 ;
        RECT 512.400 225.600 513.600 238.050 ;
        RECT 517.950 236.850 520.050 238.950 ;
        RECT 520.950 238.050 523.050 240.150 ;
        RECT 523.950 238.950 525.000 245.400 ;
        RECT 539.400 246.300 541.200 251.400 ;
        RECT 545.400 246.300 547.200 251.400 ;
        RECT 539.400 244.950 547.200 246.300 ;
        RECT 548.400 245.400 550.200 251.400 ;
        RECT 548.400 243.300 549.600 245.400 ;
        RECT 545.850 242.250 549.600 243.300 ;
        RECT 560.100 243.000 561.900 251.400 ;
        RECT 576.000 244.200 577.800 251.400 ;
        RECT 589.800 248.400 591.600 251.400 ;
        RECT 576.000 243.300 579.600 244.200 ;
        RECT 526.950 240.150 528.750 241.950 ;
        RECT 542.100 240.150 543.900 241.950 ;
        RECT 523.950 236.850 526.050 238.950 ;
        RECT 526.950 238.050 529.050 240.150 ;
        RECT 529.950 236.850 532.050 238.950 ;
        RECT 538.950 236.850 541.050 238.950 ;
        RECT 541.950 238.050 544.050 240.150 ;
        RECT 545.850 238.950 547.050 242.250 ;
        RECT 560.100 241.350 564.300 243.000 ;
        RECT 556.950 240.450 559.050 241.050 ;
        RECT 544.950 236.850 547.050 238.950 ;
        RECT 551.550 239.550 559.050 240.450 ;
        RECT 518.250 235.050 520.050 236.850 ;
        RECT 525.150 233.400 526.050 236.850 ;
        RECT 530.100 235.050 531.900 236.850 ;
        RECT 539.100 235.050 540.900 236.850 ;
        RECT 525.150 232.500 529.200 233.400 ;
        RECT 518.400 230.400 526.200 231.300 ;
        RECT 512.400 219.600 514.200 225.600 ;
        RECT 518.400 219.600 520.200 230.400 ;
        RECT 524.400 220.500 526.200 230.400 ;
        RECT 527.400 221.400 529.200 232.500 ;
        RECT 544.950 231.600 546.150 236.850 ;
        RECT 547.950 233.850 550.050 235.950 ;
        RECT 547.950 232.050 549.750 233.850 ;
        RECT 551.550 232.050 552.450 239.550 ;
        RECT 556.950 238.950 559.050 239.550 ;
        RECT 563.400 237.150 564.300 241.350 ;
        RECT 565.950 240.450 568.050 241.050 ;
        RECT 565.950 239.550 573.450 240.450 ;
        RECT 565.950 238.950 568.050 239.550 ;
        RECT 553.950 233.850 556.050 235.950 ;
        RECT 559.950 233.850 562.050 235.950 ;
        RECT 562.950 235.050 565.050 237.150 ;
        RECT 568.950 235.950 571.050 238.050 ;
        RECT 554.100 232.050 555.900 233.850 ;
        RECT 530.400 220.500 532.200 231.600 ;
        RECT 524.400 219.600 532.200 220.500 ;
        RECT 544.500 219.600 546.300 231.600 ;
        RECT 550.950 229.950 553.050 232.050 ;
        RECT 556.950 230.850 559.050 232.950 ;
        RECT 560.250 232.050 562.050 233.850 ;
        RECT 557.100 229.050 558.900 230.850 ;
        RECT 563.400 226.800 564.300 235.050 ;
        RECT 557.700 225.900 564.300 226.800 ;
        RECT 569.550 226.050 570.450 235.950 ;
        RECT 572.550 231.450 573.450 239.550 ;
        RECT 575.100 237.150 576.900 238.950 ;
        RECT 574.950 235.050 577.050 237.150 ;
        RECT 578.400 235.950 579.600 243.300 ;
        RECT 580.950 243.450 583.050 244.050 ;
        RECT 580.950 242.550 585.450 243.450 ;
        RECT 580.950 241.950 583.050 242.550 ;
        RECT 581.100 237.150 582.900 238.950 ;
        RECT 584.550 238.050 585.450 242.550 ;
        RECT 589.950 241.950 591.000 248.400 ;
        RECT 603.000 244.200 604.800 251.400 ;
        RECT 614.400 248.400 616.200 251.400 ;
        RECT 615.300 244.200 616.200 248.400 ;
        RECT 620.400 245.400 622.200 251.400 ;
        RECT 636.000 247.050 637.800 251.400 ;
        RECT 632.400 245.400 637.800 247.050 ;
        RECT 603.000 243.300 606.600 244.200 ;
        RECT 615.300 243.300 618.750 244.200 ;
        RECT 589.950 239.850 592.050 241.950 ;
        RECT 577.950 233.850 580.050 235.950 ;
        RECT 580.950 235.050 583.050 237.150 ;
        RECT 583.950 235.950 586.050 238.050 ;
        RECT 586.950 236.850 589.050 238.950 ;
        RECT 587.100 235.050 588.900 236.850 ;
        RECT 574.950 231.450 577.050 232.050 ;
        RECT 572.550 230.550 577.050 231.450 ;
        RECT 574.950 229.950 577.050 230.550 ;
        RECT 557.700 225.600 559.200 225.900 ;
        RECT 557.400 219.600 559.200 225.600 ;
        RECT 563.400 225.600 564.300 225.900 ;
        RECT 563.400 219.600 565.200 225.600 ;
        RECT 568.950 223.950 571.050 226.050 ;
        RECT 578.400 225.600 579.600 233.850 ;
        RECT 589.950 232.650 591.000 239.850 ;
        RECT 592.950 236.850 595.050 238.950 ;
        RECT 602.100 237.150 603.900 238.950 ;
        RECT 593.100 235.050 594.900 236.850 ;
        RECT 601.950 235.050 604.050 237.150 ;
        RECT 605.400 235.950 606.600 243.300 ;
        RECT 616.950 242.400 618.750 243.300 ;
        RECT 610.950 239.850 613.050 241.950 ;
        RECT 608.100 237.150 609.900 238.950 ;
        RECT 611.100 238.050 612.900 239.850 ;
        RECT 604.950 233.850 607.050 235.950 ;
        RECT 607.950 235.050 610.050 237.150 ;
        RECT 613.950 236.850 616.050 238.950 ;
        RECT 614.100 235.050 615.900 236.850 ;
        RECT 617.700 234.150 618.600 242.400 ;
        RECT 621.000 240.150 622.050 245.400 ;
        RECT 616.800 234.000 618.600 234.150 ;
        RECT 577.800 219.600 579.600 225.600 ;
        RECT 588.600 231.600 591.000 232.650 ;
        RECT 588.600 219.600 590.400 231.600 ;
        RECT 605.400 225.600 606.600 233.850 ;
        RECT 604.800 219.600 606.600 225.600 ;
        RECT 611.400 232.800 618.600 234.000 ;
        RECT 611.400 231.600 612.600 232.800 ;
        RECT 616.800 232.350 618.600 232.800 ;
        RECT 619.950 238.050 622.050 240.150 ;
        RECT 632.400 238.950 633.300 245.400 ;
        RECT 648.000 244.200 649.800 251.400 ;
        RECT 648.000 243.300 651.600 244.200 ;
        RECT 635.100 240.150 636.900 241.950 ;
        RECT 611.400 219.600 613.200 231.600 ;
        RECT 619.950 231.450 621.300 238.050 ;
        RECT 631.950 236.850 634.050 238.950 ;
        RECT 634.950 238.050 637.050 240.150 ;
        RECT 637.950 239.850 640.050 241.950 ;
        RECT 641.100 240.150 642.900 241.950 ;
        RECT 638.100 238.050 639.900 239.850 ;
        RECT 640.950 238.050 643.050 240.150 ;
        RECT 647.100 237.150 648.900 238.950 ;
        RECT 632.400 231.600 633.300 236.850 ;
        RECT 646.950 235.050 649.050 237.150 ;
        RECT 650.400 235.950 651.600 243.300 ;
        RECT 656.400 243.900 658.200 251.400 ;
        RECT 663.900 246.900 665.700 251.400 ;
        RECT 663.900 245.400 667.050 246.900 ;
        RECT 676.200 245.400 678.000 251.400 ;
        RECT 691.800 245.400 693.600 251.400 ;
        RECT 662.100 243.900 663.900 244.500 ;
        RECT 656.400 242.700 663.900 243.900 ;
        RECT 653.100 237.150 654.900 238.950 ;
        RECT 649.950 233.850 652.050 235.950 ;
        RECT 652.950 235.050 655.050 237.150 ;
        RECT 655.950 236.850 658.050 238.950 ;
        RECT 656.100 235.050 657.900 236.850 ;
        RECT 618.900 230.100 621.300 231.450 ;
        RECT 618.900 219.600 620.700 230.100 ;
        RECT 631.800 219.600 633.600 231.600 ;
        RECT 634.800 230.700 642.600 231.600 ;
        RECT 634.800 219.600 636.600 230.700 ;
        RECT 640.800 219.600 642.600 230.700 ;
        RECT 650.400 225.600 651.600 233.850 ;
        RECT 659.550 225.600 660.600 242.700 ;
        RECT 666.000 238.950 667.050 245.400 ;
        RECT 674.250 240.150 676.050 241.950 ;
        RECT 662.100 237.150 663.900 238.950 ;
        RECT 661.950 235.050 664.050 237.150 ;
        RECT 664.950 236.850 667.050 238.950 ;
        RECT 670.950 236.850 673.050 238.950 ;
        RECT 673.950 238.050 676.050 240.150 ;
        RECT 676.950 238.950 678.000 245.400 ;
        RECT 682.950 243.450 685.050 244.050 ;
        RECT 682.950 242.550 690.450 243.450 ;
        RECT 682.950 241.950 685.050 242.550 ;
        RECT 679.950 240.150 681.750 241.950 ;
        RECT 676.950 236.850 679.050 238.950 ;
        RECT 679.950 238.050 682.050 240.150 ;
        RECT 682.950 236.850 685.050 238.950 ;
        RECT 666.000 231.600 667.050 236.850 ;
        RECT 671.250 235.050 673.050 236.850 ;
        RECT 678.150 233.400 679.050 236.850 ;
        RECT 683.100 235.050 684.900 236.850 ;
        RECT 678.150 232.500 682.200 233.400 ;
        RECT 649.800 219.600 651.600 225.600 ;
        RECT 659.400 219.600 661.200 225.600 ;
        RECT 666.000 219.600 667.800 231.600 ;
        RECT 671.400 230.400 679.200 231.300 ;
        RECT 671.400 219.600 673.200 230.400 ;
        RECT 677.400 220.500 679.200 230.400 ;
        RECT 680.400 221.400 682.200 232.500 ;
        RECT 683.400 220.500 685.200 231.600 ;
        RECT 689.550 228.450 690.450 242.550 ;
        RECT 692.400 243.300 693.600 245.400 ;
        RECT 694.800 246.300 696.600 251.400 ;
        RECT 700.800 246.300 702.600 251.400 ;
        RECT 694.800 244.950 702.600 246.300 ;
        RECT 704.400 246.300 706.200 251.400 ;
        RECT 710.400 246.300 712.200 251.400 ;
        RECT 704.400 244.950 712.200 246.300 ;
        RECT 713.400 245.400 715.200 251.400 ;
        RECT 713.400 243.300 714.600 245.400 ;
        RECT 692.400 242.250 696.150 243.300 ;
        RECT 694.950 238.950 696.150 242.250 ;
        RECT 710.850 242.250 714.600 243.300 ;
        RECT 725.100 243.000 726.900 251.400 ;
        RECT 743.100 243.000 744.900 251.400 ;
        RECT 761.100 243.000 762.900 251.400 ;
        RECT 698.100 240.150 699.900 241.950 ;
        RECT 707.100 240.150 708.900 241.950 ;
        RECT 694.950 236.850 697.050 238.950 ;
        RECT 697.950 238.050 700.050 240.150 ;
        RECT 700.950 236.850 703.050 238.950 ;
        RECT 703.950 236.850 706.050 238.950 ;
        RECT 706.950 238.050 709.050 240.150 ;
        RECT 710.850 238.950 712.050 242.250 ;
        RECT 725.100 241.350 729.300 243.000 ;
        RECT 743.100 241.350 747.300 243.000 ;
        RECT 721.950 240.450 724.050 241.050 ;
        RECT 709.950 236.850 712.050 238.950 ;
        RECT 716.550 239.550 724.050 240.450 ;
        RECT 691.950 233.850 694.050 235.950 ;
        RECT 692.250 232.050 694.050 233.850 ;
        RECT 695.850 231.600 697.050 236.850 ;
        RECT 701.100 235.050 702.900 236.850 ;
        RECT 704.100 235.050 705.900 236.850 ;
        RECT 709.950 231.600 711.150 236.850 ;
        RECT 712.950 233.850 715.050 235.950 ;
        RECT 712.950 232.050 714.750 233.850 ;
        RECT 716.550 232.050 717.450 239.550 ;
        RECT 721.950 238.950 724.050 239.550 ;
        RECT 728.400 237.150 729.300 241.350 ;
        RECT 733.950 240.450 736.050 241.050 ;
        RECT 739.950 240.450 742.050 241.050 ;
        RECT 733.950 239.550 742.050 240.450 ;
        RECT 733.950 238.950 736.050 239.550 ;
        RECT 739.950 238.950 742.050 239.550 ;
        RECT 746.400 237.150 747.300 241.350 ;
        RECT 758.700 241.350 762.900 243.000 ;
        RECT 748.950 238.950 751.050 241.050 ;
        RECT 718.950 233.850 721.050 235.950 ;
        RECT 724.950 233.850 727.050 235.950 ;
        RECT 727.950 235.050 730.050 237.150 ;
        RECT 719.100 232.050 720.900 233.850 ;
        RECT 691.950 228.450 694.050 229.050 ;
        RECT 689.550 227.550 694.050 228.450 ;
        RECT 691.950 226.950 694.050 227.550 ;
        RECT 677.400 219.600 685.200 220.500 ;
        RECT 695.700 219.600 697.500 231.600 ;
        RECT 709.500 219.600 711.300 231.600 ;
        RECT 715.950 229.950 718.050 232.050 ;
        RECT 721.950 230.850 724.050 232.950 ;
        RECT 725.250 232.050 727.050 233.850 ;
        RECT 722.100 229.050 723.900 230.850 ;
        RECT 728.400 226.800 729.300 235.050 ;
        RECT 736.950 233.850 739.050 235.950 ;
        RECT 742.950 233.850 745.050 235.950 ;
        RECT 745.950 235.050 748.050 237.150 ;
        RECT 737.100 232.050 738.900 233.850 ;
        RECT 730.950 229.950 733.050 232.050 ;
        RECT 739.950 230.850 742.050 232.950 ;
        RECT 743.250 232.050 745.050 233.850 ;
        RECT 731.550 228.450 732.450 229.950 ;
        RECT 740.100 229.050 741.900 230.850 ;
        RECT 733.950 228.450 736.050 229.050 ;
        RECT 731.550 227.550 736.050 228.450 ;
        RECT 733.950 226.950 736.050 227.550 ;
        RECT 746.400 226.800 747.300 235.050 ;
        RECT 749.550 229.050 750.450 238.950 ;
        RECT 758.700 237.150 759.600 241.350 ;
        RECT 757.950 235.050 760.050 237.150 ;
        RECT 748.950 226.950 751.050 229.050 ;
        RECT 722.700 225.900 729.300 226.800 ;
        RECT 722.700 225.600 724.200 225.900 ;
        RECT 722.400 219.600 724.200 225.600 ;
        RECT 728.400 225.600 729.300 225.900 ;
        RECT 740.700 225.900 747.300 226.800 ;
        RECT 740.700 225.600 742.200 225.900 ;
        RECT 728.400 219.600 730.200 225.600 ;
        RECT 740.400 219.600 742.200 225.600 ;
        RECT 746.400 225.600 747.300 225.900 ;
        RECT 758.700 226.800 759.600 235.050 ;
        RECT 760.950 233.850 763.050 235.950 ;
        RECT 766.950 233.850 769.050 235.950 ;
        RECT 760.950 232.050 762.750 233.850 ;
        RECT 763.950 230.850 766.050 232.950 ;
        RECT 767.100 232.050 768.900 233.850 ;
        RECT 764.100 229.050 765.900 230.850 ;
        RECT 758.700 225.900 765.300 226.800 ;
        RECT 758.700 225.600 759.600 225.900 ;
        RECT 746.400 219.600 748.200 225.600 ;
        RECT 757.800 219.600 759.600 225.600 ;
        RECT 763.800 225.600 765.300 225.900 ;
        RECT 763.800 219.600 765.600 225.600 ;
        RECT 1.950 205.950 4.050 208.050 ;
        RECT 2.550 195.450 3.450 205.950 ;
        RECT 8.700 203.400 10.500 215.400 ;
        RECT 19.800 209.400 21.600 215.400 ;
        RECT 5.250 201.150 7.050 202.950 ;
        RECT 4.950 199.050 7.050 201.150 ;
        RECT 8.850 198.150 10.050 203.400 ;
        RECT 14.100 198.150 15.900 199.950 ;
        RECT 7.950 196.050 10.050 198.150 ;
        RECT 4.950 195.450 7.050 196.050 ;
        RECT 2.550 194.550 7.050 195.450 ;
        RECT 4.950 193.950 7.050 194.550 ;
        RECT 7.950 192.750 9.150 196.050 ;
        RECT 10.950 194.850 13.050 196.950 ;
        RECT 13.950 196.050 16.050 198.150 ;
        RECT 20.400 196.950 21.600 209.400 ;
        RECT 31.500 203.400 33.300 215.400 ;
        RECT 44.400 209.400 46.200 215.400 ;
        RECT 44.700 209.100 46.200 209.400 ;
        RECT 50.400 209.400 52.200 215.400 ;
        RECT 61.800 209.400 63.600 215.400 ;
        RECT 50.400 209.100 51.300 209.400 ;
        RECT 44.700 208.200 51.300 209.100 ;
        RECT 44.100 204.150 45.900 205.950 ;
        RECT 26.100 198.150 27.900 199.950 ;
        RECT 31.950 198.150 33.150 203.400 ;
        RECT 34.950 201.150 36.750 202.950 ;
        RECT 41.100 201.150 42.900 202.950 ;
        RECT 43.950 202.050 46.050 204.150 ;
        RECT 47.250 201.150 49.050 202.950 ;
        RECT 34.950 199.050 37.050 201.150 ;
        RECT 40.950 199.050 43.050 201.150 ;
        RECT 46.950 199.050 49.050 201.150 ;
        RECT 50.400 199.950 51.300 208.200 ;
        RECT 19.950 194.850 22.050 196.950 ;
        RECT 23.100 195.150 24.900 196.950 ;
        RECT 25.950 196.050 28.050 198.150 ;
        RECT 11.100 193.050 12.900 194.850 ;
        RECT 5.400 191.700 9.150 192.750 ;
        RECT 5.400 189.600 6.600 191.700 ;
        RECT 4.800 183.600 6.600 189.600 ;
        RECT 7.800 188.700 15.600 190.050 ;
        RECT 7.800 183.600 9.600 188.700 ;
        RECT 13.800 183.600 15.600 188.700 ;
        RECT 20.400 186.600 21.600 194.850 ;
        RECT 22.950 193.050 25.050 195.150 ;
        RECT 28.950 194.850 31.050 196.950 ;
        RECT 31.950 196.050 34.050 198.150 ;
        RECT 49.950 197.850 52.050 199.950 ;
        RECT 29.100 193.050 30.900 194.850 ;
        RECT 32.850 192.750 34.050 196.050 ;
        RECT 50.400 193.650 51.300 197.850 ;
        RECT 62.400 196.950 63.600 209.400 ;
        RECT 70.800 203.400 72.600 215.400 ;
        RECT 73.800 204.300 75.600 215.400 ;
        RECT 79.800 204.300 81.600 215.400 ;
        RECT 73.800 203.400 81.600 204.300 ;
        RECT 86.400 209.400 88.200 215.400 ;
        RECT 71.400 198.150 72.300 203.400 ;
        RECT 86.400 201.150 87.600 209.400 ;
        RECT 104.700 203.400 106.500 215.400 ;
        RECT 120.600 203.400 122.400 215.400 ;
        RECT 130.800 209.400 132.600 215.400 ;
        RECT 101.250 201.150 103.050 202.950 ;
        RECT 61.950 194.850 64.050 196.950 ;
        RECT 65.100 195.150 66.900 196.950 ;
        RECT 70.950 196.050 73.050 198.150 ;
        RECT 82.950 197.850 85.050 199.950 ;
        RECT 85.950 199.050 88.050 201.150 ;
        RECT 32.850 191.700 36.600 192.750 ;
        RECT 19.800 183.600 21.600 186.600 ;
        RECT 26.400 188.700 34.200 190.050 ;
        RECT 26.400 183.600 28.200 188.700 ;
        RECT 32.400 183.600 34.200 188.700 ;
        RECT 35.400 189.600 36.600 191.700 ;
        RECT 47.100 192.000 51.300 193.650 ;
        RECT 35.400 183.600 37.200 189.600 ;
        RECT 47.100 183.600 48.900 192.000 ;
        RECT 62.400 186.600 63.600 194.850 ;
        RECT 64.950 193.050 67.050 195.150 ;
        RECT 71.400 189.600 72.300 196.050 ;
        RECT 73.950 194.850 76.050 196.950 ;
        RECT 77.100 195.150 78.900 196.950 ;
        RECT 74.100 193.050 75.900 194.850 ;
        RECT 76.950 193.050 79.050 195.150 ;
        RECT 79.950 194.850 82.050 196.950 ;
        RECT 83.100 196.050 84.900 197.850 ;
        RECT 80.100 193.050 81.900 194.850 ;
        RECT 86.400 191.700 87.600 199.050 ;
        RECT 88.950 197.850 91.050 199.950 ;
        RECT 100.950 199.050 103.050 201.150 ;
        RECT 104.850 198.150 106.050 203.400 ;
        RECT 120.600 202.350 123.000 203.400 ;
        RECT 110.100 198.150 111.900 199.950 ;
        RECT 119.100 198.150 120.900 199.950 ;
        RECT 89.100 196.050 90.900 197.850 ;
        RECT 103.950 196.050 106.050 198.150 ;
        RECT 103.950 192.750 105.150 196.050 ;
        RECT 106.950 194.850 109.050 196.950 ;
        RECT 109.950 196.050 112.050 198.150 ;
        RECT 118.950 196.050 121.050 198.150 ;
        RECT 121.950 195.150 123.000 202.350 ;
        RECT 125.100 198.150 126.900 199.950 ;
        RECT 124.950 196.050 127.050 198.150 ;
        RECT 131.400 196.950 132.600 209.400 ;
        RECT 139.200 203.400 141.000 215.400 ;
        RECT 145.800 209.400 147.600 215.400 ;
        RECT 133.950 201.450 136.050 202.050 ;
        RECT 133.950 200.550 138.450 201.450 ;
        RECT 133.950 199.950 136.050 200.550 ;
        RECT 107.100 193.050 108.900 194.850 ;
        RECT 121.950 193.050 124.050 195.150 ;
        RECT 130.950 194.850 133.050 196.950 ;
        RECT 134.100 195.150 135.900 196.950 ;
        RECT 101.400 191.700 105.150 192.750 ;
        RECT 86.400 190.800 90.000 191.700 ;
        RECT 71.400 187.950 76.800 189.600 ;
        RECT 61.800 183.600 63.600 186.600 ;
        RECT 75.000 183.600 76.800 187.950 ;
        RECT 88.200 183.600 90.000 190.800 ;
        RECT 101.400 189.600 102.600 191.700 ;
        RECT 100.800 183.600 102.600 189.600 ;
        RECT 103.800 188.700 111.600 190.050 ;
        RECT 103.800 183.600 105.600 188.700 ;
        RECT 109.800 183.600 111.600 188.700 ;
        RECT 121.950 186.600 123.000 193.050 ;
        RECT 131.400 186.600 132.600 194.850 ;
        RECT 133.950 193.050 136.050 195.150 ;
        RECT 137.550 193.050 138.450 200.550 ;
        RECT 139.950 198.150 141.000 203.400 ;
        RECT 139.950 196.050 142.050 198.150 ;
        RECT 142.950 197.850 145.050 199.950 ;
        RECT 143.100 196.050 144.900 197.850 ;
        RECT 136.950 190.950 139.050 193.050 ;
        RECT 139.950 189.600 141.000 196.050 ;
        RECT 146.400 192.300 147.450 209.400 ;
        RECT 157.500 203.400 159.300 215.400 ;
        RECT 149.100 198.150 150.900 199.950 ;
        RECT 152.100 198.150 153.900 199.950 ;
        RECT 157.950 198.150 159.150 203.400 ;
        RECT 166.950 202.950 169.050 205.050 ;
        RECT 171.600 203.400 173.400 215.400 ;
        RECT 183.900 203.400 187.200 215.400 ;
        RECT 200.400 209.400 202.200 215.400 ;
        RECT 212.400 209.400 214.200 215.400 ;
        RECT 224.400 209.400 226.200 215.400 ;
        RECT 160.950 201.150 162.750 202.950 ;
        RECT 160.950 199.050 163.050 201.150 ;
        RECT 148.950 196.050 151.050 198.150 ;
        RECT 151.950 196.050 154.050 198.150 ;
        RECT 154.950 194.850 157.050 196.950 ;
        RECT 157.950 196.050 160.050 198.150 ;
        RECT 155.100 193.050 156.900 194.850 ;
        RECT 158.850 192.750 160.050 196.050 ;
        RECT 160.950 195.450 163.050 196.050 ;
        RECT 167.550 195.450 168.450 202.950 ;
        RECT 171.600 202.350 174.000 203.400 ;
        RECT 170.100 198.150 171.900 199.950 ;
        RECT 169.950 196.050 172.050 198.150 ;
        RECT 160.950 194.550 168.450 195.450 ;
        RECT 172.950 195.150 174.000 202.350 ;
        RECT 176.100 198.150 177.900 199.950 ;
        RECT 179.100 198.150 180.900 199.950 ;
        RECT 185.400 198.150 186.600 203.400 ;
        RECT 200.400 201.150 201.600 209.400 ;
        RECT 212.400 201.150 213.600 209.400 ;
        RECT 224.400 201.150 225.600 209.400 ;
        RECT 233.400 204.600 235.200 215.400 ;
        RECT 239.400 214.500 247.200 215.400 ;
        RECT 239.400 204.600 241.200 214.500 ;
        RECT 233.400 203.700 241.200 204.600 ;
        RECT 242.400 202.500 244.200 213.600 ;
        RECT 245.400 203.400 247.200 214.500 ;
        RECT 253.800 203.400 255.600 215.400 ;
        RECT 256.800 204.300 258.600 215.400 ;
        RECT 262.800 204.300 264.600 215.400 ;
        RECT 268.800 209.400 270.600 215.400 ;
        RECT 269.700 209.100 270.600 209.400 ;
        RECT 274.800 209.400 276.600 215.400 ;
        RECT 284.400 209.400 286.200 215.400 ;
        RECT 299.400 209.400 301.200 215.400 ;
        RECT 311.400 209.400 313.200 215.400 ;
        RECT 274.800 209.100 276.300 209.400 ;
        RECT 269.700 208.200 276.300 209.100 ;
        RECT 256.800 203.400 264.600 204.300 ;
        RECT 240.150 201.600 244.200 202.500 ;
        RECT 190.950 198.150 192.750 199.950 ;
        RECT 175.950 196.050 178.050 198.150 ;
        RECT 178.950 196.050 181.050 198.150 ;
        RECT 160.950 193.950 163.050 194.550 ;
        RECT 172.950 193.050 175.050 195.150 ;
        RECT 181.950 194.850 184.050 196.950 ;
        RECT 184.950 196.050 187.050 198.150 ;
        RECT 182.100 193.050 183.900 194.850 ;
        RECT 143.100 191.100 150.600 192.300 ;
        RECT 158.850 191.700 162.600 192.750 ;
        RECT 143.100 190.500 144.900 191.100 ;
        RECT 139.950 188.100 143.100 189.600 ;
        RECT 121.800 183.600 123.600 186.600 ;
        RECT 130.800 183.600 132.600 186.600 ;
        RECT 141.300 183.600 143.100 188.100 ;
        RECT 148.800 183.600 150.600 191.100 ;
        RECT 152.400 188.700 160.200 190.050 ;
        RECT 152.400 183.600 154.200 188.700 ;
        RECT 158.400 183.600 160.200 188.700 ;
        RECT 161.400 189.600 162.600 191.700 ;
        RECT 161.400 183.600 163.200 189.600 ;
        RECT 172.950 186.600 174.000 193.050 ;
        RECT 185.400 192.150 186.600 196.050 ;
        RECT 187.950 194.850 190.050 196.950 ;
        RECT 190.950 196.050 193.050 198.150 ;
        RECT 196.950 197.850 199.050 199.950 ;
        RECT 199.950 199.050 202.050 201.150 ;
        RECT 197.100 196.050 198.900 197.850 ;
        RECT 187.500 193.050 189.300 194.850 ;
        RECT 185.400 191.100 189.600 192.150 ;
        RECT 179.400 189.000 187.200 189.900 ;
        RECT 188.700 189.600 189.600 191.100 ;
        RECT 200.400 191.700 201.600 199.050 ;
        RECT 202.950 197.850 205.050 199.950 ;
        RECT 208.950 197.850 211.050 199.950 ;
        RECT 211.950 199.050 214.050 201.150 ;
        RECT 203.100 196.050 204.900 197.850 ;
        RECT 209.100 196.050 210.900 197.850 ;
        RECT 212.400 191.700 213.600 199.050 ;
        RECT 214.950 197.850 217.050 199.950 ;
        RECT 220.950 197.850 223.050 199.950 ;
        RECT 223.950 199.050 226.050 201.150 ;
        RECT 215.100 196.050 216.900 197.850 ;
        RECT 221.100 196.050 222.900 197.850 ;
        RECT 224.400 191.700 225.600 199.050 ;
        RECT 226.950 197.850 229.050 199.950 ;
        RECT 233.250 198.150 235.050 199.950 ;
        RECT 240.150 198.150 241.050 201.600 ;
        RECT 245.100 198.150 246.900 199.950 ;
        RECT 254.400 198.150 255.300 203.400 ;
        RECT 265.950 202.950 268.050 205.050 ;
        RECT 259.950 201.450 262.050 202.050 ;
        RECT 266.550 201.450 267.450 202.950 ;
        RECT 259.950 200.550 267.450 201.450 ;
        RECT 259.950 199.950 262.050 200.550 ;
        RECT 269.700 199.950 270.600 208.200 ;
        RECT 275.100 204.150 276.900 205.950 ;
        RECT 271.950 201.150 273.750 202.950 ;
        RECT 274.950 202.050 277.050 204.150 ;
        RECT 278.100 201.150 279.900 202.950 ;
        RECT 284.400 201.150 285.600 209.400 ;
        RECT 299.400 201.150 300.600 209.400 ;
        RECT 227.100 196.050 228.900 197.850 ;
        RECT 232.950 196.050 235.050 198.150 ;
        RECT 235.950 194.850 238.050 196.950 ;
        RECT 236.250 193.050 238.050 194.850 ;
        RECT 238.950 196.050 241.050 198.150 ;
        RECT 200.400 190.800 204.000 191.700 ;
        RECT 212.400 190.800 216.000 191.700 ;
        RECT 224.400 190.800 228.000 191.700 ;
        RECT 172.800 183.600 174.600 186.600 ;
        RECT 179.400 183.600 181.200 189.000 ;
        RECT 185.400 184.500 187.200 189.000 ;
        RECT 188.400 185.400 190.200 189.600 ;
        RECT 191.400 184.500 193.200 189.600 ;
        RECT 185.400 183.600 193.200 184.500 ;
        RECT 202.200 183.600 204.000 190.800 ;
        RECT 214.200 183.600 216.000 190.800 ;
        RECT 226.200 183.600 228.000 190.800 ;
        RECT 238.950 189.600 240.000 196.050 ;
        RECT 241.950 194.850 244.050 196.950 ;
        RECT 244.950 196.050 247.050 198.150 ;
        RECT 253.950 196.050 256.050 198.150 ;
        RECT 268.950 197.850 271.050 199.950 ;
        RECT 271.950 199.050 274.050 201.150 ;
        RECT 277.950 199.050 280.050 201.150 ;
        RECT 280.950 197.850 283.050 199.950 ;
        RECT 283.950 199.050 286.050 201.150 ;
        RECT 241.950 193.050 243.750 194.850 ;
        RECT 238.200 183.600 240.000 189.600 ;
        RECT 254.400 189.600 255.300 196.050 ;
        RECT 256.950 194.850 259.050 196.950 ;
        RECT 260.100 195.150 261.900 196.950 ;
        RECT 257.100 193.050 258.900 194.850 ;
        RECT 259.950 193.050 262.050 195.150 ;
        RECT 262.950 194.850 265.050 196.950 ;
        RECT 263.100 193.050 264.900 194.850 ;
        RECT 269.700 193.650 270.600 197.850 ;
        RECT 281.100 196.050 282.900 197.850 ;
        RECT 269.700 192.000 273.900 193.650 ;
        RECT 254.400 187.950 259.800 189.600 ;
        RECT 258.000 183.600 259.800 187.950 ;
        RECT 272.100 183.600 273.900 192.000 ;
        RECT 284.400 191.700 285.600 199.050 ;
        RECT 286.950 197.850 289.050 199.950 ;
        RECT 295.950 197.850 298.050 199.950 ;
        RECT 298.950 199.050 301.050 201.150 ;
        RECT 287.100 196.050 288.900 197.850 ;
        RECT 296.100 196.050 297.900 197.850 ;
        RECT 299.400 191.700 300.600 199.050 ;
        RECT 301.950 197.850 304.050 199.950 ;
        RECT 308.100 198.150 309.900 199.950 ;
        RECT 302.100 196.050 303.900 197.850 ;
        RECT 307.950 196.050 310.050 198.150 ;
        RECT 311.550 192.300 312.600 209.400 ;
        RECT 318.000 203.400 319.800 215.400 ;
        RECT 328.800 209.400 330.600 215.400 ;
        RECT 325.950 204.450 328.050 205.050 ;
        RECT 323.550 203.550 328.050 204.450 ;
        RECT 313.950 197.850 316.050 199.950 ;
        RECT 318.000 198.150 319.050 203.400 ;
        RECT 314.100 196.050 315.900 197.850 ;
        RECT 316.950 196.050 319.050 198.150 ;
        RECT 319.950 198.450 322.050 199.050 ;
        RECT 323.550 198.450 324.450 203.550 ;
        RECT 325.950 202.950 328.050 203.550 ;
        RECT 329.400 201.150 330.600 209.400 ;
        RECT 344.700 203.400 346.500 215.400 ;
        RECT 356.400 209.400 358.200 215.400 ;
        RECT 356.700 209.100 358.200 209.400 ;
        RECT 362.400 209.400 364.200 215.400 ;
        RECT 362.400 209.100 363.300 209.400 ;
        RECT 356.700 208.200 363.300 209.100 ;
        RECT 356.100 204.150 357.900 205.950 ;
        RECT 341.250 201.150 343.050 202.950 ;
        RECT 319.950 197.550 324.450 198.450 ;
        RECT 325.950 197.850 328.050 199.950 ;
        RECT 328.950 199.050 331.050 201.150 ;
        RECT 319.950 196.950 322.050 197.550 ;
        RECT 326.100 196.050 327.900 197.850 ;
        RECT 284.400 190.800 288.000 191.700 ;
        RECT 299.400 190.800 303.000 191.700 ;
        RECT 286.200 183.600 288.000 190.800 ;
        RECT 301.200 183.600 303.000 190.800 ;
        RECT 308.400 191.100 315.900 192.300 ;
        RECT 308.400 183.600 310.200 191.100 ;
        RECT 314.100 190.500 315.900 191.100 ;
        RECT 318.000 189.600 319.050 196.050 ;
        RECT 329.400 191.700 330.600 199.050 ;
        RECT 331.950 197.850 334.050 199.950 ;
        RECT 340.950 199.050 343.050 201.150 ;
        RECT 344.850 198.150 346.050 203.400 ;
        RECT 353.100 201.150 354.900 202.950 ;
        RECT 355.950 202.050 358.050 204.150 ;
        RECT 359.250 201.150 361.050 202.950 ;
        RECT 350.100 198.150 351.900 199.950 ;
        RECT 352.950 199.050 355.050 201.150 ;
        RECT 358.950 199.050 361.050 201.150 ;
        RECT 362.400 199.950 363.300 208.200 ;
        RECT 367.950 205.950 370.050 208.050 ;
        RECT 364.950 202.950 367.050 205.050 ;
        RECT 332.100 196.050 333.900 197.850 ;
        RECT 343.950 196.050 346.050 198.150 ;
        RECT 343.950 192.750 345.150 196.050 ;
        RECT 346.950 194.850 349.050 196.950 ;
        RECT 349.950 196.050 352.050 198.150 ;
        RECT 361.950 197.850 364.050 199.950 ;
        RECT 347.100 193.050 348.900 194.850 ;
        RECT 362.400 193.650 363.300 197.850 ;
        RECT 365.550 196.050 366.450 202.950 ;
        RECT 368.550 196.050 369.450 205.950 ;
        RECT 374.700 203.400 376.500 215.400 ;
        RECT 387.600 203.400 389.400 215.400 ;
        RECT 397.800 203.400 399.600 215.400 ;
        RECT 400.800 204.300 402.600 215.400 ;
        RECT 406.800 204.300 408.600 215.400 ;
        RECT 400.800 203.400 408.600 204.300 ;
        RECT 414.600 203.400 416.400 215.400 ;
        RECT 421.950 208.950 424.050 211.050 ;
        RECT 371.250 201.150 373.050 202.950 ;
        RECT 370.950 199.050 373.050 201.150 ;
        RECT 374.850 198.150 376.050 203.400 ;
        RECT 387.600 202.350 390.000 203.400 ;
        RECT 382.950 199.950 385.050 202.050 ;
        RECT 380.100 198.150 381.900 199.950 ;
        RECT 373.950 196.050 376.050 198.150 ;
        RECT 364.950 193.950 367.050 196.050 ;
        RECT 367.950 193.950 370.050 196.050 ;
        RECT 315.900 188.100 319.050 189.600 ;
        RECT 327.000 190.800 330.600 191.700 ;
        RECT 341.400 191.700 345.150 192.750 ;
        RECT 359.100 192.000 363.300 193.650 ;
        RECT 373.950 192.750 375.150 196.050 ;
        RECT 376.950 194.850 379.050 196.950 ;
        RECT 379.950 196.050 382.050 198.150 ;
        RECT 377.100 193.050 378.900 194.850 ;
        RECT 315.900 183.600 317.700 188.100 ;
        RECT 327.000 183.600 328.800 190.800 ;
        RECT 341.400 189.600 342.600 191.700 ;
        RECT 340.800 183.600 342.600 189.600 ;
        RECT 343.800 188.700 351.600 190.050 ;
        RECT 343.800 183.600 345.600 188.700 ;
        RECT 349.800 183.600 351.600 188.700 ;
        RECT 359.100 183.600 360.900 192.000 ;
        RECT 371.400 191.700 375.150 192.750 ;
        RECT 379.950 192.450 382.050 193.050 ;
        RECT 383.550 192.450 384.450 199.950 ;
        RECT 386.100 198.150 387.900 199.950 ;
        RECT 385.950 196.050 388.050 198.150 ;
        RECT 371.400 189.600 372.600 191.700 ;
        RECT 379.950 191.550 384.450 192.450 ;
        RECT 388.950 195.150 390.000 202.350 ;
        RECT 392.100 198.150 393.900 199.950 ;
        RECT 398.400 198.150 399.300 203.400 ;
        RECT 414.600 202.350 417.000 203.400 ;
        RECT 400.950 201.450 403.050 202.050 ;
        RECT 400.950 200.550 411.450 201.450 ;
        RECT 400.950 199.950 403.050 200.550 ;
        RECT 391.950 196.050 394.050 198.150 ;
        RECT 397.950 196.050 400.050 198.150 ;
        RECT 388.950 193.050 391.050 195.150 ;
        RECT 379.950 190.950 382.050 191.550 ;
        RECT 370.800 183.600 372.600 189.600 ;
        RECT 373.800 188.700 381.600 190.050 ;
        RECT 373.800 183.600 375.600 188.700 ;
        RECT 379.800 183.600 381.600 188.700 ;
        RECT 388.950 186.600 390.000 193.050 ;
        RECT 398.400 189.600 399.300 196.050 ;
        RECT 400.950 194.850 403.050 196.950 ;
        RECT 404.100 195.150 405.900 196.950 ;
        RECT 401.100 193.050 402.900 194.850 ;
        RECT 403.950 193.050 406.050 195.150 ;
        RECT 406.950 194.850 409.050 196.950 ;
        RECT 407.100 193.050 408.900 194.850 ;
        RECT 410.550 193.050 411.450 200.550 ;
        RECT 413.100 198.150 414.900 199.950 ;
        RECT 412.950 196.050 415.050 198.150 ;
        RECT 415.950 195.150 417.000 202.350 ;
        RECT 419.100 198.150 420.900 199.950 ;
        RECT 418.950 196.050 421.050 198.150 ;
        RECT 415.950 193.050 418.050 195.150 ;
        RECT 409.950 190.950 412.050 193.050 ;
        RECT 398.400 187.950 403.800 189.600 ;
        RECT 388.800 183.600 390.600 186.600 ;
        RECT 402.000 183.600 403.800 187.950 ;
        RECT 415.950 186.600 417.000 193.050 ;
        RECT 418.950 192.450 421.050 193.050 ;
        RECT 422.550 192.450 423.450 208.950 ;
        RECT 427.500 203.400 429.300 215.400 ;
        RECT 433.800 209.400 435.600 215.400 ;
        RECT 418.950 191.550 423.450 192.450 ;
        RECT 427.800 198.150 429.000 203.400 ;
        RECT 434.400 202.500 435.600 209.400 ;
        RECT 445.500 203.400 447.300 215.400 ;
        RECT 460.800 209.400 462.600 215.400 ;
        RECT 470.400 209.400 472.200 215.400 ;
        RECT 429.900 201.600 435.600 202.500 ;
        RECT 429.900 200.700 431.850 201.600 ;
        RECT 427.800 196.050 430.050 198.150 ;
        RECT 418.950 190.950 421.050 191.550 ;
        RECT 427.800 189.600 429.000 196.050 ;
        RECT 430.950 192.300 431.850 200.700 ;
        RECT 434.100 198.150 435.900 199.950 ;
        RECT 440.100 198.150 441.900 199.950 ;
        RECT 445.950 198.150 447.150 203.400 ;
        RECT 448.950 201.150 450.750 202.950 ;
        RECT 461.400 201.150 462.600 209.400 ;
        RECT 470.700 209.100 472.200 209.400 ;
        RECT 476.400 209.400 478.200 215.400 ;
        RECT 476.400 209.100 477.300 209.400 ;
        RECT 470.700 208.200 477.300 209.100 ;
        RECT 470.100 204.150 471.900 205.950 ;
        RECT 467.100 201.150 468.900 202.950 ;
        RECT 469.950 202.050 472.050 204.150 ;
        RECT 473.250 201.150 475.050 202.950 ;
        RECT 448.950 199.050 451.050 201.150 ;
        RECT 433.950 196.050 436.050 198.150 ;
        RECT 439.950 196.050 442.050 198.150 ;
        RECT 442.950 194.850 445.050 196.950 ;
        RECT 445.950 196.050 448.050 198.150 ;
        RECT 457.950 197.850 460.050 199.950 ;
        RECT 460.950 199.050 463.050 201.150 ;
        RECT 458.100 196.050 459.900 197.850 ;
        RECT 443.100 193.050 444.900 194.850 ;
        RECT 429.900 191.400 431.850 192.300 ;
        RECT 446.850 192.750 448.050 196.050 ;
        RECT 446.850 191.700 450.600 192.750 ;
        RECT 461.400 191.700 462.600 199.050 ;
        RECT 463.950 197.850 466.050 199.950 ;
        RECT 466.950 199.050 469.050 201.150 ;
        RECT 472.950 199.050 475.050 201.150 ;
        RECT 476.400 199.950 477.300 208.200 ;
        RECT 487.500 203.400 489.300 215.400 ;
        RECT 490.950 207.450 493.050 208.050 ;
        RECT 490.950 206.550 495.450 207.450 ;
        RECT 490.950 205.950 493.050 206.550 ;
        RECT 475.950 197.850 478.050 199.950 ;
        RECT 482.100 198.150 483.900 199.950 ;
        RECT 487.950 198.150 489.150 203.400 ;
        RECT 490.950 201.150 492.750 202.950 ;
        RECT 490.950 199.050 493.050 201.150 ;
        RECT 464.100 196.050 465.900 197.850 ;
        RECT 476.400 193.650 477.300 197.850 ;
        RECT 481.950 196.050 484.050 198.150 ;
        RECT 484.950 194.850 487.050 196.950 ;
        RECT 487.950 196.050 490.050 198.150 ;
        RECT 494.550 196.050 495.450 206.550 ;
        RECT 502.500 203.400 504.300 215.400 ;
        RECT 518.400 209.400 520.200 215.400 ;
        RECT 527.400 209.400 529.200 215.400 ;
        RECT 536.400 209.400 538.200 215.400 ;
        RECT 497.100 198.150 498.900 199.950 ;
        RECT 502.950 198.150 504.150 203.400 ;
        RECT 505.950 201.150 507.750 202.950 ;
        RECT 505.950 199.050 508.050 201.150 ;
        RECT 496.950 196.050 499.050 198.150 ;
        RECT 429.900 190.500 435.000 191.400 ;
        RECT 415.800 183.600 417.600 186.600 ;
        RECT 427.500 183.600 429.300 189.600 ;
        RECT 433.800 186.600 435.000 190.500 ;
        RECT 440.400 188.700 448.200 190.050 ;
        RECT 433.800 183.600 435.600 186.600 ;
        RECT 440.400 183.600 442.200 188.700 ;
        RECT 446.400 183.600 448.200 188.700 ;
        RECT 449.400 189.600 450.600 191.700 ;
        RECT 459.000 190.800 462.600 191.700 ;
        RECT 473.100 192.000 477.300 193.650 ;
        RECT 485.100 193.050 486.900 194.850 ;
        RECT 488.850 192.750 490.050 196.050 ;
        RECT 493.950 193.950 496.050 196.050 ;
        RECT 499.950 194.850 502.050 196.950 ;
        RECT 502.950 196.050 505.050 198.150 ;
        RECT 518.400 196.950 519.600 209.400 ;
        RECT 527.400 196.950 528.600 209.400 ;
        RECT 536.700 209.100 538.200 209.400 ;
        RECT 542.400 209.400 544.200 215.400 ;
        RECT 553.800 209.400 555.600 215.400 ;
        RECT 563.400 209.400 565.200 215.400 ;
        RECT 542.400 209.100 543.300 209.400 ;
        RECT 536.700 208.200 543.300 209.100 ;
        RECT 536.100 204.150 537.900 205.950 ;
        RECT 529.950 199.950 532.050 202.050 ;
        RECT 533.100 201.150 534.900 202.950 ;
        RECT 535.950 202.050 538.050 204.150 ;
        RECT 539.250 201.150 541.050 202.950 ;
        RECT 500.100 193.050 501.900 194.850 ;
        RECT 503.850 192.750 505.050 196.050 ;
        RECT 515.100 195.150 516.900 196.950 ;
        RECT 514.950 193.050 517.050 195.150 ;
        RECT 517.950 194.850 520.050 196.950 ;
        RECT 524.100 195.150 525.900 196.950 ;
        RECT 449.400 183.600 451.200 189.600 ;
        RECT 459.000 183.600 460.800 190.800 ;
        RECT 473.100 183.600 474.900 192.000 ;
        RECT 488.850 191.700 492.600 192.750 ;
        RECT 503.850 191.700 507.600 192.750 ;
        RECT 482.400 188.700 490.200 190.050 ;
        RECT 482.400 183.600 484.200 188.700 ;
        RECT 488.400 183.600 490.200 188.700 ;
        RECT 491.400 189.600 492.600 191.700 ;
        RECT 491.400 183.600 493.200 189.600 ;
        RECT 497.400 188.700 505.200 190.050 ;
        RECT 497.400 183.600 499.200 188.700 ;
        RECT 503.400 183.600 505.200 188.700 ;
        RECT 506.400 189.600 507.600 191.700 ;
        RECT 506.400 183.600 508.200 189.600 ;
        RECT 518.400 186.600 519.600 194.850 ;
        RECT 523.950 193.050 526.050 195.150 ;
        RECT 526.950 194.850 529.050 196.950 ;
        RECT 530.550 195.450 531.450 199.950 ;
        RECT 532.950 199.050 535.050 201.150 ;
        RECT 538.950 199.050 541.050 201.150 ;
        RECT 542.400 199.950 543.300 208.200 ;
        RECT 550.950 207.450 553.050 208.050 ;
        RECT 545.550 206.550 553.050 207.450 ;
        RECT 541.950 197.850 544.050 199.950 ;
        RECT 535.950 195.450 538.050 196.050 ;
        RECT 527.400 186.600 528.600 194.850 ;
        RECT 530.550 194.550 538.050 195.450 ;
        RECT 535.950 193.950 538.050 194.550 ;
        RECT 542.400 193.650 543.300 197.850 ;
        RECT 545.550 196.050 546.450 206.550 ;
        RECT 550.950 205.950 553.050 206.550 ;
        RECT 554.400 201.150 555.600 209.400 ;
        RECT 550.950 197.850 553.050 199.950 ;
        RECT 553.950 199.050 556.050 201.150 ;
        RECT 551.100 196.050 552.900 197.850 ;
        RECT 544.950 193.950 547.050 196.050 ;
        RECT 539.100 192.000 543.300 193.650 ;
        RECT 518.400 183.600 520.200 186.600 ;
        RECT 527.400 183.600 529.200 186.600 ;
        RECT 539.100 183.600 540.900 192.000 ;
        RECT 554.400 191.700 555.600 199.050 ;
        RECT 556.950 197.850 559.050 199.950 ;
        RECT 560.100 198.150 561.900 199.950 ;
        RECT 557.100 196.050 558.900 197.850 ;
        RECT 559.950 196.050 562.050 198.150 ;
        RECT 563.550 192.300 564.600 209.400 ;
        RECT 570.000 203.400 571.800 215.400 ;
        RECT 575.400 204.600 577.200 215.400 ;
        RECT 581.400 214.500 589.200 215.400 ;
        RECT 581.400 204.600 583.200 214.500 ;
        RECT 575.400 203.700 583.200 204.600 ;
        RECT 565.950 197.850 568.050 199.950 ;
        RECT 570.000 198.150 571.050 203.400 ;
        RECT 584.400 202.500 586.200 213.600 ;
        RECT 587.400 203.400 589.200 214.500 ;
        RECT 599.400 209.400 601.200 215.400 ;
        RECT 595.950 204.450 598.050 205.050 ;
        RECT 593.550 203.550 598.050 204.450 ;
        RECT 582.150 201.600 586.200 202.500 ;
        RECT 575.250 198.150 577.050 199.950 ;
        RECT 582.150 198.150 583.050 201.600 ;
        RECT 593.550 201.450 594.450 203.550 ;
        RECT 595.950 202.950 598.050 203.550 ;
        RECT 590.550 200.550 594.450 201.450 ;
        RECT 587.100 198.150 588.900 199.950 ;
        RECT 566.100 196.050 567.900 197.850 ;
        RECT 568.950 196.050 571.050 198.150 ;
        RECT 574.950 196.050 577.050 198.150 ;
        RECT 552.000 190.800 555.600 191.700 ;
        RECT 560.400 191.100 567.900 192.300 ;
        RECT 552.000 183.600 553.800 190.800 ;
        RECT 560.400 183.600 562.200 191.100 ;
        RECT 566.100 190.500 567.900 191.100 ;
        RECT 570.000 189.600 571.050 196.050 ;
        RECT 577.950 194.850 580.050 196.950 ;
        RECT 578.250 193.050 580.050 194.850 ;
        RECT 580.950 196.050 583.050 198.150 ;
        RECT 580.950 189.600 582.000 196.050 ;
        RECT 583.950 194.850 586.050 196.950 ;
        RECT 586.950 196.050 589.050 198.150 ;
        RECT 583.950 193.050 585.750 194.850 ;
        RECT 586.950 192.450 589.050 193.050 ;
        RECT 590.550 192.450 591.450 200.550 ;
        RECT 596.100 198.150 597.900 199.950 ;
        RECT 595.950 196.050 598.050 198.150 ;
        RECT 586.950 191.550 591.450 192.450 ;
        RECT 599.550 192.300 600.600 209.400 ;
        RECT 606.000 203.400 607.800 215.400 ;
        RECT 616.500 203.400 618.300 215.400 ;
        RECT 629.400 209.400 631.200 215.400 ;
        RECT 638.400 209.400 640.200 215.400 ;
        RECT 650.400 209.400 652.200 215.400 ;
        RECT 601.950 197.850 604.050 199.950 ;
        RECT 606.000 198.150 607.050 203.400 ;
        RECT 611.100 198.150 612.900 199.950 ;
        RECT 616.950 198.150 618.150 203.400 ;
        RECT 619.950 201.150 621.750 202.950 ;
        RECT 619.950 199.050 622.050 201.150 ;
        RECT 602.100 196.050 603.900 197.850 ;
        RECT 604.950 196.050 607.050 198.150 ;
        RECT 610.950 196.050 613.050 198.150 ;
        RECT 586.950 190.950 589.050 191.550 ;
        RECT 596.400 191.100 603.900 192.300 ;
        RECT 567.900 188.100 571.050 189.600 ;
        RECT 567.900 183.600 569.700 188.100 ;
        RECT 580.200 183.600 582.000 189.600 ;
        RECT 596.400 183.600 598.200 191.100 ;
        RECT 602.100 190.500 603.900 191.100 ;
        RECT 606.000 189.600 607.050 196.050 ;
        RECT 613.950 194.850 616.050 196.950 ;
        RECT 616.950 196.050 619.050 198.150 ;
        RECT 629.400 196.950 630.600 209.400 ;
        RECT 634.950 204.450 637.050 205.050 ;
        RECT 632.550 203.550 637.050 204.450 ;
        RECT 614.100 193.050 615.900 194.850 ;
        RECT 617.850 192.750 619.050 196.050 ;
        RECT 626.100 195.150 627.900 196.950 ;
        RECT 625.950 193.050 628.050 195.150 ;
        RECT 628.950 194.850 631.050 196.950 ;
        RECT 617.850 191.700 621.600 192.750 ;
        RECT 603.900 188.100 607.050 189.600 ;
        RECT 611.400 188.700 619.200 190.050 ;
        RECT 603.900 183.600 605.700 188.100 ;
        RECT 611.400 183.600 613.200 188.700 ;
        RECT 617.400 183.600 619.200 188.700 ;
        RECT 620.400 189.600 621.600 191.700 ;
        RECT 620.400 183.600 622.200 189.600 ;
        RECT 629.400 186.600 630.600 194.850 ;
        RECT 632.550 193.050 633.450 203.550 ;
        RECT 634.950 202.950 637.050 203.550 ;
        RECT 638.400 201.150 639.600 209.400 ;
        RECT 650.700 209.100 652.200 209.400 ;
        RECT 656.400 209.400 658.200 215.400 ;
        RECT 656.400 209.100 657.300 209.400 ;
        RECT 650.700 208.200 657.300 209.100 ;
        RECT 650.100 204.150 651.900 205.950 ;
        RECT 647.100 201.150 648.900 202.950 ;
        RECT 649.950 202.050 652.050 204.150 ;
        RECT 653.250 201.150 655.050 202.950 ;
        RECT 634.950 197.850 637.050 199.950 ;
        RECT 637.950 199.050 640.050 201.150 ;
        RECT 635.100 196.050 636.900 197.850 ;
        RECT 631.950 190.950 634.050 193.050 ;
        RECT 638.400 191.700 639.600 199.050 ;
        RECT 640.950 197.850 643.050 199.950 ;
        RECT 646.950 199.050 649.050 201.150 ;
        RECT 652.950 199.050 655.050 201.150 ;
        RECT 656.400 199.950 657.300 208.200 ;
        RECT 665.400 204.300 667.200 215.400 ;
        RECT 671.400 204.300 673.200 215.400 ;
        RECT 665.400 203.400 673.200 204.300 ;
        RECT 674.400 203.400 676.200 215.400 ;
        RECT 683.400 209.400 685.200 215.400 ;
        RECT 683.700 209.100 685.200 209.400 ;
        RECT 689.400 209.400 691.200 215.400 ;
        RECT 689.400 209.100 690.300 209.400 ;
        RECT 683.700 208.200 690.300 209.100 ;
        RECT 683.100 204.150 684.900 205.950 ;
        RECT 655.950 197.850 658.050 199.950 ;
        RECT 674.700 198.150 675.600 203.400 ;
        RECT 680.100 201.150 681.900 202.950 ;
        RECT 682.950 202.050 685.050 204.150 ;
        RECT 686.250 201.150 688.050 202.950 ;
        RECT 679.950 199.050 682.050 201.150 ;
        RECT 685.950 199.050 688.050 201.150 ;
        RECT 689.400 199.950 690.300 208.200 ;
        RECT 695.400 204.300 697.200 215.400 ;
        RECT 701.400 204.300 703.200 215.400 ;
        RECT 695.400 203.400 703.200 204.300 ;
        RECT 704.400 203.400 706.200 215.400 ;
        RECT 715.500 203.400 717.300 215.400 ;
        RECT 728.400 209.400 730.200 215.400 ;
        RECT 728.700 209.100 730.200 209.400 ;
        RECT 734.400 209.400 736.200 215.400 ;
        RECT 743.400 209.400 745.200 215.400 ;
        RECT 734.400 209.100 735.300 209.400 ;
        RECT 728.700 208.200 735.300 209.100 ;
        RECT 743.700 209.100 745.200 209.400 ;
        RECT 749.400 209.400 751.200 215.400 ;
        RECT 749.400 209.100 750.300 209.400 ;
        RECT 743.700 208.200 750.300 209.100 ;
        RECT 724.950 207.450 727.050 208.050 ;
        RECT 722.550 206.550 727.050 207.450 ;
        RECT 641.100 196.050 642.900 197.850 ;
        RECT 656.400 193.650 657.300 197.850 ;
        RECT 664.950 194.850 667.050 196.950 ;
        RECT 668.100 195.150 669.900 196.950 ;
        RECT 653.100 192.000 657.300 193.650 ;
        RECT 665.100 193.050 666.900 194.850 ;
        RECT 667.950 193.050 670.050 195.150 ;
        RECT 670.950 194.850 673.050 196.950 ;
        RECT 673.950 196.050 676.050 198.150 ;
        RECT 688.950 197.850 691.050 199.950 ;
        RECT 704.700 198.150 705.600 203.400 ;
        RECT 710.100 198.150 711.900 199.950 ;
        RECT 715.950 198.150 717.150 203.400 ;
        RECT 718.950 201.150 720.750 202.950 ;
        RECT 718.950 199.050 721.050 201.150 ;
        RECT 671.100 193.050 672.900 194.850 ;
        RECT 638.400 190.800 642.000 191.700 ;
        RECT 629.400 183.600 631.200 186.600 ;
        RECT 640.200 183.600 642.000 190.800 ;
        RECT 653.100 183.600 654.900 192.000 ;
        RECT 674.700 189.600 675.600 196.050 ;
        RECT 689.400 193.650 690.300 197.850 ;
        RECT 694.950 194.850 697.050 196.950 ;
        RECT 698.100 195.150 699.900 196.950 ;
        RECT 670.200 187.950 675.600 189.600 ;
        RECT 686.100 192.000 690.300 193.650 ;
        RECT 695.100 193.050 696.900 194.850 ;
        RECT 697.950 193.050 700.050 195.150 ;
        RECT 700.950 194.850 703.050 196.950 ;
        RECT 703.950 196.050 706.050 198.150 ;
        RECT 709.950 196.050 712.050 198.150 ;
        RECT 701.100 193.050 702.900 194.850 ;
        RECT 670.200 183.600 672.000 187.950 ;
        RECT 686.100 183.600 687.900 192.000 ;
        RECT 704.700 189.600 705.600 196.050 ;
        RECT 712.950 194.850 715.050 196.950 ;
        RECT 715.950 196.050 718.050 198.150 ;
        RECT 713.100 193.050 714.900 194.850 ;
        RECT 716.850 192.750 718.050 196.050 ;
        RECT 718.950 195.450 721.050 196.050 ;
        RECT 722.550 195.450 723.450 206.550 ;
        RECT 724.950 205.950 727.050 206.550 ;
        RECT 728.100 204.150 729.900 205.950 ;
        RECT 725.100 201.150 726.900 202.950 ;
        RECT 727.950 202.050 730.050 204.150 ;
        RECT 731.250 201.150 733.050 202.950 ;
        RECT 724.950 199.050 727.050 201.150 ;
        RECT 730.950 199.050 733.050 201.150 ;
        RECT 734.400 199.950 735.300 208.200 ;
        RECT 743.100 204.150 744.900 205.950 ;
        RECT 740.100 201.150 741.900 202.950 ;
        RECT 742.950 202.050 745.050 204.150 ;
        RECT 746.250 201.150 748.050 202.950 ;
        RECT 733.950 197.850 736.050 199.950 ;
        RECT 739.950 199.050 742.050 201.150 ;
        RECT 745.950 199.050 748.050 201.150 ;
        RECT 749.400 199.950 750.300 208.200 ;
        RECT 761.700 203.400 763.500 215.400 ;
        RECT 758.250 201.150 760.050 202.950 ;
        RECT 748.950 197.850 751.050 199.950 ;
        RECT 757.950 199.050 760.050 201.150 ;
        RECT 761.850 198.150 763.050 203.400 ;
        RECT 767.100 198.150 768.900 199.950 ;
        RECT 718.950 194.550 723.450 195.450 ;
        RECT 718.950 193.950 721.050 194.550 ;
        RECT 734.400 193.650 735.300 197.850 ;
        RECT 749.400 193.650 750.300 197.850 ;
        RECT 716.850 191.700 720.600 192.750 ;
        RECT 700.200 187.950 705.600 189.600 ;
        RECT 710.400 188.700 718.200 190.050 ;
        RECT 700.200 183.600 702.000 187.950 ;
        RECT 710.400 183.600 712.200 188.700 ;
        RECT 716.400 183.600 718.200 188.700 ;
        RECT 719.400 189.600 720.600 191.700 ;
        RECT 731.100 192.000 735.300 193.650 ;
        RECT 746.100 192.000 750.300 193.650 ;
        RECT 760.950 196.050 763.050 198.150 ;
        RECT 760.950 192.750 762.150 196.050 ;
        RECT 763.950 194.850 766.050 196.950 ;
        RECT 766.950 196.050 769.050 198.150 ;
        RECT 764.100 193.050 765.900 194.850 ;
        RECT 719.400 183.600 721.200 189.600 ;
        RECT 731.100 183.600 732.900 192.000 ;
        RECT 746.100 183.600 747.900 192.000 ;
        RECT 758.400 191.700 762.150 192.750 ;
        RECT 758.400 189.600 759.600 191.700 ;
        RECT 757.800 183.600 759.600 189.600 ;
        RECT 760.800 188.700 768.600 190.050 ;
        RECT 760.800 183.600 762.600 188.700 ;
        RECT 766.800 183.600 768.600 188.700 ;
        RECT 10.800 176.400 12.600 179.400 ;
        RECT 20.400 176.400 22.200 179.400 ;
        RECT 10.950 169.950 12.000 176.400 ;
        RECT 21.300 172.200 22.200 176.400 ;
        RECT 26.400 173.400 28.200 179.400 ;
        RECT 21.300 171.300 24.750 172.200 ;
        RECT 22.950 170.400 24.750 171.300 ;
        RECT 10.950 167.850 13.050 169.950 ;
        RECT 16.950 167.850 19.050 169.950 ;
        RECT 7.950 164.850 10.050 166.950 ;
        RECT 8.100 163.050 9.900 164.850 ;
        RECT 10.950 160.650 12.000 167.850 ;
        RECT 13.950 164.850 16.050 166.950 ;
        RECT 17.100 166.050 18.900 167.850 ;
        RECT 19.950 164.850 22.050 166.950 ;
        RECT 14.100 163.050 15.900 164.850 ;
        RECT 20.100 163.050 21.900 164.850 ;
        RECT 23.700 162.150 24.600 170.400 ;
        RECT 27.000 168.150 28.050 173.400 ;
        RECT 41.100 171.000 42.900 179.400 ;
        RECT 22.800 162.000 24.600 162.150 ;
        RECT 9.600 159.600 12.000 160.650 ;
        RECT 17.400 160.800 24.600 162.000 ;
        RECT 17.400 159.600 18.600 160.800 ;
        RECT 22.800 160.350 24.600 160.800 ;
        RECT 25.950 166.050 28.050 168.150 ;
        RECT 38.700 169.350 42.900 171.000 ;
        RECT 53.400 176.400 55.200 179.400 ;
        RECT 9.600 147.600 11.400 159.600 ;
        RECT 17.400 147.600 19.200 159.600 ;
        RECT 25.950 159.450 27.300 166.050 ;
        RECT 38.700 165.150 39.600 169.350 ;
        RECT 49.950 167.850 52.050 169.950 ;
        RECT 53.400 168.150 54.600 176.400 ;
        RECT 59.400 174.300 61.200 179.400 ;
        RECT 65.400 174.300 67.200 179.400 ;
        RECT 59.400 172.950 67.200 174.300 ;
        RECT 68.400 173.400 70.200 179.400 ;
        RECT 76.800 173.400 78.600 179.400 ;
        RECT 82.800 176.400 84.600 179.400 ;
        RECT 68.400 171.300 69.600 173.400 ;
        RECT 65.850 170.250 69.600 171.300 ;
        RECT 62.100 168.150 63.900 169.950 ;
        RECT 50.100 166.050 51.900 167.850 ;
        RECT 52.950 166.050 55.050 168.150 ;
        RECT 37.950 163.050 40.050 165.150 ;
        RECT 24.900 158.100 27.300 159.450 ;
        RECT 24.900 147.600 26.700 158.100 ;
        RECT 38.700 154.800 39.600 163.050 ;
        RECT 40.950 161.850 43.050 163.950 ;
        RECT 46.950 161.850 49.050 163.950 ;
        RECT 40.950 160.050 42.750 161.850 ;
        RECT 43.950 158.850 46.050 160.950 ;
        RECT 47.100 160.050 48.900 161.850 ;
        RECT 44.100 157.050 45.900 158.850 ;
        RECT 38.700 153.900 45.300 154.800 ;
        RECT 38.700 153.600 39.600 153.900 ;
        RECT 37.800 147.600 39.600 153.600 ;
        RECT 43.800 153.600 45.300 153.900 ;
        RECT 53.400 153.600 54.600 166.050 ;
        RECT 58.950 164.850 61.050 166.950 ;
        RECT 61.950 166.050 64.050 168.150 ;
        RECT 65.850 166.950 67.050 170.250 ;
        RECT 64.950 164.850 67.050 166.950 ;
        RECT 76.950 168.150 78.000 173.400 ;
        RECT 82.800 172.200 83.700 176.400 ;
        RECT 94.200 172.200 96.000 179.400 ;
        RECT 80.250 171.300 83.700 172.200 ;
        RECT 92.400 171.300 96.000 172.200 ;
        RECT 80.250 170.400 82.050 171.300 ;
        RECT 76.950 166.050 79.050 168.150 ;
        RECT 59.100 163.050 60.900 164.850 ;
        RECT 64.950 159.600 66.150 164.850 ;
        RECT 67.950 161.850 70.050 163.950 ;
        RECT 67.950 160.050 69.750 161.850 ;
        RECT 43.800 147.600 45.600 153.600 ;
        RECT 53.400 147.600 55.200 153.600 ;
        RECT 64.500 147.600 66.300 159.600 ;
        RECT 77.700 159.450 79.050 166.050 ;
        RECT 80.400 162.150 81.300 170.400 ;
        RECT 85.950 167.850 88.050 169.950 ;
        RECT 82.950 164.850 85.050 166.950 ;
        RECT 86.100 166.050 87.900 167.850 ;
        RECT 89.100 165.150 90.900 166.950 ;
        RECT 83.100 163.050 84.900 164.850 ;
        RECT 88.950 163.050 91.050 165.150 ;
        RECT 92.400 163.950 93.600 171.300 ;
        RECT 110.100 171.000 111.900 179.400 ;
        RECT 124.800 176.400 126.600 179.400 ;
        RECT 133.800 176.400 135.600 179.400 ;
        RECT 107.700 169.350 111.900 171.000 ;
        RECT 95.100 165.150 96.900 166.950 ;
        RECT 107.700 165.150 108.600 169.350 ;
        RECT 125.400 168.150 126.600 176.400 ;
        RECT 124.950 166.050 127.050 168.150 ;
        RECT 127.950 167.850 130.050 169.950 ;
        RECT 134.400 168.150 135.600 176.400 ;
        RECT 144.000 172.200 145.800 179.400 ;
        RECT 157.800 176.400 159.600 179.400 ;
        RECT 144.000 171.300 147.600 172.200 ;
        RECT 128.100 166.050 129.900 167.850 ;
        RECT 133.950 166.050 136.050 168.150 ;
        RECT 136.950 167.850 139.050 169.950 ;
        RECT 137.100 166.050 138.900 167.850 ;
        RECT 80.400 162.000 82.200 162.150 ;
        RECT 80.400 160.800 87.600 162.000 ;
        RECT 91.950 161.850 94.050 163.950 ;
        RECT 94.950 163.050 97.050 165.150 ;
        RECT 106.950 163.050 109.050 165.150 ;
        RECT 80.400 160.350 82.200 160.800 ;
        RECT 86.400 159.600 87.600 160.800 ;
        RECT 77.700 158.100 80.100 159.450 ;
        RECT 78.300 147.600 80.100 158.100 ;
        RECT 85.800 147.600 87.600 159.600 ;
        RECT 92.400 153.600 93.600 161.850 ;
        RECT 107.700 154.800 108.600 163.050 ;
        RECT 109.950 161.850 112.050 163.950 ;
        RECT 115.950 161.850 118.050 163.950 ;
        RECT 109.950 160.050 111.750 161.850 ;
        RECT 112.950 158.850 115.050 160.950 ;
        RECT 116.100 160.050 117.900 161.850 ;
        RECT 113.100 157.050 114.900 158.850 ;
        RECT 107.700 153.900 114.300 154.800 ;
        RECT 107.700 153.600 108.600 153.900 ;
        RECT 92.400 147.600 94.200 153.600 ;
        RECT 106.800 147.600 108.600 153.600 ;
        RECT 112.800 153.600 114.300 153.900 ;
        RECT 125.400 153.600 126.600 166.050 ;
        RECT 134.400 153.600 135.600 166.050 ;
        RECT 143.100 165.150 144.900 166.950 ;
        RECT 142.950 163.050 145.050 165.150 ;
        RECT 146.400 163.950 147.600 171.300 ;
        RECT 158.400 168.150 159.600 176.400 ;
        RECT 164.400 174.300 166.200 179.400 ;
        RECT 170.400 174.300 172.200 179.400 ;
        RECT 164.400 172.950 172.200 174.300 ;
        RECT 173.400 173.400 175.200 179.400 ;
        RECT 181.800 173.400 183.600 179.400 ;
        RECT 173.400 171.300 174.600 173.400 ;
        RECT 170.850 170.250 174.600 171.300 ;
        RECT 182.400 171.300 183.600 173.400 ;
        RECT 184.800 174.300 186.600 179.400 ;
        RECT 190.800 174.300 192.600 179.400 ;
        RECT 184.800 172.950 192.600 174.300 ;
        RECT 200.400 176.400 202.200 179.400 ;
        RECT 209.400 176.400 211.200 179.400 ;
        RECT 182.400 170.250 186.150 171.300 ;
        RECT 149.100 165.150 150.900 166.950 ;
        RECT 157.950 166.050 160.050 168.150 ;
        RECT 160.950 167.850 163.050 169.950 ;
        RECT 167.100 168.150 168.900 169.950 ;
        RECT 161.100 166.050 162.900 167.850 ;
        RECT 145.950 161.850 148.050 163.950 ;
        RECT 148.950 163.050 151.050 165.150 ;
        RECT 146.400 153.600 147.600 161.850 ;
        RECT 158.400 153.600 159.600 166.050 ;
        RECT 163.950 164.850 166.050 166.950 ;
        RECT 166.950 166.050 169.050 168.150 ;
        RECT 170.850 166.950 172.050 170.250 ;
        RECT 169.950 164.850 172.050 166.950 ;
        RECT 184.950 166.950 186.150 170.250 ;
        RECT 188.100 168.150 189.900 169.950 ;
        RECT 184.950 164.850 187.050 166.950 ;
        RECT 187.950 166.050 190.050 168.150 ;
        RECT 196.950 167.850 199.050 169.950 ;
        RECT 200.400 168.150 201.600 176.400 ;
        RECT 190.950 164.850 193.050 166.950 ;
        RECT 197.100 166.050 198.900 167.850 ;
        RECT 199.950 166.050 202.050 168.150 ;
        RECT 205.950 167.850 208.050 169.950 ;
        RECT 209.400 168.150 210.600 176.400 ;
        RECT 220.200 175.050 222.000 179.400 ;
        RECT 220.200 173.400 225.600 175.050 ;
        RECT 215.100 168.150 216.900 169.950 ;
        RECT 206.100 166.050 207.900 167.850 ;
        RECT 208.950 166.050 211.050 168.150 ;
        RECT 214.950 166.050 217.050 168.150 ;
        RECT 217.950 167.850 220.050 169.950 ;
        RECT 221.100 168.150 222.900 169.950 ;
        RECT 218.100 166.050 219.900 167.850 ;
        RECT 220.950 166.050 223.050 168.150 ;
        RECT 224.700 166.950 225.600 173.400 ;
        RECT 239.100 171.000 240.900 179.400 ;
        RECT 254.100 171.000 255.900 179.400 ;
        RECT 266.400 176.400 268.200 179.400 ;
        RECT 277.800 176.400 279.600 179.400 ;
        RECT 239.100 169.350 243.300 171.000 ;
        RECT 164.100 163.050 165.900 164.850 ;
        RECT 169.950 159.600 171.150 164.850 ;
        RECT 172.950 161.850 175.050 163.950 ;
        RECT 181.950 161.850 184.050 163.950 ;
        RECT 172.950 160.050 174.750 161.850 ;
        RECT 182.250 160.050 184.050 161.850 ;
        RECT 185.850 159.600 187.050 164.850 ;
        RECT 191.100 163.050 192.900 164.850 ;
        RECT 112.800 147.600 114.600 153.600 ;
        RECT 124.800 147.600 126.600 153.600 ;
        RECT 133.800 147.600 135.600 153.600 ;
        RECT 145.800 147.600 147.600 153.600 ;
        RECT 157.800 147.600 159.600 153.600 ;
        RECT 169.500 147.600 171.300 159.600 ;
        RECT 185.700 147.600 187.500 159.600 ;
        RECT 200.400 153.600 201.600 166.050 ;
        RECT 209.400 153.600 210.600 166.050 ;
        RECT 223.950 164.850 226.050 166.950 ;
        RECT 242.400 165.150 243.300 169.350 ;
        RECT 251.700 169.350 255.900 171.000 ;
        RECT 267.000 169.950 268.050 176.400 ;
        RECT 251.700 165.150 252.600 169.350 ;
        RECT 265.950 167.850 268.050 169.950 ;
        RECT 278.400 168.150 279.600 176.400 ;
        RECT 289.800 173.400 291.600 179.400 ;
        RECT 290.400 171.300 291.600 173.400 ;
        RECT 292.800 174.300 294.600 179.400 ;
        RECT 298.800 174.300 300.600 179.400 ;
        RECT 292.800 172.950 300.600 174.300 ;
        RECT 305.400 176.400 307.200 179.400 ;
        RECT 313.800 176.400 315.600 179.400 ;
        RECT 290.400 170.250 294.150 171.300 ;
        RECT 224.700 159.600 225.600 164.850 ;
        RECT 232.950 161.850 235.050 163.950 ;
        RECT 238.950 161.850 241.050 163.950 ;
        RECT 241.950 163.050 244.050 165.150 ;
        RECT 250.950 163.050 253.050 165.150 ;
        RECT 262.950 164.850 265.050 166.950 ;
        RECT 233.100 160.050 234.900 161.850 ;
        RECT 215.400 158.700 223.200 159.600 ;
        RECT 200.400 147.600 202.200 153.600 ;
        RECT 209.400 147.600 211.200 153.600 ;
        RECT 215.400 147.600 217.200 158.700 ;
        RECT 221.400 147.600 223.200 158.700 ;
        RECT 224.400 147.600 226.200 159.600 ;
        RECT 235.950 158.850 238.050 160.950 ;
        RECT 239.250 160.050 241.050 161.850 ;
        RECT 236.100 157.050 237.900 158.850 ;
        RECT 242.400 154.800 243.300 163.050 ;
        RECT 236.700 153.900 243.300 154.800 ;
        RECT 236.700 153.600 238.200 153.900 ;
        RECT 236.400 147.600 238.200 153.600 ;
        RECT 242.400 153.600 243.300 153.900 ;
        RECT 251.700 154.800 252.600 163.050 ;
        RECT 253.950 161.850 256.050 163.950 ;
        RECT 259.950 161.850 262.050 163.950 ;
        RECT 263.100 163.050 264.900 164.850 ;
        RECT 253.950 160.050 255.750 161.850 ;
        RECT 256.950 158.850 259.050 160.950 ;
        RECT 260.100 160.050 261.900 161.850 ;
        RECT 267.000 160.650 268.050 167.850 ;
        RECT 268.950 164.850 271.050 166.950 ;
        RECT 277.950 166.050 280.050 168.150 ;
        RECT 280.950 167.850 283.050 169.950 ;
        RECT 281.100 166.050 282.900 167.850 ;
        RECT 292.950 166.950 294.150 170.250 ;
        RECT 296.100 168.150 297.900 169.950 ;
        RECT 269.100 163.050 270.900 164.850 ;
        RECT 267.000 159.600 269.400 160.650 ;
        RECT 257.100 157.050 258.900 158.850 ;
        RECT 251.700 153.900 258.300 154.800 ;
        RECT 251.700 153.600 252.600 153.900 ;
        RECT 242.400 147.600 244.200 153.600 ;
        RECT 250.800 147.600 252.600 153.600 ;
        RECT 256.800 153.600 258.300 153.900 ;
        RECT 256.800 147.600 258.600 153.600 ;
        RECT 267.600 147.600 269.400 159.600 ;
        RECT 278.400 153.600 279.600 166.050 ;
        RECT 292.950 164.850 295.050 166.950 ;
        RECT 295.950 166.050 298.050 168.150 ;
        RECT 301.950 167.850 304.050 169.950 ;
        RECT 305.400 168.150 306.600 176.400 ;
        RECT 314.400 168.150 315.600 176.400 ;
        RECT 326.100 171.000 327.900 179.400 ;
        RECT 339.000 172.200 340.800 179.400 ;
        RECT 350.400 176.400 352.200 179.400 ;
        RECT 339.000 171.300 342.600 172.200 ;
        RECT 298.950 164.850 301.050 166.950 ;
        RECT 302.100 166.050 303.900 167.850 ;
        RECT 304.950 166.050 307.050 168.150 ;
        RECT 313.950 166.050 316.050 168.150 ;
        RECT 316.950 167.850 319.050 169.950 ;
        RECT 326.100 169.350 330.300 171.000 ;
        RECT 317.100 166.050 318.900 167.850 ;
        RECT 289.950 161.850 292.050 163.950 ;
        RECT 290.250 160.050 292.050 161.850 ;
        RECT 293.850 159.600 295.050 164.850 ;
        RECT 299.100 163.050 300.900 164.850 ;
        RECT 277.800 147.600 279.600 153.600 ;
        RECT 293.700 147.600 295.500 159.600 ;
        RECT 305.400 153.600 306.600 166.050 ;
        RECT 314.400 153.600 315.600 166.050 ;
        RECT 329.400 165.150 330.300 169.350 ;
        RECT 338.100 165.150 339.900 166.950 ;
        RECT 319.950 161.850 322.050 163.950 ;
        RECT 325.950 161.850 328.050 163.950 ;
        RECT 328.950 163.050 331.050 165.150 ;
        RECT 337.950 163.050 340.050 165.150 ;
        RECT 341.400 163.950 342.600 171.300 ;
        RECT 346.950 167.850 349.050 169.950 ;
        RECT 350.400 168.150 351.600 176.400 ;
        RECT 361.800 173.400 363.600 179.400 ;
        RECT 362.400 171.300 363.600 173.400 ;
        RECT 364.800 174.300 366.600 179.400 ;
        RECT 370.800 174.300 372.600 179.400 ;
        RECT 364.800 172.950 372.600 174.300 ;
        RECT 384.000 173.400 385.800 179.400 ;
        RECT 362.400 170.250 366.150 171.300 ;
        RECT 361.950 168.450 364.050 169.050 ;
        RECT 344.100 165.150 345.900 166.950 ;
        RECT 347.100 166.050 348.900 167.850 ;
        RECT 349.950 166.050 352.050 168.150 ;
        RECT 359.550 167.550 364.050 168.450 ;
        RECT 320.100 160.050 321.900 161.850 ;
        RECT 322.950 158.850 325.050 160.950 ;
        RECT 326.250 160.050 328.050 161.850 ;
        RECT 323.100 157.050 324.900 158.850 ;
        RECT 329.400 154.800 330.300 163.050 ;
        RECT 340.950 161.850 343.050 163.950 ;
        RECT 343.950 163.050 346.050 165.150 ;
        RECT 323.700 153.900 330.300 154.800 ;
        RECT 323.700 153.600 325.200 153.900 ;
        RECT 305.400 147.600 307.200 153.600 ;
        RECT 313.800 147.600 315.600 153.600 ;
        RECT 323.400 147.600 325.200 153.600 ;
        RECT 329.400 153.600 330.300 153.900 ;
        RECT 341.400 153.600 342.600 161.850 ;
        RECT 329.400 147.600 331.200 153.600 ;
        RECT 340.800 147.600 342.600 153.600 ;
        RECT 350.400 153.600 351.600 166.050 ;
        RECT 359.550 156.450 360.450 167.550 ;
        RECT 361.950 166.950 364.050 167.550 ;
        RECT 364.950 166.950 366.150 170.250 ;
        RECT 368.100 168.150 369.900 169.950 ;
        RECT 380.250 168.150 382.050 169.950 ;
        RECT 364.950 164.850 367.050 166.950 ;
        RECT 367.950 166.050 370.050 168.150 ;
        RECT 370.950 164.850 373.050 166.950 ;
        RECT 376.950 164.850 379.050 166.950 ;
        RECT 379.950 166.050 382.050 168.150 ;
        RECT 384.000 166.950 385.050 173.400 ;
        RECT 392.400 171.900 394.200 179.400 ;
        RECT 399.900 174.900 401.700 179.400 ;
        RECT 412.800 176.400 414.600 179.400 ;
        RECT 399.900 173.400 403.050 174.900 ;
        RECT 398.100 171.900 399.900 172.500 ;
        RECT 392.400 170.700 399.900 171.900 ;
        RECT 382.950 164.850 385.050 166.950 ;
        RECT 385.950 168.150 387.750 169.950 ;
        RECT 385.950 166.050 388.050 168.150 ;
        RECT 388.950 164.850 391.050 166.950 ;
        RECT 391.950 164.850 394.050 166.950 ;
        RECT 361.950 161.850 364.050 163.950 ;
        RECT 362.250 160.050 364.050 161.850 ;
        RECT 365.850 159.600 367.050 164.850 ;
        RECT 371.100 163.050 372.900 164.850 ;
        RECT 377.100 163.050 378.900 164.850 ;
        RECT 382.950 161.400 383.850 164.850 ;
        RECT 388.950 163.050 390.750 164.850 ;
        RECT 392.100 163.050 393.900 164.850 ;
        RECT 379.800 160.500 383.850 161.400 ;
        RECT 361.950 156.450 364.050 157.050 ;
        RECT 359.550 155.550 364.050 156.450 ;
        RECT 361.950 154.950 364.050 155.550 ;
        RECT 350.400 147.600 352.200 153.600 ;
        RECT 365.700 147.600 367.500 159.600 ;
        RECT 376.800 148.500 378.600 159.600 ;
        RECT 379.800 149.400 381.600 160.500 ;
        RECT 382.800 158.400 390.600 159.300 ;
        RECT 382.800 148.500 384.600 158.400 ;
        RECT 376.800 147.600 384.600 148.500 ;
        RECT 388.800 147.600 390.600 158.400 ;
        RECT 395.550 153.600 396.600 170.700 ;
        RECT 402.000 166.950 403.050 173.400 ;
        RECT 413.400 168.150 414.600 176.400 ;
        RECT 422.400 174.300 424.200 179.400 ;
        RECT 428.400 174.300 430.200 179.400 ;
        RECT 422.400 172.950 430.200 174.300 ;
        RECT 431.400 173.400 433.200 179.400 ;
        RECT 431.400 171.300 432.600 173.400 ;
        RECT 441.000 172.200 442.800 179.400 ;
        RECT 455.400 176.400 457.200 179.400 ;
        RECT 441.000 171.300 444.600 172.200 ;
        RECT 428.850 170.250 432.600 171.300 ;
        RECT 398.100 165.150 399.900 166.950 ;
        RECT 397.950 163.050 400.050 165.150 ;
        RECT 400.950 164.850 403.050 166.950 ;
        RECT 412.950 166.050 415.050 168.150 ;
        RECT 415.950 167.850 418.050 169.950 ;
        RECT 425.100 168.150 426.900 169.950 ;
        RECT 416.100 166.050 417.900 167.850 ;
        RECT 402.000 159.600 403.050 164.850 ;
        RECT 395.400 147.600 397.200 153.600 ;
        RECT 402.000 147.600 403.800 159.600 ;
        RECT 413.400 153.600 414.600 166.050 ;
        RECT 421.950 164.850 424.050 166.950 ;
        RECT 424.950 166.050 427.050 168.150 ;
        RECT 428.850 166.950 430.050 170.250 ;
        RECT 427.950 164.850 430.050 166.950 ;
        RECT 440.100 165.150 441.900 166.950 ;
        RECT 422.100 163.050 423.900 164.850 ;
        RECT 427.950 159.600 429.150 164.850 ;
        RECT 430.950 161.850 433.050 163.950 ;
        RECT 439.950 163.050 442.050 165.150 ;
        RECT 443.400 163.950 444.600 171.300 ;
        RECT 456.000 169.950 457.050 176.400 ;
        RECT 469.200 172.200 471.000 179.400 ;
        RECT 454.950 167.850 457.050 169.950 ;
        RECT 446.100 165.150 447.900 166.950 ;
        RECT 442.950 161.850 445.050 163.950 ;
        RECT 445.950 163.050 448.050 165.150 ;
        RECT 451.950 164.850 454.050 166.950 ;
        RECT 452.100 163.050 453.900 164.850 ;
        RECT 430.950 160.050 432.750 161.850 ;
        RECT 412.800 147.600 414.600 153.600 ;
        RECT 427.500 147.600 429.300 159.600 ;
        RECT 443.400 153.600 444.600 161.850 ;
        RECT 456.000 160.650 457.050 167.850 ;
        RECT 467.400 171.300 471.000 172.200 ;
        RECT 486.000 173.400 487.800 179.400 ;
        RECT 457.950 164.850 460.050 166.950 ;
        RECT 464.100 165.150 465.900 166.950 ;
        RECT 458.100 163.050 459.900 164.850 ;
        RECT 463.950 163.050 466.050 165.150 ;
        RECT 467.400 163.950 468.600 171.300 ;
        RECT 482.250 168.150 484.050 169.950 ;
        RECT 470.100 165.150 471.900 166.950 ;
        RECT 466.950 161.850 469.050 163.950 ;
        RECT 469.950 163.050 472.050 165.150 ;
        RECT 478.950 164.850 481.050 166.950 ;
        RECT 481.950 166.050 484.050 168.150 ;
        RECT 486.000 166.950 487.050 173.400 ;
        RECT 500.100 171.000 501.900 179.400 ;
        RECT 515.400 176.400 517.200 179.400 ;
        RECT 484.950 164.850 487.050 166.950 ;
        RECT 487.950 168.150 489.750 169.950 ;
        RECT 500.100 169.350 504.300 171.000 ;
        RECT 487.950 166.050 490.050 168.150 ;
        RECT 490.950 164.850 493.050 166.950 ;
        RECT 503.400 165.150 504.300 169.350 ;
        RECT 511.950 167.850 514.050 169.950 ;
        RECT 515.400 168.150 516.600 176.400 ;
        RECT 529.200 172.200 531.000 179.400 ;
        RECT 527.400 171.300 531.000 172.200 ;
        RECT 540.000 172.200 541.800 179.400 ;
        RECT 540.000 171.300 543.600 172.200 ;
        RECT 512.100 166.050 513.900 167.850 ;
        RECT 514.950 166.050 517.050 168.150 ;
        RECT 479.100 163.050 480.900 164.850 ;
        RECT 456.000 159.600 458.400 160.650 ;
        RECT 442.800 147.600 444.600 153.600 ;
        RECT 456.600 147.600 458.400 159.600 ;
        RECT 467.400 153.600 468.600 161.850 ;
        RECT 484.950 161.400 485.850 164.850 ;
        RECT 490.950 163.050 492.750 164.850 ;
        RECT 493.950 161.850 496.050 163.950 ;
        RECT 499.950 161.850 502.050 163.950 ;
        RECT 502.950 163.050 505.050 165.150 ;
        RECT 481.800 160.500 485.850 161.400 ;
        RECT 467.400 147.600 469.200 153.600 ;
        RECT 478.800 148.500 480.600 159.600 ;
        RECT 481.800 149.400 483.600 160.500 ;
        RECT 494.100 160.050 495.900 161.850 ;
        RECT 484.800 158.400 492.600 159.300 ;
        RECT 496.950 158.850 499.050 160.950 ;
        RECT 500.250 160.050 502.050 161.850 ;
        RECT 484.800 148.500 486.600 158.400 ;
        RECT 478.800 147.600 486.600 148.500 ;
        RECT 490.800 147.600 492.600 158.400 ;
        RECT 497.100 157.050 498.900 158.850 ;
        RECT 503.400 154.800 504.300 163.050 ;
        RECT 497.700 153.900 504.300 154.800 ;
        RECT 497.700 153.600 499.200 153.900 ;
        RECT 497.400 147.600 499.200 153.600 ;
        RECT 503.400 153.600 504.300 153.900 ;
        RECT 515.400 153.600 516.600 166.050 ;
        RECT 524.100 165.150 525.900 166.950 ;
        RECT 523.950 163.050 526.050 165.150 ;
        RECT 527.400 163.950 528.600 171.300 ;
        RECT 530.100 165.150 531.900 166.950 ;
        RECT 539.100 165.150 540.900 166.950 ;
        RECT 526.950 161.850 529.050 163.950 ;
        RECT 529.950 163.050 532.050 165.150 ;
        RECT 538.950 163.050 541.050 165.150 ;
        RECT 542.400 163.950 543.600 171.300 ;
        RECT 544.950 171.450 547.050 172.050 ;
        RECT 544.950 170.550 549.450 171.450 ;
        RECT 554.100 171.000 555.900 179.400 ;
        RECT 568.800 173.400 570.600 179.400 ;
        RECT 544.950 169.950 547.050 170.550 ;
        RECT 545.100 165.150 546.900 166.950 ;
        RECT 541.950 161.850 544.050 163.950 ;
        RECT 544.950 163.050 547.050 165.150 ;
        RECT 527.400 153.600 528.600 161.850 ;
        RECT 542.400 153.600 543.600 161.850 ;
        RECT 544.950 159.450 547.050 160.050 ;
        RECT 548.550 159.450 549.450 170.550 ;
        RECT 551.700 169.350 555.900 171.000 ;
        RECT 569.400 171.300 570.600 173.400 ;
        RECT 571.800 174.300 573.600 179.400 ;
        RECT 577.800 174.300 579.600 179.400 ;
        RECT 571.800 172.950 579.600 174.300 ;
        RECT 569.400 170.250 573.150 171.300 ;
        RECT 587.100 171.000 588.900 179.400 ;
        RECT 601.200 175.050 603.000 179.400 ;
        RECT 601.200 173.400 606.600 175.050 ;
        RECT 551.700 165.150 552.600 169.350 ;
        RECT 571.950 166.950 573.150 170.250 ;
        RECT 575.100 168.150 576.900 169.950 ;
        RECT 584.700 169.350 588.900 171.000 ;
        RECT 562.950 165.450 565.050 166.050 ;
        RECT 550.950 163.050 553.050 165.150 ;
        RECT 562.950 164.550 567.450 165.450 ;
        RECT 571.950 164.850 574.050 166.950 ;
        RECT 574.950 166.050 577.050 168.150 ;
        RECT 577.950 164.850 580.050 166.950 ;
        RECT 584.700 165.150 585.600 169.350 ;
        RECT 596.100 168.150 597.900 169.950 ;
        RECT 595.950 166.050 598.050 168.150 ;
        RECT 598.950 167.850 601.050 169.950 ;
        RECT 602.100 168.150 603.900 169.950 ;
        RECT 599.100 166.050 600.900 167.850 ;
        RECT 601.950 166.050 604.050 168.150 ;
        RECT 605.700 166.950 606.600 173.400 ;
        RECT 611.400 174.300 613.200 179.400 ;
        RECT 617.400 174.300 619.200 179.400 ;
        RECT 611.400 172.950 619.200 174.300 ;
        RECT 620.400 173.400 622.200 179.400 ;
        RECT 628.800 176.400 630.600 179.400 ;
        RECT 620.400 171.300 621.600 173.400 ;
        RECT 617.850 170.250 621.600 171.300 ;
        RECT 614.100 168.150 615.900 169.950 ;
        RECT 562.950 163.950 565.050 164.550 ;
        RECT 544.950 158.550 549.450 159.450 ;
        RECT 544.950 157.950 547.050 158.550 ;
        RECT 551.700 154.800 552.600 163.050 ;
        RECT 553.950 161.850 556.050 163.950 ;
        RECT 559.950 161.850 562.050 163.950 ;
        RECT 553.950 160.050 555.750 161.850 ;
        RECT 556.950 158.850 559.050 160.950 ;
        RECT 560.100 160.050 561.900 161.850 ;
        RECT 557.100 157.050 558.900 158.850 ;
        RECT 566.550 156.450 567.450 164.550 ;
        RECT 568.950 161.850 571.050 163.950 ;
        RECT 569.250 160.050 571.050 161.850 ;
        RECT 572.850 159.600 574.050 164.850 ;
        RECT 578.100 163.050 579.900 164.850 ;
        RECT 583.950 163.050 586.050 165.150 ;
        RECT 604.950 164.850 607.050 166.950 ;
        RECT 610.950 164.850 613.050 166.950 ;
        RECT 613.950 166.050 616.050 168.150 ;
        RECT 617.850 166.950 619.050 170.250 ;
        RECT 629.400 168.150 630.600 176.400 ;
        RECT 640.800 173.400 642.600 179.400 ;
        RECT 641.400 171.300 642.600 173.400 ;
        RECT 643.800 174.300 645.600 179.400 ;
        RECT 649.800 174.300 651.600 179.400 ;
        RECT 643.800 172.950 651.600 174.300 ;
        RECT 655.800 173.400 657.600 179.400 ;
        RECT 656.400 171.300 657.600 173.400 ;
        RECT 658.800 174.300 660.600 179.400 ;
        RECT 664.800 174.300 666.600 179.400 ;
        RECT 658.800 172.950 666.600 174.300 ;
        RECT 641.400 170.250 645.150 171.300 ;
        RECT 656.400 170.250 660.150 171.300 ;
        RECT 616.950 164.850 619.050 166.950 ;
        RECT 628.950 166.050 631.050 168.150 ;
        RECT 631.950 167.850 634.050 169.950 ;
        RECT 632.100 166.050 633.900 167.850 ;
        RECT 643.950 166.950 645.150 170.250 ;
        RECT 647.100 168.150 648.900 169.950 ;
        RECT 568.950 156.450 571.050 157.050 ;
        RECT 566.550 155.550 571.050 156.450 ;
        RECT 568.950 154.950 571.050 155.550 ;
        RECT 551.700 153.900 558.300 154.800 ;
        RECT 551.700 153.600 552.600 153.900 ;
        RECT 503.400 147.600 505.200 153.600 ;
        RECT 515.400 147.600 517.200 153.600 ;
        RECT 527.400 147.600 529.200 153.600 ;
        RECT 541.800 147.600 543.600 153.600 ;
        RECT 550.800 147.600 552.600 153.600 ;
        RECT 556.800 153.600 558.300 153.900 ;
        RECT 556.800 147.600 558.600 153.600 ;
        RECT 572.700 147.600 574.500 159.600 ;
        RECT 584.700 154.800 585.600 163.050 ;
        RECT 586.950 161.850 589.050 163.950 ;
        RECT 592.950 161.850 595.050 163.950 ;
        RECT 586.950 160.050 588.750 161.850 ;
        RECT 589.950 158.850 592.050 160.950 ;
        RECT 593.100 160.050 594.900 161.850 ;
        RECT 605.700 159.600 606.600 164.850 ;
        RECT 611.100 163.050 612.900 164.850 ;
        RECT 616.950 159.600 618.150 164.850 ;
        RECT 619.950 161.850 622.050 163.950 ;
        RECT 619.950 160.050 621.750 161.850 ;
        RECT 590.100 157.050 591.900 158.850 ;
        RECT 596.400 158.700 604.200 159.600 ;
        RECT 584.700 153.900 591.300 154.800 ;
        RECT 584.700 153.600 585.600 153.900 ;
        RECT 583.800 147.600 585.600 153.600 ;
        RECT 589.800 153.600 591.300 153.900 ;
        RECT 589.800 147.600 591.600 153.600 ;
        RECT 596.400 147.600 598.200 158.700 ;
        RECT 602.400 147.600 604.200 158.700 ;
        RECT 605.400 147.600 607.200 159.600 ;
        RECT 616.500 147.600 618.300 159.600 ;
        RECT 629.400 153.600 630.600 166.050 ;
        RECT 643.950 164.850 646.050 166.950 ;
        RECT 646.950 166.050 649.050 168.150 ;
        RECT 658.950 166.950 660.150 170.250 ;
        RECT 677.100 171.000 678.900 179.400 ;
        RECT 694.200 175.050 696.000 179.400 ;
        RECT 694.200 173.400 699.600 175.050 ;
        RECT 662.100 168.150 663.900 169.950 ;
        RECT 677.100 169.350 681.300 171.000 ;
        RECT 649.950 164.850 652.050 166.950 ;
        RECT 658.950 164.850 661.050 166.950 ;
        RECT 661.950 166.050 664.050 168.150 ;
        RECT 664.950 164.850 667.050 166.950 ;
        RECT 680.400 165.150 681.300 169.350 ;
        RECT 689.100 168.150 690.900 169.950 ;
        RECT 688.950 166.050 691.050 168.150 ;
        RECT 691.950 167.850 694.050 169.950 ;
        RECT 695.100 168.150 696.900 169.950 ;
        RECT 692.100 166.050 693.900 167.850 ;
        RECT 694.950 166.050 697.050 168.150 ;
        RECT 698.700 166.950 699.600 173.400 ;
        RECT 704.400 174.300 706.200 179.400 ;
        RECT 710.400 174.300 712.200 179.400 ;
        RECT 704.400 172.950 712.200 174.300 ;
        RECT 713.400 173.400 715.200 179.400 ;
        RECT 729.000 175.050 730.800 179.400 ;
        RECT 725.400 173.400 730.800 175.050 ;
        RECT 713.400 171.300 714.600 173.400 ;
        RECT 710.850 170.250 714.600 171.300 ;
        RECT 707.100 168.150 708.900 169.950 ;
        RECT 640.950 161.850 643.050 163.950 ;
        RECT 641.250 160.050 643.050 161.850 ;
        RECT 644.850 159.600 646.050 164.850 ;
        RECT 650.100 163.050 651.900 164.850 ;
        RECT 655.950 161.850 658.050 163.950 ;
        RECT 656.250 160.050 658.050 161.850 ;
        RECT 659.850 159.600 661.050 164.850 ;
        RECT 665.100 163.050 666.900 164.850 ;
        RECT 670.950 161.850 673.050 163.950 ;
        RECT 676.950 161.850 679.050 163.950 ;
        RECT 679.950 163.050 682.050 165.150 ;
        RECT 697.950 164.850 700.050 166.950 ;
        RECT 703.950 164.850 706.050 166.950 ;
        RECT 706.950 166.050 709.050 168.150 ;
        RECT 710.850 166.950 712.050 170.250 ;
        RECT 725.400 166.950 726.300 173.400 ;
        RECT 746.100 171.000 747.900 179.400 ;
        RECT 728.100 168.150 729.900 169.950 ;
        RECT 709.950 164.850 712.050 166.950 ;
        RECT 724.950 164.850 727.050 166.950 ;
        RECT 727.950 166.050 730.050 168.150 ;
        RECT 730.950 167.850 733.050 169.950 ;
        RECT 734.100 168.150 735.900 169.950 ;
        RECT 743.700 169.350 747.900 171.000 ;
        RECT 731.100 166.050 732.900 167.850 ;
        RECT 733.950 166.050 736.050 168.150 ;
        RECT 743.700 165.150 744.600 169.350 ;
        RECT 671.100 160.050 672.900 161.850 ;
        RECT 628.800 147.600 630.600 153.600 ;
        RECT 644.700 147.600 646.500 159.600 ;
        RECT 659.700 147.600 661.500 159.600 ;
        RECT 673.950 158.850 676.050 160.950 ;
        RECT 677.250 160.050 679.050 161.850 ;
        RECT 674.100 157.050 675.900 158.850 ;
        RECT 680.400 154.800 681.300 163.050 ;
        RECT 698.700 159.600 699.600 164.850 ;
        RECT 704.100 163.050 705.900 164.850 ;
        RECT 709.950 159.600 711.150 164.850 ;
        RECT 712.950 161.850 715.050 163.950 ;
        RECT 712.950 160.050 714.750 161.850 ;
        RECT 725.400 159.600 726.300 164.850 ;
        RECT 742.950 163.050 745.050 165.150 ;
        RECT 674.700 153.900 681.300 154.800 ;
        RECT 674.700 153.600 676.200 153.900 ;
        RECT 674.400 147.600 676.200 153.600 ;
        RECT 680.400 153.600 681.300 153.900 ;
        RECT 689.400 158.700 697.200 159.600 ;
        RECT 680.400 147.600 682.200 153.600 ;
        RECT 689.400 147.600 691.200 158.700 ;
        RECT 695.400 147.600 697.200 158.700 ;
        RECT 698.400 147.600 700.200 159.600 ;
        RECT 709.500 147.600 711.300 159.600 ;
        RECT 724.800 147.600 726.600 159.600 ;
        RECT 727.800 158.700 735.600 159.600 ;
        RECT 727.800 147.600 729.600 158.700 ;
        RECT 733.800 147.600 735.600 158.700 ;
        RECT 743.700 154.800 744.600 163.050 ;
        RECT 745.950 161.850 748.050 163.950 ;
        RECT 751.950 161.850 754.050 163.950 ;
        RECT 745.950 160.050 747.750 161.850 ;
        RECT 748.950 158.850 751.050 160.950 ;
        RECT 752.100 160.050 753.900 161.850 ;
        RECT 749.100 157.050 750.900 158.850 ;
        RECT 743.700 153.900 750.300 154.800 ;
        RECT 743.700 153.600 744.600 153.900 ;
        RECT 742.800 147.600 744.600 153.600 ;
        RECT 748.800 153.600 750.300 153.900 ;
        RECT 748.800 147.600 750.600 153.600 ;
        RECT 4.800 137.400 6.600 143.400 ;
        RECT 13.800 137.400 15.600 143.400 ;
        RECT 22.800 137.400 24.600 143.400 ;
        RECT 5.400 124.950 6.600 137.400 ;
        RECT 14.400 124.950 15.600 137.400 ;
        RECT 23.700 137.100 24.600 137.400 ;
        RECT 28.800 137.400 30.600 143.400 ;
        RECT 28.800 137.100 30.300 137.400 ;
        RECT 23.700 136.200 30.300 137.100 ;
        RECT 23.700 127.950 24.600 136.200 ;
        RECT 29.100 132.150 30.900 133.950 ;
        RECT 38.400 132.300 40.200 143.400 ;
        RECT 44.400 132.300 46.200 143.400 ;
        RECT 25.950 129.150 27.750 130.950 ;
        RECT 28.950 130.050 31.050 132.150 ;
        RECT 38.400 131.400 46.200 132.300 ;
        RECT 47.400 131.400 49.200 143.400 ;
        RECT 58.800 137.400 60.600 143.400 ;
        RECT 32.100 129.150 33.900 130.950 ;
        RECT 22.950 125.850 25.050 127.950 ;
        RECT 25.950 127.050 28.050 129.150 ;
        RECT 31.950 127.050 34.050 129.150 ;
        RECT 47.700 126.150 48.600 131.400 ;
        RECT 59.400 129.150 60.600 137.400 ;
        RECT 71.700 131.400 73.500 143.400 ;
        RECT 84.600 131.400 86.400 143.400 ;
        RECT 94.800 137.400 96.600 143.400 ;
        RECT 68.250 129.150 70.050 130.950 ;
        RECT 4.950 122.850 7.050 124.950 ;
        RECT 8.100 123.150 9.900 124.950 ;
        RECT 5.400 114.600 6.600 122.850 ;
        RECT 7.950 121.050 10.050 123.150 ;
        RECT 13.950 122.850 16.050 124.950 ;
        RECT 17.100 123.150 18.900 124.950 ;
        RECT 14.400 114.600 15.600 122.850 ;
        RECT 16.950 121.050 19.050 123.150 ;
        RECT 23.700 121.650 24.600 125.850 ;
        RECT 37.950 122.850 40.050 124.950 ;
        RECT 41.100 123.150 42.900 124.950 ;
        RECT 23.700 120.000 27.900 121.650 ;
        RECT 38.100 121.050 39.900 122.850 ;
        RECT 40.950 121.050 43.050 123.150 ;
        RECT 43.950 122.850 46.050 124.950 ;
        RECT 46.950 124.050 49.050 126.150 ;
        RECT 55.950 125.850 58.050 127.950 ;
        RECT 58.950 127.050 61.050 129.150 ;
        RECT 56.100 124.050 57.900 125.850 ;
        RECT 44.100 121.050 45.900 122.850 ;
        RECT 4.800 111.600 6.600 114.600 ;
        RECT 13.800 111.600 15.600 114.600 ;
        RECT 26.100 111.600 27.900 120.000 ;
        RECT 47.700 117.600 48.600 124.050 ;
        RECT 59.400 119.700 60.600 127.050 ;
        RECT 61.950 125.850 64.050 127.950 ;
        RECT 67.950 127.050 70.050 129.150 ;
        RECT 71.850 126.150 73.050 131.400 ;
        RECT 84.000 130.350 86.400 131.400 ;
        RECT 95.700 137.100 96.600 137.400 ;
        RECT 100.800 137.400 102.600 143.400 ;
        RECT 112.800 137.400 114.600 143.400 ;
        RECT 124.800 137.400 126.600 143.400 ;
        RECT 100.800 137.100 102.300 137.400 ;
        RECT 95.700 136.200 102.300 137.100 ;
        RECT 77.100 126.150 78.900 127.950 ;
        RECT 80.100 126.150 81.900 127.950 ;
        RECT 62.100 124.050 63.900 125.850 ;
        RECT 70.950 124.050 73.050 126.150 ;
        RECT 70.950 120.750 72.150 124.050 ;
        RECT 73.950 122.850 76.050 124.950 ;
        RECT 76.950 124.050 79.050 126.150 ;
        RECT 79.950 124.050 82.050 126.150 ;
        RECT 84.000 123.150 85.050 130.350 ;
        RECT 95.700 127.950 96.600 136.200 ;
        RECT 101.100 132.150 102.900 133.950 ;
        RECT 97.950 129.150 99.750 130.950 ;
        RECT 100.950 130.050 103.050 132.150 ;
        RECT 104.100 129.150 105.900 130.950 ;
        RECT 113.400 129.150 114.600 137.400 ;
        RECT 125.400 129.150 126.600 137.400 ;
        RECT 133.800 131.400 135.600 143.400 ;
        RECT 145.800 137.400 147.600 143.400 ;
        RECT 160.800 137.400 162.600 143.400 ;
        RECT 175.800 137.400 177.600 143.400 ;
        RECT 86.100 126.150 87.900 127.950 ;
        RECT 85.950 124.050 88.050 126.150 ;
        RECT 94.950 125.850 97.050 127.950 ;
        RECT 97.950 127.050 100.050 129.150 ;
        RECT 103.950 127.050 106.050 129.150 ;
        RECT 109.950 125.850 112.050 127.950 ;
        RECT 112.950 127.050 115.050 129.150 ;
        RECT 74.100 121.050 75.900 122.850 ;
        RECT 82.950 121.050 85.050 123.150 ;
        RECT 43.200 115.950 48.600 117.600 ;
        RECT 57.000 118.800 60.600 119.700 ;
        RECT 68.400 119.700 72.150 120.750 ;
        RECT 43.200 111.600 45.000 115.950 ;
        RECT 57.000 111.600 58.800 118.800 ;
        RECT 68.400 117.600 69.600 119.700 ;
        RECT 67.800 111.600 69.600 117.600 ;
        RECT 70.800 116.700 78.600 118.050 ;
        RECT 70.800 111.600 72.600 116.700 ;
        RECT 76.800 111.600 78.600 116.700 ;
        RECT 84.000 114.600 85.050 121.050 ;
        RECT 95.700 121.650 96.600 125.850 ;
        RECT 110.100 124.050 111.900 125.850 ;
        RECT 95.700 120.000 99.900 121.650 ;
        RECT 83.400 111.600 85.200 114.600 ;
        RECT 98.100 111.600 99.900 120.000 ;
        RECT 113.400 119.700 114.600 127.050 ;
        RECT 115.950 125.850 118.050 127.950 ;
        RECT 121.950 125.850 124.050 127.950 ;
        RECT 124.950 127.050 127.050 129.150 ;
        RECT 116.100 124.050 117.900 125.850 ;
        RECT 122.100 124.050 123.900 125.850 ;
        RECT 125.400 119.700 126.600 127.050 ;
        RECT 127.950 125.850 130.050 127.950 ;
        RECT 134.400 126.150 135.600 131.400 ;
        RECT 146.400 129.150 147.600 137.400 ;
        RECT 161.400 129.150 162.600 137.400 ;
        RECT 176.400 129.150 177.600 137.400 ;
        RECT 188.700 131.400 190.500 143.400 ;
        RECT 202.200 131.400 204.000 143.400 ;
        RECT 208.800 137.400 210.600 143.400 ;
        RECT 220.800 137.400 222.600 143.400 ;
        RECT 229.800 137.400 231.600 143.400 ;
        RECT 185.250 129.150 187.050 130.950 ;
        RECT 128.100 124.050 129.900 125.850 ;
        RECT 133.950 124.050 136.050 126.150 ;
        RECT 142.950 125.850 145.050 127.950 ;
        RECT 145.950 127.050 148.050 129.150 ;
        RECT 111.000 118.800 114.600 119.700 ;
        RECT 123.000 118.800 126.600 119.700 ;
        RECT 111.000 111.600 112.800 118.800 ;
        RECT 123.000 111.600 124.800 118.800 ;
        RECT 134.400 117.600 135.600 124.050 ;
        RECT 136.950 122.850 139.050 124.950 ;
        RECT 143.100 124.050 144.900 125.850 ;
        RECT 137.100 121.050 138.900 122.850 ;
        RECT 146.400 119.700 147.600 127.050 ;
        RECT 148.950 125.850 151.050 127.950 ;
        RECT 157.950 125.850 160.050 127.950 ;
        RECT 160.950 127.050 163.050 129.150 ;
        RECT 149.100 124.050 150.900 125.850 ;
        RECT 158.100 124.050 159.900 125.850 ;
        RECT 161.400 119.700 162.600 127.050 ;
        RECT 163.950 125.850 166.050 127.950 ;
        RECT 172.950 125.850 175.050 127.950 ;
        RECT 175.950 127.050 178.050 129.150 ;
        RECT 164.100 124.050 165.900 125.850 ;
        RECT 173.100 124.050 174.900 125.850 ;
        RECT 176.400 119.700 177.600 127.050 ;
        RECT 178.950 125.850 181.050 127.950 ;
        RECT 184.950 127.050 187.050 129.150 ;
        RECT 188.850 126.150 190.050 131.400 ;
        RECT 194.100 126.150 195.900 127.950 ;
        RECT 202.950 126.150 204.000 131.400 ;
        RECT 179.100 124.050 180.900 125.850 ;
        RECT 187.950 124.050 190.050 126.150 ;
        RECT 187.950 120.750 189.150 124.050 ;
        RECT 190.950 122.850 193.050 124.950 ;
        RECT 193.950 124.050 196.050 126.150 ;
        RECT 202.950 124.050 205.050 126.150 ;
        RECT 205.950 125.850 208.050 127.950 ;
        RECT 206.100 124.050 207.900 125.850 ;
        RECT 191.100 121.050 192.900 122.850 ;
        RECT 133.800 111.600 135.600 117.600 ;
        RECT 144.000 118.800 147.600 119.700 ;
        RECT 159.000 118.800 162.600 119.700 ;
        RECT 174.000 118.800 177.600 119.700 ;
        RECT 185.400 119.700 189.150 120.750 ;
        RECT 144.000 111.600 145.800 118.800 ;
        RECT 159.000 111.600 160.800 118.800 ;
        RECT 174.000 111.600 175.800 118.800 ;
        RECT 185.400 117.600 186.600 119.700 ;
        RECT 184.800 111.600 186.600 117.600 ;
        RECT 187.800 116.700 195.600 118.050 ;
        RECT 187.800 111.600 189.600 116.700 ;
        RECT 193.800 111.600 195.600 116.700 ;
        RECT 202.950 117.600 204.000 124.050 ;
        RECT 209.400 120.300 210.450 137.400 ;
        RECT 221.400 129.150 222.600 137.400 ;
        RECT 212.100 126.150 213.900 127.950 ;
        RECT 211.950 124.050 214.050 126.150 ;
        RECT 217.950 125.850 220.050 127.950 ;
        RECT 220.950 127.050 223.050 129.150 ;
        RECT 218.100 124.050 219.900 125.850 ;
        RECT 206.100 119.100 213.600 120.300 ;
        RECT 221.400 119.700 222.600 127.050 ;
        RECT 223.950 125.850 226.050 127.950 ;
        RECT 224.100 124.050 225.900 125.850 ;
        RECT 230.400 124.950 231.600 137.400 ;
        RECT 244.800 131.400 248.100 143.400 ;
        RECT 259.800 137.400 261.600 143.400 ;
        RECT 239.250 126.150 241.050 127.950 ;
        RECT 245.400 126.150 246.600 131.400 ;
        RECT 260.400 129.150 261.600 137.400 ;
        RECT 269.400 132.300 271.200 143.400 ;
        RECT 275.400 132.300 277.200 143.400 ;
        RECT 269.400 131.400 277.200 132.300 ;
        RECT 278.400 131.400 280.200 143.400 ;
        RECT 290.700 131.400 292.500 143.400 ;
        RECT 303.600 131.400 305.400 143.400 ;
        RECT 316.800 137.400 318.600 143.400 ;
        RECT 251.100 126.150 252.900 127.950 ;
        RECT 229.950 122.850 232.050 124.950 ;
        RECT 233.100 123.150 234.900 124.950 ;
        RECT 238.950 124.050 241.050 126.150 ;
        RECT 206.100 118.500 207.900 119.100 ;
        RECT 202.950 116.100 206.100 117.600 ;
        RECT 204.300 111.600 206.100 116.100 ;
        RECT 211.800 111.600 213.600 119.100 ;
        RECT 219.000 118.800 222.600 119.700 ;
        RECT 219.000 111.600 220.800 118.800 ;
        RECT 230.400 114.600 231.600 122.850 ;
        RECT 232.950 121.050 235.050 123.150 ;
        RECT 241.950 122.850 244.050 124.950 ;
        RECT 244.950 124.050 247.050 126.150 ;
        RECT 242.700 121.050 244.500 122.850 ;
        RECT 245.400 120.150 246.600 124.050 ;
        RECT 247.950 122.850 250.050 124.950 ;
        RECT 250.950 124.050 253.050 126.150 ;
        RECT 256.950 125.850 259.050 127.950 ;
        RECT 259.950 127.050 262.050 129.150 ;
        RECT 257.100 124.050 258.900 125.850 ;
        RECT 248.100 121.050 249.900 122.850 ;
        RECT 242.400 119.100 246.600 120.150 ;
        RECT 260.400 119.700 261.600 127.050 ;
        RECT 262.950 125.850 265.050 127.950 ;
        RECT 278.700 126.150 279.600 131.400 ;
        RECT 287.250 129.150 289.050 130.950 ;
        RECT 286.950 127.050 289.050 129.150 ;
        RECT 290.850 126.150 292.050 131.400 ;
        RECT 303.000 130.350 305.400 131.400 ;
        RECT 296.100 126.150 297.900 127.950 ;
        RECT 299.100 126.150 300.900 127.950 ;
        RECT 263.100 124.050 264.900 125.850 ;
        RECT 268.950 122.850 271.050 124.950 ;
        RECT 272.100 123.150 273.900 124.950 ;
        RECT 269.100 121.050 270.900 122.850 ;
        RECT 271.950 121.050 274.050 123.150 ;
        RECT 274.950 122.850 277.050 124.950 ;
        RECT 277.950 124.050 280.050 126.150 ;
        RECT 289.950 124.050 292.050 126.150 ;
        RECT 275.100 121.050 276.900 122.850 ;
        RECT 242.400 117.600 243.300 119.100 ;
        RECT 258.000 118.800 261.600 119.700 ;
        RECT 229.800 111.600 231.600 114.600 ;
        RECT 238.800 112.500 240.600 117.600 ;
        RECT 241.800 113.400 243.600 117.600 ;
        RECT 244.800 117.000 252.600 117.900 ;
        RECT 244.800 112.500 246.600 117.000 ;
        RECT 238.800 111.600 246.600 112.500 ;
        RECT 250.800 111.600 252.600 117.000 ;
        RECT 258.000 111.600 259.800 118.800 ;
        RECT 278.700 117.600 279.600 124.050 ;
        RECT 289.950 120.750 291.150 124.050 ;
        RECT 292.950 122.850 295.050 124.950 ;
        RECT 295.950 124.050 298.050 126.150 ;
        RECT 298.950 124.050 301.050 126.150 ;
        RECT 303.000 123.150 304.050 130.350 ;
        RECT 317.400 129.150 318.600 137.400 ;
        RECT 326.400 137.400 328.200 143.400 ;
        RECT 326.400 129.150 327.600 137.400 ;
        RECT 328.950 135.450 331.050 136.050 ;
        RECT 337.950 135.450 340.050 136.050 ;
        RECT 328.950 134.550 340.050 135.450 ;
        RECT 328.950 133.950 331.050 134.550 ;
        RECT 337.950 133.950 340.050 134.550 ;
        RECT 331.950 130.950 334.050 133.050 ;
        RECT 342.600 131.400 344.400 143.400 ;
        RECT 353.400 137.400 355.200 143.400 ;
        RECT 367.800 137.400 369.600 143.400 ;
        RECT 305.100 126.150 306.900 127.950 ;
        RECT 304.950 124.050 307.050 126.150 ;
        RECT 313.950 125.850 316.050 127.950 ;
        RECT 316.950 127.050 319.050 129.150 ;
        RECT 314.100 124.050 315.900 125.850 ;
        RECT 293.100 121.050 294.900 122.850 ;
        RECT 301.950 121.050 304.050 123.150 ;
        RECT 287.400 119.700 291.150 120.750 ;
        RECT 287.400 117.600 288.600 119.700 ;
        RECT 274.200 115.950 279.600 117.600 ;
        RECT 274.200 111.600 276.000 115.950 ;
        RECT 286.800 111.600 288.600 117.600 ;
        RECT 289.800 116.700 297.600 118.050 ;
        RECT 289.800 111.600 291.600 116.700 ;
        RECT 295.800 111.600 297.600 116.700 ;
        RECT 303.000 114.600 304.050 121.050 ;
        RECT 317.400 119.700 318.600 127.050 ;
        RECT 319.950 125.850 322.050 127.950 ;
        RECT 322.950 125.850 325.050 127.950 ;
        RECT 325.950 127.050 328.050 129.150 ;
        RECT 320.100 124.050 321.900 125.850 ;
        RECT 323.100 124.050 324.900 125.850 ;
        RECT 315.000 118.800 318.600 119.700 ;
        RECT 326.400 119.700 327.600 127.050 ;
        RECT 328.950 125.850 331.050 127.950 ;
        RECT 329.100 124.050 330.900 125.850 ;
        RECT 326.400 118.800 330.000 119.700 ;
        RECT 302.400 111.600 304.200 114.600 ;
        RECT 315.000 111.600 316.800 118.800 ;
        RECT 328.200 111.600 330.000 118.800 ;
        RECT 332.550 118.050 333.450 130.950 ;
        RECT 342.600 130.350 345.000 131.400 ;
        RECT 341.100 126.150 342.900 127.950 ;
        RECT 340.950 124.050 343.050 126.150 ;
        RECT 343.950 123.150 345.000 130.350 ;
        RECT 353.400 129.150 354.600 137.400 ;
        RECT 368.400 129.150 369.600 137.400 ;
        RECT 377.400 137.400 379.200 143.400 ;
        RECT 377.400 129.150 378.600 137.400 ;
        RECT 388.800 131.400 390.600 143.400 ;
        RECT 391.800 132.300 393.600 143.400 ;
        RECT 397.800 132.300 399.600 143.400 ;
        RECT 404.400 137.400 406.200 143.400 ;
        RECT 404.700 137.100 406.200 137.400 ;
        RECT 410.400 137.400 412.200 143.400 ;
        RECT 421.800 137.400 423.600 143.400 ;
        RECT 410.400 137.100 411.300 137.400 ;
        RECT 404.700 136.200 411.300 137.100 ;
        RECT 391.800 131.400 399.600 132.300 ;
        RECT 404.100 132.150 405.900 133.950 ;
        RECT 347.100 126.150 348.900 127.950 ;
        RECT 346.950 124.050 349.050 126.150 ;
        RECT 349.950 125.850 352.050 127.950 ;
        RECT 352.950 127.050 355.050 129.150 ;
        RECT 350.100 124.050 351.900 125.850 ;
        RECT 343.950 121.050 346.050 123.150 ;
        RECT 331.950 115.950 334.050 118.050 ;
        RECT 343.950 114.600 345.000 121.050 ;
        RECT 353.400 119.700 354.600 127.050 ;
        RECT 355.950 125.850 358.050 127.950 ;
        RECT 364.950 125.850 367.050 127.950 ;
        RECT 367.950 127.050 370.050 129.150 ;
        RECT 356.100 124.050 357.900 125.850 ;
        RECT 365.100 124.050 366.900 125.850 ;
        RECT 368.400 119.700 369.600 127.050 ;
        RECT 370.950 125.850 373.050 127.950 ;
        RECT 373.950 125.850 376.050 127.950 ;
        RECT 376.950 127.050 379.050 129.150 ;
        RECT 371.100 124.050 372.900 125.850 ;
        RECT 374.100 124.050 375.900 125.850 ;
        RECT 353.400 118.800 357.000 119.700 ;
        RECT 343.800 111.600 345.600 114.600 ;
        RECT 355.200 111.600 357.000 118.800 ;
        RECT 366.000 118.800 369.600 119.700 ;
        RECT 377.400 119.700 378.600 127.050 ;
        RECT 379.950 125.850 382.050 127.950 ;
        RECT 389.400 126.150 390.300 131.400 ;
        RECT 401.100 129.150 402.900 130.950 ;
        RECT 403.950 130.050 406.050 132.150 ;
        RECT 407.250 129.150 409.050 130.950 ;
        RECT 400.950 127.050 403.050 129.150 ;
        RECT 406.950 127.050 409.050 129.150 ;
        RECT 410.400 127.950 411.300 136.200 ;
        RECT 422.700 137.100 423.600 137.400 ;
        RECT 427.800 137.400 429.600 143.400 ;
        RECT 427.800 137.100 429.300 137.400 ;
        RECT 422.700 136.200 429.300 137.100 ;
        RECT 422.700 127.950 423.600 136.200 ;
        RECT 428.100 132.150 429.900 133.950 ;
        RECT 424.950 129.150 426.750 130.950 ;
        RECT 427.950 130.050 430.050 132.150 ;
        RECT 443.700 131.400 445.500 143.400 ;
        RECT 454.800 131.400 456.600 143.400 ;
        RECT 457.800 132.300 459.600 143.400 ;
        RECT 463.800 132.300 465.600 143.400 ;
        RECT 457.800 131.400 465.600 132.300 ;
        RECT 472.800 131.400 474.600 143.400 ;
        RECT 475.800 132.300 477.600 143.400 ;
        RECT 481.800 132.300 483.600 143.400 ;
        RECT 490.800 137.400 492.600 143.400 ;
        RECT 475.800 131.400 483.600 132.300 ;
        RECT 431.100 129.150 432.900 130.950 ;
        RECT 380.100 124.050 381.900 125.850 ;
        RECT 388.950 124.050 391.050 126.150 ;
        RECT 409.950 125.850 412.050 127.950 ;
        RECT 421.950 125.850 424.050 127.950 ;
        RECT 424.950 127.050 427.050 129.150 ;
        RECT 430.950 127.050 433.050 129.150 ;
        RECT 433.950 127.950 436.050 130.050 ;
        RECT 440.250 129.150 442.050 130.950 ;
        RECT 377.400 118.800 381.000 119.700 ;
        RECT 366.000 111.600 367.800 118.800 ;
        RECT 379.200 111.600 381.000 118.800 ;
        RECT 389.400 117.600 390.300 124.050 ;
        RECT 391.950 122.850 394.050 124.950 ;
        RECT 395.100 123.150 396.900 124.950 ;
        RECT 392.100 121.050 393.900 122.850 ;
        RECT 394.950 121.050 397.050 123.150 ;
        RECT 397.950 122.850 400.050 124.950 ;
        RECT 398.100 121.050 399.900 122.850 ;
        RECT 410.400 121.650 411.300 125.850 ;
        RECT 407.100 120.000 411.300 121.650 ;
        RECT 422.700 121.650 423.600 125.850 ;
        RECT 430.950 123.450 433.050 124.050 ;
        RECT 434.550 123.450 435.450 127.950 ;
        RECT 439.950 127.050 442.050 129.150 ;
        RECT 443.850 126.150 445.050 131.400 ;
        RECT 449.100 126.150 450.900 127.950 ;
        RECT 455.400 126.150 456.300 131.400 ;
        RECT 473.400 126.150 474.300 131.400 ;
        RECT 491.400 129.150 492.600 137.400 ;
        RECT 500.400 137.400 502.200 143.400 ;
        RECT 430.950 122.550 435.450 123.450 ;
        RECT 442.950 124.050 445.050 126.150 ;
        RECT 430.950 121.950 433.050 122.550 ;
        RECT 422.700 120.000 426.900 121.650 ;
        RECT 442.950 120.750 444.150 124.050 ;
        RECT 445.950 122.850 448.050 124.950 ;
        RECT 448.950 124.050 451.050 126.150 ;
        RECT 454.950 124.050 457.050 126.150 ;
        RECT 446.100 121.050 447.900 122.850 ;
        RECT 389.400 115.950 394.800 117.600 ;
        RECT 393.000 111.600 394.800 115.950 ;
        RECT 407.100 111.600 408.900 120.000 ;
        RECT 425.100 111.600 426.900 120.000 ;
        RECT 440.400 119.700 444.150 120.750 ;
        RECT 440.400 117.600 441.600 119.700 ;
        RECT 439.800 111.600 441.600 117.600 ;
        RECT 442.800 116.700 450.600 118.050 ;
        RECT 442.800 111.600 444.600 116.700 ;
        RECT 448.800 111.600 450.600 116.700 ;
        RECT 455.400 117.600 456.300 124.050 ;
        RECT 457.950 122.850 460.050 124.950 ;
        RECT 461.100 123.150 462.900 124.950 ;
        RECT 458.100 121.050 459.900 122.850 ;
        RECT 460.950 121.050 463.050 123.150 ;
        RECT 463.950 122.850 466.050 124.950 ;
        RECT 472.950 124.050 475.050 126.150 ;
        RECT 487.950 125.850 490.050 127.950 ;
        RECT 490.950 127.050 493.050 129.150 ;
        RECT 464.100 121.050 465.900 122.850 ;
        RECT 473.400 117.600 474.300 124.050 ;
        RECT 475.950 122.850 478.050 124.950 ;
        RECT 479.100 123.150 480.900 124.950 ;
        RECT 476.100 121.050 477.900 122.850 ;
        RECT 478.950 121.050 481.050 123.150 ;
        RECT 481.950 122.850 484.050 124.950 ;
        RECT 488.100 124.050 489.900 125.850 ;
        RECT 482.100 121.050 483.900 122.850 ;
        RECT 491.400 119.700 492.600 127.050 ;
        RECT 493.950 125.850 496.050 127.950 ;
        RECT 494.100 124.050 495.900 125.850 ;
        RECT 500.400 124.950 501.600 137.400 ;
        RECT 512.700 131.400 514.500 143.400 ;
        RECT 527.700 131.400 529.500 143.400 ;
        RECT 541.500 131.400 543.300 143.400 ;
        RECT 554.400 137.400 556.200 143.400 ;
        RECT 554.700 137.100 556.200 137.400 ;
        RECT 560.400 137.400 562.200 143.400 ;
        RECT 572.400 137.400 574.200 143.400 ;
        RECT 560.400 137.100 561.300 137.400 ;
        RECT 554.700 136.200 561.300 137.100 ;
        RECT 572.700 137.100 574.200 137.400 ;
        RECT 578.400 137.400 580.200 143.400 ;
        RECT 586.800 142.500 594.600 143.400 ;
        RECT 578.400 137.100 579.300 137.400 ;
        RECT 572.700 136.200 579.300 137.100 ;
        RECT 544.950 135.450 547.050 136.050 ;
        RECT 544.950 134.550 549.450 135.450 ;
        RECT 544.950 133.950 547.050 134.550 ;
        RECT 509.250 129.150 511.050 130.950 ;
        RECT 508.950 127.050 511.050 129.150 ;
        RECT 512.850 126.150 514.050 131.400 ;
        RECT 524.250 129.150 526.050 130.950 ;
        RECT 518.100 126.150 519.900 127.950 ;
        RECT 523.950 127.050 526.050 129.150 ;
        RECT 527.850 126.150 529.050 131.400 ;
        RECT 533.100 126.150 534.900 127.950 ;
        RECT 536.100 126.150 537.900 127.950 ;
        RECT 541.950 126.150 543.150 131.400 ;
        RECT 544.950 129.150 546.750 130.950 ;
        RECT 544.950 127.050 547.050 129.150 ;
        RECT 497.100 123.150 498.900 124.950 ;
        RECT 496.950 121.050 499.050 123.150 ;
        RECT 499.950 122.850 502.050 124.950 ;
        RECT 511.950 124.050 514.050 126.150 ;
        RECT 489.000 118.800 492.600 119.700 ;
        RECT 455.400 115.950 460.800 117.600 ;
        RECT 473.400 115.950 478.800 117.600 ;
        RECT 459.000 111.600 460.800 115.950 ;
        RECT 477.000 111.600 478.800 115.950 ;
        RECT 489.000 111.600 490.800 118.800 ;
        RECT 500.400 114.600 501.600 122.850 ;
        RECT 511.950 120.750 513.150 124.050 ;
        RECT 514.950 122.850 517.050 124.950 ;
        RECT 517.950 124.050 520.050 126.150 ;
        RECT 526.950 124.050 529.050 126.150 ;
        RECT 515.100 121.050 516.900 122.850 ;
        RECT 526.950 120.750 528.150 124.050 ;
        RECT 529.950 122.850 532.050 124.950 ;
        RECT 532.950 124.050 535.050 126.150 ;
        RECT 535.950 124.050 538.050 126.150 ;
        RECT 538.950 122.850 541.050 124.950 ;
        RECT 541.950 124.050 544.050 126.150 ;
        RECT 530.100 121.050 531.900 122.850 ;
        RECT 539.100 121.050 540.900 122.850 ;
        RECT 509.400 119.700 513.150 120.750 ;
        RECT 524.400 119.700 528.150 120.750 ;
        RECT 542.850 120.750 544.050 124.050 ;
        RECT 544.950 123.450 547.050 124.050 ;
        RECT 548.550 123.450 549.450 134.550 ;
        RECT 554.100 132.150 555.900 133.950 ;
        RECT 551.100 129.150 552.900 130.950 ;
        RECT 553.950 130.050 556.050 132.150 ;
        RECT 557.250 129.150 559.050 130.950 ;
        RECT 550.950 127.050 553.050 129.150 ;
        RECT 556.950 127.050 559.050 129.150 ;
        RECT 560.400 127.950 561.300 136.200 ;
        RECT 572.100 132.150 573.900 133.950 ;
        RECT 569.100 129.150 570.900 130.950 ;
        RECT 571.950 130.050 574.050 132.150 ;
        RECT 575.250 129.150 577.050 130.950 ;
        RECT 559.950 125.850 562.050 127.950 ;
        RECT 568.950 127.050 571.050 129.150 ;
        RECT 574.950 127.050 577.050 129.150 ;
        RECT 578.400 127.950 579.300 136.200 ;
        RECT 586.800 131.400 588.600 142.500 ;
        RECT 589.800 130.500 591.600 141.600 ;
        RECT 592.800 132.600 594.600 142.500 ;
        RECT 598.800 132.600 600.600 143.400 ;
        RECT 605.400 137.400 607.200 143.400 ;
        RECT 605.700 137.100 607.200 137.400 ;
        RECT 611.400 137.400 613.200 143.400 ;
        RECT 620.400 137.400 622.200 143.400 ;
        RECT 611.400 137.100 612.300 137.400 ;
        RECT 605.700 136.200 612.300 137.100 ;
        RECT 620.700 137.100 622.200 137.400 ;
        RECT 626.400 137.400 628.200 143.400 ;
        RECT 626.400 137.100 627.300 137.400 ;
        RECT 620.700 136.200 627.300 137.100 ;
        RECT 592.800 131.700 600.600 132.600 ;
        RECT 605.100 132.150 606.900 133.950 ;
        RECT 589.800 129.600 593.850 130.500 ;
        RECT 577.950 125.850 580.050 127.950 ;
        RECT 587.100 126.150 588.900 127.950 ;
        RECT 592.950 126.150 593.850 129.600 ;
        RECT 602.100 129.150 603.900 130.950 ;
        RECT 604.950 130.050 607.050 132.150 ;
        RECT 608.250 129.150 610.050 130.950 ;
        RECT 598.950 126.150 600.750 127.950 ;
        RECT 601.950 127.050 604.050 129.150 ;
        RECT 607.950 127.050 610.050 129.150 ;
        RECT 611.400 127.950 612.300 136.200 ;
        RECT 620.100 132.150 621.900 133.950 ;
        RECT 617.100 129.150 618.900 130.950 ;
        RECT 619.950 130.050 622.050 132.150 ;
        RECT 623.250 129.150 625.050 130.950 ;
        RECT 544.950 122.550 549.450 123.450 ;
        RECT 544.950 121.950 547.050 122.550 ;
        RECT 560.400 121.650 561.300 125.850 ;
        RECT 578.400 121.650 579.300 125.850 ;
        RECT 586.950 124.050 589.050 126.150 ;
        RECT 589.950 122.850 592.050 124.950 ;
        RECT 592.950 124.050 595.050 126.150 ;
        RECT 542.850 119.700 546.600 120.750 ;
        RECT 509.400 117.600 510.600 119.700 ;
        RECT 500.400 111.600 502.200 114.600 ;
        RECT 508.800 111.600 510.600 117.600 ;
        RECT 511.800 116.700 519.600 118.050 ;
        RECT 524.400 117.600 525.600 119.700 ;
        RECT 511.800 111.600 513.600 116.700 ;
        RECT 517.800 111.600 519.600 116.700 ;
        RECT 523.800 111.600 525.600 117.600 ;
        RECT 526.800 116.700 534.600 118.050 ;
        RECT 526.800 111.600 528.600 116.700 ;
        RECT 532.800 111.600 534.600 116.700 ;
        RECT 536.400 116.700 544.200 118.050 ;
        RECT 536.400 111.600 538.200 116.700 ;
        RECT 542.400 111.600 544.200 116.700 ;
        RECT 545.400 117.600 546.600 119.700 ;
        RECT 557.100 120.000 561.300 121.650 ;
        RECT 575.100 120.000 579.300 121.650 ;
        RECT 590.250 121.050 592.050 122.850 ;
        RECT 545.400 111.600 547.200 117.600 ;
        RECT 557.100 111.600 558.900 120.000 ;
        RECT 575.100 111.600 576.900 120.000 ;
        RECT 594.000 117.600 595.050 124.050 ;
        RECT 595.950 122.850 598.050 124.950 ;
        RECT 598.950 124.050 601.050 126.150 ;
        RECT 610.950 125.850 613.050 127.950 ;
        RECT 616.950 127.050 619.050 129.150 ;
        RECT 622.950 127.050 625.050 129.150 ;
        RECT 626.400 127.950 627.300 136.200 ;
        RECT 632.400 132.300 634.200 143.400 ;
        RECT 638.400 132.300 640.200 143.400 ;
        RECT 632.400 131.400 640.200 132.300 ;
        RECT 641.400 131.400 643.200 143.400 ;
        RECT 652.800 131.400 654.600 143.400 ;
        RECT 655.800 132.300 657.600 143.400 ;
        RECT 661.800 132.300 663.600 143.400 ;
        RECT 668.400 137.400 670.200 143.400 ;
        RECT 668.700 137.100 670.200 137.400 ;
        RECT 674.400 137.400 676.200 143.400 ;
        RECT 682.800 137.400 684.600 143.400 ;
        RECT 674.400 137.100 675.300 137.400 ;
        RECT 668.700 136.200 675.300 137.100 ;
        RECT 655.800 131.400 663.600 132.300 ;
        RECT 668.100 132.150 669.900 133.950 ;
        RECT 625.950 125.850 628.050 127.950 ;
        RECT 641.700 126.150 642.600 131.400 ;
        RECT 653.400 126.150 654.300 131.400 ;
        RECT 665.100 129.150 666.900 130.950 ;
        RECT 667.950 130.050 670.050 132.150 ;
        RECT 671.250 129.150 673.050 130.950 ;
        RECT 664.950 127.050 667.050 129.150 ;
        RECT 670.950 127.050 673.050 129.150 ;
        RECT 674.400 127.950 675.300 136.200 ;
        RECT 683.700 137.100 684.600 137.400 ;
        RECT 688.800 137.400 690.600 143.400 ;
        RECT 688.800 137.100 690.300 137.400 ;
        RECT 683.700 136.200 690.300 137.100 ;
        RECT 683.700 127.950 684.600 136.200 ;
        RECT 689.100 132.150 690.900 133.950 ;
        RECT 685.950 129.150 687.750 130.950 ;
        RECT 688.950 130.050 691.050 132.150 ;
        RECT 700.500 131.400 702.300 143.400 ;
        RECT 712.800 131.400 714.600 143.400 ;
        RECT 715.800 132.300 717.600 143.400 ;
        RECT 721.800 132.300 723.600 143.400 ;
        RECT 728.400 137.400 730.200 143.400 ;
        RECT 728.700 137.100 730.200 137.400 ;
        RECT 734.400 137.400 736.200 143.400 ;
        RECT 734.400 137.100 735.300 137.400 ;
        RECT 728.700 136.200 735.300 137.100 ;
        RECT 715.800 131.400 723.600 132.300 ;
        RECT 728.100 132.150 729.900 133.950 ;
        RECT 692.100 129.150 693.900 130.950 ;
        RECT 595.950 121.050 597.750 122.850 ;
        RECT 611.400 121.650 612.300 125.850 ;
        RECT 626.400 121.650 627.300 125.850 ;
        RECT 631.950 122.850 634.050 124.950 ;
        RECT 635.100 123.150 636.900 124.950 ;
        RECT 608.100 120.000 612.300 121.650 ;
        RECT 623.100 120.000 627.300 121.650 ;
        RECT 632.100 121.050 633.900 122.850 ;
        RECT 634.950 121.050 637.050 123.150 ;
        RECT 637.950 122.850 640.050 124.950 ;
        RECT 640.950 124.050 643.050 126.150 ;
        RECT 652.950 124.050 655.050 126.150 ;
        RECT 673.950 125.850 676.050 127.950 ;
        RECT 682.950 125.850 685.050 127.950 ;
        RECT 685.950 127.050 688.050 129.150 ;
        RECT 691.950 127.050 694.050 129.150 ;
        RECT 695.100 126.150 696.900 127.950 ;
        RECT 700.950 126.150 702.150 131.400 ;
        RECT 703.950 129.150 705.750 130.950 ;
        RECT 703.950 127.050 706.050 129.150 ;
        RECT 713.400 126.150 714.300 131.400 ;
        RECT 725.100 129.150 726.900 130.950 ;
        RECT 727.950 130.050 730.050 132.150 ;
        RECT 731.250 129.150 733.050 130.950 ;
        RECT 724.950 127.050 727.050 129.150 ;
        RECT 730.950 127.050 733.050 129.150 ;
        RECT 734.400 127.950 735.300 136.200 ;
        RECT 745.800 131.400 747.600 143.400 ;
        RECT 748.800 132.300 750.600 143.400 ;
        RECT 754.800 132.300 756.600 143.400 ;
        RECT 748.800 131.400 756.600 132.300 ;
        RECT 638.100 121.050 639.900 122.850 ;
        RECT 594.000 111.600 595.800 117.600 ;
        RECT 608.100 111.600 609.900 120.000 ;
        RECT 623.100 111.600 624.900 120.000 ;
        RECT 641.700 117.600 642.600 124.050 ;
        RECT 637.200 115.950 642.600 117.600 ;
        RECT 653.400 117.600 654.300 124.050 ;
        RECT 655.950 122.850 658.050 124.950 ;
        RECT 659.100 123.150 660.900 124.950 ;
        RECT 656.100 121.050 657.900 122.850 ;
        RECT 658.950 121.050 661.050 123.150 ;
        RECT 661.950 122.850 664.050 124.950 ;
        RECT 662.100 121.050 663.900 122.850 ;
        RECT 674.400 121.650 675.300 125.850 ;
        RECT 671.100 120.000 675.300 121.650 ;
        RECT 683.700 121.650 684.600 125.850 ;
        RECT 694.950 124.050 697.050 126.150 ;
        RECT 697.950 122.850 700.050 124.950 ;
        RECT 700.950 124.050 703.050 126.150 ;
        RECT 712.950 124.050 715.050 126.150 ;
        RECT 733.950 125.850 736.050 127.950 ;
        RECT 746.400 126.150 747.300 131.400 ;
        RECT 683.700 120.000 687.900 121.650 ;
        RECT 698.100 121.050 699.900 122.850 ;
        RECT 653.400 115.950 658.800 117.600 ;
        RECT 637.200 111.600 639.000 115.950 ;
        RECT 657.000 111.600 658.800 115.950 ;
        RECT 671.100 111.600 672.900 120.000 ;
        RECT 686.100 111.600 687.900 120.000 ;
        RECT 701.850 120.750 703.050 124.050 ;
        RECT 701.850 119.700 705.600 120.750 ;
        RECT 695.400 116.700 703.200 118.050 ;
        RECT 695.400 111.600 697.200 116.700 ;
        RECT 701.400 111.600 703.200 116.700 ;
        RECT 704.400 117.600 705.600 119.700 ;
        RECT 713.400 117.600 714.300 124.050 ;
        RECT 715.950 122.850 718.050 124.950 ;
        RECT 719.100 123.150 720.900 124.950 ;
        RECT 716.100 121.050 717.900 122.850 ;
        RECT 718.950 121.050 721.050 123.150 ;
        RECT 721.950 122.850 724.050 124.950 ;
        RECT 722.100 121.050 723.900 122.850 ;
        RECT 734.400 121.650 735.300 125.850 ;
        RECT 745.950 124.050 748.050 126.150 ;
        RECT 731.100 120.000 735.300 121.650 ;
        RECT 704.400 111.600 706.200 117.600 ;
        RECT 713.400 115.950 718.800 117.600 ;
        RECT 717.000 111.600 718.800 115.950 ;
        RECT 731.100 111.600 732.900 120.000 ;
        RECT 746.400 117.600 747.300 124.050 ;
        RECT 748.950 122.850 751.050 124.950 ;
        RECT 752.100 123.150 753.900 124.950 ;
        RECT 749.100 121.050 750.900 122.850 ;
        RECT 751.950 121.050 754.050 123.150 ;
        RECT 754.950 122.850 757.050 124.950 ;
        RECT 755.100 121.050 756.900 122.850 ;
        RECT 746.400 115.950 751.800 117.600 ;
        RECT 750.000 111.600 751.800 115.950 ;
        RECT 11.100 99.000 12.900 107.400 ;
        RECT 20.400 102.300 22.200 107.400 ;
        RECT 26.400 102.300 28.200 107.400 ;
        RECT 20.400 100.950 28.200 102.300 ;
        RECT 29.400 101.400 31.200 107.400 ;
        RECT 29.400 99.300 30.600 101.400 ;
        RECT 8.700 97.350 12.900 99.000 ;
        RECT 26.850 98.250 30.600 99.300 ;
        RECT 41.100 99.000 42.900 107.400 ;
        RECT 50.400 102.300 52.200 107.400 ;
        RECT 56.400 102.300 58.200 107.400 ;
        RECT 50.400 100.950 58.200 102.300 ;
        RECT 59.400 101.400 61.200 107.400 ;
        RECT 71.400 104.400 73.200 107.400 ;
        RECT 59.400 99.300 60.600 101.400 ;
        RECT 8.700 93.150 9.600 97.350 ;
        RECT 23.100 96.150 24.900 97.950 ;
        RECT 7.950 91.050 10.050 93.150 ;
        RECT 19.950 92.850 22.050 94.950 ;
        RECT 22.950 94.050 25.050 96.150 ;
        RECT 26.850 94.950 28.050 98.250 ;
        RECT 41.100 97.350 45.300 99.000 ;
        RECT 56.850 98.250 60.600 99.300 ;
        RECT 28.950 96.450 31.050 97.050 ;
        RECT 34.950 96.450 37.050 97.050 ;
        RECT 28.950 95.550 37.050 96.450 ;
        RECT 28.950 94.950 31.050 95.550 ;
        RECT 34.950 94.950 37.050 95.550 ;
        RECT 25.950 92.850 28.050 94.950 ;
        RECT 44.400 93.150 45.300 97.350 ;
        RECT 53.100 96.150 54.900 97.950 ;
        RECT 8.700 82.800 9.600 91.050 ;
        RECT 10.950 89.850 13.050 91.950 ;
        RECT 16.950 89.850 19.050 91.950 ;
        RECT 20.100 91.050 21.900 92.850 ;
        RECT 10.950 88.050 12.750 89.850 ;
        RECT 13.950 86.850 16.050 88.950 ;
        RECT 17.100 88.050 18.900 89.850 ;
        RECT 25.950 87.600 27.150 92.850 ;
        RECT 28.950 89.850 31.050 91.950 ;
        RECT 34.950 89.850 37.050 91.950 ;
        RECT 40.950 89.850 43.050 91.950 ;
        RECT 43.950 91.050 46.050 93.150 ;
        RECT 49.950 92.850 52.050 94.950 ;
        RECT 52.950 94.050 55.050 96.150 ;
        RECT 56.850 94.950 58.050 98.250 ;
        RECT 67.950 95.850 70.050 97.950 ;
        RECT 71.400 96.150 72.600 104.400 ;
        RECT 83.100 99.000 84.900 107.400 ;
        RECT 97.800 101.400 99.600 107.400 ;
        RECT 98.400 99.300 99.600 101.400 ;
        RECT 100.800 102.300 102.600 107.400 ;
        RECT 106.800 102.300 108.600 107.400 ;
        RECT 100.800 100.950 108.600 102.300 ;
        RECT 113.400 104.400 115.200 107.400 ;
        RECT 83.100 97.350 87.300 99.000 ;
        RECT 98.400 98.250 102.150 99.300 ;
        RECT 55.950 92.850 58.050 94.950 ;
        RECT 68.100 94.050 69.900 95.850 ;
        RECT 70.950 94.050 73.050 96.150 ;
        RECT 50.100 91.050 51.900 92.850 ;
        RECT 28.950 88.050 30.750 89.850 ;
        RECT 35.100 88.050 36.900 89.850 ;
        RECT 14.100 85.050 15.900 86.850 ;
        RECT 8.700 81.900 15.300 82.800 ;
        RECT 8.700 81.600 9.600 81.900 ;
        RECT 7.800 75.600 9.600 81.600 ;
        RECT 13.800 81.600 15.300 81.900 ;
        RECT 13.800 75.600 15.600 81.600 ;
        RECT 25.500 75.600 27.300 87.600 ;
        RECT 37.950 86.850 40.050 88.950 ;
        RECT 41.250 88.050 43.050 89.850 ;
        RECT 38.100 85.050 39.900 86.850 ;
        RECT 44.400 82.800 45.300 91.050 ;
        RECT 55.950 87.600 57.150 92.850 ;
        RECT 58.950 89.850 61.050 91.950 ;
        RECT 58.950 88.050 60.750 89.850 ;
        RECT 38.700 81.900 45.300 82.800 ;
        RECT 38.700 81.600 40.200 81.900 ;
        RECT 38.400 75.600 40.200 81.600 ;
        RECT 44.400 81.600 45.300 81.900 ;
        RECT 44.400 75.600 46.200 81.600 ;
        RECT 55.500 75.600 57.300 87.600 ;
        RECT 71.400 81.600 72.600 94.050 ;
        RECT 86.400 93.150 87.300 97.350 ;
        RECT 100.950 94.950 102.150 98.250 ;
        RECT 104.100 96.150 105.900 97.950 ;
        RECT 76.950 89.850 79.050 91.950 ;
        RECT 82.950 89.850 85.050 91.950 ;
        RECT 85.950 91.050 88.050 93.150 ;
        RECT 100.950 92.850 103.050 94.950 ;
        RECT 103.950 94.050 106.050 96.150 ;
        RECT 109.950 95.850 112.050 97.950 ;
        RECT 113.400 96.150 114.600 104.400 ;
        RECT 129.000 103.050 130.800 107.400 ;
        RECT 125.400 101.400 130.800 103.050 ;
        RECT 139.800 101.400 141.600 107.400 ;
        RECT 145.800 104.400 147.600 107.400 ;
        RECT 106.950 92.850 109.050 94.950 ;
        RECT 110.100 94.050 111.900 95.850 ;
        RECT 112.950 94.050 115.050 96.150 ;
        RECT 125.400 94.950 126.300 101.400 ;
        RECT 128.100 96.150 129.900 97.950 ;
        RECT 77.100 88.050 78.900 89.850 ;
        RECT 79.950 86.850 82.050 88.950 ;
        RECT 83.250 88.050 85.050 89.850 ;
        RECT 80.100 85.050 81.900 86.850 ;
        RECT 86.400 82.800 87.300 91.050 ;
        RECT 97.950 89.850 100.050 91.950 ;
        RECT 98.250 88.050 100.050 89.850 ;
        RECT 101.850 87.600 103.050 92.850 ;
        RECT 107.100 91.050 108.900 92.850 ;
        RECT 80.700 81.900 87.300 82.800 ;
        RECT 80.700 81.600 82.200 81.900 ;
        RECT 71.400 75.600 73.200 81.600 ;
        RECT 80.400 75.600 82.200 81.600 ;
        RECT 86.400 81.600 87.300 81.900 ;
        RECT 86.400 75.600 88.200 81.600 ;
        RECT 101.700 75.600 103.500 87.600 ;
        RECT 113.400 81.600 114.600 94.050 ;
        RECT 124.950 92.850 127.050 94.950 ;
        RECT 127.950 94.050 130.050 96.150 ;
        RECT 130.950 95.850 133.050 97.950 ;
        RECT 134.100 96.150 135.900 97.950 ;
        RECT 139.950 96.150 141.000 101.400 ;
        RECT 145.800 100.200 146.700 104.400 ;
        RECT 159.000 103.050 160.800 107.400 ;
        RECT 143.250 99.300 146.700 100.200 ;
        RECT 155.400 101.400 160.800 103.050 ;
        RECT 143.250 98.400 145.050 99.300 ;
        RECT 131.100 94.050 132.900 95.850 ;
        RECT 133.950 94.050 136.050 96.150 ;
        RECT 139.950 94.050 142.050 96.150 ;
        RECT 125.400 87.600 126.300 92.850 ;
        RECT 113.400 75.600 115.200 81.600 ;
        RECT 124.800 75.600 126.600 87.600 ;
        RECT 127.800 86.700 135.600 87.600 ;
        RECT 127.800 75.600 129.600 86.700 ;
        RECT 133.800 75.600 135.600 86.700 ;
        RECT 140.700 87.450 142.050 94.050 ;
        RECT 143.400 90.150 144.300 98.400 ;
        RECT 148.950 95.850 151.050 97.950 ;
        RECT 145.950 92.850 148.050 94.950 ;
        RECT 149.100 94.050 150.900 95.850 ;
        RECT 155.400 94.950 156.300 101.400 ;
        RECT 176.100 99.000 177.900 107.400 ;
        RECT 188.400 102.300 190.200 107.400 ;
        RECT 194.400 102.300 196.200 107.400 ;
        RECT 188.400 100.950 196.200 102.300 ;
        RECT 197.400 101.400 199.200 107.400 ;
        RECT 206.400 104.400 208.200 107.400 ;
        RECT 197.400 99.300 198.600 101.400 ;
        RECT 158.100 96.150 159.900 97.950 ;
        RECT 154.950 92.850 157.050 94.950 ;
        RECT 157.950 94.050 160.050 96.150 ;
        RECT 160.950 95.850 163.050 97.950 ;
        RECT 164.100 96.150 165.900 97.950 ;
        RECT 173.700 97.350 177.900 99.000 ;
        RECT 194.850 98.250 198.600 99.300 ;
        RECT 161.100 94.050 162.900 95.850 ;
        RECT 163.950 94.050 166.050 96.150 ;
        RECT 173.700 93.150 174.600 97.350 ;
        RECT 191.100 96.150 192.900 97.950 ;
        RECT 146.100 91.050 147.900 92.850 ;
        RECT 143.400 90.000 145.200 90.150 ;
        RECT 143.400 88.800 150.600 90.000 ;
        RECT 143.400 88.350 145.200 88.800 ;
        RECT 149.400 87.600 150.600 88.800 ;
        RECT 155.400 87.600 156.300 92.850 ;
        RECT 172.950 91.050 175.050 93.150 ;
        RECT 187.950 92.850 190.050 94.950 ;
        RECT 190.950 94.050 193.050 96.150 ;
        RECT 194.850 94.950 196.050 98.250 ;
        RECT 202.950 95.850 205.050 97.950 ;
        RECT 206.400 96.150 207.600 104.400 ;
        RECT 217.200 100.200 219.000 107.400 ;
        RECT 215.400 99.300 219.000 100.200 ;
        RECT 193.950 92.850 196.050 94.950 ;
        RECT 203.100 94.050 204.900 95.850 ;
        RECT 205.950 94.050 208.050 96.150 ;
        RECT 140.700 86.100 143.100 87.450 ;
        RECT 141.300 75.600 143.100 86.100 ;
        RECT 148.800 75.600 150.600 87.600 ;
        RECT 154.800 75.600 156.600 87.600 ;
        RECT 157.800 86.700 165.600 87.600 ;
        RECT 157.800 75.600 159.600 86.700 ;
        RECT 163.800 75.600 165.600 86.700 ;
        RECT 173.700 82.800 174.600 91.050 ;
        RECT 175.950 89.850 178.050 91.950 ;
        RECT 181.950 89.850 184.050 91.950 ;
        RECT 188.100 91.050 189.900 92.850 ;
        RECT 175.950 88.050 177.750 89.850 ;
        RECT 178.950 86.850 181.050 88.950 ;
        RECT 182.100 88.050 183.900 89.850 ;
        RECT 193.950 87.600 195.150 92.850 ;
        RECT 196.950 89.850 199.050 91.950 ;
        RECT 196.950 88.050 198.750 89.850 ;
        RECT 179.100 85.050 180.900 86.850 ;
        RECT 173.700 81.900 180.300 82.800 ;
        RECT 173.700 81.600 174.600 81.900 ;
        RECT 172.800 75.600 174.600 81.600 ;
        RECT 178.800 81.600 180.300 81.900 ;
        RECT 178.800 75.600 180.600 81.600 ;
        RECT 193.500 75.600 195.300 87.600 ;
        RECT 206.400 81.600 207.600 94.050 ;
        RECT 212.100 93.150 213.900 94.950 ;
        RECT 211.950 91.050 214.050 93.150 ;
        RECT 215.400 91.950 216.600 99.300 ;
        RECT 230.100 99.000 231.900 107.400 ;
        RECT 244.800 104.400 246.600 107.400 ;
        RECT 230.100 97.350 234.300 99.000 ;
        RECT 218.100 93.150 219.900 94.950 ;
        RECT 233.400 93.150 234.300 97.350 ;
        RECT 244.950 97.950 246.000 104.400 ;
        RECT 253.800 101.400 255.600 107.400 ;
        RECT 259.800 104.400 261.600 107.400 ;
        RECT 244.950 95.850 247.050 97.950 ;
        RECT 253.950 96.150 255.000 101.400 ;
        RECT 259.800 100.200 260.700 104.400 ;
        RECT 257.250 99.300 260.700 100.200 ;
        RECT 257.250 98.400 259.050 99.300 ;
        RECT 272.100 99.000 273.900 107.400 ;
        RECT 291.000 103.050 292.800 107.400 ;
        RECT 214.950 89.850 217.050 91.950 ;
        RECT 217.950 91.050 220.050 93.150 ;
        RECT 223.950 89.850 226.050 91.950 ;
        RECT 229.950 89.850 232.050 91.950 ;
        RECT 232.950 91.050 235.050 93.150 ;
        RECT 241.950 92.850 244.050 94.950 ;
        RECT 242.100 91.050 243.900 92.850 ;
        RECT 215.400 81.600 216.600 89.850 ;
        RECT 224.100 88.050 225.900 89.850 ;
        RECT 226.950 86.850 229.050 88.950 ;
        RECT 230.250 88.050 232.050 89.850 ;
        RECT 227.100 85.050 228.900 86.850 ;
        RECT 233.400 82.800 234.300 91.050 ;
        RECT 244.950 88.650 246.000 95.850 ;
        RECT 247.950 92.850 250.050 94.950 ;
        RECT 253.950 94.050 256.050 96.150 ;
        RECT 248.100 91.050 249.900 92.850 ;
        RECT 227.700 81.900 234.300 82.800 ;
        RECT 227.700 81.600 229.200 81.900 ;
        RECT 206.400 75.600 208.200 81.600 ;
        RECT 215.400 75.600 217.200 81.600 ;
        RECT 227.400 75.600 229.200 81.600 ;
        RECT 233.400 81.600 234.300 81.900 ;
        RECT 243.600 87.600 246.000 88.650 ;
        RECT 233.400 75.600 235.200 81.600 ;
        RECT 243.600 75.600 245.400 87.600 ;
        RECT 254.700 87.450 256.050 94.050 ;
        RECT 257.400 90.150 258.300 98.400 ;
        RECT 262.950 95.850 265.050 97.950 ;
        RECT 269.700 97.350 273.900 99.000 ;
        RECT 287.400 101.400 292.800 103.050 ;
        RECT 259.950 92.850 262.050 94.950 ;
        RECT 263.100 94.050 264.900 95.850 ;
        RECT 269.700 93.150 270.600 97.350 ;
        RECT 287.400 94.950 288.300 101.400 ;
        RECT 305.100 99.000 306.900 107.400 ;
        RECT 316.800 101.400 318.600 107.400 ;
        RECT 317.400 99.300 318.600 101.400 ;
        RECT 319.800 102.300 321.600 107.400 ;
        RECT 325.800 102.300 327.600 107.400 ;
        RECT 336.000 103.050 337.800 107.400 ;
        RECT 319.800 100.950 327.600 102.300 ;
        RECT 332.400 101.400 337.800 103.050 ;
        RECT 351.300 102.900 353.100 107.400 ;
        RECT 349.950 101.400 353.100 102.900 ;
        RECT 290.100 96.150 291.900 97.950 ;
        RECT 260.100 91.050 261.900 92.850 ;
        RECT 268.950 91.050 271.050 93.150 ;
        RECT 286.950 92.850 289.050 94.950 ;
        RECT 289.950 94.050 292.050 96.150 ;
        RECT 292.950 95.850 295.050 97.950 ;
        RECT 296.100 96.150 297.900 97.950 ;
        RECT 305.100 97.350 309.300 99.000 ;
        RECT 317.400 98.250 321.150 99.300 ;
        RECT 293.100 94.050 294.900 95.850 ;
        RECT 295.950 94.050 298.050 96.150 ;
        RECT 308.400 93.150 309.300 97.350 ;
        RECT 319.950 94.950 321.150 98.250 ;
        RECT 323.100 96.150 324.900 97.950 ;
        RECT 257.400 90.000 259.200 90.150 ;
        RECT 257.400 88.800 264.600 90.000 ;
        RECT 257.400 88.350 259.200 88.800 ;
        RECT 263.400 87.600 264.600 88.800 ;
        RECT 254.700 86.100 257.100 87.450 ;
        RECT 255.300 75.600 257.100 86.100 ;
        RECT 262.800 75.600 264.600 87.600 ;
        RECT 269.700 82.800 270.600 91.050 ;
        RECT 271.950 89.850 274.050 91.950 ;
        RECT 277.950 89.850 280.050 91.950 ;
        RECT 271.950 88.050 273.750 89.850 ;
        RECT 274.950 86.850 277.050 88.950 ;
        RECT 278.100 88.050 279.900 89.850 ;
        RECT 287.400 87.600 288.300 92.850 ;
        RECT 298.950 89.850 301.050 91.950 ;
        RECT 304.950 89.850 307.050 91.950 ;
        RECT 307.950 91.050 310.050 93.150 ;
        RECT 319.950 92.850 322.050 94.950 ;
        RECT 322.950 94.050 325.050 96.150 ;
        RECT 332.400 94.950 333.300 101.400 ;
        RECT 335.100 96.150 336.900 97.950 ;
        RECT 325.950 92.850 328.050 94.950 ;
        RECT 331.950 92.850 334.050 94.950 ;
        RECT 334.950 94.050 337.050 96.150 ;
        RECT 337.950 95.850 340.050 97.950 ;
        RECT 341.100 96.150 342.900 97.950 ;
        RECT 338.100 94.050 339.900 95.850 ;
        RECT 340.950 94.050 343.050 96.150 ;
        RECT 349.950 94.950 351.000 101.400 ;
        RECT 353.100 99.900 354.900 100.500 ;
        RECT 358.800 99.900 360.600 107.400 ;
        RECT 367.200 101.400 369.000 107.400 ;
        RECT 353.100 98.700 360.600 99.900 ;
        RECT 349.950 92.850 352.050 94.950 ;
        RECT 353.100 93.150 354.900 94.950 ;
        RECT 299.100 88.050 300.900 89.850 ;
        RECT 275.100 85.050 276.900 86.850 ;
        RECT 269.700 81.900 276.300 82.800 ;
        RECT 269.700 81.600 270.600 81.900 ;
        RECT 268.800 75.600 270.600 81.600 ;
        RECT 274.800 81.600 276.300 81.900 ;
        RECT 274.800 75.600 276.600 81.600 ;
        RECT 286.800 75.600 288.600 87.600 ;
        RECT 289.800 86.700 297.600 87.600 ;
        RECT 301.950 86.850 304.050 88.950 ;
        RECT 305.250 88.050 307.050 89.850 ;
        RECT 289.800 75.600 291.600 86.700 ;
        RECT 295.800 75.600 297.600 86.700 ;
        RECT 302.100 85.050 303.900 86.850 ;
        RECT 308.400 82.800 309.300 91.050 ;
        RECT 316.950 89.850 319.050 91.950 ;
        RECT 317.250 88.050 319.050 89.850 ;
        RECT 320.850 87.600 322.050 92.850 ;
        RECT 326.100 91.050 327.900 92.850 ;
        RECT 332.400 87.600 333.300 92.850 ;
        RECT 349.950 87.600 351.000 92.850 ;
        RECT 352.950 91.050 355.050 93.150 ;
        RECT 302.700 81.900 309.300 82.800 ;
        RECT 302.700 81.600 304.200 81.900 ;
        RECT 302.400 75.600 304.200 81.600 ;
        RECT 308.400 81.600 309.300 81.900 ;
        RECT 308.400 75.600 310.200 81.600 ;
        RECT 320.700 75.600 322.500 87.600 ;
        RECT 331.800 75.600 333.600 87.600 ;
        RECT 334.800 86.700 342.600 87.600 ;
        RECT 334.800 75.600 336.600 86.700 ;
        RECT 340.800 75.600 342.600 86.700 ;
        RECT 349.200 75.600 351.000 87.600 ;
        RECT 356.400 81.600 357.450 98.700 ;
        RECT 365.250 96.150 367.050 97.950 ;
        RECT 358.950 92.850 361.050 94.950 ;
        RECT 361.950 92.850 364.050 94.950 ;
        RECT 364.950 94.050 367.050 96.150 ;
        RECT 367.950 94.950 369.000 101.400 ;
        RECT 386.100 99.000 387.900 107.400 ;
        RECT 401.100 99.000 402.900 107.400 ;
        RECT 415.200 103.050 417.000 107.400 ;
        RECT 415.200 101.400 420.600 103.050 ;
        RECT 370.950 96.150 372.750 97.950 ;
        RECT 386.100 97.350 390.300 99.000 ;
        RECT 367.950 92.850 370.050 94.950 ;
        RECT 370.950 94.050 373.050 96.150 ;
        RECT 373.950 92.850 376.050 94.950 ;
        RECT 389.400 93.150 390.300 97.350 ;
        RECT 398.700 97.350 402.900 99.000 ;
        RECT 398.700 93.150 399.600 97.350 ;
        RECT 410.100 96.150 411.900 97.950 ;
        RECT 409.950 94.050 412.050 96.150 ;
        RECT 412.950 95.850 415.050 97.950 ;
        RECT 416.100 96.150 417.900 97.950 ;
        RECT 413.100 94.050 414.900 95.850 ;
        RECT 415.950 94.050 418.050 96.150 ;
        RECT 419.700 94.950 420.600 101.400 ;
        RECT 435.000 101.400 436.800 107.400 ;
        RECT 431.250 96.150 433.050 97.950 ;
        RECT 359.100 91.050 360.900 92.850 ;
        RECT 362.250 91.050 364.050 92.850 ;
        RECT 369.150 89.400 370.050 92.850 ;
        RECT 374.100 91.050 375.900 92.850 ;
        RECT 379.950 89.850 382.050 91.950 ;
        RECT 385.950 89.850 388.050 91.950 ;
        RECT 388.950 91.050 391.050 93.150 ;
        RECT 397.950 91.050 400.050 93.150 ;
        RECT 418.950 92.850 421.050 94.950 ;
        RECT 427.950 92.850 430.050 94.950 ;
        RECT 430.950 94.050 433.050 96.150 ;
        RECT 435.000 94.950 436.050 101.400 ;
        RECT 452.100 99.000 453.900 107.400 ;
        RECT 468.000 103.050 469.800 107.400 ;
        RECT 478.800 104.400 480.600 107.400 ;
        RECT 464.400 101.400 469.800 103.050 ;
        RECT 433.950 92.850 436.050 94.950 ;
        RECT 436.950 96.150 438.750 97.950 ;
        RECT 452.100 97.350 456.300 99.000 ;
        RECT 445.950 96.450 448.050 97.050 ;
        RECT 436.950 94.050 439.050 96.150 ;
        RECT 443.550 95.550 448.050 96.450 ;
        RECT 439.950 92.850 442.050 94.950 ;
        RECT 369.150 88.500 373.200 89.400 ;
        RECT 362.400 86.400 370.200 87.300 ;
        RECT 355.800 75.600 357.600 81.600 ;
        RECT 362.400 75.600 364.200 86.400 ;
        RECT 368.400 76.500 370.200 86.400 ;
        RECT 371.400 77.400 373.200 88.500 ;
        RECT 380.100 88.050 381.900 89.850 ;
        RECT 374.400 76.500 376.200 87.600 ;
        RECT 382.950 86.850 385.050 88.950 ;
        RECT 386.250 88.050 388.050 89.850 ;
        RECT 383.100 85.050 384.900 86.850 ;
        RECT 389.400 82.800 390.300 91.050 ;
        RECT 383.700 81.900 390.300 82.800 ;
        RECT 383.700 81.600 385.200 81.900 ;
        RECT 368.400 75.600 376.200 76.500 ;
        RECT 383.400 75.600 385.200 81.600 ;
        RECT 389.400 81.600 390.300 81.900 ;
        RECT 398.700 82.800 399.600 91.050 ;
        RECT 400.950 89.850 403.050 91.950 ;
        RECT 406.950 89.850 409.050 91.950 ;
        RECT 400.950 88.050 402.750 89.850 ;
        RECT 403.950 86.850 406.050 88.950 ;
        RECT 407.100 88.050 408.900 89.850 ;
        RECT 419.700 87.600 420.600 92.850 ;
        RECT 428.100 91.050 429.900 92.850 ;
        RECT 433.950 89.400 434.850 92.850 ;
        RECT 439.950 91.050 441.750 92.850 ;
        RECT 430.800 88.500 434.850 89.400 ;
        RECT 404.100 85.050 405.900 86.850 ;
        RECT 410.400 86.700 418.200 87.600 ;
        RECT 398.700 81.900 405.300 82.800 ;
        RECT 398.700 81.600 399.600 81.900 ;
        RECT 389.400 75.600 391.200 81.600 ;
        RECT 397.800 75.600 399.600 81.600 ;
        RECT 403.800 81.600 405.300 81.900 ;
        RECT 403.800 75.600 405.600 81.600 ;
        RECT 410.400 75.600 412.200 86.700 ;
        RECT 416.400 75.600 418.200 86.700 ;
        RECT 419.400 75.600 421.200 87.600 ;
        RECT 427.800 76.500 429.600 87.600 ;
        RECT 430.800 77.400 432.600 88.500 ;
        RECT 433.800 86.400 441.600 87.300 ;
        RECT 433.800 76.500 435.600 86.400 ;
        RECT 427.800 75.600 435.600 76.500 ;
        RECT 439.800 75.600 441.600 86.400 ;
        RECT 443.550 84.450 444.450 95.550 ;
        RECT 445.950 94.950 448.050 95.550 ;
        RECT 455.400 93.150 456.300 97.350 ;
        RECT 464.400 94.950 465.300 101.400 ;
        RECT 467.100 96.150 468.900 97.950 ;
        RECT 445.950 89.850 448.050 91.950 ;
        RECT 451.950 89.850 454.050 91.950 ;
        RECT 454.950 91.050 457.050 93.150 ;
        RECT 463.950 92.850 466.050 94.950 ;
        RECT 466.950 94.050 469.050 96.150 ;
        RECT 469.950 95.850 472.050 97.950 ;
        RECT 473.100 96.150 474.900 97.950 ;
        RECT 479.400 96.150 480.600 104.400 ;
        RECT 491.100 99.000 492.900 107.400 ;
        RECT 505.800 101.400 507.600 107.400 ;
        RECT 470.100 94.050 471.900 95.850 ;
        RECT 472.950 94.050 475.050 96.150 ;
        RECT 478.950 94.050 481.050 96.150 ;
        RECT 481.950 95.850 484.050 97.950 ;
        RECT 488.700 97.350 492.900 99.000 ;
        RECT 506.400 99.300 507.600 101.400 ;
        RECT 508.800 102.300 510.600 107.400 ;
        RECT 514.800 102.300 516.600 107.400 ;
        RECT 508.800 100.950 516.600 102.300 ;
        RECT 506.400 98.250 510.150 99.300 ;
        RECT 524.100 99.000 525.900 107.400 ;
        RECT 540.000 103.050 541.800 107.400 ;
        RECT 555.000 103.050 556.800 107.400 ;
        RECT 482.100 94.050 483.900 95.850 ;
        RECT 446.100 88.050 447.900 89.850 ;
        RECT 448.950 86.850 451.050 88.950 ;
        RECT 452.250 88.050 454.050 89.850 ;
        RECT 449.100 85.050 450.900 86.850 ;
        RECT 445.950 84.450 448.050 85.050 ;
        RECT 443.550 83.550 448.050 84.450 ;
        RECT 445.950 82.950 448.050 83.550 ;
        RECT 455.400 82.800 456.300 91.050 ;
        RECT 464.400 87.600 465.300 92.850 ;
        RECT 449.700 81.900 456.300 82.800 ;
        RECT 449.700 81.600 451.200 81.900 ;
        RECT 449.400 75.600 451.200 81.600 ;
        RECT 455.400 81.600 456.300 81.900 ;
        RECT 455.400 75.600 457.200 81.600 ;
        RECT 463.800 75.600 465.600 87.600 ;
        RECT 466.800 86.700 474.600 87.600 ;
        RECT 466.800 75.600 468.600 86.700 ;
        RECT 472.800 75.600 474.600 86.700 ;
        RECT 479.400 81.600 480.600 94.050 ;
        RECT 488.700 93.150 489.600 97.350 ;
        RECT 508.950 94.950 510.150 98.250 ;
        RECT 512.100 96.150 513.900 97.950 ;
        RECT 521.700 97.350 525.900 99.000 ;
        RECT 536.400 101.400 541.800 103.050 ;
        RECT 551.400 101.400 556.800 103.050 ;
        RECT 487.950 91.050 490.050 93.150 ;
        RECT 508.950 92.850 511.050 94.950 ;
        RECT 511.950 94.050 514.050 96.150 ;
        RECT 514.950 92.850 517.050 94.950 ;
        RECT 521.700 93.150 522.600 97.350 ;
        RECT 536.400 94.950 537.300 101.400 ;
        RECT 539.100 96.150 540.900 97.950 ;
        RECT 488.700 82.800 489.600 91.050 ;
        RECT 490.950 89.850 493.050 91.950 ;
        RECT 496.950 89.850 499.050 91.950 ;
        RECT 505.950 89.850 508.050 91.950 ;
        RECT 490.950 88.050 492.750 89.850 ;
        RECT 493.950 86.850 496.050 88.950 ;
        RECT 497.100 88.050 498.900 89.850 ;
        RECT 506.250 88.050 508.050 89.850 ;
        RECT 509.850 87.600 511.050 92.850 ;
        RECT 515.100 91.050 516.900 92.850 ;
        RECT 520.950 91.050 523.050 93.150 ;
        RECT 535.950 92.850 538.050 94.950 ;
        RECT 538.950 94.050 541.050 96.150 ;
        RECT 541.950 95.850 544.050 97.950 ;
        RECT 545.100 96.150 546.900 97.950 ;
        RECT 542.100 94.050 543.900 95.850 ;
        RECT 544.950 94.050 547.050 96.150 ;
        RECT 551.400 94.950 552.300 101.400 ;
        RECT 569.100 99.000 570.900 107.400 ;
        RECT 581.400 104.400 583.200 107.400 ;
        RECT 593.400 104.400 595.200 107.400 ;
        RECT 554.100 96.150 555.900 97.950 ;
        RECT 550.950 92.850 553.050 94.950 ;
        RECT 553.950 94.050 556.050 96.150 ;
        RECT 556.950 95.850 559.050 97.950 ;
        RECT 560.100 96.150 561.900 97.950 ;
        RECT 569.100 97.350 573.300 99.000 ;
        RECT 557.100 94.050 558.900 95.850 ;
        RECT 559.950 94.050 562.050 96.150 ;
        RECT 572.400 93.150 573.300 97.350 ;
        RECT 577.950 95.850 580.050 97.950 ;
        RECT 581.400 96.150 582.600 104.400 ;
        RECT 578.100 94.050 579.900 95.850 ;
        RECT 580.950 94.050 583.050 96.150 ;
        RECT 589.950 95.850 592.050 97.950 ;
        RECT 593.400 96.150 594.600 104.400 ;
        RECT 606.000 100.200 607.800 107.400 ;
        RECT 606.000 99.300 609.600 100.200 ;
        RECT 590.100 94.050 591.900 95.850 ;
        RECT 592.950 94.050 595.050 96.150 ;
        RECT 494.100 85.050 495.900 86.850 ;
        RECT 488.700 81.900 495.300 82.800 ;
        RECT 488.700 81.600 489.600 81.900 ;
        RECT 478.800 75.600 480.600 81.600 ;
        RECT 487.800 75.600 489.600 81.600 ;
        RECT 493.800 81.600 495.300 81.900 ;
        RECT 493.800 75.600 495.600 81.600 ;
        RECT 509.700 75.600 511.500 87.600 ;
        RECT 521.700 82.800 522.600 91.050 ;
        RECT 523.950 89.850 526.050 91.950 ;
        RECT 529.950 89.850 532.050 91.950 ;
        RECT 523.950 88.050 525.750 89.850 ;
        RECT 526.950 86.850 529.050 88.950 ;
        RECT 530.100 88.050 531.900 89.850 ;
        RECT 536.400 87.600 537.300 92.850 ;
        RECT 551.400 87.600 552.300 92.850 ;
        RECT 562.950 89.850 565.050 91.950 ;
        RECT 568.950 89.850 571.050 91.950 ;
        RECT 571.950 91.050 574.050 93.150 ;
        RECT 563.100 88.050 564.900 89.850 ;
        RECT 527.100 85.050 528.900 86.850 ;
        RECT 521.700 81.900 528.300 82.800 ;
        RECT 521.700 81.600 522.600 81.900 ;
        RECT 520.800 75.600 522.600 81.600 ;
        RECT 526.800 81.600 528.300 81.900 ;
        RECT 526.800 75.600 528.600 81.600 ;
        RECT 535.800 75.600 537.600 87.600 ;
        RECT 538.800 86.700 546.600 87.600 ;
        RECT 538.800 75.600 540.600 86.700 ;
        RECT 544.800 75.600 546.600 86.700 ;
        RECT 550.800 75.600 552.600 87.600 ;
        RECT 553.800 86.700 561.600 87.600 ;
        RECT 565.950 86.850 568.050 88.950 ;
        RECT 569.250 88.050 571.050 89.850 ;
        RECT 553.800 75.600 555.600 86.700 ;
        RECT 559.800 75.600 561.600 86.700 ;
        RECT 566.100 85.050 567.900 86.850 ;
        RECT 572.400 82.800 573.300 91.050 ;
        RECT 566.700 81.900 573.300 82.800 ;
        RECT 566.700 81.600 568.200 81.900 ;
        RECT 566.400 75.600 568.200 81.600 ;
        RECT 572.400 81.600 573.300 81.900 ;
        RECT 581.400 81.600 582.600 94.050 ;
        RECT 593.400 81.600 594.600 94.050 ;
        RECT 605.100 93.150 606.900 94.950 ;
        RECT 604.950 91.050 607.050 93.150 ;
        RECT 608.400 91.950 609.600 99.300 ;
        RECT 614.400 99.900 616.200 107.400 ;
        RECT 621.900 102.900 623.700 107.400 ;
        RECT 636.000 103.050 637.800 107.400 ;
        RECT 621.900 101.400 625.050 102.900 ;
        RECT 620.100 99.900 621.900 100.500 ;
        RECT 614.400 98.700 621.900 99.900 ;
        RECT 611.100 93.150 612.900 94.950 ;
        RECT 607.950 89.850 610.050 91.950 ;
        RECT 610.950 91.050 613.050 93.150 ;
        RECT 613.950 92.850 616.050 94.950 ;
        RECT 614.100 91.050 615.900 92.850 ;
        RECT 608.400 81.600 609.600 89.850 ;
        RECT 617.550 81.600 618.600 98.700 ;
        RECT 624.000 94.950 625.050 101.400 ;
        RECT 632.400 101.400 637.800 103.050 ;
        RECT 646.800 101.400 648.600 107.400 ;
        RECT 632.400 94.950 633.300 101.400 ;
        RECT 647.400 99.300 648.600 101.400 ;
        RECT 649.800 102.300 651.600 107.400 ;
        RECT 655.800 102.300 657.600 107.400 ;
        RECT 649.800 100.950 657.600 102.300 ;
        RECT 662.400 102.300 664.200 107.400 ;
        RECT 668.400 102.300 670.200 107.400 ;
        RECT 662.400 100.950 670.200 102.300 ;
        RECT 671.400 101.400 673.200 107.400 ;
        RECT 677.400 102.300 679.200 107.400 ;
        RECT 683.400 102.300 685.200 107.400 ;
        RECT 655.950 99.450 658.050 100.050 ;
        RECT 647.400 98.250 651.150 99.300 ;
        RECT 635.100 96.150 636.900 97.950 ;
        RECT 620.100 93.150 621.900 94.950 ;
        RECT 619.950 91.050 622.050 93.150 ;
        RECT 622.950 92.850 625.050 94.950 ;
        RECT 631.950 92.850 634.050 94.950 ;
        RECT 634.950 94.050 637.050 96.150 ;
        RECT 637.950 95.850 640.050 97.950 ;
        RECT 641.100 96.150 642.900 97.950 ;
        RECT 638.100 94.050 639.900 95.850 ;
        RECT 640.950 94.050 643.050 96.150 ;
        RECT 649.950 94.950 651.150 98.250 ;
        RECT 655.950 98.550 660.450 99.450 ;
        RECT 671.400 99.300 672.600 101.400 ;
        RECT 677.400 100.950 685.200 102.300 ;
        RECT 686.400 101.400 688.200 107.400 ;
        RECT 686.400 99.300 687.600 101.400 ;
        RECT 655.950 97.950 658.050 98.550 ;
        RECT 653.100 96.150 654.900 97.950 ;
        RECT 649.950 92.850 652.050 94.950 ;
        RECT 652.950 94.050 655.050 96.150 ;
        RECT 655.950 92.850 658.050 94.950 ;
        RECT 624.000 87.600 625.050 92.850 ;
        RECT 632.400 87.600 633.300 92.850 ;
        RECT 646.950 89.850 649.050 91.950 ;
        RECT 647.250 88.050 649.050 89.850 ;
        RECT 650.850 87.600 652.050 92.850 ;
        RECT 656.100 91.050 657.900 92.850 ;
        RECT 572.400 75.600 574.200 81.600 ;
        RECT 581.400 75.600 583.200 81.600 ;
        RECT 593.400 75.600 595.200 81.600 ;
        RECT 607.800 75.600 609.600 81.600 ;
        RECT 617.400 75.600 619.200 81.600 ;
        RECT 624.000 75.600 625.800 87.600 ;
        RECT 631.800 75.600 633.600 87.600 ;
        RECT 634.800 86.700 642.600 87.600 ;
        RECT 634.800 75.600 636.600 86.700 ;
        RECT 640.800 75.600 642.600 86.700 ;
        RECT 650.700 75.600 652.500 87.600 ;
        RECT 659.550 85.050 660.450 98.550 ;
        RECT 668.850 98.250 672.600 99.300 ;
        RECT 683.850 98.250 687.600 99.300 ;
        RECT 698.100 99.000 699.900 107.400 ;
        RECT 716.100 99.000 717.900 107.400 ;
        RECT 732.000 103.050 733.800 107.400 ;
        RECT 728.400 101.400 733.800 103.050 ;
        RECT 665.100 96.150 666.900 97.950 ;
        RECT 661.950 92.850 664.050 94.950 ;
        RECT 664.950 94.050 667.050 96.150 ;
        RECT 668.850 94.950 670.050 98.250 ;
        RECT 680.100 96.150 681.900 97.950 ;
        RECT 667.950 92.850 670.050 94.950 ;
        RECT 676.950 92.850 679.050 94.950 ;
        RECT 679.950 94.050 682.050 96.150 ;
        RECT 683.850 94.950 685.050 98.250 ;
        RECT 698.100 97.350 702.300 99.000 ;
        RECT 716.100 97.350 720.300 99.000 ;
        RECT 682.950 92.850 685.050 94.950 ;
        RECT 701.400 93.150 702.300 97.350 ;
        RECT 719.400 93.150 720.300 97.350 ;
        RECT 728.400 94.950 729.300 101.400 ;
        RECT 746.100 99.000 747.900 107.400 ;
        RECT 731.100 96.150 732.900 97.950 ;
        RECT 662.100 91.050 663.900 92.850 ;
        RECT 667.950 87.600 669.150 92.850 ;
        RECT 670.950 89.850 673.050 91.950 ;
        RECT 677.100 91.050 678.900 92.850 ;
        RECT 670.950 88.050 672.750 89.850 ;
        RECT 682.950 87.600 684.150 92.850 ;
        RECT 685.950 89.850 688.050 91.950 ;
        RECT 691.950 89.850 694.050 91.950 ;
        RECT 697.950 89.850 700.050 91.950 ;
        RECT 700.950 91.050 703.050 93.150 ;
        RECT 685.950 88.050 687.750 89.850 ;
        RECT 692.100 88.050 693.900 89.850 ;
        RECT 658.950 82.950 661.050 85.050 ;
        RECT 667.500 75.600 669.300 87.600 ;
        RECT 682.500 75.600 684.300 87.600 ;
        RECT 694.950 86.850 697.050 88.950 ;
        RECT 698.250 88.050 700.050 89.850 ;
        RECT 695.100 85.050 696.900 86.850 ;
        RECT 701.400 82.800 702.300 91.050 ;
        RECT 709.950 89.850 712.050 91.950 ;
        RECT 715.950 89.850 718.050 91.950 ;
        RECT 718.950 91.050 721.050 93.150 ;
        RECT 727.950 92.850 730.050 94.950 ;
        RECT 730.950 94.050 733.050 96.150 ;
        RECT 733.950 95.850 736.050 97.950 ;
        RECT 737.100 96.150 738.900 97.950 ;
        RECT 746.100 97.350 750.300 99.000 ;
        RECT 734.100 94.050 735.900 95.850 ;
        RECT 736.950 94.050 739.050 96.150 ;
        RECT 749.400 93.150 750.300 97.350 ;
        RECT 710.100 88.050 711.900 89.850 ;
        RECT 712.950 86.850 715.050 88.950 ;
        RECT 716.250 88.050 718.050 89.850 ;
        RECT 713.100 85.050 714.900 86.850 ;
        RECT 719.400 82.800 720.300 91.050 ;
        RECT 728.400 87.600 729.300 92.850 ;
        RECT 739.950 89.850 742.050 91.950 ;
        RECT 745.950 89.850 748.050 91.950 ;
        RECT 748.950 91.050 751.050 93.150 ;
        RECT 740.100 88.050 741.900 89.850 ;
        RECT 695.700 81.900 702.300 82.800 ;
        RECT 695.700 81.600 697.200 81.900 ;
        RECT 695.400 75.600 697.200 81.600 ;
        RECT 701.400 81.600 702.300 81.900 ;
        RECT 713.700 81.900 720.300 82.800 ;
        RECT 713.700 81.600 715.200 81.900 ;
        RECT 701.400 75.600 703.200 81.600 ;
        RECT 713.400 75.600 715.200 81.600 ;
        RECT 719.400 81.600 720.300 81.900 ;
        RECT 719.400 75.600 721.200 81.600 ;
        RECT 727.800 75.600 729.600 87.600 ;
        RECT 730.800 86.700 738.600 87.600 ;
        RECT 742.950 86.850 745.050 88.950 ;
        RECT 746.250 88.050 748.050 89.850 ;
        RECT 730.800 75.600 732.600 86.700 ;
        RECT 736.800 75.600 738.600 86.700 ;
        RECT 743.100 85.050 744.900 86.850 ;
        RECT 749.400 82.800 750.300 91.050 ;
        RECT 743.700 81.900 750.300 82.800 ;
        RECT 743.700 81.600 745.200 81.900 ;
        RECT 743.400 75.600 745.200 81.600 ;
        RECT 749.400 81.600 750.300 81.900 ;
        RECT 749.400 75.600 751.200 81.600 ;
        RECT 7.800 65.400 9.600 71.400 ;
        RECT 16.800 65.400 18.600 71.400 ;
        RECT 4.950 63.450 7.050 64.050 ;
        RECT 2.550 62.550 7.050 63.450 ;
        RECT 2.550 49.050 3.450 62.550 ;
        RECT 4.950 61.950 7.050 62.550 ;
        RECT 8.400 57.150 9.600 65.400 ;
        RECT 17.700 65.100 18.600 65.400 ;
        RECT 22.800 65.400 24.600 71.400 ;
        RECT 22.800 65.100 24.300 65.400 ;
        RECT 17.700 64.200 24.300 65.100 ;
        RECT 4.950 53.850 7.050 55.950 ;
        RECT 7.950 55.050 10.050 57.150 ;
        RECT 17.700 55.950 18.600 64.200 ;
        RECT 23.100 60.150 24.900 61.950 ;
        RECT 19.950 57.150 21.750 58.950 ;
        RECT 22.950 58.050 25.050 60.150 ;
        RECT 34.500 59.400 36.300 71.400 ;
        RECT 49.800 65.400 51.600 71.400 ;
        RECT 61.800 65.400 63.600 71.400 ;
        RECT 71.400 65.400 73.200 71.400 ;
        RECT 26.100 57.150 27.900 58.950 ;
        RECT 5.100 52.050 6.900 53.850 ;
        RECT 1.950 46.950 4.050 49.050 ;
        RECT 8.400 47.700 9.600 55.050 ;
        RECT 10.950 53.850 13.050 55.950 ;
        RECT 16.950 53.850 19.050 55.950 ;
        RECT 19.950 55.050 22.050 57.150 ;
        RECT 25.950 55.050 28.050 57.150 ;
        RECT 29.100 54.150 30.900 55.950 ;
        RECT 34.950 54.150 36.150 59.400 ;
        RECT 37.950 57.150 39.750 58.950 ;
        RECT 50.400 57.150 51.600 65.400 ;
        RECT 37.950 55.050 40.050 57.150 ;
        RECT 11.100 52.050 12.900 53.850 ;
        RECT 17.700 49.650 18.600 53.850 ;
        RECT 28.950 52.050 31.050 54.150 ;
        RECT 31.950 50.850 34.050 52.950 ;
        RECT 34.950 52.050 37.050 54.150 ;
        RECT 46.950 53.850 49.050 55.950 ;
        RECT 49.950 55.050 52.050 57.150 ;
        RECT 47.100 52.050 48.900 53.850 ;
        RECT 17.700 48.000 21.900 49.650 ;
        RECT 32.100 49.050 33.900 50.850 ;
        RECT 6.000 46.800 9.600 47.700 ;
        RECT 6.000 39.600 7.800 46.800 ;
        RECT 20.100 39.600 21.900 48.000 ;
        RECT 35.850 48.750 37.050 52.050 ;
        RECT 35.850 47.700 39.600 48.750 ;
        RECT 50.400 47.700 51.600 55.050 ;
        RECT 52.950 53.850 55.050 55.950 ;
        RECT 53.100 52.050 54.900 53.850 ;
        RECT 62.400 52.950 63.600 65.400 ;
        RECT 71.700 65.100 73.200 65.400 ;
        RECT 77.400 65.400 79.200 71.400 ;
        RECT 77.400 65.100 78.300 65.400 ;
        RECT 71.700 64.200 78.300 65.100 ;
        RECT 71.100 60.150 72.900 61.950 ;
        RECT 68.100 57.150 69.900 58.950 ;
        RECT 70.950 58.050 73.050 60.150 ;
        RECT 74.250 57.150 76.050 58.950 ;
        RECT 67.950 55.050 70.050 57.150 ;
        RECT 73.950 55.050 76.050 57.150 ;
        RECT 77.400 55.950 78.300 64.200 ;
        RECT 90.300 60.900 92.100 71.400 ;
        RECT 89.700 59.550 92.100 60.900 ;
        RECT 76.950 53.850 79.050 55.950 ;
        RECT 61.950 50.850 64.050 52.950 ;
        RECT 65.100 51.150 66.900 52.950 ;
        RECT 29.400 44.700 37.200 46.050 ;
        RECT 29.400 39.600 31.200 44.700 ;
        RECT 35.400 39.600 37.200 44.700 ;
        RECT 38.400 45.600 39.600 47.700 ;
        RECT 48.000 46.800 51.600 47.700 ;
        RECT 38.400 39.600 40.200 45.600 ;
        RECT 48.000 39.600 49.800 46.800 ;
        RECT 62.400 42.600 63.600 50.850 ;
        RECT 64.950 49.050 67.050 51.150 ;
        RECT 77.400 49.650 78.300 53.850 ;
        RECT 89.700 52.950 91.050 59.550 ;
        RECT 97.800 59.400 99.600 71.400 ;
        RECT 101.400 60.300 103.200 71.400 ;
        RECT 107.400 60.300 109.200 71.400 ;
        RECT 101.400 59.400 109.200 60.300 ;
        RECT 110.400 59.400 112.200 71.400 ;
        RECT 121.500 59.400 123.300 71.400 ;
        RECT 136.800 65.400 138.600 71.400 ;
        RECT 146.400 65.400 148.200 71.400 ;
        RECT 61.800 39.600 63.600 42.600 ;
        RECT 74.100 48.000 78.300 49.650 ;
        RECT 88.950 50.850 91.050 52.950 ;
        RECT 92.400 58.200 94.200 58.650 ;
        RECT 98.400 58.200 99.600 59.400 ;
        RECT 92.400 57.000 99.600 58.200 ;
        RECT 92.400 56.850 94.200 57.000 ;
        RECT 74.100 39.600 75.900 48.000 ;
        RECT 88.950 45.600 90.000 50.850 ;
        RECT 92.400 48.600 93.300 56.850 ;
        RECT 95.100 54.150 96.900 55.950 ;
        RECT 110.700 54.150 111.600 59.400 ;
        RECT 116.100 54.150 117.900 55.950 ;
        RECT 121.950 54.150 123.150 59.400 ;
        RECT 124.950 57.150 126.750 58.950 ;
        RECT 137.400 57.150 138.600 65.400 ;
        RECT 146.700 65.100 148.200 65.400 ;
        RECT 152.400 65.400 154.200 71.400 ;
        RECT 163.800 65.400 165.600 71.400 ;
        RECT 152.400 65.100 153.300 65.400 ;
        RECT 146.700 64.200 153.300 65.100 ;
        RECT 146.100 60.150 147.900 61.950 ;
        RECT 143.100 57.150 144.900 58.950 ;
        RECT 145.950 58.050 148.050 60.150 ;
        RECT 149.250 57.150 151.050 58.950 ;
        RECT 124.950 55.050 127.050 57.150 ;
        RECT 94.950 52.050 97.050 54.150 ;
        RECT 98.100 51.150 99.900 52.950 ;
        RECT 97.950 49.050 100.050 51.150 ;
        RECT 100.950 50.850 103.050 52.950 ;
        RECT 104.100 51.150 105.900 52.950 ;
        RECT 101.100 49.050 102.900 50.850 ;
        RECT 103.950 49.050 106.050 51.150 ;
        RECT 106.950 50.850 109.050 52.950 ;
        RECT 109.950 52.050 112.050 54.150 ;
        RECT 115.950 52.050 118.050 54.150 ;
        RECT 107.100 49.050 108.900 50.850 ;
        RECT 92.250 47.700 94.050 48.600 ;
        RECT 92.250 46.800 95.700 47.700 ;
        RECT 88.800 39.600 90.600 45.600 ;
        RECT 94.800 42.600 95.700 46.800 ;
        RECT 110.700 45.600 111.600 52.050 ;
        RECT 118.950 50.850 121.050 52.950 ;
        RECT 121.950 52.050 124.050 54.150 ;
        RECT 133.950 53.850 136.050 55.950 ;
        RECT 136.950 55.050 139.050 57.150 ;
        RECT 134.100 52.050 135.900 53.850 ;
        RECT 119.100 49.050 120.900 50.850 ;
        RECT 122.850 48.750 124.050 52.050 ;
        RECT 122.850 47.700 126.600 48.750 ;
        RECT 137.400 47.700 138.600 55.050 ;
        RECT 139.950 53.850 142.050 55.950 ;
        RECT 142.950 55.050 145.050 57.150 ;
        RECT 148.950 55.050 151.050 57.150 ;
        RECT 152.400 55.950 153.300 64.200 ;
        RECT 164.700 65.100 165.600 65.400 ;
        RECT 169.800 65.400 171.600 71.400 ;
        RECT 178.800 65.400 180.600 71.400 ;
        RECT 169.800 65.100 171.300 65.400 ;
        RECT 164.700 64.200 171.300 65.100 ;
        RECT 179.700 65.100 180.600 65.400 ;
        RECT 184.800 65.400 186.600 71.400 ;
        RECT 194.400 65.400 196.200 71.400 ;
        RECT 203.400 65.400 205.200 71.400 ;
        RECT 215.400 65.400 217.200 71.400 ;
        RECT 184.800 65.100 186.300 65.400 ;
        RECT 179.700 64.200 186.300 65.100 ;
        RECT 164.700 55.950 165.600 64.200 ;
        RECT 170.100 60.150 171.900 61.950 ;
        RECT 166.950 57.150 168.750 58.950 ;
        RECT 169.950 58.050 172.050 60.150 ;
        RECT 173.100 57.150 174.900 58.950 ;
        RECT 151.950 53.850 154.050 55.950 ;
        RECT 163.950 53.850 166.050 55.950 ;
        RECT 166.950 55.050 169.050 57.150 ;
        RECT 172.950 55.050 175.050 57.150 ;
        RECT 179.700 55.950 180.600 64.200 ;
        RECT 185.100 60.150 186.900 61.950 ;
        RECT 181.950 57.150 183.750 58.950 ;
        RECT 184.950 58.050 187.050 60.150 ;
        RECT 188.100 57.150 189.900 58.950 ;
        RECT 178.950 53.850 181.050 55.950 ;
        RECT 181.950 55.050 184.050 57.150 ;
        RECT 187.950 55.050 190.050 57.150 ;
        RECT 140.100 52.050 141.900 53.850 ;
        RECT 152.400 49.650 153.300 53.850 ;
        RECT 106.200 43.950 111.600 45.600 ;
        RECT 116.400 44.700 124.200 46.050 ;
        RECT 94.800 39.600 96.600 42.600 ;
        RECT 106.200 39.600 108.000 43.950 ;
        RECT 116.400 39.600 118.200 44.700 ;
        RECT 122.400 39.600 124.200 44.700 ;
        RECT 125.400 45.600 126.600 47.700 ;
        RECT 135.000 46.800 138.600 47.700 ;
        RECT 149.100 48.000 153.300 49.650 ;
        RECT 164.700 49.650 165.600 53.850 ;
        RECT 179.700 49.650 180.600 53.850 ;
        RECT 194.400 52.950 195.600 65.400 ;
        RECT 203.400 57.150 204.600 65.400 ;
        RECT 215.700 65.100 217.200 65.400 ;
        RECT 221.400 65.400 223.200 71.400 ;
        RECT 230.400 65.400 232.200 71.400 ;
        RECT 242.400 65.400 244.200 71.400 ;
        RECT 221.400 65.100 222.300 65.400 ;
        RECT 215.700 64.200 222.300 65.100 ;
        RECT 215.100 60.150 216.900 61.950 ;
        RECT 212.100 57.150 213.900 58.950 ;
        RECT 214.950 58.050 217.050 60.150 ;
        RECT 218.250 57.150 220.050 58.950 ;
        RECT 199.950 53.850 202.050 55.950 ;
        RECT 202.950 55.050 205.050 57.150 ;
        RECT 191.100 51.150 192.900 52.950 ;
        RECT 164.700 48.000 168.900 49.650 ;
        RECT 179.700 48.000 183.900 49.650 ;
        RECT 190.950 49.050 193.050 51.150 ;
        RECT 193.950 50.850 196.050 52.950 ;
        RECT 200.100 52.050 201.900 53.850 ;
        RECT 125.400 39.600 127.200 45.600 ;
        RECT 135.000 39.600 136.800 46.800 ;
        RECT 149.100 39.600 150.900 48.000 ;
        RECT 167.100 39.600 168.900 48.000 ;
        RECT 182.100 39.600 183.900 48.000 ;
        RECT 194.400 42.600 195.600 50.850 ;
        RECT 203.400 47.700 204.600 55.050 ;
        RECT 205.950 53.850 208.050 55.950 ;
        RECT 211.950 55.050 214.050 57.150 ;
        RECT 217.950 55.050 220.050 57.150 ;
        RECT 221.400 55.950 222.300 64.200 ;
        RECT 230.400 57.150 231.600 65.400 ;
        RECT 220.950 53.850 223.050 55.950 ;
        RECT 226.950 53.850 229.050 55.950 ;
        RECT 229.950 55.050 232.050 57.150 ;
        RECT 206.100 52.050 207.900 53.850 ;
        RECT 221.400 49.650 222.300 53.850 ;
        RECT 227.100 52.050 228.900 53.850 ;
        RECT 218.100 48.000 222.300 49.650 ;
        RECT 203.400 46.800 207.000 47.700 ;
        RECT 194.400 39.600 196.200 42.600 ;
        RECT 205.200 39.600 207.000 46.800 ;
        RECT 218.100 39.600 219.900 48.000 ;
        RECT 230.400 47.700 231.600 55.050 ;
        RECT 232.950 53.850 235.050 55.950 ;
        RECT 239.100 54.150 240.900 55.950 ;
        RECT 233.100 52.050 234.900 53.850 ;
        RECT 238.950 52.050 241.050 54.150 ;
        RECT 242.550 48.300 243.600 65.400 ;
        RECT 249.000 59.400 250.800 71.400 ;
        RECT 262.800 65.400 264.600 71.400 ;
        RECT 244.950 53.850 247.050 55.950 ;
        RECT 249.000 54.150 250.050 59.400 ;
        RECT 263.400 57.150 264.600 65.400 ;
        RECT 276.600 59.400 278.400 71.400 ;
        RECT 286.800 65.400 288.600 71.400 ;
        RECT 276.000 58.350 278.400 59.400 ;
        RECT 287.700 65.100 288.600 65.400 ;
        RECT 292.800 65.400 294.600 71.400 ;
        RECT 292.800 65.100 294.300 65.400 ;
        RECT 287.700 64.200 294.300 65.100 ;
        RECT 245.100 52.050 246.900 53.850 ;
        RECT 247.950 52.050 250.050 54.150 ;
        RECT 259.950 53.850 262.050 55.950 ;
        RECT 262.950 55.050 265.050 57.150 ;
        RECT 260.100 52.050 261.900 53.850 ;
        RECT 230.400 46.800 234.000 47.700 ;
        RECT 232.200 39.600 234.000 46.800 ;
        RECT 239.400 47.100 246.900 48.300 ;
        RECT 239.400 39.600 241.200 47.100 ;
        RECT 245.100 46.500 246.900 47.100 ;
        RECT 249.000 45.600 250.050 52.050 ;
        RECT 263.400 47.700 264.600 55.050 ;
        RECT 265.950 53.850 268.050 55.950 ;
        RECT 272.100 54.150 273.900 55.950 ;
        RECT 266.100 52.050 267.900 53.850 ;
        RECT 271.950 52.050 274.050 54.150 ;
        RECT 276.000 51.150 277.050 58.350 ;
        RECT 287.700 55.950 288.600 64.200 ;
        RECT 293.100 60.150 294.900 61.950 ;
        RECT 289.950 57.150 291.750 58.950 ;
        RECT 292.950 58.050 295.050 60.150 ;
        RECT 305.700 59.400 307.500 71.400 ;
        RECT 317.400 60.300 319.200 71.400 ;
        RECT 323.400 60.300 325.200 71.400 ;
        RECT 317.400 59.400 325.200 60.300 ;
        RECT 326.400 59.400 328.200 71.400 ;
        RECT 334.800 65.400 336.600 71.400 ;
        RECT 335.700 65.100 336.600 65.400 ;
        RECT 340.800 65.400 342.600 71.400 ;
        RECT 353.400 65.400 355.200 71.400 ;
        RECT 340.800 65.100 342.300 65.400 ;
        RECT 335.700 64.200 342.300 65.100 ;
        RECT 353.700 65.100 355.200 65.400 ;
        RECT 359.400 65.400 361.200 71.400 ;
        RECT 367.800 65.400 369.600 71.400 ;
        RECT 377.400 65.400 379.200 71.400 ;
        RECT 359.400 65.100 360.300 65.400 ;
        RECT 353.700 64.200 360.300 65.100 ;
        RECT 296.100 57.150 297.900 58.950 ;
        RECT 302.250 57.150 304.050 58.950 ;
        RECT 278.100 54.150 279.900 55.950 ;
        RECT 277.950 52.050 280.050 54.150 ;
        RECT 286.950 53.850 289.050 55.950 ;
        RECT 289.950 55.050 292.050 57.150 ;
        RECT 295.950 55.050 298.050 57.150 ;
        RECT 301.950 55.050 304.050 57.150 ;
        RECT 305.850 54.150 307.050 59.400 ;
        RECT 311.100 54.150 312.900 55.950 ;
        RECT 326.700 54.150 327.600 59.400 ;
        RECT 335.700 55.950 336.600 64.200 ;
        RECT 341.100 60.150 342.900 61.950 ;
        RECT 353.100 60.150 354.900 61.950 ;
        RECT 337.950 57.150 339.750 58.950 ;
        RECT 340.950 58.050 343.050 60.150 ;
        RECT 344.100 57.150 345.900 58.950 ;
        RECT 350.100 57.150 351.900 58.950 ;
        RECT 352.950 58.050 355.050 60.150 ;
        RECT 356.250 57.150 358.050 58.950 ;
        RECT 274.950 49.050 277.050 51.150 ;
        RECT 246.900 44.100 250.050 45.600 ;
        RECT 261.000 46.800 264.600 47.700 ;
        RECT 246.900 39.600 248.700 44.100 ;
        RECT 261.000 39.600 262.800 46.800 ;
        RECT 276.000 42.600 277.050 49.050 ;
        RECT 287.700 49.650 288.600 53.850 ;
        RECT 304.950 52.050 307.050 54.150 ;
        RECT 287.700 48.000 291.900 49.650 ;
        RECT 304.950 48.750 306.150 52.050 ;
        RECT 307.950 50.850 310.050 52.950 ;
        RECT 310.950 52.050 313.050 54.150 ;
        RECT 316.950 50.850 319.050 52.950 ;
        RECT 320.100 51.150 321.900 52.950 ;
        RECT 308.100 49.050 309.900 50.850 ;
        RECT 317.100 49.050 318.900 50.850 ;
        RECT 319.950 49.050 322.050 51.150 ;
        RECT 322.950 50.850 325.050 52.950 ;
        RECT 325.950 52.050 328.050 54.150 ;
        RECT 334.950 53.850 337.050 55.950 ;
        RECT 337.950 55.050 340.050 57.150 ;
        RECT 343.950 55.050 346.050 57.150 ;
        RECT 349.950 55.050 352.050 57.150 ;
        RECT 355.950 55.050 358.050 57.150 ;
        RECT 359.400 55.950 360.300 64.200 ;
        RECT 358.950 53.850 361.050 55.950 ;
        RECT 323.100 49.050 324.900 50.850 ;
        RECT 275.400 39.600 277.200 42.600 ;
        RECT 290.100 39.600 291.900 48.000 ;
        RECT 302.400 47.700 306.150 48.750 ;
        RECT 302.400 45.600 303.600 47.700 ;
        RECT 301.800 39.600 303.600 45.600 ;
        RECT 304.800 44.700 312.600 46.050 ;
        RECT 326.700 45.600 327.600 52.050 ;
        RECT 335.700 49.650 336.600 53.850 ;
        RECT 359.400 49.650 360.300 53.850 ;
        RECT 368.400 52.950 369.600 65.400 ;
        RECT 377.700 65.100 379.200 65.400 ;
        RECT 383.400 65.400 385.200 71.400 ;
        RECT 392.400 65.400 394.200 71.400 ;
        RECT 383.400 65.100 384.300 65.400 ;
        RECT 377.700 64.200 384.300 65.100 ;
        RECT 392.700 65.100 394.200 65.400 ;
        RECT 398.400 65.400 400.200 71.400 ;
        RECT 398.400 65.100 399.300 65.400 ;
        RECT 392.700 64.200 399.300 65.100 ;
        RECT 377.100 60.150 378.900 61.950 ;
        RECT 374.100 57.150 375.900 58.950 ;
        RECT 376.950 58.050 379.050 60.150 ;
        RECT 380.250 57.150 382.050 58.950 ;
        RECT 373.950 55.050 376.050 57.150 ;
        RECT 379.950 55.050 382.050 57.150 ;
        RECT 383.400 55.950 384.300 64.200 ;
        RECT 385.950 58.950 388.050 61.050 ;
        RECT 392.100 60.150 393.900 61.950 ;
        RECT 382.950 53.850 385.050 55.950 ;
        RECT 367.950 50.850 370.050 52.950 ;
        RECT 371.100 51.150 372.900 52.950 ;
        RECT 335.700 48.000 339.900 49.650 ;
        RECT 304.800 39.600 306.600 44.700 ;
        RECT 310.800 39.600 312.600 44.700 ;
        RECT 322.200 43.950 327.600 45.600 ;
        RECT 322.200 39.600 324.000 43.950 ;
        RECT 338.100 39.600 339.900 48.000 ;
        RECT 356.100 48.000 360.300 49.650 ;
        RECT 356.100 39.600 357.900 48.000 ;
        RECT 368.400 42.600 369.600 50.850 ;
        RECT 370.950 49.050 373.050 51.150 ;
        RECT 383.400 49.650 384.300 53.850 ;
        RECT 386.550 51.450 387.450 58.950 ;
        RECT 389.100 57.150 390.900 58.950 ;
        RECT 391.950 58.050 394.050 60.150 ;
        RECT 395.250 57.150 397.050 58.950 ;
        RECT 388.950 55.050 391.050 57.150 ;
        RECT 394.950 55.050 397.050 57.150 ;
        RECT 398.400 55.950 399.300 64.200 ;
        RECT 412.500 59.400 414.300 71.400 ;
        RECT 422.400 60.300 424.200 71.400 ;
        RECT 428.400 60.300 430.200 71.400 ;
        RECT 422.400 59.400 430.200 60.300 ;
        RECT 431.400 59.400 433.200 71.400 ;
        RECT 442.500 59.400 444.300 71.400 ;
        RECT 455.400 65.400 457.200 71.400 ;
        RECT 455.700 65.100 457.200 65.400 ;
        RECT 461.400 65.400 463.200 71.400 ;
        RECT 469.800 65.400 471.600 71.400 ;
        RECT 461.400 65.100 462.300 65.400 ;
        RECT 455.700 64.200 462.300 65.100 ;
        RECT 455.100 60.150 456.900 61.950 ;
        RECT 397.950 53.850 400.050 55.950 ;
        RECT 407.100 54.150 408.900 55.950 ;
        RECT 412.950 54.150 414.150 59.400 ;
        RECT 415.950 57.150 417.750 58.950 ;
        RECT 415.950 55.050 418.050 57.150 ;
        RECT 431.700 54.150 432.600 59.400 ;
        RECT 437.100 54.150 438.900 55.950 ;
        RECT 442.950 54.150 444.150 59.400 ;
        RECT 445.950 57.150 447.750 58.950 ;
        RECT 452.100 57.150 453.900 58.950 ;
        RECT 454.950 58.050 457.050 60.150 ;
        RECT 458.250 57.150 460.050 58.950 ;
        RECT 445.950 55.050 448.050 57.150 ;
        RECT 451.950 55.050 454.050 57.150 ;
        RECT 457.950 55.050 460.050 57.150 ;
        RECT 461.400 55.950 462.300 64.200 ;
        RECT 470.700 65.100 471.600 65.400 ;
        RECT 475.800 65.400 477.600 71.400 ;
        RECT 488.400 65.400 490.200 71.400 ;
        RECT 475.800 65.100 477.300 65.400 ;
        RECT 470.700 64.200 477.300 65.100 ;
        RECT 488.700 65.100 490.200 65.400 ;
        RECT 494.400 65.400 496.200 71.400 ;
        RECT 494.400 65.100 495.300 65.400 ;
        RECT 488.700 64.200 495.300 65.100 ;
        RECT 470.700 55.950 471.600 64.200 ;
        RECT 476.100 60.150 477.900 61.950 ;
        RECT 488.100 60.150 489.900 61.950 ;
        RECT 472.950 57.150 474.750 58.950 ;
        RECT 475.950 58.050 478.050 60.150 ;
        RECT 479.100 57.150 480.900 58.950 ;
        RECT 485.100 57.150 486.900 58.950 ;
        RECT 487.950 58.050 490.050 60.150 ;
        RECT 491.250 57.150 493.050 58.950 ;
        RECT 391.950 51.450 394.050 52.050 ;
        RECT 386.550 50.550 394.050 51.450 ;
        RECT 391.950 49.950 394.050 50.550 ;
        RECT 398.400 49.650 399.300 53.850 ;
        RECT 406.950 52.050 409.050 54.150 ;
        RECT 409.950 50.850 412.050 52.950 ;
        RECT 412.950 52.050 415.050 54.150 ;
        RECT 367.800 39.600 369.600 42.600 ;
        RECT 380.100 48.000 384.300 49.650 ;
        RECT 395.100 48.000 399.300 49.650 ;
        RECT 410.100 49.050 411.900 50.850 ;
        RECT 413.850 48.750 415.050 52.050 ;
        RECT 421.950 50.850 424.050 52.950 ;
        RECT 425.100 51.150 426.900 52.950 ;
        RECT 422.100 49.050 423.900 50.850 ;
        RECT 424.950 49.050 427.050 51.150 ;
        RECT 427.950 50.850 430.050 52.950 ;
        RECT 430.950 52.050 433.050 54.150 ;
        RECT 436.950 52.050 439.050 54.150 ;
        RECT 428.100 49.050 429.900 50.850 ;
        RECT 380.100 39.600 381.900 48.000 ;
        RECT 395.100 39.600 396.900 48.000 ;
        RECT 413.850 47.700 417.600 48.750 ;
        RECT 407.400 44.700 415.200 46.050 ;
        RECT 407.400 39.600 409.200 44.700 ;
        RECT 413.400 39.600 415.200 44.700 ;
        RECT 416.400 45.600 417.600 47.700 ;
        RECT 431.700 45.600 432.600 52.050 ;
        RECT 439.950 50.850 442.050 52.950 ;
        RECT 442.950 52.050 445.050 54.150 ;
        RECT 460.950 53.850 463.050 55.950 ;
        RECT 469.950 53.850 472.050 55.950 ;
        RECT 472.950 55.050 475.050 57.150 ;
        RECT 478.950 55.050 481.050 57.150 ;
        RECT 484.950 55.050 487.050 57.150 ;
        RECT 490.950 55.050 493.050 57.150 ;
        RECT 494.400 55.950 495.300 64.200 ;
        RECT 500.400 60.300 502.200 71.400 ;
        RECT 506.400 60.300 508.200 71.400 ;
        RECT 500.400 59.400 508.200 60.300 ;
        RECT 509.400 59.400 511.200 71.400 ;
        RECT 518.400 65.400 520.200 71.400 ;
        RECT 518.700 65.100 520.200 65.400 ;
        RECT 524.400 65.400 526.200 71.400 ;
        RECT 524.400 65.100 525.300 65.400 ;
        RECT 518.700 64.200 525.300 65.100 ;
        RECT 518.100 60.150 519.900 61.950 ;
        RECT 493.950 53.850 496.050 55.950 ;
        RECT 509.700 54.150 510.600 59.400 ;
        RECT 515.100 57.150 516.900 58.950 ;
        RECT 517.950 58.050 520.050 60.150 ;
        RECT 521.250 57.150 523.050 58.950 ;
        RECT 514.950 55.050 517.050 57.150 ;
        RECT 520.950 55.050 523.050 57.150 ;
        RECT 524.400 55.950 525.300 64.200 ;
        RECT 535.500 59.400 537.300 71.400 ;
        RECT 548.400 65.400 550.200 71.400 ;
        RECT 548.700 65.100 550.200 65.400 ;
        RECT 554.400 65.400 556.200 71.400 ;
        RECT 554.400 65.100 555.300 65.400 ;
        RECT 548.700 64.200 555.300 65.100 ;
        RECT 544.950 63.450 547.050 64.050 ;
        RECT 542.550 62.550 547.050 63.450 ;
        RECT 440.100 49.050 441.900 50.850 ;
        RECT 443.850 48.750 445.050 52.050 ;
        RECT 461.400 49.650 462.300 53.850 ;
        RECT 443.850 47.700 447.600 48.750 ;
        RECT 416.400 39.600 418.200 45.600 ;
        RECT 427.200 43.950 432.600 45.600 ;
        RECT 437.400 44.700 445.200 46.050 ;
        RECT 427.200 39.600 429.000 43.950 ;
        RECT 437.400 39.600 439.200 44.700 ;
        RECT 443.400 39.600 445.200 44.700 ;
        RECT 446.400 45.600 447.600 47.700 ;
        RECT 458.100 48.000 462.300 49.650 ;
        RECT 470.700 49.650 471.600 53.850 ;
        RECT 475.950 51.450 478.050 52.050 ;
        RECT 487.950 51.450 490.050 52.050 ;
        RECT 475.950 50.550 490.050 51.450 ;
        RECT 475.950 49.950 478.050 50.550 ;
        RECT 487.950 49.950 490.050 50.550 ;
        RECT 494.400 49.650 495.300 53.850 ;
        RECT 499.950 50.850 502.050 52.950 ;
        RECT 503.100 51.150 504.900 52.950 ;
        RECT 470.700 48.000 474.900 49.650 ;
        RECT 446.400 39.600 448.200 45.600 ;
        RECT 458.100 39.600 459.900 48.000 ;
        RECT 473.100 39.600 474.900 48.000 ;
        RECT 491.100 48.000 495.300 49.650 ;
        RECT 500.100 49.050 501.900 50.850 ;
        RECT 502.950 49.050 505.050 51.150 ;
        RECT 505.950 50.850 508.050 52.950 ;
        RECT 508.950 52.050 511.050 54.150 ;
        RECT 523.950 53.850 526.050 55.950 ;
        RECT 530.100 54.150 531.900 55.950 ;
        RECT 535.950 54.150 537.150 59.400 ;
        RECT 538.950 57.150 540.750 58.950 ;
        RECT 538.950 55.050 541.050 57.150 ;
        RECT 506.100 49.050 507.900 50.850 ;
        RECT 491.100 39.600 492.900 48.000 ;
        RECT 509.700 45.600 510.600 52.050 ;
        RECT 524.400 49.650 525.300 53.850 ;
        RECT 529.950 52.050 532.050 54.150 ;
        RECT 532.950 50.850 535.050 52.950 ;
        RECT 535.950 52.050 538.050 54.150 ;
        RECT 505.200 43.950 510.600 45.600 ;
        RECT 521.100 48.000 525.300 49.650 ;
        RECT 533.100 49.050 534.900 50.850 ;
        RECT 536.850 48.750 538.050 52.050 ;
        RECT 538.950 51.450 541.050 52.050 ;
        RECT 542.550 51.450 543.450 62.550 ;
        RECT 544.950 61.950 547.050 62.550 ;
        RECT 548.100 60.150 549.900 61.950 ;
        RECT 545.100 57.150 546.900 58.950 ;
        RECT 547.950 58.050 550.050 60.150 ;
        RECT 551.250 57.150 553.050 58.950 ;
        RECT 544.950 55.050 547.050 57.150 ;
        RECT 550.950 55.050 553.050 57.150 ;
        RECT 554.400 55.950 555.300 64.200 ;
        RECT 565.500 59.400 567.300 71.400 ;
        RECT 581.400 65.400 583.200 71.400 ;
        RECT 553.950 53.850 556.050 55.950 ;
        RECT 560.100 54.150 561.900 55.950 ;
        RECT 565.950 54.150 567.150 59.400 ;
        RECT 568.950 57.150 570.750 58.950 ;
        RECT 581.400 57.150 582.600 65.400 ;
        RECT 583.950 60.450 586.050 61.050 ;
        RECT 583.950 59.550 588.450 60.450 ;
        RECT 583.950 58.950 586.050 59.550 ;
        RECT 568.950 55.050 571.050 57.150 ;
        RECT 538.950 50.550 543.450 51.450 ;
        RECT 538.950 49.950 541.050 50.550 ;
        RECT 554.400 49.650 555.300 53.850 ;
        RECT 559.950 52.050 562.050 54.150 ;
        RECT 562.950 50.850 565.050 52.950 ;
        RECT 565.950 52.050 568.050 54.150 ;
        RECT 577.950 53.850 580.050 55.950 ;
        RECT 580.950 55.050 583.050 57.150 ;
        RECT 578.100 52.050 579.900 53.850 ;
        RECT 505.200 39.600 507.000 43.950 ;
        RECT 521.100 39.600 522.900 48.000 ;
        RECT 536.850 47.700 540.600 48.750 ;
        RECT 530.400 44.700 538.200 46.050 ;
        RECT 530.400 39.600 532.200 44.700 ;
        RECT 536.400 39.600 538.200 44.700 ;
        RECT 539.400 45.600 540.600 47.700 ;
        RECT 551.100 48.000 555.300 49.650 ;
        RECT 563.100 49.050 564.900 50.850 ;
        RECT 566.850 48.750 568.050 52.050 ;
        RECT 539.400 39.600 541.200 45.600 ;
        RECT 551.100 39.600 552.900 48.000 ;
        RECT 566.850 47.700 570.600 48.750 ;
        RECT 560.400 44.700 568.200 46.050 ;
        RECT 560.400 39.600 562.200 44.700 ;
        RECT 566.400 39.600 568.200 44.700 ;
        RECT 569.400 45.600 570.600 47.700 ;
        RECT 581.400 47.700 582.600 55.050 ;
        RECT 583.950 53.850 586.050 55.950 ;
        RECT 584.100 52.050 585.900 53.850 ;
        RECT 587.550 49.050 588.450 59.550 ;
        RECT 594.600 59.400 596.400 71.400 ;
        RECT 594.000 58.350 596.400 59.400 ;
        RECT 609.600 59.400 611.400 71.400 ;
        RECT 623.700 59.400 625.500 71.400 ;
        RECT 638.400 65.400 640.200 71.400 ;
        RECT 650.400 65.400 652.200 71.400 ;
        RECT 609.600 58.350 612.000 59.400 ;
        RECT 590.100 54.150 591.900 55.950 ;
        RECT 589.950 52.050 592.050 54.150 ;
        RECT 594.000 51.150 595.050 58.350 ;
        RECT 596.100 54.150 597.900 55.950 ;
        RECT 608.100 54.150 609.900 55.950 ;
        RECT 595.950 52.050 598.050 54.150 ;
        RECT 607.950 52.050 610.050 54.150 ;
        RECT 592.950 49.050 595.050 51.150 ;
        RECT 581.400 46.800 585.000 47.700 ;
        RECT 586.950 46.950 589.050 49.050 ;
        RECT 569.400 39.600 571.200 45.600 ;
        RECT 583.200 39.600 585.000 46.800 ;
        RECT 594.000 42.600 595.050 49.050 ;
        RECT 610.950 51.150 612.000 58.350 ;
        RECT 620.250 57.150 622.050 58.950 ;
        RECT 614.100 54.150 615.900 55.950 ;
        RECT 619.950 55.050 622.050 57.150 ;
        RECT 623.850 54.150 625.050 59.400 ;
        RECT 638.400 57.150 639.600 65.400 ;
        RECT 629.100 54.150 630.900 55.950 ;
        RECT 613.950 52.050 616.050 54.150 ;
        RECT 622.950 52.050 625.050 54.150 ;
        RECT 610.950 49.050 613.050 51.150 ;
        RECT 610.950 42.600 612.000 49.050 ;
        RECT 622.950 48.750 624.150 52.050 ;
        RECT 625.950 50.850 628.050 52.950 ;
        RECT 628.950 52.050 631.050 54.150 ;
        RECT 634.950 53.850 637.050 55.950 ;
        RECT 637.950 55.050 640.050 57.150 ;
        RECT 635.100 52.050 636.900 53.850 ;
        RECT 626.100 49.050 627.900 50.850 ;
        RECT 620.400 47.700 624.150 48.750 ;
        RECT 638.400 47.700 639.600 55.050 ;
        RECT 640.950 53.850 643.050 55.950 ;
        RECT 641.100 52.050 642.900 53.850 ;
        RECT 650.400 52.950 651.600 65.400 ;
        RECT 661.500 59.400 663.300 71.400 ;
        RECT 673.800 59.400 675.600 71.400 ;
        RECT 676.800 60.300 678.600 71.400 ;
        RECT 682.800 60.300 684.600 71.400 ;
        RECT 676.800 59.400 684.600 60.300 ;
        RECT 688.800 59.400 690.600 71.400 ;
        RECT 691.800 60.300 693.600 71.400 ;
        RECT 697.800 60.300 699.600 71.400 ;
        RECT 704.400 65.400 706.200 71.400 ;
        RECT 704.700 65.100 706.200 65.400 ;
        RECT 710.400 65.400 712.200 71.400 ;
        RECT 721.800 65.400 723.600 71.400 ;
        RECT 710.400 65.100 711.300 65.400 ;
        RECT 704.700 64.200 711.300 65.100 ;
        RECT 691.800 59.400 699.600 60.300 ;
        RECT 704.100 60.150 705.900 61.950 ;
        RECT 656.100 54.150 657.900 55.950 ;
        RECT 661.950 54.150 663.150 59.400 ;
        RECT 664.950 57.150 666.750 58.950 ;
        RECT 664.950 55.050 667.050 57.150 ;
        RECT 674.400 54.150 675.300 59.400 ;
        RECT 689.400 54.150 690.300 59.400 ;
        RECT 701.100 57.150 702.900 58.950 ;
        RECT 703.950 58.050 706.050 60.150 ;
        RECT 707.250 57.150 709.050 58.950 ;
        RECT 700.950 55.050 703.050 57.150 ;
        RECT 706.950 55.050 709.050 57.150 ;
        RECT 710.400 55.950 711.300 64.200 ;
        RECT 722.700 65.100 723.600 65.400 ;
        RECT 727.800 65.400 729.600 71.400 ;
        RECT 737.400 65.400 739.200 71.400 ;
        RECT 727.800 65.100 729.300 65.400 ;
        RECT 722.700 64.200 729.300 65.100 ;
        RECT 737.700 65.100 739.200 65.400 ;
        RECT 743.400 65.400 745.200 71.400 ;
        RECT 743.400 65.100 744.300 65.400 ;
        RECT 737.700 64.200 744.300 65.100 ;
        RECT 722.700 55.950 723.600 64.200 ;
        RECT 728.100 60.150 729.900 61.950 ;
        RECT 737.100 60.150 738.900 61.950 ;
        RECT 724.950 57.150 726.750 58.950 ;
        RECT 727.950 58.050 730.050 60.150 ;
        RECT 731.100 57.150 732.900 58.950 ;
        RECT 734.100 57.150 735.900 58.950 ;
        RECT 736.950 58.050 739.050 60.150 ;
        RECT 740.250 57.150 742.050 58.950 ;
        RECT 647.100 51.150 648.900 52.950 ;
        RECT 646.950 49.050 649.050 51.150 ;
        RECT 649.950 50.850 652.050 52.950 ;
        RECT 655.950 52.050 658.050 54.150 ;
        RECT 658.950 50.850 661.050 52.950 ;
        RECT 661.950 52.050 664.050 54.150 ;
        RECT 673.950 52.050 676.050 54.150 ;
        RECT 620.400 45.600 621.600 47.700 ;
        RECT 638.400 46.800 642.000 47.700 ;
        RECT 593.400 39.600 595.200 42.600 ;
        RECT 610.800 39.600 612.600 42.600 ;
        RECT 619.800 39.600 621.600 45.600 ;
        RECT 622.800 44.700 630.600 46.050 ;
        RECT 622.800 39.600 624.600 44.700 ;
        RECT 628.800 39.600 630.600 44.700 ;
        RECT 640.200 39.600 642.000 46.800 ;
        RECT 650.400 42.600 651.600 50.850 ;
        RECT 659.100 49.050 660.900 50.850 ;
        RECT 662.850 48.750 664.050 52.050 ;
        RECT 662.850 47.700 666.600 48.750 ;
        RECT 656.400 44.700 664.200 46.050 ;
        RECT 650.400 39.600 652.200 42.600 ;
        RECT 656.400 39.600 658.200 44.700 ;
        RECT 662.400 39.600 664.200 44.700 ;
        RECT 665.400 45.600 666.600 47.700 ;
        RECT 674.400 45.600 675.300 52.050 ;
        RECT 676.950 50.850 679.050 52.950 ;
        RECT 680.100 51.150 681.900 52.950 ;
        RECT 677.100 49.050 678.900 50.850 ;
        RECT 679.950 49.050 682.050 51.150 ;
        RECT 682.950 50.850 685.050 52.950 ;
        RECT 688.950 52.050 691.050 54.150 ;
        RECT 709.950 53.850 712.050 55.950 ;
        RECT 721.950 53.850 724.050 55.950 ;
        RECT 724.950 55.050 727.050 57.150 ;
        RECT 730.950 55.050 733.050 57.150 ;
        RECT 733.950 55.050 736.050 57.150 ;
        RECT 739.950 55.050 742.050 57.150 ;
        RECT 743.400 55.950 744.300 64.200 ;
        RECT 749.400 60.300 751.200 71.400 ;
        RECT 755.400 60.300 757.200 71.400 ;
        RECT 749.400 59.400 757.200 60.300 ;
        RECT 758.400 59.400 760.200 71.400 ;
        RECT 742.950 53.850 745.050 55.950 ;
        RECT 758.700 54.150 759.600 59.400 ;
        RECT 683.100 49.050 684.900 50.850 ;
        RECT 689.400 45.600 690.300 52.050 ;
        RECT 691.950 50.850 694.050 52.950 ;
        RECT 695.100 51.150 696.900 52.950 ;
        RECT 692.100 49.050 693.900 50.850 ;
        RECT 694.950 49.050 697.050 51.150 ;
        RECT 697.950 50.850 700.050 52.950 ;
        RECT 698.100 49.050 699.900 50.850 ;
        RECT 710.400 49.650 711.300 53.850 ;
        RECT 707.100 48.000 711.300 49.650 ;
        RECT 722.700 49.650 723.600 53.850 ;
        RECT 743.400 49.650 744.300 53.850 ;
        RECT 748.950 50.850 751.050 52.950 ;
        RECT 752.100 51.150 753.900 52.950 ;
        RECT 722.700 48.000 726.900 49.650 ;
        RECT 665.400 39.600 667.200 45.600 ;
        RECT 674.400 43.950 679.800 45.600 ;
        RECT 689.400 43.950 694.800 45.600 ;
        RECT 678.000 39.600 679.800 43.950 ;
        RECT 693.000 39.600 694.800 43.950 ;
        RECT 707.100 39.600 708.900 48.000 ;
        RECT 725.100 39.600 726.900 48.000 ;
        RECT 740.100 48.000 744.300 49.650 ;
        RECT 749.100 49.050 750.900 50.850 ;
        RECT 751.950 49.050 754.050 51.150 ;
        RECT 754.950 50.850 757.050 52.950 ;
        RECT 757.950 52.050 760.050 54.150 ;
        RECT 755.100 49.050 756.900 50.850 ;
        RECT 740.100 39.600 741.900 48.000 ;
        RECT 758.700 45.600 759.600 52.050 ;
        RECT 754.200 43.950 759.600 45.600 ;
        RECT 754.200 39.600 756.000 43.950 ;
        RECT 7.800 32.400 9.600 35.400 ;
        RECT 7.950 25.950 9.000 32.400 ;
        RECT 14.400 27.900 16.200 35.400 ;
        RECT 21.900 30.900 23.700 35.400 ;
        RECT 21.900 29.400 25.050 30.900 ;
        RECT 20.100 27.900 21.900 28.500 ;
        RECT 14.400 26.700 21.900 27.900 ;
        RECT 7.950 23.850 10.050 25.950 ;
        RECT 4.950 20.850 7.050 22.950 ;
        RECT 5.100 19.050 6.900 20.850 ;
        RECT 7.950 16.650 9.000 23.850 ;
        RECT 10.950 20.850 13.050 22.950 ;
        RECT 13.950 20.850 16.050 22.950 ;
        RECT 11.100 19.050 12.900 20.850 ;
        RECT 14.100 19.050 15.900 20.850 ;
        RECT 6.600 15.600 9.000 16.650 ;
        RECT 6.600 3.600 8.400 15.600 ;
        RECT 17.550 9.600 18.600 26.700 ;
        RECT 24.000 22.950 25.050 29.400 ;
        RECT 32.400 30.300 34.200 35.400 ;
        RECT 38.400 30.300 40.200 35.400 ;
        RECT 32.400 28.950 40.200 30.300 ;
        RECT 41.400 29.400 43.200 35.400 ;
        RECT 51.300 30.900 53.100 35.400 ;
        RECT 49.950 29.400 53.100 30.900 ;
        RECT 41.400 27.300 42.600 29.400 ;
        RECT 38.850 26.250 42.600 27.300 ;
        RECT 35.100 24.150 36.900 25.950 ;
        RECT 20.100 21.150 21.900 22.950 ;
        RECT 19.950 19.050 22.050 21.150 ;
        RECT 22.950 20.850 25.050 22.950 ;
        RECT 31.950 20.850 34.050 22.950 ;
        RECT 34.950 22.050 37.050 24.150 ;
        RECT 38.850 22.950 40.050 26.250 ;
        RECT 37.950 20.850 40.050 22.950 ;
        RECT 49.950 22.950 51.000 29.400 ;
        RECT 53.100 27.900 54.900 28.500 ;
        RECT 58.800 27.900 60.600 35.400 ;
        RECT 53.100 26.700 60.600 27.900 ;
        RECT 66.000 28.200 67.800 35.400 ;
        RECT 79.200 29.400 81.000 35.400 ;
        RECT 66.000 27.300 69.600 28.200 ;
        RECT 49.950 20.850 52.050 22.950 ;
        RECT 53.100 21.150 54.900 22.950 ;
        RECT 24.000 15.600 25.050 20.850 ;
        RECT 32.100 19.050 33.900 20.850 ;
        RECT 37.950 15.600 39.150 20.850 ;
        RECT 40.950 17.850 43.050 19.950 ;
        RECT 40.950 16.050 42.750 17.850 ;
        RECT 49.950 15.600 51.000 20.850 ;
        RECT 52.950 19.050 55.050 21.150 ;
        RECT 17.400 3.600 19.200 9.600 ;
        RECT 24.000 3.600 25.800 15.600 ;
        RECT 37.500 3.600 39.300 15.600 ;
        RECT 49.200 3.600 51.000 15.600 ;
        RECT 56.400 9.600 57.450 26.700 ;
        RECT 58.950 20.850 61.050 22.950 ;
        RECT 65.100 21.150 66.900 22.950 ;
        RECT 59.100 19.050 60.900 20.850 ;
        RECT 64.950 19.050 67.050 21.150 ;
        RECT 68.400 19.950 69.600 27.300 ;
        RECT 77.250 24.150 79.050 25.950 ;
        RECT 71.100 21.150 72.900 22.950 ;
        RECT 67.950 17.850 70.050 19.950 ;
        RECT 70.950 19.050 73.050 21.150 ;
        RECT 73.950 20.850 76.050 22.950 ;
        RECT 76.950 22.050 79.050 24.150 ;
        RECT 79.950 22.950 81.000 29.400 ;
        RECT 98.100 27.000 99.900 35.400 ;
        RECT 114.000 31.050 115.800 35.400 ;
        RECT 110.400 29.400 115.800 31.050 ;
        RECT 82.950 24.150 84.750 25.950 ;
        RECT 98.100 25.350 102.300 27.000 ;
        RECT 79.950 20.850 82.050 22.950 ;
        RECT 82.950 22.050 85.050 24.150 ;
        RECT 85.950 20.850 88.050 22.950 ;
        RECT 101.400 21.150 102.300 25.350 ;
        RECT 110.400 22.950 111.300 29.400 ;
        RECT 128.100 27.000 129.900 35.400 ;
        RECT 139.800 29.400 141.600 35.400 ;
        RECT 140.400 27.300 141.600 29.400 ;
        RECT 142.800 30.300 144.600 35.400 ;
        RECT 148.800 30.300 150.600 35.400 ;
        RECT 142.800 28.950 150.600 30.300 ;
        RECT 152.400 30.300 154.200 35.400 ;
        RECT 158.400 30.300 160.200 35.400 ;
        RECT 152.400 28.950 160.200 30.300 ;
        RECT 161.400 29.400 163.200 35.400 ;
        RECT 170.400 30.300 172.200 35.400 ;
        RECT 176.400 30.300 178.200 35.400 ;
        RECT 161.400 27.300 162.600 29.400 ;
        RECT 170.400 28.950 178.200 30.300 ;
        RECT 179.400 29.400 181.200 35.400 ;
        RECT 179.400 27.300 180.600 29.400 ;
        RECT 113.100 24.150 114.900 25.950 ;
        RECT 74.250 19.050 76.050 20.850 ;
        RECT 68.400 9.600 69.600 17.850 ;
        RECT 81.150 17.400 82.050 20.850 ;
        RECT 86.100 19.050 87.900 20.850 ;
        RECT 91.950 17.850 94.050 19.950 ;
        RECT 97.950 17.850 100.050 19.950 ;
        RECT 100.950 19.050 103.050 21.150 ;
        RECT 109.950 20.850 112.050 22.950 ;
        RECT 112.950 22.050 115.050 24.150 ;
        RECT 115.950 23.850 118.050 25.950 ;
        RECT 119.100 24.150 120.900 25.950 ;
        RECT 128.100 25.350 132.300 27.000 ;
        RECT 140.400 26.250 144.150 27.300 ;
        RECT 116.100 22.050 117.900 23.850 ;
        RECT 118.950 22.050 121.050 24.150 ;
        RECT 131.400 21.150 132.300 25.350 ;
        RECT 142.950 22.950 144.150 26.250 ;
        RECT 158.850 26.250 162.600 27.300 ;
        RECT 176.850 26.250 180.600 27.300 ;
        RECT 191.100 27.000 192.900 35.400 ;
        RECT 206.100 27.000 207.900 35.400 ;
        RECT 220.800 29.400 222.600 35.400 ;
        RECT 221.400 27.300 222.600 29.400 ;
        RECT 223.800 30.300 225.600 35.400 ;
        RECT 229.800 30.300 231.600 35.400 ;
        RECT 240.000 31.050 241.800 35.400 ;
        RECT 223.800 28.950 231.600 30.300 ;
        RECT 236.400 29.400 241.800 31.050 ;
        RECT 146.100 24.150 147.900 25.950 ;
        RECT 155.100 24.150 156.900 25.950 ;
        RECT 81.150 16.500 85.200 17.400 ;
        RECT 55.800 3.600 57.600 9.600 ;
        RECT 67.800 3.600 69.600 9.600 ;
        RECT 74.400 14.400 82.200 15.300 ;
        RECT 74.400 3.600 76.200 14.400 ;
        RECT 80.400 4.500 82.200 14.400 ;
        RECT 83.400 5.400 85.200 16.500 ;
        RECT 92.100 16.050 93.900 17.850 ;
        RECT 86.400 4.500 88.200 15.600 ;
        RECT 94.950 14.850 97.050 16.950 ;
        RECT 98.250 16.050 100.050 17.850 ;
        RECT 95.100 13.050 96.900 14.850 ;
        RECT 101.400 10.800 102.300 19.050 ;
        RECT 110.400 15.600 111.300 20.850 ;
        RECT 121.950 17.850 124.050 19.950 ;
        RECT 127.950 17.850 130.050 19.950 ;
        RECT 130.950 19.050 133.050 21.150 ;
        RECT 142.950 20.850 145.050 22.950 ;
        RECT 145.950 22.050 148.050 24.150 ;
        RECT 148.950 20.850 151.050 22.950 ;
        RECT 151.950 20.850 154.050 22.950 ;
        RECT 154.950 22.050 157.050 24.150 ;
        RECT 158.850 22.950 160.050 26.250 ;
        RECT 173.100 24.150 174.900 25.950 ;
        RECT 157.950 20.850 160.050 22.950 ;
        RECT 169.950 20.850 172.050 22.950 ;
        RECT 172.950 22.050 175.050 24.150 ;
        RECT 176.850 22.950 178.050 26.250 ;
        RECT 191.100 25.350 195.300 27.000 ;
        RECT 206.100 25.350 210.300 27.000 ;
        RECT 221.400 26.250 225.150 27.300 ;
        RECT 175.950 20.850 178.050 22.950 ;
        RECT 194.400 21.150 195.300 25.350 ;
        RECT 209.400 21.150 210.300 25.350 ;
        RECT 223.950 22.950 225.150 26.250 ;
        RECT 227.100 24.150 228.900 25.950 ;
        RECT 122.100 16.050 123.900 17.850 ;
        RECT 95.700 9.900 102.300 10.800 ;
        RECT 95.700 9.600 97.200 9.900 ;
        RECT 80.400 3.600 88.200 4.500 ;
        RECT 95.400 3.600 97.200 9.600 ;
        RECT 101.400 9.600 102.300 9.900 ;
        RECT 101.400 3.600 103.200 9.600 ;
        RECT 109.800 3.600 111.600 15.600 ;
        RECT 112.800 14.700 120.600 15.600 ;
        RECT 124.950 14.850 127.050 16.950 ;
        RECT 128.250 16.050 130.050 17.850 ;
        RECT 112.800 3.600 114.600 14.700 ;
        RECT 118.800 3.600 120.600 14.700 ;
        RECT 125.100 13.050 126.900 14.850 ;
        RECT 131.400 10.800 132.300 19.050 ;
        RECT 139.950 17.850 142.050 19.950 ;
        RECT 140.250 16.050 142.050 17.850 ;
        RECT 143.850 15.600 145.050 20.850 ;
        RECT 149.100 19.050 150.900 20.850 ;
        RECT 152.100 19.050 153.900 20.850 ;
        RECT 157.950 15.600 159.150 20.850 ;
        RECT 160.950 17.850 163.050 19.950 ;
        RECT 170.100 19.050 171.900 20.850 ;
        RECT 160.950 16.050 162.750 17.850 ;
        RECT 175.950 15.600 177.150 20.850 ;
        RECT 178.950 17.850 181.050 19.950 ;
        RECT 184.950 17.850 187.050 19.950 ;
        RECT 190.950 17.850 193.050 19.950 ;
        RECT 193.950 19.050 196.050 21.150 ;
        RECT 178.950 16.050 180.750 17.850 ;
        RECT 185.100 16.050 186.900 17.850 ;
        RECT 125.700 9.900 132.300 10.800 ;
        RECT 125.700 9.600 127.200 9.900 ;
        RECT 125.400 3.600 127.200 9.600 ;
        RECT 131.400 9.600 132.300 9.900 ;
        RECT 131.400 3.600 133.200 9.600 ;
        RECT 143.700 3.600 145.500 15.600 ;
        RECT 157.500 3.600 159.300 15.600 ;
        RECT 175.500 3.600 177.300 15.600 ;
        RECT 187.950 14.850 190.050 16.950 ;
        RECT 191.250 16.050 193.050 17.850 ;
        RECT 188.100 13.050 189.900 14.850 ;
        RECT 194.400 10.800 195.300 19.050 ;
        RECT 199.950 17.850 202.050 19.950 ;
        RECT 205.950 17.850 208.050 19.950 ;
        RECT 208.950 19.050 211.050 21.150 ;
        RECT 223.950 20.850 226.050 22.950 ;
        RECT 226.950 22.050 229.050 24.150 ;
        RECT 236.400 22.950 237.300 29.400 ;
        RECT 254.100 27.000 255.900 35.400 ;
        RECT 268.200 31.050 270.000 35.400 ;
        RECT 268.200 29.400 273.600 31.050 ;
        RECT 239.100 24.150 240.900 25.950 ;
        RECT 229.950 20.850 232.050 22.950 ;
        RECT 235.950 20.850 238.050 22.950 ;
        RECT 238.950 22.050 241.050 24.150 ;
        RECT 241.950 23.850 244.050 25.950 ;
        RECT 245.100 24.150 246.900 25.950 ;
        RECT 254.100 25.350 258.300 27.000 ;
        RECT 242.100 22.050 243.900 23.850 ;
        RECT 244.950 22.050 247.050 24.150 ;
        RECT 257.400 21.150 258.300 25.350 ;
        RECT 263.100 24.150 264.900 25.950 ;
        RECT 262.950 22.050 265.050 24.150 ;
        RECT 265.950 23.850 268.050 25.950 ;
        RECT 269.100 24.150 270.900 25.950 ;
        RECT 266.100 22.050 267.900 23.850 ;
        RECT 268.950 22.050 271.050 24.150 ;
        RECT 272.700 22.950 273.600 29.400 ;
        RECT 278.400 30.300 280.200 35.400 ;
        RECT 284.400 30.300 286.200 35.400 ;
        RECT 278.400 28.950 286.200 30.300 ;
        RECT 287.400 29.400 289.200 35.400 ;
        RECT 287.400 27.300 288.600 29.400 ;
        RECT 284.850 26.250 288.600 27.300 ;
        RECT 299.100 27.000 300.900 35.400 ;
        RECT 318.000 31.050 319.800 35.400 ;
        RECT 314.400 29.400 319.800 31.050 ;
        RECT 281.100 24.150 282.900 25.950 ;
        RECT 200.100 16.050 201.900 17.850 ;
        RECT 202.950 14.850 205.050 16.950 ;
        RECT 206.250 16.050 208.050 17.850 ;
        RECT 203.100 13.050 204.900 14.850 ;
        RECT 209.400 10.800 210.300 19.050 ;
        RECT 220.950 17.850 223.050 19.950 ;
        RECT 221.250 16.050 223.050 17.850 ;
        RECT 224.850 15.600 226.050 20.850 ;
        RECT 230.100 19.050 231.900 20.850 ;
        RECT 236.400 15.600 237.300 20.850 ;
        RECT 247.950 17.850 250.050 19.950 ;
        RECT 253.950 17.850 256.050 19.950 ;
        RECT 256.950 19.050 259.050 21.150 ;
        RECT 271.950 20.850 274.050 22.950 ;
        RECT 277.950 20.850 280.050 22.950 ;
        RECT 280.950 22.050 283.050 24.150 ;
        RECT 284.850 22.950 286.050 26.250 ;
        RECT 299.100 25.350 303.300 27.000 ;
        RECT 283.950 20.850 286.050 22.950 ;
        RECT 302.400 21.150 303.300 25.350 ;
        RECT 314.400 22.950 315.300 29.400 ;
        RECT 335.100 27.000 336.900 35.400 ;
        RECT 346.800 29.400 348.600 35.400 ;
        RECT 347.400 27.300 348.600 29.400 ;
        RECT 349.800 30.300 351.600 35.400 ;
        RECT 355.800 30.300 357.600 35.400 ;
        RECT 349.800 28.950 357.600 30.300 ;
        RECT 359.400 30.300 361.200 35.400 ;
        RECT 365.400 30.300 367.200 35.400 ;
        RECT 359.400 28.950 367.200 30.300 ;
        RECT 368.400 29.400 370.200 35.400 ;
        RECT 380.400 32.400 382.200 35.400 ;
        RECT 386.400 32.400 388.200 35.400 ;
        RECT 381.150 31.500 382.200 32.400 ;
        RECT 387.150 31.500 388.200 32.400 ;
        RECT 381.150 30.600 391.950 31.500 ;
        RECT 368.400 27.300 369.600 29.400 ;
        RECT 317.100 24.150 318.900 25.950 ;
        RECT 248.100 16.050 249.900 17.850 ;
        RECT 188.700 9.900 195.300 10.800 ;
        RECT 188.700 9.600 190.200 9.900 ;
        RECT 188.400 3.600 190.200 9.600 ;
        RECT 194.400 9.600 195.300 9.900 ;
        RECT 203.700 9.900 210.300 10.800 ;
        RECT 203.700 9.600 205.200 9.900 ;
        RECT 194.400 3.600 196.200 9.600 ;
        RECT 203.400 3.600 205.200 9.600 ;
        RECT 209.400 9.600 210.300 9.900 ;
        RECT 209.400 3.600 211.200 9.600 ;
        RECT 224.700 3.600 226.500 15.600 ;
        RECT 235.800 3.600 237.600 15.600 ;
        RECT 238.800 14.700 246.600 15.600 ;
        RECT 250.950 14.850 253.050 16.950 ;
        RECT 254.250 16.050 256.050 17.850 ;
        RECT 238.800 3.600 240.600 14.700 ;
        RECT 244.800 3.600 246.600 14.700 ;
        RECT 251.100 13.050 252.900 14.850 ;
        RECT 257.400 10.800 258.300 19.050 ;
        RECT 259.950 18.450 262.050 19.050 ;
        RECT 265.950 18.450 268.050 19.050 ;
        RECT 259.950 17.550 268.050 18.450 ;
        RECT 259.950 16.950 262.050 17.550 ;
        RECT 265.950 16.950 268.050 17.550 ;
        RECT 272.700 15.600 273.600 20.850 ;
        RECT 278.100 19.050 279.900 20.850 ;
        RECT 283.950 15.600 285.150 20.850 ;
        RECT 286.950 17.850 289.050 19.950 ;
        RECT 292.950 17.850 295.050 19.950 ;
        RECT 298.950 17.850 301.050 19.950 ;
        RECT 301.950 19.050 304.050 21.150 ;
        RECT 313.950 20.850 316.050 22.950 ;
        RECT 316.950 22.050 319.050 24.150 ;
        RECT 319.950 23.850 322.050 25.950 ;
        RECT 323.100 24.150 324.900 25.950 ;
        RECT 335.100 25.350 339.300 27.000 ;
        RECT 347.400 26.250 351.150 27.300 ;
        RECT 320.100 22.050 321.900 23.850 ;
        RECT 322.950 22.050 325.050 24.150 ;
        RECT 338.400 21.150 339.300 25.350 ;
        RECT 349.950 22.950 351.150 26.250 ;
        RECT 365.850 26.250 369.600 27.300 ;
        RECT 353.100 24.150 354.900 25.950 ;
        RECT 362.100 24.150 363.900 25.950 ;
        RECT 286.950 16.050 288.750 17.850 ;
        RECT 293.100 16.050 294.900 17.850 ;
        RECT 251.700 9.900 258.300 10.800 ;
        RECT 251.700 9.600 253.200 9.900 ;
        RECT 251.400 3.600 253.200 9.600 ;
        RECT 257.400 9.600 258.300 9.900 ;
        RECT 263.400 14.700 271.200 15.600 ;
        RECT 257.400 3.600 259.200 9.600 ;
        RECT 263.400 3.600 265.200 14.700 ;
        RECT 269.400 3.600 271.200 14.700 ;
        RECT 272.400 3.600 274.200 15.600 ;
        RECT 283.500 3.600 285.300 15.600 ;
        RECT 295.950 14.850 298.050 16.950 ;
        RECT 299.250 16.050 301.050 17.850 ;
        RECT 296.100 13.050 297.900 14.850 ;
        RECT 302.400 10.800 303.300 19.050 ;
        RECT 314.400 15.600 315.300 20.850 ;
        RECT 328.950 17.850 331.050 19.950 ;
        RECT 334.950 17.850 337.050 19.950 ;
        RECT 337.950 19.050 340.050 21.150 ;
        RECT 349.950 20.850 352.050 22.950 ;
        RECT 352.950 22.050 355.050 24.150 ;
        RECT 355.950 20.850 358.050 22.950 ;
        RECT 358.950 20.850 361.050 22.950 ;
        RECT 361.950 22.050 364.050 24.150 ;
        RECT 365.850 22.950 367.050 26.250 ;
        RECT 383.100 24.300 384.900 26.100 ;
        RECT 390.750 24.300 391.950 30.600 ;
        RECT 404.400 30.300 406.200 35.400 ;
        RECT 410.400 30.300 412.200 35.400 ;
        RECT 404.400 28.950 412.200 30.300 ;
        RECT 413.400 29.400 415.200 35.400 ;
        RECT 429.000 31.050 430.800 35.400 ;
        RECT 425.400 29.400 430.800 31.050 ;
        RECT 441.300 30.900 443.100 35.400 ;
        RECT 439.950 29.400 443.100 30.900 ;
        RECT 413.400 27.300 414.600 29.400 ;
        RECT 410.850 26.250 414.600 27.300 ;
        RECT 364.950 20.850 367.050 22.950 ;
        RECT 376.950 21.000 379.050 23.100 ;
        RECT 382.950 22.200 385.050 24.300 ;
        RECT 385.950 21.000 388.050 23.100 ;
        RECT 390.750 22.200 394.050 24.300 ;
        RECT 407.100 24.150 408.900 25.950 ;
        RECT 329.100 16.050 330.900 17.850 ;
        RECT 296.700 9.900 303.300 10.800 ;
        RECT 296.700 9.600 298.200 9.900 ;
        RECT 296.400 3.600 298.200 9.600 ;
        RECT 302.400 9.600 303.300 9.900 ;
        RECT 302.400 3.600 304.200 9.600 ;
        RECT 313.800 3.600 315.600 15.600 ;
        RECT 316.800 14.700 324.600 15.600 ;
        RECT 331.950 14.850 334.050 16.950 ;
        RECT 335.250 16.050 337.050 17.850 ;
        RECT 316.800 3.600 318.600 14.700 ;
        RECT 322.800 3.600 324.600 14.700 ;
        RECT 332.100 13.050 333.900 14.850 ;
        RECT 338.400 10.800 339.300 19.050 ;
        RECT 346.950 17.850 349.050 19.950 ;
        RECT 347.250 16.050 349.050 17.850 ;
        RECT 350.850 15.600 352.050 20.850 ;
        RECT 356.100 19.050 357.900 20.850 ;
        RECT 359.100 19.050 360.900 20.850 ;
        RECT 364.950 15.600 366.150 20.850 ;
        RECT 367.950 17.850 370.050 19.950 ;
        RECT 377.100 19.200 378.900 21.000 ;
        RECT 386.100 19.200 387.900 21.000 ;
        RECT 367.950 16.050 369.750 17.850 ;
        RECT 390.750 16.800 391.950 22.200 ;
        RECT 403.950 20.850 406.050 22.950 ;
        RECT 406.950 22.050 409.050 24.150 ;
        RECT 410.850 22.950 412.050 26.250 ;
        RECT 425.400 22.950 426.300 29.400 ;
        RECT 428.100 24.150 429.900 25.950 ;
        RECT 409.950 20.850 412.050 22.950 ;
        RECT 424.950 20.850 427.050 22.950 ;
        RECT 427.950 22.050 430.050 24.150 ;
        RECT 430.950 23.850 433.050 25.950 ;
        RECT 434.100 24.150 435.900 25.950 ;
        RECT 431.100 22.050 432.900 23.850 ;
        RECT 433.950 22.050 436.050 24.150 ;
        RECT 439.950 22.950 441.000 29.400 ;
        RECT 443.100 27.900 444.900 28.500 ;
        RECT 448.800 27.900 450.600 35.400 ;
        RECT 443.100 26.700 450.600 27.900 ;
        RECT 465.000 29.400 466.800 35.400 ;
        RECT 439.950 20.850 442.050 22.950 ;
        RECT 443.100 21.150 444.900 22.950 ;
        RECT 404.100 19.050 405.900 20.850 ;
        RECT 390.750 15.600 394.200 16.800 ;
        RECT 409.950 15.600 411.150 20.850 ;
        RECT 412.950 17.850 415.050 19.950 ;
        RECT 412.950 16.050 414.750 17.850 ;
        RECT 425.400 15.600 426.300 20.850 ;
        RECT 439.950 15.600 441.000 20.850 ;
        RECT 442.950 19.050 445.050 21.150 ;
        RECT 332.700 9.900 339.300 10.800 ;
        RECT 332.700 9.600 334.200 9.900 ;
        RECT 332.400 3.600 334.200 9.600 ;
        RECT 338.400 9.600 339.300 9.900 ;
        RECT 338.400 3.600 340.200 9.600 ;
        RECT 350.700 3.600 352.500 15.600 ;
        RECT 364.500 3.600 366.300 15.600 ;
        RECT 374.400 13.500 382.200 14.400 ;
        RECT 374.400 3.600 376.200 13.500 ;
        RECT 380.400 4.500 382.200 13.500 ;
        RECT 383.400 13.200 391.800 14.100 ;
        RECT 383.400 5.400 385.200 13.200 ;
        RECT 386.400 4.500 388.200 12.300 ;
        RECT 380.400 3.600 388.200 4.500 ;
        RECT 390.000 4.500 391.800 13.200 ;
        RECT 393.000 13.200 394.200 15.600 ;
        RECT 393.000 5.400 394.800 13.200 ;
        RECT 396.000 4.500 397.800 13.800 ;
        RECT 390.000 3.600 397.800 4.500 ;
        RECT 409.500 3.600 411.300 15.600 ;
        RECT 424.800 3.600 426.600 15.600 ;
        RECT 427.800 14.700 435.600 15.600 ;
        RECT 427.800 3.600 429.600 14.700 ;
        RECT 433.800 3.600 435.600 14.700 ;
        RECT 439.200 3.600 441.000 15.600 ;
        RECT 446.400 9.600 447.450 26.700 ;
        RECT 461.250 24.150 463.050 25.950 ;
        RECT 448.950 20.850 451.050 22.950 ;
        RECT 457.950 20.850 460.050 22.950 ;
        RECT 460.950 22.050 463.050 24.150 ;
        RECT 465.000 22.950 466.050 29.400 ;
        RECT 478.200 28.200 480.000 35.400 ;
        RECT 487.800 29.400 489.600 35.400 ;
        RECT 476.400 27.300 480.000 28.200 ;
        RECT 488.400 27.300 489.600 29.400 ;
        RECT 490.800 30.300 492.600 35.400 ;
        RECT 496.800 30.300 498.600 35.400 ;
        RECT 504.300 30.900 506.100 35.400 ;
        RECT 490.800 28.950 498.600 30.300 ;
        RECT 502.950 29.400 506.100 30.900 ;
        RECT 463.950 20.850 466.050 22.950 ;
        RECT 466.950 24.150 468.750 25.950 ;
        RECT 466.950 22.050 469.050 24.150 ;
        RECT 469.950 20.850 472.050 22.950 ;
        RECT 473.100 21.150 474.900 22.950 ;
        RECT 449.100 19.050 450.900 20.850 ;
        RECT 458.100 19.050 459.900 20.850 ;
        RECT 463.950 17.400 464.850 20.850 ;
        RECT 469.950 19.050 471.750 20.850 ;
        RECT 472.950 19.050 475.050 21.150 ;
        RECT 476.400 19.950 477.600 27.300 ;
        RECT 488.400 26.250 492.150 27.300 ;
        RECT 490.950 22.950 492.150 26.250 ;
        RECT 494.100 24.150 495.900 25.950 ;
        RECT 479.100 21.150 480.900 22.950 ;
        RECT 475.950 17.850 478.050 19.950 ;
        RECT 478.950 19.050 481.050 21.150 ;
        RECT 490.950 20.850 493.050 22.950 ;
        RECT 493.950 22.050 496.050 24.150 ;
        RECT 502.950 22.950 504.000 29.400 ;
        RECT 506.100 27.900 507.900 28.500 ;
        RECT 511.800 27.900 513.600 35.400 ;
        RECT 523.800 32.400 525.600 35.400 ;
        RECT 506.100 26.700 513.600 27.900 ;
        RECT 496.950 20.850 499.050 22.950 ;
        RECT 502.950 20.850 505.050 22.950 ;
        RECT 506.100 21.150 507.900 22.950 ;
        RECT 487.950 17.850 490.050 19.950 ;
        RECT 460.800 16.500 464.850 17.400 ;
        RECT 445.800 3.600 447.600 9.600 ;
        RECT 457.800 4.500 459.600 15.600 ;
        RECT 460.800 5.400 462.600 16.500 ;
        RECT 463.800 14.400 471.600 15.300 ;
        RECT 463.800 4.500 465.600 14.400 ;
        RECT 457.800 3.600 465.600 4.500 ;
        RECT 469.800 3.600 471.600 14.400 ;
        RECT 476.400 9.600 477.600 17.850 ;
        RECT 488.250 16.050 490.050 17.850 ;
        RECT 491.850 15.600 493.050 20.850 ;
        RECT 497.100 19.050 498.900 20.850 ;
        RECT 502.950 15.600 504.000 20.850 ;
        RECT 505.950 19.050 508.050 21.150 ;
        RECT 476.400 3.600 478.200 9.600 ;
        RECT 491.700 3.600 493.500 15.600 ;
        RECT 502.200 3.600 504.000 15.600 ;
        RECT 509.400 9.600 510.450 26.700 ;
        RECT 523.950 25.950 525.000 32.400 ;
        RECT 530.400 30.300 532.200 35.400 ;
        RECT 536.400 30.300 538.200 35.400 ;
        RECT 530.400 28.950 538.200 30.300 ;
        RECT 539.400 29.400 541.200 35.400 ;
        RECT 551.400 32.400 553.200 35.400 ;
        RECT 539.400 27.300 540.600 29.400 ;
        RECT 536.850 26.250 540.600 27.300 ;
        RECT 523.950 23.850 526.050 25.950 ;
        RECT 533.100 24.150 534.900 25.950 ;
        RECT 511.950 20.850 514.050 22.950 ;
        RECT 520.950 20.850 523.050 22.950 ;
        RECT 512.100 19.050 513.900 20.850 ;
        RECT 521.100 19.050 522.900 20.850 ;
        RECT 523.950 16.650 525.000 23.850 ;
        RECT 526.950 20.850 529.050 22.950 ;
        RECT 529.950 20.850 532.050 22.950 ;
        RECT 532.950 22.050 535.050 24.150 ;
        RECT 536.850 22.950 538.050 26.250 ;
        RECT 547.950 23.850 550.050 25.950 ;
        RECT 551.400 24.150 552.600 32.400 ;
        RECT 563.100 27.000 564.900 35.400 ;
        RECT 574.800 29.400 576.600 35.400 ;
        RECT 580.800 32.400 582.600 35.400 ;
        RECT 563.100 25.350 567.300 27.000 ;
        RECT 535.950 20.850 538.050 22.950 ;
        RECT 548.100 22.050 549.900 23.850 ;
        RECT 550.950 22.050 553.050 24.150 ;
        RECT 527.100 19.050 528.900 20.850 ;
        RECT 530.100 19.050 531.900 20.850 ;
        RECT 522.600 15.600 525.000 16.650 ;
        RECT 535.950 15.600 537.150 20.850 ;
        RECT 538.950 17.850 541.050 19.950 ;
        RECT 538.950 16.050 540.750 17.850 ;
        RECT 508.800 3.600 510.600 9.600 ;
        RECT 522.600 3.600 524.400 15.600 ;
        RECT 535.500 3.600 537.300 15.600 ;
        RECT 551.400 9.600 552.600 22.050 ;
        RECT 566.400 21.150 567.300 25.350 ;
        RECT 574.950 24.150 576.000 29.400 ;
        RECT 580.800 28.200 581.700 32.400 ;
        RECT 578.250 27.300 581.700 28.200 ;
        RECT 591.000 28.200 592.800 35.400 ;
        RECT 603.000 28.200 604.800 35.400 ;
        RECT 591.000 27.300 594.600 28.200 ;
        RECT 603.000 27.300 606.600 28.200 ;
        RECT 578.250 26.400 580.050 27.300 ;
        RECT 574.950 22.050 577.050 24.150 ;
        RECT 556.950 17.850 559.050 19.950 ;
        RECT 562.950 17.850 565.050 19.950 ;
        RECT 565.950 19.050 568.050 21.150 ;
        RECT 557.100 16.050 558.900 17.850 ;
        RECT 559.950 14.850 562.050 16.950 ;
        RECT 563.250 16.050 565.050 17.850 ;
        RECT 560.100 13.050 561.900 14.850 ;
        RECT 566.400 10.800 567.300 19.050 ;
        RECT 575.700 15.450 577.050 22.050 ;
        RECT 578.400 18.150 579.300 26.400 ;
        RECT 583.950 23.850 586.050 25.950 ;
        RECT 580.950 20.850 583.050 22.950 ;
        RECT 584.100 22.050 585.900 23.850 ;
        RECT 590.100 21.150 591.900 22.950 ;
        RECT 581.100 19.050 582.900 20.850 ;
        RECT 589.950 19.050 592.050 21.150 ;
        RECT 593.400 19.950 594.600 27.300 ;
        RECT 596.100 21.150 597.900 22.950 ;
        RECT 602.100 21.150 603.900 22.950 ;
        RECT 578.400 18.000 580.200 18.150 ;
        RECT 578.400 16.800 585.600 18.000 ;
        RECT 592.950 17.850 595.050 19.950 ;
        RECT 595.950 19.050 598.050 21.150 ;
        RECT 601.950 19.050 604.050 21.150 ;
        RECT 605.400 19.950 606.600 27.300 ;
        RECT 617.100 27.000 618.900 35.400 ;
        RECT 614.700 25.350 618.900 27.000 ;
        RECT 632.100 27.000 633.900 35.400 ;
        RECT 646.200 28.200 648.000 35.400 ;
        RECT 644.400 27.300 648.000 28.200 ;
        RECT 632.100 25.350 636.300 27.000 ;
        RECT 608.100 21.150 609.900 22.950 ;
        RECT 614.700 21.150 615.600 25.350 ;
        RECT 635.400 21.150 636.300 25.350 ;
        RECT 641.100 21.150 642.900 22.950 ;
        RECT 604.950 17.850 607.050 19.950 ;
        RECT 607.950 19.050 610.050 21.150 ;
        RECT 613.950 19.050 616.050 21.150 ;
        RECT 578.400 16.350 580.200 16.800 ;
        RECT 584.400 15.600 585.600 16.800 ;
        RECT 575.700 14.100 578.100 15.450 ;
        RECT 560.700 9.900 567.300 10.800 ;
        RECT 560.700 9.600 562.200 9.900 ;
        RECT 551.400 3.600 553.200 9.600 ;
        RECT 560.400 3.600 562.200 9.600 ;
        RECT 566.400 9.600 567.300 9.900 ;
        RECT 566.400 3.600 568.200 9.600 ;
        RECT 576.300 3.600 578.100 14.100 ;
        RECT 583.800 3.600 585.600 15.600 ;
        RECT 593.400 9.600 594.600 17.850 ;
        RECT 605.400 9.600 606.600 17.850 ;
        RECT 614.700 10.800 615.600 19.050 ;
        RECT 616.950 17.850 619.050 19.950 ;
        RECT 622.950 17.850 625.050 19.950 ;
        RECT 625.950 17.850 628.050 19.950 ;
        RECT 631.950 17.850 634.050 19.950 ;
        RECT 634.950 19.050 637.050 21.150 ;
        RECT 640.950 19.050 643.050 21.150 ;
        RECT 644.400 19.950 645.600 27.300 ;
        RECT 659.100 27.000 660.900 35.400 ;
        RECT 656.700 25.350 660.900 27.000 ;
        RECT 674.400 32.400 676.200 35.400 ;
        RECT 647.100 21.150 648.900 22.950 ;
        RECT 656.700 21.150 657.600 25.350 ;
        RECT 670.950 23.850 673.050 25.950 ;
        RECT 674.400 24.150 675.600 32.400 ;
        RECT 689.100 27.000 690.900 35.400 ;
        RECT 703.200 28.200 705.000 35.400 ;
        RECT 710.400 30.300 712.200 35.400 ;
        RECT 716.400 30.300 718.200 35.400 ;
        RECT 710.400 28.950 718.200 30.300 ;
        RECT 719.400 29.400 721.200 35.400 ;
        RECT 727.800 29.400 729.600 35.400 ;
        RECT 701.400 27.300 705.000 28.200 ;
        RECT 719.400 27.300 720.600 29.400 ;
        RECT 689.100 25.350 693.300 27.000 ;
        RECT 671.100 22.050 672.900 23.850 ;
        RECT 673.950 22.050 676.050 24.150 ;
        RECT 616.950 16.050 618.750 17.850 ;
        RECT 619.950 14.850 622.050 16.950 ;
        RECT 623.100 16.050 624.900 17.850 ;
        RECT 626.100 16.050 627.900 17.850 ;
        RECT 628.950 14.850 631.050 16.950 ;
        RECT 632.250 16.050 634.050 17.850 ;
        RECT 620.100 13.050 621.900 14.850 ;
        RECT 629.100 13.050 630.900 14.850 ;
        RECT 635.400 10.800 636.300 19.050 ;
        RECT 643.950 17.850 646.050 19.950 ;
        RECT 646.950 19.050 649.050 21.150 ;
        RECT 655.950 19.050 658.050 21.150 ;
        RECT 614.700 9.900 621.300 10.800 ;
        RECT 614.700 9.600 615.600 9.900 ;
        RECT 592.800 3.600 594.600 9.600 ;
        RECT 604.800 3.600 606.600 9.600 ;
        RECT 613.800 3.600 615.600 9.600 ;
        RECT 619.800 9.600 621.300 9.900 ;
        RECT 629.700 9.900 636.300 10.800 ;
        RECT 629.700 9.600 631.200 9.900 ;
        RECT 619.800 3.600 621.600 9.600 ;
        RECT 629.400 3.600 631.200 9.600 ;
        RECT 635.400 9.600 636.300 9.900 ;
        RECT 644.400 9.600 645.600 17.850 ;
        RECT 646.950 15.450 649.050 16.050 ;
        RECT 652.950 15.450 655.050 16.050 ;
        RECT 646.950 14.550 655.050 15.450 ;
        RECT 646.950 13.950 649.050 14.550 ;
        RECT 652.950 13.950 655.050 14.550 ;
        RECT 656.700 10.800 657.600 19.050 ;
        RECT 658.950 17.850 661.050 19.950 ;
        RECT 664.950 17.850 667.050 19.950 ;
        RECT 658.950 16.050 660.750 17.850 ;
        RECT 661.950 14.850 664.050 16.950 ;
        RECT 665.100 16.050 666.900 17.850 ;
        RECT 662.100 13.050 663.900 14.850 ;
        RECT 656.700 9.900 663.300 10.800 ;
        RECT 656.700 9.600 657.600 9.900 ;
        RECT 635.400 3.600 637.200 9.600 ;
        RECT 644.400 3.600 646.200 9.600 ;
        RECT 655.800 3.600 657.600 9.600 ;
        RECT 661.800 9.600 663.300 9.900 ;
        RECT 674.400 9.600 675.600 22.050 ;
        RECT 692.400 21.150 693.300 25.350 ;
        RECT 698.100 21.150 699.900 22.950 ;
        RECT 682.950 17.850 685.050 19.950 ;
        RECT 688.950 17.850 691.050 19.950 ;
        RECT 691.950 19.050 694.050 21.150 ;
        RECT 697.950 19.050 700.050 21.150 ;
        RECT 701.400 19.950 702.600 27.300 ;
        RECT 716.850 26.250 720.600 27.300 ;
        RECT 728.400 27.300 729.600 29.400 ;
        RECT 730.800 30.300 732.600 35.400 ;
        RECT 736.800 30.300 738.600 35.400 ;
        RECT 730.800 28.950 738.600 30.300 ;
        RECT 740.400 30.300 742.200 35.400 ;
        RECT 746.400 30.300 748.200 35.400 ;
        RECT 740.400 28.950 748.200 30.300 ;
        RECT 749.400 29.400 751.200 35.400 ;
        RECT 749.400 27.300 750.600 29.400 ;
        RECT 728.400 26.250 732.150 27.300 ;
        RECT 713.100 24.150 714.900 25.950 ;
        RECT 704.100 21.150 705.900 22.950 ;
        RECT 683.100 16.050 684.900 17.850 ;
        RECT 685.950 14.850 688.050 16.950 ;
        RECT 689.250 16.050 691.050 17.850 ;
        RECT 686.100 13.050 687.900 14.850 ;
        RECT 692.400 10.800 693.300 19.050 ;
        RECT 700.950 17.850 703.050 19.950 ;
        RECT 703.950 19.050 706.050 21.150 ;
        RECT 709.950 20.850 712.050 22.950 ;
        RECT 712.950 22.050 715.050 24.150 ;
        RECT 716.850 22.950 718.050 26.250 ;
        RECT 715.950 20.850 718.050 22.950 ;
        RECT 730.950 22.950 732.150 26.250 ;
        RECT 746.850 26.250 750.600 27.300 ;
        RECT 734.100 24.150 735.900 25.950 ;
        RECT 743.100 24.150 744.900 25.950 ;
        RECT 730.950 20.850 733.050 22.950 ;
        RECT 733.950 22.050 736.050 24.150 ;
        RECT 736.950 20.850 739.050 22.950 ;
        RECT 739.950 20.850 742.050 22.950 ;
        RECT 742.950 22.050 745.050 24.150 ;
        RECT 746.850 22.950 748.050 26.250 ;
        RECT 745.950 20.850 748.050 22.950 ;
        RECT 710.100 19.050 711.900 20.850 ;
        RECT 686.700 9.900 693.300 10.800 ;
        RECT 686.700 9.600 688.200 9.900 ;
        RECT 661.800 3.600 663.600 9.600 ;
        RECT 674.400 3.600 676.200 9.600 ;
        RECT 686.400 3.600 688.200 9.600 ;
        RECT 692.400 9.600 693.300 9.900 ;
        RECT 701.400 9.600 702.600 17.850 ;
        RECT 715.950 15.600 717.150 20.850 ;
        RECT 718.950 17.850 721.050 19.950 ;
        RECT 727.950 17.850 730.050 19.950 ;
        RECT 718.950 16.050 720.750 17.850 ;
        RECT 728.250 16.050 730.050 17.850 ;
        RECT 731.850 15.600 733.050 20.850 ;
        RECT 737.100 19.050 738.900 20.850 ;
        RECT 740.100 19.050 741.900 20.850 ;
        RECT 745.950 15.600 747.150 20.850 ;
        RECT 748.950 17.850 751.050 19.950 ;
        RECT 748.950 16.050 750.750 17.850 ;
        RECT 692.400 3.600 694.200 9.600 ;
        RECT 701.400 3.600 703.200 9.600 ;
        RECT 715.500 3.600 717.300 15.600 ;
        RECT 731.700 3.600 733.500 15.600 ;
        RECT 745.500 3.600 747.300 15.600 ;
      LAYER metal2 ;
        RECT 103.950 712.950 106.050 715.050 ;
        RECT 115.950 712.950 118.050 715.050 ;
        RECT 370.950 712.950 373.050 715.050 ;
        RECT 31.950 706.950 34.050 709.050 ;
        RECT 25.950 704.250 28.050 705.150 ;
        RECT 32.400 703.050 33.450 706.950 ;
        RECT 58.950 704.250 61.050 705.150 ;
        RECT 67.950 704.250 70.050 705.150 ;
        RECT 97.950 704.250 100.050 705.150 ;
        RECT 104.400 703.050 105.450 712.950 ;
        RECT 109.950 706.950 112.050 709.050 ;
        RECT 110.400 703.050 111.450 706.950 ;
        RECT 7.950 702.450 10.050 703.050 ;
        RECT 16.950 702.450 19.050 703.050 ;
        RECT 4.950 701.250 6.750 702.150 ;
        RECT 7.950 701.400 12.450 702.450 ;
        RECT 7.950 700.950 10.050 701.400 ;
        RECT 4.950 697.950 7.050 700.050 ;
        RECT 8.250 698.850 10.050 699.750 ;
        RECT 5.400 697.050 6.450 697.950 ;
        RECT 4.950 694.950 7.050 697.050 ;
        RECT 7.950 673.950 10.050 676.050 ;
        RECT 8.400 670.050 9.450 673.950 ;
        RECT 11.400 673.050 12.450 701.400 ;
        RECT 13.950 701.250 15.750 702.150 ;
        RECT 16.950 701.400 21.450 702.450 ;
        RECT 16.950 700.950 19.050 701.400 ;
        RECT 13.950 697.950 16.050 700.050 ;
        RECT 17.250 698.850 19.050 699.750 ;
        RECT 20.400 688.050 21.450 701.400 ;
        RECT 25.950 700.950 28.050 703.050 ;
        RECT 29.250 701.250 30.750 702.150 ;
        RECT 31.950 700.950 34.050 703.050 ;
        RECT 35.250 701.250 37.050 702.150 ;
        RECT 40.950 700.950 43.050 703.050 ;
        RECT 46.950 700.950 49.050 703.050 ;
        RECT 49.950 701.250 51.750 702.150 ;
        RECT 52.950 700.950 55.050 703.050 ;
        RECT 56.250 701.250 57.750 702.150 ;
        RECT 58.950 700.950 61.050 703.050 ;
        RECT 67.950 700.950 70.050 703.050 ;
        RECT 71.250 701.250 72.750 702.150 ;
        RECT 73.950 700.950 76.050 703.050 ;
        RECT 77.250 701.250 79.050 702.150 ;
        RECT 79.950 700.950 82.050 703.050 ;
        RECT 82.950 701.250 84.750 702.150 ;
        RECT 85.950 700.950 88.050 703.050 ;
        RECT 91.950 702.450 94.050 703.050 ;
        RECT 91.950 701.400 96.450 702.450 ;
        RECT 91.950 700.950 94.050 701.400 ;
        RECT 26.400 700.050 27.450 700.950 ;
        RECT 25.950 697.950 28.050 700.050 ;
        RECT 28.950 697.950 31.050 700.050 ;
        RECT 32.250 698.850 33.750 699.750 ;
        RECT 34.950 697.950 37.050 700.050 ;
        RECT 40.950 698.850 43.050 699.750 ;
        RECT 43.950 698.250 46.050 699.150 ;
        RECT 29.400 697.050 30.450 697.950 ;
        RECT 35.400 697.050 36.450 697.950 ;
        RECT 28.950 694.950 31.050 697.050 ;
        RECT 34.950 694.950 37.050 697.050 ;
        RECT 43.950 696.450 46.050 697.050 ;
        RECT 47.400 696.450 48.450 700.950 ;
        RECT 59.400 700.050 60.450 700.950 ;
        RECT 49.950 697.950 52.050 700.050 ;
        RECT 53.250 698.850 54.750 699.750 ;
        RECT 55.950 697.950 58.050 700.050 ;
        RECT 58.950 697.950 61.050 700.050 ;
        RECT 43.950 695.400 48.450 696.450 ;
        RECT 43.950 694.950 46.050 695.400 ;
        RECT 50.400 688.050 51.450 697.950 ;
        RECT 19.950 685.950 22.050 688.050 ;
        RECT 49.950 685.950 52.050 688.050 ;
        RECT 56.400 684.450 57.450 697.950 ;
        RECT 53.400 683.400 57.450 684.450 ;
        RECT 19.950 679.950 22.050 682.050 ;
        RECT 16.950 673.950 19.050 676.050 ;
        RECT 10.950 670.950 13.050 673.050 ;
        RECT 13.950 670.950 16.050 673.050 ;
        RECT 4.950 668.250 6.750 669.150 ;
        RECT 7.950 667.950 10.050 670.050 ;
        RECT 11.250 668.250 13.050 669.150 ;
        RECT 4.950 664.950 7.050 667.050 ;
        RECT 8.250 665.850 9.750 666.750 ;
        RECT 10.950 664.950 13.050 667.050 ;
        RECT 5.400 664.050 6.450 664.950 ;
        RECT 4.950 661.950 7.050 664.050 ;
        RECT 7.950 661.950 10.050 664.050 ;
        RECT 8.400 631.050 9.450 661.950 ;
        RECT 11.400 634.050 12.450 664.950 ;
        RECT 14.400 664.050 15.450 670.950 ;
        RECT 17.400 667.050 18.450 673.950 ;
        RECT 20.400 670.050 21.450 679.950 ;
        RECT 28.950 676.950 31.050 679.050 ;
        RECT 29.400 673.050 30.450 676.950 ;
        RECT 22.950 670.950 25.050 673.050 ;
        RECT 26.250 671.250 27.750 672.150 ;
        RECT 28.950 670.950 31.050 673.050 ;
        RECT 19.950 667.950 22.050 670.050 ;
        RECT 23.250 668.850 24.750 669.750 ;
        RECT 25.950 667.950 28.050 670.050 ;
        RECT 29.250 668.850 31.050 669.750 ;
        RECT 31.950 668.250 33.750 669.150 ;
        RECT 34.950 667.950 37.050 670.050 ;
        RECT 38.250 668.250 40.050 669.150 ;
        RECT 40.950 667.950 43.050 670.050 ;
        RECT 46.950 668.250 48.750 669.150 ;
        RECT 49.950 667.950 52.050 670.050 ;
        RECT 16.950 664.950 19.050 667.050 ;
        RECT 19.950 665.850 22.050 666.750 ;
        RECT 13.950 661.950 16.050 664.050 ;
        RECT 26.400 658.050 27.450 667.950 ;
        RECT 31.950 664.950 34.050 667.050 ;
        RECT 35.250 665.850 36.750 666.750 ;
        RECT 37.950 664.950 40.050 667.050 ;
        RECT 25.950 655.950 28.050 658.050 ;
        RECT 32.400 634.050 33.450 664.950 ;
        RECT 37.950 637.950 40.050 640.050 ;
        RECT 38.400 634.050 39.450 637.950 ;
        RECT 41.400 637.050 42.450 667.950 ;
        RECT 53.400 667.050 54.450 683.400 ;
        RECT 55.950 679.950 58.050 682.050 ;
        RECT 56.400 670.050 57.450 679.950 ;
        RECT 55.950 667.950 58.050 670.050 ;
        RECT 46.950 664.950 49.050 667.050 ;
        RECT 50.250 665.850 51.750 666.750 ;
        RECT 52.950 664.950 55.050 667.050 ;
        RECT 56.250 665.850 58.050 666.750 ;
        RECT 52.950 662.850 55.050 663.750 ;
        RECT 59.400 640.050 60.450 697.950 ;
        RECT 68.400 688.050 69.450 700.950 ;
        RECT 70.950 697.950 73.050 700.050 ;
        RECT 74.250 698.850 75.750 699.750 ;
        RECT 76.950 697.950 79.050 700.050 ;
        RECT 67.950 685.950 70.050 688.050 ;
        RECT 77.400 676.050 78.450 697.950 ;
        RECT 80.400 691.050 81.450 700.950 ;
        RECT 95.400 700.050 96.450 701.400 ;
        RECT 97.950 700.950 100.050 703.050 ;
        RECT 101.250 701.250 102.750 702.150 ;
        RECT 103.950 700.950 106.050 703.050 ;
        RECT 107.250 701.250 109.050 702.150 ;
        RECT 109.950 700.950 112.050 703.050 ;
        RECT 112.950 700.950 115.050 703.050 ;
        RECT 82.950 697.950 85.050 700.050 ;
        RECT 86.250 698.850 88.050 699.750 ;
        RECT 88.950 698.250 91.050 699.150 ;
        RECT 91.950 698.850 94.050 699.750 ;
        RECT 94.950 699.450 97.050 700.050 ;
        RECT 94.950 698.400 99.450 699.450 ;
        RECT 94.950 697.950 97.050 698.400 ;
        RECT 88.950 694.950 91.050 697.050 ;
        RECT 91.950 694.950 94.050 697.050 ;
        RECT 98.400 696.450 99.450 698.400 ;
        RECT 100.950 697.950 103.050 700.050 ;
        RECT 104.250 698.850 105.750 699.750 ;
        RECT 106.950 697.950 109.050 700.050 ;
        RECT 109.950 698.250 112.050 699.150 ;
        RECT 112.950 698.850 115.050 699.750 ;
        RECT 107.400 697.050 108.450 697.950 ;
        RECT 100.950 696.450 103.050 697.050 ;
        RECT 98.400 695.400 103.050 696.450 ;
        RECT 100.950 694.950 103.050 695.400 ;
        RECT 106.950 694.950 109.050 697.050 ;
        RECT 109.950 694.950 112.050 697.050 ;
        RECT 89.400 694.050 90.450 694.950 ;
        RECT 88.950 691.950 91.050 694.050 ;
        RECT 92.400 691.050 93.450 694.950 ;
        RECT 79.950 688.950 82.050 691.050 ;
        RECT 91.950 688.950 94.050 691.050 ;
        RECT 88.950 679.950 91.050 682.050 ;
        RECT 85.950 676.950 88.050 679.050 ;
        RECT 76.950 673.950 79.050 676.050 ;
        RECT 73.950 670.950 76.050 673.050 ;
        RECT 61.950 668.250 63.750 669.150 ;
        RECT 64.950 667.950 67.050 670.050 ;
        RECT 68.250 668.250 70.050 669.150 ;
        RECT 70.950 667.950 73.050 670.050 ;
        RECT 61.950 664.950 64.050 667.050 ;
        RECT 65.250 665.850 66.750 666.750 ;
        RECT 67.950 666.450 70.050 667.050 ;
        RECT 71.400 666.450 72.450 667.950 ;
        RECT 67.950 665.400 72.450 666.450 ;
        RECT 74.400 666.450 75.450 670.950 ;
        RECT 76.950 668.250 78.750 669.150 ;
        RECT 79.950 667.950 82.050 670.050 ;
        RECT 83.250 668.250 85.050 669.150 ;
        RECT 86.400 667.050 87.450 676.950 ;
        RECT 89.400 670.050 90.450 679.950 ;
        RECT 110.400 679.050 111.450 694.950 ;
        RECT 116.400 694.050 117.450 712.950 ;
        RECT 238.950 709.950 241.050 712.050 ;
        RECT 358.950 709.950 361.050 712.050 ;
        RECT 148.950 706.950 151.050 709.050 ;
        RECT 217.950 706.950 220.050 709.050 ;
        RECT 142.950 704.250 145.050 705.150 ;
        RECT 149.400 703.050 150.450 706.950 ;
        RECT 166.950 703.950 169.050 706.050 ;
        RECT 172.950 703.950 175.050 706.050 ;
        RECT 181.950 703.950 184.050 706.050 ;
        RECT 187.950 703.950 190.050 706.050 ;
        RECT 193.950 704.250 196.050 705.150 ;
        RECT 196.950 703.950 199.050 706.050 ;
        RECT 202.950 705.450 205.050 706.050 ;
        RECT 200.400 704.400 205.050 705.450 ;
        RECT 208.950 705.450 211.050 706.050 ;
        RECT 121.950 702.450 124.050 703.050 ;
        RECT 130.950 702.450 133.050 703.050 ;
        RECT 119.400 701.400 124.050 702.450 ;
        RECT 115.950 691.950 118.050 694.050 ;
        RECT 119.400 691.050 120.450 701.400 ;
        RECT 121.950 700.950 124.050 701.400 ;
        RECT 125.250 701.250 127.050 702.150 ;
        RECT 128.400 701.400 133.050 702.450 ;
        RECT 121.950 698.850 123.750 699.750 ;
        RECT 124.950 697.950 127.050 700.050 ;
        RECT 112.950 688.950 115.050 691.050 ;
        RECT 118.950 688.950 121.050 691.050 ;
        RECT 100.950 676.950 103.050 679.050 ;
        RECT 109.950 676.950 112.050 679.050 ;
        RECT 101.400 673.050 102.450 676.950 ;
        RECT 103.950 675.450 106.050 676.050 ;
        RECT 103.950 674.400 111.450 675.450 ;
        RECT 103.950 673.950 106.050 674.400 ;
        RECT 91.950 670.950 94.050 673.050 ;
        RECT 95.250 671.250 96.750 672.150 ;
        RECT 97.950 670.950 100.050 673.050 ;
        RECT 100.950 670.950 103.050 673.050 ;
        RECT 104.250 671.850 105.750 672.750 ;
        RECT 106.950 670.950 109.050 673.050 ;
        RECT 88.950 667.950 91.050 670.050 ;
        RECT 92.250 668.850 93.750 669.750 ;
        RECT 94.950 667.950 97.050 670.050 ;
        RECT 98.250 668.850 100.050 669.750 ;
        RECT 100.950 668.850 103.050 669.750 ;
        RECT 106.950 668.850 109.050 669.750 ;
        RECT 110.400 667.050 111.450 674.400 ;
        RECT 113.400 673.050 114.450 688.950 ;
        RECT 118.950 679.950 121.050 682.050 ;
        RECT 115.950 676.950 118.050 679.050 ;
        RECT 116.400 673.050 117.450 676.950 ;
        RECT 119.400 673.050 120.450 679.950 ;
        RECT 124.950 673.950 127.050 676.050 ;
        RECT 125.400 673.050 126.450 673.950 ;
        RECT 128.400 673.050 129.450 701.400 ;
        RECT 130.950 700.950 133.050 701.400 ;
        RECT 134.250 701.250 136.050 702.150 ;
        RECT 142.950 700.950 145.050 703.050 ;
        RECT 146.250 701.250 147.750 702.150 ;
        RECT 148.950 700.950 151.050 703.050 ;
        RECT 152.250 701.250 154.050 702.150 ;
        RECT 154.950 701.250 157.050 702.150 ;
        RECT 160.950 701.250 163.050 702.150 ;
        RECT 130.950 698.850 132.750 699.750 ;
        RECT 133.950 697.950 136.050 700.050 ;
        RECT 145.950 697.950 148.050 700.050 ;
        RECT 149.250 698.850 150.750 699.750 ;
        RECT 151.950 697.950 154.050 700.050 ;
        RECT 160.950 697.950 163.050 700.050 ;
        RECT 152.400 697.050 153.450 697.950 ;
        RECT 151.950 694.950 154.050 697.050 ;
        RECT 167.400 694.050 168.450 703.950 ;
        RECT 173.400 703.050 174.450 703.950 ;
        RECT 169.950 701.250 171.750 702.150 ;
        RECT 172.950 700.950 175.050 703.050 ;
        RECT 178.950 700.950 181.050 703.050 ;
        RECT 169.950 697.950 172.050 700.050 ;
        RECT 173.250 698.850 175.050 699.750 ;
        RECT 175.950 698.250 178.050 699.150 ;
        RECT 178.950 698.850 181.050 699.750 ;
        RECT 170.400 696.450 171.450 697.950 ;
        RECT 182.400 697.050 183.450 703.950 ;
        RECT 188.400 703.050 189.450 703.950 ;
        RECT 184.950 701.250 186.750 702.150 ;
        RECT 187.950 700.950 190.050 703.050 ;
        RECT 191.250 701.250 192.750 702.150 ;
        RECT 193.950 700.950 196.050 703.050 ;
        RECT 194.400 700.050 195.450 700.950 ;
        RECT 184.950 697.950 187.050 700.050 ;
        RECT 188.250 698.850 189.750 699.750 ;
        RECT 190.950 697.950 193.050 700.050 ;
        RECT 193.950 697.950 196.050 700.050 ;
        RECT 191.400 697.050 192.450 697.950 ;
        RECT 170.400 695.400 174.450 696.450 ;
        RECT 166.950 691.950 169.050 694.050 ;
        RECT 169.950 691.950 172.050 694.050 ;
        RECT 154.950 688.950 157.050 691.050 ;
        RECT 139.950 682.950 142.050 685.050 ;
        RECT 148.950 682.950 151.050 685.050 ;
        RECT 112.950 670.950 115.050 673.050 ;
        RECT 115.950 670.950 118.050 673.050 ;
        RECT 118.950 670.950 121.050 673.050 ;
        RECT 122.250 671.250 123.750 672.150 ;
        RECT 124.950 670.950 127.050 673.050 ;
        RECT 127.950 670.950 130.050 673.050 ;
        RECT 113.400 669.450 114.450 670.950 ;
        RECT 115.950 669.450 118.050 670.050 ;
        RECT 113.400 668.400 118.050 669.450 ;
        RECT 119.250 668.850 120.750 669.750 ;
        RECT 76.950 666.450 79.050 667.050 ;
        RECT 74.400 665.400 79.050 666.450 ;
        RECT 80.250 665.850 81.750 666.750 ;
        RECT 67.950 664.950 70.050 665.400 ;
        RECT 76.950 664.950 79.050 665.400 ;
        RECT 82.950 664.950 85.050 667.050 ;
        RECT 85.950 664.950 88.050 667.050 ;
        RECT 88.950 665.850 91.050 666.750 ;
        RECT 109.950 664.950 112.050 667.050 ;
        RECT 62.400 661.050 63.450 664.950 ;
        RECT 64.950 661.950 67.050 664.050 ;
        RECT 61.950 658.950 64.050 661.050 ;
        RECT 58.950 637.950 61.050 640.050 ;
        RECT 40.950 634.950 43.050 637.050 ;
        RECT 43.950 635.250 46.050 636.150 ;
        RECT 10.950 631.950 13.050 634.050 ;
        RECT 16.950 631.950 19.050 634.050 ;
        RECT 19.950 631.950 22.050 634.050 ;
        RECT 31.950 633.450 34.050 634.050 ;
        RECT 29.400 632.400 34.050 633.450 ;
        RECT 4.950 629.250 7.050 630.150 ;
        RECT 7.950 628.950 10.050 631.050 ;
        RECT 10.950 629.250 13.050 630.150 ;
        RECT 13.950 629.250 16.050 630.150 ;
        RECT 4.950 625.950 7.050 628.050 ;
        RECT 8.250 626.250 9.750 627.150 ;
        RECT 10.950 625.950 13.050 628.050 ;
        RECT 13.950 625.950 16.050 628.050 ;
        RECT 11.400 625.050 12.450 625.950 ;
        RECT 17.400 625.050 18.450 631.950 ;
        RECT 19.950 629.850 22.050 630.750 ;
        RECT 22.950 629.250 25.050 630.150 ;
        RECT 29.400 628.050 30.450 632.400 ;
        RECT 31.950 631.950 34.050 632.400 ;
        RECT 35.250 632.250 36.750 633.150 ;
        RECT 37.950 631.950 40.050 634.050 ;
        RECT 40.950 632.250 42.750 633.150 ;
        RECT 43.950 631.950 46.050 634.050 ;
        RECT 49.950 633.450 52.050 634.050 ;
        RECT 47.250 632.250 48.750 633.150 ;
        RECT 49.950 632.400 54.450 633.450 ;
        RECT 49.950 631.950 52.050 632.400 ;
        RECT 31.950 629.850 33.750 630.750 ;
        RECT 34.950 628.950 37.050 631.050 ;
        RECT 38.250 629.850 40.050 630.750 ;
        RECT 40.950 628.950 43.050 631.050 ;
        RECT 43.950 628.950 46.050 631.050 ;
        RECT 46.950 628.950 49.050 631.050 ;
        RECT 50.250 629.850 52.050 630.750 ;
        RECT 22.950 625.950 25.050 628.050 ;
        RECT 28.950 625.950 31.050 628.050 ;
        RECT 7.950 622.950 10.050 625.050 ;
        RECT 10.950 622.950 13.050 625.050 ;
        RECT 16.950 622.950 19.050 625.050 ;
        RECT 8.400 603.450 9.450 622.950 ;
        RECT 13.950 604.950 16.050 607.050 ;
        RECT 5.400 602.400 9.450 603.450 ;
        RECT 5.400 601.050 6.450 602.400 ;
        RECT 4.950 598.950 7.050 601.050 ;
        RECT 8.250 599.250 9.750 600.150 ;
        RECT 10.950 598.950 13.050 601.050 ;
        RECT 14.400 598.050 15.450 604.950 ;
        RECT 19.950 598.950 22.050 601.050 ;
        RECT 4.950 596.850 6.750 597.750 ;
        RECT 7.950 595.950 10.050 598.050 ;
        RECT 11.250 596.850 12.750 597.750 ;
        RECT 13.950 595.950 16.050 598.050 ;
        RECT 13.950 593.850 16.050 594.750 ;
        RECT 20.400 589.050 21.450 598.950 ;
        RECT 23.400 598.050 24.450 625.950 ;
        RECT 35.400 622.050 36.450 628.950 ;
        RECT 34.950 619.950 37.050 622.050 ;
        RECT 41.400 604.050 42.450 628.950 ;
        RECT 28.950 601.950 31.050 604.050 ;
        RECT 40.950 601.950 43.050 604.050 ;
        RECT 25.950 599.250 28.050 600.150 ;
        RECT 28.950 599.850 31.050 600.750 ;
        RECT 31.950 598.950 34.050 601.050 ;
        RECT 35.250 599.250 36.750 600.150 ;
        RECT 37.950 598.950 40.050 601.050 ;
        RECT 22.950 595.950 25.050 598.050 ;
        RECT 25.950 595.950 28.050 598.050 ;
        RECT 31.950 596.850 33.750 597.750 ;
        RECT 34.950 595.950 37.050 598.050 ;
        RECT 38.250 596.850 39.750 597.750 ;
        RECT 40.950 597.450 43.050 598.050 ;
        RECT 44.400 597.450 45.450 628.950 ;
        RECT 47.400 628.050 48.450 628.950 ;
        RECT 46.950 625.950 49.050 628.050 ;
        RECT 53.400 604.050 54.450 632.400 ;
        RECT 55.950 631.950 58.050 634.050 ;
        RECT 56.400 624.450 57.450 631.950 ;
        RECT 61.950 628.950 64.050 631.050 ;
        RECT 58.950 626.250 61.050 627.150 ;
        RECT 61.950 626.850 64.050 627.750 ;
        RECT 58.950 624.450 61.050 625.050 ;
        RECT 56.400 623.400 61.050 624.450 ;
        RECT 58.950 622.950 61.050 623.400 ;
        RECT 61.950 613.950 64.050 616.050 ;
        RECT 52.950 601.950 55.050 604.050 ;
        RECT 49.950 598.950 52.050 601.050 ;
        RECT 40.950 596.400 45.450 597.450 ;
        RECT 40.950 595.950 43.050 596.400 ;
        RECT 23.400 595.050 24.450 595.950 ;
        RECT 35.400 595.050 36.450 595.950 ;
        RECT 22.950 592.950 25.050 595.050 ;
        RECT 34.950 592.950 37.050 595.050 ;
        RECT 40.950 593.850 43.050 594.750 ;
        RECT 50.400 594.450 51.450 598.950 ;
        RECT 52.950 596.250 54.750 597.150 ;
        RECT 55.950 595.950 58.050 598.050 ;
        RECT 59.250 596.250 61.050 597.150 ;
        RECT 52.950 594.450 55.050 595.050 ;
        RECT 50.400 593.400 55.050 594.450 ;
        RECT 56.250 593.850 57.750 594.750 ;
        RECT 52.950 592.950 55.050 593.400 ;
        RECT 58.950 592.950 61.050 595.050 ;
        RECT 19.950 586.950 22.050 589.050 ;
        RECT 16.950 580.950 19.050 583.050 ;
        RECT 17.400 558.450 18.450 580.950 ;
        RECT 62.400 568.050 63.450 613.950 ;
        RECT 65.400 607.050 66.450 661.950 ;
        RECT 83.400 658.050 84.450 664.950 ;
        RECT 113.400 664.050 114.450 668.400 ;
        RECT 115.950 667.950 118.050 668.400 ;
        RECT 121.950 667.950 124.050 670.050 ;
        RECT 125.250 668.850 127.050 669.750 ;
        RECT 127.950 668.250 129.750 669.150 ;
        RECT 130.950 667.950 133.050 670.050 ;
        RECT 134.250 668.250 136.050 669.150 ;
        RECT 136.950 667.950 139.050 670.050 ;
        RECT 115.950 665.850 118.050 666.750 ;
        RECT 127.950 664.950 130.050 667.050 ;
        RECT 131.250 665.850 132.750 666.750 ;
        RECT 133.950 664.950 136.050 667.050 ;
        RECT 112.950 661.950 115.050 664.050 ;
        RECT 137.400 661.050 138.450 667.950 ;
        RECT 140.400 667.050 141.450 682.950 ;
        RECT 145.950 679.950 148.050 682.050 ;
        RECT 142.950 673.950 145.050 676.050 ;
        RECT 139.950 664.950 142.050 667.050 ;
        RECT 136.950 658.950 139.050 661.050 ;
        RECT 82.950 655.950 85.050 658.050 ;
        RECT 82.950 637.950 85.050 640.050 ;
        RECT 139.950 637.950 142.050 640.050 ;
        RECT 74.400 632.400 81.450 633.450 ;
        RECT 74.400 631.050 75.450 632.400 ;
        RECT 80.400 631.050 81.450 632.400 ;
        RECT 67.950 628.950 70.050 631.050 ;
        RECT 73.950 628.950 76.050 631.050 ;
        RECT 77.250 629.250 79.050 630.150 ;
        RECT 79.950 628.950 82.050 631.050 ;
        RECT 67.950 626.850 70.050 627.750 ;
        RECT 70.950 626.250 73.050 627.150 ;
        RECT 73.950 626.850 75.750 627.750 ;
        RECT 76.950 625.950 79.050 628.050 ;
        RECT 70.950 622.950 73.050 625.050 ;
        RECT 64.950 604.950 67.050 607.050 ;
        RECT 67.950 601.950 70.050 604.050 ;
        RECT 64.950 598.950 67.050 601.050 ;
        RECT 65.400 598.050 66.450 598.950 ;
        RECT 64.950 595.950 67.050 598.050 ;
        RECT 68.400 595.050 69.450 601.950 ;
        RECT 70.950 598.950 73.050 601.050 ;
        RECT 71.400 598.050 72.450 598.950 ;
        RECT 70.950 595.950 73.050 598.050 ;
        RECT 74.250 596.250 76.050 597.150 ;
        RECT 64.950 593.850 66.750 594.750 ;
        RECT 67.950 592.950 70.050 595.050 ;
        RECT 71.250 593.850 72.750 594.750 ;
        RECT 73.950 592.950 76.050 595.050 ;
        RECT 67.950 590.850 70.050 591.750 ;
        RECT 46.950 565.950 49.050 568.050 ;
        RECT 61.950 565.950 64.050 568.050 ;
        RECT 19.950 560.250 22.050 561.150 ;
        RECT 40.950 560.250 43.050 561.150 ;
        RECT 19.950 558.450 22.050 559.050 ;
        RECT 4.950 557.250 7.050 558.150 ;
        RECT 10.950 557.250 13.050 558.150 ;
        RECT 17.400 557.400 22.050 558.450 ;
        RECT 19.950 556.950 22.050 557.400 ;
        RECT 23.250 557.250 24.750 558.150 ;
        RECT 25.950 556.950 28.050 559.050 ;
        RECT 29.250 557.250 31.050 558.150 ;
        RECT 31.950 557.250 33.750 558.150 ;
        RECT 34.950 556.950 37.050 559.050 ;
        RECT 38.250 557.250 39.750 558.150 ;
        RECT 40.950 556.950 43.050 559.050 ;
        RECT 20.400 556.050 21.450 556.950 ;
        RECT 10.950 553.950 13.050 556.050 ;
        RECT 19.950 553.950 22.050 556.050 ;
        RECT 22.950 553.950 25.050 556.050 ;
        RECT 26.250 554.850 27.750 555.750 ;
        RECT 28.950 553.950 31.050 556.050 ;
        RECT 31.950 553.950 34.050 556.050 ;
        RECT 35.250 554.850 36.750 555.750 ;
        RECT 37.950 553.950 40.050 556.050 ;
        RECT 11.400 544.050 12.450 553.950 ;
        RECT 23.400 553.050 24.450 553.950 ;
        RECT 22.950 550.950 25.050 553.050 ;
        RECT 10.950 541.950 13.050 544.050 ;
        RECT 23.400 532.050 24.450 550.950 ;
        RECT 29.400 550.050 30.450 553.950 ;
        RECT 28.950 547.950 31.050 550.050 ;
        RECT 38.400 535.050 39.450 553.950 ;
        RECT 41.400 553.050 42.450 556.950 ;
        RECT 47.400 553.050 48.450 565.950 ;
        RECT 58.950 562.950 61.050 565.050 ;
        RECT 52.950 559.950 55.050 562.050 ;
        RECT 53.400 559.050 54.450 559.950 ;
        RECT 59.400 559.050 60.450 562.950 ;
        RECT 62.400 561.450 63.450 565.950 ;
        RECT 62.400 560.400 66.450 561.450 ;
        RECT 65.400 559.050 66.450 560.400 ;
        RECT 70.950 560.250 73.050 561.150 ;
        RECT 49.950 557.250 51.750 558.150 ;
        RECT 52.950 556.950 55.050 559.050 ;
        RECT 58.950 556.950 61.050 559.050 ;
        RECT 61.950 557.250 63.750 558.150 ;
        RECT 64.950 556.950 67.050 559.050 ;
        RECT 68.250 557.250 69.750 558.150 ;
        RECT 70.950 556.950 73.050 559.050 ;
        RECT 74.400 558.450 75.450 592.950 ;
        RECT 77.400 565.050 78.450 625.950 ;
        RECT 83.400 612.450 84.450 637.950 ;
        RECT 106.950 634.950 109.050 637.050 ;
        RECT 121.950 634.950 124.050 637.050 ;
        RECT 91.950 631.950 94.050 634.050 ;
        RECT 94.950 632.250 97.050 633.150 ;
        RECT 85.950 628.950 88.050 631.050 ;
        RECT 92.400 628.050 93.450 631.950 ;
        RECT 94.950 628.950 97.050 631.050 ;
        RECT 98.250 629.250 99.750 630.150 ;
        RECT 100.950 628.950 103.050 631.050 ;
        RECT 104.250 629.250 106.050 630.150 ;
        RECT 85.950 626.850 88.050 627.750 ;
        RECT 88.950 626.250 91.050 627.150 ;
        RECT 91.950 625.950 94.050 628.050 ;
        RECT 95.400 625.050 96.450 628.950 ;
        RECT 97.950 625.950 100.050 628.050 ;
        RECT 101.250 626.850 102.750 627.750 ;
        RECT 103.950 625.950 106.050 628.050 ;
        RECT 88.950 622.950 91.050 625.050 ;
        RECT 94.950 622.950 97.050 625.050 ;
        RECT 104.400 622.050 105.450 625.950 ;
        RECT 103.950 619.950 106.050 622.050 ;
        RECT 80.400 611.400 84.450 612.450 ;
        RECT 80.400 586.050 81.450 611.400 ;
        RECT 107.400 610.050 108.450 634.950 ;
        RECT 109.950 632.250 112.050 633.150 ;
        RECT 109.950 628.950 112.050 631.050 ;
        RECT 113.250 629.250 114.750 630.150 ;
        RECT 115.950 628.950 118.050 631.050 ;
        RECT 119.250 629.250 121.050 630.150 ;
        RECT 110.400 622.050 111.450 628.950 ;
        RECT 112.950 625.950 115.050 628.050 ;
        RECT 116.250 626.850 117.750 627.750 ;
        RECT 118.950 627.450 121.050 628.050 ;
        RECT 122.400 627.450 123.450 634.950 ;
        RECT 127.950 631.950 130.050 634.050 ;
        RECT 133.950 631.950 136.050 634.050 ;
        RECT 128.400 631.050 129.450 631.950 ;
        RECT 134.400 631.050 135.450 631.950 ;
        RECT 124.950 629.250 126.750 630.150 ;
        RECT 127.950 628.950 130.050 631.050 ;
        RECT 133.950 628.950 136.050 631.050 ;
        RECT 136.950 628.950 139.050 631.050 ;
        RECT 140.400 630.450 141.450 637.950 ;
        RECT 143.400 637.050 144.450 673.950 ;
        RECT 146.400 673.050 147.450 679.950 ;
        RECT 149.400 673.050 150.450 682.950 ;
        RECT 155.400 673.050 156.450 688.950 ;
        RECT 163.950 679.950 166.050 682.050 ;
        RECT 166.950 679.950 169.050 682.050 ;
        RECT 164.400 676.050 165.450 679.950 ;
        RECT 163.950 673.950 166.050 676.050 ;
        RECT 167.400 673.050 168.450 679.950 ;
        RECT 145.950 670.950 148.050 673.050 ;
        RECT 148.950 670.950 151.050 673.050 ;
        RECT 152.250 671.250 153.750 672.150 ;
        RECT 154.950 670.950 157.050 673.050 ;
        RECT 160.950 670.950 163.050 673.050 ;
        RECT 164.250 671.850 165.750 672.750 ;
        RECT 166.950 670.950 169.050 673.050 ;
        RECT 145.950 667.950 148.050 670.050 ;
        RECT 149.250 668.850 150.750 669.750 ;
        RECT 151.950 667.950 154.050 670.050 ;
        RECT 155.250 668.850 157.050 669.750 ;
        RECT 160.950 668.850 163.050 669.750 ;
        RECT 166.950 668.850 169.050 669.750 ;
        RECT 145.950 665.850 148.050 666.750 ;
        RECT 170.400 655.050 171.450 691.950 ;
        RECT 173.400 679.050 174.450 695.400 ;
        RECT 175.950 694.950 178.050 697.050 ;
        RECT 181.950 694.950 184.050 697.050 ;
        RECT 190.950 694.950 193.050 697.050 ;
        RECT 176.400 694.050 177.450 694.950 ;
        RECT 175.950 691.950 178.050 694.050 ;
        RECT 193.950 691.950 196.050 694.050 ;
        RECT 187.950 679.950 190.050 682.050 ;
        RECT 172.950 676.950 175.050 679.050 ;
        RECT 175.950 676.950 178.050 679.050 ;
        RECT 176.400 673.050 177.450 676.950 ;
        RECT 184.950 673.950 187.050 676.050 ;
        RECT 185.400 673.050 186.450 673.950 ;
        RECT 172.950 670.950 175.050 673.050 ;
        RECT 175.950 670.950 178.050 673.050 ;
        RECT 178.950 670.950 181.050 673.050 ;
        RECT 182.250 671.250 183.750 672.150 ;
        RECT 184.950 670.950 187.050 673.050 ;
        RECT 173.400 667.050 174.450 670.950 ;
        RECT 175.950 667.950 178.050 670.050 ;
        RECT 179.250 668.850 180.750 669.750 ;
        RECT 181.950 667.950 184.050 670.050 ;
        RECT 185.250 668.850 187.050 669.750 ;
        RECT 182.400 667.050 183.450 667.950 ;
        RECT 188.400 667.050 189.450 679.950 ;
        RECT 194.400 673.050 195.450 691.950 ;
        RECT 197.400 676.050 198.450 703.950 ;
        RECT 200.400 703.050 201.450 704.400 ;
        RECT 202.950 703.950 205.050 704.400 ;
        RECT 206.250 704.250 207.750 705.150 ;
        RECT 208.950 704.400 213.450 705.450 ;
        RECT 208.950 703.950 211.050 704.400 ;
        RECT 199.950 700.950 202.050 703.050 ;
        RECT 202.950 701.850 204.750 702.750 ;
        RECT 205.950 700.950 208.050 703.050 ;
        RECT 209.250 701.850 211.050 702.750 ;
        RECT 202.950 697.950 205.050 700.050 ;
        RECT 196.950 673.950 199.050 676.050 ;
        RECT 199.950 673.950 202.050 676.050 ;
        RECT 200.400 673.050 201.450 673.950 ;
        RECT 190.950 670.950 193.050 673.050 ;
        RECT 193.950 670.950 196.050 673.050 ;
        RECT 197.250 671.250 198.750 672.150 ;
        RECT 199.950 670.950 202.050 673.050 ;
        RECT 191.400 670.050 192.450 670.950 ;
        RECT 190.950 667.950 193.050 670.050 ;
        RECT 194.250 668.850 195.750 669.750 ;
        RECT 196.950 667.950 199.050 670.050 ;
        RECT 200.250 668.850 202.050 669.750 ;
        RECT 197.400 667.050 198.450 667.950 ;
        RECT 203.400 667.050 204.450 697.950 ;
        RECT 206.400 679.050 207.450 700.950 ;
        RECT 212.400 697.050 213.450 704.400 ;
        RECT 214.950 700.950 217.050 703.050 ;
        RECT 218.400 700.050 219.450 706.950 ;
        RECT 220.950 701.250 223.050 702.150 ;
        RECT 229.950 700.950 232.050 703.050 ;
        RECT 214.950 698.850 217.050 699.750 ;
        RECT 217.950 697.950 220.050 700.050 ;
        RECT 220.950 697.950 223.050 700.050 ;
        RECT 224.250 698.250 226.050 699.150 ;
        RECT 229.950 698.850 232.050 699.750 ;
        RECT 232.950 698.250 235.050 699.150 ;
        RECT 211.950 694.950 214.050 697.050 ;
        RECT 221.400 691.050 222.450 697.950 ;
        RECT 223.950 694.950 226.050 697.050 ;
        RECT 232.950 694.950 235.050 697.050 ;
        RECT 224.400 694.050 225.450 694.950 ;
        RECT 223.950 691.950 226.050 694.050 ;
        RECT 220.950 688.950 223.050 691.050 ;
        RECT 223.950 682.950 226.050 685.050 ;
        RECT 208.950 679.950 211.050 682.050 ;
        RECT 205.950 676.950 208.050 679.050 ;
        RECT 209.400 676.050 210.450 679.950 ;
        RECT 208.950 673.950 211.050 676.050 ;
        RECT 224.400 673.050 225.450 682.950 ;
        RECT 239.400 678.450 240.450 709.950 ;
        RECT 277.950 706.950 280.050 709.050 ;
        RECT 298.950 706.950 301.050 709.050 ;
        RECT 307.950 706.950 310.050 709.050 ;
        RECT 328.950 706.950 331.050 709.050 ;
        RECT 241.950 704.250 244.050 705.150 ;
        RECT 262.950 703.950 265.050 706.050 ;
        RECT 241.950 700.950 244.050 703.050 ;
        RECT 245.250 701.250 246.750 702.150 ;
        RECT 247.950 700.950 250.050 703.050 ;
        RECT 251.250 701.250 253.050 702.150 ;
        RECT 253.950 701.250 256.050 702.150 ;
        RECT 259.950 701.250 262.050 702.150 ;
        RECT 242.400 694.050 243.450 700.950 ;
        RECT 244.950 697.950 247.050 700.050 ;
        RECT 248.250 698.850 249.750 699.750 ;
        RECT 257.250 698.250 258.750 699.150 ;
        RECT 259.950 697.950 262.050 700.050 ;
        RECT 263.400 697.050 264.450 703.950 ;
        RECT 278.400 703.050 279.450 706.950 ;
        RECT 283.950 704.250 286.050 705.150 ;
        RECT 268.950 702.450 271.050 703.050 ;
        RECT 266.400 701.400 271.050 702.450 ;
        RECT 266.400 700.050 267.450 701.400 ;
        RECT 268.950 700.950 271.050 701.400 ;
        RECT 274.950 701.250 276.750 702.150 ;
        RECT 277.950 700.950 280.050 703.050 ;
        RECT 281.250 701.250 282.750 702.150 ;
        RECT 289.950 701.250 292.050 702.150 ;
        RECT 295.950 701.250 298.050 702.150 ;
        RECT 265.950 697.950 268.050 700.050 ;
        RECT 268.950 698.850 271.050 699.750 ;
        RECT 271.950 698.250 274.050 699.150 ;
        RECT 274.950 697.950 277.050 700.050 ;
        RECT 278.250 698.850 279.750 699.750 ;
        RECT 280.950 697.950 283.050 700.050 ;
        RECT 289.950 697.950 292.050 700.050 ;
        RECT 293.250 698.250 294.750 699.150 ;
        RECT 295.950 697.950 298.050 700.050 ;
        RECT 256.950 694.950 259.050 697.050 ;
        RECT 262.950 694.950 265.050 697.050 ;
        RECT 271.950 694.950 274.050 697.050 ;
        RECT 241.950 691.950 244.050 694.050 ;
        RECT 239.400 677.400 243.450 678.450 ;
        RECT 226.950 673.950 229.050 676.050 ;
        RECT 238.950 673.950 241.050 676.050 ;
        RECT 227.400 673.050 228.450 673.950 ;
        RECT 239.400 673.050 240.450 673.950 ;
        RECT 205.950 671.250 208.050 672.150 ;
        RECT 208.950 671.850 211.050 672.750 ;
        RECT 211.950 670.950 214.050 673.050 ;
        RECT 214.950 672.450 217.050 673.050 ;
        RECT 217.950 672.450 220.050 673.050 ;
        RECT 214.950 671.400 220.050 672.450 ;
        RECT 214.950 670.950 217.050 671.400 ;
        RECT 217.950 670.950 220.050 671.400 ;
        RECT 221.250 671.250 222.750 672.150 ;
        RECT 223.950 670.950 226.050 673.050 ;
        RECT 226.950 670.950 229.050 673.050 ;
        RECT 230.250 671.250 231.750 672.150 ;
        RECT 232.950 670.950 235.050 673.050 ;
        RECT 236.250 671.250 237.750 672.150 ;
        RECT 238.950 670.950 241.050 673.050 ;
        RECT 205.950 667.950 208.050 670.050 ;
        RECT 172.950 664.950 175.050 667.050 ;
        RECT 175.950 665.850 178.050 666.750 ;
        RECT 181.950 664.950 184.050 667.050 ;
        RECT 187.950 664.950 190.050 667.050 ;
        RECT 190.950 665.850 193.050 666.750 ;
        RECT 196.950 664.950 199.050 667.050 ;
        RECT 202.950 664.950 205.050 667.050 ;
        RECT 208.950 664.950 211.050 667.050 ;
        RECT 172.950 661.950 175.050 664.050 ;
        RECT 169.950 652.950 172.050 655.050 ;
        RECT 169.950 640.950 172.050 643.050 ;
        RECT 142.950 634.950 145.050 637.050 ;
        RECT 142.950 632.250 145.050 633.150 ;
        RECT 154.950 631.950 157.050 634.050 ;
        RECT 157.950 632.250 160.050 633.150 ;
        RECT 142.950 630.450 145.050 631.050 ;
        RECT 140.400 629.400 145.050 630.450 ;
        RECT 142.950 628.950 145.050 629.400 ;
        RECT 146.250 629.250 147.750 630.150 ;
        RECT 148.950 628.950 151.050 631.050 ;
        RECT 152.250 629.250 154.050 630.150 ;
        RECT 118.950 626.400 123.450 627.450 ;
        RECT 118.950 625.950 121.050 626.400 ;
        RECT 113.400 625.050 114.450 625.950 ;
        RECT 112.950 622.950 115.050 625.050 ;
        RECT 109.950 619.950 112.050 622.050 ;
        RECT 94.950 607.950 97.050 610.050 ;
        RECT 106.950 607.950 109.050 610.050 ;
        RECT 115.950 607.950 118.050 610.050 ;
        RECT 88.950 604.950 91.050 607.050 ;
        RECT 89.400 604.050 90.450 604.950 ;
        RECT 88.950 601.950 91.050 604.050 ;
        RECT 82.950 598.950 85.050 601.050 ;
        RECT 86.250 599.250 88.050 600.150 ;
        RECT 88.950 599.850 91.050 600.750 ;
        RECT 91.950 599.250 94.050 600.150 ;
        RECT 82.950 596.850 84.750 597.750 ;
        RECT 85.950 595.950 88.050 598.050 ;
        RECT 88.950 595.950 91.050 598.050 ;
        RECT 91.950 597.450 94.050 598.050 ;
        RECT 95.400 597.450 96.450 607.950 ;
        RECT 116.400 604.050 117.450 607.950 ;
        RECT 115.950 601.950 118.050 604.050 ;
        RECT 97.950 599.250 100.050 600.150 ;
        RECT 100.950 599.850 103.050 600.750 ;
        RECT 115.950 599.850 118.050 600.750 ;
        RECT 118.950 599.250 121.050 600.150 ;
        RECT 91.950 596.400 96.450 597.450 ;
        RECT 91.950 595.950 94.050 596.400 ;
        RECT 97.950 595.950 100.050 598.050 ;
        RECT 100.950 595.950 103.050 598.050 ;
        RECT 103.950 596.250 105.750 597.150 ;
        RECT 106.950 595.950 109.050 598.050 ;
        RECT 110.250 596.250 112.050 597.150 ;
        RECT 118.950 595.950 121.050 598.050 ;
        RECT 86.400 595.050 87.450 595.950 ;
        RECT 85.950 592.950 88.050 595.050 ;
        RECT 79.950 583.950 82.050 586.050 ;
        RECT 80.400 571.050 81.450 583.950 ;
        RECT 89.400 577.050 90.450 595.950 ;
        RECT 98.400 595.050 99.450 595.950 ;
        RECT 97.950 592.950 100.050 595.050 ;
        RECT 88.950 574.950 91.050 577.050 ;
        RECT 79.950 568.950 82.050 571.050 ;
        RECT 88.950 568.950 91.050 571.050 ;
        RECT 76.950 562.950 79.050 565.050 ;
        RECT 80.400 559.050 81.450 568.950 ;
        RECT 89.400 559.050 90.450 568.950 ;
        RECT 91.950 562.950 94.050 565.050 ;
        RECT 76.950 558.450 79.050 559.050 ;
        RECT 74.400 557.400 79.050 558.450 ;
        RECT 76.950 556.950 79.050 557.400 ;
        RECT 79.950 556.950 82.050 559.050 ;
        RECT 82.950 556.950 85.050 559.050 ;
        RECT 86.250 557.250 88.050 558.150 ;
        RECT 88.950 556.950 91.050 559.050 ;
        RECT 92.400 558.450 93.450 562.950 ;
        RECT 94.950 560.250 97.050 561.150 ;
        RECT 101.400 559.050 102.450 595.950 ;
        RECT 107.250 593.850 108.750 594.750 ;
        RECT 109.950 592.950 112.050 595.050 ;
        RECT 110.400 589.050 111.450 592.950 ;
        RECT 109.950 586.950 112.050 589.050 ;
        RECT 119.400 580.050 120.450 595.950 ;
        RECT 118.950 577.950 121.050 580.050 ;
        RECT 106.950 574.950 109.050 577.050 ;
        RECT 107.400 571.050 108.450 574.950 ;
        RECT 106.950 568.950 109.050 571.050 ;
        RECT 94.950 558.450 97.050 559.050 ;
        RECT 92.400 557.400 97.050 558.450 ;
        RECT 49.950 553.950 52.050 556.050 ;
        RECT 53.250 554.850 55.050 555.750 ;
        RECT 55.950 554.250 58.050 555.150 ;
        RECT 58.950 554.850 61.050 555.750 ;
        RECT 61.950 553.950 64.050 556.050 ;
        RECT 65.250 554.850 66.750 555.750 ;
        RECT 67.950 553.950 70.050 556.050 ;
        RECT 76.950 554.850 79.050 555.750 ;
        RECT 79.950 554.250 82.050 555.150 ;
        RECT 82.950 554.850 84.750 555.750 ;
        RECT 85.950 553.950 88.050 556.050 ;
        RECT 40.950 550.950 43.050 553.050 ;
        RECT 46.950 550.950 49.050 553.050 ;
        RECT 55.950 550.950 58.050 553.050 ;
        RECT 79.950 550.950 82.050 553.050 ;
        RECT 86.400 541.050 87.450 553.950 ;
        RECT 92.400 553.050 93.450 557.400 ;
        RECT 94.950 556.950 97.050 557.400 ;
        RECT 98.250 557.250 99.750 558.150 ;
        RECT 100.950 556.950 103.050 559.050 ;
        RECT 104.250 557.250 106.050 558.150 ;
        RECT 97.950 553.950 100.050 556.050 ;
        RECT 101.250 554.850 102.750 555.750 ;
        RECT 103.950 555.450 106.050 556.050 ;
        RECT 107.400 555.450 108.450 568.950 ;
        RECT 122.400 562.050 123.450 626.400 ;
        RECT 124.950 625.950 127.050 628.050 ;
        RECT 128.250 626.850 130.050 627.750 ;
        RECT 130.950 626.250 133.050 627.150 ;
        RECT 133.950 626.850 136.050 627.750 ;
        RECT 137.400 625.050 138.450 628.950 ;
        RECT 142.950 627.450 145.050 628.050 ;
        RECT 145.950 627.450 148.050 628.050 ;
        RECT 142.950 626.400 148.050 627.450 ;
        RECT 149.250 626.850 150.750 627.750 ;
        RECT 151.950 627.450 154.050 628.050 ;
        RECT 155.400 627.450 156.450 631.950 ;
        RECT 157.950 628.950 160.050 631.050 ;
        RECT 161.250 629.250 162.750 630.150 ;
        RECT 163.950 628.950 166.050 631.050 ;
        RECT 167.250 629.250 169.050 630.150 ;
        RECT 142.950 625.950 145.050 626.400 ;
        RECT 145.950 625.950 148.050 626.400 ;
        RECT 151.950 626.400 156.450 627.450 ;
        RECT 151.950 625.950 154.050 626.400 ;
        RECT 130.950 622.950 133.050 625.050 ;
        RECT 136.950 622.950 139.050 625.050 ;
        RECT 152.400 619.050 153.450 625.950 ;
        RECT 145.950 616.950 148.050 619.050 ;
        RECT 151.950 616.950 154.050 619.050 ;
        RECT 146.400 601.050 147.450 616.950 ;
        RECT 127.950 600.450 130.050 601.050 ;
        RECT 125.400 599.400 130.050 600.450 ;
        RECT 125.400 565.050 126.450 599.400 ;
        RECT 127.950 598.950 130.050 599.400 ;
        RECT 145.950 598.950 148.050 601.050 ;
        RECT 127.950 596.850 130.050 597.750 ;
        RECT 133.950 596.850 136.050 597.750 ;
        RECT 139.950 596.850 142.050 597.750 ;
        RECT 145.950 596.850 148.050 597.750 ;
        RECT 139.950 571.950 142.050 574.050 ;
        RECT 124.950 562.950 127.050 565.050 ;
        RECT 125.400 562.050 126.450 562.950 ;
        RECT 109.950 560.250 112.050 561.150 ;
        RECT 121.950 559.950 124.050 562.050 ;
        RECT 124.950 559.950 127.050 562.050 ;
        RECT 127.950 559.950 130.050 562.050 ;
        RECT 133.950 560.250 136.050 561.150 ;
        RECT 128.400 559.050 129.450 559.950 ;
        RECT 140.400 559.050 141.450 571.950 ;
        RECT 152.400 568.050 153.450 616.950 ;
        RECT 158.400 598.050 159.450 628.950 ;
        RECT 160.950 625.950 163.050 628.050 ;
        RECT 164.250 626.850 165.750 627.750 ;
        RECT 166.950 625.950 169.050 628.050 ;
        RECT 161.400 622.050 162.450 625.950 ;
        RECT 167.400 622.050 168.450 625.950 ;
        RECT 160.950 619.950 163.050 622.050 ;
        RECT 166.950 619.950 169.050 622.050 ;
        RECT 170.400 613.050 171.450 640.950 ;
        RECT 173.400 637.050 174.450 661.950 ;
        RECT 203.400 640.050 204.450 664.950 ;
        RECT 209.400 661.050 210.450 664.950 ;
        RECT 208.950 658.950 211.050 661.050 ;
        RECT 212.400 658.050 213.450 670.950 ;
        RECT 214.950 667.950 217.050 670.050 ;
        RECT 218.250 668.850 219.750 669.750 ;
        RECT 220.950 667.950 223.050 670.050 ;
        RECT 224.250 668.850 226.050 669.750 ;
        RECT 226.950 668.850 228.750 669.750 ;
        RECT 229.950 667.950 232.050 670.050 ;
        RECT 233.250 668.850 234.750 669.750 ;
        RECT 235.950 667.950 238.050 670.050 ;
        RECT 239.250 668.850 241.050 669.750 ;
        RECT 221.400 667.050 222.450 667.950 ;
        RECT 214.950 665.850 217.050 666.750 ;
        RECT 220.950 664.950 223.050 667.050 ;
        RECT 230.400 661.050 231.450 667.950 ;
        RECT 232.950 661.950 235.050 664.050 ;
        RECT 229.950 658.950 232.050 661.050 ;
        RECT 211.950 655.950 214.050 658.050 ;
        RECT 217.950 655.950 220.050 658.050 ;
        RECT 202.950 637.950 205.050 640.050 ;
        RECT 205.950 637.950 208.050 640.050 ;
        RECT 172.950 634.950 175.050 637.050 ;
        RECT 181.950 636.450 184.050 637.050 ;
        RECT 184.950 636.450 187.050 637.050 ;
        RECT 181.950 635.400 187.050 636.450 ;
        RECT 181.950 634.950 184.050 635.400 ;
        RECT 184.950 634.950 187.050 635.400 ;
        RECT 187.950 633.450 190.050 634.050 ;
        RECT 172.950 632.250 175.050 633.150 ;
        RECT 185.400 632.400 190.050 633.450 ;
        RECT 193.950 633.450 196.050 634.050 ;
        RECT 172.950 628.950 175.050 631.050 ;
        RECT 176.250 629.250 177.750 630.150 ;
        RECT 178.950 628.950 181.050 631.050 ;
        RECT 182.250 629.250 184.050 630.150 ;
        RECT 172.950 625.950 175.050 628.050 ;
        RECT 175.950 625.950 178.050 628.050 ;
        RECT 179.250 626.850 180.750 627.750 ;
        RECT 181.950 625.950 184.050 628.050 ;
        RECT 173.400 619.050 174.450 625.950 ;
        RECT 176.400 622.050 177.450 625.950 ;
        RECT 182.400 625.050 183.450 625.950 ;
        RECT 185.400 625.050 186.450 632.400 ;
        RECT 187.950 631.950 190.050 632.400 ;
        RECT 191.250 632.250 192.750 633.150 ;
        RECT 193.950 632.400 198.450 633.450 ;
        RECT 193.950 631.950 196.050 632.400 ;
        RECT 197.400 631.050 198.450 632.400 ;
        RECT 206.400 631.050 207.450 637.950 ;
        RECT 211.950 634.950 214.050 637.050 ;
        RECT 212.400 631.050 213.450 634.950 ;
        RECT 218.400 634.050 219.450 655.950 ;
        RECT 229.950 637.950 232.050 640.050 ;
        RECT 223.950 634.950 226.050 637.050 ;
        RECT 224.400 634.050 225.450 634.950 ;
        RECT 230.400 634.050 231.450 637.950 ;
        RECT 217.950 631.950 220.050 634.050 ;
        RECT 223.950 631.950 226.050 634.050 ;
        RECT 229.950 631.950 232.050 634.050 ;
        RECT 187.950 629.850 189.750 630.750 ;
        RECT 190.950 628.950 193.050 631.050 ;
        RECT 194.250 629.850 196.050 630.750 ;
        RECT 196.950 628.950 199.050 631.050 ;
        RECT 199.950 628.950 202.050 631.050 ;
        RECT 202.950 629.250 204.750 630.150 ;
        RECT 205.950 628.950 208.050 631.050 ;
        RECT 209.250 629.250 210.750 630.150 ;
        RECT 211.950 628.950 214.050 631.050 ;
        RECT 215.250 629.250 217.050 630.150 ;
        RECT 181.950 622.950 184.050 625.050 ;
        RECT 184.950 622.950 187.050 625.050 ;
        RECT 187.950 622.950 190.050 625.050 ;
        RECT 175.950 619.950 178.050 622.050 ;
        RECT 172.950 616.950 175.050 619.050 ;
        RECT 169.950 610.950 172.050 613.050 ;
        RECT 188.400 604.050 189.450 622.950 ;
        RECT 191.400 622.050 192.450 628.950 ;
        RECT 197.400 625.050 198.450 628.950 ;
        RECT 200.400 628.050 201.450 628.950 ;
        RECT 199.950 625.950 202.050 628.050 ;
        RECT 202.950 625.950 205.050 628.050 ;
        RECT 206.250 626.850 207.750 627.750 ;
        RECT 208.950 625.950 211.050 628.050 ;
        RECT 212.250 626.850 213.750 627.750 ;
        RECT 214.950 625.950 217.050 628.050 ;
        RECT 193.950 622.950 196.050 625.050 ;
        RECT 196.950 622.950 199.050 625.050 ;
        RECT 190.950 619.950 193.050 622.050 ;
        RECT 169.950 601.950 172.050 604.050 ;
        RECT 181.950 601.950 184.050 604.050 ;
        RECT 187.950 601.950 190.050 604.050 ;
        RECT 166.950 600.450 169.050 601.050 ;
        RECT 164.400 599.400 169.050 600.450 ;
        RECT 170.250 599.850 171.750 600.750 ;
        RECT 172.950 600.450 175.050 601.050 ;
        RECT 154.950 596.250 156.750 597.150 ;
        RECT 157.950 595.950 160.050 598.050 ;
        RECT 161.250 596.250 163.050 597.150 ;
        RECT 164.400 595.050 165.450 599.400 ;
        RECT 166.950 598.950 169.050 599.400 ;
        RECT 172.950 599.400 177.450 600.450 ;
        RECT 172.950 598.950 175.050 599.400 ;
        RECT 166.950 596.850 169.050 597.750 ;
        RECT 169.950 595.950 172.050 598.050 ;
        RECT 172.950 596.850 175.050 597.750 ;
        RECT 176.400 597.450 177.450 599.400 ;
        RECT 178.950 599.250 181.050 600.150 ;
        RECT 181.950 599.850 184.050 600.750 ;
        RECT 178.950 597.450 181.050 598.050 ;
        RECT 176.400 596.400 181.050 597.450 ;
        RECT 178.950 595.950 181.050 596.400 ;
        RECT 184.950 596.250 186.750 597.150 ;
        RECT 187.950 595.950 190.050 598.050 ;
        RECT 191.250 596.250 193.050 597.150 ;
        RECT 154.950 592.950 157.050 595.050 ;
        RECT 158.250 593.850 159.750 594.750 ;
        RECT 163.950 592.950 166.050 595.050 ;
        RECT 166.950 592.950 169.050 595.050 ;
        RECT 155.400 577.050 156.450 592.950 ;
        RECT 163.950 583.950 166.050 586.050 ;
        RECT 154.950 574.950 157.050 577.050 ;
        RECT 151.950 565.950 154.050 568.050 ;
        RECT 154.950 565.950 157.050 568.050 ;
        RECT 142.950 560.250 145.050 561.150 ;
        RECT 148.950 559.950 151.050 562.050 ;
        RECT 149.400 559.050 150.450 559.950 ;
        RECT 109.950 556.950 112.050 559.050 ;
        RECT 113.250 557.250 114.750 558.150 ;
        RECT 115.950 556.950 118.050 559.050 ;
        RECT 119.250 557.250 121.050 558.150 ;
        RECT 121.950 556.950 124.050 559.050 ;
        RECT 124.950 557.250 126.750 558.150 ;
        RECT 127.950 556.950 130.050 559.050 ;
        RECT 131.250 557.250 132.750 558.150 ;
        RECT 133.950 556.950 136.050 559.050 ;
        RECT 139.950 556.950 142.050 559.050 ;
        RECT 142.950 556.950 145.050 559.050 ;
        RECT 146.250 557.250 147.750 558.150 ;
        RECT 148.950 556.950 151.050 559.050 ;
        RECT 152.250 557.250 154.050 558.150 ;
        RECT 103.950 554.400 108.450 555.450 ;
        RECT 103.950 553.950 106.050 554.400 ;
        RECT 112.950 553.950 115.050 556.050 ;
        RECT 116.250 554.850 117.750 555.750 ;
        RECT 118.950 553.950 121.050 556.050 ;
        RECT 91.950 550.950 94.050 553.050 ;
        RECT 88.950 547.950 91.050 550.050 ;
        RECT 85.950 538.950 88.050 541.050 ;
        RECT 37.950 532.950 40.050 535.050 ;
        RECT 43.950 532.950 46.050 535.050 ;
        RECT 58.950 532.950 61.050 535.050 ;
        RECT 73.950 532.950 76.050 535.050 ;
        RECT 44.400 532.050 45.450 532.950 ;
        RECT 22.950 529.950 25.050 532.050 ;
        RECT 28.950 529.950 31.050 532.050 ;
        RECT 43.950 529.950 46.050 532.050 ;
        RECT 49.950 529.950 52.050 532.050 ;
        RECT 13.950 528.450 16.050 529.050 ;
        RECT 22.950 528.450 25.050 529.050 ;
        RECT 13.950 527.400 18.450 528.450 ;
        RECT 13.950 526.950 16.050 527.400 ;
        RECT 7.950 524.850 10.050 525.750 ;
        RECT 13.950 524.850 16.050 525.750 ;
        RECT 17.400 505.050 18.450 527.400 ;
        RECT 20.400 527.400 25.050 528.450 ;
        RECT 16.950 502.950 19.050 505.050 ;
        RECT 20.400 496.050 21.450 527.400 ;
        RECT 22.950 526.950 25.050 527.400 ;
        RECT 26.250 527.250 28.050 528.150 ;
        RECT 28.950 527.850 31.050 528.750 ;
        RECT 31.950 527.250 34.050 528.150 ;
        RECT 40.950 527.250 43.050 528.150 ;
        RECT 43.950 527.850 46.050 528.750 ;
        RECT 50.400 526.050 51.450 529.950 ;
        RECT 59.400 529.050 60.450 532.950 ;
        RECT 52.950 526.950 55.050 529.050 ;
        RECT 56.250 527.250 57.750 528.150 ;
        RECT 58.950 526.950 61.050 529.050 ;
        RECT 61.950 528.450 64.050 529.050 ;
        RECT 64.950 528.450 67.050 529.050 ;
        RECT 61.950 527.400 67.050 528.450 ;
        RECT 61.950 526.950 64.050 527.400 ;
        RECT 64.950 526.950 67.050 527.400 ;
        RECT 22.950 524.850 24.750 525.750 ;
        RECT 25.950 523.950 28.050 526.050 ;
        RECT 31.950 523.950 34.050 526.050 ;
        RECT 40.950 523.950 43.050 526.050 ;
        RECT 43.950 523.950 46.050 526.050 ;
        RECT 49.950 523.950 52.050 526.050 ;
        RECT 53.250 524.850 54.750 525.750 ;
        RECT 55.950 523.950 58.050 526.050 ;
        RECT 59.250 524.850 61.050 525.750 ;
        RECT 61.950 523.950 64.050 526.050 ;
        RECT 64.950 524.250 66.750 525.150 ;
        RECT 67.950 523.950 70.050 526.050 ;
        RECT 71.250 524.250 73.050 525.150 ;
        RECT 13.950 493.950 16.050 496.050 ;
        RECT 19.950 493.950 22.050 496.050 ;
        RECT 7.950 487.950 10.050 490.050 ;
        RECT 8.400 487.050 9.450 487.950 ;
        RECT 7.950 484.950 10.050 487.050 ;
        RECT 7.950 482.850 10.050 483.750 ;
        RECT 10.950 482.250 13.050 483.150 ;
        RECT 10.950 478.950 13.050 481.050 ;
        RECT 11.400 478.050 12.450 478.950 ;
        RECT 10.950 475.950 13.050 478.050 ;
        RECT 7.950 457.950 10.050 460.050 ;
        RECT 14.400 457.050 15.450 493.950 ;
        RECT 16.950 490.950 19.050 493.050 ;
        RECT 17.400 490.050 18.450 490.950 ;
        RECT 16.950 487.950 19.050 490.050 ;
        RECT 20.250 488.250 21.750 489.150 ;
        RECT 22.950 487.950 25.050 490.050 ;
        RECT 26.400 487.050 27.450 523.950 ;
        RECT 32.400 517.050 33.450 523.950 ;
        RECT 41.400 520.050 42.450 523.950 ;
        RECT 40.950 517.950 43.050 520.050 ;
        RECT 31.950 514.950 34.050 517.050 ;
        RECT 40.950 514.950 43.050 517.050 ;
        RECT 41.400 487.050 42.450 514.950 ;
        RECT 16.950 485.850 18.750 486.750 ;
        RECT 19.950 484.950 22.050 487.050 ;
        RECT 23.250 485.850 25.050 486.750 ;
        RECT 25.950 484.950 28.050 487.050 ;
        RECT 28.950 484.950 31.050 487.050 ;
        RECT 31.950 485.250 33.750 486.150 ;
        RECT 34.950 484.950 37.050 487.050 ;
        RECT 40.950 484.950 43.050 487.050 ;
        RECT 29.400 478.050 30.450 484.950 ;
        RECT 31.950 481.950 34.050 484.050 ;
        RECT 35.250 482.850 37.050 483.750 ;
        RECT 37.950 482.250 40.050 483.150 ;
        RECT 40.950 482.850 43.050 483.750 ;
        RECT 28.950 475.950 31.050 478.050 ;
        RECT 16.950 460.950 19.050 463.050 ;
        RECT 25.950 460.950 28.050 463.050 ;
        RECT 17.400 457.050 18.450 460.950 ;
        RECT 26.400 457.050 27.450 460.950 ;
        RECT 4.950 455.250 7.050 456.150 ;
        RECT 7.950 455.850 10.050 456.750 ;
        RECT 13.950 454.950 16.050 457.050 ;
        RECT 16.950 454.950 19.050 457.050 ;
        RECT 20.250 455.250 21.750 456.150 ;
        RECT 22.950 454.950 25.050 457.050 ;
        RECT 25.950 454.950 28.050 457.050 ;
        RECT 32.400 456.450 33.450 481.950 ;
        RECT 44.400 481.050 45.450 523.950 ;
        RECT 49.950 521.850 52.050 522.750 ;
        RECT 55.950 520.950 58.050 523.050 ;
        RECT 58.950 520.950 61.050 523.050 ;
        RECT 62.400 522.450 63.450 523.950 ;
        RECT 74.400 523.050 75.450 532.950 ;
        RECT 86.400 532.050 87.450 538.950 ;
        RECT 85.950 529.950 88.050 532.050 ;
        RECT 79.950 526.950 82.050 529.050 ;
        RECT 83.250 527.250 84.750 528.150 ;
        RECT 85.950 526.950 88.050 529.050 ;
        RECT 76.950 523.950 79.050 526.050 ;
        RECT 80.250 524.850 81.750 525.750 ;
        RECT 82.950 523.950 85.050 526.050 ;
        RECT 86.250 524.850 88.050 525.750 ;
        RECT 64.950 522.450 67.050 523.050 ;
        RECT 62.400 521.400 67.050 522.450 ;
        RECT 68.250 521.850 69.750 522.750 ;
        RECT 64.950 520.950 67.050 521.400 ;
        RECT 70.950 520.950 73.050 523.050 ;
        RECT 73.950 520.950 76.050 523.050 ;
        RECT 76.950 521.850 79.050 522.750 ;
        RECT 46.950 496.950 49.050 499.050 ;
        RECT 47.400 490.050 48.450 496.950 ;
        RECT 56.400 496.050 57.450 520.950 ;
        RECT 59.400 514.050 60.450 520.950 ;
        RECT 61.950 517.950 64.050 520.050 ;
        RECT 62.400 517.050 63.450 517.950 ;
        RECT 65.400 517.050 66.450 520.950 ;
        RECT 71.400 520.050 72.450 520.950 ;
        RECT 70.950 517.950 73.050 520.050 ;
        RECT 61.950 514.950 64.050 517.050 ;
        RECT 64.950 514.950 67.050 517.050 ;
        RECT 58.950 511.950 61.050 514.050 ;
        RECT 62.400 499.050 63.450 514.950 ;
        RECT 89.400 502.050 90.450 547.950 ;
        RECT 98.400 538.050 99.450 553.950 ;
        RECT 97.950 535.950 100.050 538.050 ;
        RECT 100.950 531.450 103.050 532.050 ;
        RECT 92.400 530.400 103.050 531.450 ;
        RECT 92.400 529.050 93.450 530.400 ;
        RECT 100.950 529.950 103.050 530.400 ;
        RECT 101.400 529.050 102.450 529.950 ;
        RECT 91.950 526.950 94.050 529.050 ;
        RECT 94.950 526.950 97.050 529.050 ;
        RECT 98.250 527.250 99.750 528.150 ;
        RECT 100.950 526.950 103.050 529.050 ;
        RECT 113.400 526.050 114.450 553.950 ;
        RECT 122.400 547.050 123.450 556.950 ;
        RECT 124.950 553.950 127.050 556.050 ;
        RECT 128.250 554.850 129.750 555.750 ;
        RECT 130.950 553.950 133.050 556.050 ;
        RECT 125.400 553.050 126.450 553.950 ;
        RECT 124.950 550.950 127.050 553.050 ;
        RECT 125.400 550.050 126.450 550.950 ;
        RECT 124.950 547.950 127.050 550.050 ;
        RECT 131.400 547.050 132.450 553.950 ;
        RECT 140.400 553.050 141.450 556.950 ;
        RECT 143.400 556.050 144.450 556.950 ;
        RECT 142.950 553.950 145.050 556.050 ;
        RECT 145.950 553.950 148.050 556.050 ;
        RECT 149.250 554.850 150.750 555.750 ;
        RECT 151.950 553.950 154.050 556.050 ;
        RECT 139.950 550.950 142.050 553.050 ;
        RECT 146.400 550.050 147.450 553.950 ;
        RECT 152.400 553.050 153.450 553.950 ;
        RECT 151.950 550.950 154.050 553.050 ;
        RECT 139.950 547.950 142.050 550.050 ;
        RECT 145.950 547.950 148.050 550.050 ;
        RECT 118.950 544.950 121.050 547.050 ;
        RECT 121.950 544.950 124.050 547.050 ;
        RECT 127.950 544.950 130.050 547.050 ;
        RECT 130.950 544.950 133.050 547.050 ;
        RECT 136.950 544.950 139.050 547.050 ;
        RECT 119.400 532.050 120.450 544.950 ;
        RECT 128.400 532.050 129.450 544.950 ;
        RECT 137.400 532.050 138.450 544.950 ;
        RECT 118.950 529.950 121.050 532.050 ;
        RECT 127.950 529.950 130.050 532.050 ;
        RECT 130.950 529.950 133.050 532.050 ;
        RECT 136.950 529.950 139.050 532.050 ;
        RECT 115.950 527.250 118.050 528.150 ;
        RECT 118.950 527.850 121.050 528.750 ;
        RECT 124.950 528.450 127.050 529.050 ;
        RECT 121.950 527.250 123.750 528.150 ;
        RECT 124.950 527.400 129.450 528.450 ;
        RECT 124.950 526.950 127.050 527.400 ;
        RECT 91.950 523.950 94.050 526.050 ;
        RECT 95.250 524.850 96.750 525.750 ;
        RECT 97.950 523.950 100.050 526.050 ;
        RECT 101.250 524.850 103.050 525.750 ;
        RECT 103.950 524.250 105.750 525.150 ;
        RECT 106.950 523.950 109.050 526.050 ;
        RECT 110.250 524.250 112.050 525.150 ;
        RECT 112.950 523.950 115.050 526.050 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 121.950 523.950 124.050 526.050 ;
        RECT 125.250 524.850 127.050 525.750 ;
        RECT 91.950 521.850 94.050 522.750 ;
        RECT 103.950 520.950 106.050 523.050 ;
        RECT 107.250 521.850 108.750 522.750 ;
        RECT 109.950 520.950 112.050 523.050 ;
        RECT 112.950 520.950 115.050 523.050 ;
        RECT 110.400 514.050 111.450 520.950 ;
        RECT 109.950 511.950 112.050 514.050 ;
        RECT 88.950 499.950 91.050 502.050 ;
        RECT 58.950 496.950 61.050 499.050 ;
        RECT 61.950 496.950 64.050 499.050 ;
        RECT 76.950 496.950 79.050 499.050 ;
        RECT 59.400 496.050 60.450 496.950 ;
        RECT 55.950 493.950 58.050 496.050 ;
        RECT 58.950 493.950 61.050 496.050 ;
        RECT 61.950 493.950 64.050 496.050 ;
        RECT 52.950 491.250 55.050 492.150 ;
        RECT 58.950 490.950 61.050 493.050 ;
        RECT 46.950 487.950 49.050 490.050 ;
        RECT 50.250 488.250 51.750 489.150 ;
        RECT 52.950 487.950 55.050 490.050 ;
        RECT 56.250 488.250 58.050 489.150 ;
        RECT 46.950 485.850 48.750 486.750 ;
        RECT 49.950 484.950 52.050 487.050 ;
        RECT 55.950 486.450 58.050 487.050 ;
        RECT 59.400 486.450 60.450 490.950 ;
        RECT 62.400 490.050 63.450 493.950 ;
        RECT 77.400 493.050 78.450 496.950 ;
        RECT 103.950 493.950 106.050 496.050 ;
        RECT 67.950 490.950 70.050 493.050 ;
        RECT 73.950 491.250 76.050 492.150 ;
        RECT 76.950 490.950 79.050 493.050 ;
        RECT 68.400 490.050 69.450 490.950 ;
        RECT 104.400 490.050 105.450 493.950 ;
        RECT 113.400 493.050 114.450 520.950 ;
        RECT 116.400 520.050 117.450 523.950 ;
        RECT 118.950 520.950 121.050 523.050 ;
        RECT 115.950 517.950 118.050 520.050 ;
        RECT 119.400 517.050 120.450 520.950 ;
        RECT 118.950 514.950 121.050 517.050 ;
        RECT 112.950 490.950 115.050 493.050 ;
        RECT 128.400 490.050 129.450 527.400 ;
        RECT 131.400 526.050 132.450 529.950 ;
        RECT 133.950 527.250 136.050 528.150 ;
        RECT 136.950 527.850 139.050 528.750 ;
        RECT 130.950 523.950 133.050 526.050 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 140.400 523.050 141.450 547.950 ;
        RECT 148.950 544.950 151.050 547.050 ;
        RECT 149.400 532.050 150.450 544.950 ;
        RECT 151.950 535.950 154.050 538.050 ;
        RECT 152.400 532.050 153.450 535.950 ;
        RECT 155.400 535.050 156.450 565.950 ;
        RECT 164.400 562.050 165.450 583.950 ;
        RECT 167.400 583.050 168.450 592.950 ;
        RECT 170.400 583.050 171.450 595.950 ;
        RECT 166.950 580.950 169.050 583.050 ;
        RECT 169.950 580.950 172.050 583.050 ;
        RECT 179.400 574.050 180.450 595.950 ;
        RECT 188.250 593.850 189.750 594.750 ;
        RECT 190.950 592.950 193.050 595.050 ;
        RECT 187.950 580.950 190.050 583.050 ;
        RECT 190.950 580.950 193.050 583.050 ;
        RECT 184.950 577.950 187.050 580.050 ;
        RECT 169.950 571.950 172.050 574.050 ;
        RECT 178.950 571.950 181.050 574.050 ;
        RECT 170.400 568.050 171.450 571.950 ;
        RECT 166.950 565.950 169.050 568.050 ;
        RECT 169.950 565.950 172.050 568.050 ;
        RECT 163.950 559.950 166.050 562.050 ;
        RECT 167.400 559.050 168.450 565.950 ;
        RECT 181.950 562.950 184.050 565.050 ;
        RECT 178.950 560.250 181.050 561.150 ;
        RECT 157.950 557.250 159.750 558.150 ;
        RECT 160.950 556.950 163.050 559.050 ;
        RECT 166.950 556.950 169.050 559.050 ;
        RECT 169.950 557.250 171.750 558.150 ;
        RECT 172.950 556.950 175.050 559.050 ;
        RECT 176.250 557.250 177.750 558.150 ;
        RECT 178.950 556.950 181.050 559.050 ;
        RECT 179.400 556.050 180.450 556.950 ;
        RECT 157.950 553.950 160.050 556.050 ;
        RECT 161.250 554.850 163.050 555.750 ;
        RECT 163.950 554.250 166.050 555.150 ;
        RECT 166.950 554.850 169.050 555.750 ;
        RECT 169.950 553.950 172.050 556.050 ;
        RECT 173.250 554.850 174.750 555.750 ;
        RECT 175.950 553.950 178.050 556.050 ;
        RECT 178.950 553.950 181.050 556.050 ;
        RECT 163.950 550.950 166.050 553.050 ;
        RECT 169.950 552.450 172.050 553.050 ;
        RECT 176.400 552.450 177.450 553.950 ;
        RECT 169.950 551.400 177.450 552.450 ;
        RECT 169.950 550.950 172.050 551.400 ;
        RECT 164.400 550.050 165.450 550.950 ;
        RECT 163.950 547.950 166.050 550.050 ;
        RECT 175.950 547.950 178.050 550.050 ;
        RECT 160.950 544.950 163.050 547.050 ;
        RECT 166.950 544.950 169.050 547.050 ;
        RECT 154.950 532.950 157.050 535.050 ;
        RECT 161.400 532.050 162.450 544.950 ;
        RECT 167.400 532.050 168.450 544.950 ;
        RECT 148.950 529.950 151.050 532.050 ;
        RECT 151.950 529.950 154.050 532.050 ;
        RECT 154.950 529.950 157.050 532.050 ;
        RECT 160.950 529.950 163.050 532.050 ;
        RECT 166.950 529.950 169.050 532.050 ;
        RECT 142.950 526.950 145.050 529.050 ;
        RECT 146.250 527.250 148.050 528.150 ;
        RECT 148.950 527.850 151.050 528.750 ;
        RECT 151.950 527.250 154.050 528.150 ;
        RECT 154.950 527.850 157.050 528.750 ;
        RECT 157.950 527.250 160.050 528.150 ;
        RECT 142.950 524.850 144.750 525.750 ;
        RECT 145.950 523.950 148.050 526.050 ;
        RECT 151.950 523.950 154.050 526.050 ;
        RECT 157.950 525.450 160.050 526.050 ;
        RECT 161.400 525.450 162.450 529.950 ;
        RECT 163.950 527.250 166.050 528.150 ;
        RECT 166.950 527.850 169.050 528.750 ;
        RECT 169.950 527.250 171.750 528.150 ;
        RECT 172.950 526.950 175.050 529.050 ;
        RECT 157.950 524.400 162.450 525.450 ;
        RECT 157.950 523.950 160.050 524.400 ;
        RECT 163.950 523.950 166.050 526.050 ;
        RECT 166.950 523.950 169.050 526.050 ;
        RECT 169.950 523.950 172.050 526.050 ;
        RECT 173.250 524.850 175.050 525.750 ;
        RECT 130.950 520.950 133.050 523.050 ;
        RECT 139.950 520.950 142.050 523.050 ;
        RECT 131.400 514.050 132.450 520.950 ;
        RECT 130.950 511.950 133.050 514.050 ;
        RECT 160.950 505.950 163.050 508.050 ;
        RECT 142.950 499.950 145.050 502.050 ;
        RECT 61.950 487.950 64.050 490.050 ;
        RECT 65.250 488.250 66.750 489.150 ;
        RECT 67.950 487.950 70.050 490.050 ;
        RECT 70.950 488.250 72.750 489.150 ;
        RECT 73.950 487.950 76.050 490.050 ;
        RECT 77.250 488.250 78.750 489.150 ;
        RECT 79.950 487.950 82.050 490.050 ;
        RECT 94.950 488.250 97.050 489.150 ;
        RECT 100.950 487.950 103.050 490.050 ;
        RECT 103.950 487.950 106.050 490.050 ;
        RECT 109.950 489.450 112.050 490.050 ;
        RECT 107.250 488.250 108.750 489.150 ;
        RECT 109.950 488.400 114.450 489.450 ;
        RECT 109.950 487.950 112.050 488.400 ;
        RECT 55.950 485.400 60.450 486.450 ;
        RECT 61.950 485.850 63.750 486.750 ;
        RECT 55.950 484.950 58.050 485.400 ;
        RECT 64.950 484.950 67.050 487.050 ;
        RECT 68.250 485.850 70.050 486.750 ;
        RECT 70.950 484.950 73.050 487.050 ;
        RECT 76.950 484.950 79.050 487.050 ;
        RECT 80.250 485.850 82.050 486.750 ;
        RECT 82.950 484.950 85.050 487.050 ;
        RECT 85.950 485.250 87.750 486.150 ;
        RECT 88.950 484.950 91.050 487.050 ;
        RECT 92.250 485.250 93.750 486.150 ;
        RECT 94.950 484.950 97.050 487.050 ;
        RECT 46.950 481.950 49.050 484.050 ;
        RECT 52.950 481.950 55.050 484.050 ;
        RECT 37.950 478.950 40.050 481.050 ;
        RECT 43.950 478.950 46.050 481.050 ;
        RECT 47.400 477.450 48.450 481.950 ;
        RECT 44.400 476.400 48.450 477.450 ;
        RECT 40.950 466.950 43.050 469.050 ;
        RECT 29.400 455.400 33.450 456.450 ;
        RECT 34.950 456.450 37.050 457.050 ;
        RECT 34.950 455.400 39.450 456.450 ;
        RECT 4.950 451.950 7.050 454.050 ;
        RECT 13.950 451.950 16.050 454.050 ;
        RECT 17.250 452.850 18.750 453.750 ;
        RECT 19.950 451.950 22.050 454.050 ;
        RECT 23.250 452.850 25.050 453.750 ;
        RECT 25.950 452.850 28.050 453.750 ;
        RECT 13.950 449.850 16.050 450.750 ;
        RECT 25.950 430.950 28.050 433.050 ;
        RECT 10.950 421.950 13.050 424.050 ;
        RECT 4.950 412.950 7.050 415.050 ;
        RECT 4.950 410.850 7.050 411.750 ;
        RECT 7.950 410.250 10.050 411.150 ;
        RECT 7.950 408.450 10.050 409.050 ;
        RECT 11.400 408.450 12.450 421.950 ;
        RECT 13.950 416.250 16.050 417.150 ;
        RECT 13.950 412.950 16.050 415.050 ;
        RECT 17.250 413.250 18.750 414.150 ;
        RECT 19.950 412.950 22.050 415.050 ;
        RECT 23.250 413.250 25.050 414.150 ;
        RECT 16.950 409.950 19.050 412.050 ;
        RECT 20.250 410.850 21.750 411.750 ;
        RECT 22.950 409.950 25.050 412.050 ;
        RECT 7.950 407.400 12.450 408.450 ;
        RECT 7.950 406.950 10.050 407.400 ;
        RECT 17.400 406.050 18.450 409.950 ;
        RECT 16.950 403.950 19.050 406.050 ;
        RECT 26.400 391.050 27.450 430.950 ;
        RECT 29.400 417.450 30.450 455.400 ;
        RECT 34.950 454.950 37.050 455.400 ;
        RECT 31.950 452.250 34.050 453.150 ;
        RECT 34.950 452.850 37.050 453.750 ;
        RECT 31.950 448.950 34.050 451.050 ;
        RECT 38.400 430.050 39.450 455.400 ;
        RECT 37.950 427.950 40.050 430.050 ;
        RECT 29.400 416.400 33.450 417.450 ;
        RECT 32.400 415.050 33.450 416.400 ;
        RECT 37.950 416.250 40.050 417.150 ;
        RECT 28.950 413.250 30.750 414.150 ;
        RECT 31.950 412.950 34.050 415.050 ;
        RECT 37.950 414.450 40.050 415.050 ;
        RECT 41.400 414.450 42.450 466.950 ;
        RECT 44.400 436.050 45.450 476.400 ;
        RECT 49.950 453.450 52.050 454.050 ;
        RECT 53.400 453.450 54.450 481.950 ;
        RECT 55.950 460.950 58.050 463.050 ;
        RECT 56.400 460.050 57.450 460.950 ;
        RECT 55.950 457.950 58.050 460.050 ;
        RECT 58.950 457.950 61.050 460.050 ;
        RECT 56.400 454.050 57.450 457.950 ;
        RECT 58.950 455.850 61.050 456.750 ;
        RECT 61.950 455.250 64.050 456.150 ;
        RECT 65.400 454.050 66.450 484.950 ;
        RECT 71.400 481.050 72.450 484.950 ;
        RECT 70.950 478.950 73.050 481.050 ;
        RECT 79.950 478.950 82.050 481.050 ;
        RECT 73.950 466.950 76.050 469.050 ;
        RECT 74.400 460.050 75.450 466.950 ;
        RECT 73.950 457.950 76.050 460.050 ;
        RECT 70.950 455.250 73.050 456.150 ;
        RECT 73.950 455.850 76.050 456.750 ;
        RECT 80.400 454.050 81.450 478.950 ;
        RECT 83.400 469.050 84.450 484.950 ;
        RECT 85.950 481.950 88.050 484.050 ;
        RECT 89.250 482.850 90.750 483.750 ;
        RECT 91.950 481.950 94.050 484.050 ;
        RECT 86.400 481.050 87.450 481.950 ;
        RECT 85.950 478.950 88.050 481.050 ;
        RECT 82.950 466.950 85.050 469.050 ;
        RECT 46.950 452.250 48.750 453.150 ;
        RECT 49.950 452.400 54.450 453.450 ;
        RECT 49.950 451.950 52.050 452.400 ;
        RECT 55.950 451.950 58.050 454.050 ;
        RECT 61.950 451.950 64.050 454.050 ;
        RECT 64.950 451.950 67.050 454.050 ;
        RECT 70.950 451.950 73.050 454.050 ;
        RECT 79.950 453.450 82.050 454.050 ;
        RECT 77.400 452.400 82.050 453.450 ;
        RECT 62.400 451.050 63.450 451.950 ;
        RECT 46.950 448.950 49.050 451.050 ;
        RECT 50.250 449.850 51.750 450.750 ;
        RECT 52.950 448.950 55.050 451.050 ;
        RECT 56.250 449.850 58.050 450.750 ;
        RECT 61.950 448.950 64.050 451.050 ;
        RECT 52.950 446.850 55.050 447.750 ;
        RECT 43.950 433.950 46.050 436.050 ;
        RECT 44.400 418.050 45.450 433.950 ;
        RECT 52.950 424.950 55.050 427.050 ;
        RECT 53.400 421.050 54.450 424.950 ;
        RECT 65.400 421.050 66.450 451.950 ;
        RECT 71.400 436.050 72.450 451.950 ;
        RECT 70.950 433.950 73.050 436.050 ;
        RECT 77.400 424.050 78.450 452.400 ;
        RECT 79.950 451.950 82.050 452.400 ;
        RECT 83.400 451.050 84.450 466.950 ;
        RECT 92.400 460.050 93.450 481.950 ;
        RECT 95.400 475.050 96.450 484.950 ;
        RECT 94.950 472.950 97.050 475.050 ;
        RECT 101.400 460.050 102.450 487.950 ;
        RECT 103.950 485.850 105.750 486.750 ;
        RECT 106.950 484.950 109.050 487.050 ;
        RECT 110.250 485.850 112.050 486.750 ;
        RECT 91.950 457.950 94.050 460.050 ;
        RECT 97.950 459.450 100.050 460.050 ;
        RECT 95.400 458.400 100.050 459.450 ;
        RECT 85.950 451.950 88.050 454.050 ;
        RECT 89.250 452.250 91.050 453.150 ;
        RECT 79.950 449.850 81.750 450.750 ;
        RECT 82.950 448.950 85.050 451.050 ;
        RECT 86.250 449.850 87.750 450.750 ;
        RECT 88.950 448.950 91.050 451.050 ;
        RECT 82.950 446.850 85.050 447.750 ;
        RECT 79.950 439.950 82.050 442.050 ;
        RECT 76.950 421.950 79.050 424.050 ;
        RECT 80.400 421.050 81.450 439.950 ;
        RECT 89.400 421.050 90.450 448.950 ;
        RECT 95.400 442.050 96.450 458.400 ;
        RECT 97.950 457.950 100.050 458.400 ;
        RECT 100.950 457.950 103.050 460.050 ;
        RECT 107.400 457.050 108.450 484.950 ;
        RECT 113.400 484.050 114.450 488.400 ;
        RECT 115.950 488.250 118.050 489.150 ;
        RECT 121.950 487.950 124.050 490.050 ;
        RECT 127.950 487.950 130.050 490.050 ;
        RECT 133.950 487.950 136.050 490.050 ;
        RECT 139.950 488.250 142.050 489.150 ;
        RECT 122.400 487.050 123.450 487.950 ;
        RECT 134.400 487.050 135.450 487.950 ;
        RECT 115.950 484.950 118.050 487.050 ;
        RECT 119.250 485.250 120.750 486.150 ;
        RECT 121.950 484.950 124.050 487.050 ;
        RECT 125.250 485.250 127.050 486.150 ;
        RECT 127.950 484.950 130.050 487.050 ;
        RECT 130.950 485.250 132.750 486.150 ;
        RECT 133.950 484.950 136.050 487.050 ;
        RECT 137.250 485.250 138.750 486.150 ;
        RECT 139.950 484.950 142.050 487.050 ;
        RECT 112.950 481.950 115.050 484.050 ;
        RECT 113.400 478.050 114.450 481.950 ;
        RECT 116.400 481.050 117.450 484.950 ;
        RECT 118.950 481.950 121.050 484.050 ;
        RECT 122.250 482.850 123.750 483.750 ;
        RECT 124.950 481.950 127.050 484.050 ;
        RECT 115.950 478.950 118.050 481.050 ;
        RECT 125.400 478.050 126.450 481.950 ;
        RECT 112.950 475.950 115.050 478.050 ;
        RECT 124.950 475.950 127.050 478.050 ;
        RECT 128.400 472.050 129.450 484.950 ;
        RECT 130.950 481.950 133.050 484.050 ;
        RECT 134.250 482.850 135.750 483.750 ;
        RECT 136.950 481.950 139.050 484.050 ;
        RECT 131.400 481.050 132.450 481.950 ;
        RECT 130.950 478.950 133.050 481.050 ;
        RECT 127.950 469.950 130.050 472.050 ;
        RECT 131.400 463.050 132.450 478.950 ;
        RECT 140.400 478.050 141.450 484.950 ;
        RECT 143.400 481.050 144.450 499.950 ;
        RECT 154.950 490.950 157.050 493.050 ;
        RECT 148.950 488.250 151.050 489.150 ;
        RECT 155.400 487.050 156.450 490.950 ;
        RECT 148.950 484.950 151.050 487.050 ;
        RECT 152.250 485.250 153.750 486.150 ;
        RECT 154.950 484.950 157.050 487.050 ;
        RECT 158.250 485.250 160.050 486.150 ;
        RECT 149.400 481.050 150.450 484.950 ;
        RECT 151.950 481.950 154.050 484.050 ;
        RECT 155.250 482.850 156.750 483.750 ;
        RECT 157.950 481.950 160.050 484.050 ;
        RECT 142.950 478.950 145.050 481.050 ;
        RECT 148.950 478.950 151.050 481.050 ;
        RECT 139.950 475.950 142.050 478.050 ;
        RECT 149.400 475.050 150.450 478.950 ;
        RECT 148.950 472.950 151.050 475.050 ;
        RECT 136.950 469.950 139.050 472.050 ;
        RECT 142.950 469.950 145.050 472.050 ;
        RECT 130.950 460.950 133.050 463.050 ;
        RECT 137.400 460.050 138.450 469.950 ;
        RECT 118.950 457.950 121.050 460.050 ;
        RECT 136.950 457.950 139.050 460.050 ;
        RECT 97.950 455.850 100.050 456.750 ;
        RECT 100.950 455.250 103.050 456.150 ;
        RECT 106.950 454.950 109.050 457.050 ;
        RECT 100.950 451.950 103.050 454.050 ;
        RECT 94.950 439.950 97.050 442.050 ;
        RECT 101.400 421.050 102.450 451.950 ;
        RECT 107.400 450.450 108.450 454.950 ;
        RECT 119.400 454.050 120.450 457.950 ;
        RECT 121.950 454.950 124.050 457.050 ;
        RECT 136.950 455.850 139.050 456.750 ;
        RECT 143.400 456.450 144.450 469.950 ;
        RECT 152.400 469.050 153.450 481.950 ;
        RECT 151.950 466.950 154.050 469.050 ;
        RECT 161.400 468.450 162.450 505.950 ;
        RECT 167.400 493.050 168.450 523.950 ;
        RECT 176.400 499.050 177.450 547.950 ;
        RECT 182.400 529.050 183.450 562.950 ;
        RECT 185.400 553.050 186.450 577.950 ;
        RECT 188.400 562.050 189.450 580.950 ;
        RECT 191.400 577.050 192.450 580.950 ;
        RECT 190.950 574.950 193.050 577.050 ;
        RECT 194.400 573.450 195.450 622.950 ;
        RECT 200.400 613.050 201.450 625.950 ;
        RECT 203.400 622.050 204.450 625.950 ;
        RECT 202.950 619.950 205.050 622.050 ;
        RECT 209.400 619.050 210.450 625.950 ;
        RECT 215.400 619.050 216.450 625.950 ;
        RECT 208.950 616.950 211.050 619.050 ;
        RECT 211.950 616.950 214.050 619.050 ;
        RECT 214.950 616.950 217.050 619.050 ;
        RECT 196.950 610.950 199.050 613.050 ;
        RECT 199.950 610.950 202.050 613.050 ;
        RECT 197.400 595.050 198.450 610.950 ;
        RECT 208.950 607.950 211.050 610.050 ;
        RECT 209.400 601.050 210.450 607.950 ;
        RECT 212.400 601.050 213.450 616.950 ;
        RECT 218.400 604.050 219.450 631.950 ;
        RECT 220.950 629.250 223.050 630.150 ;
        RECT 223.950 629.850 226.050 630.750 ;
        RECT 229.950 629.250 232.050 630.150 ;
        RECT 220.950 625.950 223.050 628.050 ;
        RECT 229.950 625.950 232.050 628.050 ;
        RECT 221.400 625.050 222.450 625.950 ;
        RECT 230.400 625.050 231.450 625.950 ;
        RECT 220.950 622.950 223.050 625.050 ;
        RECT 229.950 622.950 232.050 625.050 ;
        RECT 233.400 622.050 234.450 661.950 ;
        RECT 242.400 646.050 243.450 677.400 ;
        RECT 244.950 673.950 247.050 676.050 ;
        RECT 253.950 673.950 256.050 676.050 ;
        RECT 245.400 661.050 246.450 673.950 ;
        RECT 254.400 670.050 255.450 673.950 ;
        RECT 257.400 670.050 258.450 694.950 ;
        RECT 272.400 685.050 273.450 694.950 ;
        RECT 290.400 685.050 291.450 697.950 ;
        RECT 292.950 694.950 295.050 697.050 ;
        RECT 296.400 694.050 297.450 697.950 ;
        RECT 299.400 694.050 300.450 706.950 ;
        RECT 308.400 703.050 309.450 706.950 ;
        RECT 325.950 704.250 328.050 705.150 ;
        RECT 304.950 701.250 306.750 702.150 ;
        RECT 307.950 700.950 310.050 703.050 ;
        RECT 313.950 700.950 316.050 703.050 ;
        RECT 316.950 701.250 318.750 702.150 ;
        RECT 319.950 700.950 322.050 703.050 ;
        RECT 323.250 701.250 324.750 702.150 ;
        RECT 325.950 700.950 328.050 703.050 ;
        RECT 304.950 699.450 307.050 700.050 ;
        RECT 302.400 698.400 307.050 699.450 ;
        RECT 308.250 698.850 310.050 699.750 ;
        RECT 295.950 691.950 298.050 694.050 ;
        RECT 298.950 691.950 301.050 694.050 ;
        RECT 271.950 682.950 274.050 685.050 ;
        RECT 289.950 682.950 292.050 685.050 ;
        RECT 302.400 684.450 303.450 698.400 ;
        RECT 304.950 697.950 307.050 698.400 ;
        RECT 310.950 698.250 313.050 699.150 ;
        RECT 313.950 698.850 316.050 699.750 ;
        RECT 316.950 697.950 319.050 700.050 ;
        RECT 320.250 698.850 321.750 699.750 ;
        RECT 322.950 697.950 325.050 700.050 ;
        RECT 304.950 694.950 307.050 697.050 ;
        RECT 310.950 694.950 313.050 697.050 ;
        RECT 317.400 696.450 318.450 697.950 ;
        RECT 317.400 695.400 321.450 696.450 ;
        RECT 299.400 683.400 303.450 684.450 ;
        RECT 299.400 682.050 300.450 683.400 ;
        RECT 298.950 679.950 301.050 682.050 ;
        RECT 301.950 679.950 304.050 682.050 ;
        RECT 274.950 676.950 277.050 679.050 ;
        RECT 262.950 673.950 265.050 676.050 ;
        RECT 250.950 668.250 252.750 669.150 ;
        RECT 253.950 667.950 256.050 670.050 ;
        RECT 256.950 667.950 259.050 670.050 ;
        RECT 259.950 667.950 262.050 670.050 ;
        RECT 250.950 664.950 253.050 667.050 ;
        RECT 254.250 665.850 255.750 666.750 ;
        RECT 256.950 664.950 259.050 667.050 ;
        RECT 260.250 665.850 262.050 666.750 ;
        RECT 251.400 661.050 252.450 664.950 ;
        RECT 256.950 662.850 259.050 663.750 ;
        RECT 263.400 661.050 264.450 673.950 ;
        RECT 265.950 668.250 267.750 669.150 ;
        RECT 268.950 667.950 271.050 670.050 ;
        RECT 272.250 668.250 274.050 669.150 ;
        RECT 269.250 665.850 270.750 666.750 ;
        RECT 271.950 664.950 274.050 667.050 ;
        RECT 272.400 664.050 273.450 664.950 ;
        RECT 271.950 661.950 274.050 664.050 ;
        RECT 244.950 658.950 247.050 661.050 ;
        RECT 250.950 658.950 253.050 661.050 ;
        RECT 262.950 658.950 265.050 661.050 ;
        RECT 275.400 658.050 276.450 676.950 ;
        RECT 302.400 673.050 303.450 679.950 ;
        RECT 283.950 670.950 286.050 673.050 ;
        RECT 287.250 671.250 288.750 672.150 ;
        RECT 289.950 670.950 292.050 673.050 ;
        RECT 301.950 670.950 304.050 673.050 ;
        RECT 280.950 667.950 283.050 670.050 ;
        RECT 284.250 668.850 285.750 669.750 ;
        RECT 286.950 667.950 289.050 670.050 ;
        RECT 290.250 668.850 292.050 669.750 ;
        RECT 292.950 668.250 294.750 669.150 ;
        RECT 295.950 667.950 298.050 670.050 ;
        RECT 299.250 668.250 301.050 669.150 ;
        RECT 280.950 665.850 283.050 666.750 ;
        RECT 292.950 664.950 295.050 667.050 ;
        RECT 296.250 665.850 297.750 666.750 ;
        RECT 298.950 664.950 301.050 667.050 ;
        RECT 286.950 661.950 289.050 664.050 ;
        RECT 274.950 655.950 277.050 658.050 ;
        RECT 262.950 652.950 265.050 655.050 ;
        RECT 268.950 652.950 271.050 655.050 ;
        RECT 235.950 643.950 238.050 646.050 ;
        RECT 241.950 643.950 244.050 646.050 ;
        RECT 236.400 634.050 237.450 643.950 ;
        RECT 253.950 634.950 256.050 637.050 ;
        RECT 235.950 631.950 238.050 634.050 ;
        RECT 239.250 632.250 240.750 633.150 ;
        RECT 247.950 632.250 250.050 633.150 ;
        RECT 254.400 631.050 255.450 634.950 ;
        RECT 263.400 631.050 264.450 652.950 ;
        RECT 269.400 640.050 270.450 652.950 ;
        RECT 268.950 637.950 271.050 640.050 ;
        RECT 269.400 631.050 270.450 637.950 ;
        RECT 274.950 634.950 277.050 637.050 ;
        RECT 235.950 629.850 237.750 630.750 ;
        RECT 238.950 628.950 241.050 631.050 ;
        RECT 242.250 629.850 244.050 630.750 ;
        RECT 247.950 628.950 250.050 631.050 ;
        RECT 251.250 629.250 252.750 630.150 ;
        RECT 253.950 628.950 256.050 631.050 ;
        RECT 257.250 629.250 259.050 630.150 ;
        RECT 259.950 629.250 261.750 630.150 ;
        RECT 262.950 628.950 265.050 631.050 ;
        RECT 266.250 629.250 267.750 630.150 ;
        RECT 268.950 628.950 271.050 631.050 ;
        RECT 272.250 629.250 274.050 630.150 ;
        RECT 235.950 625.950 238.050 628.050 ;
        RECT 241.950 625.950 244.050 628.050 ;
        RECT 250.950 625.950 253.050 628.050 ;
        RECT 254.250 626.850 255.750 627.750 ;
        RECT 256.950 625.950 259.050 628.050 ;
        RECT 259.950 625.950 262.050 628.050 ;
        RECT 263.250 626.850 264.750 627.750 ;
        RECT 265.950 625.950 268.050 628.050 ;
        RECT 269.250 626.850 270.750 627.750 ;
        RECT 271.950 625.950 274.050 628.050 ;
        RECT 232.950 619.950 235.050 622.050 ;
        RECT 217.950 601.950 220.050 604.050 ;
        RECT 236.400 601.050 237.450 625.950 ;
        RECT 238.950 616.950 241.050 619.050 ;
        RECT 202.950 598.950 205.050 601.050 ;
        RECT 206.250 599.250 207.750 600.150 ;
        RECT 208.950 598.950 211.050 601.050 ;
        RECT 211.950 598.950 214.050 601.050 ;
        RECT 215.250 599.250 216.750 600.150 ;
        RECT 217.950 598.950 220.050 601.050 ;
        RECT 221.250 599.250 222.750 600.150 ;
        RECT 223.950 598.950 226.050 601.050 ;
        RECT 232.950 598.950 235.050 601.050 ;
        RECT 235.950 598.950 238.050 601.050 ;
        RECT 233.400 598.050 234.450 598.950 ;
        RECT 199.950 595.950 202.050 598.050 ;
        RECT 203.250 596.850 204.750 597.750 ;
        RECT 205.950 595.950 208.050 598.050 ;
        RECT 209.250 596.850 211.050 597.750 ;
        RECT 211.950 596.850 213.750 597.750 ;
        RECT 214.950 595.950 217.050 598.050 ;
        RECT 218.250 596.850 219.750 597.750 ;
        RECT 220.950 595.950 223.050 598.050 ;
        RECT 224.250 596.850 226.050 597.750 ;
        RECT 229.950 596.250 231.750 597.150 ;
        RECT 232.950 595.950 235.050 598.050 ;
        RECT 236.250 596.250 238.050 597.150 ;
        RECT 196.950 592.950 199.050 595.050 ;
        RECT 199.950 593.850 202.050 594.750 ;
        RECT 208.950 592.950 211.050 595.050 ;
        RECT 191.400 572.400 195.450 573.450 ;
        RECT 191.400 565.050 192.450 572.400 ;
        RECT 193.950 568.950 196.050 571.050 ;
        RECT 190.950 562.950 193.050 565.050 ;
        RECT 194.400 562.050 195.450 568.950 ;
        RECT 196.950 565.950 199.050 568.050 ;
        RECT 187.950 559.950 190.050 562.050 ;
        RECT 191.250 560.250 192.750 561.150 ;
        RECT 193.950 559.950 196.050 562.050 ;
        RECT 187.950 557.850 189.750 558.750 ;
        RECT 190.950 556.950 193.050 559.050 ;
        RECT 194.250 557.850 196.050 558.750 ;
        RECT 197.400 556.050 198.450 565.950 ;
        RECT 199.950 557.250 202.050 558.150 ;
        RECT 205.950 557.250 208.050 558.150 ;
        RECT 190.950 553.950 193.050 556.050 ;
        RECT 193.950 553.950 196.050 556.050 ;
        RECT 196.950 553.950 199.050 556.050 ;
        RECT 199.950 553.950 202.050 556.050 ;
        RECT 203.250 554.250 204.750 555.150 ;
        RECT 184.950 550.950 187.050 553.050 ;
        RECT 181.950 528.450 184.050 529.050 ;
        RECT 179.400 527.400 184.050 528.450 ;
        RECT 179.400 520.050 180.450 527.400 ;
        RECT 181.950 526.950 184.050 527.400 ;
        RECT 185.250 527.250 186.750 528.150 ;
        RECT 187.950 526.950 190.050 529.050 ;
        RECT 191.400 526.050 192.450 553.950 ;
        RECT 181.950 524.850 183.750 525.750 ;
        RECT 184.950 523.950 187.050 526.050 ;
        RECT 188.250 524.850 189.750 525.750 ;
        RECT 190.950 523.950 193.050 526.050 ;
        RECT 178.950 517.950 181.050 520.050 ;
        RECT 185.400 508.050 186.450 523.950 ;
        RECT 190.950 521.850 193.050 522.750 ;
        RECT 184.950 505.950 187.050 508.050 ;
        RECT 175.950 496.950 178.050 499.050 ;
        RECT 194.400 493.050 195.450 553.950 ;
        RECT 200.400 553.050 201.450 553.950 ;
        RECT 199.950 550.950 202.050 553.050 ;
        RECT 202.950 550.950 205.050 553.050 ;
        RECT 203.400 535.050 204.450 550.950 ;
        RECT 209.400 550.050 210.450 592.950 ;
        RECT 215.400 592.050 216.450 595.950 ;
        RECT 214.950 589.950 217.050 592.050 ;
        RECT 221.400 570.450 222.450 595.950 ;
        RECT 229.950 592.950 232.050 595.050 ;
        RECT 233.250 593.850 234.750 594.750 ;
        RECT 235.950 592.950 238.050 595.050 ;
        RECT 221.400 569.400 225.450 570.450 ;
        RECT 214.950 559.950 217.050 562.050 ;
        RECT 218.250 560.250 219.750 561.150 ;
        RECT 214.950 557.850 216.750 558.750 ;
        RECT 217.950 556.950 220.050 559.050 ;
        RECT 221.250 557.850 223.050 558.750 ;
        RECT 224.400 555.450 225.450 569.400 ;
        RECT 230.400 562.050 231.450 592.950 ;
        RECT 236.400 589.050 237.450 592.950 ;
        RECT 235.950 586.950 238.050 589.050 ;
        RECT 232.950 574.950 235.050 577.050 ;
        RECT 226.950 560.250 229.050 561.150 ;
        RECT 229.950 559.950 232.050 562.050 ;
        RECT 233.400 559.050 234.450 574.950 ;
        RECT 239.400 562.050 240.450 616.950 ;
        RECT 242.400 616.050 243.450 625.950 ;
        RECT 251.400 622.050 252.450 625.950 ;
        RECT 253.950 622.950 256.050 625.050 ;
        RECT 250.950 619.950 253.050 622.050 ;
        RECT 241.950 613.950 244.050 616.050 ;
        RECT 244.950 613.950 247.050 616.050 ;
        RECT 245.400 601.050 246.450 613.950 ;
        RECT 254.400 610.050 255.450 622.950 ;
        RECT 257.400 622.050 258.450 625.950 ;
        RECT 256.950 619.950 259.050 622.050 ;
        RECT 260.400 619.050 261.450 625.950 ;
        RECT 262.950 622.950 265.050 625.050 ;
        RECT 259.950 616.950 262.050 619.050 ;
        RECT 250.950 607.950 253.050 610.050 ;
        RECT 253.950 607.950 256.050 610.050 ;
        RECT 251.400 601.050 252.450 607.950 ;
        RECT 259.950 604.950 262.050 607.050 ;
        RECT 256.950 601.950 259.050 604.050 ;
        RECT 244.950 600.450 247.050 601.050 ;
        RECT 242.400 599.400 247.050 600.450 ;
        RECT 242.400 595.050 243.450 599.400 ;
        RECT 244.950 598.950 247.050 599.400 ;
        RECT 248.250 599.250 249.750 600.150 ;
        RECT 250.950 598.950 253.050 601.050 ;
        RECT 244.950 596.850 246.750 597.750 ;
        RECT 247.950 595.950 250.050 598.050 ;
        RECT 251.250 596.850 252.750 597.750 ;
        RECT 253.950 597.450 256.050 598.050 ;
        RECT 257.400 597.450 258.450 601.950 ;
        RECT 253.950 596.400 258.450 597.450 ;
        RECT 253.950 595.950 256.050 596.400 ;
        RECT 241.950 592.950 244.050 595.050 ;
        RECT 244.950 592.950 247.050 595.050 ;
        RECT 242.400 582.450 243.450 592.950 ;
        RECT 245.400 585.450 246.450 592.950 ;
        RECT 248.400 589.050 249.450 595.950 ;
        RECT 253.950 593.850 256.050 594.750 ;
        RECT 247.950 586.950 250.050 589.050 ;
        RECT 257.400 586.050 258.450 596.400 ;
        RECT 245.400 584.400 249.450 585.450 ;
        RECT 242.400 581.400 246.450 582.450 ;
        RECT 241.950 565.950 244.050 568.050 ;
        RECT 238.950 559.950 241.050 562.050 ;
        RECT 242.400 559.050 243.450 565.950 ;
        RECT 245.400 562.050 246.450 581.400 ;
        RECT 244.950 559.950 247.050 562.050 ;
        RECT 248.400 559.050 249.450 584.400 ;
        RECT 256.950 583.950 259.050 586.050 ;
        RECT 260.400 583.050 261.450 604.950 ;
        RECT 263.400 595.050 264.450 622.950 ;
        RECT 266.400 622.050 267.450 625.950 ;
        RECT 265.950 619.950 268.050 622.050 ;
        RECT 265.950 598.950 268.050 601.050 ;
        RECT 265.950 596.850 268.050 597.750 ;
        RECT 268.950 596.250 271.050 597.150 ;
        RECT 272.400 595.050 273.450 625.950 ;
        RECT 275.400 622.050 276.450 634.950 ;
        RECT 281.250 632.250 282.750 633.150 ;
        RECT 287.400 631.050 288.450 661.950 ;
        RECT 293.400 658.050 294.450 664.950 ;
        RECT 292.950 655.950 295.050 658.050 ;
        RECT 289.950 634.950 292.050 637.050 ;
        RECT 277.950 629.850 279.750 630.750 ;
        RECT 280.950 628.950 283.050 631.050 ;
        RECT 284.250 629.850 286.050 630.750 ;
        RECT 286.950 628.950 289.050 631.050 ;
        RECT 274.950 619.950 277.050 622.050 ;
        RECT 274.950 607.950 277.050 610.050 ;
        RECT 275.400 601.050 276.450 607.950 ;
        RECT 274.950 598.950 277.050 601.050 ;
        RECT 281.400 600.450 282.450 628.950 ;
        RECT 286.950 625.950 289.050 628.050 ;
        RECT 290.400 627.450 291.450 634.950 ;
        RECT 292.950 629.250 294.750 630.150 ;
        RECT 299.400 628.050 300.450 664.950 ;
        RECT 305.400 655.050 306.450 694.950 ;
        RECT 311.400 685.050 312.450 694.950 ;
        RECT 310.950 682.950 313.050 685.050 ;
        RECT 316.950 676.950 319.050 679.050 ;
        RECT 310.950 670.950 313.050 673.050 ;
        RECT 311.400 670.050 312.450 670.950 ;
        RECT 317.400 670.050 318.450 676.950 ;
        RECT 320.400 676.050 321.450 695.400 ;
        RECT 326.400 694.050 327.450 700.950 ;
        RECT 329.400 700.050 330.450 706.950 ;
        RECT 334.950 703.950 337.050 706.050 ;
        RECT 352.950 705.450 355.050 706.050 ;
        RECT 350.250 704.250 351.750 705.150 ;
        RECT 352.950 704.400 357.450 705.450 ;
        RECT 352.950 703.950 355.050 704.400 ;
        RECT 335.400 700.050 336.450 703.950 ;
        RECT 337.950 700.950 340.050 703.050 ;
        RECT 346.950 701.850 348.750 702.750 ;
        RECT 349.950 700.950 352.050 703.050 ;
        RECT 353.250 701.850 355.050 702.750 ;
        RECT 350.400 700.050 351.450 700.950 ;
        RECT 328.950 697.950 331.050 700.050 ;
        RECT 334.950 697.950 337.050 700.050 ;
        RECT 337.950 698.850 340.050 699.750 ;
        RECT 343.950 698.850 346.050 699.750 ;
        RECT 349.950 697.950 352.050 700.050 ;
        RECT 325.950 691.950 328.050 694.050 ;
        RECT 319.950 673.950 322.050 676.050 ;
        RECT 307.950 668.250 309.750 669.150 ;
        RECT 310.950 667.950 313.050 670.050 ;
        RECT 316.950 667.950 319.050 670.050 ;
        RECT 320.400 667.050 321.450 673.950 ;
        RECT 335.400 673.050 336.450 697.950 ;
        RECT 356.400 697.050 357.450 704.400 ;
        RECT 349.950 694.950 352.050 697.050 ;
        RECT 355.950 694.950 358.050 697.050 ;
        RECT 340.950 679.950 343.050 682.050 ;
        RECT 341.400 673.050 342.450 679.950 ;
        RECT 346.950 673.950 349.050 676.050 ;
        RECT 347.400 673.050 348.450 673.950 ;
        RECT 331.950 670.950 334.050 673.050 ;
        RECT 334.950 670.950 337.050 673.050 ;
        RECT 338.250 671.250 339.750 672.150 ;
        RECT 340.950 670.950 343.050 673.050 ;
        RECT 344.250 671.250 345.750 672.150 ;
        RECT 346.950 670.950 349.050 673.050 ;
        RECT 322.950 668.250 324.750 669.150 ;
        RECT 325.950 667.950 328.050 670.050 ;
        RECT 329.250 668.250 331.050 669.150 ;
        RECT 332.400 667.050 333.450 670.950 ;
        RECT 334.950 668.850 336.750 669.750 ;
        RECT 337.950 667.950 340.050 670.050 ;
        RECT 341.250 668.850 342.750 669.750 ;
        RECT 343.950 667.950 346.050 670.050 ;
        RECT 347.250 668.850 349.050 669.750 ;
        RECT 307.950 664.950 310.050 667.050 ;
        RECT 311.250 665.850 312.750 666.750 ;
        RECT 313.950 664.950 316.050 667.050 ;
        RECT 317.250 665.850 319.050 666.750 ;
        RECT 319.950 664.950 322.050 667.050 ;
        RECT 322.950 664.950 325.050 667.050 ;
        RECT 326.250 665.850 327.750 666.750 ;
        RECT 328.950 664.950 331.050 667.050 ;
        RECT 331.950 664.950 334.050 667.050 ;
        RECT 343.950 664.950 346.050 667.050 ;
        RECT 346.950 664.950 349.050 667.050 ;
        RECT 308.400 661.050 309.450 664.950 ;
        RECT 313.950 662.850 316.050 663.750 ;
        RECT 323.400 663.450 324.450 664.950 ;
        RECT 323.400 662.400 327.450 663.450 ;
        RECT 307.950 658.950 310.050 661.050 ;
        RECT 304.950 652.950 307.050 655.050 ;
        RECT 322.950 646.950 325.050 649.050 ;
        RECT 301.950 632.250 304.050 633.150 ;
        RECT 301.950 628.950 304.050 631.050 ;
        RECT 305.250 629.250 306.750 630.150 ;
        RECT 307.950 628.950 310.050 631.050 ;
        RECT 311.250 629.250 313.050 630.150 ;
        RECT 316.950 628.950 319.050 631.050 ;
        RECT 292.950 627.450 295.050 628.050 ;
        RECT 290.400 626.400 295.050 627.450 ;
        RECT 296.250 626.850 298.050 627.750 ;
        RECT 292.950 625.950 295.050 626.400 ;
        RECT 298.950 625.950 301.050 628.050 ;
        RECT 287.400 607.050 288.450 625.950 ;
        RECT 289.950 622.950 292.050 625.050 ;
        RECT 286.950 604.950 289.050 607.050 ;
        RECT 278.400 599.400 282.450 600.450 ;
        RECT 274.950 596.850 277.050 597.750 ;
        RECT 262.950 592.950 265.050 595.050 ;
        RECT 268.950 592.950 271.050 595.050 ;
        RECT 271.950 592.950 274.050 595.050 ;
        RECT 263.400 592.050 264.450 592.950 ;
        RECT 262.950 589.950 265.050 592.050 ;
        RECT 256.950 580.950 259.050 583.050 ;
        RECT 259.950 580.950 262.050 583.050 ;
        RECT 253.950 574.950 256.050 577.050 ;
        RECT 226.950 556.950 229.050 559.050 ;
        RECT 230.250 557.250 231.750 558.150 ;
        RECT 232.950 556.950 235.050 559.050 ;
        RECT 236.250 557.250 238.050 558.150 ;
        RECT 238.950 557.250 240.750 558.150 ;
        RECT 241.950 556.950 244.050 559.050 ;
        RECT 245.250 557.250 246.750 558.150 ;
        RECT 247.950 556.950 250.050 559.050 ;
        RECT 251.250 557.250 253.050 558.150 ;
        RECT 221.400 554.400 225.450 555.450 ;
        RECT 208.950 547.950 211.050 550.050 ;
        RECT 211.950 538.950 214.050 541.050 ;
        RECT 205.950 535.950 208.050 538.050 ;
        RECT 202.950 532.950 205.050 535.050 ;
        RECT 199.950 529.950 202.050 532.050 ;
        RECT 202.950 529.950 205.050 532.050 ;
        RECT 200.400 529.050 201.450 529.950 ;
        RECT 206.400 529.050 207.450 535.950 ;
        RECT 208.950 532.950 211.050 535.050 ;
        RECT 199.950 526.950 202.050 529.050 ;
        RECT 203.250 527.850 204.750 528.750 ;
        RECT 205.950 526.950 208.050 529.050 ;
        RECT 199.950 524.850 202.050 525.750 ;
        RECT 205.950 524.850 208.050 525.750 ;
        RECT 199.950 499.950 202.050 502.050 ;
        RECT 166.950 490.950 169.050 493.050 ;
        RECT 184.950 490.950 187.050 493.050 ;
        RECT 193.950 490.950 196.050 493.050 ;
        RECT 167.400 489.450 168.450 490.950 ;
        RECT 163.950 488.250 166.050 489.150 ;
        RECT 167.400 488.400 171.450 489.450 ;
        RECT 170.400 487.050 171.450 488.400 ;
        RECT 163.950 484.950 166.050 487.050 ;
        RECT 167.250 485.250 168.750 486.150 ;
        RECT 169.950 484.950 172.050 487.050 ;
        RECT 178.950 486.450 181.050 487.050 ;
        RECT 173.250 485.250 175.050 486.150 ;
        RECT 178.950 485.400 183.450 486.450 ;
        RECT 178.950 484.950 181.050 485.400 ;
        RECT 164.400 484.050 165.450 484.950 ;
        RECT 163.950 481.950 166.050 484.050 ;
        RECT 166.950 481.950 169.050 484.050 ;
        RECT 170.250 482.850 171.750 483.750 ;
        RECT 172.950 481.950 175.050 484.050 ;
        RECT 175.950 482.250 178.050 483.150 ;
        RECT 178.950 482.850 181.050 483.750 ;
        RECT 167.400 481.050 168.450 481.950 ;
        RECT 166.950 478.950 169.050 481.050 ;
        RECT 158.400 467.400 162.450 468.450 ;
        RECT 145.950 456.450 148.050 457.050 ;
        RECT 139.950 455.250 142.050 456.150 ;
        RECT 143.400 455.400 148.050 456.450 ;
        RECT 145.950 454.950 148.050 455.400 ;
        RECT 149.250 455.250 150.750 456.150 ;
        RECT 151.950 454.950 154.050 457.050 ;
        RECT 109.950 452.250 111.750 453.150 ;
        RECT 112.950 451.950 115.050 454.050 ;
        RECT 116.250 452.250 118.050 453.150 ;
        RECT 118.950 451.950 121.050 454.050 ;
        RECT 122.400 451.050 123.450 454.950 ;
        RECT 124.950 451.950 127.050 454.050 ;
        RECT 128.250 452.250 130.050 453.150 ;
        RECT 139.950 451.950 142.050 454.050 ;
        RECT 142.950 451.950 145.050 454.050 ;
        RECT 145.950 452.850 147.750 453.750 ;
        RECT 148.950 451.950 151.050 454.050 ;
        RECT 152.250 452.850 153.750 453.750 ;
        RECT 109.950 450.450 112.050 451.050 ;
        RECT 107.400 449.400 112.050 450.450 ;
        RECT 113.250 449.850 114.750 450.750 ;
        RECT 109.950 448.950 112.050 449.400 ;
        RECT 115.950 448.950 118.050 451.050 ;
        RECT 118.950 449.850 120.750 450.750 ;
        RECT 121.950 448.950 124.050 451.050 ;
        RECT 125.250 449.850 126.750 450.750 ;
        RECT 127.950 448.950 130.050 451.050 ;
        RECT 121.950 446.850 124.050 447.750 ;
        RECT 52.950 418.950 55.050 421.050 ;
        RECT 64.950 418.950 67.050 421.050 ;
        RECT 67.950 419.250 70.050 420.150 ;
        RECT 76.950 419.250 79.050 420.150 ;
        RECT 79.950 418.950 82.050 421.050 ;
        RECT 88.950 418.950 91.050 421.050 ;
        RECT 97.950 418.950 100.050 421.050 ;
        RECT 100.950 418.950 103.050 421.050 ;
        RECT 103.950 419.250 106.050 420.150 ;
        RECT 133.950 418.950 136.050 421.050 ;
        RECT 98.400 418.050 99.450 418.950 ;
        RECT 43.950 415.950 46.050 418.050 ;
        RECT 49.950 417.450 52.050 418.050 ;
        RECT 47.400 416.400 52.050 417.450 ;
        RECT 35.250 413.250 36.750 414.150 ;
        RECT 37.950 413.400 42.450 414.450 ;
        RECT 37.950 412.950 40.050 413.400 ;
        RECT 44.400 412.050 45.450 415.950 ;
        RECT 28.950 409.950 31.050 412.050 ;
        RECT 32.250 410.850 33.750 411.750 ;
        RECT 34.950 409.950 37.050 412.050 ;
        RECT 43.950 409.950 46.050 412.050 ;
        RECT 35.400 409.050 36.450 409.950 ;
        RECT 47.400 409.050 48.450 416.400 ;
        RECT 49.950 415.950 52.050 416.400 ;
        RECT 53.250 416.250 54.750 417.150 ;
        RECT 55.950 415.950 58.050 418.050 ;
        RECT 58.950 415.950 61.050 418.050 ;
        RECT 61.950 415.950 64.050 418.050 ;
        RECT 65.250 416.250 66.750 417.150 ;
        RECT 67.950 415.950 70.050 418.050 ;
        RECT 71.250 416.250 73.050 417.150 ;
        RECT 73.950 416.250 75.750 417.150 ;
        RECT 76.950 415.950 79.050 418.050 ;
        RECT 82.950 417.450 85.050 418.050 ;
        RECT 91.950 417.450 94.050 418.050 ;
        RECT 80.250 416.250 81.750 417.150 ;
        RECT 82.950 416.400 87.450 417.450 ;
        RECT 82.950 415.950 85.050 416.400 ;
        RECT 49.950 413.850 51.750 414.750 ;
        RECT 52.950 412.950 55.050 415.050 ;
        RECT 56.250 413.850 58.050 414.750 ;
        RECT 34.950 406.950 37.050 409.050 ;
        RECT 46.950 406.950 49.050 409.050 ;
        RECT 59.400 408.450 60.450 415.950 ;
        RECT 61.950 413.850 63.750 414.750 ;
        RECT 64.950 412.950 67.050 415.050 ;
        RECT 68.400 412.050 69.450 415.950 ;
        RECT 70.950 412.950 73.050 415.050 ;
        RECT 73.950 412.950 76.050 415.050 ;
        RECT 79.950 412.950 82.050 415.050 ;
        RECT 83.250 413.850 85.050 414.750 ;
        RECT 67.950 409.950 70.050 412.050 ;
        RECT 74.400 411.450 75.450 412.950 ;
        RECT 71.400 410.400 75.450 411.450 ;
        RECT 71.400 408.450 72.450 410.400 ;
        RECT 80.400 409.050 81.450 412.950 ;
        RECT 86.400 409.050 87.450 416.400 ;
        RECT 89.400 416.400 94.050 417.450 ;
        RECT 59.400 407.400 72.450 408.450 ;
        RECT 79.950 406.950 82.050 409.050 ;
        RECT 85.950 406.950 88.050 409.050 ;
        RECT 89.400 406.050 90.450 416.400 ;
        RECT 91.950 415.950 94.050 416.400 ;
        RECT 95.250 416.250 96.750 417.150 ;
        RECT 97.950 415.950 100.050 418.050 ;
        RECT 100.950 416.250 102.750 417.150 ;
        RECT 103.950 415.950 106.050 418.050 ;
        RECT 107.250 416.250 108.750 417.150 ;
        RECT 109.950 415.950 112.050 418.050 ;
        RECT 118.950 415.950 121.050 418.050 ;
        RECT 124.950 417.450 127.050 418.050 ;
        RECT 122.250 416.250 123.750 417.150 ;
        RECT 124.950 416.400 129.450 417.450 ;
        RECT 124.950 415.950 127.050 416.400 ;
        RECT 91.950 413.850 93.750 414.750 ;
        RECT 94.950 412.950 97.050 415.050 ;
        RECT 98.250 413.850 100.050 414.750 ;
        RECT 100.950 412.950 103.050 415.050 ;
        RECT 106.950 412.950 109.050 415.050 ;
        RECT 110.250 413.850 112.050 414.750 ;
        RECT 118.950 413.850 120.750 414.750 ;
        RECT 121.950 412.950 124.050 415.050 ;
        RECT 125.250 413.850 127.050 414.750 ;
        RECT 95.400 412.050 96.450 412.950 ;
        RECT 94.950 409.950 97.050 412.050 ;
        RECT 107.400 406.050 108.450 412.950 ;
        RECT 122.400 406.050 123.450 412.950 ;
        RECT 128.400 409.050 129.450 416.400 ;
        RECT 130.950 413.250 133.050 414.150 ;
        RECT 130.950 409.950 133.050 412.050 ;
        RECT 134.400 411.450 135.450 418.950 ;
        RECT 136.950 415.950 139.050 418.050 ;
        RECT 143.400 415.050 144.450 451.950 ;
        RECT 149.400 448.050 150.450 451.950 ;
        RECT 154.950 449.850 157.050 450.750 ;
        RECT 148.950 445.950 151.050 448.050 ;
        RECT 149.400 445.050 150.450 445.950 ;
        RECT 148.950 442.950 151.050 445.050 ;
        RECT 158.400 433.050 159.450 467.400 ;
        RECT 160.950 463.950 163.050 466.050 ;
        RECT 161.400 436.050 162.450 463.950 ;
        RECT 173.400 463.050 174.450 481.950 ;
        RECT 182.400 481.050 183.450 485.400 ;
        RECT 175.950 478.950 178.050 481.050 ;
        RECT 181.950 478.950 184.050 481.050 ;
        RECT 185.400 463.050 186.450 490.950 ;
        RECT 200.400 490.050 201.450 499.950 ;
        RECT 205.950 493.950 208.050 496.050 ;
        RECT 206.400 490.050 207.450 493.950 ;
        RECT 209.400 490.050 210.450 532.950 ;
        RECT 212.400 529.050 213.450 538.950 ;
        RECT 221.400 532.050 222.450 554.400 ;
        RECT 229.950 553.950 232.050 556.050 ;
        RECT 233.250 554.850 234.750 555.750 ;
        RECT 235.950 553.950 238.050 556.050 ;
        RECT 238.950 553.950 241.050 556.050 ;
        RECT 242.250 554.850 243.750 555.750 ;
        RECT 244.950 553.950 247.050 556.050 ;
        RECT 248.250 554.850 249.750 555.750 ;
        RECT 250.950 553.950 253.050 556.050 ;
        RECT 223.950 550.950 226.050 553.050 ;
        RECT 214.950 529.950 217.050 532.050 ;
        RECT 220.950 529.950 223.050 532.050 ;
        RECT 211.950 526.950 214.050 529.050 ;
        RECT 215.250 527.850 216.750 528.750 ;
        RECT 217.950 528.450 220.050 529.050 ;
        RECT 217.950 527.400 222.450 528.450 ;
        RECT 217.950 526.950 220.050 527.400 ;
        RECT 211.950 524.850 214.050 525.750 ;
        RECT 214.950 523.950 217.050 526.050 ;
        RECT 217.950 524.850 220.050 525.750 ;
        RECT 215.400 522.450 216.450 523.950 ;
        RECT 221.400 523.050 222.450 527.400 ;
        RECT 212.400 521.400 216.450 522.450 ;
        RECT 199.950 487.950 202.050 490.050 ;
        RECT 203.250 488.250 204.750 489.150 ;
        RECT 205.950 487.950 208.050 490.050 ;
        RECT 208.950 487.950 211.050 490.050 ;
        RECT 187.950 485.250 189.750 486.150 ;
        RECT 190.950 484.950 193.050 487.050 ;
        RECT 196.950 484.950 199.050 487.050 ;
        RECT 199.950 485.850 201.750 486.750 ;
        RECT 202.950 484.950 205.050 487.050 ;
        RECT 206.250 485.850 208.050 486.750 ;
        RECT 187.950 481.950 190.050 484.050 ;
        RECT 191.250 482.850 193.050 483.750 ;
        RECT 193.950 482.250 196.050 483.150 ;
        RECT 196.950 482.850 199.050 483.750 ;
        RECT 172.950 460.950 175.050 463.050 ;
        RECT 184.950 460.950 187.050 463.050 ;
        RECT 175.950 457.950 178.050 460.050 ;
        RECT 184.950 457.950 187.050 460.050 ;
        RECT 166.950 454.950 169.050 457.050 ;
        RECT 167.400 451.050 168.450 454.950 ;
        RECT 169.950 451.950 172.050 454.050 ;
        RECT 173.250 452.250 175.050 453.150 ;
        RECT 163.950 449.850 165.750 450.750 ;
        RECT 166.950 448.950 169.050 451.050 ;
        RECT 170.250 449.850 171.750 450.750 ;
        RECT 172.950 448.950 175.050 451.050 ;
        RECT 166.950 446.850 169.050 447.750 ;
        RECT 169.950 445.950 172.050 448.050 ;
        RECT 160.950 433.950 163.050 436.050 ;
        RECT 170.400 433.050 171.450 445.950 ;
        RECT 157.950 430.950 160.050 433.050 ;
        RECT 169.950 430.950 172.050 433.050 ;
        RECT 151.950 427.950 154.050 430.050 ;
        RECT 152.400 418.050 153.450 427.950 ;
        RECT 170.400 427.050 171.450 430.950 ;
        RECT 169.950 424.950 172.050 427.050 ;
        RECT 169.950 421.950 172.050 424.050 ;
        RECT 166.950 418.950 169.050 421.050 ;
        RECT 167.400 418.050 168.450 418.950 ;
        RECT 151.950 415.950 154.050 418.050 ;
        RECT 160.950 417.450 163.050 418.050 ;
        RECT 154.950 416.250 157.050 417.150 ;
        RECT 158.400 416.400 163.050 417.450 ;
        RECT 136.950 413.850 139.050 414.750 ;
        RECT 139.950 413.250 142.050 414.150 ;
        RECT 142.950 412.950 145.050 415.050 ;
        RECT 145.950 413.250 147.750 414.150 ;
        RECT 148.950 412.950 151.050 415.050 ;
        RECT 152.250 413.250 153.750 414.150 ;
        RECT 154.950 412.950 157.050 415.050 ;
        RECT 155.400 412.050 156.450 412.950 ;
        RECT 139.950 411.450 142.050 412.050 ;
        RECT 134.400 410.400 142.050 411.450 ;
        RECT 139.950 409.950 142.050 410.400 ;
        RECT 145.950 409.950 148.050 412.050 ;
        RECT 149.250 410.850 150.750 411.750 ;
        RECT 151.950 409.950 154.050 412.050 ;
        RECT 154.950 409.950 157.050 412.050 ;
        RECT 131.400 409.050 132.450 409.950 ;
        RECT 152.400 409.050 153.450 409.950 ;
        RECT 158.400 409.050 159.450 416.400 ;
        RECT 160.950 415.950 163.050 416.400 ;
        RECT 164.250 416.250 165.750 417.150 ;
        RECT 166.950 415.950 169.050 418.050 ;
        RECT 160.950 413.850 162.750 414.750 ;
        RECT 163.950 412.950 166.050 415.050 ;
        RECT 167.250 413.850 169.050 414.750 ;
        RECT 170.400 411.450 171.450 421.950 ;
        RECT 173.400 421.050 174.450 448.950 ;
        RECT 176.400 442.050 177.450 457.950 ;
        RECT 188.400 457.050 189.450 481.950 ;
        RECT 193.950 478.950 196.050 481.050 ;
        RECT 194.400 475.050 195.450 478.950 ;
        RECT 193.950 472.950 196.050 475.050 ;
        RECT 193.950 457.950 196.050 460.050 ;
        RECT 178.950 454.950 181.050 457.050 ;
        RECT 181.950 454.950 184.050 457.050 ;
        RECT 185.250 455.850 186.750 456.750 ;
        RECT 187.950 454.950 190.050 457.050 ;
        RECT 190.950 454.950 193.050 457.050 ;
        RECT 194.250 455.850 195.750 456.750 ;
        RECT 196.950 454.950 199.050 457.050 ;
        RECT 179.400 448.050 180.450 454.950 ;
        RECT 181.950 452.850 184.050 453.750 ;
        RECT 187.950 452.850 190.050 453.750 ;
        RECT 190.950 452.850 193.050 453.750 ;
        RECT 193.950 451.950 196.050 454.050 ;
        RECT 196.950 452.850 199.050 453.750 ;
        RECT 178.950 445.950 181.050 448.050 ;
        RECT 175.950 439.950 178.050 442.050 ;
        RECT 194.400 439.050 195.450 451.950 ;
        RECT 203.400 447.450 204.450 484.950 ;
        RECT 208.950 481.950 211.050 484.050 ;
        RECT 209.400 478.050 210.450 481.950 ;
        RECT 208.950 475.950 211.050 478.050 ;
        RECT 212.400 463.050 213.450 521.400 ;
        RECT 220.950 520.950 223.050 523.050 ;
        RECT 220.950 514.950 223.050 517.050 ;
        RECT 221.400 514.050 222.450 514.950 ;
        RECT 220.950 511.950 223.050 514.050 ;
        RECT 217.950 484.950 220.050 487.050 ;
        RECT 214.950 482.250 217.050 483.150 ;
        RECT 217.950 482.850 220.050 483.750 ;
        RECT 214.950 478.950 217.050 481.050 ;
        RECT 214.950 472.950 217.050 475.050 ;
        RECT 211.950 460.950 214.050 463.050 ;
        RECT 215.400 457.050 216.450 472.950 ;
        RECT 221.400 466.050 222.450 511.950 ;
        RECT 224.400 508.050 225.450 550.950 ;
        RECT 229.950 538.950 232.050 541.050 ;
        RECT 226.950 535.950 229.050 538.050 ;
        RECT 227.400 529.050 228.450 535.950 ;
        RECT 230.400 532.050 231.450 538.950 ;
        RECT 236.400 538.050 237.450 553.950 ;
        RECT 235.950 535.950 238.050 538.050 ;
        RECT 239.400 532.050 240.450 553.950 ;
        RECT 245.400 550.050 246.450 553.950 ;
        RECT 251.400 553.050 252.450 553.950 ;
        RECT 250.950 550.950 253.050 553.050 ;
        RECT 254.400 550.050 255.450 574.950 ;
        RECT 257.400 562.050 258.450 580.950 ;
        RECT 278.400 577.050 279.450 599.400 ;
        RECT 283.950 598.950 286.050 601.050 ;
        RECT 284.400 598.050 285.450 598.950 ;
        RECT 280.950 596.250 282.750 597.150 ;
        RECT 283.950 595.950 286.050 598.050 ;
        RECT 287.400 595.050 288.450 604.950 ;
        RECT 290.400 601.050 291.450 622.950 ;
        RECT 289.950 598.950 292.050 601.050 ;
        RECT 290.400 598.050 291.450 598.950 ;
        RECT 293.400 598.050 294.450 625.950 ;
        RECT 298.950 619.950 301.050 622.050 ;
        RECT 295.950 601.950 298.050 604.050 ;
        RECT 296.400 598.050 297.450 601.950 ;
        RECT 299.400 601.050 300.450 619.950 ;
        RECT 302.400 610.050 303.450 628.950 ;
        RECT 304.950 625.950 307.050 628.050 ;
        RECT 308.250 626.850 309.750 627.750 ;
        RECT 316.950 626.850 319.050 627.750 ;
        RECT 319.950 626.250 322.050 627.150 ;
        RECT 319.950 622.950 322.050 625.050 ;
        RECT 320.400 622.050 321.450 622.950 ;
        RECT 319.950 619.950 322.050 622.050 ;
        RECT 323.400 616.050 324.450 646.950 ;
        RECT 326.400 637.050 327.450 662.400 ;
        RECT 329.400 658.050 330.450 664.950 ;
        RECT 328.950 655.950 331.050 658.050 ;
        RECT 325.950 634.950 328.050 637.050 ;
        RECT 325.950 631.950 328.050 634.050 ;
        RECT 331.950 633.450 334.050 634.050 ;
        RECT 329.250 632.250 330.750 633.150 ;
        RECT 331.950 632.400 336.450 633.450 ;
        RECT 331.950 631.950 334.050 632.400 ;
        RECT 325.950 629.850 327.750 630.750 ;
        RECT 328.950 628.950 331.050 631.050 ;
        RECT 332.250 629.850 334.050 630.750 ;
        RECT 329.400 625.050 330.450 628.950 ;
        RECT 325.950 622.950 328.050 625.050 ;
        RECT 328.950 622.950 331.050 625.050 ;
        RECT 335.400 624.450 336.450 632.400 ;
        RECT 341.250 629.250 343.050 630.150 ;
        RECT 337.950 626.850 339.750 627.750 ;
        RECT 340.950 625.950 343.050 628.050 ;
        RECT 344.400 625.050 345.450 664.950 ;
        RECT 347.400 661.050 348.450 664.950 ;
        RECT 346.950 658.950 349.050 661.050 ;
        RECT 350.400 636.450 351.450 694.950 ;
        RECT 359.400 693.450 360.450 709.950 ;
        RECT 371.400 703.050 372.450 712.950 ;
        RECT 448.950 710.400 451.050 712.500 ;
        RECT 469.950 711.300 472.050 713.400 ;
        RECT 547.950 711.300 550.050 713.400 ;
        RECT 631.950 713.100 634.050 715.200 ;
        RECT 382.950 703.950 385.050 706.050 ;
        RECT 388.950 704.250 391.050 705.150 ;
        RECT 398.250 704.250 399.750 705.150 ;
        RECT 400.950 703.950 403.050 706.050 ;
        RECT 383.400 703.050 384.450 703.950 ;
        RECT 361.950 701.250 363.750 702.150 ;
        RECT 364.950 700.950 367.050 703.050 ;
        RECT 368.250 701.250 369.750 702.150 ;
        RECT 370.950 700.950 373.050 703.050 ;
        RECT 374.250 701.250 376.050 702.150 ;
        RECT 376.950 700.950 379.050 703.050 ;
        RECT 379.950 701.250 381.750 702.150 ;
        RECT 382.950 700.950 385.050 703.050 ;
        RECT 386.250 701.250 387.750 702.150 ;
        RECT 388.950 700.950 391.050 703.050 ;
        RECT 394.950 701.850 396.750 702.750 ;
        RECT 397.950 700.950 400.050 703.050 ;
        RECT 401.250 701.850 403.050 702.750 ;
        RECT 412.950 702.450 415.050 703.050 ;
        RECT 412.950 701.400 417.450 702.450 ;
        RECT 412.950 700.950 415.050 701.400 ;
        RECT 361.950 697.950 364.050 700.050 ;
        RECT 365.250 698.850 366.750 699.750 ;
        RECT 367.950 697.950 370.050 700.050 ;
        RECT 371.250 698.850 372.750 699.750 ;
        RECT 373.950 697.950 376.050 700.050 ;
        RECT 362.400 696.450 363.450 697.950 ;
        RECT 362.400 695.400 369.450 696.450 ;
        RECT 359.400 692.400 363.450 693.450 ;
        RECT 355.950 688.950 358.050 691.050 ;
        RECT 352.950 676.950 355.050 679.050 ;
        RECT 353.400 673.050 354.450 676.950 ;
        RECT 356.400 673.050 357.450 688.950 ;
        RECT 362.400 673.050 363.450 692.400 ;
        RECT 352.950 670.950 355.050 673.050 ;
        RECT 355.950 670.950 358.050 673.050 ;
        RECT 359.250 671.250 360.750 672.150 ;
        RECT 361.950 670.950 364.050 673.050 ;
        RECT 368.400 670.050 369.450 695.400 ;
        RECT 373.950 694.950 376.050 697.050 ;
        RECT 374.400 691.050 375.450 694.950 ;
        RECT 377.400 691.050 378.450 700.950 ;
        RECT 379.950 697.950 382.050 700.050 ;
        RECT 383.250 698.850 384.750 699.750 ;
        RECT 385.950 697.950 388.050 700.050 ;
        RECT 409.950 698.250 412.050 699.150 ;
        RECT 412.950 698.850 415.050 699.750 ;
        RECT 380.400 697.050 381.450 697.950 ;
        RECT 379.950 694.950 382.050 697.050 ;
        RECT 373.950 688.950 376.050 691.050 ;
        RECT 376.950 688.950 379.050 691.050 ;
        RECT 386.400 688.050 387.450 697.950 ;
        RECT 416.400 694.050 417.450 701.400 ;
        RECT 424.950 701.250 426.750 702.150 ;
        RECT 430.950 701.250 433.050 702.150 ;
        RECT 436.950 701.250 439.050 702.150 ;
        RECT 424.950 697.950 427.050 700.050 ;
        RECT 428.250 698.850 430.050 699.750 ;
        RECT 436.950 697.950 439.050 700.050 ;
        RECT 442.950 697.950 445.050 700.050 ;
        RECT 415.950 691.950 418.050 694.050 ;
        RECT 421.950 691.950 424.050 694.050 ;
        RECT 391.950 688.950 394.050 691.050 ;
        RECT 385.950 685.950 388.050 688.050 ;
        RECT 392.400 676.050 393.450 688.950 ;
        RECT 406.950 676.950 409.050 679.050 ;
        RECT 373.950 673.950 376.050 676.050 ;
        RECT 382.950 673.950 385.050 676.050 ;
        RECT 391.950 673.950 394.050 676.050 ;
        RECT 352.950 667.950 355.050 670.050 ;
        RECT 356.250 668.850 357.750 669.750 ;
        RECT 358.950 667.950 361.050 670.050 ;
        RECT 362.250 668.850 364.050 669.750 ;
        RECT 364.950 668.250 366.750 669.150 ;
        RECT 367.950 667.950 370.050 670.050 ;
        RECT 371.250 668.250 373.050 669.150 ;
        RECT 352.950 665.850 355.050 666.750 ;
        RECT 364.950 664.950 367.050 667.050 ;
        RECT 368.250 665.850 369.750 666.750 ;
        RECT 370.950 666.450 373.050 667.050 ;
        RECT 374.400 666.450 375.450 673.950 ;
        RECT 383.250 671.850 384.750 672.750 ;
        RECT 385.950 672.450 388.050 673.050 ;
        RECT 385.950 671.400 390.450 672.450 ;
        RECT 391.950 671.850 394.050 672.750 ;
        RECT 385.950 670.950 388.050 671.400 ;
        RECT 389.400 670.050 390.450 671.400 ;
        RECT 394.950 671.250 397.050 672.150 ;
        RECT 407.400 670.050 408.450 676.950 ;
        RECT 415.950 671.850 418.050 672.750 ;
        RECT 418.950 671.250 421.050 672.150 ;
        RECT 379.950 668.850 382.050 669.750 ;
        RECT 385.950 668.850 388.050 669.750 ;
        RECT 388.950 667.950 391.050 670.050 ;
        RECT 394.950 667.950 397.050 670.050 ;
        RECT 403.950 668.250 405.750 669.150 ;
        RECT 406.950 667.950 409.050 670.050 ;
        RECT 410.250 668.250 412.050 669.150 ;
        RECT 418.950 667.950 421.050 670.050 ;
        RECT 370.950 665.400 375.450 666.450 ;
        RECT 370.950 664.950 373.050 665.400 ;
        RECT 403.950 664.950 406.050 667.050 ;
        RECT 407.250 665.850 408.750 666.750 ;
        RECT 365.400 643.050 366.450 664.950 ;
        RECT 397.950 661.950 400.050 664.050 ;
        RECT 404.400 663.450 405.450 664.950 ;
        RECT 404.400 662.400 408.450 663.450 ;
        RECT 382.950 655.950 385.050 658.050 ;
        RECT 361.950 640.950 364.050 643.050 ;
        RECT 364.950 640.950 367.050 643.050 ;
        RECT 362.400 637.050 363.450 640.950 ;
        RECT 350.400 635.400 354.450 636.450 ;
        RECT 346.950 631.950 349.050 634.050 ;
        RECT 347.400 631.050 348.450 631.950 ;
        RECT 346.950 628.950 349.050 631.050 ;
        RECT 350.250 629.250 352.050 630.150 ;
        RECT 346.950 626.850 348.750 627.750 ;
        RECT 335.400 623.400 339.450 624.450 ;
        RECT 326.400 616.050 327.450 622.950 ;
        RECT 322.950 613.950 325.050 616.050 ;
        RECT 325.950 613.950 328.050 616.050 ;
        RECT 301.950 607.950 304.050 610.050 ;
        RECT 322.950 607.950 325.050 610.050 ;
        RECT 331.950 607.950 334.050 610.050 ;
        RECT 310.950 601.950 313.050 604.050 ;
        RECT 319.950 601.950 322.050 604.050 ;
        RECT 298.950 598.950 301.050 601.050 ;
        RECT 302.250 599.250 303.750 600.150 ;
        RECT 304.950 598.950 307.050 601.050 ;
        RECT 311.250 599.850 312.750 600.750 ;
        RECT 313.950 600.450 316.050 601.050 ;
        RECT 313.950 599.400 318.450 600.450 ;
        RECT 313.950 598.950 316.050 599.400 ;
        RECT 317.400 598.050 318.450 599.400 ;
        RECT 289.950 595.950 292.050 598.050 ;
        RECT 292.950 595.950 295.050 598.050 ;
        RECT 295.950 595.950 298.050 598.050 ;
        RECT 299.250 596.850 300.750 597.750 ;
        RECT 301.950 595.950 304.050 598.050 ;
        RECT 305.250 596.850 307.050 597.750 ;
        RECT 307.950 596.850 310.050 597.750 ;
        RECT 313.950 596.850 316.050 597.750 ;
        RECT 316.950 595.950 319.050 598.050 ;
        RECT 280.950 592.950 283.050 595.050 ;
        RECT 284.250 593.850 285.750 594.750 ;
        RECT 286.950 592.950 289.050 595.050 ;
        RECT 290.250 593.850 292.050 594.750 ;
        RECT 292.950 592.950 295.050 595.050 ;
        RECT 295.950 593.850 298.050 594.750 ;
        RECT 286.950 590.850 289.050 591.750 ;
        RECT 286.950 583.950 289.050 586.050 ;
        RECT 262.950 574.950 265.050 577.050 ;
        RECT 274.950 574.950 277.050 577.050 ;
        RECT 277.950 574.950 280.050 577.050 ;
        RECT 283.950 574.950 286.050 577.050 ;
        RECT 263.400 562.050 264.450 574.950 ;
        RECT 265.950 565.950 268.050 568.050 ;
        RECT 256.950 559.950 259.050 562.050 ;
        RECT 260.250 560.250 261.750 561.150 ;
        RECT 262.950 559.950 265.050 562.050 ;
        RECT 256.950 557.850 258.750 558.750 ;
        RECT 259.950 556.950 262.050 559.050 ;
        RECT 263.250 557.850 265.050 558.750 ;
        RECT 256.950 552.450 259.050 553.050 ;
        RECT 260.400 552.450 261.450 556.950 ;
        RECT 262.950 553.950 265.050 556.050 ;
        RECT 256.950 551.400 261.450 552.450 ;
        RECT 256.950 550.950 259.050 551.400 ;
        RECT 241.950 547.950 244.050 550.050 ;
        RECT 244.950 547.950 247.050 550.050 ;
        RECT 253.950 547.950 256.050 550.050 ;
        RECT 242.400 535.050 243.450 547.950 ;
        RECT 263.400 546.450 264.450 553.950 ;
        RECT 266.400 550.050 267.450 565.950 ;
        RECT 268.950 559.950 271.050 562.050 ;
        RECT 269.400 555.450 270.450 559.950 ;
        RECT 275.400 559.050 276.450 574.950 ;
        RECT 280.950 560.250 283.050 561.150 ;
        RECT 271.950 557.250 273.750 558.150 ;
        RECT 274.950 556.950 277.050 559.050 ;
        RECT 278.250 557.250 279.750 558.150 ;
        RECT 280.950 556.950 283.050 559.050 ;
        RECT 271.950 555.450 274.050 556.050 ;
        RECT 269.400 554.400 274.050 555.450 ;
        RECT 275.250 554.850 276.750 555.750 ;
        RECT 271.950 553.950 274.050 554.400 ;
        RECT 277.950 553.950 280.050 556.050 ;
        RECT 265.950 547.950 268.050 550.050 ;
        RECT 274.950 547.950 277.050 550.050 ;
        RECT 263.400 545.400 267.450 546.450 ;
        RECT 241.950 532.950 244.050 535.050 ;
        RECT 250.950 532.950 253.050 535.050 ;
        RECT 229.950 529.950 232.050 532.050 ;
        RECT 238.950 531.450 241.050 532.050 ;
        RECT 236.400 530.400 241.050 531.450 ;
        RECT 236.400 529.050 237.450 530.400 ;
        RECT 238.950 529.950 241.050 530.400 ;
        RECT 226.950 526.950 229.050 529.050 ;
        RECT 230.250 527.850 231.750 528.750 ;
        RECT 235.950 526.950 238.050 529.050 ;
        RECT 239.250 527.250 240.750 528.150 ;
        RECT 241.950 526.950 244.050 529.050 ;
        RECT 245.250 527.250 246.750 528.150 ;
        RECT 247.950 526.950 250.050 529.050 ;
        RECT 226.950 524.850 229.050 525.750 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 232.950 524.850 235.050 525.750 ;
        RECT 235.950 524.850 237.750 525.750 ;
        RECT 238.950 523.950 241.050 526.050 ;
        RECT 242.250 524.850 243.750 525.750 ;
        RECT 244.950 523.950 247.050 526.050 ;
        RECT 248.250 524.850 250.050 525.750 ;
        RECT 230.400 520.050 231.450 523.950 ;
        RECT 239.400 523.050 240.450 523.950 ;
        RECT 232.950 520.950 235.050 523.050 ;
        RECT 238.950 520.950 241.050 523.050 ;
        RECT 229.950 517.950 232.050 520.050 ;
        RECT 223.950 505.950 226.050 508.050 ;
        RECT 233.400 487.050 234.450 520.950 ;
        RECT 239.400 517.050 240.450 520.950 ;
        RECT 245.400 520.050 246.450 523.950 ;
        RECT 251.400 520.050 252.450 532.950 ;
        RECT 256.950 526.950 259.050 529.050 ;
        RECT 262.950 526.950 265.050 529.050 ;
        RECT 257.400 526.050 258.450 526.950 ;
        RECT 253.950 524.250 255.750 525.150 ;
        RECT 256.950 523.950 259.050 526.050 ;
        RECT 260.250 524.250 262.050 525.150 ;
        RECT 253.950 520.950 256.050 523.050 ;
        RECT 257.250 521.850 258.750 522.750 ;
        RECT 259.950 522.450 262.050 523.050 ;
        RECT 263.400 522.450 264.450 526.950 ;
        RECT 259.950 521.400 264.450 522.450 ;
        RECT 259.950 520.950 262.050 521.400 ;
        RECT 254.400 520.050 255.450 520.950 ;
        RECT 244.950 517.950 247.050 520.050 ;
        RECT 250.950 517.950 253.050 520.050 ;
        RECT 253.950 517.950 256.050 520.050 ;
        RECT 259.950 517.950 262.050 520.050 ;
        RECT 245.400 517.050 246.450 517.950 ;
        RECT 238.950 514.950 241.050 517.050 ;
        RECT 244.950 514.950 247.050 517.050 ;
        RECT 241.950 508.950 244.050 511.050 ;
        RECT 223.950 485.250 225.750 486.150 ;
        RECT 226.950 484.950 229.050 487.050 ;
        RECT 230.250 485.250 231.750 486.150 ;
        RECT 232.950 484.950 235.050 487.050 ;
        RECT 236.250 485.250 238.050 486.150 ;
        RECT 223.950 481.950 226.050 484.050 ;
        RECT 227.250 482.850 228.750 483.750 ;
        RECT 229.950 481.950 232.050 484.050 ;
        RECT 233.250 482.850 234.750 483.750 ;
        RECT 235.950 481.950 238.050 484.050 ;
        RECT 224.400 466.050 225.450 481.950 ;
        RECT 236.400 478.050 237.450 481.950 ;
        RECT 242.400 480.450 243.450 508.950 ;
        RECT 244.950 487.950 247.050 490.050 ;
        RECT 247.950 488.250 250.050 489.150 ;
        RECT 253.950 487.950 256.050 490.050 ;
        RECT 245.400 484.050 246.450 487.950 ;
        RECT 254.400 487.050 255.450 487.950 ;
        RECT 247.950 484.950 250.050 487.050 ;
        RECT 251.250 485.250 252.750 486.150 ;
        RECT 253.950 484.950 256.050 487.050 ;
        RECT 257.250 485.250 259.050 486.150 ;
        RECT 244.950 481.950 247.050 484.050 ;
        RECT 242.400 479.400 246.450 480.450 ;
        RECT 235.950 475.950 238.050 478.050 ;
        RECT 220.950 463.950 223.050 466.050 ;
        RECT 223.950 463.950 226.050 466.050 ;
        RECT 223.950 460.950 226.050 463.050 ;
        RECT 217.950 457.950 220.050 460.050 ;
        RECT 220.950 457.950 223.050 460.050 ;
        RECT 218.400 457.050 219.450 457.950 ;
        RECT 224.400 457.050 225.450 460.950 ;
        RECT 232.950 457.950 235.050 460.050 ;
        RECT 241.950 457.950 244.050 460.050 ;
        RECT 242.400 457.050 243.450 457.950 ;
        RECT 205.950 456.450 208.050 457.050 ;
        RECT 205.950 455.400 210.450 456.450 ;
        RECT 205.950 454.950 208.050 455.400 ;
        RECT 209.400 454.050 210.450 455.400 ;
        RECT 214.950 454.950 217.050 457.050 ;
        RECT 217.950 454.950 220.050 457.050 ;
        RECT 221.250 455.850 222.750 456.750 ;
        RECT 223.950 456.450 226.050 457.050 ;
        RECT 223.950 455.400 228.450 456.450 ;
        RECT 223.950 454.950 226.050 455.400 ;
        RECT 205.950 452.250 207.750 453.150 ;
        RECT 208.950 451.950 211.050 454.050 ;
        RECT 212.250 452.250 214.050 453.150 ;
        RECT 214.950 451.950 217.050 454.050 ;
        RECT 217.950 452.850 220.050 453.750 ;
        RECT 223.950 452.850 226.050 453.750 ;
        RECT 205.950 448.950 208.050 451.050 ;
        RECT 209.250 449.850 210.750 450.750 ;
        RECT 211.950 448.950 214.050 451.050 ;
        RECT 212.400 447.450 213.450 448.950 ;
        RECT 215.400 448.050 216.450 451.950 ;
        RECT 227.400 448.050 228.450 455.400 ;
        RECT 229.950 454.950 232.050 457.050 ;
        RECT 233.250 455.850 234.750 456.750 ;
        RECT 235.950 456.450 238.050 457.050 ;
        RECT 235.950 455.400 240.450 456.450 ;
        RECT 235.950 454.950 238.050 455.400 ;
        RECT 229.950 452.850 232.050 453.750 ;
        RECT 232.950 451.950 235.050 454.050 ;
        RECT 235.950 452.850 238.050 453.750 ;
        RECT 203.400 446.400 213.450 447.450 ;
        RECT 214.950 445.950 217.050 448.050 ;
        RECT 226.950 445.950 229.050 448.050 ;
        RECT 193.950 436.950 196.050 439.050 ;
        RECT 194.400 424.050 195.450 436.950 ;
        RECT 199.950 433.950 202.050 436.050 ;
        RECT 193.950 421.950 196.050 424.050 ;
        RECT 172.950 418.950 175.050 421.050 ;
        RECT 175.950 419.250 178.050 420.150 ;
        RECT 184.950 418.950 187.050 421.050 ;
        RECT 172.950 416.250 174.750 417.150 ;
        RECT 175.950 415.950 178.050 418.050 ;
        RECT 179.250 416.250 180.750 417.150 ;
        RECT 181.950 415.950 184.050 418.050 ;
        RECT 172.950 412.950 175.050 415.050 ;
        RECT 178.950 412.950 181.050 415.050 ;
        RECT 182.250 413.850 184.050 414.750 ;
        RECT 173.400 412.050 174.450 412.950 ;
        RECT 167.400 410.400 171.450 411.450 ;
        RECT 127.950 406.950 130.050 409.050 ;
        RECT 130.950 406.950 133.050 409.050 ;
        RECT 151.950 406.950 154.050 409.050 ;
        RECT 157.950 406.950 160.050 409.050 ;
        RECT 88.950 403.950 91.050 406.050 ;
        RECT 106.950 403.950 109.050 406.050 ;
        RECT 121.950 403.950 124.050 406.050 ;
        RECT 130.950 397.950 133.050 400.050 ;
        RECT 1.950 388.950 4.050 391.050 ;
        RECT 25.950 388.950 28.050 391.050 ;
        RECT 43.950 388.950 46.050 391.050 ;
        RECT 94.950 388.950 97.050 391.050 ;
        RECT 2.400 211.050 3.450 388.950 ;
        RECT 44.400 388.050 45.450 388.950 ;
        RECT 13.950 387.450 16.050 388.050 ;
        RECT 25.950 387.450 28.050 388.050 ;
        RECT 13.950 386.400 18.450 387.450 ;
        RECT 13.950 385.950 16.050 386.400 ;
        RECT 4.950 383.250 7.050 384.150 ;
        RECT 10.950 382.950 13.050 385.050 ;
        RECT 14.250 383.850 16.050 384.750 ;
        RECT 4.950 379.950 7.050 382.050 ;
        RECT 10.950 380.850 13.050 381.750 ;
        RECT 5.400 379.050 6.450 379.950 ;
        RECT 4.950 376.950 7.050 379.050 ;
        RECT 17.400 378.450 18.450 386.400 ;
        RECT 23.400 386.400 28.050 387.450 ;
        RECT 23.400 382.050 24.450 386.400 ;
        RECT 25.950 385.950 28.050 386.400 ;
        RECT 34.950 385.950 37.050 388.050 ;
        RECT 43.950 385.950 46.050 388.050 ;
        RECT 67.950 385.950 70.050 388.050 ;
        RECT 73.950 385.950 76.050 388.050 ;
        RECT 82.950 385.950 85.050 388.050 ;
        RECT 88.950 385.950 91.050 388.050 ;
        RECT 28.950 382.950 31.050 385.050 ;
        RECT 19.950 380.250 21.750 381.150 ;
        RECT 22.950 379.950 25.050 382.050 ;
        RECT 26.250 380.250 28.050 381.150 ;
        RECT 19.950 378.450 22.050 379.050 ;
        RECT 17.400 377.400 22.050 378.450 ;
        RECT 23.250 377.850 24.750 378.750 ;
        RECT 25.950 378.450 28.050 379.050 ;
        RECT 29.400 378.450 30.450 382.950 ;
        RECT 35.400 382.050 36.450 385.950 ;
        RECT 43.950 383.850 46.050 384.750 ;
        RECT 46.950 383.250 49.050 384.150 ;
        RECT 58.950 382.950 61.050 385.050 ;
        RECT 64.950 384.450 67.050 385.050 ;
        RECT 68.400 384.450 69.450 385.950 ;
        RECT 89.400 385.050 90.450 385.950 ;
        RECT 62.250 383.250 63.750 384.150 ;
        RECT 64.950 383.400 69.450 384.450 ;
        RECT 64.950 382.950 67.050 383.400 ;
        RECT 31.950 380.250 33.750 381.150 ;
        RECT 34.950 379.950 37.050 382.050 ;
        RECT 38.250 380.250 40.050 381.150 ;
        RECT 46.950 379.950 49.050 382.050 ;
        RECT 55.950 379.950 58.050 382.050 ;
        RECT 59.250 380.850 60.750 381.750 ;
        RECT 61.950 379.950 64.050 382.050 ;
        RECT 65.250 380.850 67.050 381.750 ;
        RECT 17.400 343.050 18.450 377.400 ;
        RECT 19.950 376.950 22.050 377.400 ;
        RECT 25.950 377.400 30.450 378.450 ;
        RECT 25.950 376.950 28.050 377.400 ;
        RECT 31.950 376.950 34.050 379.050 ;
        RECT 35.250 377.850 36.750 378.750 ;
        RECT 37.950 376.950 40.050 379.050 ;
        RECT 55.950 377.850 58.050 378.750 ;
        RECT 22.950 344.250 25.050 345.150 ;
        RECT 7.950 340.950 10.050 343.050 ;
        RECT 13.950 341.250 15.750 342.150 ;
        RECT 16.950 340.950 19.050 343.050 ;
        RECT 20.250 341.250 21.750 342.150 ;
        RECT 22.950 340.950 25.050 343.050 ;
        RECT 7.950 338.850 10.050 339.750 ;
        RECT 10.950 338.250 13.050 339.150 ;
        RECT 13.950 337.950 16.050 340.050 ;
        RECT 17.250 338.850 18.750 339.750 ;
        RECT 19.950 337.950 22.050 340.050 ;
        RECT 4.950 334.950 7.050 337.050 ;
        RECT 10.950 334.950 13.050 337.050 ;
        RECT 5.400 303.450 6.450 334.950 ;
        RECT 20.400 334.050 21.450 337.950 ;
        RECT 19.950 331.950 22.050 334.050 ;
        RECT 23.400 319.050 24.450 340.950 ;
        RECT 26.400 340.050 27.450 376.950 ;
        RECT 32.400 376.050 33.450 376.950 ;
        RECT 31.950 373.950 34.050 376.050 ;
        RECT 62.400 372.450 63.450 379.950 ;
        RECT 59.400 371.400 63.450 372.450 ;
        RECT 52.950 349.950 55.050 352.050 ;
        RECT 53.400 346.050 54.450 349.950 ;
        RECT 52.950 343.950 55.050 346.050 ;
        RECT 31.950 340.950 34.050 343.050 ;
        RECT 37.950 341.250 40.050 342.150 ;
        RECT 46.950 341.250 49.050 342.150 ;
        RECT 52.950 341.850 55.050 342.750 ;
        RECT 55.950 341.250 58.050 342.150 ;
        RECT 25.950 337.950 28.050 340.050 ;
        RECT 31.950 338.850 34.050 339.750 ;
        RECT 34.950 337.950 37.050 340.050 ;
        RECT 37.950 337.950 40.050 340.050 ;
        RECT 41.250 338.250 43.050 339.150 ;
        RECT 46.950 337.950 49.050 340.050 ;
        RECT 55.950 337.950 58.050 340.050 ;
        RECT 22.950 316.950 25.050 319.050 ;
        RECT 10.950 315.450 13.050 316.050 ;
        RECT 10.950 314.400 15.450 315.450 ;
        RECT 10.950 313.950 13.050 314.400 ;
        RECT 14.400 313.050 15.450 314.400 ;
        RECT 19.950 313.950 22.050 316.050 ;
        RECT 7.950 311.250 10.050 312.150 ;
        RECT 10.950 311.850 13.050 312.750 ;
        RECT 13.950 310.950 16.050 313.050 ;
        RECT 7.950 307.950 10.050 310.050 ;
        RECT 8.400 307.050 9.450 307.950 ;
        RECT 7.950 304.950 10.050 307.050 ;
        RECT 5.400 302.400 9.450 303.450 ;
        RECT 8.400 274.050 9.450 302.400 ;
        RECT 14.400 274.050 15.450 310.950 ;
        RECT 20.400 310.050 21.450 313.950 ;
        RECT 16.950 308.250 18.750 309.150 ;
        RECT 19.950 307.950 22.050 310.050 ;
        RECT 23.250 308.250 25.050 309.150 ;
        RECT 25.950 308.250 27.750 309.150 ;
        RECT 28.950 307.950 31.050 310.050 ;
        RECT 32.250 308.250 34.050 309.150 ;
        RECT 16.950 304.950 19.050 307.050 ;
        RECT 20.250 305.850 21.750 306.750 ;
        RECT 22.950 304.950 25.050 307.050 ;
        RECT 25.950 304.950 28.050 307.050 ;
        RECT 29.250 305.850 30.750 306.750 ;
        RECT 31.950 304.950 34.050 307.050 ;
        RECT 26.400 277.050 27.450 304.950 ;
        RECT 32.400 304.050 33.450 304.950 ;
        RECT 31.950 301.950 34.050 304.050 ;
        RECT 35.400 298.050 36.450 337.950 ;
        RECT 38.400 331.050 39.450 337.950 ;
        RECT 59.400 337.050 60.450 371.400 ;
        RECT 68.400 364.050 69.450 383.400 ;
        RECT 70.950 383.250 73.050 384.150 ;
        RECT 73.950 383.850 76.050 384.750 ;
        RECT 76.950 382.950 79.050 385.050 ;
        RECT 79.950 383.250 82.050 384.150 ;
        RECT 82.950 383.850 85.050 384.750 ;
        RECT 85.950 383.250 87.750 384.150 ;
        RECT 88.950 382.950 91.050 385.050 ;
        RECT 91.950 382.950 94.050 385.050 ;
        RECT 70.950 379.950 73.050 382.050 ;
        RECT 71.400 379.050 72.450 379.950 ;
        RECT 70.950 376.950 73.050 379.050 ;
        RECT 77.400 373.050 78.450 382.950 ;
        RECT 79.950 379.950 82.050 382.050 ;
        RECT 85.950 379.950 88.050 382.050 ;
        RECT 89.250 380.850 91.050 381.750 ;
        RECT 80.400 376.050 81.450 379.950 ;
        RECT 92.400 376.050 93.450 382.950 ;
        RECT 95.400 382.050 96.450 388.950 ;
        RECT 131.400 388.050 132.450 397.950 ;
        RECT 136.950 391.950 139.050 394.050 ;
        RECT 97.950 385.950 100.050 388.050 ;
        RECT 130.950 385.950 133.050 388.050 ;
        RECT 98.400 382.050 99.450 385.950 ;
        RECT 100.950 382.950 103.050 385.050 ;
        RECT 115.950 382.950 118.050 385.050 ;
        RECT 121.950 382.950 124.050 385.050 ;
        RECT 127.950 383.250 130.050 384.150 ;
        RECT 130.950 383.850 133.050 384.750 ;
        RECT 101.400 382.050 102.450 382.950 ;
        RECT 116.400 382.050 117.450 382.950 ;
        RECT 94.950 379.950 97.050 382.050 ;
        RECT 97.950 379.950 100.050 382.050 ;
        RECT 100.950 379.950 103.050 382.050 ;
        RECT 104.250 380.250 106.050 381.150 ;
        RECT 106.950 379.950 109.050 382.050 ;
        RECT 109.950 379.950 112.050 382.050 ;
        RECT 115.950 379.950 118.050 382.050 ;
        RECT 119.250 380.250 121.050 381.150 ;
        RECT 94.950 377.850 96.750 378.750 ;
        RECT 97.950 376.950 100.050 379.050 ;
        RECT 101.250 377.850 102.750 378.750 ;
        RECT 103.950 376.950 106.050 379.050 ;
        RECT 79.950 373.950 82.050 376.050 ;
        RECT 88.950 373.950 91.050 376.050 ;
        RECT 91.950 373.950 94.050 376.050 ;
        RECT 94.950 373.950 97.050 376.050 ;
        RECT 97.950 374.850 100.050 375.750 ;
        RECT 76.950 370.950 79.050 373.050 ;
        RECT 67.950 361.950 70.050 364.050 ;
        RECT 73.950 361.950 76.050 364.050 ;
        RECT 64.950 347.250 67.050 348.150 ;
        RECT 61.950 344.250 63.750 345.150 ;
        RECT 64.950 343.950 67.050 346.050 ;
        RECT 68.250 344.250 69.750 345.150 ;
        RECT 70.950 343.950 73.050 346.050 ;
        RECT 61.950 340.950 64.050 343.050 ;
        RECT 40.950 334.950 43.050 337.050 ;
        RECT 58.950 334.950 61.050 337.050 ;
        RECT 37.950 328.950 40.050 331.050 ;
        RECT 41.400 325.050 42.450 334.950 ;
        RECT 62.400 331.050 63.450 340.950 ;
        RECT 61.950 328.950 64.050 331.050 ;
        RECT 40.950 322.950 43.050 325.050 ;
        RECT 58.950 322.950 61.050 325.050 ;
        RECT 52.950 313.950 55.050 316.050 ;
        RECT 46.950 310.950 49.050 313.050 ;
        RECT 47.400 310.050 48.450 310.950 ;
        RECT 40.950 309.450 43.050 310.050 ;
        RECT 38.400 308.400 43.050 309.450 ;
        RECT 38.400 307.050 39.450 308.400 ;
        RECT 40.950 307.950 43.050 308.400 ;
        RECT 46.950 307.950 49.050 310.050 ;
        RECT 50.250 308.250 52.050 309.150 ;
        RECT 37.950 304.950 40.050 307.050 ;
        RECT 40.950 305.850 42.750 306.750 ;
        RECT 43.950 304.950 46.050 307.050 ;
        RECT 47.250 305.850 48.750 306.750 ;
        RECT 49.950 306.450 52.050 307.050 ;
        RECT 53.400 306.450 54.450 313.950 ;
        RECT 59.400 310.050 60.450 322.950 ;
        RECT 62.400 316.050 63.450 328.950 ;
        RECT 65.400 325.050 66.450 343.950 ;
        RECT 67.950 340.950 70.050 343.050 ;
        RECT 71.250 341.850 73.050 342.750 ;
        RECT 64.950 322.950 67.050 325.050 ;
        RECT 70.950 322.950 73.050 325.050 ;
        RECT 64.950 316.950 67.050 319.050 ;
        RECT 61.950 313.950 64.050 316.050 ;
        RECT 55.950 308.250 57.750 309.150 ;
        RECT 58.950 307.950 61.050 310.050 ;
        RECT 62.250 308.250 64.050 309.150 ;
        RECT 49.950 305.400 54.450 306.450 ;
        RECT 49.950 304.950 52.050 305.400 ;
        RECT 55.950 304.950 58.050 307.050 ;
        RECT 59.250 305.850 60.750 306.750 ;
        RECT 61.950 304.950 64.050 307.050 ;
        RECT 43.950 302.850 46.050 303.750 ;
        RECT 46.950 301.950 49.050 304.050 ;
        RECT 40.950 298.950 43.050 301.050 ;
        RECT 34.950 295.950 37.050 298.050 ;
        RECT 25.950 274.950 28.050 277.050 ;
        RECT 34.950 275.250 37.050 276.150 ;
        RECT 41.400 274.050 42.450 298.950 ;
        RECT 43.950 274.950 46.050 277.050 ;
        RECT 4.950 272.250 7.050 273.150 ;
        RECT 7.950 271.950 10.050 274.050 ;
        RECT 13.950 271.950 16.050 274.050 ;
        RECT 19.950 273.450 22.050 274.050 ;
        RECT 17.400 272.400 22.050 273.450 ;
        RECT 25.950 273.450 28.050 274.050 ;
        RECT 17.400 271.050 18.450 272.400 ;
        RECT 19.950 271.950 22.050 272.400 ;
        RECT 23.250 272.250 24.750 273.150 ;
        RECT 25.950 272.400 30.450 273.450 ;
        RECT 25.950 271.950 28.050 272.400 ;
        RECT 4.950 268.950 7.050 271.050 ;
        RECT 8.250 269.250 9.750 270.150 ;
        RECT 10.950 268.950 13.050 271.050 ;
        RECT 14.250 269.250 16.050 270.150 ;
        RECT 16.950 268.950 19.050 271.050 ;
        RECT 19.950 269.850 21.750 270.750 ;
        RECT 22.950 268.950 25.050 271.050 ;
        RECT 26.250 269.850 28.050 270.750 ;
        RECT 5.400 265.050 6.450 268.950 ;
        RECT 7.950 265.950 10.050 268.050 ;
        RECT 11.250 266.850 12.750 267.750 ;
        RECT 13.950 265.950 16.050 268.050 ;
        RECT 14.400 265.050 15.450 265.950 ;
        RECT 4.950 262.950 7.050 265.050 ;
        RECT 10.950 262.950 13.050 265.050 ;
        RECT 13.950 262.950 16.050 265.050 ;
        RECT 4.950 259.950 7.050 262.050 ;
        RECT 5.400 237.450 6.450 259.950 ;
        RECT 7.950 239.250 10.050 240.150 ;
        RECT 7.950 237.450 10.050 238.050 ;
        RECT 5.400 236.400 10.050 237.450 ;
        RECT 7.950 235.950 10.050 236.400 ;
        RECT 11.400 235.050 12.450 262.950 ;
        RECT 14.400 241.050 15.450 262.950 ;
        RECT 17.400 244.050 18.450 268.950 ;
        RECT 19.950 265.950 22.050 268.050 ;
        RECT 22.950 265.950 25.050 268.050 ;
        RECT 16.950 241.950 19.050 244.050 ;
        RECT 13.950 238.950 16.050 241.050 ;
        RECT 17.250 239.850 19.050 240.750 ;
        RECT 13.950 236.850 16.050 237.750 ;
        RECT 20.400 237.450 21.450 265.950 ;
        RECT 23.400 241.050 24.450 265.950 ;
        RECT 29.400 265.050 30.450 272.400 ;
        RECT 31.950 272.250 33.750 273.150 ;
        RECT 34.950 271.950 37.050 274.050 ;
        RECT 38.250 272.250 39.750 273.150 ;
        RECT 40.950 271.950 43.050 274.050 ;
        RECT 31.950 268.950 34.050 271.050 ;
        RECT 31.950 265.950 34.050 268.050 ;
        RECT 28.950 262.950 31.050 265.050 ;
        RECT 25.950 241.950 28.050 244.050 ;
        RECT 22.950 238.950 25.050 241.050 ;
        RECT 26.400 238.050 27.450 241.950 ;
        RECT 32.400 241.050 33.450 265.950 ;
        RECT 35.400 262.050 36.450 271.950 ;
        RECT 37.950 268.950 40.050 271.050 ;
        RECT 41.250 269.850 43.050 270.750 ;
        RECT 37.950 265.950 40.050 268.050 ;
        RECT 34.950 259.950 37.050 262.050 ;
        RECT 31.950 238.950 34.050 241.050 ;
        RECT 34.950 239.250 37.050 240.150 ;
        RECT 17.400 236.400 21.450 237.450 ;
        RECT 7.950 232.950 10.050 235.050 ;
        RECT 10.950 232.950 13.050 235.050 ;
        RECT 1.950 208.950 4.050 211.050 ;
        RECT 1.950 205.950 4.050 208.050 ;
        RECT 2.400 205.050 3.450 205.950 ;
        RECT 1.950 202.950 4.050 205.050 ;
        RECT 8.400 202.050 9.450 232.950 ;
        RECT 10.950 202.950 13.050 205.050 ;
        RECT 1.950 199.950 4.050 202.050 ;
        RECT 4.950 200.250 7.050 201.150 ;
        RECT 7.950 199.950 10.050 202.050 ;
        RECT 2.400 196.050 3.450 199.950 ;
        RECT 11.400 199.050 12.450 202.950 ;
        RECT 4.950 196.950 7.050 199.050 ;
        RECT 8.250 197.250 9.750 198.150 ;
        RECT 10.950 196.950 13.050 199.050 ;
        RECT 14.250 197.250 16.050 198.150 ;
        RECT 1.950 193.950 4.050 196.050 ;
        RECT 4.950 193.950 7.050 196.050 ;
        RECT 7.950 193.950 10.050 196.050 ;
        RECT 11.250 194.850 12.750 195.750 ;
        RECT 13.950 193.950 16.050 196.050 ;
        RECT 5.400 193.050 6.450 193.950 ;
        RECT 4.950 190.950 7.050 193.050 ;
        RECT 10.950 190.950 13.050 193.050 ;
        RECT 1.950 184.950 4.050 187.050 ;
        RECT 2.400 166.050 3.450 184.950 ;
        RECT 7.950 181.950 10.050 184.050 ;
        RECT 4.950 175.950 7.050 178.050 ;
        RECT 1.950 163.950 4.050 166.050 ;
        RECT 5.400 127.050 6.450 175.950 ;
        RECT 8.400 169.050 9.450 181.950 ;
        RECT 11.400 172.050 12.450 190.950 ;
        RECT 14.400 190.050 15.450 193.950 ;
        RECT 13.950 187.950 16.050 190.050 ;
        RECT 17.400 187.050 18.450 236.400 ;
        RECT 22.950 236.250 24.750 237.150 ;
        RECT 25.950 235.950 28.050 238.050 ;
        RECT 29.250 236.250 31.050 237.150 ;
        RECT 31.950 235.950 34.050 238.050 ;
        RECT 34.950 235.950 37.050 238.050 ;
        RECT 22.950 232.950 25.050 235.050 ;
        RECT 26.250 233.850 27.750 234.750 ;
        RECT 28.950 234.450 31.050 235.050 ;
        RECT 32.400 234.450 33.450 235.950 ;
        RECT 35.400 235.050 36.450 235.950 ;
        RECT 28.950 233.400 33.450 234.450 ;
        RECT 28.950 232.950 31.050 233.400 ;
        RECT 34.950 232.950 37.050 235.050 ;
        RECT 31.950 229.950 34.050 232.050 ;
        RECT 32.400 202.050 33.450 229.950 ;
        RECT 31.950 199.950 34.050 202.050 ;
        RECT 34.950 200.250 37.050 201.150 ;
        RECT 38.400 199.050 39.450 265.950 ;
        RECT 44.400 262.050 45.450 274.950 ;
        RECT 47.400 262.050 48.450 301.950 ;
        RECT 56.400 301.050 57.450 304.950 ;
        RECT 62.400 301.050 63.450 304.950 ;
        RECT 55.950 298.950 58.050 301.050 ;
        RECT 61.950 298.950 64.050 301.050 ;
        RECT 55.950 277.950 58.050 280.050 ;
        RECT 49.950 274.950 52.050 277.050 ;
        RECT 50.400 274.050 51.450 274.950 ;
        RECT 56.400 274.050 57.450 277.950 ;
        RECT 65.400 277.050 66.450 316.950 ;
        RECT 71.400 313.050 72.450 322.950 ;
        RECT 74.400 313.050 75.450 361.950 ;
        RECT 85.950 352.950 88.050 355.050 ;
        RECT 79.950 347.250 82.050 348.150 ;
        RECT 86.400 346.050 87.450 352.950 ;
        RECT 76.950 344.250 78.750 345.150 ;
        RECT 79.950 343.950 82.050 346.050 ;
        RECT 83.250 344.250 84.750 345.150 ;
        RECT 85.950 343.950 88.050 346.050 ;
        RECT 80.400 343.050 81.450 343.950 ;
        RECT 76.950 340.950 79.050 343.050 ;
        RECT 79.950 340.950 82.050 343.050 ;
        RECT 82.950 340.950 85.050 343.050 ;
        RECT 86.250 341.850 88.050 342.750 ;
        RECT 77.400 340.050 78.450 340.950 ;
        RECT 89.400 340.050 90.450 373.950 ;
        RECT 95.400 343.050 96.450 373.950 ;
        RECT 107.400 352.050 108.450 379.950 ;
        RECT 109.950 377.850 111.750 378.750 ;
        RECT 112.950 376.950 115.050 379.050 ;
        RECT 116.250 377.850 117.750 378.750 ;
        RECT 118.950 376.950 121.050 379.050 ;
        RECT 112.950 374.850 115.050 375.750 ;
        RECT 122.400 373.050 123.450 382.950 ;
        RECT 127.950 379.950 130.050 382.050 ;
        RECT 137.400 379.050 138.450 391.950 ;
        RECT 152.400 391.050 153.450 406.950 ;
        RECT 145.950 388.950 148.050 391.050 ;
        RECT 151.950 388.950 154.050 391.050 ;
        RECT 154.950 388.950 157.050 391.050 ;
        RECT 146.400 385.050 147.450 388.950 ;
        RECT 139.950 383.250 142.050 384.150 ;
        RECT 145.950 382.950 148.050 385.050 ;
        RECT 149.250 383.850 151.050 384.750 ;
        RECT 139.950 379.950 142.050 382.050 ;
        RECT 145.950 380.850 148.050 381.750 ;
        RECT 151.950 381.450 154.050 382.050 ;
        RECT 155.400 381.450 156.450 388.950 ;
        RECT 151.950 380.400 156.450 381.450 ;
        RECT 151.950 379.950 154.050 380.400 ;
        RECT 157.950 379.950 160.050 382.050 ;
        RECT 161.250 380.250 163.050 381.150 ;
        RECT 140.400 379.050 141.450 379.950 ;
        RECT 136.950 376.950 139.050 379.050 ;
        RECT 139.950 376.950 142.050 379.050 ;
        RECT 151.950 377.850 153.750 378.750 ;
        RECT 154.950 376.950 157.050 379.050 ;
        RECT 158.250 377.850 159.750 378.750 ;
        RECT 160.950 376.950 163.050 379.050 ;
        RECT 154.950 374.850 157.050 375.750 ;
        RECT 160.950 373.950 163.050 376.050 ;
        RECT 121.950 370.950 124.050 373.050 ;
        RECT 106.950 349.950 109.050 352.050 ;
        RECT 100.950 344.250 103.050 345.150 ;
        RECT 107.400 343.050 108.450 349.950 ;
        RECT 112.950 346.950 115.050 349.050 ;
        RECT 118.950 347.250 121.050 348.150 ;
        RECT 113.400 346.050 114.450 346.950 ;
        RECT 112.950 343.950 115.050 346.050 ;
        RECT 116.250 344.250 117.750 345.150 ;
        RECT 118.950 343.950 121.050 346.050 ;
        RECT 122.250 344.250 124.050 345.150 ;
        RECT 157.950 344.250 160.050 345.150 ;
        RECT 91.950 341.250 93.750 342.150 ;
        RECT 94.950 340.950 97.050 343.050 ;
        RECT 98.250 341.250 99.750 342.150 ;
        RECT 100.950 340.950 103.050 343.050 ;
        RECT 106.950 340.950 109.050 343.050 ;
        RECT 112.950 341.850 114.750 342.750 ;
        RECT 115.950 340.950 118.050 343.050 ;
        RECT 76.950 337.950 79.050 340.050 ;
        RECT 88.950 337.950 91.050 340.050 ;
        RECT 91.950 337.950 94.050 340.050 ;
        RECT 95.250 338.850 96.750 339.750 ;
        RECT 97.950 337.950 100.050 340.050 ;
        RECT 100.950 337.950 103.050 340.050 ;
        RECT 92.400 334.050 93.450 337.950 ;
        RECT 91.950 331.950 94.050 334.050 ;
        RECT 98.400 331.050 99.450 337.950 ;
        RECT 97.950 328.950 100.050 331.050 ;
        RECT 97.950 322.950 100.050 325.050 ;
        RECT 98.400 322.050 99.450 322.950 ;
        RECT 97.950 319.950 100.050 322.050 ;
        RECT 79.950 313.950 82.050 316.050 ;
        RECT 85.950 313.950 88.050 316.050 ;
        RECT 94.950 313.950 97.050 316.050 ;
        RECT 80.400 313.050 81.450 313.950 ;
        RECT 67.950 310.950 70.050 313.050 ;
        RECT 70.950 310.950 73.050 313.050 ;
        RECT 73.950 310.950 76.050 313.050 ;
        RECT 77.250 311.250 78.750 312.150 ;
        RECT 79.950 310.950 82.050 313.050 ;
        RECT 68.400 304.050 69.450 310.950 ;
        RECT 86.400 310.050 87.450 313.950 ;
        RECT 98.400 313.050 99.450 319.950 ;
        RECT 94.950 311.850 96.750 312.750 ;
        RECT 97.950 310.950 100.050 313.050 ;
        RECT 70.950 307.950 73.050 310.050 ;
        RECT 74.250 308.850 75.750 309.750 ;
        RECT 76.950 307.950 79.050 310.050 ;
        RECT 80.250 308.850 82.050 309.750 ;
        RECT 82.950 308.250 84.750 309.150 ;
        RECT 85.950 307.950 88.050 310.050 ;
        RECT 89.250 308.250 91.050 309.150 ;
        RECT 97.950 308.850 100.050 309.750 ;
        RECT 70.950 305.850 73.050 306.750 ;
        RECT 82.950 304.950 85.050 307.050 ;
        RECT 86.250 305.850 87.750 306.750 ;
        RECT 88.950 304.950 91.050 307.050 ;
        RECT 89.400 304.050 90.450 304.950 ;
        RECT 101.400 304.050 102.450 337.950 ;
        RECT 116.400 325.050 117.450 340.950 ;
        RECT 119.400 328.050 120.450 343.950 ;
        RECT 121.950 340.950 124.050 343.050 ;
        RECT 127.950 340.950 130.050 343.050 ;
        RECT 133.950 342.450 136.050 343.050 ;
        RECT 131.400 341.400 136.050 342.450 ;
        RECT 124.950 338.250 127.050 339.150 ;
        RECT 127.950 338.850 130.050 339.750 ;
        RECT 124.950 334.950 127.050 337.050 ;
        RECT 118.950 325.950 121.050 328.050 ;
        RECT 115.950 322.950 118.050 325.050 ;
        RECT 118.950 316.950 121.050 319.050 ;
        RECT 103.950 311.250 106.050 312.150 ;
        RECT 119.400 310.050 120.450 316.950 ;
        RECT 125.400 316.050 126.450 334.950 ;
        RECT 131.400 325.050 132.450 341.400 ;
        RECT 133.950 340.950 136.050 341.400 ;
        RECT 139.950 340.950 142.050 343.050 ;
        RECT 143.250 341.250 145.050 342.150 ;
        RECT 148.950 341.250 150.750 342.150 ;
        RECT 151.950 340.950 154.050 343.050 ;
        RECT 155.250 341.250 156.750 342.150 ;
        RECT 133.950 338.850 136.050 339.750 ;
        RECT 136.950 338.250 139.050 339.150 ;
        RECT 139.950 338.850 141.750 339.750 ;
        RECT 142.950 337.950 145.050 340.050 ;
        RECT 148.950 337.950 151.050 340.050 ;
        RECT 152.250 338.850 153.750 339.750 ;
        RECT 154.950 339.450 157.050 340.050 ;
        RECT 161.400 339.450 162.450 373.950 ;
        RECT 154.950 338.400 162.450 339.450 ;
        RECT 154.950 337.950 157.050 338.400 ;
        RECT 136.950 334.950 139.050 337.050 ;
        RECT 157.950 334.950 160.050 337.050 ;
        RECT 137.400 328.050 138.450 334.950 ;
        RECT 148.950 331.950 151.050 334.050 ;
        RECT 136.950 325.950 139.050 328.050 ;
        RECT 130.950 322.950 133.050 325.050 ;
        RECT 124.950 313.950 127.050 316.050 ;
        RECT 125.400 313.050 126.450 313.950 ;
        RECT 124.950 310.950 127.050 313.050 ;
        RECT 131.400 310.050 132.450 322.950 ;
        RECT 133.950 313.950 136.050 316.050 ;
        RECT 103.950 307.950 106.050 310.050 ;
        RECT 115.950 308.250 117.750 309.150 ;
        RECT 118.950 307.950 121.050 310.050 ;
        RECT 122.250 308.250 124.050 309.150 ;
        RECT 127.950 308.250 129.750 309.150 ;
        RECT 130.950 307.950 133.050 310.050 ;
        RECT 134.400 307.050 135.450 313.950 ;
        RECT 137.400 310.050 138.450 325.950 ;
        RECT 139.950 319.950 142.050 322.050 ;
        RECT 140.400 313.050 141.450 319.950 ;
        RECT 142.950 313.950 145.050 316.050 ;
        RECT 139.950 310.950 142.050 313.050 ;
        RECT 143.250 311.850 144.750 312.750 ;
        RECT 145.950 310.950 148.050 313.050 ;
        RECT 136.950 307.950 139.050 310.050 ;
        RECT 139.950 308.850 142.050 309.750 ;
        RECT 145.950 308.850 148.050 309.750 ;
        RECT 106.950 304.950 109.050 307.050 ;
        RECT 115.950 304.950 118.050 307.050 ;
        RECT 119.250 305.850 120.750 306.750 ;
        RECT 121.950 304.950 124.050 307.050 ;
        RECT 127.950 304.950 130.050 307.050 ;
        RECT 131.250 305.850 132.750 306.750 ;
        RECT 133.950 304.950 136.050 307.050 ;
        RECT 137.250 305.850 139.050 306.750 ;
        RECT 67.950 301.950 70.050 304.050 ;
        RECT 88.950 301.950 91.050 304.050 ;
        RECT 100.950 301.950 103.050 304.050 ;
        RECT 67.950 298.950 70.050 301.050 ;
        RECT 61.950 275.250 64.050 276.150 ;
        RECT 64.950 274.950 67.050 277.050 ;
        RECT 68.400 274.050 69.450 298.950 ;
        RECT 100.950 295.950 103.050 298.050 ;
        RECT 73.950 274.950 76.050 277.050 ;
        RECT 91.950 274.950 94.050 277.050 ;
        RECT 49.950 271.950 52.050 274.050 ;
        RECT 53.250 272.250 54.750 273.150 ;
        RECT 55.950 271.950 58.050 274.050 ;
        RECT 58.950 272.250 60.750 273.150 ;
        RECT 61.950 271.950 64.050 274.050 ;
        RECT 65.250 272.250 66.750 273.150 ;
        RECT 67.950 271.950 70.050 274.050 ;
        RECT 49.950 269.850 51.750 270.750 ;
        RECT 52.950 268.950 55.050 271.050 ;
        RECT 56.250 269.850 58.050 270.750 ;
        RECT 58.950 268.950 61.050 271.050 ;
        RECT 59.400 268.050 60.450 268.950 ;
        RECT 58.950 265.950 61.050 268.050 ;
        RECT 62.400 262.050 63.450 271.950 ;
        RECT 64.950 268.950 67.050 271.050 ;
        RECT 68.250 269.850 70.050 270.750 ;
        RECT 43.950 259.950 46.050 262.050 ;
        RECT 46.950 259.950 49.050 262.050 ;
        RECT 49.950 259.950 52.050 262.050 ;
        RECT 61.950 259.950 64.050 262.050 ;
        RECT 40.950 244.950 43.050 247.050 ;
        RECT 41.400 241.050 42.450 244.950 ;
        RECT 43.950 241.950 46.050 244.050 ;
        RECT 40.950 238.950 43.050 241.050 ;
        RECT 44.250 239.850 46.050 240.750 ;
        RECT 40.950 236.850 43.050 237.750 ;
        RECT 43.950 203.250 46.050 204.150 ;
        RECT 50.400 202.050 51.450 259.950 ;
        RECT 64.950 250.950 67.050 253.050 ;
        RECT 61.950 247.950 64.050 250.050 ;
        RECT 52.950 244.950 55.050 247.050 ;
        RECT 53.400 238.050 54.450 244.950 ;
        RECT 62.400 241.050 63.450 247.950 ;
        RECT 55.950 238.950 58.050 241.050 ;
        RECT 59.250 239.250 60.750 240.150 ;
        RECT 61.950 238.950 64.050 241.050 ;
        RECT 52.950 235.950 55.050 238.050 ;
        RECT 56.250 236.850 57.750 237.750 ;
        RECT 58.950 235.950 61.050 238.050 ;
        RECT 62.250 236.850 64.050 237.750 ;
        RECT 52.950 233.850 55.050 234.750 ;
        RECT 59.400 226.050 60.450 235.950 ;
        RECT 58.950 223.950 61.050 226.050 ;
        RECT 52.950 208.950 55.050 211.050 ;
        RECT 40.950 200.250 42.750 201.150 ;
        RECT 43.950 199.950 46.050 202.050 ;
        RECT 47.250 200.250 48.750 201.150 ;
        RECT 49.950 199.950 52.050 202.050 ;
        RECT 44.400 199.050 45.450 199.950 ;
        RECT 19.950 196.950 22.050 199.050 ;
        RECT 25.950 197.250 27.750 198.150 ;
        RECT 28.950 196.950 31.050 199.050 ;
        RECT 32.250 197.250 33.750 198.150 ;
        RECT 34.950 196.950 37.050 199.050 ;
        RECT 37.950 196.950 40.050 199.050 ;
        RECT 40.950 196.950 43.050 199.050 ;
        RECT 43.950 196.950 46.050 199.050 ;
        RECT 46.950 196.950 49.050 199.050 ;
        RECT 50.250 197.850 52.050 198.750 ;
        RECT 19.950 194.850 22.050 195.750 ;
        RECT 22.950 194.250 25.050 195.150 ;
        RECT 25.950 193.950 28.050 196.050 ;
        RECT 29.250 194.850 30.750 195.750 ;
        RECT 31.950 193.950 34.050 196.050 ;
        RECT 22.950 190.950 25.050 193.050 ;
        RECT 23.400 187.050 24.450 190.950 ;
        RECT 16.950 184.950 19.050 187.050 ;
        RECT 22.950 184.950 25.050 187.050 ;
        RECT 16.950 181.950 19.050 184.050 ;
        RECT 17.400 172.050 18.450 181.950 ;
        RECT 10.950 169.950 13.050 172.050 ;
        RECT 16.950 169.950 19.050 172.050 ;
        RECT 7.950 166.950 10.050 169.050 ;
        RECT 11.250 167.850 12.750 168.750 ;
        RECT 13.950 166.950 16.050 169.050 ;
        RECT 16.950 167.850 18.750 168.750 ;
        RECT 19.950 168.450 22.050 169.050 ;
        RECT 19.950 167.400 24.450 168.450 ;
        RECT 19.950 166.950 22.050 167.400 ;
        RECT 7.950 164.850 10.050 165.750 ;
        RECT 10.950 163.950 13.050 166.050 ;
        RECT 13.950 164.850 16.050 165.750 ;
        RECT 19.950 164.850 22.050 165.750 ;
        RECT 4.950 126.450 7.050 127.050 ;
        RECT 2.400 125.400 7.050 126.450 ;
        RECT 2.400 82.050 3.450 125.400 ;
        RECT 4.950 124.950 7.050 125.400 ;
        RECT 4.950 122.850 7.050 123.750 ;
        RECT 7.950 122.250 10.050 123.150 ;
        RECT 7.950 118.950 10.050 121.050 ;
        RECT 11.400 108.450 12.450 163.950 ;
        RECT 23.400 130.050 24.450 167.400 ;
        RECT 25.950 167.250 28.050 168.150 ;
        RECT 35.400 166.050 36.450 196.950 ;
        RECT 41.400 187.050 42.450 196.950 ;
        RECT 40.950 184.950 43.050 187.050 ;
        RECT 41.400 169.050 42.450 184.950 ;
        RECT 53.400 184.050 54.450 208.950 ;
        RECT 65.400 205.050 66.450 250.950 ;
        RECT 70.950 247.950 73.050 250.050 ;
        RECT 71.400 244.050 72.450 247.950 ;
        RECT 70.950 241.950 73.050 244.050 ;
        RECT 74.400 241.050 75.450 274.950 ;
        RECT 92.400 274.050 93.450 274.950 ;
        RECT 85.950 271.950 88.050 274.050 ;
        RECT 91.950 271.950 94.050 274.050 ;
        RECT 95.250 272.250 96.750 273.150 ;
        RECT 97.950 271.950 100.050 274.050 ;
        RECT 86.400 271.050 87.450 271.950 ;
        RECT 76.950 269.250 78.750 270.150 ;
        RECT 79.950 268.950 82.050 271.050 ;
        RECT 85.950 268.950 88.050 271.050 ;
        RECT 88.950 268.950 91.050 271.050 ;
        RECT 91.950 269.850 93.750 270.750 ;
        RECT 94.950 268.950 97.050 271.050 ;
        RECT 98.250 269.850 100.050 270.750 ;
        RECT 76.950 265.950 79.050 268.050 ;
        RECT 80.250 266.850 82.050 267.750 ;
        RECT 82.950 266.250 85.050 267.150 ;
        RECT 85.950 266.850 88.050 267.750 ;
        RECT 77.400 265.050 78.450 265.950 ;
        RECT 76.950 262.950 79.050 265.050 ;
        RECT 82.950 262.950 85.050 265.050 ;
        RECT 83.400 262.050 84.450 262.950 ;
        RECT 82.950 259.950 85.050 262.050 ;
        RECT 89.400 259.050 90.450 268.950 ;
        RECT 88.950 256.950 91.050 259.050 ;
        RECT 76.950 253.950 79.050 256.050 ;
        RECT 67.950 239.250 70.050 240.150 ;
        RECT 70.950 239.850 73.050 240.750 ;
        RECT 73.950 238.950 76.050 241.050 ;
        RECT 67.950 235.950 70.050 238.050 ;
        RECT 70.950 235.950 73.050 238.050 ;
        RECT 73.950 235.950 76.050 238.050 ;
        RECT 68.400 235.050 69.450 235.950 ;
        RECT 67.950 232.950 70.050 235.050 ;
        RECT 71.400 232.050 72.450 235.950 ;
        RECT 77.400 235.050 78.450 253.950 ;
        RECT 95.400 244.050 96.450 268.950 ;
        RECT 101.400 265.050 102.450 295.950 ;
        RECT 103.950 274.950 106.050 277.050 ;
        RECT 100.950 262.950 103.050 265.050 ;
        RECT 104.400 262.050 105.450 274.950 ;
        RECT 107.400 271.050 108.450 304.950 ;
        RECT 128.400 304.050 129.450 304.950 ;
        RECT 127.950 301.950 130.050 304.050 ;
        RECT 133.950 302.850 136.050 303.750 ;
        RECT 127.950 286.950 130.050 289.050 ;
        RECT 118.950 271.950 121.050 274.050 ;
        RECT 121.950 272.250 124.050 273.150 ;
        RECT 106.950 268.950 109.050 271.050 ;
        RECT 109.950 269.250 112.050 270.150 ;
        RECT 115.950 269.250 118.050 270.150 ;
        RECT 107.400 264.450 108.450 268.950 ;
        RECT 119.400 268.050 120.450 271.950 ;
        RECT 128.400 271.050 129.450 286.950 ;
        RECT 136.950 271.950 139.050 274.050 ;
        RECT 137.400 271.050 138.450 271.950 ;
        RECT 121.950 268.950 124.050 271.050 ;
        RECT 125.250 269.250 126.750 270.150 ;
        RECT 127.950 268.950 130.050 271.050 ;
        RECT 131.250 269.250 133.050 270.150 ;
        RECT 133.950 269.250 135.750 270.150 ;
        RECT 136.950 268.950 139.050 271.050 ;
        RECT 140.250 269.250 141.750 270.150 ;
        RECT 142.950 268.950 145.050 271.050 ;
        RECT 146.250 269.250 148.050 270.150 ;
        RECT 109.950 265.950 112.050 268.050 ;
        RECT 113.250 266.250 114.750 267.150 ;
        RECT 115.950 265.950 118.050 268.050 ;
        RECT 118.950 265.950 121.050 268.050 ;
        RECT 121.950 265.950 124.050 268.050 ;
        RECT 124.950 265.950 127.050 268.050 ;
        RECT 128.250 266.850 129.750 267.750 ;
        RECT 130.950 265.950 133.050 268.050 ;
        RECT 133.950 265.950 136.050 268.050 ;
        RECT 137.250 266.850 138.750 267.750 ;
        RECT 139.950 265.950 142.050 268.050 ;
        RECT 143.250 266.850 144.750 267.750 ;
        RECT 145.950 265.950 148.050 268.050 ;
        RECT 107.400 263.400 111.450 264.450 ;
        RECT 103.950 259.950 106.050 262.050 ;
        RECT 100.950 253.950 103.050 256.050 ;
        RECT 79.950 241.950 82.050 244.050 ;
        RECT 88.950 241.950 91.050 244.050 ;
        RECT 94.950 241.950 97.050 244.050 ;
        RECT 80.400 238.050 81.450 241.950 ;
        RECT 85.950 238.950 88.050 241.050 ;
        RECT 79.950 235.950 82.050 238.050 ;
        RECT 83.250 236.250 85.050 237.150 ;
        RECT 73.950 233.850 75.750 234.750 ;
        RECT 76.950 232.950 79.050 235.050 ;
        RECT 80.250 233.850 81.750 234.750 ;
        RECT 82.950 232.950 85.050 235.050 ;
        RECT 83.400 232.050 84.450 232.950 ;
        RECT 70.950 229.950 73.050 232.050 ;
        RECT 76.950 230.850 79.050 231.750 ;
        RECT 82.950 229.950 85.050 232.050 ;
        RECT 64.950 202.950 67.050 205.050 ;
        RECT 83.400 202.050 84.450 229.950 ;
        RECT 86.400 229.050 87.450 238.950 ;
        RECT 89.400 234.450 90.450 241.950 ;
        RECT 91.950 236.250 93.750 237.150 ;
        RECT 94.950 235.950 97.050 238.050 ;
        RECT 98.250 236.250 100.050 237.150 ;
        RECT 91.950 234.450 94.050 235.050 ;
        RECT 89.400 233.400 94.050 234.450 ;
        RECT 95.250 233.850 96.750 234.750 ;
        RECT 97.950 234.450 100.050 235.050 ;
        RECT 101.400 234.450 102.450 253.950 ;
        RECT 110.400 247.050 111.450 263.400 ;
        RECT 112.950 262.950 115.050 265.050 ;
        RECT 113.400 262.050 114.450 262.950 ;
        RECT 116.400 262.050 117.450 265.950 ;
        RECT 112.950 259.950 115.050 262.050 ;
        RECT 115.950 259.950 118.050 262.050 ;
        RECT 116.400 253.050 117.450 259.950 ;
        RECT 115.950 250.950 118.050 253.050 ;
        RECT 106.950 244.950 109.050 247.050 ;
        RECT 109.950 244.950 112.050 247.050 ;
        RECT 115.950 244.950 118.050 247.050 ;
        RECT 107.400 238.050 108.450 244.950 ;
        RECT 116.400 244.050 117.450 244.950 ;
        RECT 115.950 241.950 118.050 244.050 ;
        RECT 119.400 241.050 120.450 265.950 ;
        RECT 122.400 244.050 123.450 265.950 ;
        RECT 125.400 265.050 126.450 265.950 ;
        RECT 124.950 262.950 127.050 265.050 ;
        RECT 131.400 250.050 132.450 265.950 ;
        RECT 134.400 262.050 135.450 265.950 ;
        RECT 133.950 259.950 136.050 262.050 ;
        RECT 140.400 256.050 141.450 265.950 ;
        RECT 146.400 265.050 147.450 265.950 ;
        RECT 145.950 262.950 148.050 265.050 ;
        RECT 145.950 259.950 148.050 262.050 ;
        RECT 146.400 259.050 147.450 259.950 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 139.950 253.950 142.050 256.050 ;
        RECT 130.950 247.950 133.050 250.050 ;
        RECT 136.950 247.950 139.050 250.050 ;
        RECT 124.950 244.950 127.050 247.050 ;
        RECT 121.950 241.950 124.050 244.050 ;
        RECT 125.400 241.050 126.450 244.950 ;
        RECT 137.400 241.050 138.450 247.950 ;
        RECT 146.400 244.050 147.450 256.950 ;
        RECT 149.400 244.050 150.450 331.950 ;
        RECT 158.400 313.050 159.450 334.950 ;
        RECT 167.400 334.050 168.450 410.400 ;
        RECT 172.950 409.950 175.050 412.050 ;
        RECT 175.950 409.950 178.050 412.050 ;
        RECT 172.950 383.400 175.050 384.300 ;
        RECT 172.950 381.450 175.050 382.200 ;
        RECT 176.400 381.450 177.450 409.950 ;
        RECT 179.400 406.050 180.450 412.950 ;
        RECT 178.950 403.950 181.050 406.050 ;
        RECT 185.400 391.050 186.450 418.950 ;
        RECT 187.950 415.950 190.050 418.050 ;
        RECT 191.250 416.250 192.750 417.150 ;
        RECT 193.950 415.950 196.050 418.050 ;
        RECT 187.950 413.850 189.750 414.750 ;
        RECT 190.950 412.950 193.050 415.050 ;
        RECT 194.250 413.850 196.050 414.750 ;
        RECT 191.400 409.050 192.450 412.950 ;
        RECT 190.950 406.950 193.050 409.050 ;
        RECT 184.950 388.950 187.050 391.050 ;
        RECT 193.950 387.450 196.050 388.050 ;
        RECT 191.400 386.400 196.050 387.450 ;
        RECT 178.950 382.950 181.050 385.200 ;
        RECT 182.250 383.400 184.050 384.300 ;
        RECT 187.950 382.950 190.050 385.200 ;
        RECT 172.950 380.400 177.450 381.450 ;
        RECT 178.950 381.000 180.750 381.900 ;
        RECT 172.950 380.100 175.050 380.400 ;
        RECT 181.950 379.950 184.050 382.200 ;
        RECT 191.400 382.050 192.450 386.400 ;
        RECT 193.950 385.950 196.050 386.400 ;
        RECT 193.950 383.850 196.050 384.750 ;
        RECT 196.950 383.250 199.050 384.150 ;
        RECT 187.950 381.000 190.050 381.900 ;
        RECT 190.950 379.950 193.050 382.050 ;
        RECT 193.950 379.950 196.050 382.050 ;
        RECT 196.950 379.950 199.050 382.050 ;
        RECT 169.950 340.950 172.050 343.050 ;
        RECT 181.950 341.250 184.050 342.150 ;
        RECT 187.950 341.250 190.050 342.150 ;
        RECT 169.950 338.850 172.050 339.750 ;
        RECT 172.950 338.250 175.050 339.150 ;
        RECT 175.950 337.950 178.050 340.050 ;
        RECT 181.950 337.950 184.050 340.050 ;
        RECT 187.950 339.450 190.050 340.050 ;
        RECT 191.400 339.450 192.450 379.950 ;
        RECT 194.400 343.050 195.450 379.950 ;
        RECT 193.950 340.950 196.050 343.050 ;
        RECT 185.250 338.250 186.750 339.150 ;
        RECT 187.950 338.400 192.450 339.450 ;
        RECT 193.950 338.850 196.050 339.750 ;
        RECT 187.950 337.950 190.050 338.400 ;
        RECT 196.950 338.250 199.050 339.150 ;
        RECT 172.950 334.950 175.050 337.050 ;
        RECT 166.950 331.950 169.050 334.050 ;
        RECT 169.950 331.950 172.050 334.050 ;
        RECT 163.950 319.950 166.050 322.050 ;
        RECT 164.400 316.050 165.450 319.950 ;
        RECT 163.950 313.950 166.050 316.050 ;
        RECT 157.950 310.950 160.050 313.050 ;
        RECT 161.250 311.250 163.050 312.150 ;
        RECT 163.950 311.850 166.050 312.750 ;
        RECT 166.950 311.250 169.050 312.150 ;
        RECT 157.950 308.850 159.750 309.750 ;
        RECT 160.950 307.950 163.050 310.050 ;
        RECT 166.950 307.950 169.050 310.050 ;
        RECT 167.400 307.050 168.450 307.950 ;
        RECT 160.950 304.950 163.050 307.050 ;
        RECT 166.950 304.950 169.050 307.050 ;
        RECT 151.950 274.950 154.050 277.050 ;
        RECT 152.400 267.450 153.450 274.950 ;
        RECT 161.400 271.050 162.450 304.950 ;
        RECT 170.400 286.050 171.450 331.950 ;
        RECT 173.400 316.050 174.450 334.950 ;
        RECT 172.950 313.950 175.050 316.050 ;
        RECT 173.400 292.050 174.450 313.950 ;
        RECT 176.400 313.050 177.450 337.950 ;
        RECT 182.400 337.050 183.450 337.950 ;
        RECT 181.950 334.950 184.050 337.050 ;
        RECT 184.950 334.950 187.050 337.050 ;
        RECT 181.950 319.950 184.050 322.050 ;
        RECT 182.400 316.050 183.450 319.950 ;
        RECT 185.400 319.050 186.450 334.950 ;
        RECT 184.950 316.950 187.050 319.050 ;
        RECT 188.400 316.050 189.450 337.950 ;
        RECT 196.950 334.950 199.050 337.050 ;
        RECT 193.950 325.950 196.050 328.050 ;
        RECT 181.950 313.950 184.050 316.050 ;
        RECT 187.950 313.950 190.050 316.050 ;
        RECT 194.400 313.050 195.450 325.950 ;
        RECT 197.400 324.450 198.450 334.950 ;
        RECT 200.400 334.050 201.450 433.950 ;
        RECT 223.950 427.950 226.050 430.050 ;
        RECT 208.950 415.950 211.050 418.050 ;
        RECT 214.950 415.950 217.050 418.050 ;
        RECT 220.950 416.250 223.050 417.150 ;
        RECT 205.950 412.950 208.050 415.050 ;
        RECT 202.950 410.250 205.050 411.150 ;
        RECT 205.950 410.850 208.050 411.750 ;
        RECT 202.950 406.950 205.050 409.050 ;
        RECT 209.400 408.450 210.450 415.950 ;
        RECT 215.400 415.050 216.450 415.950 ;
        RECT 211.950 413.250 213.750 414.150 ;
        RECT 214.950 412.950 217.050 415.050 ;
        RECT 218.250 413.250 219.750 414.150 ;
        RECT 220.950 412.950 223.050 415.050 ;
        RECT 211.950 409.950 214.050 412.050 ;
        RECT 215.250 410.850 216.750 411.750 ;
        RECT 217.950 409.950 220.050 412.050 ;
        RECT 209.400 407.400 213.450 408.450 ;
        RECT 212.400 385.050 213.450 407.400 ;
        RECT 218.400 403.050 219.450 409.950 ;
        RECT 224.400 408.450 225.450 427.950 ;
        RECT 229.950 421.950 232.050 424.050 ;
        RECT 230.400 415.050 231.450 421.950 ;
        RECT 233.400 418.050 234.450 451.950 ;
        RECT 239.400 436.050 240.450 455.400 ;
        RECT 241.950 454.950 244.050 457.050 ;
        RECT 245.400 454.050 246.450 479.400 ;
        RECT 248.400 466.050 249.450 484.950 ;
        RECT 250.950 481.950 253.050 484.050 ;
        RECT 254.250 482.850 255.750 483.750 ;
        RECT 256.950 483.450 259.050 484.050 ;
        RECT 260.400 483.450 261.450 517.950 ;
        RECT 263.400 490.050 264.450 521.400 ;
        RECT 266.400 511.050 267.450 545.400 ;
        RECT 268.950 526.950 271.050 529.050 ;
        RECT 268.950 524.850 271.050 525.750 ;
        RECT 271.950 524.250 274.050 525.150 ;
        RECT 268.950 520.950 271.050 523.050 ;
        RECT 271.950 520.950 274.050 523.050 ;
        RECT 269.400 511.050 270.450 520.950 ;
        RECT 275.400 519.450 276.450 547.950 ;
        RECT 278.400 538.050 279.450 553.950 ;
        RECT 280.950 547.950 283.050 550.050 ;
        RECT 281.400 544.050 282.450 547.950 ;
        RECT 280.950 541.950 283.050 544.050 ;
        RECT 277.950 535.950 280.050 538.050 ;
        RECT 280.950 532.950 283.050 535.050 ;
        RECT 277.950 526.950 280.050 529.050 ;
        RECT 277.950 524.850 280.050 525.750 ;
        RECT 281.400 523.050 282.450 532.950 ;
        RECT 284.400 526.050 285.450 574.950 ;
        RECT 287.400 559.050 288.450 583.950 ;
        RECT 293.400 568.050 294.450 592.950 ;
        RECT 302.400 592.050 303.450 595.950 ;
        RECT 320.400 592.050 321.450 601.950 ;
        RECT 295.950 589.950 298.050 592.050 ;
        RECT 301.950 589.950 304.050 592.050 ;
        RECT 319.950 589.950 322.050 592.050 ;
        RECT 296.400 568.050 297.450 589.950 ;
        RECT 323.400 589.050 324.450 607.950 ;
        RECT 328.950 604.950 331.050 607.050 ;
        RECT 329.400 604.050 330.450 604.950 ;
        RECT 328.950 601.950 331.050 604.050 ;
        RECT 332.400 601.050 333.450 607.950 ;
        RECT 338.400 601.050 339.450 623.400 ;
        RECT 343.950 622.950 346.050 625.050 ;
        RECT 353.400 619.050 354.450 635.400 ;
        RECT 361.950 634.950 364.050 637.050 ;
        RECT 361.950 631.950 364.050 634.050 ;
        RECT 370.950 631.950 373.050 634.050 ;
        RECT 374.250 632.250 375.750 633.150 ;
        RECT 376.950 631.950 379.050 634.050 ;
        RECT 358.950 629.250 361.050 630.150 ;
        RECT 358.950 625.950 361.050 628.050 ;
        RECT 362.400 627.450 363.450 631.950 ;
        RECT 364.950 629.250 367.050 630.150 ;
        RECT 370.950 629.850 372.750 630.750 ;
        RECT 373.950 628.950 376.050 631.050 ;
        RECT 377.250 629.850 379.050 630.750 ;
        RECT 364.950 627.450 367.050 628.050 ;
        RECT 362.400 626.400 367.050 627.450 ;
        RECT 352.950 616.950 355.050 619.050 ;
        RECT 343.950 601.950 346.050 604.050 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 325.950 599.250 328.050 600.150 ;
        RECT 328.950 599.850 331.050 600.750 ;
        RECT 331.950 598.950 334.050 601.050 ;
        RECT 335.250 599.250 336.750 600.150 ;
        RECT 337.950 598.950 340.050 601.050 ;
        RECT 340.950 598.950 343.050 601.050 ;
        RECT 341.400 598.050 342.450 598.950 ;
        RECT 325.950 595.950 328.050 598.050 ;
        RECT 331.950 596.850 333.750 597.750 ;
        RECT 334.950 595.950 337.050 598.050 ;
        RECT 338.250 596.850 339.750 597.750 ;
        RECT 340.950 595.950 343.050 598.050 ;
        RECT 340.950 593.850 343.050 594.750 ;
        RECT 344.400 592.050 345.450 601.950 ;
        RECT 346.950 599.850 349.050 600.750 ;
        RECT 349.950 599.250 352.050 600.150 ;
        RECT 353.400 598.050 354.450 616.950 ;
        RECT 355.950 601.950 358.050 604.050 ;
        RECT 349.950 595.950 352.050 598.050 ;
        RECT 352.950 595.950 355.050 598.050 ;
        RECT 346.950 592.950 349.050 595.050 ;
        RECT 331.950 589.950 334.050 592.050 ;
        RECT 343.950 589.950 346.050 592.050 ;
        RECT 322.950 586.950 325.050 589.050 ;
        RECT 325.950 586.950 328.050 589.050 ;
        RECT 304.950 574.950 307.050 577.050 ;
        RECT 292.950 565.950 295.050 568.050 ;
        RECT 295.950 565.950 298.050 568.050 ;
        RECT 293.400 562.050 294.450 565.950 ;
        RECT 292.950 559.950 295.050 562.050 ;
        RECT 286.950 556.950 289.050 559.050 ;
        RECT 289.950 557.250 292.050 558.150 ;
        RECT 292.950 557.850 295.050 558.750 ;
        RECT 289.950 553.950 292.050 556.050 ;
        RECT 296.400 555.450 297.450 565.950 ;
        RECT 305.400 562.050 306.450 574.950 ;
        RECT 310.950 571.950 313.050 574.050 ;
        RECT 311.400 562.050 312.450 571.950 ;
        RECT 304.950 559.950 307.050 562.050 ;
        RECT 310.950 559.950 313.050 562.050 ;
        RECT 319.950 560.250 322.050 561.150 ;
        RECT 322.950 559.950 325.050 562.050 ;
        RECT 319.950 558.450 322.050 559.050 ;
        RECT 323.400 558.450 324.450 559.950 ;
        RECT 298.950 557.250 301.050 558.150 ;
        RECT 304.950 557.250 306.750 558.150 ;
        RECT 310.950 557.250 312.750 558.150 ;
        RECT 317.250 557.250 318.750 558.150 ;
        RECT 319.950 557.400 324.450 558.450 ;
        RECT 319.950 556.950 322.050 557.400 ;
        RECT 298.950 555.450 301.050 556.050 ;
        RECT 296.400 554.400 301.050 555.450 ;
        RECT 298.950 553.950 301.050 554.400 ;
        RECT 304.950 553.950 307.050 556.050 ;
        RECT 308.250 554.850 310.050 555.750 ;
        RECT 310.950 553.950 313.050 556.050 ;
        RECT 314.250 554.850 315.750 555.750 ;
        RECT 316.950 553.950 319.050 556.050 ;
        RECT 319.950 553.950 322.050 556.050 ;
        RECT 301.950 532.950 304.050 535.050 ;
        RECT 295.950 529.950 298.050 532.050 ;
        RECT 296.400 529.050 297.450 529.950 ;
        RECT 302.400 529.050 303.450 532.950 ;
        RECT 305.400 532.050 306.450 553.950 ;
        RECT 317.400 544.050 318.450 553.950 ;
        RECT 316.950 541.950 319.050 544.050 ;
        RECT 313.950 535.950 316.050 538.050 ;
        RECT 310.950 532.950 313.050 535.050 ;
        RECT 304.950 529.950 307.050 532.050 ;
        RECT 286.950 526.950 289.050 529.050 ;
        RECT 290.250 527.250 291.750 528.150 ;
        RECT 292.950 526.950 295.050 529.050 ;
        RECT 295.950 526.950 298.050 529.050 ;
        RECT 299.250 527.250 300.750 528.150 ;
        RECT 301.950 526.950 304.050 529.050 ;
        RECT 305.250 527.250 306.750 528.150 ;
        RECT 307.950 526.950 310.050 529.050 ;
        RECT 283.950 523.950 286.050 526.050 ;
        RECT 287.250 524.850 288.750 525.750 ;
        RECT 289.950 523.950 292.050 526.050 ;
        RECT 293.250 524.850 295.050 525.750 ;
        RECT 295.950 524.850 297.750 525.750 ;
        RECT 298.950 523.950 301.050 526.050 ;
        RECT 302.250 524.850 303.750 525.750 ;
        RECT 304.950 523.950 307.050 526.050 ;
        RECT 308.250 524.850 310.050 525.750 ;
        RECT 290.400 523.050 291.450 523.950 ;
        RECT 280.950 520.950 283.050 523.050 ;
        RECT 283.950 521.850 286.050 522.750 ;
        RECT 289.950 520.950 292.050 523.050 ;
        RECT 292.950 520.950 295.050 523.050 ;
        RECT 299.400 522.450 300.450 523.950 ;
        RECT 299.400 521.400 303.450 522.450 ;
        RECT 272.400 518.400 276.450 519.450 ;
        RECT 265.950 508.950 268.050 511.050 ;
        RECT 268.950 508.950 271.050 511.050 ;
        RECT 265.950 502.950 268.050 505.050 ;
        RECT 266.400 490.050 267.450 502.950 ;
        RECT 272.400 499.050 273.450 518.400 ;
        RECT 274.950 502.950 277.050 505.050 ;
        RECT 271.950 496.950 274.050 499.050 ;
        RECT 275.400 496.050 276.450 502.950 ;
        RECT 277.950 499.950 280.050 502.050 ;
        RECT 274.950 493.950 277.050 496.050 ;
        RECT 274.950 490.950 277.050 493.050 ;
        RECT 262.950 487.950 265.050 490.050 ;
        RECT 265.950 487.950 268.050 490.050 ;
        RECT 265.950 485.250 268.050 486.150 ;
        RECT 271.950 485.250 274.050 486.150 ;
        RECT 256.950 482.400 261.450 483.450 ;
        RECT 256.950 481.950 259.050 482.400 ;
        RECT 265.950 481.950 268.050 484.050 ;
        RECT 271.950 483.450 274.050 484.050 ;
        RECT 275.400 483.450 276.450 490.950 ;
        RECT 269.250 482.250 270.750 483.150 ;
        RECT 271.950 482.400 276.450 483.450 ;
        RECT 271.950 481.950 274.050 482.400 ;
        RECT 251.400 478.050 252.450 481.950 ;
        RECT 253.950 478.950 256.050 481.050 ;
        RECT 254.400 478.050 255.450 478.950 ;
        RECT 250.950 475.950 253.050 478.050 ;
        RECT 253.950 475.950 256.050 478.050 ;
        RECT 247.950 463.950 250.050 466.050 ;
        RECT 247.950 460.950 250.050 463.050 ;
        RECT 248.400 457.050 249.450 460.950 ;
        RECT 247.950 454.950 250.050 457.050 ;
        RECT 250.950 454.950 253.050 457.050 ;
        RECT 241.950 452.850 244.050 453.750 ;
        RECT 244.950 451.950 247.050 454.050 ;
        RECT 247.950 452.250 250.050 453.150 ;
        RECT 250.950 452.850 253.050 453.750 ;
        RECT 247.950 448.950 250.050 451.050 ;
        RECT 241.950 439.950 244.050 442.050 ;
        RECT 238.950 433.950 241.050 436.050 ;
        RECT 239.400 433.050 240.450 433.950 ;
        RECT 238.950 430.950 241.050 433.050 ;
        RECT 242.400 426.450 243.450 439.950 ;
        RECT 254.400 439.050 255.450 475.950 ;
        RECT 257.400 442.050 258.450 481.950 ;
        RECT 266.400 466.050 267.450 481.950 ;
        RECT 268.950 478.950 271.050 481.050 ;
        RECT 269.400 469.050 270.450 478.950 ;
        RECT 268.950 466.950 271.050 469.050 ;
        RECT 265.950 463.950 268.050 466.050 ;
        RECT 262.950 457.950 265.050 460.050 ;
        RECT 271.950 457.950 274.050 460.050 ;
        RECT 274.950 457.950 277.050 460.050 ;
        RECT 272.400 457.050 273.450 457.950 ;
        RECT 278.400 457.050 279.450 499.950 ;
        RECT 293.400 496.050 294.450 520.950 ;
        RECT 295.950 517.950 298.050 520.050 ;
        RECT 296.400 496.050 297.450 517.950 ;
        RECT 302.400 514.050 303.450 521.400 ;
        RECT 305.400 517.050 306.450 523.950 ;
        RECT 307.950 520.950 310.050 523.050 ;
        RECT 304.950 514.950 307.050 517.050 ;
        RECT 301.950 511.950 304.050 514.050 ;
        RECT 302.400 508.050 303.450 511.950 ;
        RECT 301.950 505.950 304.050 508.050 ;
        RECT 301.950 502.950 304.050 505.050 ;
        RECT 292.950 493.950 295.050 496.050 ;
        RECT 295.950 493.950 298.050 496.050 ;
        RECT 302.400 487.050 303.450 502.950 ;
        RECT 280.950 485.250 283.050 486.150 ;
        RECT 286.950 485.250 289.050 486.150 ;
        RECT 292.950 485.250 294.750 486.150 ;
        RECT 295.950 484.950 298.050 487.050 ;
        RECT 299.250 485.250 300.750 486.150 ;
        RECT 301.950 484.950 304.050 487.050 ;
        RECT 305.250 485.250 307.050 486.150 ;
        RECT 280.950 481.950 283.050 484.050 ;
        RECT 284.250 482.250 285.750 483.150 ;
        RECT 286.950 481.950 289.050 484.050 ;
        RECT 289.950 481.950 292.050 484.050 ;
        RECT 292.950 481.950 295.050 484.050 ;
        RECT 296.250 482.850 297.750 483.750 ;
        RECT 298.950 481.950 301.050 484.050 ;
        RECT 302.250 482.850 303.750 483.750 ;
        RECT 304.950 481.950 307.050 484.050 ;
        RECT 287.400 481.050 288.450 481.950 ;
        RECT 280.950 480.450 283.050 481.050 ;
        RECT 283.950 480.450 286.050 481.050 ;
        RECT 280.950 479.400 286.050 480.450 ;
        RECT 280.950 478.950 283.050 479.400 ;
        RECT 283.950 478.950 286.050 479.400 ;
        RECT 286.950 478.950 289.050 481.050 ;
        RECT 290.400 475.050 291.450 481.950 ;
        RECT 283.950 472.950 286.050 475.050 ;
        RECT 289.950 472.950 292.050 475.050 ;
        RECT 280.950 466.950 283.050 469.050 ;
        RECT 259.950 454.950 262.050 457.050 ;
        RECT 263.250 455.850 264.750 456.750 ;
        RECT 268.950 454.950 271.050 457.050 ;
        RECT 271.950 454.950 274.050 457.050 ;
        RECT 275.250 455.850 276.750 456.750 ;
        RECT 277.950 454.950 280.050 457.050 ;
        RECT 259.950 452.850 262.050 453.750 ;
        RECT 265.950 452.850 268.050 453.750 ;
        RECT 256.950 439.950 259.050 442.050 ;
        RECT 253.950 436.950 256.050 439.050 ;
        RECT 253.950 433.950 256.050 436.050 ;
        RECT 239.400 425.400 243.450 426.450 ;
        RECT 232.950 415.950 235.050 418.050 ;
        RECT 235.950 416.250 238.050 417.150 ;
        RECT 226.950 413.250 228.750 414.150 ;
        RECT 229.950 412.950 232.050 415.050 ;
        RECT 233.250 413.250 234.750 414.150 ;
        RECT 235.950 412.950 238.050 415.050 ;
        RECT 226.950 409.950 229.050 412.050 ;
        RECT 230.250 410.850 231.750 411.750 ;
        RECT 232.950 409.950 235.050 412.050 ;
        RECT 224.400 407.400 228.450 408.450 ;
        RECT 217.950 400.950 220.050 403.050 ;
        RECT 217.950 385.950 220.050 388.050 ;
        RECT 205.950 382.950 208.050 385.050 ;
        RECT 209.250 383.250 210.750 384.150 ;
        RECT 211.950 382.950 214.050 385.050 ;
        RECT 218.400 384.450 219.450 385.950 ;
        RECT 227.400 385.050 228.450 407.400 ;
        RECT 236.400 400.050 237.450 412.950 ;
        RECT 235.950 397.950 238.050 400.050 ;
        RECT 239.400 396.450 240.450 425.400 ;
        RECT 254.400 418.050 255.450 433.950 ;
        RECT 259.950 427.950 262.050 430.050 ;
        RECT 260.400 418.050 261.450 427.950 ;
        RECT 269.400 424.050 270.450 454.950 ;
        RECT 271.950 452.850 274.050 453.750 ;
        RECT 277.950 452.850 280.050 453.750 ;
        RECT 281.400 433.050 282.450 466.950 ;
        RECT 284.400 442.050 285.450 472.950 ;
        RECT 286.950 469.950 289.050 472.050 ;
        RECT 287.400 460.050 288.450 469.950 ;
        RECT 293.400 469.050 294.450 481.950 ;
        RECT 295.950 478.950 298.050 481.050 ;
        RECT 301.950 478.950 304.050 481.050 ;
        RECT 292.950 466.950 295.050 469.050 ;
        RECT 296.400 460.050 297.450 478.950 ;
        RECT 302.400 469.050 303.450 478.950 ;
        RECT 305.400 475.050 306.450 481.950 ;
        RECT 308.400 478.050 309.450 520.950 ;
        RECT 311.400 517.050 312.450 532.950 ;
        RECT 314.400 520.050 315.450 535.950 ;
        RECT 320.400 535.050 321.450 553.950 ;
        RECT 326.400 535.050 327.450 586.950 ;
        RECT 328.950 557.250 331.050 558.150 ;
        RECT 328.950 555.450 331.050 556.050 ;
        RECT 332.400 555.450 333.450 589.950 ;
        RECT 347.400 580.050 348.450 592.950 ;
        RECT 350.400 592.050 351.450 595.950 ;
        RECT 349.950 589.950 352.050 592.050 ;
        RECT 356.400 583.050 357.450 601.950 ;
        RECT 359.400 598.050 360.450 625.950 ;
        RECT 362.400 613.050 363.450 626.400 ;
        RECT 364.950 625.950 367.050 626.400 ;
        RECT 383.400 622.050 384.450 655.950 ;
        RECT 398.400 649.050 399.450 661.950 ;
        RECT 407.400 649.050 408.450 662.400 ;
        RECT 397.950 646.950 400.050 649.050 ;
        RECT 406.950 646.950 409.050 649.050 ;
        RECT 385.950 632.250 388.050 633.150 ;
        RECT 391.950 631.950 394.050 634.050 ;
        RECT 392.400 631.050 393.450 631.950 ;
        RECT 385.950 628.950 388.050 631.050 ;
        RECT 389.250 629.250 390.750 630.150 ;
        RECT 391.950 628.950 394.050 631.050 ;
        RECT 395.250 629.250 397.050 630.150 ;
        RECT 403.950 629.250 406.050 630.150 ;
        RECT 388.950 625.950 391.050 628.050 ;
        RECT 392.250 626.850 393.750 627.750 ;
        RECT 394.950 625.950 397.050 628.050 ;
        RECT 403.950 625.950 406.050 628.050 ;
        RECT 382.950 619.950 385.050 622.050 ;
        RECT 361.950 610.950 364.050 613.050 ;
        RECT 373.950 610.950 376.050 613.050 ;
        RECT 364.950 607.950 367.050 610.050 ;
        RECT 365.400 604.050 366.450 607.950 ;
        RECT 364.950 601.950 367.050 604.050 ;
        RECT 374.400 601.050 375.450 610.950 ;
        RECT 382.950 605.400 385.050 607.500 ;
        RECT 361.950 599.250 364.050 600.150 ;
        RECT 364.950 599.850 367.050 600.750 ;
        RECT 367.950 599.850 370.050 600.750 ;
        RECT 370.950 599.250 373.050 600.150 ;
        RECT 373.950 598.950 376.050 601.050 ;
        RECT 358.950 595.950 361.050 598.050 ;
        RECT 361.950 595.950 364.050 598.050 ;
        RECT 367.950 595.950 370.050 598.050 ;
        RECT 370.950 595.950 373.050 598.050 ;
        RECT 362.400 589.050 363.450 595.950 ;
        RECT 368.400 589.050 369.450 595.950 ;
        RECT 361.950 586.950 364.050 589.050 ;
        RECT 367.950 586.950 370.050 589.050 ;
        RECT 383.400 588.600 384.600 605.400 ;
        RECT 389.400 601.050 390.450 625.950 ;
        RECT 404.400 622.050 405.450 625.950 ;
        RECT 403.950 619.950 406.050 622.050 ;
        RECT 407.400 610.050 408.450 646.950 ;
        RECT 418.950 639.300 421.050 641.400 ;
        RECT 415.950 634.950 418.050 637.050 ;
        RECT 419.550 635.700 420.750 639.300 ;
        RECT 409.950 629.250 412.050 630.150 ;
        RECT 416.400 628.050 417.450 634.950 ;
        RECT 418.950 633.600 421.050 635.700 ;
        RECT 409.950 625.950 412.050 628.050 ;
        RECT 415.950 625.950 418.050 628.050 ;
        RECT 410.400 619.050 411.450 625.950 ;
        RECT 415.950 623.850 418.050 624.750 ;
        RECT 419.550 621.600 420.750 633.600 ;
        RECT 422.400 628.050 423.450 691.950 ;
        RECT 437.400 685.050 438.450 697.950 ;
        RECT 436.950 682.950 439.050 685.050 ;
        RECT 437.400 676.050 438.450 682.950 ;
        RECT 430.950 673.950 433.050 676.050 ;
        RECT 436.950 673.950 439.050 676.050 ;
        RECT 431.400 670.050 432.450 673.950 ;
        RECT 436.950 671.850 439.050 672.750 ;
        RECT 439.950 671.250 442.050 672.150 ;
        RECT 427.950 668.250 429.750 669.150 ;
        RECT 430.950 667.950 433.050 670.050 ;
        RECT 434.250 668.250 436.050 669.150 ;
        RECT 439.950 667.950 442.050 670.050 ;
        RECT 427.950 664.950 430.050 667.050 ;
        RECT 431.250 665.850 432.750 666.750 ;
        RECT 433.950 664.950 436.050 667.050 ;
        RECT 428.400 634.050 429.450 664.950 ;
        RECT 434.400 663.450 435.450 664.950 ;
        RECT 431.400 662.400 435.450 663.450 ;
        RECT 427.950 631.950 430.050 634.050 ;
        RECT 427.950 629.250 430.050 630.150 ;
        RECT 421.950 625.950 424.050 628.050 ;
        RECT 427.950 625.950 430.050 628.050 ;
        RECT 428.400 625.050 429.450 625.950 ;
        RECT 427.950 622.950 430.050 625.050 ;
        RECT 418.950 619.500 421.050 621.600 ;
        RECT 409.950 616.950 412.050 619.050 ;
        RECT 406.950 607.950 409.050 610.050 ;
        RECT 403.950 605.400 406.050 607.500 ;
        RECT 418.950 605.400 421.050 607.500 ;
        RECT 388.950 598.950 391.050 601.050 ;
        RECT 394.950 598.950 397.050 601.050 ;
        RECT 388.950 596.850 391.050 597.750 ;
        RECT 394.950 596.850 397.050 597.750 ;
        RECT 400.950 592.950 403.050 595.050 ;
        RECT 404.250 593.400 405.450 605.400 ;
        RECT 406.950 602.250 409.050 603.150 ;
        RECT 415.950 602.250 418.050 603.150 ;
        RECT 406.950 598.950 409.050 601.050 ;
        RECT 415.950 598.950 418.050 601.050 ;
        RECT 355.950 580.950 358.050 583.050 ;
        RECT 346.950 577.950 349.050 580.050 ;
        RECT 352.950 571.950 355.050 574.050 ;
        RECT 343.950 567.300 346.050 569.400 ;
        RECT 344.550 563.700 345.750 567.300 ;
        RECT 346.950 565.950 349.050 568.050 ;
        RECT 343.950 561.600 346.050 563.700 ;
        RECT 334.950 557.250 337.050 558.150 ;
        RECT 328.950 554.400 333.450 555.450 ;
        RECT 334.950 555.450 337.050 556.050 ;
        RECT 334.950 554.400 339.450 555.450 ;
        RECT 328.950 553.950 331.050 554.400 ;
        RECT 334.950 553.950 337.050 554.400 ;
        RECT 338.400 538.050 339.450 554.400 ;
        RECT 340.950 553.950 343.050 556.050 ;
        RECT 340.950 551.850 343.050 552.750 ;
        RECT 344.550 549.600 345.750 561.600 ;
        RECT 343.950 547.500 346.050 549.600 ;
        RECT 334.950 535.950 337.050 538.050 ;
        RECT 337.950 535.950 340.050 538.050 ;
        RECT 319.950 532.950 322.050 535.050 ;
        RECT 322.950 532.950 325.050 535.050 ;
        RECT 325.950 532.950 328.050 535.050 ;
        RECT 335.400 534.450 336.450 535.950 ;
        RECT 335.400 533.400 339.450 534.450 ;
        RECT 323.400 529.050 324.450 532.950 ;
        RECT 325.950 529.950 328.050 532.050 ;
        RECT 328.950 529.950 331.050 532.050 ;
        RECT 319.950 526.950 322.050 529.050 ;
        RECT 322.950 526.950 325.050 529.050 ;
        RECT 320.400 526.050 321.450 526.950 ;
        RECT 316.950 524.250 318.750 525.150 ;
        RECT 319.950 523.950 322.050 526.050 ;
        RECT 323.250 524.250 325.050 525.150 ;
        RECT 316.950 520.950 319.050 523.050 ;
        RECT 320.250 521.850 321.750 522.750 ;
        RECT 322.950 520.950 325.050 523.050 ;
        RECT 323.400 520.050 324.450 520.950 ;
        RECT 326.400 520.050 327.450 529.950 ;
        RECT 329.400 529.050 330.450 529.950 ;
        RECT 338.400 529.050 339.450 533.400 ;
        RECT 347.400 532.050 348.450 565.950 ;
        RECT 353.400 562.050 354.450 571.950 ;
        RECT 364.950 566.400 367.050 568.500 ;
        RECT 352.950 559.950 355.050 562.050 ;
        RECT 361.950 559.950 364.050 562.050 ;
        RECT 352.950 557.250 355.050 558.150 ;
        RECT 358.950 557.250 361.050 558.150 ;
        RECT 349.950 553.950 352.050 556.050 ;
        RECT 352.950 555.450 355.050 556.050 ;
        RECT 358.950 555.450 361.050 556.050 ;
        RECT 362.400 555.450 363.450 559.950 ;
        RECT 352.950 554.400 357.450 555.450 ;
        RECT 352.950 553.950 355.050 554.400 ;
        RECT 350.400 550.050 351.450 553.950 ;
        RECT 349.950 547.950 352.050 550.050 ;
        RECT 349.950 532.950 352.050 535.050 ;
        RECT 340.950 529.950 343.050 532.050 ;
        RECT 346.950 529.950 349.050 532.050 ;
        RECT 328.950 526.950 331.050 529.050 ;
        RECT 337.950 526.950 340.050 529.050 ;
        RECT 328.950 524.850 331.050 525.750 ;
        RECT 334.950 524.250 337.050 525.150 ;
        RECT 337.950 524.850 340.050 525.750 ;
        RECT 334.950 522.450 337.050 523.050 ;
        RECT 334.950 521.400 339.450 522.450 ;
        RECT 334.950 520.950 337.050 521.400 ;
        RECT 313.950 517.950 316.050 520.050 ;
        RECT 322.950 517.950 325.050 520.050 ;
        RECT 325.950 517.950 328.050 520.050 ;
        RECT 328.950 517.950 331.050 520.050 ;
        RECT 310.950 514.950 313.050 517.050 ;
        RECT 316.950 514.950 319.050 517.050 ;
        RECT 319.950 514.950 322.050 517.050 ;
        RECT 313.950 495.300 316.050 497.400 ;
        RECT 314.550 491.700 315.750 495.300 ;
        RECT 310.950 487.950 313.050 490.050 ;
        RECT 313.950 489.600 316.050 491.700 ;
        RECT 311.400 484.050 312.450 487.950 ;
        RECT 310.950 481.950 313.050 484.050 ;
        RECT 310.950 479.850 313.050 480.750 ;
        RECT 307.950 475.950 310.050 478.050 ;
        RECT 314.550 477.600 315.750 489.600 ;
        RECT 313.950 475.500 316.050 477.600 ;
        RECT 304.950 472.950 307.050 475.050 ;
        RECT 317.400 471.450 318.450 514.950 ;
        RECT 320.400 483.450 321.450 514.950 ;
        RECT 323.400 505.050 324.450 517.950 ;
        RECT 322.950 502.950 325.050 505.050 ;
        RECT 322.950 485.250 325.050 486.150 ;
        RECT 322.950 483.450 325.050 484.050 ;
        RECT 320.400 482.400 325.050 483.450 ;
        RECT 322.950 481.950 325.050 482.400 ;
        RECT 322.950 478.950 325.050 481.050 ;
        RECT 314.400 470.400 318.450 471.450 ;
        RECT 301.950 466.950 304.050 469.050 ;
        RECT 307.950 466.950 310.050 469.050 ;
        RECT 308.400 460.050 309.450 466.950 ;
        RECT 286.950 457.950 289.050 460.050 ;
        RECT 295.950 457.950 298.050 460.050 ;
        RECT 307.950 457.950 310.050 460.050 ;
        RECT 286.950 455.850 289.050 456.750 ;
        RECT 289.950 455.250 292.050 456.150 ;
        RECT 307.950 455.850 310.050 456.750 ;
        RECT 310.950 455.250 313.050 456.150 ;
        RECT 289.950 451.950 292.050 454.050 ;
        RECT 292.950 451.950 295.050 454.050 ;
        RECT 295.950 452.250 297.750 453.150 ;
        RECT 298.950 451.950 301.050 454.050 ;
        RECT 302.250 452.250 304.050 453.150 ;
        RECT 310.950 451.950 313.050 454.050 ;
        RECT 283.950 439.950 286.050 442.050 ;
        RECT 280.950 430.950 283.050 433.050 ;
        RECT 277.950 427.950 280.050 430.050 ;
        RECT 268.950 421.950 271.050 424.050 ;
        RECT 241.950 415.950 244.050 418.050 ;
        RECT 253.950 415.950 256.050 418.050 ;
        RECT 257.250 416.250 258.750 417.150 ;
        RECT 259.950 415.950 262.050 418.050 ;
        RECT 242.400 412.050 243.450 415.950 ;
        RECT 269.400 415.050 270.450 421.950 ;
        RECT 274.950 416.250 277.050 417.150 ;
        RECT 247.950 414.450 250.050 415.050 ;
        RECT 247.950 413.400 252.450 414.450 ;
        RECT 253.950 413.850 255.750 414.750 ;
        RECT 247.950 412.950 250.050 413.400 ;
        RECT 241.950 409.950 244.050 412.050 ;
        RECT 244.950 410.250 247.050 411.150 ;
        RECT 247.950 410.850 250.050 411.750 ;
        RECT 251.400 409.050 252.450 413.400 ;
        RECT 256.950 412.950 259.050 415.050 ;
        RECT 260.250 413.850 262.050 414.750 ;
        RECT 265.950 413.250 267.750 414.150 ;
        RECT 268.950 412.950 271.050 415.050 ;
        RECT 272.250 413.250 273.750 414.150 ;
        RECT 274.950 412.950 277.050 415.050 ;
        RECT 253.950 409.950 256.050 412.050 ;
        RECT 244.950 406.950 247.050 409.050 ;
        RECT 250.950 406.950 253.050 409.050 ;
        RECT 236.400 395.400 240.450 396.450 ;
        RECT 220.950 384.450 223.050 385.050 ;
        RECT 218.400 383.400 223.050 384.450 ;
        RECT 205.950 380.850 207.750 381.750 ;
        RECT 208.950 379.950 211.050 382.050 ;
        RECT 212.250 380.850 213.750 381.750 ;
        RECT 209.400 343.050 210.450 379.950 ;
        RECT 214.950 377.850 217.050 378.750 ;
        RECT 218.400 358.050 219.450 383.400 ;
        RECT 220.950 382.950 223.050 383.400 ;
        RECT 224.250 383.250 225.750 384.150 ;
        RECT 226.950 382.950 229.050 385.050 ;
        RECT 232.950 382.950 235.050 385.050 ;
        RECT 220.950 380.850 222.750 381.750 ;
        RECT 223.950 379.950 226.050 382.050 ;
        RECT 227.250 380.850 228.750 381.750 ;
        RECT 217.950 355.950 220.050 358.050 ;
        RECT 202.950 341.250 204.750 342.150 ;
        RECT 205.950 340.950 208.050 343.050 ;
        RECT 208.950 340.950 211.050 343.050 ;
        RECT 211.950 340.950 214.050 343.050 ;
        RECT 214.950 341.250 217.050 342.150 ;
        RECT 220.950 341.250 223.050 342.150 ;
        RECT 202.950 337.950 205.050 340.050 ;
        RECT 206.250 338.850 208.050 339.750 ;
        RECT 208.950 338.250 211.050 339.150 ;
        RECT 211.950 338.850 214.050 339.750 ;
        RECT 214.950 337.950 217.050 340.050 ;
        RECT 218.250 338.250 219.750 339.150 ;
        RECT 220.950 337.950 223.050 340.050 ;
        RECT 215.400 337.050 216.450 337.950 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 214.950 334.950 217.050 337.050 ;
        RECT 217.950 334.950 220.050 337.050 ;
        RECT 221.400 334.050 222.450 337.950 ;
        RECT 224.400 337.050 225.450 379.950 ;
        RECT 229.950 377.850 232.050 378.750 ;
        RECT 226.950 355.950 229.050 358.050 ;
        RECT 223.950 334.950 226.050 337.050 ;
        RECT 227.400 336.450 228.450 355.950 ;
        RECT 233.400 343.050 234.450 382.950 ;
        RECT 236.400 373.050 237.450 395.400 ;
        RECT 238.950 385.950 241.050 388.050 ;
        RECT 247.950 385.950 250.050 388.050 ;
        RECT 239.400 379.050 240.450 385.950 ;
        RECT 241.950 382.950 244.050 385.050 ;
        RECT 245.250 383.250 247.050 384.150 ;
        RECT 247.950 383.850 250.050 384.750 ;
        RECT 250.950 383.250 253.050 384.150 ;
        RECT 241.950 380.850 243.750 381.750 ;
        RECT 244.950 379.950 247.050 382.050 ;
        RECT 250.950 379.950 253.050 382.050 ;
        RECT 238.950 376.950 241.050 379.050 ;
        RECT 235.950 370.950 238.050 373.050 ;
        RECT 245.400 367.050 246.450 379.950 ;
        RECT 238.950 364.950 241.050 367.050 ;
        RECT 244.950 364.950 247.050 367.050 ;
        RECT 239.400 343.050 240.450 364.950 ;
        RECT 229.950 341.250 231.750 342.150 ;
        RECT 232.950 340.950 235.050 343.050 ;
        RECT 236.250 341.250 237.750 342.150 ;
        RECT 238.950 340.950 241.050 343.050 ;
        RECT 247.950 342.450 250.050 343.050 ;
        RECT 242.250 341.250 244.050 342.150 ;
        RECT 245.400 341.400 250.050 342.450 ;
        RECT 229.950 337.950 232.050 340.050 ;
        RECT 233.250 338.850 234.750 339.750 ;
        RECT 235.950 337.950 238.050 340.050 ;
        RECT 239.250 338.850 240.750 339.750 ;
        RECT 241.950 339.450 244.050 340.050 ;
        RECT 245.400 339.450 246.450 341.400 ;
        RECT 247.950 340.950 250.050 341.400 ;
        RECT 241.950 338.400 246.450 339.450 ;
        RECT 247.950 338.850 250.050 339.750 ;
        RECT 241.950 337.950 244.050 338.400 ;
        RECT 250.950 338.250 253.050 339.150 ;
        RECT 227.400 335.400 231.450 336.450 ;
        RECT 199.950 331.950 202.050 334.050 ;
        RECT 220.950 331.950 223.050 334.050 ;
        RECT 197.400 323.400 201.450 324.450 ;
        RECT 175.950 310.950 178.050 313.050 ;
        RECT 179.250 311.250 181.050 312.150 ;
        RECT 181.950 311.850 184.050 312.750 ;
        RECT 184.950 311.250 187.050 312.150 ;
        RECT 187.950 310.950 190.050 313.050 ;
        RECT 191.250 311.250 192.750 312.150 ;
        RECT 193.950 310.950 196.050 313.050 ;
        RECT 175.950 308.850 177.750 309.750 ;
        RECT 178.950 307.950 181.050 310.050 ;
        RECT 184.950 307.950 187.050 310.050 ;
        RECT 187.950 308.850 189.750 309.750 ;
        RECT 190.950 307.950 193.050 310.050 ;
        RECT 194.250 308.850 195.750 309.750 ;
        RECT 196.950 307.950 199.050 310.050 ;
        RECT 185.400 307.050 186.450 307.950 ;
        RECT 184.950 304.950 187.050 307.050 ;
        RECT 172.950 289.950 175.050 292.050 ;
        RECT 187.950 286.950 190.050 289.050 ;
        RECT 163.950 283.950 166.050 286.050 ;
        RECT 169.950 283.950 172.050 286.050 ;
        RECT 164.400 271.050 165.450 283.950 ;
        RECT 175.950 271.950 178.050 274.050 ;
        RECT 154.950 269.250 156.750 270.150 ;
        RECT 157.950 268.950 160.050 271.050 ;
        RECT 160.950 268.950 163.050 271.050 ;
        RECT 163.950 268.950 166.050 271.050 ;
        RECT 166.950 269.250 169.050 270.150 ;
        RECT 172.950 269.250 175.050 270.150 ;
        RECT 154.950 267.450 157.050 268.050 ;
        RECT 152.400 266.400 157.050 267.450 ;
        RECT 158.250 266.850 160.050 267.750 ;
        RECT 154.950 265.950 157.050 266.400 ;
        RECT 160.950 266.250 163.050 267.150 ;
        RECT 163.950 266.850 166.050 267.750 ;
        RECT 166.950 265.950 169.050 268.050 ;
        RECT 170.250 266.250 171.750 267.150 ;
        RECT 172.950 265.950 175.050 268.050 ;
        RECT 160.950 262.950 163.050 265.050 ;
        RECT 169.950 262.950 172.050 265.050 ;
        RECT 161.400 262.050 162.450 262.950 ;
        RECT 173.400 262.050 174.450 265.950 ;
        RECT 160.950 259.950 163.050 262.050 ;
        RECT 163.950 259.950 166.050 262.050 ;
        RECT 172.950 259.950 175.050 262.050 ;
        RECT 151.950 247.950 154.050 250.050 ;
        RECT 139.950 241.950 142.050 244.050 ;
        RECT 142.950 241.950 145.050 244.050 ;
        RECT 145.950 241.950 148.050 244.050 ;
        RECT 148.950 241.950 151.050 244.050 ;
        RECT 112.950 238.950 115.050 241.050 ;
        RECT 116.250 239.850 117.750 240.750 ;
        RECT 118.950 240.450 121.050 241.050 ;
        RECT 118.950 239.400 123.450 240.450 ;
        RECT 118.950 238.950 121.050 239.400 ;
        RECT 103.950 236.250 105.750 237.150 ;
        RECT 106.950 235.950 109.050 238.050 ;
        RECT 110.250 236.250 112.050 237.150 ;
        RECT 112.950 236.850 115.050 237.750 ;
        RECT 115.950 235.950 118.050 238.050 ;
        RECT 118.950 236.850 121.050 237.750 ;
        RECT 91.950 232.950 94.050 233.400 ;
        RECT 97.950 233.400 102.450 234.450 ;
        RECT 97.950 232.950 100.050 233.400 ;
        RECT 103.950 232.950 106.050 235.050 ;
        RECT 107.250 233.850 108.750 234.750 ;
        RECT 109.950 232.950 112.050 235.050 ;
        RECT 97.950 229.950 100.050 232.050 ;
        RECT 85.950 226.950 88.050 229.050 ;
        RECT 98.400 226.050 99.450 229.950 ;
        RECT 104.400 229.050 105.450 232.950 ;
        RECT 112.950 229.950 115.050 232.050 ;
        RECT 103.950 226.950 106.050 229.050 ;
        RECT 97.950 223.950 100.050 226.050 ;
        RECT 94.950 202.950 97.050 205.050 ;
        RECT 67.950 199.950 70.050 202.050 ;
        RECT 82.950 199.950 85.050 202.050 ;
        RECT 88.950 201.450 91.050 202.050 ;
        RECT 86.250 200.250 87.750 201.150 ;
        RECT 88.950 200.400 93.450 201.450 ;
        RECT 88.950 199.950 91.050 200.400 ;
        RECT 61.950 196.950 64.050 199.050 ;
        RECT 58.950 193.950 61.050 196.050 ;
        RECT 61.950 194.850 64.050 195.750 ;
        RECT 64.950 194.250 67.050 195.150 ;
        RECT 52.950 181.950 55.050 184.050 ;
        RECT 59.400 178.050 60.450 193.950 ;
        RECT 68.400 193.050 69.450 199.950 ;
        RECT 92.400 199.050 93.450 200.400 ;
        RECT 70.950 197.250 72.750 198.150 ;
        RECT 73.950 196.950 76.050 199.050 ;
        RECT 79.950 196.950 82.050 199.050 ;
        RECT 82.950 197.850 84.750 198.750 ;
        RECT 85.950 196.950 88.050 199.050 ;
        RECT 89.250 197.850 91.050 198.750 ;
        RECT 91.950 196.950 94.050 199.050 ;
        RECT 70.950 193.950 73.050 196.050 ;
        RECT 74.250 194.850 76.050 195.750 ;
        RECT 76.950 194.250 79.050 195.150 ;
        RECT 79.950 194.850 82.050 195.750 ;
        RECT 64.950 190.950 67.050 193.050 ;
        RECT 67.950 190.950 70.050 193.050 ;
        RECT 65.400 190.050 66.450 190.950 ;
        RECT 71.400 190.050 72.450 193.950 ;
        RECT 76.950 190.950 79.050 193.050 ;
        RECT 64.950 187.950 67.050 190.050 ;
        RECT 70.950 187.950 73.050 190.050 ;
        RECT 73.950 187.950 76.050 190.050 ;
        RECT 58.950 175.950 61.050 178.050 ;
        RECT 49.950 172.950 52.050 175.050 ;
        RECT 58.950 172.950 61.050 175.050 ;
        RECT 50.400 172.050 51.450 172.950 ;
        RECT 49.950 169.950 52.050 172.050 ;
        RECT 59.400 169.050 60.450 172.950 ;
        RECT 40.950 166.950 43.050 169.050 ;
        RECT 49.950 167.850 52.050 168.750 ;
        RECT 52.950 167.250 55.050 168.150 ;
        RECT 58.950 166.950 61.050 169.050 ;
        RECT 62.250 167.250 63.750 168.150 ;
        RECT 64.950 166.950 67.050 169.050 ;
        RECT 25.950 163.950 28.050 166.050 ;
        RECT 34.950 163.950 37.050 166.050 ;
        RECT 37.950 164.250 39.750 165.150 ;
        RECT 40.950 163.950 43.050 166.050 ;
        RECT 46.950 165.450 49.050 166.050 ;
        RECT 52.950 165.450 55.050 166.050 ;
        RECT 46.950 164.400 55.050 165.450 ;
        RECT 46.950 163.950 49.050 164.400 ;
        RECT 52.950 163.950 55.050 164.400 ;
        RECT 55.950 163.950 58.050 166.050 ;
        RECT 58.950 164.850 60.750 165.750 ;
        RECT 61.950 163.950 64.050 166.050 ;
        RECT 65.250 164.850 66.750 165.750 ;
        RECT 67.950 163.950 70.050 166.050 ;
        RECT 37.950 160.950 40.050 163.050 ;
        RECT 41.250 161.850 42.750 162.750 ;
        RECT 43.950 160.950 46.050 163.050 ;
        RECT 47.250 161.850 49.050 162.750 ;
        RECT 28.950 131.250 31.050 132.150 ;
        RECT 38.400 130.050 39.450 160.950 ;
        RECT 43.950 158.850 46.050 159.750 ;
        RECT 43.950 142.950 46.050 145.050 ;
        RECT 49.950 142.950 52.050 145.050 ;
        RECT 22.950 129.450 25.050 130.050 ;
        RECT 20.400 128.400 25.050 129.450 ;
        RECT 13.950 124.950 16.050 127.050 ;
        RECT 13.950 122.850 16.050 123.750 ;
        RECT 16.950 122.250 19.050 123.150 ;
        RECT 20.400 121.050 21.450 128.400 ;
        RECT 22.950 127.950 25.050 128.400 ;
        RECT 26.250 128.250 27.750 129.150 ;
        RECT 28.950 127.950 31.050 130.050 ;
        RECT 32.250 128.250 34.050 129.150 ;
        RECT 34.950 127.950 37.050 130.050 ;
        RECT 37.950 127.950 40.050 130.050 ;
        RECT 22.950 125.850 24.750 126.750 ;
        RECT 25.950 124.950 28.050 127.050 ;
        RECT 28.950 124.950 31.050 127.050 ;
        RECT 31.950 124.950 34.050 127.050 ;
        RECT 26.400 124.050 27.450 124.950 ;
        RECT 25.950 121.950 28.050 124.050 ;
        RECT 16.950 118.950 19.050 121.050 ;
        RECT 19.950 118.950 22.050 121.050 ;
        RECT 17.400 115.050 18.450 118.950 ;
        RECT 16.950 112.950 19.050 115.050 ;
        RECT 20.400 108.450 21.450 118.950 ;
        RECT 11.400 107.400 15.450 108.450 ;
        RECT 10.950 97.950 13.050 100.050 ;
        RECT 4.950 94.950 7.050 97.050 ;
        RECT 1.950 79.950 4.050 82.050 ;
        RECT 1.950 76.950 4.050 79.050 ;
        RECT 2.400 55.050 3.450 76.950 ;
        RECT 5.400 64.050 6.450 94.950 ;
        RECT 11.400 94.050 12.450 97.950 ;
        RECT 14.400 94.050 15.450 107.400 ;
        RECT 17.400 107.400 21.450 108.450 ;
        RECT 17.400 94.050 18.450 107.400 ;
        RECT 19.950 103.950 22.050 106.050 ;
        RECT 20.400 97.050 21.450 103.950 ;
        RECT 29.400 100.050 30.450 124.950 ;
        RECT 32.400 118.050 33.450 124.950 ;
        RECT 35.400 121.050 36.450 127.950 ;
        RECT 44.400 127.050 45.450 142.950 ;
        RECT 37.950 124.950 40.050 127.050 ;
        RECT 43.950 124.950 46.050 127.050 ;
        RECT 47.250 125.250 49.050 126.150 ;
        RECT 37.950 122.850 40.050 123.750 ;
        RECT 40.950 122.250 43.050 123.150 ;
        RECT 43.950 122.850 45.750 123.750 ;
        RECT 46.950 121.950 49.050 124.050 ;
        RECT 34.950 118.950 37.050 121.050 ;
        RECT 40.950 118.950 43.050 121.050 ;
        RECT 31.950 115.950 34.050 118.050 ;
        RECT 47.400 115.050 48.450 121.950 ;
        RECT 50.400 118.050 51.450 142.950 ;
        RECT 56.400 133.050 57.450 163.950 ;
        RECT 62.400 162.450 63.450 163.950 ;
        RECT 62.400 161.400 66.450 162.450 ;
        RECT 67.950 161.850 70.050 162.750 ;
        RECT 61.950 157.950 64.050 160.050 ;
        RECT 55.950 130.950 58.050 133.050 ;
        RECT 56.400 130.050 57.450 130.950 ;
        RECT 62.400 130.050 63.450 157.950 ;
        RECT 55.950 127.950 58.050 130.050 ;
        RECT 59.250 128.250 60.750 129.150 ;
        RECT 61.950 127.950 64.050 130.050 ;
        RECT 65.400 127.050 66.450 161.400 ;
        RECT 67.950 128.250 70.050 129.150 ;
        RECT 74.400 127.050 75.450 187.950 ;
        RECT 86.400 187.050 87.450 196.950 ;
        RECT 92.400 196.050 93.450 196.950 ;
        RECT 91.950 193.950 94.050 196.050 ;
        RECT 95.400 193.050 96.450 202.950 ;
        RECT 98.400 198.450 99.450 223.950 ;
        RECT 100.950 200.250 103.050 201.150 ;
        RECT 100.950 198.450 103.050 199.050 ;
        RECT 98.400 197.400 103.050 198.450 ;
        RECT 100.950 196.950 103.050 197.400 ;
        RECT 104.250 197.250 105.750 198.150 ;
        RECT 106.950 196.950 109.050 199.050 ;
        RECT 110.250 197.250 112.050 198.150 ;
        RECT 103.950 193.950 106.050 196.050 ;
        RECT 107.250 194.850 108.750 195.750 ;
        RECT 109.950 193.950 112.050 196.050 ;
        RECT 94.950 190.950 97.050 193.050 ;
        RECT 113.400 190.050 114.450 229.950 ;
        RECT 116.400 196.050 117.450 235.950 ;
        RECT 122.400 232.050 123.450 239.400 ;
        RECT 124.950 238.950 127.050 241.050 ;
        RECT 128.250 239.250 129.750 240.150 ;
        RECT 130.950 238.950 133.050 241.050 ;
        RECT 134.250 239.250 135.750 240.150 ;
        RECT 136.950 238.950 139.050 241.050 ;
        RECT 124.950 236.850 126.750 237.750 ;
        RECT 127.950 235.950 130.050 238.050 ;
        RECT 131.250 236.850 132.750 237.750 ;
        RECT 133.950 235.950 136.050 238.050 ;
        RECT 137.250 236.850 139.050 237.750 ;
        RECT 128.400 235.050 129.450 235.950 ;
        RECT 127.950 232.950 130.050 235.050 ;
        RECT 121.950 229.950 124.050 232.050 ;
        RECT 118.950 197.250 121.050 198.150 ;
        RECT 124.950 197.250 127.050 198.150 ;
        RECT 128.400 196.050 129.450 232.950 ;
        RECT 134.400 232.050 135.450 235.950 ;
        RECT 140.400 235.050 141.450 241.950 ;
        RECT 143.400 241.050 144.450 241.950 ;
        RECT 142.950 238.950 145.050 241.050 ;
        RECT 146.250 239.850 147.750 240.750 ;
        RECT 148.950 238.950 151.050 241.050 ;
        RECT 142.950 236.850 145.050 237.750 ;
        RECT 148.950 236.850 151.050 237.750 ;
        RECT 139.950 232.950 142.050 235.050 ;
        RECT 133.950 229.950 136.050 232.050 ;
        RECT 133.950 220.950 136.050 223.050 ;
        RECT 134.400 202.050 135.450 220.950 ;
        RECT 152.400 202.050 153.450 247.950 ;
        RECT 157.950 244.950 160.050 247.050 ;
        RECT 154.950 241.950 157.050 244.050 ;
        RECT 155.400 226.050 156.450 241.950 ;
        RECT 158.400 235.050 159.450 244.950 ;
        RECT 164.400 244.050 165.450 259.950 ;
        RECT 176.400 259.050 177.450 271.950 ;
        RECT 178.950 269.250 181.050 270.150 ;
        RECT 184.950 269.250 187.050 270.150 ;
        RECT 178.950 265.950 181.050 268.050 ;
        RECT 184.950 267.450 187.050 268.050 ;
        RECT 188.400 267.450 189.450 286.950 ;
        RECT 191.400 271.050 192.450 307.950 ;
        RECT 196.950 305.850 199.050 306.750 ;
        RECT 200.400 283.050 201.450 323.400 ;
        RECT 226.950 316.950 229.050 319.050 ;
        RECT 227.400 313.050 228.450 316.950 ;
        RECT 214.950 312.450 217.050 313.050 ;
        RECT 212.400 311.400 217.050 312.450 ;
        RECT 202.950 308.250 204.750 309.150 ;
        RECT 205.950 307.950 208.050 310.050 ;
        RECT 209.250 308.250 211.050 309.150 ;
        RECT 202.950 304.950 205.050 307.050 ;
        RECT 206.250 305.850 207.750 306.750 ;
        RECT 208.950 304.950 211.050 307.050 ;
        RECT 203.400 304.050 204.450 304.950 ;
        RECT 202.950 301.950 205.050 304.050 ;
        RECT 199.950 280.950 202.050 283.050 ;
        RECT 193.950 271.950 196.050 274.050 ;
        RECT 199.950 273.450 202.050 274.050 ;
        RECT 203.400 273.450 204.450 301.950 ;
        RECT 209.400 277.050 210.450 304.950 ;
        RECT 212.400 304.050 213.450 311.400 ;
        RECT 214.950 310.950 217.050 311.400 ;
        RECT 218.250 311.250 219.750 312.150 ;
        RECT 220.950 310.950 223.050 313.050 ;
        RECT 224.250 311.250 225.750 312.150 ;
        RECT 226.950 310.950 229.050 313.050 ;
        RECT 214.950 308.850 216.750 309.750 ;
        RECT 217.950 307.950 220.050 310.050 ;
        RECT 221.250 308.850 222.750 309.750 ;
        RECT 223.950 307.950 226.050 310.050 ;
        RECT 227.250 308.850 229.050 309.750 ;
        RECT 218.400 307.050 219.450 307.950 ;
        RECT 224.400 307.050 225.450 307.950 ;
        RECT 217.950 304.950 220.050 307.050 ;
        RECT 223.950 304.950 226.050 307.050 ;
        RECT 211.950 301.950 214.050 304.050 ;
        RECT 230.400 298.050 231.450 335.400 ;
        RECT 232.950 334.950 235.050 337.050 ;
        RECT 250.950 334.950 253.050 337.050 ;
        RECT 233.400 331.050 234.450 334.950 ;
        RECT 232.950 328.950 235.050 331.050 ;
        RECT 250.950 328.950 253.050 331.050 ;
        RECT 232.950 313.950 235.050 316.050 ;
        RECT 238.950 313.950 241.050 316.050 ;
        RECT 233.400 310.050 234.450 313.950 ;
        RECT 235.950 311.250 238.050 312.150 ;
        RECT 238.950 311.850 241.050 312.750 ;
        RECT 241.950 311.250 243.750 312.150 ;
        RECT 244.950 310.950 247.050 313.050 ;
        RECT 232.950 307.950 235.050 310.050 ;
        RECT 235.950 307.950 238.050 310.050 ;
        RECT 241.950 307.950 244.050 310.050 ;
        RECT 245.250 308.850 247.050 309.750 ;
        RECT 236.400 304.050 237.450 307.950 ;
        RECT 242.400 307.050 243.450 307.950 ;
        RECT 241.950 304.950 244.050 307.050 ;
        RECT 235.950 301.950 238.050 304.050 ;
        RECT 241.950 298.950 244.050 301.050 ;
        RECT 229.950 295.950 232.050 298.050 ;
        RECT 211.950 280.950 214.050 283.050 ;
        RECT 232.950 280.950 235.050 283.050 ;
        RECT 208.950 274.950 211.050 277.050 ;
        RECT 212.400 274.050 213.450 280.950 ;
        RECT 220.950 277.950 223.050 280.050 ;
        RECT 217.950 274.950 220.050 277.050 ;
        RECT 197.250 272.250 198.750 273.150 ;
        RECT 199.950 272.400 204.450 273.450 ;
        RECT 199.950 271.950 202.050 272.400 ;
        RECT 190.950 268.950 193.050 271.050 ;
        RECT 193.950 269.850 195.750 270.750 ;
        RECT 196.950 268.950 199.050 271.050 ;
        RECT 200.250 269.850 202.050 270.750 ;
        RECT 203.400 267.450 204.450 272.400 ;
        RECT 205.950 271.950 208.050 274.050 ;
        RECT 209.250 272.250 210.750 273.150 ;
        RECT 211.950 271.950 214.050 274.050 ;
        RECT 214.950 271.950 217.050 274.050 ;
        RECT 205.950 269.850 207.750 270.750 ;
        RECT 208.950 268.950 211.050 271.050 ;
        RECT 212.250 269.850 214.050 270.750 ;
        RECT 182.250 266.250 183.750 267.150 ;
        RECT 184.950 266.400 189.450 267.450 ;
        RECT 200.400 266.400 204.450 267.450 ;
        RECT 184.950 265.950 187.050 266.400 ;
        RECT 166.950 256.950 169.050 259.050 ;
        RECT 175.950 256.950 178.050 259.050 ;
        RECT 163.950 241.950 166.050 244.050 ;
        RECT 160.950 239.250 163.050 240.150 ;
        RECT 163.950 239.850 166.050 240.750 ;
        RECT 160.950 235.950 163.050 238.050 ;
        RECT 157.950 232.950 160.050 235.050 ;
        RECT 154.950 223.950 157.050 226.050 ;
        RECT 161.400 205.050 162.450 235.950 ;
        RECT 167.400 205.050 168.450 256.950 ;
        RECT 175.950 253.950 178.050 256.050 ;
        RECT 176.400 247.050 177.450 253.950 ;
        RECT 179.400 250.050 180.450 265.950 ;
        RECT 181.950 262.950 184.050 265.050 ;
        RECT 184.950 259.950 187.050 262.050 ;
        RECT 181.950 250.950 184.050 253.050 ;
        RECT 178.950 247.950 181.050 250.050 ;
        RECT 172.950 244.950 175.050 247.050 ;
        RECT 175.950 244.950 178.050 247.050 ;
        RECT 182.400 246.450 183.450 250.950 ;
        RECT 179.400 245.400 183.450 246.450 ;
        RECT 173.400 244.050 174.450 244.950 ;
        RECT 172.950 241.950 175.050 244.050 ;
        RECT 175.950 241.950 178.050 244.050 ;
        RECT 169.950 239.250 172.050 240.150 ;
        RECT 172.950 239.850 175.050 240.750 ;
        RECT 169.950 235.950 172.050 238.050 ;
        RECT 172.950 235.950 175.050 238.050 ;
        RECT 170.400 235.050 171.450 235.950 ;
        RECT 173.400 235.050 174.450 235.950 ;
        RECT 169.950 232.950 172.050 235.050 ;
        RECT 172.950 232.950 175.050 235.050 ;
        RECT 160.950 202.950 163.050 205.050 ;
        RECT 166.950 202.950 169.050 205.050 ;
        RECT 176.400 202.050 177.450 241.950 ;
        RECT 179.400 241.050 180.450 245.400 ;
        RECT 181.950 243.450 184.050 244.050 ;
        RECT 185.400 243.450 186.450 259.950 ;
        RECT 187.950 253.950 190.050 256.050 ;
        RECT 181.950 242.400 186.450 243.450 ;
        RECT 181.950 241.950 184.050 242.400 ;
        RECT 188.400 241.050 189.450 253.950 ;
        RECT 190.950 250.950 193.050 253.050 ;
        RECT 178.950 238.950 181.050 241.050 ;
        RECT 182.250 239.850 183.750 240.750 ;
        RECT 184.950 238.950 187.050 241.050 ;
        RECT 187.950 238.950 190.050 241.050 ;
        RECT 191.400 238.050 192.450 250.950 ;
        RECT 178.950 236.850 181.050 237.750 ;
        RECT 184.950 236.850 187.050 237.750 ;
        RECT 187.950 236.250 189.750 237.150 ;
        RECT 190.950 235.950 193.050 238.050 ;
        RECT 194.250 236.250 196.050 237.150 ;
        RECT 187.950 232.950 190.050 235.050 ;
        RECT 191.250 233.850 192.750 234.750 ;
        RECT 193.950 232.950 196.050 235.050 ;
        RECT 188.400 226.050 189.450 232.950 ;
        RECT 187.950 223.950 190.050 226.050 ;
        RECT 190.950 223.950 193.050 226.050 ;
        RECT 191.400 202.050 192.450 223.950 ;
        RECT 194.400 223.050 195.450 232.950 ;
        RECT 200.400 229.050 201.450 266.400 ;
        RECT 215.400 265.050 216.450 271.950 ;
        RECT 202.950 262.950 205.050 265.050 ;
        RECT 214.950 262.950 217.050 265.050 ;
        RECT 203.400 244.050 204.450 262.950 ;
        RECT 214.950 244.950 217.050 247.050 ;
        RECT 202.950 241.950 205.050 244.050 ;
        RECT 203.400 241.050 204.450 241.950 ;
        RECT 215.400 241.050 216.450 244.950 ;
        RECT 202.950 238.950 205.050 241.050 ;
        RECT 206.250 239.250 207.750 240.150 ;
        RECT 208.950 238.950 211.050 241.050 ;
        RECT 212.250 239.250 213.750 240.150 ;
        RECT 214.950 238.950 217.050 241.050 ;
        RECT 202.950 236.850 204.750 237.750 ;
        RECT 205.950 235.950 208.050 238.050 ;
        RECT 209.250 236.850 210.750 237.750 ;
        RECT 211.950 235.950 214.050 238.050 ;
        RECT 215.250 236.850 217.050 237.750 ;
        RECT 206.400 232.050 207.450 235.950 ;
        RECT 202.950 229.950 205.050 232.050 ;
        RECT 205.950 229.950 208.050 232.050 ;
        RECT 199.950 226.950 202.050 229.050 ;
        RECT 193.950 220.950 196.050 223.050 ;
        RECT 193.950 217.950 196.050 220.050 ;
        RECT 133.950 199.950 136.050 202.050 ;
        RECT 136.950 199.950 139.050 202.050 ;
        RECT 142.950 199.950 145.050 202.050 ;
        RECT 151.950 199.950 154.050 202.050 ;
        RECT 160.950 200.250 163.050 201.150 ;
        RECT 166.950 199.950 169.050 202.050 ;
        RECT 175.950 199.950 178.050 202.050 ;
        RECT 187.950 199.950 190.050 202.050 ;
        RECT 190.950 199.950 193.050 202.050 ;
        RECT 130.950 196.950 133.050 199.050 ;
        RECT 137.400 196.050 138.450 199.950 ;
        RECT 139.950 197.250 142.050 198.150 ;
        RECT 142.950 197.850 145.050 198.750 ;
        RECT 145.950 196.950 148.050 199.050 ;
        RECT 148.950 197.250 151.050 198.150 ;
        RECT 151.950 197.250 153.750 198.150 ;
        RECT 154.950 196.950 157.050 199.050 ;
        RECT 158.250 197.250 159.750 198.150 ;
        RECT 160.950 196.950 163.050 199.050 ;
        RECT 115.950 193.950 118.050 196.050 ;
        RECT 118.950 193.950 121.050 196.050 ;
        RECT 122.250 194.250 123.750 195.150 ;
        RECT 124.950 193.950 127.050 196.050 ;
        RECT 127.950 193.950 130.050 196.050 ;
        RECT 130.950 194.850 133.050 195.750 ;
        RECT 133.950 194.250 136.050 195.150 ;
        RECT 136.950 193.950 139.050 196.050 ;
        RECT 139.950 193.950 142.050 196.050 ;
        RECT 142.950 193.950 145.050 196.050 ;
        RECT 112.950 187.950 115.050 190.050 ;
        RECT 85.950 184.950 88.050 187.050 ;
        RECT 79.950 181.950 82.050 184.050 ;
        RECT 85.950 181.950 88.050 184.050 ;
        RECT 97.950 181.950 100.050 184.050 ;
        RECT 76.950 167.250 79.050 168.150 ;
        RECT 76.950 163.950 79.050 166.050 ;
        RECT 77.400 133.050 78.450 163.950 ;
        RECT 80.400 157.050 81.450 181.950 ;
        RECT 82.950 175.950 85.050 178.050 ;
        RECT 83.400 169.050 84.450 175.950 ;
        RECT 86.400 172.050 87.450 181.950 ;
        RECT 85.950 169.950 88.050 172.050 ;
        RECT 82.950 166.950 85.050 169.050 ;
        RECT 86.250 167.850 88.050 168.750 ;
        RECT 82.950 164.850 85.050 165.750 ;
        RECT 85.950 163.950 88.050 166.050 ;
        RECT 88.950 164.250 90.750 165.150 ;
        RECT 91.950 163.950 94.050 166.050 ;
        RECT 95.250 164.250 97.050 165.150 ;
        RECT 86.400 162.450 87.450 163.950 ;
        RECT 88.950 162.450 91.050 163.050 ;
        RECT 86.400 161.400 91.050 162.450 ;
        RECT 92.250 161.850 93.750 162.750 ;
        RECT 94.950 162.450 97.050 163.050 ;
        RECT 98.400 162.450 99.450 181.950 ;
        RECT 109.950 166.950 112.050 169.050 ;
        RECT 110.400 166.050 111.450 166.950 ;
        RECT 106.950 164.250 108.750 165.150 ;
        RECT 109.950 163.950 112.050 166.050 ;
        RECT 115.950 163.950 118.050 166.050 ;
        RECT 88.950 160.950 91.050 161.400 ;
        RECT 94.950 161.400 99.450 162.450 ;
        RECT 94.950 160.950 97.050 161.400 ;
        RECT 106.950 160.950 109.050 163.050 ;
        RECT 110.250 161.850 111.750 162.750 ;
        RECT 112.950 160.950 115.050 163.050 ;
        RECT 116.250 161.850 118.050 162.750 ;
        RECT 79.950 154.950 82.050 157.050 ;
        RECT 88.950 133.950 91.050 136.050 ;
        RECT 76.950 130.950 79.050 133.050 ;
        RECT 55.950 125.850 57.750 126.750 ;
        RECT 58.950 124.950 61.050 127.050 ;
        RECT 62.250 125.850 64.050 126.750 ;
        RECT 64.950 124.950 67.050 127.050 ;
        RECT 67.950 124.950 70.050 127.050 ;
        RECT 71.250 125.250 72.750 126.150 ;
        RECT 73.950 124.950 76.050 127.050 ;
        RECT 77.250 125.250 79.050 126.150 ;
        RECT 79.950 125.250 82.050 126.150 ;
        RECT 85.950 125.250 88.050 126.150 ;
        RECT 70.950 121.950 73.050 124.050 ;
        RECT 74.250 122.850 75.750 123.750 ;
        RECT 76.950 121.950 79.050 124.050 ;
        RECT 79.950 121.950 82.050 124.050 ;
        RECT 85.950 123.450 88.050 124.050 ;
        RECT 89.400 123.450 90.450 133.950 ;
        RECT 100.950 131.250 103.050 132.150 ;
        RECT 94.950 129.450 97.050 130.050 ;
        RECT 83.250 122.250 84.750 123.150 ;
        RECT 85.950 122.400 90.450 123.450 ;
        RECT 92.400 128.400 97.050 129.450 ;
        RECT 85.950 121.950 88.050 122.400 ;
        RECT 77.400 121.050 78.450 121.950 ;
        RECT 80.400 121.050 81.450 121.950 ;
        RECT 76.950 118.950 79.050 121.050 ;
        RECT 79.950 118.950 82.050 121.050 ;
        RECT 82.950 118.950 85.050 121.050 ;
        RECT 49.950 115.950 52.050 118.050 ;
        RECT 46.950 112.950 49.050 115.050 ;
        RECT 47.400 106.050 48.450 112.950 ;
        RECT 46.950 105.450 49.050 106.050 ;
        RECT 46.950 104.400 51.450 105.450 ;
        RECT 46.950 103.950 49.050 104.400 ;
        RECT 46.950 100.950 49.050 103.050 ;
        RECT 28.950 97.950 31.050 100.050 ;
        RECT 29.400 97.050 30.450 97.950 ;
        RECT 19.950 94.950 22.050 97.050 ;
        RECT 23.250 95.250 24.750 96.150 ;
        RECT 25.950 94.950 28.050 97.050 ;
        RECT 28.950 94.950 31.050 97.050 ;
        RECT 31.950 94.950 34.050 97.050 ;
        RECT 34.950 94.950 37.050 97.050 ;
        RECT 40.950 94.950 43.050 97.050 ;
        RECT 7.950 92.250 9.750 93.150 ;
        RECT 10.950 91.950 13.050 94.050 ;
        RECT 13.950 91.950 16.050 94.050 ;
        RECT 16.950 91.950 19.050 94.050 ;
        RECT 19.950 92.850 21.750 93.750 ;
        RECT 22.950 91.950 25.050 94.050 ;
        RECT 26.250 92.850 27.750 93.750 ;
        RECT 28.950 93.450 31.050 94.050 ;
        RECT 32.400 93.450 33.450 94.950 ;
        RECT 35.400 94.050 36.450 94.950 ;
        RECT 41.400 94.050 42.450 94.950 ;
        RECT 28.950 92.400 33.450 93.450 ;
        RECT 28.950 91.950 31.050 92.400 ;
        RECT 7.950 88.950 10.050 91.050 ;
        RECT 11.250 89.850 12.750 90.750 ;
        RECT 13.950 88.950 16.050 91.050 ;
        RECT 17.250 89.850 19.050 90.750 ;
        RECT 8.400 87.450 9.450 88.950 ;
        RECT 8.400 86.400 12.450 87.450 ;
        RECT 13.950 86.850 16.050 87.750 ;
        RECT 7.950 82.950 10.050 85.050 ;
        RECT 8.400 79.050 9.450 82.950 ;
        RECT 7.950 76.950 10.050 79.050 ;
        RECT 4.950 61.950 7.050 64.050 ;
        RECT 4.950 58.950 7.050 61.050 ;
        RECT 5.400 58.050 6.450 58.950 ;
        RECT 11.400 58.050 12.450 86.400 ;
        RECT 23.400 82.050 24.450 91.950 ;
        RECT 28.950 89.850 31.050 90.750 ;
        RECT 22.950 79.950 25.050 82.050 ;
        RECT 32.400 79.050 33.450 92.400 ;
        RECT 34.950 91.950 37.050 94.050 ;
        RECT 37.950 91.950 40.050 94.050 ;
        RECT 40.950 91.950 43.050 94.050 ;
        RECT 44.250 92.250 46.050 93.150 ;
        RECT 38.400 91.050 39.450 91.950 ;
        RECT 34.950 89.850 36.750 90.750 ;
        RECT 37.950 88.950 40.050 91.050 ;
        RECT 41.250 89.850 42.750 90.750 ;
        RECT 43.950 88.950 46.050 91.050 ;
        RECT 37.950 86.850 40.050 87.750 ;
        RECT 31.950 76.950 34.050 79.050 ;
        RECT 40.950 73.950 43.050 76.050 ;
        RECT 13.950 61.950 16.050 64.050 ;
        RECT 4.950 55.950 7.050 58.050 ;
        RECT 8.250 56.250 9.750 57.150 ;
        RECT 10.950 55.950 13.050 58.050 ;
        RECT 1.950 52.950 4.050 55.050 ;
        RECT 4.950 53.850 6.750 54.750 ;
        RECT 7.950 52.950 10.050 55.050 ;
        RECT 11.250 53.850 13.050 54.750 ;
        RECT 1.950 49.950 4.050 52.050 ;
        RECT 2.400 49.050 3.450 49.950 ;
        RECT 1.950 46.950 4.050 49.050 ;
        RECT 10.950 37.950 13.050 40.050 ;
        RECT 7.950 25.950 10.050 28.050 ;
        RECT 11.400 25.050 12.450 37.950 ;
        RECT 14.400 25.050 15.450 61.950 ;
        RECT 16.950 58.950 19.050 61.050 ;
        RECT 22.950 59.250 25.050 60.150 ;
        RECT 17.400 58.050 18.450 58.950 ;
        RECT 41.400 58.050 42.450 73.950 ;
        RECT 43.950 61.950 46.050 64.050 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 20.250 56.250 21.750 57.150 ;
        RECT 22.950 55.950 25.050 58.050 ;
        RECT 26.250 56.250 28.050 57.150 ;
        RECT 37.950 56.250 40.050 57.150 ;
        RECT 40.950 55.950 43.050 58.050 ;
        RECT 44.400 57.450 45.450 61.950 ;
        RECT 47.400 61.050 48.450 100.950 ;
        RECT 50.400 97.050 51.450 104.400 ;
        RECT 83.400 103.050 84.450 118.950 ;
        RECT 82.950 100.950 85.050 103.050 ;
        RECT 67.950 97.950 70.050 100.050 ;
        RECT 49.950 94.950 52.050 97.050 ;
        RECT 53.250 95.250 54.750 96.150 ;
        RECT 55.950 94.950 58.050 97.050 ;
        RECT 64.950 94.950 67.050 97.050 ;
        RECT 67.950 95.850 70.050 96.750 ;
        RECT 70.950 95.250 73.050 96.150 ;
        RECT 73.950 94.950 76.050 97.050 ;
        RECT 79.950 94.950 82.050 97.050 ;
        RECT 88.950 94.950 91.050 97.050 ;
        RECT 49.950 92.850 51.750 93.750 ;
        RECT 52.950 91.950 55.050 94.050 ;
        RECT 56.250 92.850 57.750 93.750 ;
        RECT 58.950 93.450 61.050 94.050 ;
        RECT 58.950 92.400 63.450 93.450 ;
        RECT 58.950 91.950 61.050 92.400 ;
        RECT 53.400 82.050 54.450 91.950 ;
        RECT 58.950 89.850 61.050 90.750 ;
        RECT 62.400 88.050 63.450 92.400 ;
        RECT 61.950 85.950 64.050 88.050 ;
        RECT 65.400 85.050 66.450 94.950 ;
        RECT 67.950 91.950 70.050 94.050 ;
        RECT 70.950 91.950 73.050 94.050 ;
        RECT 64.950 82.950 67.050 85.050 ;
        RECT 52.950 79.950 55.050 82.050 ;
        RECT 68.400 76.050 69.450 91.950 ;
        RECT 74.400 85.050 75.450 94.950 ;
        RECT 76.950 91.950 79.050 94.050 ;
        RECT 80.400 91.050 81.450 94.950 ;
        RECT 82.950 91.950 85.050 94.050 ;
        RECT 86.250 92.250 88.050 93.150 ;
        RECT 76.950 89.850 78.750 90.750 ;
        RECT 79.950 88.950 82.050 91.050 ;
        RECT 83.250 89.850 84.750 90.750 ;
        RECT 85.950 88.950 88.050 91.050 ;
        RECT 79.950 86.850 82.050 87.750 ;
        RECT 73.950 82.950 76.050 85.050 ;
        RECT 67.950 73.950 70.050 76.050 ;
        RECT 86.400 73.050 87.450 88.950 ;
        RECT 89.400 88.050 90.450 94.950 ;
        RECT 92.400 94.050 93.450 128.400 ;
        RECT 94.950 127.950 97.050 128.400 ;
        RECT 98.250 128.250 99.750 129.150 ;
        RECT 100.950 127.950 103.050 130.050 ;
        RECT 107.400 129.450 108.450 160.950 ;
        RECT 112.950 158.850 115.050 159.750 ;
        RECT 119.400 136.050 120.450 193.950 ;
        RECT 125.400 193.050 126.450 193.950 ;
        RECT 121.950 190.950 124.050 193.050 ;
        RECT 124.950 190.950 127.050 193.050 ;
        RECT 133.950 192.450 136.050 193.050 ;
        RECT 136.950 192.450 139.050 193.050 ;
        RECT 133.950 191.400 139.050 192.450 ;
        RECT 133.950 190.950 136.050 191.400 ;
        RECT 136.950 190.950 139.050 191.400 ;
        RECT 122.400 178.050 123.450 190.950 ;
        RECT 121.950 175.950 124.050 178.050 ;
        RECT 127.950 175.950 130.050 178.050 ;
        RECT 128.400 172.050 129.450 175.950 ;
        RECT 127.950 169.950 130.050 172.050 ;
        RECT 136.950 169.950 139.050 172.050 ;
        RECT 121.950 166.950 124.050 169.050 ;
        RECT 124.950 167.250 127.050 168.150 ;
        RECT 127.950 167.850 130.050 168.750 ;
        RECT 133.950 167.250 136.050 168.150 ;
        RECT 136.950 167.850 139.050 168.750 ;
        RECT 118.950 133.950 121.050 136.050 ;
        RECT 122.400 133.050 123.450 166.950 ;
        RECT 124.950 163.950 127.050 166.050 ;
        RECT 133.950 163.950 136.050 166.050 ;
        RECT 134.400 160.050 135.450 163.950 ;
        RECT 133.950 157.950 136.050 160.050 ;
        RECT 140.400 145.050 141.450 193.950 ;
        RECT 143.400 190.050 144.450 193.950 ;
        RECT 146.400 193.050 147.450 196.950 ;
        RECT 148.950 193.950 151.050 196.050 ;
        RECT 151.950 193.950 154.050 196.050 ;
        RECT 155.250 194.850 156.750 195.750 ;
        RECT 157.950 193.950 160.050 196.050 ;
        RECT 160.950 193.950 163.050 196.050 ;
        RECT 145.950 190.950 148.050 193.050 ;
        RECT 158.400 190.050 159.450 193.950 ;
        RECT 161.400 193.050 162.450 193.950 ;
        RECT 160.950 190.950 163.050 193.050 ;
        RECT 142.950 187.950 145.050 190.050 ;
        RECT 157.950 187.950 160.050 190.050 ;
        RECT 154.950 184.950 157.050 187.050 ;
        RECT 151.950 175.950 154.050 178.050 ;
        RECT 145.950 172.950 148.050 175.050 ;
        RECT 146.400 166.050 147.450 172.950 ;
        RECT 152.400 166.050 153.450 175.950 ;
        RECT 142.950 164.250 144.750 165.150 ;
        RECT 145.950 163.950 148.050 166.050 ;
        RECT 149.250 164.250 151.050 165.150 ;
        RECT 151.950 163.950 154.050 166.050 ;
        RECT 142.950 160.950 145.050 163.050 ;
        RECT 146.250 161.850 147.750 162.750 ;
        RECT 148.950 160.950 151.050 163.050 ;
        RECT 143.400 157.050 144.450 160.950 ;
        RECT 149.400 160.050 150.450 160.950 ;
        RECT 155.400 160.050 156.450 184.950 ;
        RECT 160.950 178.950 163.050 181.050 ;
        RECT 161.400 172.050 162.450 178.950 ;
        RECT 160.950 169.950 163.050 172.050 ;
        RECT 163.950 171.450 166.050 172.050 ;
        RECT 167.400 171.450 168.450 199.950 ;
        RECT 188.400 199.050 189.450 199.950 ;
        RECT 169.950 197.250 172.050 198.150 ;
        RECT 175.950 197.250 178.050 198.150 ;
        RECT 178.950 197.250 180.750 198.150 ;
        RECT 181.950 196.950 184.050 199.050 ;
        RECT 185.250 197.250 186.750 198.150 ;
        RECT 187.950 196.950 190.050 199.050 ;
        RECT 191.250 197.250 193.050 198.150 ;
        RECT 169.950 193.950 172.050 196.050 ;
        RECT 175.950 195.450 178.050 196.050 ;
        RECT 178.950 195.450 181.050 196.050 ;
        RECT 173.250 194.250 174.750 195.150 ;
        RECT 175.950 194.400 181.050 195.450 ;
        RECT 182.250 194.850 183.750 195.750 ;
        RECT 175.950 193.950 178.050 194.400 ;
        RECT 178.950 193.950 181.050 194.400 ;
        RECT 184.950 193.950 187.050 196.050 ;
        RECT 188.250 194.850 189.750 195.750 ;
        RECT 190.950 193.950 193.050 196.050 ;
        RECT 172.950 190.950 175.050 193.050 ;
        RECT 175.950 190.950 178.050 193.050 ;
        RECT 173.400 183.450 174.450 190.950 ;
        RECT 170.400 182.400 174.450 183.450 ;
        RECT 170.400 178.050 171.450 182.400 ;
        RECT 172.950 178.950 175.050 181.050 ;
        RECT 169.950 175.950 172.050 178.050 ;
        RECT 163.950 170.400 168.450 171.450 ;
        RECT 163.950 169.950 166.050 170.400 ;
        RECT 164.400 169.050 165.450 169.950 ;
        RECT 157.950 167.250 160.050 168.150 ;
        RECT 160.950 167.850 163.050 168.750 ;
        RECT 163.950 166.950 166.050 169.050 ;
        RECT 167.250 167.250 168.750 168.150 ;
        RECT 169.950 166.950 172.050 169.050 ;
        RECT 173.400 166.050 174.450 178.950 ;
        RECT 157.950 163.950 160.050 166.050 ;
        RECT 163.950 164.850 165.750 165.750 ;
        RECT 166.950 163.950 169.050 166.050 ;
        RECT 170.250 164.850 171.750 165.750 ;
        RECT 172.950 163.950 175.050 166.050 ;
        RECT 158.400 163.050 159.450 163.950 ;
        RECT 176.400 163.050 177.450 190.950 ;
        RECT 179.400 187.050 180.450 193.950 ;
        RECT 181.950 187.950 184.050 190.050 ;
        RECT 178.950 184.950 181.050 187.050 ;
        RECT 178.950 175.950 181.050 178.050 ;
        RECT 157.950 160.950 160.050 163.050 ;
        RECT 169.950 160.950 172.050 163.050 ;
        RECT 172.950 161.850 175.050 162.750 ;
        RECT 175.950 160.950 178.050 163.050 ;
        RECT 148.950 157.950 151.050 160.050 ;
        RECT 154.950 157.950 157.050 160.050 ;
        RECT 142.950 154.950 145.050 157.050 ;
        RECT 139.950 142.950 142.050 145.050 ;
        RECT 139.950 139.950 142.050 142.050 ;
        RECT 115.950 130.950 118.050 133.050 ;
        RECT 121.950 130.950 124.050 133.050 ;
        RECT 116.400 130.050 117.450 130.950 ;
        RECT 109.950 129.450 112.050 130.050 ;
        RECT 104.250 128.250 106.050 129.150 ;
        RECT 107.400 128.400 112.050 129.450 ;
        RECT 94.950 125.850 96.750 126.750 ;
        RECT 97.950 124.950 100.050 127.050 ;
        RECT 103.950 126.450 106.050 127.050 ;
        RECT 107.400 126.450 108.450 128.400 ;
        RECT 109.950 127.950 112.050 128.400 ;
        RECT 113.250 128.250 114.750 129.150 ;
        RECT 115.950 127.950 118.050 130.050 ;
        RECT 121.950 129.450 124.050 130.050 ;
        RECT 119.400 128.400 124.050 129.450 ;
        RECT 103.950 125.400 108.450 126.450 ;
        RECT 109.950 125.850 111.750 126.750 ;
        RECT 103.950 124.950 106.050 125.400 ;
        RECT 112.950 124.950 115.050 127.050 ;
        RECT 116.250 125.850 118.050 126.750 ;
        RECT 98.400 115.050 99.450 124.950 ;
        RECT 97.950 112.950 100.050 115.050 ;
        RECT 113.400 103.050 114.450 124.950 ;
        RECT 119.400 115.050 120.450 128.400 ;
        RECT 121.950 127.950 124.050 128.400 ;
        RECT 125.250 128.250 126.750 129.150 ;
        RECT 127.950 127.950 130.050 130.050 ;
        RECT 136.950 127.950 139.050 130.050 ;
        RECT 137.400 127.050 138.450 127.950 ;
        RECT 121.950 125.850 123.750 126.750 ;
        RECT 124.950 124.950 127.050 127.050 ;
        RECT 128.250 125.850 130.050 126.750 ;
        RECT 133.950 125.250 135.750 126.150 ;
        RECT 136.950 124.950 139.050 127.050 ;
        RECT 118.950 112.950 121.050 115.050 ;
        RECT 112.950 100.950 115.050 103.050 ;
        RECT 125.400 100.050 126.450 124.950 ;
        RECT 133.950 121.950 136.050 124.050 ;
        RECT 137.250 122.850 139.050 123.750 ;
        RECT 140.400 121.050 141.450 139.950 ;
        RECT 143.400 130.050 144.450 154.950 ;
        RECT 148.950 136.950 151.050 139.050 ;
        RECT 149.400 130.050 150.450 136.950 ;
        RECT 142.950 127.950 145.050 130.050 ;
        RECT 146.250 128.250 147.750 129.150 ;
        RECT 148.950 127.950 151.050 130.050 ;
        RECT 157.950 129.450 160.050 130.050 ;
        RECT 155.400 128.400 160.050 129.450 ;
        RECT 163.950 129.450 166.050 130.050 ;
        RECT 142.950 125.850 144.750 126.750 ;
        RECT 145.950 124.950 148.050 127.050 ;
        RECT 149.250 125.850 151.050 126.750 ;
        RECT 139.950 118.950 142.050 121.050 ;
        RECT 146.400 105.450 147.450 124.950 ;
        RECT 148.950 112.950 151.050 115.050 ;
        RECT 143.400 104.400 147.450 105.450 ;
        RECT 109.950 97.950 112.050 100.050 ;
        RECT 115.950 97.950 118.050 100.050 ;
        RECT 124.950 97.950 127.050 100.050 ;
        RECT 130.950 97.950 133.050 100.050 ;
        RECT 100.950 94.950 103.050 97.050 ;
        RECT 104.250 95.250 105.750 96.150 ;
        RECT 106.950 94.950 109.050 97.050 ;
        RECT 109.950 95.850 112.050 96.750 ;
        RECT 112.950 95.250 115.050 96.150 ;
        RECT 91.950 91.950 94.050 94.050 ;
        RECT 97.950 91.950 100.050 94.050 ;
        RECT 101.250 92.850 102.750 93.750 ;
        RECT 103.950 91.950 106.050 94.050 ;
        RECT 107.250 92.850 109.050 93.750 ;
        RECT 112.950 93.450 115.050 94.050 ;
        RECT 110.400 92.400 115.050 93.450 ;
        RECT 88.950 85.950 91.050 88.050 ;
        RECT 85.950 70.950 88.050 73.050 ;
        RECT 82.950 64.950 85.050 67.050 ;
        RECT 46.950 58.950 49.050 61.050 ;
        RECT 52.950 58.950 55.050 61.050 ;
        RECT 58.950 58.950 61.050 61.050 ;
        RECT 70.950 59.250 73.050 60.150 ;
        RECT 53.400 58.050 54.450 58.950 ;
        RECT 46.950 57.450 49.050 58.050 ;
        RECT 44.400 56.400 49.050 57.450 ;
        RECT 46.950 55.950 49.050 56.400 ;
        RECT 50.250 56.250 51.750 57.150 ;
        RECT 52.950 55.950 55.050 58.050 ;
        RECT 16.950 53.850 18.750 54.750 ;
        RECT 19.950 52.950 22.050 55.050 ;
        RECT 25.950 52.950 28.050 55.050 ;
        RECT 28.950 53.250 30.750 54.150 ;
        RECT 31.950 52.950 34.050 55.050 ;
        RECT 35.250 53.250 36.750 54.150 ;
        RECT 37.950 52.950 40.050 55.050 ;
        RECT 20.400 52.050 21.450 52.950 ;
        RECT 41.400 52.050 42.450 55.950 ;
        RECT 46.950 53.850 48.750 54.750 ;
        RECT 49.950 52.950 52.050 55.050 ;
        RECT 53.250 53.850 55.050 54.750 ;
        RECT 19.950 49.950 22.050 52.050 ;
        RECT 25.950 49.950 28.050 52.050 ;
        RECT 28.950 49.950 31.050 52.050 ;
        RECT 32.250 50.850 33.750 51.750 ;
        RECT 34.950 49.950 37.050 52.050 ;
        RECT 40.950 49.950 43.050 52.050 ;
        RECT 16.950 37.950 19.050 40.050 ;
        RECT 4.950 22.950 7.050 25.050 ;
        RECT 8.250 23.850 9.750 24.750 ;
        RECT 10.950 22.950 13.050 25.050 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 4.950 20.850 7.050 21.750 ;
        RECT 10.950 20.850 13.050 21.750 ;
        RECT 13.950 20.850 16.050 21.750 ;
        RECT 17.400 18.450 18.450 37.950 ;
        RECT 26.400 28.050 27.450 49.950 ;
        RECT 29.400 49.050 30.450 49.950 ;
        RECT 28.950 46.950 31.050 49.050 ;
        RECT 40.950 46.950 43.050 49.050 ;
        RECT 25.950 25.950 28.050 28.050 ;
        RECT 31.950 25.950 34.050 28.050 ;
        RECT 32.400 25.050 33.450 25.950 ;
        RECT 22.950 22.950 25.050 25.050 ;
        RECT 31.950 22.950 34.050 25.050 ;
        RECT 35.250 23.250 36.750 24.150 ;
        RECT 37.950 22.950 40.050 25.050 ;
        RECT 41.400 22.050 42.450 46.950 ;
        RECT 50.400 46.050 51.450 52.950 ;
        RECT 59.400 52.050 60.450 58.950 ;
        RECT 67.950 56.250 69.750 57.150 ;
        RECT 70.950 55.950 73.050 58.050 ;
        RECT 76.950 57.450 79.050 58.050 ;
        RECT 74.250 56.250 75.750 57.150 ;
        RECT 76.950 56.400 81.450 57.450 ;
        RECT 76.950 55.950 79.050 56.400 ;
        RECT 61.950 52.950 64.050 55.050 ;
        RECT 67.950 52.950 70.050 55.050 ;
        RECT 58.950 49.950 61.050 52.050 ;
        RECT 61.950 50.850 64.050 51.750 ;
        RECT 64.950 50.250 67.050 51.150 ;
        RECT 49.950 43.950 52.050 46.050 ;
        RECT 59.400 40.050 60.450 49.950 ;
        RECT 64.950 46.950 67.050 49.050 ;
        RECT 71.400 46.050 72.450 55.950 ;
        RECT 73.950 52.950 76.050 55.050 ;
        RECT 77.250 53.850 79.050 54.750 ;
        RECT 70.950 43.950 73.050 46.050 ;
        RECT 67.950 40.950 70.050 43.050 ;
        RECT 58.950 37.950 61.050 40.050 ;
        RECT 58.950 34.950 61.050 37.050 ;
        RECT 49.950 25.950 52.050 28.050 ;
        RECT 50.400 25.050 51.450 25.950 ;
        RECT 59.400 25.050 60.450 34.950 ;
        RECT 49.950 22.950 52.050 25.050 ;
        RECT 55.950 22.950 58.050 25.050 ;
        RECT 58.950 24.450 61.050 25.050 ;
        RECT 58.950 23.400 63.450 24.450 ;
        RECT 58.950 22.950 61.050 23.400 ;
        RECT 19.950 20.250 22.050 21.150 ;
        RECT 22.950 20.850 25.050 21.750 ;
        RECT 31.950 20.850 33.750 21.750 ;
        RECT 34.950 19.950 37.050 22.050 ;
        RECT 38.250 20.850 39.750 21.750 ;
        RECT 40.950 19.950 43.050 22.050 ;
        RECT 49.950 20.850 52.050 21.750 ;
        RECT 52.950 20.250 55.050 21.150 ;
        RECT 56.400 19.050 57.450 22.950 ;
        RECT 58.950 20.850 61.050 21.750 ;
        RECT 19.950 18.450 22.050 19.050 ;
        RECT 17.400 17.400 22.050 18.450 ;
        RECT 40.950 17.850 43.050 18.750 ;
        RECT 52.950 18.450 55.050 19.050 ;
        RECT 55.950 18.450 58.050 19.050 ;
        RECT 19.950 16.950 22.050 17.400 ;
        RECT 52.950 17.400 58.050 18.450 ;
        RECT 62.400 18.450 63.450 23.400 ;
        RECT 68.400 22.050 69.450 40.950 ;
        RECT 80.400 37.050 81.450 56.400 ;
        RECT 83.400 49.050 84.450 64.950 ;
        RECT 88.950 52.950 91.050 55.050 ;
        RECT 88.950 50.850 91.050 51.750 ;
        RECT 82.950 46.950 85.050 49.050 ;
        RECT 73.950 34.950 76.050 37.050 ;
        RECT 79.950 34.950 82.050 37.050 ;
        RECT 74.400 25.050 75.450 34.950 ;
        RECT 79.950 31.950 82.050 34.050 ;
        RECT 80.400 25.050 81.450 31.950 ;
        RECT 92.400 25.050 93.450 91.950 ;
        RECT 104.400 91.050 105.450 91.950 ;
        RECT 110.400 91.050 111.450 92.400 ;
        RECT 112.950 91.950 115.050 92.400 ;
        RECT 116.400 91.050 117.450 97.950 ;
        RECT 124.950 96.450 127.050 97.050 ;
        RECT 122.400 95.400 127.050 96.450 ;
        RECT 97.950 89.850 100.050 90.750 ;
        RECT 103.950 88.950 106.050 91.050 ;
        RECT 109.950 88.950 112.050 91.050 ;
        RECT 112.950 88.950 115.050 91.050 ;
        RECT 115.950 88.950 118.050 91.050 ;
        RECT 103.950 76.950 106.050 79.050 ;
        RECT 104.400 55.050 105.450 76.950 ;
        RECT 106.950 67.950 109.050 70.050 ;
        RECT 107.400 55.050 108.450 67.950 ;
        RECT 110.400 58.050 111.450 88.950 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 94.950 53.250 97.050 54.150 ;
        RECT 100.950 52.950 103.050 55.050 ;
        RECT 103.950 52.950 106.050 55.050 ;
        RECT 106.950 52.950 109.050 55.050 ;
        RECT 110.250 53.250 112.050 54.150 ;
        RECT 94.950 49.950 97.050 52.050 ;
        RECT 98.250 50.250 100.050 51.150 ;
        RECT 100.950 50.850 103.050 51.750 ;
        RECT 103.950 50.250 106.050 51.150 ;
        RECT 106.950 50.850 108.750 51.750 ;
        RECT 109.950 49.950 112.050 52.050 ;
        RECT 113.400 49.050 114.450 88.950 ;
        RECT 122.400 79.050 123.450 95.400 ;
        RECT 124.950 94.950 127.050 95.400 ;
        RECT 128.250 95.250 130.050 96.150 ;
        RECT 130.950 95.850 133.050 96.750 ;
        RECT 133.950 95.250 136.050 96.150 ;
        RECT 139.950 95.250 142.050 96.150 ;
        RECT 124.950 92.850 126.750 93.750 ;
        RECT 127.950 91.950 130.050 94.050 ;
        RECT 133.950 91.950 136.050 94.050 ;
        RECT 139.950 91.950 142.050 94.050 ;
        RECT 121.950 76.950 124.050 79.050 ;
        RECT 118.950 55.950 121.050 58.050 ;
        RECT 124.950 56.250 127.050 57.150 ;
        RECT 119.400 55.050 120.450 55.950 ;
        RECT 115.950 53.250 117.750 54.150 ;
        RECT 118.950 52.950 121.050 55.050 ;
        RECT 124.950 54.450 127.050 55.050 ;
        RECT 128.400 54.450 129.450 91.950 ;
        RECT 133.950 70.950 136.050 73.050 ;
        RECT 130.950 61.950 133.050 64.050 ;
        RECT 122.250 53.250 123.750 54.150 ;
        RECT 124.950 53.400 129.450 54.450 ;
        RECT 124.950 52.950 127.050 53.400 ;
        RECT 115.950 49.950 118.050 52.050 ;
        RECT 119.250 50.850 120.750 51.750 ;
        RECT 121.950 49.950 124.050 52.050 ;
        RECT 97.950 46.950 100.050 49.050 ;
        RECT 100.950 46.950 103.050 49.050 ;
        RECT 103.950 46.950 106.050 49.050 ;
        RECT 112.950 46.950 115.050 49.050 ;
        RECT 98.400 46.050 99.450 46.950 ;
        RECT 97.950 43.950 100.050 46.050 ;
        RECT 101.400 28.050 102.450 46.950 ;
        RECT 97.950 25.950 100.050 28.050 ;
        RECT 100.950 25.950 103.050 28.050 ;
        RECT 73.950 22.950 76.050 25.050 ;
        RECT 77.250 23.250 78.750 24.150 ;
        RECT 79.950 22.950 82.050 25.050 ;
        RECT 83.250 23.250 84.750 24.150 ;
        RECT 85.950 22.950 88.050 25.050 ;
        RECT 91.950 22.950 94.050 25.050 ;
        RECT 92.400 22.050 93.450 22.950 ;
        RECT 98.400 22.050 99.450 25.950 ;
        RECT 104.400 22.050 105.450 46.950 ;
        RECT 122.400 28.050 123.450 49.950 ;
        RECT 125.400 43.050 126.450 52.950 ;
        RECT 131.400 46.050 132.450 61.950 ;
        RECT 134.400 58.050 135.450 70.950 ;
        RECT 143.400 67.050 144.450 104.400 ;
        RECT 145.950 100.950 148.050 103.050 ;
        RECT 146.400 100.050 147.450 100.950 ;
        RECT 149.400 100.050 150.450 112.950 ;
        RECT 155.400 103.050 156.450 128.400 ;
        RECT 157.950 127.950 160.050 128.400 ;
        RECT 161.250 128.250 162.750 129.150 ;
        RECT 163.950 128.400 168.450 129.450 ;
        RECT 163.950 127.950 166.050 128.400 ;
        RECT 157.950 125.850 159.750 126.750 ;
        RECT 160.950 124.950 163.050 127.050 ;
        RECT 164.250 125.850 166.050 126.750 ;
        RECT 161.400 115.050 162.450 124.950 ;
        RECT 167.400 121.050 168.450 128.400 ;
        RECT 166.950 118.950 169.050 121.050 ;
        RECT 160.950 112.950 163.050 115.050 ;
        RECT 154.950 100.950 157.050 103.050 ;
        RECT 160.950 100.950 163.050 103.050 ;
        RECT 161.400 100.050 162.450 100.950 ;
        RECT 145.950 97.950 148.050 100.050 ;
        RECT 148.950 97.950 151.050 100.050 ;
        RECT 160.950 97.950 163.050 100.050 ;
        RECT 146.400 97.050 147.450 97.950 ;
        RECT 145.950 94.950 148.050 97.050 ;
        RECT 149.250 95.850 151.050 96.750 ;
        RECT 154.950 96.450 157.050 97.050 ;
        RECT 152.400 95.400 157.050 96.450 ;
        RECT 145.950 92.850 148.050 93.750 ;
        RECT 152.400 70.050 153.450 95.400 ;
        RECT 154.950 94.950 157.050 95.400 ;
        RECT 158.250 95.250 160.050 96.150 ;
        RECT 160.950 95.850 163.050 96.750 ;
        RECT 163.950 95.250 166.050 96.150 ;
        RECT 167.400 94.050 168.450 118.950 ;
        RECT 154.950 92.850 156.750 93.750 ;
        RECT 157.950 91.950 160.050 94.050 ;
        RECT 163.950 93.450 166.050 94.050 ;
        RECT 166.950 93.450 169.050 94.050 ;
        RECT 163.950 92.400 169.050 93.450 ;
        RECT 163.950 91.950 166.050 92.400 ;
        RECT 166.950 91.950 169.050 92.400 ;
        RECT 163.950 85.950 166.050 88.050 ;
        RECT 160.950 76.950 163.050 79.050 ;
        RECT 151.950 67.950 154.050 70.050 ;
        RECT 142.950 64.950 145.050 67.050 ;
        RECT 151.950 64.950 154.050 67.050 ;
        RECT 139.950 58.950 142.050 61.050 ;
        RECT 145.950 59.250 148.050 60.150 ;
        RECT 140.400 58.050 141.450 58.950 ;
        RECT 152.400 58.050 153.450 64.950 ;
        RECT 133.950 55.950 136.050 58.050 ;
        RECT 137.250 56.250 138.750 57.150 ;
        RECT 139.950 55.950 142.050 58.050 ;
        RECT 142.950 56.250 144.750 57.150 ;
        RECT 145.950 55.950 148.050 58.050 ;
        RECT 149.250 56.250 150.750 57.150 ;
        RECT 151.950 55.950 154.050 58.050 ;
        RECT 133.950 53.850 135.750 54.750 ;
        RECT 136.950 52.950 139.050 55.050 ;
        RECT 140.250 53.850 142.050 54.750 ;
        RECT 142.950 52.950 145.050 55.050 ;
        RECT 148.950 52.950 151.050 55.050 ;
        RECT 152.250 53.850 154.050 54.750 ;
        RECT 137.400 52.050 138.450 52.950 ;
        RECT 136.950 49.950 139.050 52.050 ;
        RECT 149.400 49.050 150.450 52.950 ;
        RECT 142.950 46.950 145.050 49.050 ;
        RECT 148.950 46.950 151.050 49.050 ;
        RECT 130.950 43.950 133.050 46.050 ;
        RECT 124.950 40.950 127.050 43.050 ;
        RECT 139.950 40.950 142.050 43.050 ;
        RECT 115.950 25.950 118.050 28.050 ;
        RECT 121.950 25.950 124.050 28.050 ;
        RECT 109.950 24.450 112.050 25.050 ;
        RECT 107.400 23.400 112.050 24.450 ;
        RECT 64.950 20.250 66.750 21.150 ;
        RECT 67.950 19.950 70.050 22.050 ;
        RECT 71.250 20.250 73.050 21.150 ;
        RECT 73.950 20.850 75.750 21.750 ;
        RECT 76.950 19.950 79.050 22.050 ;
        RECT 80.250 20.850 81.750 21.750 ;
        RECT 82.950 19.950 85.050 22.050 ;
        RECT 86.250 20.850 88.050 21.750 ;
        RECT 91.950 19.950 94.050 22.050 ;
        RECT 94.950 19.950 97.050 22.050 ;
        RECT 97.950 19.950 100.050 22.050 ;
        RECT 101.250 20.250 103.050 21.150 ;
        RECT 103.950 19.950 106.050 22.050 ;
        RECT 77.400 19.050 78.450 19.950 ;
        RECT 95.400 19.050 96.450 19.950 ;
        RECT 64.950 18.450 67.050 19.050 ;
        RECT 62.400 17.400 67.050 18.450 ;
        RECT 68.250 17.850 69.750 18.750 ;
        RECT 52.950 16.950 55.050 17.400 ;
        RECT 55.950 16.950 58.050 17.400 ;
        RECT 64.950 16.950 67.050 17.400 ;
        RECT 70.950 16.950 73.050 19.050 ;
        RECT 76.950 16.950 79.050 19.050 ;
        RECT 91.950 17.850 93.750 18.750 ;
        RECT 94.950 16.950 97.050 19.050 ;
        RECT 98.250 17.850 99.750 18.750 ;
        RECT 100.950 16.950 103.050 19.050 ;
        RECT 94.950 14.850 97.050 15.750 ;
        RECT 107.400 13.050 108.450 23.400 ;
        RECT 109.950 22.950 112.050 23.400 ;
        RECT 113.250 23.250 115.050 24.150 ;
        RECT 115.950 23.850 118.050 24.750 ;
        RECT 118.950 23.250 121.050 24.150 ;
        RECT 122.400 22.050 123.450 25.950 ;
        RECT 127.950 22.950 130.050 25.050 ;
        RECT 128.400 22.050 129.450 22.950 ;
        RECT 140.400 22.050 141.450 40.950 ;
        RECT 143.400 25.050 144.450 46.950 ;
        RECT 157.950 34.950 160.050 37.050 ;
        RECT 151.950 31.950 154.050 34.050 ;
        RECT 148.950 28.950 151.050 31.050 ;
        RECT 149.400 25.050 150.450 28.950 ;
        RECT 152.400 25.050 153.450 31.950 ;
        RECT 158.400 25.050 159.450 34.950 ;
        RECT 161.400 27.450 162.450 76.950 ;
        RECT 164.400 58.050 165.450 85.950 ;
        RECT 170.400 67.050 171.450 160.950 ;
        RECT 179.400 160.050 180.450 175.950 ;
        RECT 182.400 175.050 183.450 187.950 ;
        RECT 185.400 184.050 186.450 193.950 ;
        RECT 191.400 193.050 192.450 193.950 ;
        RECT 187.950 190.950 190.050 193.050 ;
        RECT 190.950 190.950 193.050 193.050 ;
        RECT 184.950 181.950 187.050 184.050 ;
        RECT 188.400 181.050 189.450 190.950 ;
        RECT 190.950 181.950 193.050 184.050 ;
        RECT 187.950 178.950 190.050 181.050 ;
        RECT 181.950 172.950 184.050 175.050 ;
        RECT 181.950 169.950 184.050 172.050 ;
        RECT 182.400 166.050 183.450 169.950 ;
        RECT 191.400 169.050 192.450 181.950 ;
        RECT 194.400 178.050 195.450 217.950 ;
        RECT 203.400 202.050 204.450 229.950 ;
        RECT 205.950 226.950 208.050 229.050 ;
        RECT 208.950 226.950 211.050 229.050 ;
        RECT 196.950 199.950 199.050 202.050 ;
        RECT 200.250 200.250 201.750 201.150 ;
        RECT 202.950 199.950 205.050 202.050 ;
        RECT 196.950 197.850 198.750 198.750 ;
        RECT 199.950 196.950 202.050 199.050 ;
        RECT 203.250 197.850 205.050 198.750 ;
        RECT 206.400 195.450 207.450 226.950 ;
        RECT 209.400 202.050 210.450 226.950 ;
        RECT 212.400 211.050 213.450 235.950 ;
        RECT 218.400 220.050 219.450 274.950 ;
        RECT 221.400 274.050 222.450 277.950 ;
        RECT 233.400 274.050 234.450 280.950 ;
        RECT 238.950 274.950 241.050 277.050 ;
        RECT 239.400 274.050 240.450 274.950 ;
        RECT 220.950 271.950 223.050 274.050 ;
        RECT 226.950 273.450 229.050 274.050 ;
        RECT 224.250 272.250 225.750 273.150 ;
        RECT 226.950 272.400 231.450 273.450 ;
        RECT 226.950 271.950 229.050 272.400 ;
        RECT 220.950 269.850 222.750 270.750 ;
        RECT 223.950 268.950 226.050 271.050 ;
        RECT 227.250 269.850 229.050 270.750 ;
        RECT 224.400 259.050 225.450 268.950 ;
        RECT 230.400 268.050 231.450 272.400 ;
        RECT 232.950 271.950 235.050 274.050 ;
        RECT 236.250 272.250 237.750 273.150 ;
        RECT 238.950 271.950 241.050 274.050 ;
        RECT 232.950 269.850 234.750 270.750 ;
        RECT 235.950 268.950 238.050 271.050 ;
        RECT 239.250 269.850 241.050 270.750 ;
        RECT 226.950 265.950 229.050 268.050 ;
        RECT 229.950 265.950 232.050 268.050 ;
        RECT 227.400 259.050 228.450 265.950 ;
        RECT 223.950 256.950 226.050 259.050 ;
        RECT 226.950 256.950 229.050 259.050 ;
        RECT 242.400 256.050 243.450 298.950 ;
        RECT 251.400 280.050 252.450 328.950 ;
        RECT 254.400 316.050 255.450 409.950 ;
        RECT 257.400 382.050 258.450 412.950 ;
        RECT 265.950 409.950 268.050 412.050 ;
        RECT 269.250 410.850 270.750 411.750 ;
        RECT 271.950 409.950 274.050 412.050 ;
        RECT 266.400 409.050 267.450 409.950 ;
        RECT 265.950 406.950 268.050 409.050 ;
        RECT 265.950 403.950 268.050 406.050 ;
        RECT 266.400 385.050 267.450 403.950 ;
        RECT 275.400 400.050 276.450 412.950 ;
        RECT 278.400 409.050 279.450 427.950 ;
        RECT 284.400 421.050 285.450 439.950 ;
        RECT 286.950 430.950 289.050 433.050 ;
        RECT 283.950 418.950 286.050 421.050 ;
        RECT 287.400 415.050 288.450 430.950 ;
        RECT 293.400 418.050 294.450 451.950 ;
        RECT 295.950 448.950 298.050 451.050 ;
        RECT 299.250 449.850 300.750 450.750 ;
        RECT 301.950 448.950 304.050 451.050 ;
        RECT 296.400 445.050 297.450 448.950 ;
        RECT 302.400 445.050 303.450 448.950 ;
        RECT 307.950 445.950 310.050 448.050 ;
        RECT 295.950 442.950 298.050 445.050 ;
        RECT 301.950 442.950 304.050 445.050 ;
        RECT 302.400 430.050 303.450 442.950 ;
        RECT 308.400 430.050 309.450 445.950 ;
        RECT 301.950 427.950 304.050 430.050 ;
        RECT 307.950 427.950 310.050 430.050 ;
        RECT 307.950 424.950 310.050 427.050 ;
        RECT 298.950 421.950 301.050 424.050 ;
        RECT 292.950 415.950 295.050 418.050 ;
        RECT 283.950 413.250 285.750 414.150 ;
        RECT 286.950 412.950 289.050 415.050 ;
        RECT 292.950 412.950 295.050 415.050 ;
        RECT 283.950 409.950 286.050 412.050 ;
        RECT 287.250 410.850 289.050 411.750 ;
        RECT 289.950 410.250 292.050 411.150 ;
        RECT 292.950 410.850 295.050 411.750 ;
        RECT 295.950 409.950 298.050 412.050 ;
        RECT 277.950 406.950 280.050 409.050 ;
        RECT 278.400 406.050 279.450 406.950 ;
        RECT 277.950 403.950 280.050 406.050 ;
        RECT 274.950 397.950 277.050 400.050 ;
        RECT 271.950 391.950 274.050 394.050 ;
        RECT 277.950 391.950 280.050 394.050 ;
        RECT 272.400 385.050 273.450 391.950 ;
        RECT 278.400 385.050 279.450 391.950 ;
        RECT 284.400 388.050 285.450 409.950 ;
        RECT 289.950 406.950 292.050 409.050 ;
        RECT 290.400 405.450 291.450 406.950 ;
        RECT 296.400 406.050 297.450 409.950 ;
        RECT 287.400 404.400 291.450 405.450 ;
        RECT 287.400 388.050 288.450 404.400 ;
        RECT 295.950 403.950 298.050 406.050 ;
        RECT 299.400 403.050 300.450 421.950 ;
        RECT 301.950 416.250 304.050 417.150 ;
        RECT 308.400 415.050 309.450 424.950 ;
        RECT 301.950 412.950 304.050 415.050 ;
        RECT 305.250 413.250 306.750 414.150 ;
        RECT 307.950 412.950 310.050 415.050 ;
        RECT 311.250 413.250 313.050 414.150 ;
        RECT 304.950 409.950 307.050 412.050 ;
        RECT 308.250 410.850 309.750 411.750 ;
        RECT 310.950 409.950 313.050 412.050 ;
        RECT 311.400 409.050 312.450 409.950 ;
        RECT 310.950 406.950 313.050 409.050 ;
        RECT 298.950 400.950 301.050 403.050 ;
        RECT 307.950 400.950 310.050 403.050 ;
        RECT 304.950 389.400 307.050 391.500 ;
        RECT 283.950 385.950 286.050 388.050 ;
        RECT 286.950 385.950 289.050 388.050 ;
        RECT 295.950 387.450 298.050 388.050 ;
        RECT 290.400 386.400 298.050 387.450 ;
        RECT 259.950 382.950 262.050 385.050 ;
        RECT 263.250 383.250 264.750 384.150 ;
        RECT 265.950 382.950 268.050 385.050 ;
        RECT 271.950 382.950 274.050 385.050 ;
        RECT 275.250 383.250 276.750 384.150 ;
        RECT 277.950 382.950 280.050 385.050 ;
        RECT 281.250 383.250 282.750 384.150 ;
        RECT 283.950 382.950 286.050 385.050 ;
        RECT 256.950 379.950 259.050 382.050 ;
        RECT 260.250 380.850 261.750 381.750 ;
        RECT 262.950 379.950 265.050 382.050 ;
        RECT 266.250 380.850 268.050 381.750 ;
        RECT 271.950 380.850 273.750 381.750 ;
        RECT 274.950 379.950 277.050 382.050 ;
        RECT 278.250 380.850 279.750 381.750 ;
        RECT 280.950 379.950 283.050 382.050 ;
        RECT 284.250 380.850 286.050 381.750 ;
        RECT 256.950 377.850 259.050 378.750 ;
        RECT 256.950 370.950 259.050 373.050 ;
        RECT 257.400 331.050 258.450 370.950 ;
        RECT 263.400 370.050 264.450 379.950 ;
        RECT 281.400 373.050 282.450 379.950 ;
        RECT 287.400 379.050 288.450 385.950 ;
        RECT 290.400 385.050 291.450 386.400 ;
        RECT 295.950 385.950 298.050 386.400 ;
        RECT 289.950 382.950 292.050 385.050 ;
        RECT 292.950 383.250 295.050 384.150 ;
        RECT 295.950 383.850 298.050 384.750 ;
        RECT 301.950 382.950 304.050 385.050 ;
        RECT 292.950 379.950 295.050 382.050 ;
        RECT 286.950 376.950 289.050 379.050 ;
        RECT 280.950 370.950 283.050 373.050 ;
        RECT 262.950 367.950 265.050 370.050 ;
        RECT 281.400 367.050 282.450 370.950 ;
        RECT 280.950 364.950 283.050 367.050 ;
        RECT 286.950 364.950 289.050 367.050 ;
        RECT 259.950 350.400 262.050 352.500 ;
        RECT 280.950 351.300 283.050 353.400 ;
        RECT 260.400 333.600 261.600 350.400 ;
        RECT 274.950 346.950 277.050 349.050 ;
        RECT 281.250 347.700 282.450 351.300 ;
        RECT 265.950 341.250 268.050 342.150 ;
        RECT 271.950 341.250 274.050 342.150 ;
        RECT 265.950 337.950 268.050 340.050 ;
        RECT 271.950 339.450 274.050 340.050 ;
        RECT 275.400 339.450 276.450 346.950 ;
        RECT 280.950 345.600 283.050 347.700 ;
        RECT 271.950 338.400 276.450 339.450 ;
        RECT 271.950 337.950 274.050 338.400 ;
        RECT 259.950 331.500 262.050 333.600 ;
        RECT 271.950 331.950 274.050 334.050 ;
        RECT 281.250 333.600 282.450 345.600 ;
        RECT 283.950 337.950 286.050 340.050 ;
        RECT 283.950 335.850 286.050 336.750 ;
        RECT 256.950 328.950 259.050 331.050 ;
        RECT 265.950 325.950 268.050 328.050 ;
        RECT 256.950 322.950 259.050 325.050 ;
        RECT 253.950 313.950 256.050 316.050 ;
        RECT 257.400 313.050 258.450 322.950 ;
        RECT 266.400 313.050 267.450 325.950 ;
        RECT 272.400 313.050 273.450 331.950 ;
        RECT 280.950 331.500 283.050 333.600 ;
        RECT 274.950 319.950 277.050 322.050 ;
        RECT 275.400 313.050 276.450 319.950 ;
        RECT 280.950 315.450 283.050 316.050 ;
        RECT 278.400 314.400 283.050 315.450 ;
        RECT 253.950 310.950 256.050 313.050 ;
        RECT 256.950 310.950 259.050 313.050 ;
        RECT 262.950 312.450 265.050 313.050 ;
        RECT 265.950 312.450 268.050 313.050 ;
        RECT 260.250 311.250 261.750 312.150 ;
        RECT 262.950 311.400 268.050 312.450 ;
        RECT 262.950 310.950 265.050 311.400 ;
        RECT 265.950 310.950 268.050 311.400 ;
        RECT 269.250 311.250 270.750 312.150 ;
        RECT 271.950 310.950 274.050 313.050 ;
        RECT 274.950 310.950 277.050 313.050 ;
        RECT 254.400 310.050 255.450 310.950 ;
        RECT 253.950 307.950 256.050 310.050 ;
        RECT 257.250 308.850 258.750 309.750 ;
        RECT 259.950 307.950 262.050 310.050 ;
        RECT 263.250 308.850 265.050 309.750 ;
        RECT 265.950 308.850 267.750 309.750 ;
        RECT 268.950 307.950 271.050 310.050 ;
        RECT 272.250 308.850 273.750 309.750 ;
        RECT 274.950 307.950 277.050 310.050 ;
        RECT 253.950 305.850 256.050 306.750 ;
        RECT 256.950 295.950 259.050 298.050 ;
        RECT 244.950 277.950 247.050 280.050 ;
        RECT 250.950 277.950 253.050 280.050 ;
        RECT 245.400 271.050 246.450 277.950 ;
        RECT 250.950 271.950 253.050 274.050 ;
        RECT 244.950 268.950 247.050 271.050 ;
        RECT 248.250 269.250 250.050 270.150 ;
        RECT 244.950 266.850 246.750 267.750 ;
        RECT 247.950 265.950 250.050 268.050 ;
        RECT 244.950 262.950 247.050 265.050 ;
        RECT 241.950 253.950 244.050 256.050 ;
        RECT 220.950 244.950 223.050 247.050 ;
        RECT 221.400 241.050 222.450 244.950 ;
        RECT 223.950 241.950 226.050 244.050 ;
        RECT 220.950 238.950 223.050 241.050 ;
        RECT 220.950 236.850 223.050 237.750 ;
        RECT 220.950 232.950 223.050 235.050 ;
        RECT 217.950 217.950 220.050 220.050 ;
        RECT 221.400 217.050 222.450 232.950 ;
        RECT 224.400 229.050 225.450 241.950 ;
        RECT 229.950 238.950 232.050 241.050 ;
        RECT 233.400 239.400 240.450 240.450 ;
        RECT 226.950 236.250 229.050 237.150 ;
        RECT 229.950 236.850 232.050 237.750 ;
        RECT 226.950 232.950 229.050 235.050 ;
        RECT 227.400 232.050 228.450 232.950 ;
        RECT 226.950 229.950 229.050 232.050 ;
        RECT 223.950 226.950 226.050 229.050 ;
        RECT 226.950 220.950 229.050 223.050 ;
        RECT 220.950 214.950 223.050 217.050 ;
        RECT 211.950 208.950 214.050 211.050 ;
        RECT 214.950 208.950 217.050 211.050 ;
        RECT 215.400 202.050 216.450 208.950 ;
        RECT 221.400 202.050 222.450 214.950 ;
        RECT 227.400 202.050 228.450 220.950 ;
        RECT 229.950 217.950 232.050 220.050 ;
        RECT 208.950 199.950 211.050 202.050 ;
        RECT 212.250 200.250 213.750 201.150 ;
        RECT 214.950 199.950 217.050 202.050 ;
        RECT 217.950 199.950 220.050 202.050 ;
        RECT 220.950 199.950 223.050 202.050 ;
        RECT 224.250 200.250 225.750 201.150 ;
        RECT 226.950 199.950 229.050 202.050 ;
        RECT 208.950 197.850 210.750 198.750 ;
        RECT 211.950 196.950 214.050 199.050 ;
        RECT 215.250 197.850 217.050 198.750 ;
        RECT 203.400 194.400 207.450 195.450 ;
        RECT 196.950 178.950 199.050 181.050 ;
        RECT 193.950 175.950 196.050 178.050 ;
        RECT 197.400 172.050 198.450 178.950 ;
        RECT 196.950 171.450 199.050 172.050 ;
        RECT 194.400 170.400 199.050 171.450 ;
        RECT 184.950 166.950 187.050 169.050 ;
        RECT 188.250 167.250 189.750 168.150 ;
        RECT 190.950 166.950 193.050 169.050 ;
        RECT 194.400 166.050 195.450 170.400 ;
        RECT 196.950 169.950 199.050 170.400 ;
        RECT 196.950 167.850 199.050 168.750 ;
        RECT 199.950 167.250 202.050 168.150 ;
        RECT 181.950 163.950 184.050 166.050 ;
        RECT 185.250 164.850 186.750 165.750 ;
        RECT 187.950 163.950 190.050 166.050 ;
        RECT 191.250 164.850 193.050 165.750 ;
        RECT 193.950 163.950 196.050 166.050 ;
        RECT 199.950 163.950 202.050 166.050 ;
        RECT 181.950 161.850 184.050 162.750 ;
        RECT 184.950 160.950 187.050 163.050 ;
        RECT 203.400 162.450 204.450 194.400 ;
        RECT 212.400 187.050 213.450 196.950 ;
        RECT 211.950 184.950 214.050 187.050 ;
        RECT 205.950 181.950 208.050 184.050 ;
        RECT 206.400 172.050 207.450 181.950 ;
        RECT 218.400 178.050 219.450 199.950 ;
        RECT 220.950 197.850 222.750 198.750 ;
        RECT 223.950 196.950 226.050 199.050 ;
        RECT 227.250 197.850 229.050 198.750 ;
        RECT 224.400 193.050 225.450 196.950 ;
        RECT 223.950 190.950 226.050 193.050 ;
        RECT 211.950 175.950 214.050 178.050 ;
        RECT 217.950 175.950 220.050 178.050 ;
        RECT 212.400 172.050 213.450 175.950 ;
        RECT 205.950 169.950 208.050 172.050 ;
        RECT 211.950 169.950 214.050 172.050 ;
        RECT 217.950 169.950 220.050 172.050 ;
        RECT 205.950 167.850 208.050 168.750 ;
        RECT 208.950 167.250 211.050 168.150 ;
        RECT 208.950 163.950 211.050 166.050 ;
        RECT 212.400 165.450 213.450 169.950 ;
        RECT 214.950 167.250 217.050 168.150 ;
        RECT 217.950 167.850 220.050 168.750 ;
        RECT 223.950 168.450 226.050 169.050 ;
        RECT 220.950 167.250 222.750 168.150 ;
        RECT 223.950 167.400 228.450 168.450 ;
        RECT 223.950 166.950 226.050 167.400 ;
        RECT 214.950 165.450 217.050 166.050 ;
        RECT 212.400 164.400 217.050 165.450 ;
        RECT 214.950 163.950 217.050 164.400 ;
        RECT 220.950 163.950 223.050 166.050 ;
        RECT 224.250 164.850 226.050 165.750 ;
        RECT 200.400 161.400 204.450 162.450 ;
        RECT 178.950 157.950 181.050 160.050 ;
        RECT 172.950 151.950 175.050 154.050 ;
        RECT 173.400 130.050 174.450 151.950 ;
        RECT 178.950 130.950 181.050 133.050 ;
        RECT 185.400 132.450 186.450 160.950 ;
        RECT 196.950 157.950 199.050 160.050 ;
        RECT 182.400 131.400 186.450 132.450 ;
        RECT 179.400 130.050 180.450 130.950 ;
        RECT 172.950 127.950 175.050 130.050 ;
        RECT 176.250 128.250 177.750 129.150 ;
        RECT 178.950 127.950 181.050 130.050 ;
        RECT 172.950 125.850 174.750 126.750 ;
        RECT 175.950 124.950 178.050 127.050 ;
        RECT 179.250 125.850 181.050 126.750 ;
        RECT 172.950 103.950 175.050 106.050 ;
        RECT 173.400 97.050 174.450 103.950 ;
        RECT 178.950 100.950 181.050 103.050 ;
        RECT 175.950 97.950 178.050 100.050 ;
        RECT 172.950 94.950 175.050 97.050 ;
        RECT 176.400 94.050 177.450 97.950 ;
        RECT 172.950 92.250 174.750 93.150 ;
        RECT 175.950 91.950 178.050 94.050 ;
        RECT 179.400 91.050 180.450 100.950 ;
        RECT 182.400 96.450 183.450 131.400 ;
        RECT 184.950 128.250 187.050 129.150 ;
        RECT 184.950 124.950 187.050 127.050 ;
        RECT 188.250 125.250 189.750 126.150 ;
        RECT 190.950 124.950 193.050 127.050 ;
        RECT 194.250 125.250 196.050 126.150 ;
        RECT 185.400 99.450 186.450 124.950 ;
        RECT 187.950 121.950 190.050 124.050 ;
        RECT 191.250 122.850 192.750 123.750 ;
        RECT 193.950 121.950 196.050 124.050 ;
        RECT 188.400 118.050 189.450 121.950 ;
        RECT 187.950 115.950 190.050 118.050 ;
        RECT 194.400 106.050 195.450 121.950 ;
        RECT 197.400 115.050 198.450 157.950 ;
        RECT 196.950 112.950 199.050 115.050 ;
        RECT 190.950 103.950 193.050 106.050 ;
        RECT 193.950 103.950 196.050 106.050 ;
        RECT 196.950 103.950 199.050 106.050 ;
        RECT 191.400 102.450 192.450 103.950 ;
        RECT 191.400 101.400 195.450 102.450 ;
        RECT 187.950 99.450 190.050 100.050 ;
        RECT 185.400 98.400 190.050 99.450 ;
        RECT 187.950 97.950 190.050 98.400 ;
        RECT 188.400 97.050 189.450 97.950 ;
        RECT 194.400 97.050 195.450 101.400 ;
        RECT 197.400 97.050 198.450 103.950 ;
        RECT 182.400 95.400 186.450 96.450 ;
        RECT 181.950 91.950 184.050 94.050 ;
        RECT 172.950 88.950 175.050 91.050 ;
        RECT 176.250 89.850 177.750 90.750 ;
        RECT 178.950 88.950 181.050 91.050 ;
        RECT 182.250 89.850 184.050 90.750 ;
        RECT 178.950 86.850 181.050 87.750 ;
        RECT 169.950 64.950 172.050 67.050 ;
        RECT 185.400 64.050 186.450 95.400 ;
        RECT 187.950 94.950 190.050 97.050 ;
        RECT 191.250 95.250 192.750 96.150 ;
        RECT 193.950 94.950 196.050 97.050 ;
        RECT 196.950 94.950 199.050 97.050 ;
        RECT 187.950 92.850 189.750 93.750 ;
        RECT 190.950 91.950 193.050 94.050 ;
        RECT 194.250 92.850 195.750 93.750 ;
        RECT 196.950 91.950 199.050 94.050 ;
        RECT 190.950 88.950 193.050 91.050 ;
        RECT 196.950 89.850 199.050 90.750 ;
        RECT 184.950 61.950 187.050 64.050 ;
        RECT 169.950 59.250 172.050 60.150 ;
        RECT 184.950 59.250 187.050 60.150 ;
        RECT 163.950 55.950 166.050 58.050 ;
        RECT 167.250 56.250 168.750 57.150 ;
        RECT 169.950 55.950 172.050 58.050 ;
        RECT 173.250 56.250 175.050 57.150 ;
        RECT 178.950 55.950 181.050 58.050 ;
        RECT 182.250 56.250 183.750 57.150 ;
        RECT 184.950 55.950 187.050 58.050 ;
        RECT 188.250 56.250 190.050 57.150 ;
        RECT 163.950 53.850 165.750 54.750 ;
        RECT 166.950 52.950 169.050 55.050 ;
        RECT 172.950 52.950 175.050 55.050 ;
        RECT 175.950 52.950 178.050 55.050 ;
        RECT 178.950 53.850 180.750 54.750 ;
        RECT 181.950 52.950 184.050 55.050 ;
        RECT 167.400 52.050 168.450 52.950 ;
        RECT 166.950 49.950 169.050 52.050 ;
        RECT 173.400 43.050 174.450 52.950 ;
        RECT 172.950 40.950 175.050 43.050 ;
        RECT 169.950 31.950 172.050 34.050 ;
        RECT 161.400 26.400 165.450 27.450 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 146.250 23.250 147.750 24.150 ;
        RECT 148.950 22.950 151.050 25.050 ;
        RECT 151.950 22.950 154.050 25.050 ;
        RECT 155.250 23.250 156.750 24.150 ;
        RECT 157.950 22.950 160.050 25.050 ;
        RECT 160.950 22.950 163.050 25.050 ;
        RECT 161.400 22.050 162.450 22.950 ;
        RECT 164.400 22.050 165.450 26.400 ;
        RECT 170.400 25.050 171.450 31.950 ;
        RECT 176.400 25.050 177.450 52.950 ;
        RECT 185.400 43.050 186.450 55.950 ;
        RECT 187.950 54.450 190.050 55.050 ;
        RECT 191.400 54.450 192.450 88.950 ;
        RECT 200.400 88.050 201.450 161.400 ;
        RECT 227.400 160.050 228.450 167.400 ;
        RECT 214.950 157.950 217.050 160.050 ;
        RECT 226.950 157.950 229.050 160.050 ;
        RECT 205.950 145.950 208.050 148.050 ;
        RECT 206.400 130.050 207.450 145.950 ;
        RECT 205.950 129.450 208.050 130.050 ;
        RECT 205.950 128.400 210.450 129.450 ;
        RECT 205.950 127.950 208.050 128.400 ;
        RECT 202.950 125.250 205.050 126.150 ;
        RECT 205.950 125.850 208.050 126.750 ;
        RECT 202.950 121.950 205.050 124.050 ;
        RECT 209.400 111.450 210.450 128.400 ;
        RECT 211.950 125.250 214.050 126.150 ;
        RECT 215.400 124.050 216.450 157.950 ;
        RECT 223.950 154.950 226.050 157.050 ;
        RECT 224.400 130.050 225.450 154.950 ;
        RECT 226.950 148.950 229.050 151.050 ;
        RECT 217.950 127.950 220.050 130.050 ;
        RECT 221.250 128.250 222.750 129.150 ;
        RECT 223.950 127.950 226.050 130.050 ;
        RECT 217.950 125.850 219.750 126.750 ;
        RECT 220.950 124.950 223.050 127.050 ;
        RECT 224.250 125.850 226.050 126.750 ;
        RECT 211.950 121.950 214.050 124.050 ;
        RECT 214.950 121.950 217.050 124.050 ;
        RECT 212.400 112.050 213.450 121.950 ;
        RECT 221.400 121.050 222.450 124.950 ;
        RECT 227.400 121.050 228.450 148.950 ;
        RECT 230.400 139.050 231.450 217.950 ;
        RECT 233.400 202.050 234.450 239.400 ;
        RECT 239.400 238.050 240.450 239.400 ;
        RECT 235.950 236.250 237.750 237.150 ;
        RECT 238.950 235.950 241.050 238.050 ;
        RECT 242.250 236.250 244.050 237.150 ;
        RECT 235.950 232.950 238.050 235.050 ;
        RECT 239.250 233.850 240.750 234.750 ;
        RECT 241.950 232.950 244.050 235.050 ;
        RECT 245.400 232.050 246.450 262.950 ;
        RECT 248.400 250.050 249.450 265.950 ;
        RECT 247.950 247.950 250.050 250.050 ;
        RECT 251.400 246.450 252.450 271.950 ;
        RECT 257.400 267.450 258.450 295.950 ;
        RECT 260.400 295.050 261.450 307.950 ;
        RECT 269.400 295.050 270.450 307.950 ;
        RECT 278.400 307.050 279.450 314.400 ;
        RECT 280.950 313.950 283.050 314.400 ;
        RECT 280.950 311.850 283.050 312.750 ;
        RECT 283.950 311.250 286.050 312.150 ;
        RECT 280.950 307.950 283.050 310.050 ;
        RECT 283.950 307.950 286.050 310.050 ;
        RECT 274.950 305.850 277.050 306.750 ;
        RECT 277.950 304.950 280.050 307.050 ;
        RECT 274.950 295.950 277.050 298.050 ;
        RECT 259.950 292.950 262.050 295.050 ;
        RECT 268.950 292.950 271.050 295.050 ;
        RECT 262.950 289.950 265.050 292.050 ;
        RECT 263.400 271.050 264.450 289.950 ;
        RECT 268.950 271.950 271.050 274.050 ;
        RECT 269.400 271.050 270.450 271.950 ;
        RECT 259.950 269.250 261.750 270.150 ;
        RECT 262.950 268.950 265.050 271.050 ;
        RECT 268.950 268.950 271.050 271.050 ;
        RECT 259.950 267.450 262.050 268.050 ;
        RECT 257.400 266.400 262.050 267.450 ;
        RECT 263.250 266.850 265.050 267.750 ;
        RECT 259.950 265.950 262.050 266.400 ;
        RECT 265.950 266.250 268.050 267.150 ;
        RECT 268.950 266.850 271.050 267.750 ;
        RECT 265.950 262.950 268.050 265.050 ;
        RECT 268.950 253.950 271.050 256.050 ;
        RECT 259.950 247.950 262.050 250.050 ;
        RECT 248.400 245.400 252.450 246.450 ;
        RECT 241.950 229.950 244.050 232.050 ;
        RECT 244.950 229.950 247.050 232.050 ;
        RECT 238.950 214.950 241.050 217.050 ;
        RECT 235.950 208.950 238.050 211.050 ;
        RECT 232.950 199.950 235.050 202.050 ;
        RECT 236.400 199.050 237.450 208.950 ;
        RECT 239.400 202.050 240.450 214.950 ;
        RECT 238.950 199.950 241.050 202.050 ;
        RECT 242.400 199.050 243.450 229.950 ;
        RECT 248.400 202.050 249.450 245.400 ;
        RECT 260.400 241.050 261.450 247.950 ;
        RECT 269.400 244.050 270.450 253.950 ;
        RECT 275.400 250.050 276.450 295.950 ;
        RECT 278.400 292.050 279.450 304.950 ;
        RECT 277.950 289.950 280.050 292.050 ;
        RECT 277.950 269.250 280.050 270.150 ;
        RECT 277.950 265.950 280.050 268.050 ;
        RECT 281.400 265.050 282.450 307.950 ;
        RECT 287.400 304.050 288.450 364.950 ;
        RECT 292.950 352.950 295.050 355.050 ;
        RECT 289.950 341.250 292.050 342.150 ;
        RECT 289.950 337.950 292.050 340.050 ;
        RECT 293.400 334.050 294.450 352.950 ;
        RECT 295.950 341.250 298.050 342.150 ;
        RECT 295.950 337.950 298.050 340.050 ;
        RECT 292.950 331.950 295.050 334.050 ;
        RECT 296.400 325.050 297.450 337.950 ;
        RECT 295.950 322.950 298.050 325.050 ;
        RECT 302.400 322.050 303.450 382.950 ;
        RECT 305.400 372.600 306.600 389.400 ;
        RECT 304.950 370.500 307.050 372.600 ;
        RECT 308.400 366.450 309.450 400.950 ;
        RECT 310.950 391.950 313.050 394.050 ;
        RECT 311.400 385.050 312.450 391.950 ;
        RECT 310.950 382.950 313.050 385.050 ;
        RECT 310.950 380.850 313.050 381.750 ;
        RECT 314.400 367.050 315.450 470.400 ;
        RECT 323.400 457.050 324.450 478.950 ;
        RECT 326.400 466.050 327.450 517.950 ;
        RECT 329.400 493.050 330.450 517.950 ;
        RECT 338.400 514.050 339.450 521.400 ;
        RECT 337.950 511.950 340.050 514.050 ;
        RECT 334.950 494.400 337.050 496.500 ;
        RECT 328.950 490.950 331.050 493.050 ;
        RECT 328.950 485.250 331.050 486.150 ;
        RECT 328.950 481.950 331.050 484.050 ;
        RECT 329.400 481.050 330.450 481.950 ;
        RECT 328.950 478.950 331.050 481.050 ;
        RECT 335.400 477.600 336.600 494.400 ;
        RECT 334.950 475.500 337.050 477.600 ;
        RECT 325.950 463.950 328.050 466.050 ;
        RECT 338.400 463.050 339.450 511.950 ;
        RECT 341.400 496.050 342.450 529.950 ;
        RECT 350.400 529.050 351.450 532.950 ;
        RECT 343.950 526.950 346.050 529.050 ;
        RECT 347.250 527.250 348.750 528.150 ;
        RECT 349.950 526.950 352.050 529.050 ;
        RECT 343.950 524.850 345.750 525.750 ;
        RECT 346.950 523.950 349.050 526.050 ;
        RECT 350.250 524.850 351.750 525.750 ;
        RECT 352.950 523.950 355.050 526.050 ;
        RECT 347.400 505.050 348.450 523.950 ;
        RECT 352.950 521.850 355.050 522.750 ;
        RECT 356.400 517.050 357.450 554.400 ;
        RECT 358.950 554.400 363.450 555.450 ;
        RECT 358.950 553.950 361.050 554.400 ;
        RECT 365.400 549.600 366.600 566.400 ;
        RECT 368.400 550.050 369.450 586.950 ;
        RECT 382.950 586.500 385.050 588.600 ;
        RECT 379.950 571.950 382.050 574.050 ;
        RECT 373.950 568.950 376.050 571.050 ;
        RECT 370.950 565.950 373.050 568.050 ;
        RECT 371.400 559.050 372.450 565.950 ;
        RECT 374.400 559.050 375.450 568.950 ;
        RECT 370.950 556.950 373.050 559.050 ;
        RECT 373.950 556.950 376.050 559.050 ;
        RECT 376.950 556.950 379.050 559.050 ;
        RECT 373.950 554.250 376.050 555.150 ;
        RECT 376.950 554.850 379.050 555.750 ;
        RECT 373.950 550.950 376.050 553.050 ;
        RECT 364.950 547.500 367.050 549.600 ;
        RECT 367.950 547.950 370.050 550.050 ;
        RECT 373.950 547.950 376.050 550.050 ;
        RECT 358.950 541.950 361.050 544.050 ;
        RECT 367.950 541.950 370.050 544.050 ;
        RECT 355.950 514.950 358.050 517.050 ;
        RECT 359.400 514.050 360.450 541.950 ;
        RECT 361.950 538.950 364.050 541.050 ;
        RECT 362.400 529.050 363.450 538.950 ;
        RECT 364.950 529.950 367.050 532.050 ;
        RECT 368.400 529.050 369.450 541.950 ;
        RECT 370.950 538.950 373.050 541.050 ;
        RECT 361.950 526.950 364.050 529.050 ;
        RECT 365.250 527.850 366.750 528.750 ;
        RECT 367.950 526.950 370.050 529.050 ;
        RECT 361.950 524.850 364.050 525.750 ;
        RECT 364.950 523.950 367.050 526.050 ;
        RECT 367.950 524.850 370.050 525.750 ;
        RECT 361.950 520.950 364.050 523.050 ;
        RECT 358.950 511.950 361.050 514.050 ;
        RECT 346.950 502.950 349.050 505.050 ;
        RECT 346.950 496.950 349.050 499.050 ;
        RECT 355.950 496.950 358.050 499.050 ;
        RECT 340.950 493.950 343.050 496.050 ;
        RECT 343.950 485.250 346.050 486.150 ;
        RECT 343.950 481.950 346.050 484.050 ;
        RECT 347.400 483.450 348.450 496.950 ;
        RECT 356.400 490.050 357.450 496.950 ;
        RECT 362.400 490.050 363.450 520.950 ;
        RECT 365.400 502.050 366.450 523.950 ;
        RECT 367.950 517.950 370.050 520.050 ;
        RECT 364.950 499.950 367.050 502.050 ;
        RECT 364.950 493.950 367.050 496.050 ;
        RECT 355.950 487.950 358.050 490.050 ;
        RECT 359.250 488.250 360.750 489.150 ;
        RECT 361.950 487.950 364.050 490.050 ;
        RECT 349.950 485.250 352.050 486.150 ;
        RECT 355.950 485.850 357.750 486.750 ;
        RECT 358.950 484.950 361.050 487.050 ;
        RECT 362.250 485.850 364.050 486.750 ;
        RECT 349.950 483.450 352.050 484.050 ;
        RECT 347.400 482.400 352.050 483.450 ;
        RECT 349.950 481.950 352.050 482.400 ;
        RECT 344.400 480.450 345.450 481.950 ;
        RECT 365.400 481.050 366.450 493.950 ;
        RECT 344.400 479.400 348.450 480.450 ;
        RECT 337.950 460.950 340.050 463.050 ;
        RECT 337.950 457.950 340.050 460.050 ;
        RECT 343.950 457.950 346.050 460.050 ;
        RECT 344.400 457.050 345.450 457.950 ;
        RECT 316.950 454.950 319.050 457.050 ;
        RECT 320.250 455.250 321.750 456.150 ;
        RECT 322.950 454.950 325.050 457.050 ;
        RECT 326.250 455.250 327.750 456.150 ;
        RECT 328.950 454.950 331.050 457.050 ;
        RECT 331.950 454.950 334.050 457.050 ;
        RECT 334.950 455.250 337.050 456.150 ;
        RECT 337.950 455.850 340.050 456.750 ;
        RECT 340.950 455.250 342.750 456.150 ;
        RECT 343.950 454.950 346.050 457.050 ;
        RECT 316.950 452.850 318.750 453.750 ;
        RECT 319.950 451.950 322.050 454.050 ;
        RECT 323.250 452.850 324.750 453.750 ;
        RECT 325.950 451.950 328.050 454.050 ;
        RECT 329.250 452.850 331.050 453.750 ;
        RECT 320.400 433.050 321.450 451.950 ;
        RECT 326.400 448.050 327.450 451.950 ;
        RECT 328.950 448.950 331.050 451.050 ;
        RECT 325.950 445.950 328.050 448.050 ;
        RECT 319.950 430.950 322.050 433.050 ;
        RECT 320.400 421.050 321.450 430.950 ;
        RECT 319.950 418.950 322.050 421.050 ;
        RECT 316.950 416.250 319.050 417.150 ;
        RECT 316.950 412.950 319.050 415.050 ;
        RECT 320.250 413.250 321.750 414.150 ;
        RECT 322.950 412.950 325.050 415.050 ;
        RECT 326.250 413.250 328.050 414.150 ;
        RECT 317.400 406.050 318.450 412.950 ;
        RECT 319.950 409.950 322.050 412.050 ;
        RECT 323.250 410.850 324.750 411.750 ;
        RECT 325.950 409.950 328.050 412.050 ;
        RECT 320.400 409.050 321.450 409.950 ;
        RECT 319.950 406.950 322.050 409.050 ;
        RECT 326.400 408.450 327.450 409.950 ;
        RECT 329.400 409.050 330.450 448.950 ;
        RECT 332.400 448.050 333.450 454.950 ;
        RECT 334.950 451.950 337.050 454.050 ;
        RECT 340.950 451.950 343.050 454.050 ;
        RECT 344.250 452.850 346.050 453.750 ;
        RECT 331.950 445.950 334.050 448.050 ;
        RECT 335.400 445.050 336.450 451.950 ;
        RECT 341.400 451.050 342.450 451.950 ;
        RECT 340.950 448.950 343.050 451.050 ;
        RECT 347.400 448.050 348.450 479.400 ;
        RECT 364.950 478.950 367.050 481.050 ;
        RECT 368.400 472.050 369.450 517.950 ;
        RECT 371.400 499.050 372.450 538.950 ;
        RECT 370.950 496.950 373.050 499.050 ;
        RECT 374.400 493.050 375.450 547.950 ;
        RECT 380.400 544.050 381.450 571.950 ;
        RECT 401.400 562.050 402.450 592.950 ;
        RECT 403.950 591.300 406.050 593.400 ;
        RECT 404.250 587.700 405.450 591.300 ;
        RECT 407.400 589.050 408.450 598.950 ;
        RECT 409.950 595.950 412.050 598.050 ;
        RECT 403.950 585.600 406.050 587.700 ;
        RECT 406.950 586.950 409.050 589.050 ;
        RECT 406.950 580.950 409.050 583.050 ;
        RECT 407.400 562.050 408.450 580.950 ;
        RECT 410.400 562.050 411.450 595.950 ;
        RECT 412.950 589.950 415.050 592.050 ;
        RECT 413.400 562.050 414.450 589.950 ;
        RECT 416.400 589.050 417.450 598.950 ;
        RECT 419.550 593.400 420.750 605.400 ;
        RECT 428.400 601.050 429.450 622.950 ;
        RECT 431.400 616.050 432.450 662.400 ;
        RECT 434.400 661.050 435.450 662.400 ;
        RECT 433.950 658.950 436.050 661.050 ;
        RECT 440.400 658.050 441.450 667.950 ;
        RECT 439.950 655.950 442.050 658.050 ;
        RECT 436.950 649.950 439.050 652.050 ;
        RECT 433.950 629.250 436.050 630.150 ;
        RECT 433.950 625.950 436.050 628.050 ;
        RECT 430.950 613.950 433.050 616.050 ;
        RECT 427.950 598.950 430.050 601.050 ;
        RECT 427.950 596.850 430.050 597.750 ;
        RECT 431.400 594.450 432.450 613.950 ;
        RECT 433.950 598.950 436.050 601.050 ;
        RECT 433.950 596.850 436.050 597.750 ;
        RECT 428.400 593.400 432.450 594.450 ;
        RECT 418.950 591.300 421.050 593.400 ;
        RECT 415.950 586.950 418.050 589.050 ;
        RECT 419.550 587.700 420.750 591.300 ;
        RECT 418.950 585.600 421.050 587.700 ;
        RECT 421.950 580.950 424.050 583.050 ;
        RECT 391.950 560.250 394.050 561.150 ;
        RECT 394.950 559.950 397.050 562.050 ;
        RECT 400.950 559.950 403.050 562.050 ;
        RECT 404.250 560.250 405.750 561.150 ;
        RECT 406.950 559.950 409.050 562.050 ;
        RECT 409.950 559.950 412.050 562.050 ;
        RECT 412.950 559.950 415.050 562.050 ;
        RECT 415.950 560.250 418.050 561.150 ;
        RECT 382.950 557.250 384.750 558.150 ;
        RECT 385.950 556.950 388.050 559.050 ;
        RECT 389.250 557.250 390.750 558.150 ;
        RECT 391.950 556.950 394.050 559.050 ;
        RECT 382.950 553.950 385.050 556.050 ;
        RECT 386.250 554.850 387.750 555.750 ;
        RECT 388.950 553.950 391.050 556.050 ;
        RECT 391.950 553.950 394.050 556.050 ;
        RECT 389.400 544.050 390.450 553.950 ;
        RECT 392.400 550.050 393.450 553.950 ;
        RECT 391.950 547.950 394.050 550.050 ;
        RECT 395.400 544.050 396.450 559.950 ;
        RECT 422.400 559.050 423.450 580.950 ;
        RECT 400.950 557.850 402.750 558.750 ;
        RECT 403.950 556.950 406.050 559.050 ;
        RECT 407.250 557.850 409.050 558.750 ;
        RECT 409.950 558.450 412.050 559.050 ;
        RECT 415.950 558.450 418.050 559.050 ;
        RECT 409.950 557.400 418.050 558.450 ;
        RECT 409.950 556.950 412.050 557.400 ;
        RECT 415.950 556.950 418.050 557.400 ;
        RECT 419.250 557.250 420.750 558.150 ;
        RECT 421.950 556.950 424.050 559.050 ;
        RECT 425.250 557.250 427.050 558.150 ;
        RECT 400.950 553.950 403.050 556.050 ;
        RECT 412.950 553.950 415.050 556.050 ;
        RECT 418.950 553.950 421.050 556.050 ;
        RECT 422.250 554.850 423.750 555.750 ;
        RECT 424.950 553.950 427.050 556.050 ;
        RECT 379.950 541.950 382.050 544.050 ;
        RECT 388.950 541.950 391.050 544.050 ;
        RECT 394.950 541.950 397.050 544.050 ;
        RECT 397.950 541.950 400.050 544.050 ;
        RECT 388.950 538.950 391.050 541.050 ;
        RECT 391.950 538.950 394.050 541.050 ;
        RECT 379.950 532.950 382.050 535.050 ;
        RECT 376.950 529.950 379.050 532.050 ;
        RECT 377.400 526.050 378.450 529.950 ;
        RECT 380.400 529.050 381.450 532.950 ;
        RECT 389.400 532.050 390.450 538.950 ;
        RECT 388.950 529.950 391.050 532.050 ;
        RECT 379.950 526.950 382.050 529.050 ;
        RECT 383.250 527.250 384.750 528.150 ;
        RECT 385.950 526.950 388.050 529.050 ;
        RECT 392.400 526.050 393.450 538.950 ;
        RECT 398.400 532.050 399.450 541.950 ;
        RECT 401.400 541.050 402.450 553.950 ;
        RECT 403.950 544.950 406.050 547.050 ;
        RECT 400.950 538.950 403.050 541.050 ;
        RECT 397.950 529.950 400.050 532.050 ;
        RECT 400.950 529.950 403.050 532.050 ;
        RECT 397.950 526.950 400.050 529.050 ;
        RECT 376.950 523.950 379.050 526.050 ;
        RECT 380.250 524.850 381.750 525.750 ;
        RECT 382.950 523.950 385.050 526.050 ;
        RECT 386.250 524.850 388.050 525.750 ;
        RECT 388.950 524.250 390.750 525.150 ;
        RECT 391.950 523.950 394.050 526.050 ;
        RECT 395.250 524.250 397.050 525.150 ;
        RECT 376.950 521.850 379.050 522.750 ;
        RECT 383.400 496.050 384.450 523.950 ;
        RECT 388.950 520.950 391.050 523.050 ;
        RECT 392.250 521.850 393.750 522.750 ;
        RECT 394.950 522.450 397.050 523.050 ;
        RECT 398.400 522.450 399.450 526.950 ;
        RECT 394.950 521.400 399.450 522.450 ;
        RECT 394.950 520.950 397.050 521.400 ;
        RECT 389.400 502.050 390.450 520.950 ;
        RECT 391.950 505.950 394.050 508.050 ;
        RECT 388.950 499.950 391.050 502.050 ;
        RECT 382.950 493.950 385.050 496.050 ;
        RECT 373.950 490.950 376.050 493.050 ;
        RECT 382.950 490.950 385.050 493.050 ;
        RECT 370.950 488.250 373.050 489.150 ;
        RECT 370.950 484.950 373.050 487.050 ;
        RECT 374.250 485.250 375.750 486.150 ;
        RECT 376.950 484.950 379.050 487.050 ;
        RECT 380.250 485.250 382.050 486.150 ;
        RECT 373.950 481.950 376.050 484.050 ;
        RECT 377.250 482.850 378.750 483.750 ;
        RECT 379.950 481.950 382.050 484.050 ;
        RECT 367.950 469.950 370.050 472.050 ;
        RECT 358.950 466.950 361.050 469.050 ;
        RECT 359.400 460.050 360.450 466.950 ;
        RECT 370.950 461.400 373.050 463.500 ;
        RECT 358.950 457.950 361.050 460.050 ;
        RECT 364.950 457.950 367.050 460.050 ;
        RECT 367.950 458.250 370.050 459.150 ;
        RECT 352.950 454.950 355.050 457.050 ;
        RECT 356.250 455.250 358.050 456.150 ;
        RECT 358.950 455.850 361.050 456.750 ;
        RECT 361.950 455.250 364.050 456.150 ;
        RECT 352.950 452.850 354.750 453.750 ;
        RECT 355.950 451.950 358.050 454.050 ;
        RECT 361.950 451.950 364.050 454.050 ;
        RECT 352.950 448.950 355.050 451.050 ;
        RECT 340.950 445.950 343.050 448.050 ;
        RECT 346.950 445.950 349.050 448.050 ;
        RECT 334.950 442.950 337.050 445.050 ;
        RECT 335.400 433.050 336.450 442.950 ;
        RECT 334.950 430.950 337.050 433.050 ;
        RECT 337.950 418.950 340.050 421.050 ;
        RECT 331.950 416.250 334.050 417.150 ;
        RECT 338.400 415.050 339.450 418.950 ;
        RECT 341.400 418.050 342.450 445.950 ;
        RECT 353.400 433.050 354.450 448.950 ;
        RECT 349.950 430.950 352.050 433.050 ;
        RECT 352.950 430.950 355.050 433.050 ;
        RECT 343.950 427.950 346.050 430.050 ;
        RECT 344.400 418.050 345.450 427.950 ;
        RECT 350.400 418.050 351.450 430.950 ;
        RECT 340.950 415.950 343.050 418.050 ;
        RECT 343.950 415.950 346.050 418.050 ;
        RECT 347.250 416.250 348.750 417.150 ;
        RECT 349.950 415.950 352.050 418.050 ;
        RECT 335.250 413.250 336.750 414.150 ;
        RECT 337.950 412.950 340.050 415.050 ;
        RECT 341.250 413.250 343.050 414.150 ;
        RECT 343.950 413.850 345.750 414.750 ;
        RECT 346.950 412.950 349.050 415.050 ;
        RECT 350.250 413.850 352.050 414.750 ;
        RECT 331.950 409.950 334.050 412.050 ;
        RECT 334.950 409.950 337.050 412.050 ;
        RECT 338.250 410.850 339.750 411.750 ;
        RECT 340.950 411.450 343.050 412.050 ;
        RECT 340.950 410.400 345.450 411.450 ;
        RECT 340.950 409.950 343.050 410.400 ;
        RECT 323.400 407.400 327.450 408.450 ;
        RECT 316.950 403.950 319.050 406.050 ;
        RECT 316.950 388.950 319.050 391.050 ;
        RECT 317.400 385.050 318.450 388.950 ;
        RECT 316.950 382.950 319.050 385.050 ;
        RECT 316.950 380.850 319.050 381.750 ;
        RECT 323.400 367.050 324.450 407.400 ;
        RECT 328.950 406.950 331.050 409.050 ;
        RECT 325.950 389.400 328.050 391.500 ;
        RECT 326.250 377.400 327.450 389.400 ;
        RECT 328.950 386.250 331.050 387.150 ;
        RECT 328.950 382.950 331.050 385.050 ;
        RECT 332.400 379.050 333.450 409.950 ;
        RECT 335.400 400.050 336.450 409.950 ;
        RECT 337.950 406.950 340.050 409.050 ;
        RECT 338.400 403.050 339.450 406.950 ;
        RECT 344.400 406.050 345.450 410.400 ;
        RECT 347.400 409.050 348.450 412.950 ;
        RECT 349.950 409.950 352.050 412.050 ;
        RECT 346.950 406.950 349.050 409.050 ;
        RECT 343.950 403.950 346.050 406.050 ;
        RECT 337.950 400.950 340.050 403.050 ;
        RECT 334.950 397.950 337.050 400.050 ;
        RECT 337.950 397.950 340.050 400.050 ;
        RECT 338.400 388.050 339.450 397.950 ;
        RECT 350.400 388.050 351.450 409.950 ;
        RECT 353.400 406.050 354.450 430.950 ;
        RECT 356.400 421.050 357.450 451.950 ;
        RECT 358.950 424.950 361.050 427.050 ;
        RECT 355.950 418.950 358.050 421.050 ;
        RECT 359.400 417.450 360.450 424.950 ;
        RECT 361.950 418.950 364.050 421.050 ;
        RECT 356.400 416.400 360.450 417.450 ;
        RECT 352.950 403.950 355.050 406.050 ;
        RECT 356.400 397.050 357.450 416.400 ;
        RECT 362.400 415.050 363.450 418.950 ;
        RECT 365.400 415.050 366.450 457.950 ;
        RECT 367.950 454.950 370.050 457.050 ;
        RECT 368.400 448.050 369.450 454.950 ;
        RECT 371.550 449.400 372.750 461.400 ;
        RECT 374.400 454.050 375.450 481.950 ;
        RECT 379.950 478.950 382.050 481.050 ;
        RECT 376.950 463.950 379.050 466.050 ;
        RECT 373.950 451.950 376.050 454.050 ;
        RECT 367.950 445.950 370.050 448.050 ;
        RECT 370.950 447.300 373.050 449.400 ;
        RECT 371.550 443.700 372.750 447.300 ;
        RECT 370.950 441.600 373.050 443.700 ;
        RECT 377.400 430.050 378.450 463.950 ;
        RECT 380.400 460.050 381.450 478.950 ;
        RECT 383.400 466.050 384.450 490.950 ;
        RECT 392.400 490.050 393.450 505.950 ;
        RECT 401.400 496.050 402.450 529.950 ;
        RECT 404.400 520.050 405.450 544.950 ;
        RECT 413.400 544.050 414.450 553.950 ;
        RECT 415.950 550.950 418.050 553.050 ;
        RECT 412.950 541.950 415.050 544.050 ;
        RECT 406.950 532.950 409.050 535.050 ;
        RECT 407.400 526.050 408.450 532.950 ;
        RECT 416.400 531.450 417.450 550.950 ;
        RECT 419.400 547.050 420.450 553.950 ;
        RECT 428.400 553.050 429.450 593.400 ;
        RECT 437.400 568.050 438.450 649.950 ;
        RECT 439.950 638.400 442.050 640.500 ;
        RECT 440.400 621.600 441.600 638.400 ;
        RECT 443.400 625.050 444.450 697.950 ;
        RECT 449.400 693.600 450.600 710.400 ;
        RECT 470.250 707.700 471.450 711.300 ;
        RECT 548.550 707.700 549.750 711.300 ;
        RECT 568.950 710.400 571.050 712.500 ;
        RECT 469.950 705.600 472.050 707.700 ;
        RECT 454.950 701.250 457.050 702.150 ;
        RECT 460.950 701.250 463.050 702.150 ;
        RECT 454.950 697.950 457.050 700.050 ;
        RECT 460.950 697.950 463.050 700.050 ;
        RECT 448.950 691.500 451.050 693.600 ;
        RECT 451.950 673.950 454.050 676.050 ;
        RECT 452.400 670.050 453.450 673.950 ;
        RECT 455.400 673.050 456.450 697.950 ;
        RECT 470.250 693.600 471.450 705.600 ;
        RECT 520.950 704.250 523.050 705.150 ;
        RECT 523.950 703.950 526.050 706.050 ;
        RECT 532.950 705.450 535.050 706.050 ;
        RECT 530.400 704.400 535.050 705.450 ;
        RECT 478.950 700.950 481.050 703.050 ;
        RECT 484.950 700.950 487.050 703.050 ;
        RECT 493.950 700.950 496.050 703.050 ;
        RECT 511.950 701.250 513.750 702.150 ;
        RECT 514.950 700.950 517.050 703.050 ;
        RECT 518.250 701.250 519.750 702.150 ;
        RECT 520.950 700.950 523.050 703.050 ;
        RECT 479.400 700.050 480.450 700.950 ;
        RECT 472.950 699.450 475.050 700.050 ;
        RECT 472.950 698.400 477.450 699.450 ;
        RECT 472.950 697.950 475.050 698.400 ;
        RECT 472.950 695.850 475.050 696.750 ;
        RECT 469.950 691.500 472.050 693.600 ;
        RECT 469.950 677.400 472.050 679.500 ;
        RECT 466.950 674.250 469.050 675.150 ;
        RECT 454.950 670.950 457.050 673.050 ;
        RECT 460.950 672.450 463.050 673.050 ;
        RECT 458.250 671.250 459.750 672.150 ;
        RECT 460.950 671.400 465.450 672.450 ;
        RECT 460.950 670.950 463.050 671.400 ;
        RECT 464.400 670.050 465.450 671.400 ;
        RECT 466.950 670.950 469.050 673.050 ;
        RECT 451.950 667.950 454.050 670.050 ;
        RECT 455.250 668.850 456.750 669.750 ;
        RECT 457.950 667.950 460.050 670.050 ;
        RECT 461.250 668.850 463.050 669.750 ;
        RECT 463.950 667.950 466.050 670.050 ;
        RECT 458.400 667.050 459.450 667.950 ;
        RECT 451.950 665.850 454.050 666.750 ;
        RECT 457.950 664.950 460.050 667.050 ;
        RECT 458.400 640.050 459.450 664.950 ;
        RECT 467.400 664.050 468.450 670.950 ;
        RECT 470.550 665.400 471.750 677.400 ;
        RECT 466.950 661.950 469.050 664.050 ;
        RECT 469.950 663.300 472.050 665.400 ;
        RECT 470.550 659.700 471.750 663.300 ;
        RECT 476.400 661.050 477.450 698.400 ;
        RECT 478.950 697.950 481.050 700.050 ;
        RECT 484.950 698.850 487.050 699.750 ;
        RECT 479.400 673.050 480.450 697.950 ;
        RECT 484.950 676.950 487.050 679.050 ;
        RECT 490.950 677.400 493.050 679.500 ;
        RECT 485.400 673.050 486.450 676.950 ;
        RECT 478.950 670.950 481.050 673.050 ;
        RECT 484.950 670.950 487.050 673.050 ;
        RECT 478.950 668.850 481.050 669.750 ;
        RECT 484.950 668.850 487.050 669.750 ;
        RECT 469.950 657.600 472.050 659.700 ;
        RECT 475.950 658.950 478.050 661.050 ;
        RECT 491.400 660.600 492.600 677.400 ;
        RECT 494.400 670.050 495.450 700.950 ;
        RECT 521.400 700.050 522.450 700.950 ;
        RECT 505.950 698.850 508.050 699.750 ;
        RECT 511.950 697.950 514.050 700.050 ;
        RECT 515.250 698.850 516.750 699.750 ;
        RECT 517.950 697.950 520.050 700.050 ;
        RECT 520.950 697.950 523.050 700.050 ;
        RECT 512.400 694.050 513.450 697.950 ;
        RECT 518.400 697.050 519.450 697.950 ;
        RECT 517.950 694.950 520.050 697.050 ;
        RECT 511.950 691.950 514.050 694.050 ;
        RECT 505.950 676.950 508.050 679.050 ;
        RECT 506.400 673.050 507.450 676.950 ;
        RECT 499.950 670.950 502.050 673.050 ;
        RECT 503.250 671.250 504.750 672.150 ;
        RECT 505.950 670.950 508.050 673.050 ;
        RECT 493.950 667.950 496.050 670.050 ;
        RECT 499.950 668.850 501.750 669.750 ;
        RECT 502.950 667.950 505.050 670.050 ;
        RECT 506.250 668.850 507.750 669.750 ;
        RECT 508.950 667.950 511.050 670.050 ;
        RECT 514.950 668.250 516.750 669.150 ;
        RECT 517.950 667.950 520.050 670.050 ;
        RECT 521.250 668.250 523.050 669.150 ;
        RECT 490.950 658.500 493.050 660.600 ;
        RECT 457.950 637.950 460.050 640.050 ;
        RECT 484.950 639.300 487.050 641.400 ;
        RECT 466.950 634.950 469.050 637.050 ;
        RECT 485.550 635.700 486.750 639.300 ;
        RECT 487.950 637.950 490.050 640.050 ;
        RECT 467.400 634.050 468.450 634.950 ;
        RECT 454.950 632.250 457.050 633.150 ;
        RECT 460.950 631.950 463.050 634.050 ;
        RECT 466.950 631.950 469.050 634.050 ;
        RECT 470.250 632.250 471.750 633.150 ;
        RECT 472.950 631.950 475.050 634.050 ;
        RECT 484.950 633.600 487.050 635.700 ;
        RECT 461.400 631.050 462.450 631.950 ;
        RECT 454.950 628.950 457.050 631.050 ;
        RECT 458.250 629.250 459.750 630.150 ;
        RECT 460.950 628.950 463.050 631.050 ;
        RECT 464.250 629.250 466.050 630.150 ;
        RECT 466.950 629.850 468.750 630.750 ;
        RECT 469.950 628.950 472.050 631.050 ;
        RECT 473.250 629.850 475.050 630.750 ;
        RECT 457.950 625.950 460.050 628.050 ;
        RECT 461.250 626.850 462.750 627.750 ;
        RECT 463.950 625.950 466.050 628.050 ;
        RECT 466.950 625.950 469.050 628.050 ;
        RECT 481.950 625.950 484.050 628.050 ;
        RECT 442.950 622.950 445.050 625.050 ;
        RECT 439.950 619.500 442.050 621.600 ;
        RECT 442.950 607.950 445.050 610.050 ;
        RECT 439.950 605.400 442.050 607.500 ;
        RECT 440.400 588.600 441.600 605.400 ;
        RECT 439.950 586.500 442.050 588.600 ;
        RECT 436.950 565.950 439.050 568.050 ;
        RECT 433.950 559.950 436.050 562.050 ;
        RECT 439.950 560.250 442.050 561.150 ;
        RECT 434.400 559.050 435.450 559.950 ;
        RECT 430.950 557.250 432.750 558.150 ;
        RECT 433.950 556.950 436.050 559.050 ;
        RECT 437.250 557.250 438.750 558.150 ;
        RECT 439.950 556.950 442.050 559.050 ;
        RECT 430.950 553.950 433.050 556.050 ;
        RECT 434.250 554.850 435.750 555.750 ;
        RECT 436.950 553.950 439.050 556.050 ;
        RECT 427.950 550.950 430.050 553.050 ;
        RECT 439.950 550.950 442.050 553.050 ;
        RECT 436.950 547.950 439.050 550.050 ;
        RECT 418.950 544.950 421.050 547.050 ;
        RECT 427.950 538.950 430.050 541.050 ;
        RECT 424.950 532.950 427.050 535.050 ;
        RECT 418.950 531.450 421.050 532.050 ;
        RECT 416.400 530.400 421.050 531.450 ;
        RECT 418.950 529.950 421.050 530.400 ;
        RECT 409.950 526.950 412.050 529.050 ;
        RECT 413.250 527.250 414.750 528.150 ;
        RECT 415.950 526.950 418.050 529.050 ;
        RECT 418.950 527.850 421.050 528.750 ;
        RECT 421.950 527.250 424.050 528.150 ;
        RECT 406.950 523.950 409.050 526.050 ;
        RECT 410.250 524.850 411.750 525.750 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 416.250 524.850 418.050 525.750 ;
        RECT 421.950 523.950 424.050 526.050 ;
        RECT 406.950 521.850 409.050 522.750 ;
        RECT 403.950 517.950 406.050 520.050 ;
        RECT 413.400 514.050 414.450 523.950 ;
        RECT 425.400 522.450 426.450 532.950 ;
        RECT 428.400 532.050 429.450 538.950 ;
        RECT 427.950 529.950 430.050 532.050 ;
        RECT 430.950 529.950 433.050 532.050 ;
        RECT 431.400 526.050 432.450 529.950 ;
        RECT 427.950 524.250 429.750 525.150 ;
        RECT 430.950 523.950 433.050 526.050 ;
        RECT 434.250 524.250 436.050 525.150 ;
        RECT 422.400 521.400 426.450 522.450 ;
        RECT 412.950 511.950 415.050 514.050 ;
        RECT 409.950 496.950 412.050 499.050 ;
        RECT 400.950 493.950 403.050 496.050 ;
        RECT 406.950 490.950 409.050 493.050 ;
        RECT 407.400 490.050 408.450 490.950 ;
        RECT 388.950 488.250 391.050 489.150 ;
        RECT 391.950 487.950 394.050 490.050 ;
        RECT 394.950 487.950 397.050 490.050 ;
        RECT 406.950 487.950 409.050 490.050 ;
        RECT 395.400 487.050 396.450 487.950 ;
        RECT 392.250 485.250 393.750 486.150 ;
        RECT 394.950 484.950 397.050 487.050 ;
        RECT 398.250 485.250 400.050 486.150 ;
        RECT 400.950 484.950 403.050 487.050 ;
        RECT 403.950 485.250 406.050 486.150 ;
        RECT 406.950 485.850 409.050 486.750 ;
        RECT 391.950 481.950 394.050 484.050 ;
        RECT 395.250 482.850 396.750 483.750 ;
        RECT 397.950 481.950 400.050 484.050 ;
        RECT 401.400 483.450 402.450 484.950 ;
        RECT 403.950 483.450 406.050 484.050 ;
        RECT 401.400 482.400 406.050 483.450 ;
        RECT 403.950 481.950 406.050 482.400 ;
        RECT 385.950 469.950 388.050 472.050 ;
        RECT 382.950 463.950 385.050 466.050 ;
        RECT 379.950 457.950 382.050 460.050 ;
        RECT 386.400 457.050 387.450 469.950 ;
        RECT 410.400 469.050 411.450 496.950 ;
        RECT 422.400 496.050 423.450 521.400 ;
        RECT 427.950 520.950 430.050 523.050 ;
        RECT 431.250 521.850 432.750 522.750 ;
        RECT 433.950 520.950 436.050 523.050 ;
        RECT 434.400 520.050 435.450 520.950 ;
        RECT 424.950 517.950 427.050 520.050 ;
        RECT 433.950 517.950 436.050 520.050 ;
        RECT 415.950 493.950 418.050 496.050 ;
        RECT 421.950 493.950 424.050 496.050 ;
        RECT 412.950 485.250 415.050 486.150 ;
        RECT 412.950 481.950 415.050 484.050 ;
        RECT 394.950 466.950 397.050 469.050 ;
        RECT 409.950 466.950 412.050 469.050 ;
        RECT 391.950 461.400 394.050 463.500 ;
        RECT 379.950 456.450 382.050 457.050 ;
        RECT 379.950 455.400 384.450 456.450 ;
        RECT 379.950 454.950 382.050 455.400 ;
        RECT 379.950 452.850 382.050 453.750 ;
        RECT 383.400 451.050 384.450 455.400 ;
        RECT 385.950 454.950 388.050 457.050 ;
        RECT 385.950 452.850 388.050 453.750 ;
        RECT 382.950 448.950 385.050 451.050 ;
        RECT 385.950 445.950 388.050 448.050 ;
        RECT 370.950 427.950 373.050 430.050 ;
        RECT 376.950 427.950 379.050 430.050 ;
        RECT 379.950 427.950 382.050 430.050 ;
        RECT 358.950 413.250 360.750 414.150 ;
        RECT 361.950 412.950 364.050 415.050 ;
        RECT 364.950 412.950 367.050 415.050 ;
        RECT 367.950 412.950 370.050 415.050 ;
        RECT 358.950 409.950 361.050 412.050 ;
        RECT 362.250 410.850 364.050 411.750 ;
        RECT 364.950 410.250 367.050 411.150 ;
        RECT 367.950 410.850 370.050 411.750 ;
        RECT 355.950 394.950 358.050 397.050 ;
        RECT 352.950 388.950 355.050 391.050 ;
        RECT 337.950 385.950 340.050 388.050 ;
        RECT 343.950 385.950 346.050 388.050 ;
        RECT 349.950 385.950 352.050 388.050 ;
        RECT 337.950 384.450 340.050 385.050 ;
        RECT 335.400 383.400 340.050 384.450 ;
        RECT 325.950 375.300 328.050 377.400 ;
        RECT 331.950 376.950 334.050 379.050 ;
        RECT 326.250 371.700 327.450 375.300 ;
        RECT 325.950 369.600 328.050 371.700 ;
        RECT 331.950 370.950 334.050 373.050 ;
        RECT 305.400 365.400 309.450 366.450 ;
        RECT 305.400 340.050 306.450 365.400 ;
        RECT 313.950 364.950 316.050 367.050 ;
        RECT 322.950 364.950 325.050 367.050 ;
        RECT 325.950 349.950 328.050 352.050 ;
        RECT 307.950 344.250 310.050 345.150 ;
        RECT 326.400 343.050 327.450 349.950 ;
        RECT 332.400 343.050 333.450 370.950 ;
        RECT 335.400 352.050 336.450 383.400 ;
        RECT 337.950 382.950 340.050 383.400 ;
        RECT 341.250 383.250 343.050 384.150 ;
        RECT 343.950 383.850 346.050 384.750 ;
        RECT 346.950 383.250 349.050 384.150 ;
        RECT 349.950 382.950 352.050 385.050 ;
        RECT 337.950 380.850 339.750 381.750 ;
        RECT 340.950 379.950 343.050 382.050 ;
        RECT 346.950 379.950 349.050 382.050 ;
        RECT 337.950 376.950 340.050 379.050 ;
        RECT 334.950 349.950 337.050 352.050 ;
        RECT 311.250 341.250 312.750 342.150 ;
        RECT 313.950 340.950 316.050 343.050 ;
        RECT 317.250 341.250 319.050 342.150 ;
        RECT 319.950 340.950 322.050 343.050 ;
        RECT 322.950 341.250 324.750 342.150 ;
        RECT 325.950 340.950 328.050 343.050 ;
        RECT 329.250 341.250 330.750 342.150 ;
        RECT 331.950 340.950 334.050 343.050 ;
        RECT 335.250 341.250 337.050 342.150 ;
        RECT 304.950 337.950 307.050 340.050 ;
        RECT 307.950 337.950 310.050 340.050 ;
        RECT 310.950 337.950 313.050 340.050 ;
        RECT 314.250 338.850 315.750 339.750 ;
        RECT 316.950 337.950 319.050 340.050 ;
        RECT 301.950 319.950 304.050 322.050 ;
        RECT 298.950 316.950 301.050 319.050 ;
        RECT 289.950 313.950 292.050 316.050 ;
        RECT 295.950 313.950 298.050 316.050 ;
        RECT 286.950 301.950 289.050 304.050 ;
        RECT 290.400 289.050 291.450 313.950 ;
        RECT 296.400 310.050 297.450 313.950 ;
        RECT 292.950 308.250 294.750 309.150 ;
        RECT 295.950 307.950 298.050 310.050 ;
        RECT 299.400 307.050 300.450 316.950 ;
        RECT 301.950 307.950 304.050 310.050 ;
        RECT 292.950 304.950 295.050 307.050 ;
        RECT 296.250 305.850 297.750 306.750 ;
        RECT 298.950 304.950 301.050 307.050 ;
        RECT 302.250 305.850 304.050 306.750 ;
        RECT 298.950 302.850 301.050 303.750 ;
        RECT 286.950 286.950 289.050 289.050 ;
        RECT 289.950 286.950 292.050 289.050 ;
        RECT 298.950 286.950 301.050 289.050 ;
        RECT 287.400 285.450 288.450 286.950 ;
        RECT 287.400 284.400 291.450 285.450 ;
        RECT 286.950 280.950 289.050 283.050 ;
        RECT 283.950 269.250 286.050 270.150 ;
        RECT 283.950 265.950 286.050 268.050 ;
        RECT 284.400 265.050 285.450 265.950 ;
        RECT 287.400 265.050 288.450 280.950 ;
        RECT 290.400 271.050 291.450 284.400 ;
        RECT 295.950 283.950 298.050 286.050 ;
        RECT 296.400 271.050 297.450 283.950 ;
        RECT 299.400 271.050 300.450 286.950 ;
        RECT 305.400 283.050 306.450 337.950 ;
        RECT 308.400 334.050 309.450 337.950 ;
        RECT 311.400 334.050 312.450 337.950 ;
        RECT 307.950 331.950 310.050 334.050 ;
        RECT 310.950 331.950 313.050 334.050 ;
        RECT 317.400 319.050 318.450 337.950 ;
        RECT 320.400 336.450 321.450 340.950 ;
        RECT 322.950 337.950 325.050 340.050 ;
        RECT 326.250 338.850 327.750 339.750 ;
        RECT 328.950 337.950 331.050 340.050 ;
        RECT 332.250 338.850 333.750 339.750 ;
        RECT 334.950 337.950 337.050 340.050 ;
        RECT 320.400 335.400 324.450 336.450 ;
        RECT 307.950 316.950 310.050 319.050 ;
        RECT 316.950 316.950 319.050 319.050 ;
        RECT 308.400 313.050 309.450 316.950 ;
        RECT 317.400 316.050 318.450 316.950 ;
        RECT 310.950 313.950 313.050 316.050 ;
        RECT 316.950 313.950 319.050 316.050 ;
        RECT 323.400 313.050 324.450 335.400 ;
        RECT 338.400 334.050 339.450 376.950 ;
        RECT 341.400 373.050 342.450 379.950 ;
        RECT 347.400 379.050 348.450 379.950 ;
        RECT 346.950 376.950 349.050 379.050 ;
        RECT 350.400 376.050 351.450 382.950 ;
        RECT 349.950 373.950 352.050 376.050 ;
        RECT 340.950 370.950 343.050 373.050 ;
        RECT 346.950 364.950 349.050 367.050 ;
        RECT 340.950 340.950 343.050 343.050 ;
        RECT 340.950 338.850 343.050 339.750 ;
        RECT 343.950 338.250 346.050 339.150 ;
        RECT 343.950 334.950 346.050 337.050 ;
        RECT 337.950 331.950 340.050 334.050 ;
        RECT 344.400 331.050 345.450 334.950 ;
        RECT 343.950 328.950 346.050 331.050 ;
        RECT 343.950 325.950 346.050 328.050 ;
        RECT 344.400 322.050 345.450 325.950 ;
        RECT 331.950 319.950 334.050 322.050 ;
        RECT 343.950 319.950 346.050 322.050 ;
        RECT 332.400 313.050 333.450 319.950 ;
        RECT 340.950 316.950 343.050 319.050 ;
        RECT 307.950 310.950 310.050 313.050 ;
        RECT 311.250 311.850 312.750 312.750 ;
        RECT 313.950 310.950 316.050 313.050 ;
        RECT 316.950 310.950 319.050 313.050 ;
        RECT 320.250 311.250 321.750 312.150 ;
        RECT 322.950 310.950 325.050 313.050 ;
        RECT 331.950 310.950 334.050 313.050 ;
        RECT 307.950 308.850 310.050 309.750 ;
        RECT 310.950 307.950 313.050 310.050 ;
        RECT 313.950 308.850 316.050 309.750 ;
        RECT 316.950 308.850 318.750 309.750 ;
        RECT 319.950 307.950 322.050 310.050 ;
        RECT 323.250 308.850 324.750 309.750 ;
        RECT 325.950 309.450 328.050 310.050 ;
        RECT 325.950 308.400 330.450 309.450 ;
        RECT 331.950 308.850 334.050 309.750 ;
        RECT 337.950 308.850 340.050 309.750 ;
        RECT 325.950 307.950 328.050 308.400 ;
        RECT 311.400 286.050 312.450 307.950 ;
        RECT 329.400 307.050 330.450 308.400 ;
        RECT 325.950 305.850 328.050 306.750 ;
        RECT 328.950 304.950 331.050 307.050 ;
        RECT 319.950 301.950 322.050 304.050 ;
        RECT 310.950 283.950 313.050 286.050 ;
        RECT 304.950 280.950 307.050 283.050 ;
        RECT 289.950 270.450 292.050 271.050 ;
        RECT 289.950 269.400 294.450 270.450 ;
        RECT 289.950 268.950 292.050 269.400 ;
        RECT 289.950 266.850 292.050 267.750 ;
        RECT 280.950 262.950 283.050 265.050 ;
        RECT 283.950 262.950 286.050 265.050 ;
        RECT 286.950 262.950 289.050 265.050 ;
        RECT 277.950 256.950 280.050 259.050 ;
        RECT 274.950 247.950 277.050 250.050 ;
        RECT 278.400 244.050 279.450 256.950 ;
        RECT 289.950 253.950 292.050 256.050 ;
        RECT 280.950 247.950 283.050 250.050 ;
        RECT 286.950 247.950 289.050 250.050 ;
        RECT 268.950 241.950 271.050 244.050 ;
        RECT 277.950 241.950 280.050 244.050 ;
        RECT 278.400 241.050 279.450 241.950 ;
        RECT 250.950 238.950 253.050 241.050 ;
        RECT 253.950 238.950 256.050 241.050 ;
        RECT 257.250 239.250 258.750 240.150 ;
        RECT 259.950 238.950 262.050 241.050 ;
        RECT 262.950 238.950 265.050 241.050 ;
        RECT 265.950 238.950 268.050 241.050 ;
        RECT 271.950 238.950 274.050 241.050 ;
        RECT 275.250 239.250 276.750 240.150 ;
        RECT 277.950 238.950 280.050 241.050 ;
        RECT 251.400 238.050 252.450 238.950 ;
        RECT 250.950 235.950 253.050 238.050 ;
        RECT 254.250 236.850 255.750 237.750 ;
        RECT 256.950 235.950 259.050 238.050 ;
        RECT 260.250 236.850 262.050 237.750 ;
        RECT 250.950 233.850 253.050 234.750 ;
        RECT 257.400 229.050 258.450 235.950 ;
        RECT 256.950 226.950 259.050 229.050 ;
        RECT 259.950 223.950 262.050 226.050 ;
        RECT 253.950 220.950 256.050 223.050 ;
        RECT 250.950 205.950 253.050 208.050 ;
        RECT 247.950 199.950 250.050 202.050 ;
        RECT 232.950 197.250 234.750 198.150 ;
        RECT 235.950 196.950 238.050 199.050 ;
        RECT 239.250 197.250 240.750 198.150 ;
        RECT 241.950 196.950 244.050 199.050 ;
        RECT 245.250 197.250 247.050 198.150 ;
        RECT 247.950 196.950 250.050 199.050 ;
        RECT 232.950 193.950 235.050 196.050 ;
        RECT 236.250 194.850 237.750 195.750 ;
        RECT 238.950 193.950 241.050 196.050 ;
        RECT 242.250 194.850 243.750 195.750 ;
        RECT 244.950 193.950 247.050 196.050 ;
        RECT 233.400 184.050 234.450 193.950 ;
        RECT 232.950 181.950 235.050 184.050 ;
        RECT 239.400 181.050 240.450 193.950 ;
        RECT 245.400 190.050 246.450 193.950 ;
        RECT 244.950 187.950 247.050 190.050 ;
        RECT 248.400 187.050 249.450 196.950 ;
        RECT 247.950 184.950 250.050 187.050 ;
        RECT 238.950 178.950 241.050 181.050 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 238.950 175.950 241.050 178.050 ;
        RECT 235.950 169.950 238.050 172.050 ;
        RECT 232.950 163.950 235.050 166.050 ;
        RECT 236.400 163.050 237.450 169.950 ;
        RECT 239.400 166.050 240.450 175.950 ;
        RECT 242.400 169.050 243.450 178.950 ;
        RECT 244.950 175.950 247.050 178.050 ;
        RECT 241.950 166.950 244.050 169.050 ;
        RECT 238.950 163.950 241.050 166.050 ;
        RECT 242.250 164.250 244.050 165.150 ;
        RECT 232.950 161.850 234.750 162.750 ;
        RECT 235.950 160.950 238.050 163.050 ;
        RECT 239.250 161.850 240.750 162.750 ;
        RECT 241.950 160.950 244.050 163.050 ;
        RECT 235.950 158.850 238.050 159.750 ;
        RECT 238.950 157.950 241.050 160.050 ;
        RECT 239.400 151.050 240.450 157.950 ;
        RECT 238.950 148.950 241.050 151.050 ;
        RECT 241.950 142.950 244.050 145.050 ;
        RECT 229.950 136.950 232.050 139.050 ;
        RECT 235.950 136.950 238.050 139.050 ;
        RECT 229.950 133.950 232.050 136.050 ;
        RECT 230.400 130.050 231.450 133.950 ;
        RECT 229.950 127.950 232.050 130.050 ;
        RECT 230.400 127.050 231.450 127.950 ;
        RECT 229.950 124.950 232.050 127.050 ;
        RECT 229.950 122.850 232.050 123.750 ;
        RECT 232.950 122.250 235.050 123.150 ;
        RECT 220.950 118.950 223.050 121.050 ;
        RECT 226.950 118.950 229.050 121.050 ;
        RECT 232.950 120.450 235.050 121.050 ;
        RECT 236.400 120.450 237.450 136.950 ;
        RECT 242.400 127.050 243.450 142.950 ;
        RECT 245.400 133.050 246.450 175.950 ;
        RECT 251.400 172.050 252.450 205.950 ;
        RECT 254.400 205.050 255.450 220.950 ;
        RECT 260.400 214.050 261.450 223.950 ;
        RECT 259.950 211.950 262.050 214.050 ;
        RECT 253.950 202.950 256.050 205.050 ;
        RECT 259.950 199.950 262.050 202.050 ;
        RECT 260.400 199.050 261.450 199.950 ;
        RECT 263.400 199.050 264.450 238.950 ;
        RECT 266.400 205.050 267.450 238.950 ;
        RECT 268.950 235.950 271.050 238.050 ;
        RECT 272.250 236.850 273.750 237.750 ;
        RECT 274.950 235.950 277.050 238.050 ;
        RECT 278.250 236.850 280.050 237.750 ;
        RECT 275.400 235.050 276.450 235.950 ;
        RECT 268.950 233.850 271.050 234.750 ;
        RECT 274.950 232.950 277.050 235.050 ;
        RECT 281.400 226.050 282.450 247.950 ;
        RECT 287.400 241.050 288.450 247.950 ;
        RECT 283.950 238.950 286.050 241.050 ;
        RECT 286.950 238.950 289.050 241.050 ;
        RECT 290.400 240.450 291.450 253.950 ;
        RECT 293.400 243.450 294.450 269.400 ;
        RECT 295.950 268.950 298.050 271.050 ;
        RECT 298.950 268.950 301.050 271.050 ;
        RECT 302.250 269.250 304.050 270.150 ;
        RECT 304.950 268.950 307.050 271.050 ;
        RECT 310.950 269.250 312.750 270.150 ;
        RECT 313.950 268.950 316.050 271.050 ;
        RECT 316.950 269.250 319.050 270.150 ;
        RECT 295.950 266.850 298.050 267.750 ;
        RECT 298.950 266.850 300.750 267.750 ;
        RECT 301.950 265.950 304.050 268.050 ;
        RECT 302.400 256.050 303.450 265.950 ;
        RECT 301.950 253.950 304.050 256.050 ;
        RECT 298.950 244.950 301.050 247.050 ;
        RECT 293.400 242.400 297.450 243.450 ;
        RECT 292.950 240.450 295.050 241.050 ;
        RECT 290.400 239.400 295.050 240.450 ;
        RECT 292.950 238.950 295.050 239.400 ;
        RECT 283.950 236.850 286.050 237.750 ;
        RECT 286.950 236.250 289.050 237.150 ;
        RECT 289.950 235.950 292.050 238.050 ;
        RECT 292.950 236.850 295.050 237.750 ;
        RECT 286.950 232.950 289.050 235.050 ;
        RECT 287.400 232.050 288.450 232.950 ;
        RECT 286.950 229.950 289.050 232.050 ;
        RECT 280.950 223.950 283.050 226.050 ;
        RECT 274.950 217.950 277.050 220.050 ;
        RECT 275.400 211.050 276.450 217.950 ;
        RECT 274.950 208.950 277.050 211.050 ;
        RECT 268.950 205.950 271.050 208.050 ;
        RECT 265.950 202.950 268.050 205.050 ;
        RECT 269.400 202.050 270.450 205.950 ;
        RECT 274.950 203.250 277.050 204.150 ;
        RECT 281.400 202.050 282.450 223.950 ;
        RECT 286.950 202.950 289.050 205.050 ;
        RECT 287.400 202.050 288.450 202.950 ;
        RECT 265.950 199.950 268.050 202.050 ;
        RECT 268.950 199.950 271.050 202.050 ;
        RECT 272.250 200.250 273.750 201.150 ;
        RECT 274.950 199.950 277.050 202.050 ;
        RECT 278.250 200.250 280.050 201.150 ;
        RECT 280.950 199.950 283.050 202.050 ;
        RECT 284.250 200.250 285.750 201.150 ;
        RECT 286.950 199.950 289.050 202.050 ;
        RECT 253.950 197.250 255.750 198.150 ;
        RECT 256.950 196.950 259.050 199.050 ;
        RECT 259.950 196.950 262.050 199.050 ;
        RECT 262.950 196.950 265.050 199.050 ;
        RECT 253.950 193.950 256.050 196.050 ;
        RECT 257.250 194.850 259.050 195.750 ;
        RECT 259.950 194.250 262.050 195.150 ;
        RECT 262.950 194.850 265.050 195.750 ;
        RECT 250.950 169.950 253.050 172.050 ;
        RECT 254.400 169.050 255.450 193.950 ;
        RECT 259.950 190.950 262.050 193.050 ;
        RECT 262.950 190.950 265.050 193.050 ;
        RECT 263.400 187.050 264.450 190.950 ;
        RECT 262.950 184.950 265.050 187.050 ;
        RECT 266.400 181.050 267.450 199.950 ;
        RECT 275.400 199.050 276.450 199.950 ;
        RECT 268.950 197.850 270.750 198.750 ;
        RECT 271.950 196.950 274.050 199.050 ;
        RECT 274.950 196.950 277.050 199.050 ;
        RECT 277.950 196.950 280.050 199.050 ;
        RECT 280.950 197.850 282.750 198.750 ;
        RECT 283.950 196.950 286.050 199.050 ;
        RECT 287.250 197.850 289.050 198.750 ;
        RECT 272.400 196.050 273.450 196.950 ;
        RECT 278.400 196.050 279.450 196.950 ;
        RECT 284.400 196.050 285.450 196.950 ;
        RECT 271.950 193.950 274.050 196.050 ;
        RECT 277.950 193.950 280.050 196.050 ;
        RECT 283.950 193.950 286.050 196.050 ;
        RECT 278.400 193.050 279.450 193.950 ;
        RECT 277.950 190.950 280.050 193.050 ;
        RECT 280.950 190.950 283.050 193.050 ;
        RECT 268.950 184.950 271.050 187.050 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 256.950 169.950 259.050 172.050 ;
        RECT 259.950 169.950 262.050 172.050 ;
        RECT 265.950 169.950 268.050 172.050 ;
        RECT 247.950 166.950 250.050 169.050 ;
        RECT 253.950 166.950 256.050 169.050 ;
        RECT 248.400 145.050 249.450 166.950 ;
        RECT 253.950 165.450 256.050 166.050 ;
        RECT 257.400 165.450 258.450 169.950 ;
        RECT 260.400 166.050 261.450 169.950 ;
        RECT 269.400 169.050 270.450 184.950 ;
        RECT 271.950 181.950 274.050 184.050 ;
        RECT 274.950 181.950 277.050 184.050 ;
        RECT 262.950 166.950 265.050 169.050 ;
        RECT 266.250 167.850 267.750 168.750 ;
        RECT 268.950 166.950 271.050 169.050 ;
        RECT 250.950 164.250 252.750 165.150 ;
        RECT 253.950 164.400 258.450 165.450 ;
        RECT 253.950 163.950 256.050 164.400 ;
        RECT 259.950 163.950 262.050 166.050 ;
        RECT 262.950 164.850 265.050 165.750 ;
        RECT 265.950 163.950 268.050 166.050 ;
        RECT 268.950 164.850 271.050 165.750 ;
        RECT 250.950 160.950 253.050 163.050 ;
        RECT 254.250 161.850 255.750 162.750 ;
        RECT 256.950 160.950 259.050 163.050 ;
        RECT 260.250 161.850 262.050 162.750 ;
        RECT 247.950 142.950 250.050 145.050 ;
        RECT 247.950 136.950 250.050 139.050 ;
        RECT 244.950 130.950 247.050 133.050 ;
        RECT 248.400 127.050 249.450 136.950 ;
        RECT 251.400 133.050 252.450 160.950 ;
        RECT 256.950 158.850 259.050 159.750 ;
        RECT 266.400 139.050 267.450 163.950 ;
        RECT 272.400 145.050 273.450 181.950 ;
        RECT 275.400 165.450 276.450 181.950 ;
        RECT 281.400 175.050 282.450 190.950 ;
        RECT 283.950 184.950 286.050 187.050 ;
        RECT 280.950 172.950 283.050 175.050 ;
        RECT 281.400 172.050 282.450 172.950 ;
        RECT 280.950 169.950 283.050 172.050 ;
        RECT 277.950 167.250 280.050 168.150 ;
        RECT 280.950 167.850 283.050 168.750 ;
        RECT 277.950 165.450 280.050 166.050 ;
        RECT 275.400 164.400 280.050 165.450 ;
        RECT 271.950 142.950 274.050 145.050 ;
        RECT 275.400 142.050 276.450 164.400 ;
        RECT 277.950 163.950 280.050 164.400 ;
        RECT 280.950 163.950 283.050 166.050 ;
        RECT 277.950 148.950 280.050 151.050 ;
        RECT 274.950 139.950 277.050 142.050 ;
        RECT 265.950 136.950 268.050 139.050 ;
        RECT 268.950 133.950 271.050 136.050 ;
        RECT 250.950 130.950 253.050 133.050 ;
        RECT 253.950 130.950 256.050 133.050 ;
        RECT 262.950 130.950 265.050 133.050 ;
        RECT 238.950 125.250 240.750 126.150 ;
        RECT 241.950 124.950 244.050 127.050 ;
        RECT 245.250 125.250 246.750 126.150 ;
        RECT 247.950 124.950 250.050 127.050 ;
        RECT 251.250 125.250 253.050 126.150 ;
        RECT 238.950 121.950 241.050 124.050 ;
        RECT 242.250 122.850 243.750 123.750 ;
        RECT 244.950 121.950 247.050 124.050 ;
        RECT 248.250 122.850 249.750 123.750 ;
        RECT 250.950 121.950 253.050 124.050 ;
        RECT 232.950 119.400 237.450 120.450 ;
        RECT 232.950 118.950 235.050 119.400 ;
        RECT 238.950 118.950 241.050 121.050 ;
        RECT 235.950 112.950 238.050 115.050 ;
        RECT 206.400 110.400 210.450 111.450 ;
        RECT 206.400 100.050 207.450 110.400 ;
        RECT 211.950 109.950 214.050 112.050 ;
        RECT 220.950 109.950 223.050 112.050 ;
        RECT 202.950 97.950 205.050 100.050 ;
        RECT 205.950 97.950 208.050 100.050 ;
        RECT 202.950 95.850 205.050 96.750 ;
        RECT 205.950 95.250 208.050 96.150 ;
        RECT 205.950 91.950 208.050 94.050 ;
        RECT 211.950 92.250 213.750 93.150 ;
        RECT 214.950 91.950 217.050 94.050 ;
        RECT 218.250 92.250 220.050 93.150 ;
        RECT 211.950 88.950 214.050 91.050 ;
        RECT 215.250 89.850 216.750 90.750 ;
        RECT 217.950 90.450 220.050 91.050 ;
        RECT 221.400 90.450 222.450 109.950 ;
        RECT 223.950 94.950 226.050 97.050 ;
        RECT 224.400 94.050 225.450 94.950 ;
        RECT 223.950 91.950 226.050 94.050 ;
        RECT 226.950 91.950 229.050 94.050 ;
        RECT 229.950 91.950 232.050 94.050 ;
        RECT 233.250 92.250 235.050 93.150 ;
        RECT 227.400 91.050 228.450 91.950 ;
        RECT 236.400 91.050 237.450 112.950 ;
        RECT 217.950 89.400 222.450 90.450 ;
        RECT 223.950 89.850 225.750 90.750 ;
        RECT 217.950 88.950 220.050 89.400 ;
        RECT 226.950 88.950 229.050 91.050 ;
        RECT 230.250 89.850 231.750 90.750 ;
        RECT 232.950 88.950 235.050 91.050 ;
        RECT 235.950 88.950 238.050 91.050 ;
        RECT 199.950 85.950 202.050 88.050 ;
        RECT 212.400 85.050 213.450 88.950 ;
        RECT 220.950 85.950 223.050 88.050 ;
        RECT 226.950 86.850 229.050 87.750 ;
        RECT 211.950 82.950 214.050 85.050 ;
        RECT 214.950 59.250 217.050 60.150 ;
        RECT 221.400 58.050 222.450 85.950 ;
        RECT 226.950 67.950 229.050 70.050 ;
        RECT 227.400 58.050 228.450 67.950 ;
        RECT 233.400 58.050 234.450 88.950 ;
        RECT 239.400 88.050 240.450 118.950 ;
        RECT 245.400 112.050 246.450 121.950 ;
        RECT 251.400 121.050 252.450 121.950 ;
        RECT 250.950 118.950 253.050 121.050 ;
        RECT 250.950 115.950 253.050 118.050 ;
        RECT 241.950 109.950 244.050 112.050 ;
        RECT 244.950 109.950 247.050 112.050 ;
        RECT 242.400 109.050 243.450 109.950 ;
        RECT 241.950 106.950 244.050 109.050 ;
        RECT 242.400 97.050 243.450 106.950 ;
        RECT 244.950 103.950 247.050 106.050 ;
        RECT 245.400 100.050 246.450 103.950 ;
        RECT 244.950 97.950 247.050 100.050 ;
        RECT 247.950 97.950 250.050 100.050 ;
        RECT 248.400 97.050 249.450 97.950 ;
        RECT 241.950 94.950 244.050 97.050 ;
        RECT 245.250 95.850 246.750 96.750 ;
        RECT 247.950 94.950 250.050 97.050 ;
        RECT 241.950 92.850 244.050 93.750 ;
        RECT 247.950 92.850 250.050 93.750 ;
        RECT 238.950 85.950 241.050 88.050 ;
        RECT 251.400 70.050 252.450 115.950 ;
        RECT 254.400 103.050 255.450 130.950 ;
        RECT 263.400 130.050 264.450 130.950 ;
        RECT 256.950 127.950 259.050 130.050 ;
        RECT 260.250 128.250 261.750 129.150 ;
        RECT 262.950 127.950 265.050 130.050 ;
        RECT 265.950 127.950 268.050 130.050 ;
        RECT 256.950 125.850 258.750 126.750 ;
        RECT 259.950 124.950 262.050 127.050 ;
        RECT 263.250 125.850 265.050 126.750 ;
        RECT 260.400 115.050 261.450 124.950 ;
        RECT 266.400 121.050 267.450 127.950 ;
        RECT 269.400 127.050 270.450 133.950 ;
        RECT 278.400 129.450 279.450 148.950 ;
        RECT 275.400 128.400 279.450 129.450 ;
        RECT 275.400 127.050 276.450 128.400 ;
        RECT 268.950 124.950 271.050 127.050 ;
        RECT 274.950 124.950 277.050 127.050 ;
        RECT 278.250 125.250 280.050 126.150 ;
        RECT 268.950 122.850 271.050 123.750 ;
        RECT 271.950 122.250 274.050 123.150 ;
        RECT 274.950 122.850 276.750 123.750 ;
        RECT 277.950 121.950 280.050 124.050 ;
        RECT 265.950 118.950 268.050 121.050 ;
        RECT 271.950 118.950 274.050 121.050 ;
        RECT 259.950 112.950 262.050 115.050 ;
        RECT 277.950 112.950 280.050 115.050 ;
        RECT 265.950 109.950 268.050 112.050 ;
        RECT 271.950 109.950 274.050 112.050 ;
        RECT 262.950 106.950 265.050 109.050 ;
        RECT 263.400 106.050 264.450 106.950 ;
        RECT 262.950 103.950 265.050 106.050 ;
        RECT 253.950 100.950 256.050 103.050 ;
        RECT 254.400 100.050 255.450 100.950 ;
        RECT 263.400 100.050 264.450 103.950 ;
        RECT 253.950 97.950 256.050 100.050 ;
        RECT 262.950 97.950 265.050 100.050 ;
        RECT 253.950 95.250 256.050 96.150 ;
        RECT 256.950 94.950 259.050 97.050 ;
        RECT 259.950 94.950 262.050 97.050 ;
        RECT 263.250 95.850 265.050 96.750 ;
        RECT 253.950 91.950 256.050 94.050 ;
        RECT 257.400 85.050 258.450 94.950 ;
        RECT 266.400 94.050 267.450 109.950 ;
        RECT 272.400 94.050 273.450 109.950 ;
        RECT 278.400 109.050 279.450 112.950 ;
        RECT 277.950 106.950 280.050 109.050 ;
        RECT 274.950 100.950 277.050 103.050 ;
        RECT 278.400 102.450 279.450 106.950 ;
        RECT 281.400 106.050 282.450 163.950 ;
        RECT 284.400 157.050 285.450 184.950 ;
        RECT 290.400 181.050 291.450 235.950 ;
        RECT 296.400 220.050 297.450 242.400 ;
        RECT 299.400 241.050 300.450 244.950 ;
        RECT 302.400 244.050 303.450 253.950 ;
        RECT 305.400 247.050 306.450 268.950 ;
        RECT 310.950 265.950 313.050 268.050 ;
        RECT 314.250 266.850 316.050 267.750 ;
        RECT 316.950 265.950 319.050 268.050 ;
        RECT 311.400 250.050 312.450 265.950 ;
        RECT 317.400 265.050 318.450 265.950 ;
        RECT 316.950 262.950 319.050 265.050 ;
        RECT 320.400 261.450 321.450 301.950 ;
        RECT 325.950 283.950 328.050 286.050 ;
        RECT 326.400 271.050 327.450 283.950 ;
        RECT 322.950 269.250 325.050 270.150 ;
        RECT 325.950 268.950 328.050 271.050 ;
        RECT 322.950 265.950 325.050 268.050 ;
        RECT 317.400 260.400 321.450 261.450 ;
        RECT 310.950 247.950 313.050 250.050 ;
        RECT 304.950 244.950 307.050 247.050 ;
        RECT 301.950 241.950 304.050 244.050 ;
        RECT 298.950 238.950 301.050 241.050 ;
        RECT 302.250 239.250 303.750 240.150 ;
        RECT 304.950 238.950 307.050 241.050 ;
        RECT 308.250 239.250 309.750 240.150 ;
        RECT 310.950 238.950 313.050 241.050 ;
        RECT 298.950 236.850 300.750 237.750 ;
        RECT 301.950 235.950 304.050 238.050 ;
        RECT 305.250 236.850 306.750 237.750 ;
        RECT 307.950 235.950 310.050 238.050 ;
        RECT 311.250 236.850 313.050 237.750 ;
        RECT 302.400 232.050 303.450 235.950 ;
        RECT 301.950 229.950 304.050 232.050 ;
        RECT 308.400 226.050 309.450 235.950 ;
        RECT 317.400 235.050 318.450 260.400 ;
        RECT 323.400 250.050 324.450 265.950 ;
        RECT 329.400 265.050 330.450 304.950 ;
        RECT 341.400 280.050 342.450 316.950 ;
        RECT 344.400 310.050 345.450 319.950 ;
        RECT 347.400 319.050 348.450 364.950 ;
        RECT 353.400 358.050 354.450 388.950 ;
        RECT 359.400 388.050 360.450 409.950 ;
        RECT 364.950 406.950 367.050 409.050 ;
        RECT 365.400 400.050 366.450 406.950 ;
        RECT 364.950 397.950 367.050 400.050 ;
        RECT 361.950 391.950 364.050 394.050 ;
        RECT 358.950 385.950 361.050 388.050 ;
        RECT 362.400 385.050 363.450 391.950 ;
        RECT 355.950 382.950 358.050 385.050 ;
        RECT 359.250 383.250 360.750 384.150 ;
        RECT 361.950 382.950 364.050 385.050 ;
        RECT 365.250 383.250 366.750 384.150 ;
        RECT 367.950 382.950 370.050 385.050 ;
        RECT 355.950 380.850 357.750 381.750 ;
        RECT 358.950 379.950 361.050 382.050 ;
        RECT 362.250 380.850 363.750 381.750 ;
        RECT 364.950 379.950 367.050 382.050 ;
        RECT 368.250 380.850 370.050 381.750 ;
        RECT 365.400 376.050 366.450 379.950 ;
        RECT 364.950 373.950 367.050 376.050 ;
        RECT 365.400 373.050 366.450 373.950 ;
        RECT 364.950 370.950 367.050 373.050 ;
        RECT 367.950 370.950 370.050 373.050 ;
        RECT 352.950 355.950 355.050 358.050 ;
        RECT 361.950 355.950 364.050 358.050 ;
        RECT 352.950 350.400 355.050 352.500 ;
        RECT 353.400 333.600 354.600 350.400 ;
        RECT 362.400 349.050 363.450 355.950 ;
        RECT 361.950 346.950 364.050 349.050 ;
        RECT 355.950 343.950 358.050 346.050 ;
        RECT 356.400 339.450 357.450 343.950 ;
        RECT 358.950 341.250 361.050 342.150 ;
        RECT 358.950 339.450 361.050 340.050 ;
        RECT 356.400 338.400 361.050 339.450 ;
        RECT 362.400 339.450 363.450 346.950 ;
        RECT 364.950 341.250 367.050 342.150 ;
        RECT 364.950 339.450 367.050 340.050 ;
        RECT 362.400 338.400 367.050 339.450 ;
        RECT 358.950 337.950 361.050 338.400 ;
        RECT 364.950 337.950 367.050 338.400 ;
        RECT 352.950 331.500 355.050 333.600 ;
        RECT 368.400 328.050 369.450 370.950 ;
        RECT 367.950 325.950 370.050 328.050 ;
        RECT 346.950 316.950 349.050 319.050 ;
        RECT 371.400 318.450 372.450 427.950 ;
        RECT 373.950 416.250 376.050 417.150 ;
        RECT 380.400 415.050 381.450 427.950 ;
        RECT 386.400 424.050 387.450 445.950 ;
        RECT 392.400 444.600 393.600 461.400 ;
        RECT 391.950 442.500 394.050 444.600 ;
        RECT 385.950 421.950 388.050 424.050 ;
        RECT 385.950 418.950 388.050 421.050 ;
        RECT 373.950 412.950 376.050 415.050 ;
        RECT 377.250 413.250 378.750 414.150 ;
        RECT 379.950 412.950 382.050 415.050 ;
        RECT 383.250 413.250 385.050 414.150 ;
        RECT 374.400 406.050 375.450 412.950 ;
        RECT 376.950 409.950 379.050 412.050 ;
        RECT 380.250 410.850 381.750 411.750 ;
        RECT 382.950 409.950 385.050 412.050 ;
        RECT 373.950 403.950 376.050 406.050 ;
        RECT 386.400 403.050 387.450 418.950 ;
        RECT 388.950 415.950 391.050 418.050 ;
        RECT 391.950 415.950 394.050 418.050 ;
        RECT 389.400 412.050 390.450 415.950 ;
        RECT 392.400 415.050 393.450 415.950 ;
        RECT 391.950 412.950 394.050 415.050 ;
        RECT 388.950 409.950 391.050 412.050 ;
        RECT 391.950 410.850 394.050 411.750 ;
        RECT 391.950 406.950 394.050 409.050 ;
        RECT 379.950 400.950 382.050 403.050 ;
        RECT 385.950 400.950 388.050 403.050 ;
        RECT 376.950 385.950 379.050 388.050 ;
        RECT 373.950 383.250 376.050 384.150 ;
        RECT 376.950 383.850 379.050 384.750 ;
        RECT 373.950 379.950 376.050 382.050 ;
        RECT 380.400 376.050 381.450 400.950 ;
        RECT 385.950 389.400 388.050 391.500 ;
        RECT 382.950 386.250 385.050 387.150 ;
        RECT 382.950 382.950 385.050 385.050 ;
        RECT 386.550 377.400 387.750 389.400 ;
        RECT 388.950 382.950 391.050 385.050 ;
        RECT 379.950 373.950 382.050 376.050 ;
        RECT 385.950 375.300 388.050 377.400 ;
        RECT 386.550 371.700 387.750 375.300 ;
        RECT 385.950 369.600 388.050 371.700 ;
        RECT 373.950 351.300 376.050 353.400 ;
        RECT 374.250 347.700 375.450 351.300 ;
        RECT 373.950 345.600 376.050 347.700 ;
        RECT 382.950 346.950 385.050 349.050 ;
        RECT 374.250 333.600 375.450 345.600 ;
        RECT 376.950 339.450 379.050 340.050 ;
        RECT 383.400 339.450 384.450 346.950 ;
        RECT 385.950 341.250 388.050 342.150 ;
        RECT 385.950 339.450 388.050 340.050 ;
        RECT 376.950 338.400 381.450 339.450 ;
        RECT 383.400 338.400 388.050 339.450 ;
        RECT 376.950 337.950 379.050 338.400 ;
        RECT 376.950 335.850 379.050 336.750 ;
        RECT 373.950 331.500 376.050 333.600 ;
        RECT 380.400 331.050 381.450 338.400 ;
        RECT 385.950 337.950 388.050 338.400 ;
        RECT 386.400 334.050 387.450 337.950 ;
        RECT 382.950 331.950 385.050 334.050 ;
        RECT 385.950 331.950 388.050 334.050 ;
        RECT 379.950 328.950 382.050 331.050 ;
        RECT 379.950 325.950 382.050 328.050 ;
        RECT 368.400 317.400 372.450 318.450 ;
        RECT 349.950 310.950 352.050 313.050 ;
        RECT 355.950 310.950 358.050 313.050 ;
        RECT 361.950 310.950 364.050 313.050 ;
        RECT 350.400 310.050 351.450 310.950 ;
        RECT 343.950 307.950 346.050 310.050 ;
        RECT 346.950 308.250 348.750 309.150 ;
        RECT 349.950 307.950 352.050 310.050 ;
        RECT 353.250 308.250 355.050 309.150 ;
        RECT 346.950 304.950 349.050 307.050 ;
        RECT 350.250 305.850 351.750 306.750 ;
        RECT 352.950 304.950 355.050 307.050 ;
        RECT 356.400 306.450 357.450 310.950 ;
        RECT 362.400 310.050 363.450 310.950 ;
        RECT 358.950 308.250 360.750 309.150 ;
        RECT 361.950 307.950 364.050 310.050 ;
        RECT 365.250 308.250 367.050 309.150 ;
        RECT 358.950 306.450 361.050 307.050 ;
        RECT 356.400 305.400 361.050 306.450 ;
        RECT 362.250 305.850 363.750 306.750 ;
        RECT 358.950 304.950 361.050 305.400 ;
        RECT 364.950 304.950 367.050 307.050 ;
        RECT 343.950 301.950 346.050 304.050 ;
        RECT 340.950 277.950 343.050 280.050 ;
        RECT 337.950 275.250 340.050 276.150 ;
        RECT 331.950 271.950 334.050 274.050 ;
        RECT 335.250 272.250 336.750 273.150 ;
        RECT 337.950 271.950 340.050 274.050 ;
        RECT 341.250 272.250 343.050 273.150 ;
        RECT 338.400 271.050 339.450 271.950 ;
        RECT 331.950 269.850 333.750 270.750 ;
        RECT 334.950 268.950 337.050 271.050 ;
        RECT 337.950 268.950 340.050 271.050 ;
        RECT 340.950 268.950 343.050 271.050 ;
        RECT 334.950 267.450 337.050 268.050 ;
        RECT 337.950 267.450 340.050 268.050 ;
        RECT 334.950 266.400 340.050 267.450 ;
        RECT 334.950 265.950 337.050 266.400 ;
        RECT 337.950 265.950 340.050 266.400 ;
        RECT 328.950 262.950 331.050 265.050 ;
        RECT 341.400 259.050 342.450 268.950 ;
        RECT 340.950 256.950 343.050 259.050 ;
        RECT 344.400 256.050 345.450 301.950 ;
        RECT 347.400 277.050 348.450 304.950 ;
        RECT 353.400 304.050 354.450 304.950 ;
        RECT 352.950 301.950 355.050 304.050 ;
        RECT 352.950 292.950 355.050 295.050 ;
        RECT 353.400 277.050 354.450 292.950 ;
        RECT 368.400 289.050 369.450 317.400 ;
        RECT 380.400 313.050 381.450 325.950 ;
        RECT 370.950 310.950 373.050 313.050 ;
        RECT 379.950 310.950 382.050 313.050 ;
        RECT 370.950 308.850 373.050 309.750 ;
        RECT 376.950 308.250 379.050 309.150 ;
        RECT 379.950 308.850 382.050 309.750 ;
        RECT 376.950 304.950 379.050 307.050 ;
        RECT 367.950 286.950 370.050 289.050 ;
        RECT 377.400 283.050 378.450 304.950 ;
        RECT 379.950 298.950 382.050 301.050 ;
        RECT 380.400 295.050 381.450 298.950 ;
        RECT 379.950 292.950 382.050 295.050 ;
        RECT 379.950 283.950 382.050 286.050 ;
        RECT 355.950 280.950 358.050 283.050 ;
        RECT 370.950 280.950 373.050 283.050 ;
        RECT 376.950 280.950 379.050 283.050 ;
        RECT 346.950 274.950 349.050 277.050 ;
        RECT 352.950 274.950 355.050 277.050 ;
        RECT 346.950 271.950 349.050 274.050 ;
        RECT 352.950 273.450 355.050 274.050 ;
        RECT 356.400 273.450 357.450 280.950 ;
        RECT 350.250 272.250 351.750 273.150 ;
        RECT 352.950 272.400 357.450 273.450 ;
        RECT 352.950 271.950 355.050 272.400 ;
        RECT 346.950 269.850 348.750 270.750 ;
        RECT 349.950 268.950 352.050 271.050 ;
        RECT 353.250 269.850 355.050 270.750 ;
        RECT 350.400 264.450 351.450 268.950 ;
        RECT 352.950 264.450 355.050 265.050 ;
        RECT 350.400 263.400 355.050 264.450 ;
        RECT 352.950 262.950 355.050 263.400 ;
        RECT 352.950 259.950 355.050 262.050 ;
        RECT 340.950 253.950 343.050 256.050 ;
        RECT 343.950 253.950 346.050 256.050 ;
        RECT 322.950 247.950 325.050 250.050 ;
        RECT 328.950 247.950 331.050 250.050 ;
        RECT 319.950 244.950 322.050 247.050 ;
        RECT 320.400 241.050 321.450 244.950 ;
        RECT 323.400 241.050 324.450 247.950 ;
        RECT 325.950 241.950 328.050 244.050 ;
        RECT 326.400 241.050 327.450 241.950 ;
        RECT 329.400 241.050 330.450 247.950 ;
        RECT 341.400 247.050 342.450 253.950 ;
        RECT 331.950 244.950 334.050 247.050 ;
        RECT 340.950 244.950 343.050 247.050 ;
        RECT 319.950 238.950 322.050 241.050 ;
        RECT 322.950 238.950 325.050 241.050 ;
        RECT 325.950 238.950 328.050 241.050 ;
        RECT 328.950 238.950 331.050 241.050 ;
        RECT 319.950 236.850 322.050 237.750 ;
        RECT 325.950 236.850 328.050 237.750 ;
        RECT 328.950 236.850 331.050 237.750 ;
        RECT 310.950 232.950 313.050 235.050 ;
        RECT 316.950 232.950 319.050 235.050 ;
        RECT 307.950 223.950 310.050 226.050 ;
        RECT 307.950 220.950 310.050 223.050 ;
        RECT 295.950 217.950 298.050 220.050 ;
        RECT 304.950 211.950 307.050 214.050 ;
        RECT 292.950 202.950 295.050 205.050 ;
        RECT 289.950 178.950 292.050 181.050 ;
        RECT 293.400 178.050 294.450 202.950 ;
        RECT 295.950 199.950 298.050 202.050 ;
        RECT 299.250 200.250 300.750 201.150 ;
        RECT 301.950 199.950 304.050 202.050 ;
        RECT 295.950 197.850 297.750 198.750 ;
        RECT 298.950 196.950 301.050 199.050 ;
        RECT 302.250 197.850 304.050 198.750 ;
        RECT 292.950 175.950 295.050 178.050 ;
        RECT 289.950 172.950 292.050 175.050 ;
        RECT 290.400 166.050 291.450 172.950 ;
        RECT 299.400 172.050 300.450 196.950 ;
        RECT 305.400 190.050 306.450 211.950 ;
        RECT 308.400 211.050 309.450 220.950 ;
        RECT 311.400 214.050 312.450 232.950 ;
        RECT 319.950 229.950 322.050 232.050 ;
        RECT 316.950 228.450 319.050 229.050 ;
        RECT 320.400 228.450 321.450 229.950 ;
        RECT 316.950 227.400 321.450 228.450 ;
        RECT 316.950 226.950 319.050 227.400 ;
        RECT 322.950 223.950 325.050 226.050 ;
        RECT 310.950 211.950 313.050 214.050 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 307.950 208.950 310.050 211.050 ;
        RECT 310.950 208.950 313.050 211.050 ;
        RECT 308.400 202.050 309.450 208.950 ;
        RECT 307.950 199.950 310.050 202.050 ;
        RECT 307.950 197.250 310.050 198.150 ;
        RECT 307.950 193.950 310.050 196.050 ;
        RECT 308.400 193.050 309.450 193.950 ;
        RECT 307.950 190.950 310.050 193.050 ;
        RECT 304.950 187.950 307.050 190.050 ;
        RECT 311.400 184.050 312.450 208.950 ;
        RECT 313.950 205.950 316.050 208.050 ;
        RECT 314.400 202.050 315.450 205.950 ;
        RECT 320.400 202.050 321.450 211.950 ;
        RECT 313.950 199.950 316.050 202.050 ;
        RECT 319.950 199.950 322.050 202.050 ;
        RECT 313.950 197.850 316.050 198.750 ;
        RECT 316.950 197.250 319.050 198.150 ;
        RECT 319.950 196.950 322.050 199.050 ;
        RECT 320.400 196.050 321.450 196.950 ;
        RECT 316.950 193.950 319.050 196.050 ;
        RECT 319.950 193.950 322.050 196.050 ;
        RECT 319.950 190.950 322.050 193.050 ;
        RECT 310.950 181.950 313.050 184.050 ;
        RECT 301.950 178.950 304.050 181.050 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 302.400 172.050 303.450 178.950 ;
        RECT 298.950 169.950 301.050 172.050 ;
        RECT 301.950 169.950 304.050 172.050 ;
        RECT 299.400 169.050 300.450 169.950 ;
        RECT 292.950 166.950 295.050 169.050 ;
        RECT 296.250 167.250 297.750 168.150 ;
        RECT 298.950 166.950 301.050 169.050 ;
        RECT 301.950 167.850 304.050 168.750 ;
        RECT 304.950 167.250 307.050 168.150 ;
        RECT 308.400 166.050 309.450 178.950 ;
        RECT 316.950 175.950 319.050 178.050 ;
        RECT 317.400 172.050 318.450 175.950 ;
        RECT 316.950 169.950 319.050 172.050 ;
        RECT 320.400 169.050 321.450 190.950 ;
        RECT 323.400 184.050 324.450 223.950 ;
        RECT 332.400 208.050 333.450 244.950 ;
        RECT 337.950 240.450 340.050 241.050 ;
        RECT 337.950 239.400 342.450 240.450 ;
        RECT 337.950 238.950 340.050 239.400 ;
        RECT 334.950 236.250 337.050 237.150 ;
        RECT 337.950 236.850 340.050 237.750 ;
        RECT 334.950 232.950 337.050 235.050 ;
        RECT 335.400 229.050 336.450 232.950 ;
        RECT 334.950 226.950 337.050 229.050 ;
        RECT 331.950 205.950 334.050 208.050 ;
        RECT 341.400 205.050 342.450 239.400 ;
        RECT 344.400 226.050 345.450 253.950 ;
        RECT 353.400 244.050 354.450 259.950 ;
        RECT 356.400 259.050 357.450 272.400 ;
        RECT 358.950 271.950 361.050 274.050 ;
        RECT 355.950 256.950 358.050 259.050 ;
        RECT 359.400 247.050 360.450 271.950 ;
        RECT 371.400 271.050 372.450 280.950 ;
        RECT 373.950 277.950 376.050 280.050 ;
        RECT 374.400 274.050 375.450 277.950 ;
        RECT 380.400 274.050 381.450 283.950 ;
        RECT 373.950 271.950 376.050 274.050 ;
        RECT 377.250 272.250 378.750 273.150 ;
        RECT 379.950 271.950 382.050 274.050 ;
        RECT 361.950 269.250 363.750 270.150 ;
        RECT 364.950 268.950 367.050 271.050 ;
        RECT 370.950 268.950 373.050 271.050 ;
        RECT 373.950 269.850 375.750 270.750 ;
        RECT 376.950 268.950 379.050 271.050 ;
        RECT 380.250 269.850 382.050 270.750 ;
        RECT 361.950 265.950 364.050 268.050 ;
        RECT 365.250 266.850 367.050 267.750 ;
        RECT 367.950 266.250 370.050 267.150 ;
        RECT 370.950 266.850 373.050 267.750 ;
        RECT 383.400 267.450 384.450 331.950 ;
        RECT 386.400 325.050 387.450 331.950 ;
        RECT 385.950 322.950 388.050 325.050 ;
        RECT 386.400 304.050 387.450 322.950 ;
        RECT 389.400 316.050 390.450 382.950 ;
        RECT 392.400 373.050 393.450 406.950 ;
        RECT 395.400 400.050 396.450 466.950 ;
        RECT 400.950 460.950 403.050 463.050 ;
        RECT 397.950 457.950 400.050 460.050 ;
        RECT 398.400 448.050 399.450 457.950 ;
        RECT 397.950 445.950 400.050 448.050 ;
        RECT 401.400 445.050 402.450 460.950 ;
        RECT 410.400 459.450 411.450 466.950 ;
        RECT 413.400 463.050 414.450 481.950 ;
        RECT 412.950 460.950 415.050 463.050 ;
        RECT 416.400 460.050 417.450 493.950 ;
        RECT 425.400 487.050 426.450 517.950 ;
        RECT 427.950 505.950 430.050 508.050 ;
        RECT 418.950 485.250 420.750 486.150 ;
        RECT 421.950 484.950 424.050 487.050 ;
        RECT 424.950 484.950 427.050 487.050 ;
        RECT 428.400 484.050 429.450 505.950 ;
        RECT 430.950 495.300 433.050 497.400 ;
        RECT 431.550 491.700 432.750 495.300 ;
        RECT 430.950 489.600 433.050 491.700 ;
        RECT 434.400 490.050 435.450 517.950 ;
        RECT 437.400 502.050 438.450 547.950 ;
        RECT 436.950 499.950 439.050 502.050 ;
        RECT 440.400 493.050 441.450 550.950 ;
        RECT 443.400 532.050 444.450 607.950 ;
        RECT 464.400 604.050 465.450 625.950 ;
        RECT 467.400 613.050 468.450 625.950 ;
        RECT 481.950 623.850 484.050 624.750 ;
        RECT 485.550 621.600 486.750 633.600 ;
        RECT 484.950 619.500 487.050 621.600 ;
        RECT 466.950 610.950 469.050 613.050 ;
        RECT 463.950 601.950 466.050 604.050 ;
        RECT 472.950 601.950 475.050 604.050 ;
        RECT 473.400 601.050 474.450 601.950 ;
        RECT 488.400 601.050 489.450 637.950 ;
        RECT 503.400 634.050 504.450 667.950 ;
        RECT 508.950 665.850 511.050 666.750 ;
        RECT 514.950 664.950 517.050 667.050 ;
        RECT 518.250 665.850 519.750 666.750 ;
        RECT 520.950 664.950 523.050 667.050 ;
        RECT 515.400 664.050 516.450 664.950 ;
        RECT 514.950 661.950 517.050 664.050 ;
        RECT 524.400 661.050 525.450 703.950 ;
        RECT 530.400 703.050 531.450 704.400 ;
        RECT 532.950 703.950 535.050 704.400 ;
        RECT 536.250 704.250 537.750 705.150 ;
        RECT 538.950 703.950 541.050 706.050 ;
        RECT 544.950 703.950 547.050 706.050 ;
        RECT 547.950 705.600 550.050 707.700 ;
        RECT 529.950 700.950 532.050 703.050 ;
        RECT 532.950 701.850 534.750 702.750 ;
        RECT 535.950 700.950 538.050 703.050 ;
        RECT 539.250 701.850 541.050 702.750 ;
        RECT 536.400 700.050 537.450 700.950 ;
        RECT 545.400 700.050 546.450 703.950 ;
        RECT 535.950 697.950 538.050 700.050 ;
        RECT 544.950 697.950 547.050 700.050 ;
        RECT 544.950 695.850 547.050 696.750 ;
        RECT 548.550 693.600 549.750 705.600 ;
        RECT 556.950 701.250 559.050 702.150 ;
        RECT 562.950 701.250 565.050 702.150 ;
        RECT 556.950 697.950 559.050 700.050 ;
        RECT 562.950 697.950 565.050 700.050 ;
        RECT 563.400 697.050 564.450 697.950 ;
        RECT 562.950 694.950 565.050 697.050 ;
        RECT 569.400 693.600 570.600 710.400 ;
        RECT 632.550 709.350 633.750 713.100 ;
        RECT 655.950 712.950 658.050 715.050 ;
        RECT 658.950 712.950 661.050 715.050 ;
        RECT 661.950 712.950 664.050 715.050 ;
        RECT 718.950 713.100 721.050 715.200 ;
        RECT 634.950 710.850 637.050 712.950 ;
        RECT 631.950 707.250 634.050 709.350 ;
        RECT 622.950 704.250 625.050 705.150 ;
        RECT 571.950 700.950 574.050 703.050 ;
        RECT 601.950 702.450 604.050 703.050 ;
        RECT 610.950 702.450 613.050 703.050 ;
        RECT 601.950 701.400 606.450 702.450 ;
        RECT 601.950 700.950 604.050 701.400 ;
        RECT 547.950 691.500 550.050 693.600 ;
        RECT 568.950 691.500 571.050 693.600 ;
        RECT 565.950 688.950 568.050 691.050 ;
        RECT 526.950 671.850 529.050 672.750 ;
        RECT 535.950 672.450 538.050 673.050 ;
        RECT 529.950 671.250 532.050 672.150 ;
        RECT 533.400 671.400 538.050 672.450 ;
        RECT 529.950 669.450 532.050 670.050 ;
        RECT 533.400 669.450 534.450 671.400 ;
        RECT 535.950 670.950 538.050 671.400 ;
        RECT 539.250 671.250 540.750 672.150 ;
        RECT 541.950 670.950 544.050 673.050 ;
        RECT 529.950 668.400 534.450 669.450 ;
        RECT 535.950 668.850 537.750 669.750 ;
        RECT 529.950 667.950 532.050 668.400 ;
        RECT 538.950 667.950 541.050 670.050 ;
        RECT 542.250 668.850 543.750 669.750 ;
        RECT 544.950 667.950 547.050 670.050 ;
        RECT 553.950 668.250 555.750 669.150 ;
        RECT 556.950 667.950 559.050 670.050 ;
        RECT 560.250 668.250 562.050 669.150 ;
        RECT 508.950 658.950 511.050 661.050 ;
        RECT 523.950 658.950 526.050 661.050 ;
        RECT 505.950 638.400 508.050 640.500 ;
        RECT 502.950 631.950 505.050 634.050 ;
        RECT 493.950 629.250 496.050 630.150 ;
        RECT 499.950 629.250 502.050 630.150 ;
        RECT 493.950 625.950 496.050 628.050 ;
        RECT 499.950 625.950 502.050 628.050 ;
        RECT 494.400 607.050 495.450 625.950 ;
        RECT 500.400 625.050 501.450 625.950 ;
        RECT 499.950 622.950 502.050 625.050 ;
        RECT 503.400 621.450 504.450 631.950 ;
        RECT 506.400 621.600 507.600 638.400 ;
        RECT 500.400 620.400 504.450 621.450 ;
        RECT 493.950 604.950 496.050 607.050 ;
        RECT 500.400 601.050 501.450 620.400 ;
        RECT 505.950 619.500 508.050 621.600 ;
        RECT 505.950 613.950 508.050 616.050 ;
        RECT 506.400 601.050 507.450 613.950 ;
        RECT 463.950 600.450 466.050 601.050 ;
        RECT 466.950 600.450 469.050 601.050 ;
        RECT 463.950 599.400 469.050 600.450 ;
        RECT 463.950 598.950 466.050 599.400 ;
        RECT 466.950 598.950 469.050 599.400 ;
        RECT 470.250 599.250 471.750 600.150 ;
        RECT 472.950 598.950 475.050 601.050 ;
        RECT 475.950 599.850 478.050 600.750 ;
        RECT 478.950 599.250 481.050 600.150 ;
        RECT 487.950 598.950 490.050 601.050 ;
        RECT 493.950 598.950 496.050 601.050 ;
        RECT 499.950 598.950 502.050 601.050 ;
        RECT 505.950 600.450 508.050 601.050 ;
        RECT 503.400 599.400 508.050 600.450 ;
        RECT 448.950 596.250 450.750 597.150 ;
        RECT 451.950 595.950 454.050 598.050 ;
        RECT 455.250 596.250 457.050 597.150 ;
        RECT 463.950 595.950 466.050 598.050 ;
        RECT 467.250 596.850 468.750 597.750 ;
        RECT 469.950 595.950 472.050 598.050 ;
        RECT 473.250 596.850 475.050 597.750 ;
        RECT 478.950 595.950 481.050 598.050 ;
        RECT 487.950 596.850 490.050 597.750 ;
        RECT 493.950 596.850 496.050 597.750 ;
        RECT 499.950 596.850 502.050 597.750 ;
        RECT 479.400 595.050 480.450 595.950 ;
        RECT 448.950 592.950 451.050 595.050 ;
        RECT 452.250 593.850 453.750 594.750 ;
        RECT 454.950 592.950 457.050 595.050 ;
        RECT 463.950 593.850 466.050 594.750 ;
        RECT 478.950 592.950 481.050 595.050 ;
        RECT 449.400 589.050 450.450 592.950 ;
        RECT 448.950 586.950 451.050 589.050 ;
        RECT 455.400 583.050 456.450 592.950 ;
        RECT 490.950 586.950 493.050 589.050 ;
        RECT 454.950 580.950 457.050 583.050 ;
        RECT 454.950 574.950 457.050 577.050 ;
        RECT 455.400 562.050 456.450 574.950 ;
        RECT 463.950 566.400 466.050 568.500 ;
        RECT 484.950 567.300 487.050 569.400 ;
        RECT 445.950 561.450 448.050 562.050 ;
        RECT 448.950 561.450 451.050 562.050 ;
        RECT 445.950 560.400 451.050 561.450 ;
        RECT 445.950 559.950 448.050 560.400 ;
        RECT 448.950 559.950 451.050 560.400 ;
        RECT 452.250 560.250 453.750 561.150 ;
        RECT 454.950 559.950 457.050 562.050 ;
        RECT 446.400 547.050 447.450 559.950 ;
        RECT 448.950 557.850 450.750 558.750 ;
        RECT 451.950 556.950 454.050 559.050 ;
        RECT 455.250 557.850 457.050 558.750 ;
        RECT 464.400 549.600 465.600 566.400 ;
        RECT 485.250 563.700 486.450 567.300 ;
        RECT 481.950 559.950 484.050 562.050 ;
        RECT 484.950 561.600 487.050 563.700 ;
        RECT 469.950 557.250 472.050 558.150 ;
        RECT 475.950 557.250 478.050 558.150 ;
        RECT 482.400 556.050 483.450 559.950 ;
        RECT 469.950 553.950 472.050 556.050 ;
        RECT 475.950 553.950 478.050 556.050 ;
        RECT 481.950 553.950 484.050 556.050 ;
        RECT 476.400 553.050 477.450 553.950 ;
        RECT 475.950 550.950 478.050 553.050 ;
        RECT 463.950 547.500 466.050 549.600 ;
        RECT 445.950 544.950 448.050 547.050 ;
        RECT 469.950 544.950 472.050 547.050 ;
        RECT 460.950 532.950 463.050 535.050 ;
        RECT 442.950 529.950 445.050 532.050 ;
        RECT 448.950 529.950 451.050 532.050 ;
        RECT 461.400 529.050 462.450 532.950 ;
        RECT 470.400 529.050 471.450 544.950 ;
        RECT 478.950 532.950 481.050 535.050 ;
        RECT 442.950 526.950 445.050 529.050 ;
        RECT 446.250 527.250 448.050 528.150 ;
        RECT 448.950 527.850 451.050 528.750 ;
        RECT 451.950 527.250 454.050 528.150 ;
        RECT 454.950 526.950 457.050 529.050 ;
        RECT 458.250 527.250 459.750 528.150 ;
        RECT 460.950 526.950 463.050 529.050 ;
        RECT 469.950 526.950 472.050 529.050 ;
        RECT 442.950 524.850 444.750 525.750 ;
        RECT 445.950 523.950 448.050 526.050 ;
        RECT 448.950 523.950 451.050 526.050 ;
        RECT 451.950 523.950 454.050 526.050 ;
        RECT 454.950 524.850 456.750 525.750 ;
        RECT 457.950 523.950 460.050 526.050 ;
        RECT 461.250 524.850 462.750 525.750 ;
        RECT 463.950 523.950 466.050 526.050 ;
        RECT 469.950 524.250 471.750 525.150 ;
        RECT 472.950 523.950 475.050 526.050 ;
        RECT 476.250 524.250 478.050 525.150 ;
        RECT 446.400 523.050 447.450 523.950 ;
        RECT 445.950 520.950 448.050 523.050 ;
        RECT 446.400 520.050 447.450 520.950 ;
        RECT 449.400 520.050 450.450 523.950 ;
        RECT 445.950 517.950 448.050 520.050 ;
        RECT 448.950 517.950 451.050 520.050 ;
        RECT 452.400 517.050 453.450 523.950 ;
        RECT 454.950 517.950 457.050 520.050 ;
        RECT 442.950 514.950 445.050 517.050 ;
        RECT 451.950 514.950 454.050 517.050 ;
        RECT 436.950 490.950 439.050 493.050 ;
        RECT 439.950 490.950 442.050 493.050 ;
        RECT 418.950 481.950 421.050 484.050 ;
        RECT 422.250 482.850 424.050 483.750 ;
        RECT 427.950 483.450 430.050 484.050 ;
        RECT 425.400 482.400 430.050 483.450 ;
        RECT 419.400 469.050 420.450 481.950 ;
        RECT 425.400 481.050 426.450 482.400 ;
        RECT 427.950 481.950 430.050 482.400 ;
        RECT 424.950 478.950 427.050 481.050 ;
        RECT 427.950 479.850 430.050 480.750 ;
        RECT 427.950 475.950 430.050 478.050 ;
        RECT 431.550 477.600 432.750 489.600 ;
        RECT 433.950 487.950 436.050 490.050 ;
        RECT 428.400 471.450 429.450 475.950 ;
        RECT 430.950 475.500 433.050 477.600 ;
        RECT 428.400 470.400 432.450 471.450 ;
        RECT 418.950 466.950 421.050 469.050 ;
        RECT 418.950 463.950 421.050 466.050 ;
        RECT 412.950 459.450 415.050 460.050 ;
        RECT 410.400 458.400 415.050 459.450 ;
        RECT 412.950 457.950 415.050 458.400 ;
        RECT 415.950 457.950 418.050 460.050 ;
        RECT 419.400 457.050 420.450 463.950 ;
        RECT 427.950 457.950 430.050 460.050 ;
        RECT 406.950 456.450 409.050 457.050 ;
        RECT 404.400 455.400 409.050 456.450 ;
        RECT 400.950 442.950 403.050 445.050 ;
        RECT 400.950 421.950 403.050 424.050 ;
        RECT 397.950 410.850 400.050 411.750 ;
        RECT 401.400 411.450 402.450 421.950 ;
        RECT 404.400 417.450 405.450 455.400 ;
        RECT 406.950 454.950 409.050 455.400 ;
        RECT 410.250 455.250 412.050 456.150 ;
        RECT 412.950 455.850 415.050 456.750 ;
        RECT 415.950 455.250 418.050 456.150 ;
        RECT 418.950 454.950 421.050 457.050 ;
        RECT 422.250 455.250 423.750 456.150 ;
        RECT 424.950 454.950 427.050 457.050 ;
        RECT 428.400 454.050 429.450 457.950 ;
        RECT 406.950 452.850 408.750 453.750 ;
        RECT 409.950 451.950 412.050 454.050 ;
        RECT 415.950 451.950 418.050 454.050 ;
        RECT 418.950 452.850 420.750 453.750 ;
        RECT 421.950 451.950 424.050 454.050 ;
        RECT 425.250 452.850 426.750 453.750 ;
        RECT 427.950 451.950 430.050 454.050 ;
        RECT 410.400 448.050 411.450 451.950 ;
        RECT 427.950 449.850 430.050 450.750 ;
        RECT 409.950 445.950 412.050 448.050 ;
        RECT 410.400 421.050 411.450 445.950 ;
        RECT 431.400 433.050 432.450 470.400 ;
        RECT 434.400 466.050 435.450 487.950 ;
        RECT 437.400 478.050 438.450 490.950 ;
        RECT 443.400 487.050 444.450 514.950 ;
        RECT 455.400 510.450 456.450 517.950 ;
        RECT 458.400 514.050 459.450 523.950 ;
        RECT 460.950 520.950 463.050 523.050 ;
        RECT 463.950 521.850 466.050 522.750 ;
        RECT 469.950 520.950 472.050 523.050 ;
        RECT 473.250 521.850 474.750 522.750 ;
        RECT 475.950 520.950 478.050 523.050 ;
        RECT 457.950 511.950 460.050 514.050 ;
        RECT 455.400 509.400 459.450 510.450 ;
        RECT 454.950 499.950 457.050 502.050 ;
        RECT 448.950 493.950 451.050 496.050 ;
        RECT 451.950 494.400 454.050 496.500 ;
        RECT 439.950 485.250 442.050 486.150 ;
        RECT 442.950 484.950 445.050 487.050 ;
        RECT 445.950 485.250 448.050 486.150 ;
        RECT 439.950 483.450 442.050 484.050 ;
        RECT 443.400 483.450 444.450 484.950 ;
        RECT 439.950 482.400 444.450 483.450 ;
        RECT 445.950 483.450 448.050 484.050 ;
        RECT 449.400 483.450 450.450 493.950 ;
        RECT 445.950 482.400 450.450 483.450 ;
        RECT 439.950 481.950 442.050 482.400 ;
        RECT 445.950 481.950 448.050 482.400 ;
        RECT 445.950 478.950 448.050 481.050 ;
        RECT 436.950 475.950 439.050 478.050 ;
        RECT 442.950 469.950 445.050 472.050 ;
        RECT 433.950 463.950 436.050 466.050 ;
        RECT 430.950 430.950 433.050 433.050 ;
        RECT 430.950 427.950 433.050 430.050 ;
        RECT 409.950 418.950 412.050 421.050 ;
        RECT 412.950 418.950 415.050 421.050 ;
        RECT 404.400 416.400 408.450 417.450 ;
        RECT 407.400 415.050 408.450 416.400 ;
        RECT 413.400 415.050 414.450 418.950 ;
        RECT 403.950 413.250 405.750 414.150 ;
        RECT 406.950 412.950 409.050 415.050 ;
        RECT 410.250 413.250 411.750 414.150 ;
        RECT 412.950 412.950 415.050 415.050 ;
        RECT 416.250 413.250 418.050 414.150 ;
        RECT 421.950 412.950 424.050 415.050 ;
        RECT 427.950 413.250 430.050 414.150 ;
        RECT 403.950 411.450 406.050 412.050 ;
        RECT 401.400 410.400 406.050 411.450 ;
        RECT 407.250 410.850 408.750 411.750 ;
        RECT 403.950 409.950 406.050 410.400 ;
        RECT 409.950 409.950 412.050 412.050 ;
        RECT 413.250 410.850 414.750 411.750 ;
        RECT 415.950 409.950 418.050 412.050 ;
        RECT 418.950 410.250 421.050 411.150 ;
        RECT 421.950 410.850 424.050 411.750 ;
        RECT 427.950 409.950 430.050 412.050 ;
        RECT 397.950 403.950 400.050 406.050 ;
        RECT 394.950 397.950 397.050 400.050 ;
        RECT 394.950 388.950 397.050 391.050 ;
        RECT 395.400 385.050 396.450 388.950 ;
        RECT 394.950 382.950 397.050 385.050 ;
        RECT 394.950 380.850 397.050 381.750 ;
        RECT 391.950 370.950 394.050 373.050 ;
        RECT 391.950 343.950 394.050 346.050 ;
        RECT 391.950 341.850 394.050 342.750 ;
        RECT 394.950 341.250 397.050 342.150 ;
        RECT 394.950 337.950 397.050 340.050 ;
        RECT 391.950 328.950 394.050 331.050 ;
        RECT 388.950 313.950 391.050 316.050 ;
        RECT 388.950 312.450 391.050 313.050 ;
        RECT 392.400 312.450 393.450 328.950 ;
        RECT 395.400 325.050 396.450 337.950 ;
        RECT 398.400 328.050 399.450 403.950 ;
        RECT 400.950 391.950 403.050 394.050 ;
        RECT 401.400 385.050 402.450 391.950 ;
        RECT 406.950 389.400 409.050 391.500 ;
        RECT 400.950 382.950 403.050 385.050 ;
        RECT 400.950 380.850 403.050 381.750 ;
        RECT 400.950 376.950 403.050 379.050 ;
        RECT 397.950 325.950 400.050 328.050 ;
        RECT 394.950 322.950 397.050 325.050 ;
        RECT 401.400 324.450 402.450 376.950 ;
        RECT 407.400 372.600 408.600 389.400 ;
        RECT 410.400 388.050 411.450 409.950 ;
        RECT 428.400 409.050 429.450 409.950 ;
        RECT 418.950 406.950 421.050 409.050 ;
        RECT 424.950 406.950 427.050 409.050 ;
        RECT 427.950 406.950 430.050 409.050 ;
        RECT 421.950 389.400 424.050 391.500 ;
        RECT 409.950 385.950 412.050 388.050 ;
        RECT 418.950 386.250 421.050 387.150 ;
        RECT 418.950 382.950 421.050 385.050 ;
        RECT 422.550 377.400 423.750 389.400 ;
        RECT 425.400 385.050 426.450 406.950 ;
        RECT 427.950 400.950 430.050 403.050 ;
        RECT 424.950 382.950 427.050 385.050 ;
        RECT 421.950 375.300 424.050 377.400 ;
        RECT 406.950 370.500 409.050 372.600 ;
        RECT 422.550 371.700 423.750 375.300 ;
        RECT 421.950 369.600 424.050 371.700 ;
        RECT 406.950 364.950 409.050 367.050 ;
        RECT 403.950 349.950 406.050 352.050 ;
        RECT 404.400 343.050 405.450 349.950 ;
        RECT 407.400 346.050 408.450 364.950 ;
        RECT 412.950 346.950 415.050 349.050 ;
        RECT 415.950 346.950 418.050 349.050 ;
        RECT 413.400 346.050 414.450 346.950 ;
        RECT 406.950 343.950 409.050 346.050 ;
        RECT 410.250 344.250 411.750 345.150 ;
        RECT 412.950 343.950 415.050 346.050 ;
        RECT 403.950 340.950 406.050 343.050 ;
        RECT 406.950 341.850 408.750 342.750 ;
        RECT 409.950 340.950 412.050 343.050 ;
        RECT 413.250 341.850 415.050 342.750 ;
        RECT 409.950 328.950 412.050 331.050 ;
        RECT 398.400 323.400 402.450 324.450 ;
        RECT 388.950 311.400 393.450 312.450 ;
        RECT 388.950 310.950 391.050 311.400 ;
        RECT 388.950 308.850 391.050 309.750 ;
        RECT 391.950 307.950 394.050 310.050 ;
        RECT 394.950 308.850 397.050 309.750 ;
        RECT 385.950 301.950 388.050 304.050 ;
        RECT 392.400 297.450 393.450 307.950 ;
        RECT 392.400 296.400 396.450 297.450 ;
        RECT 388.950 286.950 391.050 289.050 ;
        RECT 385.950 269.250 388.050 270.150 ;
        RECT 385.950 267.450 388.050 268.050 ;
        RECT 383.400 266.400 388.050 267.450 ;
        RECT 385.950 265.950 388.050 266.400 ;
        RECT 367.950 262.950 370.050 265.050 ;
        RECT 385.950 262.950 388.050 265.050 ;
        RECT 364.950 247.950 367.050 250.050 ;
        RECT 355.950 244.950 358.050 247.050 ;
        RECT 358.950 244.950 361.050 247.050 ;
        RECT 352.950 241.950 355.050 244.050 ;
        RECT 353.400 241.050 354.450 241.950 ;
        RECT 346.950 238.950 349.050 241.050 ;
        RECT 352.950 238.950 355.050 241.050 ;
        RECT 346.950 236.850 349.050 237.750 ;
        RECT 352.950 236.850 355.050 237.750 ;
        RECT 343.950 223.950 346.050 226.050 ;
        RECT 349.950 211.950 352.050 214.050 ;
        RECT 346.950 208.950 349.050 211.050 ;
        RECT 325.950 202.950 328.050 205.050 ;
        RECT 331.950 202.950 334.050 205.050 ;
        RECT 340.950 202.950 343.050 205.050 ;
        RECT 326.400 202.050 327.450 202.950 ;
        RECT 332.400 202.050 333.450 202.950 ;
        RECT 325.950 199.950 328.050 202.050 ;
        RECT 329.250 200.250 330.750 201.150 ;
        RECT 331.950 199.950 334.050 202.050 ;
        RECT 340.950 200.250 343.050 201.150 ;
        RECT 347.400 199.050 348.450 208.950 ;
        RECT 350.400 202.050 351.450 211.950 ;
        RECT 356.400 208.050 357.450 244.950 ;
        RECT 359.400 241.050 360.450 244.950 ;
        RECT 365.400 241.050 366.450 247.950 ;
        RECT 358.950 238.950 361.050 241.050 ;
        RECT 362.250 239.250 364.050 240.150 ;
        RECT 364.950 238.950 367.050 241.050 ;
        RECT 358.950 236.850 360.750 237.750 ;
        RECT 361.950 235.950 364.050 238.050 ;
        RECT 364.950 236.850 367.050 237.750 ;
        RECT 364.950 232.950 367.050 235.050 ;
        RECT 355.950 205.950 358.050 208.050 ;
        RECT 365.400 205.050 366.450 232.950 ;
        RECT 368.400 226.050 369.450 262.950 ;
        RECT 376.950 244.950 379.050 247.050 ;
        RECT 373.950 241.950 376.050 244.050 ;
        RECT 374.400 241.050 375.450 241.950 ;
        RECT 373.950 238.950 376.050 241.050 ;
        RECT 370.950 236.250 373.050 237.150 ;
        RECT 373.950 236.850 376.050 237.750 ;
        RECT 370.950 232.950 373.050 235.050 ;
        RECT 367.950 223.950 370.050 226.050 ;
        RECT 367.950 214.950 370.050 217.050 ;
        RECT 368.400 208.050 369.450 214.950 ;
        RECT 371.400 214.050 372.450 232.950 ;
        RECT 377.400 232.050 378.450 244.950 ;
        RECT 382.950 238.950 385.050 241.050 ;
        RECT 382.950 236.850 385.050 237.750 ;
        RECT 379.950 232.950 382.050 235.050 ;
        RECT 376.950 229.950 379.050 232.050 ;
        RECT 373.950 217.950 376.050 220.050 ;
        RECT 370.950 211.950 373.050 214.050 ;
        RECT 374.400 208.050 375.450 217.950 ;
        RECT 367.950 205.950 370.050 208.050 ;
        RECT 373.950 205.950 376.050 208.050 ;
        RECT 355.950 203.250 358.050 204.150 ;
        RECT 364.950 202.950 367.050 205.050 ;
        RECT 367.950 202.950 370.050 205.050 ;
        RECT 349.950 199.950 352.050 202.050 ;
        RECT 352.950 200.250 354.750 201.150 ;
        RECT 355.950 199.950 358.050 202.050 ;
        RECT 361.950 201.450 364.050 202.050 ;
        RECT 359.250 200.250 360.750 201.150 ;
        RECT 361.950 200.400 366.450 201.450 ;
        RECT 361.950 199.950 364.050 200.400 ;
        RECT 365.400 199.050 366.450 200.400 ;
        RECT 325.950 197.850 327.750 198.750 ;
        RECT 328.950 196.950 331.050 199.050 ;
        RECT 332.250 197.850 334.050 198.750 ;
        RECT 340.950 196.950 343.050 199.050 ;
        RECT 344.250 197.250 345.750 198.150 ;
        RECT 346.950 196.950 349.050 199.050 ;
        RECT 350.250 197.250 352.050 198.150 ;
        RECT 352.950 196.950 355.050 199.050 ;
        RECT 358.950 198.450 361.050 199.050 ;
        RECT 356.400 197.400 361.050 198.450 ;
        RECT 362.250 197.850 364.050 198.750 ;
        RECT 322.950 181.950 325.050 184.050 ;
        RECT 329.400 175.050 330.450 196.950 ;
        RECT 341.400 196.050 342.450 196.950 ;
        RECT 340.950 193.950 343.050 196.050 ;
        RECT 343.950 193.950 346.050 196.050 ;
        RECT 347.250 194.850 348.750 195.750 ;
        RECT 349.950 193.950 352.050 196.050 ;
        RECT 344.400 193.050 345.450 193.950 ;
        RECT 343.950 190.950 346.050 193.050 ;
        RECT 350.400 190.050 351.450 193.950 ;
        RECT 334.950 187.950 337.050 190.050 ;
        RECT 349.950 187.950 352.050 190.050 ;
        RECT 328.950 172.950 331.050 175.050 ;
        RECT 313.950 167.250 316.050 168.150 ;
        RECT 316.950 167.850 319.050 168.750 ;
        RECT 319.950 166.950 322.050 169.050 ;
        RECT 329.400 168.450 330.450 172.950 ;
        RECT 335.400 169.050 336.450 187.950 ;
        RECT 340.950 184.950 343.050 187.050 ;
        RECT 353.400 186.450 354.450 196.950 ;
        RECT 356.400 193.050 357.450 197.400 ;
        RECT 358.950 196.950 361.050 197.400 ;
        RECT 364.950 196.950 367.050 199.050 ;
        RECT 368.400 198.450 369.450 202.950 ;
        RECT 374.400 202.050 375.450 205.950 ;
        RECT 377.400 202.050 378.450 229.950 ;
        RECT 380.400 223.050 381.450 232.950 ;
        RECT 386.400 223.050 387.450 262.950 ;
        RECT 389.400 262.050 390.450 286.950 ;
        RECT 391.950 269.250 394.050 270.150 ;
        RECT 391.950 262.950 394.050 265.050 ;
        RECT 388.950 259.950 391.050 262.050 ;
        RECT 392.400 249.450 393.450 262.950 ;
        RECT 395.400 253.050 396.450 296.400 ;
        RECT 398.400 295.050 399.450 323.400 ;
        RECT 410.400 322.050 411.450 328.950 ;
        RECT 416.400 325.050 417.450 346.950 ;
        RECT 428.400 346.050 429.450 400.950 ;
        RECT 431.400 400.050 432.450 427.950 ;
        RECT 434.400 418.050 435.450 463.950 ;
        RECT 436.950 455.250 439.050 456.150 ;
        RECT 436.950 451.950 439.050 454.050 ;
        RECT 437.400 451.050 438.450 451.950 ;
        RECT 436.950 448.950 439.050 451.050 ;
        RECT 433.950 415.950 436.050 418.050 ;
        RECT 433.950 413.250 436.050 414.150 ;
        RECT 433.950 406.950 436.050 409.050 ;
        RECT 430.950 397.950 433.050 400.050 ;
        RECT 430.950 388.950 433.050 391.050 ;
        RECT 431.400 385.050 432.450 388.950 ;
        RECT 430.950 382.950 433.050 385.050 ;
        RECT 430.950 380.850 433.050 381.750 ;
        RECT 434.400 373.050 435.450 406.950 ;
        RECT 437.400 391.050 438.450 448.950 ;
        RECT 439.950 433.950 442.050 436.050 ;
        RECT 440.400 403.050 441.450 433.950 ;
        RECT 443.400 418.050 444.450 469.950 ;
        RECT 446.400 439.050 447.450 478.950 ;
        RECT 452.400 477.600 453.600 494.400 ;
        RECT 451.950 475.500 454.050 477.600 ;
        RECT 455.400 448.050 456.450 499.950 ;
        RECT 458.400 472.050 459.450 509.400 ;
        RECT 461.400 496.050 462.450 520.950 ;
        RECT 470.400 508.050 471.450 520.950 ;
        RECT 472.950 517.950 475.050 520.050 ;
        RECT 473.400 511.050 474.450 517.950 ;
        RECT 476.400 514.050 477.450 520.950 ;
        RECT 479.400 517.050 480.450 532.950 ;
        RECT 482.400 517.050 483.450 553.950 ;
        RECT 485.250 549.600 486.450 561.600 ;
        RECT 487.950 553.950 490.050 556.050 ;
        RECT 487.950 551.850 490.050 552.750 ;
        RECT 484.950 547.500 487.050 549.600 ;
        RECT 487.950 533.400 490.050 535.500 ;
        RECT 484.950 530.250 487.050 531.150 ;
        RECT 484.950 526.950 487.050 529.050 ;
        RECT 485.400 523.050 486.450 526.950 ;
        RECT 484.950 520.950 487.050 523.050 ;
        RECT 488.550 521.400 489.750 533.400 ;
        RECT 487.950 519.300 490.050 521.400 ;
        RECT 491.400 520.050 492.450 586.950 ;
        RECT 503.400 577.050 504.450 599.400 ;
        RECT 505.950 598.950 508.050 599.400 ;
        RECT 505.950 596.850 508.050 597.750 ;
        RECT 505.950 592.950 508.050 595.050 ;
        RECT 493.950 574.950 496.050 577.050 ;
        RECT 502.950 574.950 505.050 577.050 ;
        RECT 494.400 555.450 495.450 574.950 ;
        RECT 496.950 557.250 499.050 558.150 ;
        RECT 502.950 557.250 505.050 558.150 ;
        RECT 496.950 555.450 499.050 556.050 ;
        RECT 494.400 554.400 499.050 555.450 ;
        RECT 496.950 553.950 499.050 554.400 ;
        RECT 502.950 553.950 505.050 556.050 ;
        RECT 493.950 550.950 496.050 553.050 ;
        RECT 494.400 528.450 495.450 550.950 ;
        RECT 503.400 547.050 504.450 553.950 ;
        RECT 502.950 544.950 505.050 547.050 ;
        RECT 502.950 529.950 505.050 532.050 ;
        RECT 503.400 529.050 504.450 529.950 ;
        RECT 496.950 528.450 499.050 529.050 ;
        RECT 494.400 527.400 499.050 528.450 ;
        RECT 478.950 514.950 481.050 517.050 ;
        RECT 481.950 514.950 484.050 517.050 ;
        RECT 488.550 515.700 489.750 519.300 ;
        RECT 490.950 517.950 493.050 520.050 ;
        RECT 475.950 511.950 478.050 514.050 ;
        RECT 487.950 513.600 490.050 515.700 ;
        RECT 490.950 514.950 493.050 517.050 ;
        RECT 472.950 508.950 475.050 511.050 ;
        RECT 478.950 508.950 481.050 511.050 ;
        RECT 469.950 505.950 472.050 508.050 ;
        RECT 460.950 493.950 463.050 496.050 ;
        RECT 472.950 493.950 475.050 496.050 ;
        RECT 460.950 490.950 463.050 493.050 ;
        RECT 457.950 469.950 460.050 472.050 ;
        RECT 457.950 455.250 460.050 456.150 ;
        RECT 454.950 445.950 457.050 448.050 ;
        RECT 461.400 442.050 462.450 490.950 ;
        RECT 466.950 487.950 469.050 490.050 ;
        RECT 463.950 484.950 466.050 487.050 ;
        RECT 463.950 482.850 466.050 483.750 ;
        RECT 463.950 469.950 466.050 472.050 ;
        RECT 464.400 463.050 465.450 469.950 ;
        RECT 463.950 460.950 466.050 463.050 ;
        RECT 463.950 454.950 466.050 457.050 ;
        RECT 464.400 445.050 465.450 454.950 ;
        RECT 463.950 442.950 466.050 445.050 ;
        RECT 451.950 439.950 454.050 442.050 ;
        RECT 460.950 439.950 463.050 442.050 ;
        RECT 445.950 436.950 448.050 439.050 ;
        RECT 445.950 427.950 448.050 430.050 ;
        RECT 442.950 415.950 445.050 418.050 ;
        RECT 442.950 413.250 445.050 414.150 ;
        RECT 442.950 409.950 445.050 412.050 ;
        RECT 439.950 400.950 442.050 403.050 ;
        RECT 443.400 397.050 444.450 409.950 ;
        RECT 439.950 394.950 442.050 397.050 ;
        RECT 442.950 394.950 445.050 397.050 ;
        RECT 436.950 388.950 439.050 391.050 ;
        RECT 436.950 385.950 439.050 388.050 ;
        RECT 437.400 385.050 438.450 385.950 ;
        RECT 436.950 382.950 439.050 385.050 ;
        RECT 436.950 380.850 439.050 381.750 ;
        RECT 433.950 370.950 436.050 373.050 ;
        RECT 440.400 366.450 441.450 394.950 ;
        RECT 442.950 389.400 445.050 391.500 ;
        RECT 443.400 372.600 444.600 389.400 ;
        RECT 442.950 370.500 445.050 372.600 ;
        RECT 440.400 365.400 444.450 366.450 ;
        RECT 439.950 361.950 442.050 364.050 ;
        RECT 440.400 352.050 441.450 361.950 ;
        RECT 439.950 349.950 442.050 352.050 ;
        RECT 418.950 343.950 421.050 346.050 ;
        RECT 427.950 343.950 430.050 346.050 ;
        RECT 436.950 344.250 439.050 345.150 ;
        RECT 415.950 322.950 418.050 325.050 ;
        RECT 409.950 319.950 412.050 322.050 ;
        RECT 412.950 319.950 415.050 322.050 ;
        RECT 400.950 313.950 403.050 316.050 ;
        RECT 401.400 313.050 402.450 313.950 ;
        RECT 400.950 310.950 403.050 313.050 ;
        RECT 400.950 308.850 403.050 309.750 ;
        RECT 406.950 308.850 409.050 309.750 ;
        RECT 410.400 307.050 411.450 319.950 ;
        RECT 413.400 313.050 414.450 319.950 ;
        RECT 412.950 310.950 415.050 313.050 ;
        RECT 416.400 310.050 417.450 322.950 ;
        RECT 419.400 316.050 420.450 343.950 ;
        RECT 421.950 340.950 424.050 343.050 ;
        RECT 427.950 341.250 429.750 342.150 ;
        RECT 430.950 340.950 433.050 343.050 ;
        RECT 436.950 342.450 439.050 343.050 ;
        RECT 440.400 342.450 441.450 349.950 ;
        RECT 443.400 343.050 444.450 365.400 ;
        RECT 446.400 352.050 447.450 427.950 ;
        RECT 448.950 413.250 451.050 414.150 ;
        RECT 448.950 409.950 451.050 412.050 ;
        RECT 449.400 409.050 450.450 409.950 ;
        RECT 448.950 406.950 451.050 409.050 ;
        RECT 448.950 400.950 451.050 403.050 ;
        RECT 449.400 367.050 450.450 400.950 ;
        RECT 452.400 379.050 453.450 439.950 ;
        RECT 457.950 421.950 460.050 424.050 ;
        RECT 458.400 418.050 459.450 421.950 ;
        RECT 464.400 421.050 465.450 442.950 ;
        RECT 463.950 418.950 466.050 421.050 ;
        RECT 457.950 415.950 460.050 418.050 ;
        RECT 461.250 416.250 462.750 417.150 ;
        RECT 463.950 415.950 466.050 418.050 ;
        RECT 457.950 413.850 459.750 414.750 ;
        RECT 460.950 412.950 463.050 415.050 ;
        RECT 464.250 413.850 466.050 414.750 ;
        RECT 461.400 400.050 462.450 412.950 ;
        RECT 467.400 403.050 468.450 487.950 ;
        RECT 473.400 457.050 474.450 493.950 ;
        RECT 479.400 487.050 480.450 508.950 ;
        RECT 487.950 493.950 490.050 496.050 ;
        RECT 478.950 484.950 481.050 487.050 ;
        RECT 484.950 482.850 487.050 483.750 ;
        RECT 488.400 481.050 489.450 493.950 ;
        RECT 487.950 478.950 490.050 481.050 ;
        RECT 478.950 463.950 481.050 466.050 ;
        RECT 472.950 454.950 475.050 457.050 ;
        RECT 469.950 452.250 471.750 453.150 ;
        RECT 472.950 451.950 475.050 454.050 ;
        RECT 476.250 452.250 478.050 453.150 ;
        RECT 469.950 448.950 472.050 451.050 ;
        RECT 473.250 449.850 474.750 450.750 ;
        RECT 475.950 448.950 478.050 451.050 ;
        RECT 476.400 445.050 477.450 448.950 ;
        RECT 475.950 442.950 478.050 445.050 ;
        RECT 479.400 427.050 480.450 463.950 ;
        RECT 481.950 452.250 483.750 453.150 ;
        RECT 484.950 451.950 487.050 454.050 ;
        RECT 488.250 452.250 490.050 453.150 ;
        RECT 481.950 448.950 484.050 451.050 ;
        RECT 485.250 449.850 486.750 450.750 ;
        RECT 487.950 448.950 490.050 451.050 ;
        RECT 482.400 448.050 483.450 448.950 ;
        RECT 481.950 445.950 484.050 448.050 ;
        RECT 491.400 433.050 492.450 514.950 ;
        RECT 494.400 511.050 495.450 527.400 ;
        RECT 496.950 526.950 499.050 527.400 ;
        RECT 502.950 526.950 505.050 529.050 ;
        RECT 496.950 524.850 499.050 525.750 ;
        RECT 502.950 524.850 505.050 525.750 ;
        RECT 506.400 523.050 507.450 592.950 ;
        RECT 509.400 565.050 510.450 658.950 ;
        RECT 517.950 640.950 520.050 643.050 ;
        RECT 511.950 634.950 514.050 637.050 ;
        RECT 512.400 628.050 513.450 634.950 ;
        RECT 514.950 629.250 517.050 630.150 ;
        RECT 511.950 625.950 514.050 628.050 ;
        RECT 514.950 625.950 517.050 628.050 ;
        RECT 512.400 595.050 513.450 625.950 ;
        RECT 515.400 616.050 516.450 625.950 ;
        RECT 518.400 616.050 519.450 640.950 ;
        RECT 530.400 639.450 531.450 667.950 ;
        RECT 539.400 667.050 540.450 667.950 ;
        RECT 538.950 664.950 541.050 667.050 ;
        RECT 544.950 665.850 547.050 666.750 ;
        RECT 553.950 664.950 556.050 667.050 ;
        RECT 557.250 665.850 558.750 666.750 ;
        RECT 559.950 664.950 562.050 667.050 ;
        RECT 527.400 638.400 531.450 639.450 ;
        RECT 520.950 629.250 523.050 630.150 ;
        RECT 520.950 625.950 523.050 628.050 ;
        RECT 514.950 613.950 517.050 616.050 ;
        RECT 517.950 613.950 520.050 616.050 ;
        RECT 515.400 613.050 516.450 613.950 ;
        RECT 514.950 610.950 517.050 613.050 ;
        RECT 527.400 604.050 528.450 638.400 ;
        RECT 538.950 634.950 541.050 637.050 ;
        RECT 539.400 634.050 540.450 634.950 ;
        RECT 554.400 634.050 555.450 664.950 ;
        RECT 560.400 649.050 561.450 664.950 ;
        RECT 559.950 646.950 562.050 649.050 ;
        RECT 556.950 640.950 559.050 643.050 ;
        RECT 532.950 633.450 535.050 634.050 ;
        RECT 530.400 632.400 535.050 633.450 ;
        RECT 530.400 628.050 531.450 632.400 ;
        RECT 532.950 631.950 535.050 632.400 ;
        RECT 536.250 632.250 537.750 633.150 ;
        RECT 538.950 631.950 541.050 634.050 ;
        RECT 544.950 632.250 547.050 633.150 ;
        RECT 550.950 631.950 553.050 634.050 ;
        RECT 553.950 631.950 556.050 634.050 ;
        RECT 551.400 631.050 552.450 631.950 ;
        RECT 532.950 629.850 534.750 630.750 ;
        RECT 535.950 628.950 538.050 631.050 ;
        RECT 539.250 629.850 541.050 630.750 ;
        RECT 544.950 628.950 547.050 631.050 ;
        RECT 548.250 629.250 549.750 630.150 ;
        RECT 550.950 628.950 553.050 631.050 ;
        RECT 554.250 629.250 556.050 630.150 ;
        RECT 529.950 625.950 532.050 628.050 ;
        RECT 547.950 625.950 550.050 628.050 ;
        RECT 551.250 626.850 552.750 627.750 ;
        RECT 553.950 625.950 556.050 628.050 ;
        RECT 548.400 625.050 549.450 625.950 ;
        RECT 547.950 622.950 550.050 625.050 ;
        RECT 538.950 616.950 541.050 619.050 ;
        RECT 526.950 601.950 529.050 604.050 ;
        RECT 535.950 601.950 538.050 604.050 ;
        RECT 536.400 601.050 537.450 601.950 ;
        RECT 523.950 598.950 526.050 601.050 ;
        RECT 529.950 598.950 532.050 601.050 ;
        RECT 533.250 599.250 534.750 600.150 ;
        RECT 535.950 598.950 538.050 601.050 ;
        RECT 539.400 600.450 540.450 616.950 ;
        RECT 544.950 605.400 547.050 607.500 ;
        RECT 554.400 607.050 555.450 625.950 ;
        RECT 541.950 602.250 544.050 603.150 ;
        RECT 541.950 600.450 544.050 601.050 ;
        RECT 539.400 599.400 544.050 600.450 ;
        RECT 541.950 598.950 544.050 599.400 ;
        RECT 514.950 596.250 516.750 597.150 ;
        RECT 517.950 595.950 520.050 598.050 ;
        RECT 521.250 596.250 523.050 597.150 ;
        RECT 511.950 592.950 514.050 595.050 ;
        RECT 514.950 592.950 517.050 595.050 ;
        RECT 518.250 593.850 519.750 594.750 ;
        RECT 520.950 592.950 523.050 595.050 ;
        RECT 515.400 583.050 516.450 592.950 ;
        RECT 514.950 580.950 517.050 583.050 ;
        RECT 508.950 562.950 511.050 565.050 ;
        RECT 509.400 547.050 510.450 562.950 ;
        RECT 511.950 557.250 514.050 558.150 ;
        RECT 511.950 555.450 514.050 556.050 ;
        RECT 515.400 555.450 516.450 580.950 ;
        RECT 521.400 580.050 522.450 592.950 ;
        RECT 524.400 589.050 525.450 598.950 ;
        RECT 526.950 595.950 529.050 598.050 ;
        RECT 530.250 596.850 531.750 597.750 ;
        RECT 532.950 595.950 535.050 598.050 ;
        RECT 536.250 596.850 538.050 597.750 ;
        RECT 533.400 595.050 534.450 595.950 ;
        RECT 526.950 593.850 529.050 594.750 ;
        RECT 532.950 592.950 535.050 595.050 ;
        RECT 532.950 589.950 535.050 592.050 ;
        RECT 523.950 586.950 526.050 589.050 ;
        RECT 520.950 577.950 523.050 580.050 ;
        RECT 517.950 557.250 520.050 558.150 ;
        RECT 511.950 554.400 516.450 555.450 ;
        RECT 511.950 553.950 514.050 554.400 ;
        RECT 517.950 553.950 520.050 556.050 ;
        RECT 518.400 553.050 519.450 553.950 ;
        RECT 517.950 550.950 520.050 553.050 ;
        RECT 508.950 544.950 511.050 547.050 ;
        RECT 508.950 533.400 511.050 535.500 ;
        RECT 521.400 535.050 522.450 577.950 ;
        RECT 523.950 557.250 526.050 558.150 ;
        RECT 529.950 557.250 532.050 558.150 ;
        RECT 529.950 553.950 532.050 556.050 ;
        RECT 529.950 544.950 532.050 547.050 ;
        RECT 526.950 541.950 529.050 544.050 ;
        RECT 527.400 538.050 528.450 541.950 ;
        RECT 526.950 535.950 529.050 538.050 ;
        RECT 502.950 520.950 505.050 523.050 ;
        RECT 505.950 520.950 508.050 523.050 ;
        RECT 503.400 514.050 504.450 520.950 ;
        RECT 505.950 514.950 508.050 517.050 ;
        RECT 509.400 516.600 510.600 533.400 ;
        RECT 514.950 532.950 517.050 535.050 ;
        RECT 520.950 532.950 523.050 535.050 ;
        RECT 511.950 526.950 514.050 529.050 ;
        RECT 502.950 511.950 505.050 514.050 ;
        RECT 493.950 508.950 496.050 511.050 ;
        RECT 493.950 488.250 496.050 489.150 ;
        RECT 497.250 485.250 498.750 486.150 ;
        RECT 499.950 484.950 502.050 487.050 ;
        RECT 503.250 485.250 505.050 486.150 ;
        RECT 496.950 481.950 499.050 484.050 ;
        RECT 500.250 482.850 501.750 483.750 ;
        RECT 502.950 481.950 505.050 484.050 ;
        RECT 497.400 475.050 498.450 481.950 ;
        RECT 502.950 478.950 505.050 481.050 ;
        RECT 496.950 472.950 499.050 475.050 ;
        RECT 503.400 454.050 504.450 478.950 ;
        RECT 506.400 460.050 507.450 514.950 ;
        RECT 508.950 514.500 511.050 516.600 ;
        RECT 512.400 493.050 513.450 526.950 ;
        RECT 511.950 490.950 514.050 493.050 ;
        RECT 515.400 490.050 516.450 532.950 ;
        RECT 523.950 529.950 526.050 532.050 ;
        RECT 524.400 529.050 525.450 529.950 ;
        RECT 517.950 526.950 520.050 529.050 ;
        RECT 521.250 527.250 522.750 528.150 ;
        RECT 523.950 526.950 526.050 529.050 ;
        RECT 517.950 524.850 519.750 525.750 ;
        RECT 520.950 523.950 523.050 526.050 ;
        RECT 524.250 524.850 525.750 525.750 ;
        RECT 526.950 523.950 529.050 526.050 ;
        RECT 530.400 523.050 531.450 544.950 ;
        RECT 533.400 532.050 534.450 589.950 ;
        RECT 538.950 567.300 541.050 569.400 ;
        RECT 539.550 563.700 540.750 567.300 ;
        RECT 538.950 561.600 541.050 563.700 ;
        RECT 535.950 556.950 538.050 559.050 ;
        RECT 536.400 556.050 537.450 556.950 ;
        RECT 535.950 553.950 538.050 556.050 ;
        RECT 535.950 551.850 538.050 552.750 ;
        RECT 539.550 549.600 540.750 561.600 ;
        RECT 538.950 547.500 541.050 549.600 ;
        RECT 532.950 529.950 535.050 532.050 ;
        RECT 542.400 531.450 543.450 598.950 ;
        RECT 545.550 593.400 546.750 605.400 ;
        RECT 550.950 604.950 553.050 607.050 ;
        RECT 553.950 604.950 556.050 607.050 ;
        RECT 551.400 604.050 552.450 604.950 ;
        RECT 550.950 601.950 553.050 604.050 ;
        RECT 553.950 601.950 556.050 604.050 ;
        RECT 544.950 591.300 547.050 593.400 ;
        RECT 545.550 587.700 546.750 591.300 ;
        RECT 544.950 585.600 547.050 587.700 ;
        RECT 547.950 577.950 550.050 580.050 ;
        RECT 548.400 574.050 549.450 577.950 ;
        RECT 547.950 571.950 550.050 574.050 ;
        RECT 547.950 557.250 550.050 558.150 ;
        RECT 547.950 555.450 550.050 556.050 ;
        RECT 551.400 555.450 552.450 601.950 ;
        RECT 554.400 601.050 555.450 601.950 ;
        RECT 553.950 598.950 556.050 601.050 ;
        RECT 553.950 596.850 556.050 597.750 ;
        RECT 557.400 592.050 558.450 640.950 ;
        RECT 566.400 634.050 567.450 688.950 ;
        RECT 568.950 677.400 571.050 679.500 ;
        RECT 569.400 660.600 570.600 677.400 ;
        RECT 568.950 658.500 571.050 660.600 ;
        RECT 572.400 651.450 573.450 700.950 ;
        RECT 605.400 700.050 606.450 701.400 ;
        RECT 608.400 701.400 613.050 702.450 ;
        RECT 580.950 698.850 583.050 699.750 ;
        RECT 601.950 698.850 604.050 699.750 ;
        RECT 604.950 697.950 607.050 700.050 ;
        RECT 580.950 694.950 583.050 697.050 ;
        RECT 586.950 694.950 589.050 697.050 ;
        RECT 608.400 696.450 609.450 701.400 ;
        RECT 610.950 700.950 613.050 701.400 ;
        RECT 622.950 700.950 625.050 703.050 ;
        RECT 623.400 700.050 624.450 700.950 ;
        RECT 610.950 698.850 613.050 699.750 ;
        RECT 622.950 697.950 625.050 700.050 ;
        RECT 625.950 697.950 628.050 700.050 ;
        RECT 608.400 695.400 612.450 696.450 ;
        RECT 581.400 673.050 582.450 694.950 ;
        RECT 574.950 670.950 577.050 673.050 ;
        RECT 580.950 670.950 583.050 673.050 ;
        RECT 574.950 668.850 577.050 669.750 ;
        RECT 580.950 668.850 583.050 669.750 ;
        RECT 569.400 650.400 573.450 651.450 ;
        RECT 559.950 631.950 562.050 634.050 ;
        RECT 563.250 632.250 564.750 633.150 ;
        RECT 565.950 631.950 568.050 634.050 ;
        RECT 559.950 629.850 561.750 630.750 ;
        RECT 562.950 628.950 565.050 631.050 ;
        RECT 566.250 629.850 568.050 630.750 ;
        RECT 562.950 613.950 565.050 616.050 ;
        RECT 559.950 598.950 562.050 601.050 ;
        RECT 559.950 596.850 562.050 597.750 ;
        RECT 556.950 589.950 559.050 592.050 ;
        RECT 556.950 586.950 559.050 589.050 ;
        RECT 557.400 574.050 558.450 586.950 ;
        RECT 563.400 582.450 564.450 613.950 ;
        RECT 565.950 605.400 568.050 607.500 ;
        RECT 566.400 588.600 567.600 605.400 ;
        RECT 565.950 586.500 568.050 588.600 ;
        RECT 569.400 583.050 570.450 650.400 ;
        RECT 571.950 632.250 574.050 633.150 ;
        RECT 571.950 628.950 574.050 631.050 ;
        RECT 575.250 629.250 576.750 630.150 ;
        RECT 577.950 628.950 580.050 631.050 ;
        RECT 581.250 629.250 583.050 630.150 ;
        RECT 583.950 629.250 586.050 630.150 ;
        RECT 574.950 625.950 577.050 628.050 ;
        RECT 578.250 626.850 579.750 627.750 ;
        RECT 580.950 625.950 583.050 628.050 ;
        RECT 583.950 625.950 586.050 628.050 ;
        RECT 575.400 610.050 576.450 625.950 ;
        RECT 577.950 616.950 580.050 619.050 ;
        RECT 574.950 607.950 577.050 610.050 ;
        RECT 563.400 581.400 567.450 582.450 ;
        RECT 556.950 571.950 559.050 574.050 ;
        RECT 553.950 557.250 556.050 558.150 ;
        RECT 547.950 554.400 552.450 555.450 ;
        RECT 547.950 553.950 550.050 554.400 ;
        RECT 553.950 553.950 556.050 556.050 ;
        RECT 550.950 532.950 553.050 535.050 ;
        RECT 542.400 530.400 546.450 531.450 ;
        RECT 545.400 529.050 546.450 530.400 ;
        RECT 551.400 529.050 552.450 532.950 ;
        RECT 554.400 532.050 555.450 553.950 ;
        RECT 557.400 553.050 558.450 571.950 ;
        RECT 559.950 566.400 562.050 568.500 ;
        RECT 556.950 550.950 559.050 553.050 ;
        RECT 560.400 549.600 561.600 566.400 ;
        RECT 562.950 553.950 565.050 556.050 ;
        RECT 559.950 547.500 562.050 549.600 ;
        RECT 563.400 544.050 564.450 553.950 ;
        RECT 566.400 553.050 567.450 581.400 ;
        RECT 568.950 580.950 571.050 583.050 ;
        RECT 571.950 562.950 574.050 565.050 ;
        RECT 568.950 557.250 571.050 558.150 ;
        RECT 568.950 553.950 571.050 556.050 ;
        RECT 572.400 555.450 573.450 562.950 ;
        RECT 574.950 557.250 577.050 558.150 ;
        RECT 574.950 555.450 577.050 556.050 ;
        RECT 572.400 554.400 577.050 555.450 ;
        RECT 574.950 553.950 577.050 554.400 ;
        RECT 565.950 550.950 568.050 553.050 ;
        RECT 574.950 550.950 577.050 553.050 ;
        RECT 565.950 544.950 568.050 547.050 ;
        RECT 562.950 541.950 565.050 544.050 ;
        RECT 563.400 532.050 564.450 541.950 ;
        RECT 553.950 529.950 556.050 532.050 ;
        RECT 562.950 529.950 565.050 532.050 ;
        RECT 541.950 526.950 544.050 529.050 ;
        RECT 544.950 528.450 547.050 529.050 ;
        RECT 544.950 527.400 549.450 528.450 ;
        RECT 544.950 526.950 547.050 527.400 ;
        RECT 542.400 526.050 543.450 526.950 ;
        RECT 532.950 524.250 534.750 525.150 ;
        RECT 535.950 523.950 538.050 526.050 ;
        RECT 539.250 524.250 541.050 525.150 ;
        RECT 541.950 523.950 544.050 526.050 ;
        RECT 544.950 524.850 547.050 525.750 ;
        RECT 520.950 520.950 523.050 523.050 ;
        RECT 523.950 520.950 526.050 523.050 ;
        RECT 526.950 521.850 529.050 522.750 ;
        RECT 529.950 520.950 532.050 523.050 ;
        RECT 532.950 520.950 535.050 523.050 ;
        RECT 536.250 521.850 537.750 522.750 ;
        RECT 538.950 522.450 541.050 523.050 ;
        RECT 542.400 522.450 543.450 523.950 ;
        RECT 538.950 521.400 543.450 522.450 ;
        RECT 538.950 520.950 541.050 521.400 ;
        RECT 521.400 508.050 522.450 520.950 ;
        RECT 520.950 505.950 523.050 508.050 ;
        RECT 521.400 490.050 522.450 505.950 ;
        RECT 514.950 487.950 517.050 490.050 ;
        RECT 518.250 488.250 519.750 489.150 ;
        RECT 520.950 487.950 523.050 490.050 ;
        RECT 508.950 484.950 511.050 487.050 ;
        RECT 514.950 485.850 516.750 486.750 ;
        RECT 517.950 484.950 520.050 487.050 ;
        RECT 521.250 485.850 523.050 486.750 ;
        RECT 508.950 482.850 511.050 483.750 ;
        RECT 511.950 482.250 514.050 483.150 ;
        RECT 514.950 481.950 517.050 484.050 ;
        RECT 511.950 480.450 514.050 481.050 ;
        RECT 515.400 480.450 516.450 481.950 ;
        RECT 511.950 479.400 516.450 480.450 ;
        RECT 511.950 478.950 514.050 479.400 ;
        RECT 508.950 460.950 511.050 463.050 ;
        RECT 505.950 457.950 508.050 460.050 ;
        RECT 509.400 456.450 510.450 460.950 ;
        RECT 512.400 457.050 513.450 478.950 ;
        RECT 518.400 472.050 519.450 484.950 ;
        RECT 517.950 469.950 520.050 472.050 ;
        RECT 524.400 466.050 525.450 520.950 ;
        RECT 526.950 514.950 529.050 517.050 ;
        RECT 527.400 490.050 528.450 514.950 ;
        RECT 533.400 514.050 534.450 520.950 ;
        RECT 548.400 517.050 549.450 527.400 ;
        RECT 550.950 526.950 553.050 529.050 ;
        RECT 556.950 528.450 559.050 529.050 ;
        RECT 554.400 527.400 559.050 528.450 ;
        RECT 550.950 524.850 553.050 525.750 ;
        RECT 547.950 514.950 550.050 517.050 ;
        RECT 532.950 511.950 535.050 514.050 ;
        RECT 535.950 511.950 538.050 514.050 ;
        RECT 529.950 508.950 532.050 511.050 ;
        RECT 530.400 499.050 531.450 508.950 ;
        RECT 536.400 505.050 537.450 511.950 ;
        RECT 535.950 502.950 538.050 505.050 ;
        RECT 538.950 502.950 541.050 505.050 ;
        RECT 529.950 496.950 532.050 499.050 ;
        RECT 532.950 496.950 535.050 499.050 ;
        RECT 526.950 487.950 529.050 490.050 ;
        RECT 533.400 487.050 534.450 496.950 ;
        RECT 539.400 487.050 540.450 502.950 ;
        RECT 554.400 502.050 555.450 527.400 ;
        RECT 556.950 526.950 559.050 527.400 ;
        RECT 560.250 527.250 561.750 528.150 ;
        RECT 562.950 526.950 565.050 529.050 ;
        RECT 566.400 526.050 567.450 544.950 ;
        RECT 568.950 541.950 571.050 544.050 ;
        RECT 556.950 524.850 558.750 525.750 ;
        RECT 559.950 523.950 562.050 526.050 ;
        RECT 563.250 524.850 564.750 525.750 ;
        RECT 565.950 523.950 568.050 526.050 ;
        RECT 560.400 514.050 561.450 523.950 ;
        RECT 562.950 520.950 565.050 523.050 ;
        RECT 565.950 521.850 568.050 522.750 ;
        RECT 559.950 511.950 562.050 514.050 ;
        RECT 563.400 504.450 564.450 520.950 ;
        RECT 569.400 519.450 570.450 541.950 ;
        RECT 575.400 538.050 576.450 550.950 ;
        RECT 578.400 544.050 579.450 616.950 ;
        RECT 584.400 613.050 585.450 625.950 ;
        RECT 587.400 619.050 588.450 694.950 ;
        RECT 589.950 677.400 592.050 679.500 ;
        RECT 590.250 665.400 591.450 677.400 ;
        RECT 592.950 674.250 595.050 675.150 ;
        RECT 592.950 670.950 595.050 673.050 ;
        RECT 593.400 667.050 594.450 670.950 ;
        RECT 601.950 668.250 603.750 669.150 ;
        RECT 604.950 667.950 607.050 670.050 ;
        RECT 608.250 668.250 610.050 669.150 ;
        RECT 589.950 663.300 592.050 665.400 ;
        RECT 592.950 664.950 595.050 667.050 ;
        RECT 601.950 666.450 604.050 667.050 ;
        RECT 599.400 665.400 604.050 666.450 ;
        RECT 605.250 665.850 606.750 666.750 ;
        RECT 590.250 659.700 591.450 663.300 ;
        RECT 589.950 657.600 592.050 659.700 ;
        RECT 592.950 655.950 595.050 658.050 ;
        RECT 593.400 631.050 594.450 655.950 ;
        RECT 599.400 637.050 600.450 665.400 ;
        RECT 601.950 664.950 604.050 665.400 ;
        RECT 607.950 664.950 610.050 667.050 ;
        RECT 604.950 661.950 607.050 664.050 ;
        RECT 598.950 634.950 601.050 637.050 ;
        RECT 605.400 636.450 606.450 661.950 ;
        RECT 608.400 658.050 609.450 664.950 ;
        RECT 607.950 655.950 610.050 658.050 ;
        RECT 605.400 635.400 609.450 636.450 ;
        RECT 599.400 631.050 600.450 634.950 ;
        RECT 604.950 632.250 607.050 633.150 ;
        RECT 589.950 629.250 592.050 630.150 ;
        RECT 592.950 628.950 595.050 631.050 ;
        RECT 595.950 629.250 597.750 630.150 ;
        RECT 598.950 628.950 601.050 631.050 ;
        RECT 604.950 630.450 607.050 631.050 ;
        RECT 608.400 630.450 609.450 635.400 ;
        RECT 602.250 629.250 603.750 630.150 ;
        RECT 604.950 629.400 609.450 630.450 ;
        RECT 604.950 628.950 607.050 629.400 ;
        RECT 589.950 625.950 592.050 628.050 ;
        RECT 593.400 627.450 594.450 628.950 ;
        RECT 595.950 627.450 598.050 628.050 ;
        RECT 593.400 626.400 598.050 627.450 ;
        RECT 599.250 626.850 600.750 627.750 ;
        RECT 595.950 625.950 598.050 626.400 ;
        RECT 601.950 625.950 604.050 628.050 ;
        RECT 607.950 619.950 610.050 622.050 ;
        RECT 586.950 616.950 589.050 619.050 ;
        RECT 583.950 610.950 586.050 613.050 ;
        RECT 586.950 607.950 589.050 610.050 ;
        RECT 580.950 605.400 583.050 607.500 ;
        RECT 581.400 588.600 582.600 605.400 ;
        RECT 583.950 604.950 586.050 607.050 ;
        RECT 584.400 598.050 585.450 604.950 ;
        RECT 587.400 601.050 588.450 607.950 ;
        RECT 601.950 605.400 604.050 607.500 ;
        RECT 592.950 601.950 595.050 604.050 ;
        RECT 593.400 601.050 594.450 601.950 ;
        RECT 586.950 598.950 589.050 601.050 ;
        RECT 592.950 600.450 595.050 601.050 ;
        RECT 592.950 599.400 597.450 600.450 ;
        RECT 592.950 598.950 595.050 599.400 ;
        RECT 583.950 595.950 586.050 598.050 ;
        RECT 586.950 596.850 589.050 597.750 ;
        RECT 589.950 595.950 592.050 598.050 ;
        RECT 592.950 596.850 595.050 597.750 ;
        RECT 580.950 586.500 583.050 588.600 ;
        RECT 580.950 580.950 583.050 583.050 ;
        RECT 583.950 580.950 586.050 583.050 ;
        RECT 581.400 553.050 582.450 580.950 ;
        RECT 580.950 550.950 583.050 553.050 ;
        RECT 577.950 541.950 580.050 544.050 ;
        RECT 574.950 535.950 577.050 538.050 ;
        RECT 577.950 533.400 580.050 535.500 ;
        RECT 574.950 530.250 577.050 531.150 ;
        RECT 574.950 526.950 577.050 529.050 ;
        RECT 575.400 523.050 576.450 526.950 ;
        RECT 574.950 520.950 577.050 523.050 ;
        RECT 578.550 521.400 579.750 533.400 ;
        RECT 580.950 532.950 583.050 535.050 ;
        RECT 560.400 503.400 564.450 504.450 ;
        RECT 566.400 518.400 570.450 519.450 ;
        RECT 553.950 499.950 556.050 502.050 ;
        RECT 556.950 496.950 559.050 499.050 ;
        RECT 544.950 490.950 547.050 493.050 ;
        RECT 550.950 491.250 553.050 492.150 ;
        RECT 545.400 490.050 546.450 490.950 ;
        RECT 557.400 490.050 558.450 496.950 ;
        RECT 541.950 487.950 544.050 490.050 ;
        RECT 544.950 487.950 547.050 490.050 ;
        RECT 548.250 488.250 549.750 489.150 ;
        RECT 550.950 487.950 553.050 490.050 ;
        RECT 554.250 488.250 556.050 489.150 ;
        RECT 556.950 487.950 559.050 490.050 ;
        RECT 526.950 484.950 529.050 487.050 ;
        RECT 529.950 485.250 531.750 486.150 ;
        RECT 532.950 484.950 535.050 487.050 ;
        RECT 538.950 484.950 541.050 487.050 ;
        RECT 527.400 469.050 528.450 484.950 ;
        RECT 529.950 481.950 532.050 484.050 ;
        RECT 533.250 482.850 535.050 483.750 ;
        RECT 535.950 482.250 538.050 483.150 ;
        RECT 538.950 482.850 541.050 483.750 ;
        RECT 542.400 483.450 543.450 487.950 ;
        RECT 544.950 485.850 546.750 486.750 ;
        RECT 547.950 484.950 550.050 487.050 ;
        RECT 551.400 484.050 552.450 487.950 ;
        RECT 560.400 487.050 561.450 503.400 ;
        RECT 562.950 496.950 565.050 499.050 ;
        RECT 563.400 493.050 564.450 496.950 ;
        RECT 562.950 490.950 565.050 493.050 ;
        RECT 553.950 484.950 556.050 487.050 ;
        RECT 556.950 485.250 559.050 486.150 ;
        RECT 559.950 484.950 562.050 487.050 ;
        RECT 562.950 485.250 565.050 486.150 ;
        RECT 542.400 482.400 546.450 483.450 ;
        RECT 530.400 481.050 531.450 481.950 ;
        RECT 529.950 478.950 532.050 481.050 ;
        RECT 535.950 478.950 538.050 481.050 ;
        RECT 538.950 478.950 541.050 481.050 ;
        RECT 539.400 472.050 540.450 478.950 ;
        RECT 538.950 469.950 541.050 472.050 ;
        RECT 541.950 469.950 544.050 472.050 ;
        RECT 526.950 466.950 529.050 469.050 ;
        RECT 523.950 463.950 526.050 466.050 ;
        RECT 517.950 460.950 520.050 463.050 ;
        RECT 532.950 460.950 535.050 463.050 ;
        RECT 514.950 457.950 517.050 460.050 ;
        RECT 506.400 455.400 510.450 456.450 ;
        RECT 493.950 452.250 495.750 453.150 ;
        RECT 496.950 451.950 499.050 454.050 ;
        RECT 500.250 452.250 502.050 453.150 ;
        RECT 502.950 451.950 505.050 454.050 ;
        RECT 506.400 451.050 507.450 455.400 ;
        RECT 511.950 454.950 514.050 457.050 ;
        RECT 508.950 451.950 511.050 454.050 ;
        RECT 512.250 452.250 514.050 453.150 ;
        RECT 493.950 448.950 496.050 451.050 ;
        RECT 497.250 449.850 498.750 450.750 ;
        RECT 499.950 448.950 502.050 451.050 ;
        RECT 502.950 449.850 504.750 450.750 ;
        RECT 505.950 448.950 508.050 451.050 ;
        RECT 509.250 449.850 510.750 450.750 ;
        RECT 511.950 448.950 514.050 451.050 ;
        RECT 500.400 448.050 501.450 448.950 ;
        RECT 499.950 445.950 502.050 448.050 ;
        RECT 505.950 446.850 508.050 447.750 ;
        RECT 512.400 445.050 513.450 448.950 ;
        RECT 511.950 442.950 514.050 445.050 ;
        RECT 493.950 439.950 496.050 442.050 ;
        RECT 490.950 430.950 493.050 433.050 ;
        RECT 478.950 424.950 481.050 427.050 ;
        RECT 469.950 421.950 472.050 424.050 ;
        RECT 475.950 421.950 478.050 424.050 ;
        RECT 470.400 415.050 471.450 421.950 ;
        RECT 469.950 412.950 472.050 415.050 ;
        RECT 469.950 410.850 472.050 411.750 ;
        RECT 472.950 410.250 475.050 411.150 ;
        RECT 472.950 408.450 475.050 409.050 ;
        RECT 476.400 408.450 477.450 421.950 ;
        RECT 490.950 418.950 493.050 421.050 ;
        RECT 478.950 416.250 481.050 417.150 ;
        RECT 478.950 412.950 481.050 415.050 ;
        RECT 482.250 413.250 483.750 414.150 ;
        RECT 484.950 412.950 487.050 415.050 ;
        RECT 488.250 413.250 490.050 414.150 ;
        RECT 481.950 409.950 484.050 412.050 ;
        RECT 485.250 410.850 486.750 411.750 ;
        RECT 487.950 409.950 490.050 412.050 ;
        RECT 472.950 407.400 477.450 408.450 ;
        RECT 472.950 406.950 475.050 407.400 ;
        RECT 466.950 400.950 469.050 403.050 ;
        RECT 460.950 397.950 463.050 400.050 ;
        RECT 466.950 394.950 469.050 397.050 ;
        RECT 457.950 382.950 460.050 385.050 ;
        RECT 461.250 383.250 462.750 384.150 ;
        RECT 463.950 382.950 466.050 385.050 ;
        RECT 458.250 380.850 459.750 381.750 ;
        RECT 460.950 379.950 463.050 382.050 ;
        RECT 464.250 380.850 466.050 381.750 ;
        RECT 451.950 376.950 454.050 379.050 ;
        RECT 454.950 377.850 457.050 378.750 ;
        RECT 448.950 364.950 451.050 367.050 ;
        RECT 451.950 358.950 454.050 361.050 ;
        RECT 445.950 349.950 448.050 352.050 ;
        RECT 452.400 346.050 453.450 358.950 ;
        RECT 461.400 358.050 462.450 379.950 ;
        RECT 463.950 370.950 466.050 373.050 ;
        RECT 460.950 355.950 463.050 358.050 ;
        RECT 445.950 343.950 448.050 346.050 ;
        RECT 449.250 344.250 450.750 345.150 ;
        RECT 451.950 343.950 454.050 346.050 ;
        RECT 454.950 345.450 457.050 346.050 ;
        RECT 457.950 345.450 460.050 346.050 ;
        RECT 454.950 344.400 460.050 345.450 ;
        RECT 454.950 343.950 457.050 344.400 ;
        RECT 457.950 343.950 460.050 344.400 ;
        RECT 464.400 343.050 465.450 370.950 ;
        RECT 467.400 349.050 468.450 394.950 ;
        RECT 476.400 391.050 477.450 407.400 ;
        RECT 488.400 403.050 489.450 409.950 ;
        RECT 487.950 400.950 490.050 403.050 ;
        RECT 491.400 391.050 492.450 418.950 ;
        RECT 494.400 406.050 495.450 439.950 ;
        RECT 499.950 430.950 502.050 433.050 ;
        RECT 496.950 421.950 499.050 424.050 ;
        RECT 497.400 414.900 498.450 421.950 ;
        RECT 496.950 412.800 499.050 414.900 ;
        RECT 496.950 410.700 499.050 411.600 ;
        RECT 493.950 403.950 496.050 406.050 ;
        RECT 500.400 402.450 501.450 430.950 ;
        RECT 512.400 418.050 513.450 442.950 ;
        RECT 505.950 415.950 508.050 418.050 ;
        RECT 511.950 415.950 514.050 418.050 ;
        RECT 506.400 414.900 507.450 415.950 ;
        RECT 502.950 413.100 504.750 414.000 ;
        RECT 505.950 412.800 508.050 414.900 ;
        RECT 508.950 412.950 511.050 415.050 ;
        RECT 511.950 413.100 514.050 414.000 ;
        RECT 502.950 409.800 505.050 412.050 ;
        RECT 506.250 410.700 508.050 411.600 ;
        RECT 505.950 406.950 508.050 409.050 ;
        RECT 497.400 401.400 501.450 402.450 ;
        RECT 475.950 388.950 478.050 391.050 ;
        RECT 487.950 388.950 490.050 391.050 ;
        RECT 490.950 388.950 493.050 391.050 ;
        RECT 475.950 385.950 478.050 388.050 ;
        RECT 484.950 385.950 487.050 388.050 ;
        RECT 469.950 382.950 472.050 385.050 ;
        RECT 473.250 383.250 475.050 384.150 ;
        RECT 475.950 383.850 478.050 384.750 ;
        RECT 478.950 383.250 481.050 384.150 ;
        RECT 469.950 380.850 471.750 381.750 ;
        RECT 472.950 379.950 475.050 382.050 ;
        RECT 478.950 381.450 481.050 382.050 ;
        RECT 481.950 381.450 484.050 382.050 ;
        RECT 478.950 380.400 484.050 381.450 ;
        RECT 478.950 379.950 481.050 380.400 ;
        RECT 481.950 379.950 484.050 380.400 ;
        RECT 479.400 355.050 480.450 379.950 ;
        RECT 485.400 379.050 486.450 385.950 ;
        RECT 488.400 382.050 489.450 388.950 ;
        RECT 493.950 385.950 496.050 388.050 ;
        RECT 487.950 379.950 490.050 382.050 ;
        RECT 491.250 380.250 493.050 381.150 ;
        RECT 481.950 377.850 483.750 378.750 ;
        RECT 484.950 376.950 487.050 379.050 ;
        RECT 488.250 377.850 489.750 378.750 ;
        RECT 490.950 378.450 493.050 379.050 ;
        RECT 494.400 378.450 495.450 385.950 ;
        RECT 490.950 377.400 495.450 378.450 ;
        RECT 490.950 376.950 493.050 377.400 ;
        RECT 484.950 374.850 487.050 375.750 ;
        RECT 490.950 373.950 493.050 376.050 ;
        RECT 481.950 370.950 484.050 373.050 ;
        RECT 478.950 352.950 481.050 355.050 ;
        RECT 466.950 346.950 469.050 349.050 ;
        RECT 472.950 346.950 475.050 349.050 ;
        RECT 475.950 346.950 478.050 349.050 ;
        RECT 473.400 346.050 474.450 346.950 ;
        RECT 466.950 343.950 469.050 346.050 ;
        RECT 470.250 344.250 471.750 345.150 ;
        RECT 472.950 343.950 475.050 346.050 ;
        RECT 476.400 343.050 477.450 346.950 ;
        RECT 482.400 343.050 483.450 370.950 ;
        RECT 484.950 355.950 487.050 358.050 ;
        RECT 485.400 346.050 486.450 355.950 ;
        RECT 487.950 349.950 490.050 352.050 ;
        RECT 484.950 343.950 487.050 346.050 ;
        RECT 434.250 341.250 435.750 342.150 ;
        RECT 436.950 341.400 441.450 342.450 ;
        RECT 436.950 340.950 439.050 341.400 ;
        RECT 442.950 340.950 445.050 343.050 ;
        RECT 445.950 341.850 447.750 342.750 ;
        RECT 448.950 340.950 451.050 343.050 ;
        RECT 452.250 341.850 454.050 342.750 ;
        RECT 454.950 340.950 457.050 343.050 ;
        RECT 460.950 342.450 463.050 343.050 ;
        RECT 458.400 341.400 463.050 342.450 ;
        RECT 421.950 338.850 424.050 339.750 ;
        RECT 424.950 338.250 427.050 339.150 ;
        RECT 427.950 337.950 430.050 340.050 ;
        RECT 431.250 338.850 432.750 339.750 ;
        RECT 433.950 337.950 436.050 340.050 ;
        RECT 421.950 334.950 424.050 337.050 ;
        RECT 424.950 334.950 427.050 337.050 ;
        RECT 422.400 316.050 423.450 334.950 ;
        RECT 428.400 330.450 429.450 337.950 ;
        RECT 425.400 329.400 429.450 330.450 ;
        RECT 418.950 313.950 421.050 316.050 ;
        RECT 421.950 313.950 424.050 316.050 ;
        RECT 425.400 313.050 426.450 329.400 ;
        RECT 427.950 325.950 430.050 328.050 ;
        RECT 418.950 310.950 421.050 313.050 ;
        RECT 422.250 311.250 423.750 312.150 ;
        RECT 424.950 310.950 427.050 313.050 ;
        RECT 412.950 307.950 415.050 310.050 ;
        RECT 415.950 307.950 418.050 310.050 ;
        RECT 419.250 308.850 420.750 309.750 ;
        RECT 421.950 307.950 424.050 310.050 ;
        RECT 425.250 308.850 427.050 309.750 ;
        RECT 409.950 304.950 412.050 307.050 ;
        RECT 397.950 292.950 400.050 295.050 ;
        RECT 413.400 292.050 414.450 307.950 ;
        RECT 415.950 305.850 418.050 306.750 ;
        RECT 406.950 289.950 409.050 292.050 ;
        RECT 412.950 289.950 415.050 292.050 ;
        RECT 403.950 274.950 406.050 277.050 ;
        RECT 404.400 274.050 405.450 274.950 ;
        RECT 403.950 271.950 406.050 274.050 ;
        RECT 400.950 269.250 403.050 270.150 ;
        RECT 403.950 269.850 406.050 270.750 ;
        RECT 400.950 265.950 403.050 268.050 ;
        RECT 401.400 259.050 402.450 265.950 ;
        RECT 400.950 256.950 403.050 259.050 ;
        RECT 394.950 250.950 397.050 253.050 ;
        RECT 400.950 250.950 403.050 253.050 ;
        RECT 392.400 248.400 396.450 249.450 ;
        RECT 391.950 244.950 394.050 247.050 ;
        RECT 392.400 241.050 393.450 244.950 ;
        RECT 391.950 238.950 394.050 241.050 ;
        RECT 395.400 238.050 396.450 248.400 ;
        RECT 401.400 238.050 402.450 250.950 ;
        RECT 388.950 236.250 391.050 237.150 ;
        RECT 391.950 236.850 394.050 237.750 ;
        RECT 394.950 235.950 397.050 238.050 ;
        RECT 397.950 236.250 399.750 237.150 ;
        RECT 400.950 235.950 403.050 238.050 ;
        RECT 404.250 236.250 406.050 237.150 ;
        RECT 388.950 232.950 391.050 235.050 ;
        RECT 397.950 232.950 400.050 235.050 ;
        RECT 401.250 233.850 402.750 234.750 ;
        RECT 403.950 232.950 406.050 235.050 ;
        RECT 379.950 220.950 382.050 223.050 ;
        RECT 385.950 220.950 388.050 223.050 ;
        RECT 385.950 217.950 388.050 220.050 ;
        RECT 386.400 214.050 387.450 217.950 ;
        RECT 398.400 217.050 399.450 232.950 ;
        RECT 404.400 232.050 405.450 232.950 ;
        RECT 403.950 229.950 406.050 232.050 ;
        RECT 407.400 231.450 408.450 289.950 ;
        RECT 422.400 280.050 423.450 307.950 ;
        RECT 421.950 277.950 424.050 280.050 ;
        RECT 412.950 274.950 415.050 277.050 ;
        RECT 413.400 271.050 414.450 274.950 ;
        RECT 409.950 269.250 412.050 270.150 ;
        RECT 412.950 268.950 415.050 271.050 ;
        RECT 416.250 269.250 418.050 270.150 ;
        RECT 424.950 269.250 427.050 270.150 ;
        RECT 428.400 268.050 429.450 325.950 ;
        RECT 434.400 312.450 435.450 337.950 ;
        RECT 451.950 334.950 454.050 337.050 ;
        RECT 445.950 331.950 448.050 334.050 ;
        RECT 442.950 325.950 445.050 328.050 ;
        RECT 443.400 322.050 444.450 325.950 ;
        RECT 442.950 319.950 445.050 322.050 ;
        RECT 442.950 316.950 445.050 319.050 ;
        RECT 443.400 316.050 444.450 316.950 ;
        RECT 436.950 313.950 439.050 316.050 ;
        RECT 442.950 313.950 445.050 316.050 ;
        RECT 446.400 315.450 447.450 331.950 ;
        RECT 452.400 331.050 453.450 334.950 ;
        RECT 455.400 334.050 456.450 340.950 ;
        RECT 458.400 336.450 459.450 341.400 ;
        RECT 460.950 340.950 463.050 341.400 ;
        RECT 463.950 340.950 466.050 343.050 ;
        RECT 466.950 341.850 468.750 342.750 ;
        RECT 469.950 340.950 472.050 343.050 ;
        RECT 473.250 341.850 475.050 342.750 ;
        RECT 475.950 340.950 478.050 343.050 ;
        RECT 478.950 341.250 481.050 342.150 ;
        RECT 481.950 340.950 484.050 343.050 ;
        RECT 484.950 341.250 487.050 342.150 ;
        RECT 460.950 338.850 463.050 339.750 ;
        RECT 463.950 338.250 466.050 339.150 ;
        RECT 466.950 337.950 469.050 340.050 ;
        RECT 472.950 337.950 475.050 340.050 ;
        RECT 475.950 337.950 478.050 340.050 ;
        RECT 478.950 337.950 481.050 340.050 ;
        RECT 482.250 338.250 483.750 339.150 ;
        RECT 484.950 337.950 487.050 340.050 ;
        RECT 458.400 335.400 462.450 336.450 ;
        RECT 454.950 331.950 457.050 334.050 ;
        RECT 448.950 328.950 451.050 331.050 ;
        RECT 451.950 328.950 454.050 331.050 ;
        RECT 461.400 330.450 462.450 335.400 ;
        RECT 463.950 334.950 466.050 337.050 ;
        RECT 464.400 334.050 465.450 334.950 ;
        RECT 463.950 331.950 466.050 334.050 ;
        RECT 461.400 329.400 465.450 330.450 ;
        RECT 449.400 322.050 450.450 328.950 ;
        RECT 464.400 325.050 465.450 329.400 ;
        RECT 460.950 322.950 463.050 325.050 ;
        RECT 463.950 322.950 466.050 325.050 ;
        RECT 448.950 319.950 451.050 322.050 ;
        RECT 446.400 314.400 450.450 315.450 ;
        RECT 431.400 311.400 435.450 312.450 ;
        RECT 431.400 310.050 432.450 311.400 ;
        RECT 437.400 310.050 438.450 313.950 ;
        RECT 442.950 311.850 445.050 312.750 ;
        RECT 445.950 311.250 448.050 312.150 ;
        RECT 430.950 307.950 433.050 310.050 ;
        RECT 433.950 308.250 435.750 309.150 ;
        RECT 436.950 307.950 439.050 310.050 ;
        RECT 440.250 308.250 442.050 309.150 ;
        RECT 445.950 307.950 448.050 310.050 ;
        RECT 446.400 307.050 447.450 307.950 ;
        RECT 430.950 304.950 433.050 307.050 ;
        RECT 433.950 304.950 436.050 307.050 ;
        RECT 437.250 305.850 438.750 306.750 ;
        RECT 439.950 304.950 442.050 307.050 ;
        RECT 445.950 304.950 448.050 307.050 ;
        RECT 431.400 274.050 432.450 304.950 ;
        RECT 434.400 300.450 435.450 304.950 ;
        RECT 434.400 299.400 438.450 300.450 ;
        RECT 433.950 295.950 436.050 298.050 ;
        RECT 430.950 271.950 433.050 274.050 ;
        RECT 430.950 269.250 433.050 270.150 ;
        RECT 409.950 265.950 412.050 268.050 ;
        RECT 412.950 266.850 414.750 267.750 ;
        RECT 415.950 265.950 418.050 268.050 ;
        RECT 424.950 265.950 427.050 268.050 ;
        RECT 427.950 265.950 430.050 268.050 ;
        RECT 430.950 265.950 433.050 268.050 ;
        RECT 410.400 256.050 411.450 265.950 ;
        RECT 409.950 253.950 412.050 256.050 ;
        RECT 416.400 250.050 417.450 265.950 ;
        RECT 425.400 262.050 426.450 265.950 ;
        RECT 424.950 259.950 427.050 262.050 ;
        RECT 421.950 256.950 424.050 259.050 ;
        RECT 409.950 247.950 412.050 250.050 ;
        RECT 415.950 247.950 418.050 250.050 ;
        RECT 410.400 235.050 411.450 247.950 ;
        RECT 412.950 241.950 415.050 244.050 ;
        RECT 413.400 238.050 414.450 241.950 ;
        RECT 422.400 241.050 423.450 256.950 ;
        RECT 431.400 253.050 432.450 265.950 ;
        RECT 430.950 250.950 433.050 253.050 ;
        RECT 427.950 247.950 430.050 250.050 ;
        RECT 415.950 238.950 418.050 241.050 ;
        RECT 419.250 239.250 420.750 240.150 ;
        RECT 421.950 238.950 424.050 241.050 ;
        RECT 428.400 238.050 429.450 247.950 ;
        RECT 412.950 235.950 415.050 238.050 ;
        RECT 416.250 236.850 417.750 237.750 ;
        RECT 418.950 235.950 421.050 238.050 ;
        RECT 422.250 236.850 424.050 237.750 ;
        RECT 424.950 236.250 426.750 237.150 ;
        RECT 427.950 235.950 430.050 238.050 ;
        RECT 431.250 236.250 433.050 237.150 ;
        RECT 419.400 235.050 420.450 235.950 ;
        RECT 409.950 232.950 412.050 235.050 ;
        RECT 412.950 233.850 415.050 234.750 ;
        RECT 415.950 232.950 418.050 235.050 ;
        RECT 418.950 232.950 421.050 235.050 ;
        RECT 424.950 232.950 427.050 235.050 ;
        RECT 428.250 233.850 429.750 234.750 ;
        RECT 430.950 232.950 433.050 235.050 ;
        RECT 407.400 230.400 411.450 231.450 ;
        RECT 406.950 223.950 409.050 226.050 ;
        RECT 397.950 214.950 400.050 217.050 ;
        RECT 400.950 214.950 403.050 217.050 ;
        RECT 385.950 211.950 388.050 214.050 ;
        RECT 401.400 211.050 402.450 214.950 ;
        RECT 400.950 208.950 403.050 211.050 ;
        RECT 403.950 208.950 406.050 211.050 ;
        RECT 382.950 202.950 385.050 205.050 ;
        RECT 388.950 202.950 391.050 205.050 ;
        RECT 400.950 204.450 403.050 205.050 ;
        RECT 404.400 204.450 405.450 208.950 ;
        RECT 407.400 208.050 408.450 223.950 ;
        RECT 406.950 205.950 409.050 208.050 ;
        RECT 400.950 203.400 405.450 204.450 ;
        RECT 400.950 202.950 403.050 203.400 ;
        RECT 383.400 202.050 384.450 202.950 ;
        RECT 370.950 200.250 373.050 201.150 ;
        RECT 373.950 199.950 376.050 202.050 ;
        RECT 376.950 199.950 379.050 202.050 ;
        RECT 382.950 199.950 385.050 202.050 ;
        RECT 377.400 199.050 378.450 199.950 ;
        RECT 389.400 199.050 390.450 202.950 ;
        RECT 400.950 199.950 403.050 202.050 ;
        RECT 401.400 199.050 402.450 199.950 ;
        RECT 407.400 199.050 408.450 205.950 ;
        RECT 370.950 198.450 373.050 199.050 ;
        RECT 368.400 197.400 373.050 198.450 ;
        RECT 370.950 196.950 373.050 197.400 ;
        RECT 374.250 197.250 375.750 198.150 ;
        RECT 376.950 196.950 379.050 199.050 ;
        RECT 380.250 197.250 382.050 198.150 ;
        RECT 382.950 196.950 385.050 199.050 ;
        RECT 385.950 197.250 388.050 198.150 ;
        RECT 388.950 196.950 391.050 199.050 ;
        RECT 391.950 197.250 394.050 198.150 ;
        RECT 397.950 197.250 399.750 198.150 ;
        RECT 400.950 196.950 403.050 199.050 ;
        RECT 406.950 196.950 409.050 199.050 ;
        RECT 358.950 193.950 361.050 196.050 ;
        RECT 364.950 193.950 367.050 196.050 ;
        RECT 367.950 193.950 370.050 196.050 ;
        RECT 373.950 193.950 376.050 196.050 ;
        RECT 377.250 194.850 378.750 195.750 ;
        RECT 379.950 193.950 382.050 196.050 ;
        RECT 355.950 190.950 358.050 193.050 ;
        RECT 350.400 185.400 354.450 186.450 ;
        RECT 341.400 181.050 342.450 184.950 ;
        RECT 340.950 178.950 343.050 181.050 ;
        RECT 350.400 178.050 351.450 185.400 ;
        RECT 352.950 181.950 355.050 184.050 ;
        RECT 349.950 175.950 352.050 178.050 ;
        RECT 346.950 172.950 349.050 175.050 ;
        RECT 347.400 172.050 348.450 172.950 ;
        RECT 346.950 169.950 349.050 172.050 ;
        RECT 326.400 167.400 330.450 168.450 ;
        RECT 326.400 166.050 327.450 167.400 ;
        RECT 331.950 166.950 334.050 169.050 ;
        RECT 334.950 166.950 337.050 169.050 ;
        RECT 346.950 167.850 349.050 168.750 ;
        RECT 349.950 167.250 352.050 168.150 ;
        RECT 289.950 163.950 292.050 166.050 ;
        RECT 293.250 164.850 294.750 165.750 ;
        RECT 295.950 163.950 298.050 166.050 ;
        RECT 299.250 164.850 301.050 165.750 ;
        RECT 304.950 163.950 307.050 166.050 ;
        RECT 307.950 163.950 310.050 166.050 ;
        RECT 313.950 163.950 316.050 166.050 ;
        RECT 319.950 163.950 322.050 166.050 ;
        RECT 325.950 163.950 328.050 166.050 ;
        RECT 329.250 164.250 331.050 165.150 ;
        RECT 305.400 163.050 306.450 163.950 ;
        RECT 289.950 161.850 292.050 162.750 ;
        RECT 304.950 160.950 307.050 163.050 ;
        RECT 319.950 161.850 321.750 162.750 ;
        RECT 322.950 160.950 325.050 163.050 ;
        RECT 326.250 161.850 327.750 162.750 ;
        RECT 328.950 160.950 331.050 163.050 ;
        RECT 322.950 158.850 325.050 159.750 ;
        RECT 283.950 154.950 286.050 157.050 ;
        RECT 284.400 130.050 285.450 154.950 ;
        RECT 313.950 142.950 316.050 145.050 ;
        RECT 329.400 144.450 330.450 160.950 ;
        RECT 332.400 157.050 333.450 166.950 ;
        RECT 334.950 163.950 337.050 166.050 ;
        RECT 337.950 164.250 339.750 165.150 ;
        RECT 340.950 163.950 343.050 166.050 ;
        RECT 344.250 164.250 346.050 165.150 ;
        RECT 346.950 163.950 349.050 166.050 ;
        RECT 349.950 163.950 352.050 166.050 ;
        RECT 331.950 154.950 334.050 157.050 ;
        RECT 326.400 143.400 330.450 144.450 ;
        RECT 314.400 133.050 315.450 142.950 ;
        RECT 326.400 133.050 327.450 143.400 ;
        RECT 328.950 139.950 331.050 142.050 ;
        RECT 331.950 139.950 334.050 142.050 ;
        RECT 329.400 136.050 330.450 139.950 ;
        RECT 328.950 133.950 331.050 136.050 ;
        RECT 332.400 133.050 333.450 139.950 ;
        RECT 335.400 139.050 336.450 163.950 ;
        RECT 337.950 160.950 340.050 163.050 ;
        RECT 341.250 161.850 342.750 162.750 ;
        RECT 343.950 160.950 346.050 163.050 ;
        RECT 338.400 160.050 339.450 160.950 ;
        RECT 337.950 157.950 340.050 160.050 ;
        RECT 334.950 136.950 337.050 139.050 ;
        RECT 337.950 135.450 340.050 136.050 ;
        RECT 340.950 135.450 343.050 136.050 ;
        RECT 337.950 134.400 343.050 135.450 ;
        RECT 337.950 133.950 340.050 134.400 ;
        RECT 340.950 133.950 343.050 134.400 ;
        RECT 307.950 130.950 310.050 133.050 ;
        RECT 313.950 130.950 316.050 133.050 ;
        RECT 325.950 130.950 328.050 133.050 ;
        RECT 331.950 130.950 334.050 133.050 ;
        RECT 337.950 130.950 340.050 133.050 ;
        RECT 283.950 127.950 286.050 130.050 ;
        RECT 286.950 128.250 289.050 129.150 ;
        RECT 283.950 124.950 286.050 127.050 ;
        RECT 286.950 124.950 289.050 127.050 ;
        RECT 290.250 125.250 291.750 126.150 ;
        RECT 292.950 124.950 295.050 127.050 ;
        RECT 296.250 125.250 298.050 126.150 ;
        RECT 298.950 125.250 301.050 126.150 ;
        RECT 304.950 125.250 307.050 126.150 ;
        RECT 284.400 115.050 285.450 124.950 ;
        RECT 287.400 118.050 288.450 124.950 ;
        RECT 289.950 121.950 292.050 124.050 ;
        RECT 293.250 122.850 294.750 123.750 ;
        RECT 295.950 121.950 298.050 124.050 ;
        RECT 298.950 121.950 301.050 124.050 ;
        RECT 302.250 122.250 303.750 123.150 ;
        RECT 304.950 121.950 307.050 124.050 ;
        RECT 286.950 115.950 289.050 118.050 ;
        RECT 283.950 112.950 286.050 115.050 ;
        RECT 290.400 112.050 291.450 121.950 ;
        RECT 296.400 121.050 297.450 121.950 ;
        RECT 295.950 118.950 298.050 121.050 ;
        RECT 301.950 118.950 304.050 121.050 ;
        RECT 302.400 115.050 303.450 118.950 ;
        RECT 305.400 115.050 306.450 121.950 ;
        RECT 308.400 115.050 309.450 130.950 ;
        RECT 314.400 130.050 315.450 130.950 ;
        RECT 310.950 127.950 313.050 130.050 ;
        RECT 313.950 127.950 316.050 130.050 ;
        RECT 317.250 128.250 318.750 129.150 ;
        RECT 319.950 127.950 322.050 130.050 ;
        RECT 322.950 127.950 325.050 130.050 ;
        RECT 328.950 129.450 331.050 130.050 ;
        RECT 326.250 128.250 327.750 129.150 ;
        RECT 328.950 128.400 333.450 129.450 ;
        RECT 328.950 127.950 331.050 128.400 ;
        RECT 311.400 124.050 312.450 127.950 ;
        RECT 313.950 125.850 315.750 126.750 ;
        RECT 316.950 124.950 319.050 127.050 ;
        RECT 320.250 125.850 322.050 126.750 ;
        RECT 322.950 125.850 324.750 126.750 ;
        RECT 325.950 124.950 328.050 127.050 ;
        RECT 329.250 125.850 331.050 126.750 ;
        RECT 310.950 121.950 313.050 124.050 ;
        RECT 317.400 118.050 318.450 124.950 ;
        RECT 316.950 115.950 319.050 118.050 ;
        RECT 301.950 112.950 304.050 115.050 ;
        RECT 304.950 112.950 307.050 115.050 ;
        RECT 307.950 112.950 310.050 115.050 ;
        RECT 317.400 112.050 318.450 115.950 ;
        RECT 283.950 109.950 286.050 112.050 ;
        RECT 289.950 109.950 292.050 112.050 ;
        RECT 316.950 109.950 319.050 112.050 ;
        RECT 280.950 103.950 283.050 106.050 ;
        RECT 278.400 101.400 282.450 102.450 ;
        RECT 275.400 100.050 276.450 100.950 ;
        RECT 274.950 97.950 277.050 100.050 ;
        RECT 277.950 97.950 280.050 100.050 ;
        RECT 259.950 92.850 262.050 93.750 ;
        RECT 262.950 91.950 265.050 94.050 ;
        RECT 265.950 91.950 268.050 94.050 ;
        RECT 268.950 92.250 270.750 93.150 ;
        RECT 271.950 91.950 274.050 94.050 ;
        RECT 259.950 85.950 262.050 88.050 ;
        RECT 256.950 82.950 259.050 85.050 ;
        RECT 244.950 67.950 247.050 70.050 ;
        RECT 250.950 67.950 253.050 70.050 ;
        RECT 253.950 67.950 256.050 70.050 ;
        RECT 245.400 58.050 246.450 67.950 ;
        RECT 250.950 61.950 253.050 64.050 ;
        RECT 199.950 55.950 202.050 58.050 ;
        RECT 205.950 57.450 208.050 58.050 ;
        RECT 203.250 56.250 204.750 57.150 ;
        RECT 205.950 56.400 210.450 57.450 ;
        RECT 205.950 55.950 208.050 56.400 ;
        RECT 187.950 53.400 192.450 54.450 ;
        RECT 193.950 54.450 196.050 55.050 ;
        RECT 193.950 53.400 198.450 54.450 ;
        RECT 199.950 53.850 201.750 54.750 ;
        RECT 187.950 52.950 190.050 53.400 ;
        RECT 193.950 52.950 196.050 53.400 ;
        RECT 188.400 48.450 189.450 52.950 ;
        RECT 190.950 50.250 193.050 51.150 ;
        RECT 193.950 50.850 196.050 51.750 ;
        RECT 190.950 48.450 193.050 49.050 ;
        RECT 188.400 47.400 193.050 48.450 ;
        RECT 190.950 46.950 193.050 47.400 ;
        RECT 184.950 40.950 187.050 43.050 ;
        RECT 197.400 31.050 198.450 53.400 ;
        RECT 202.950 52.950 205.050 55.050 ;
        RECT 206.250 53.850 208.050 54.750 ;
        RECT 209.400 54.450 210.450 56.400 ;
        RECT 211.950 56.250 213.750 57.150 ;
        RECT 214.950 55.950 217.050 58.050 ;
        RECT 218.250 56.250 219.750 57.150 ;
        RECT 220.950 55.950 223.050 58.050 ;
        RECT 226.950 55.950 229.050 58.050 ;
        RECT 232.950 57.450 235.050 58.050 ;
        RECT 230.250 56.250 231.750 57.150 ;
        RECT 232.950 56.400 237.450 57.450 ;
        RECT 232.950 55.950 235.050 56.400 ;
        RECT 211.950 54.450 214.050 55.050 ;
        RECT 209.400 53.400 214.050 54.450 ;
        RECT 211.950 52.950 214.050 53.400 ;
        RECT 217.950 52.950 220.050 55.050 ;
        RECT 221.250 53.850 223.050 54.750 ;
        RECT 226.950 53.850 228.750 54.750 ;
        RECT 229.950 52.950 232.050 55.050 ;
        RECT 233.250 53.850 235.050 54.750 ;
        RECT 202.950 34.950 205.050 37.050 ;
        RECT 196.950 28.950 199.050 31.050 ;
        RECT 184.950 25.950 187.050 28.050 ;
        RECT 190.950 25.950 193.050 28.050 ;
        RECT 169.950 22.950 172.050 25.050 ;
        RECT 173.250 23.250 174.750 24.150 ;
        RECT 175.950 22.950 178.050 25.050 ;
        RECT 185.400 22.050 186.450 25.950 ;
        RECT 191.400 22.050 192.450 25.950 ;
        RECT 109.950 20.850 111.750 21.750 ;
        RECT 112.950 19.950 115.050 22.050 ;
        RECT 118.950 19.950 121.050 22.050 ;
        RECT 121.950 19.950 124.050 22.050 ;
        RECT 127.950 19.950 130.050 22.050 ;
        RECT 131.250 20.250 133.050 21.150 ;
        RECT 139.950 19.950 142.050 22.050 ;
        RECT 143.250 20.850 144.750 21.750 ;
        RECT 145.950 19.950 148.050 22.050 ;
        RECT 149.250 20.850 151.050 21.750 ;
        RECT 151.950 20.850 153.750 21.750 ;
        RECT 154.950 19.950 157.050 22.050 ;
        RECT 158.250 20.850 159.750 21.750 ;
        RECT 160.950 19.950 163.050 22.050 ;
        RECT 163.950 19.950 166.050 22.050 ;
        RECT 169.950 20.850 171.750 21.750 ;
        RECT 172.950 19.950 175.050 22.050 ;
        RECT 176.250 20.850 177.750 21.750 ;
        RECT 178.950 19.950 181.050 22.050 ;
        RECT 184.950 19.950 187.050 22.050 ;
        RECT 190.950 19.950 193.050 22.050 ;
        RECT 197.400 21.450 198.450 28.950 ;
        RECT 199.950 21.450 202.050 22.050 ;
        RECT 194.250 20.250 196.050 21.150 ;
        RECT 197.400 20.400 202.050 21.450 ;
        RECT 199.950 19.950 202.050 20.400 ;
        RECT 119.400 19.050 120.450 19.950 ;
        RECT 118.950 16.950 121.050 19.050 ;
        RECT 121.950 17.850 123.750 18.750 ;
        RECT 124.950 16.950 127.050 19.050 ;
        RECT 128.250 17.850 129.750 18.750 ;
        RECT 130.950 16.950 133.050 19.050 ;
        RECT 139.950 17.850 142.050 18.750 ;
        RECT 119.400 16.050 120.450 16.950 ;
        RECT 118.950 13.950 121.050 16.050 ;
        RECT 124.950 14.850 127.050 15.750 ;
        RECT 146.400 13.050 147.450 19.950 ;
        RECT 203.400 19.050 204.450 34.950 ;
        RECT 205.950 19.950 208.050 22.050 ;
        RECT 209.250 20.250 211.050 21.150 ;
        RECT 160.950 17.850 163.050 18.750 ;
        RECT 178.950 17.850 181.050 18.750 ;
        RECT 184.950 17.850 186.750 18.750 ;
        RECT 187.950 16.950 190.050 19.050 ;
        RECT 191.250 17.850 192.750 18.750 ;
        RECT 193.950 16.950 196.050 19.050 ;
        RECT 199.950 17.850 201.750 18.750 ;
        RECT 202.950 16.950 205.050 19.050 ;
        RECT 206.250 17.850 207.750 18.750 ;
        RECT 208.950 18.450 211.050 19.050 ;
        RECT 212.400 18.450 213.450 52.950 ;
        RECT 218.400 49.050 219.450 52.950 ;
        RECT 217.950 46.950 220.050 49.050 ;
        RECT 220.950 37.950 223.050 40.050 ;
        RECT 221.400 22.050 222.450 37.950 ;
        RECT 230.400 31.050 231.450 52.950 ;
        RECT 236.400 51.450 237.450 56.400 ;
        RECT 244.950 55.950 247.050 58.050 ;
        RECT 238.950 53.250 241.050 54.150 ;
        RECT 244.950 53.850 247.050 54.750 ;
        RECT 247.950 53.250 250.050 54.150 ;
        RECT 238.950 51.450 241.050 52.050 ;
        RECT 236.400 50.400 241.050 51.450 ;
        RECT 238.950 49.950 241.050 50.400 ;
        RECT 247.950 49.950 250.050 52.050 ;
        RECT 232.950 40.950 235.050 43.050 ;
        RECT 229.950 28.950 232.050 31.050 ;
        RECT 230.400 25.050 231.450 28.950 ;
        RECT 223.950 22.950 226.050 25.050 ;
        RECT 227.250 23.250 228.750 24.150 ;
        RECT 229.950 22.950 232.050 25.050 ;
        RECT 233.400 22.050 234.450 40.950 ;
        RECT 238.950 34.950 241.050 37.050 ;
        RECT 239.400 28.050 240.450 34.950 ;
        RECT 241.950 31.950 244.050 34.050 ;
        RECT 242.400 28.050 243.450 31.950 ;
        RECT 235.950 25.950 238.050 28.050 ;
        RECT 238.950 25.950 241.050 28.050 ;
        RECT 241.950 25.950 244.050 28.050 ;
        RECT 236.400 25.050 237.450 25.950 ;
        RECT 248.400 25.050 249.450 49.950 ;
        RECT 251.400 40.050 252.450 61.950 ;
        RECT 254.400 43.050 255.450 67.950 ;
        RECT 260.400 58.050 261.450 85.950 ;
        RECT 263.400 70.050 264.450 91.950 ;
        RECT 275.400 91.050 276.450 97.950 ;
        RECT 278.400 94.050 279.450 97.950 ;
        RECT 277.950 91.950 280.050 94.050 ;
        RECT 268.950 88.950 271.050 91.050 ;
        RECT 272.250 89.850 273.750 90.750 ;
        RECT 274.950 88.950 277.050 91.050 ;
        RECT 278.250 89.850 280.050 90.750 ;
        RECT 262.950 67.950 265.050 70.050 ;
        RECT 269.400 64.050 270.450 88.950 ;
        RECT 274.950 86.850 277.050 87.750 ;
        RECT 268.950 61.950 271.050 64.050 ;
        RECT 281.400 58.050 282.450 101.400 ;
        RECT 284.400 94.050 285.450 109.950 ;
        RECT 326.400 109.050 327.450 124.950 ;
        RECT 332.400 124.050 333.450 128.400 ;
        RECT 331.950 121.950 334.050 124.050 ;
        RECT 331.950 118.950 334.050 121.050 ;
        RECT 332.400 118.050 333.450 118.950 ;
        RECT 331.950 115.950 334.050 118.050 ;
        RECT 316.950 106.950 319.050 109.050 ;
        RECT 325.950 106.950 328.050 109.050 ;
        RECT 292.950 100.950 295.050 103.050 ;
        RECT 301.950 100.950 304.050 103.050 ;
        RECT 293.400 100.050 294.450 100.950 ;
        RECT 292.950 97.950 295.050 100.050 ;
        RECT 298.950 97.950 301.050 100.050 ;
        RECT 286.950 94.950 289.050 97.050 ;
        RECT 290.250 95.250 292.050 96.150 ;
        RECT 292.950 95.850 295.050 96.750 ;
        RECT 295.950 95.250 298.050 96.150 ;
        RECT 299.400 94.050 300.450 97.950 ;
        RECT 283.950 91.950 286.050 94.050 ;
        RECT 286.950 92.850 288.750 93.750 ;
        RECT 289.950 91.950 292.050 94.050 ;
        RECT 295.950 93.450 298.050 94.050 ;
        RECT 298.950 93.450 301.050 94.050 ;
        RECT 295.950 92.400 301.050 93.450 ;
        RECT 295.950 91.950 298.050 92.400 ;
        RECT 298.950 91.950 301.050 92.400 ;
        RECT 302.400 91.050 303.450 100.950 ;
        RECT 317.400 94.050 318.450 106.950 ;
        RECT 325.950 103.950 328.050 106.050 ;
        RECT 326.400 97.050 327.450 103.950 ;
        RECT 338.400 103.050 339.450 130.950 ;
        RECT 344.400 127.050 345.450 160.950 ;
        RECT 347.400 130.050 348.450 163.950 ;
        RECT 353.400 133.050 354.450 181.950 ;
        RECT 355.950 172.950 358.050 175.050 ;
        RECT 356.400 151.050 357.450 172.950 ;
        RECT 355.950 148.950 358.050 151.050 ;
        RECT 349.950 130.950 352.050 133.050 ;
        RECT 352.950 130.950 355.050 133.050 ;
        RECT 350.400 130.050 351.450 130.950 ;
        RECT 346.950 127.950 349.050 130.050 ;
        RECT 349.950 127.950 352.050 130.050 ;
        RECT 355.950 129.450 358.050 130.050 ;
        RECT 359.400 129.450 360.450 193.950 ;
        RECT 365.400 187.050 366.450 193.950 ;
        RECT 364.950 184.950 367.050 187.050 ;
        RECT 368.400 178.050 369.450 193.950 ;
        RECT 380.400 193.050 381.450 193.950 ;
        RECT 383.400 193.050 384.450 196.950 ;
        RECT 410.400 196.050 411.450 230.400 ;
        RECT 412.950 226.950 415.050 229.050 ;
        RECT 413.400 205.050 414.450 226.950 ;
        RECT 416.400 205.050 417.450 232.950 ;
        RECT 418.950 223.950 421.050 226.050 ;
        RECT 419.400 211.050 420.450 223.950 ;
        RECT 421.950 220.950 424.050 223.050 ;
        RECT 422.400 211.050 423.450 220.950 ;
        RECT 418.950 208.950 421.050 211.050 ;
        RECT 421.950 208.950 424.050 211.050 ;
        RECT 421.950 205.950 424.050 208.050 ;
        RECT 430.950 205.950 433.050 208.050 ;
        RECT 412.950 202.950 415.050 205.050 ;
        RECT 415.950 202.950 418.050 205.050 ;
        RECT 416.400 199.050 417.450 202.950 ;
        RECT 412.950 197.250 415.050 198.150 ;
        RECT 415.950 196.950 418.050 199.050 ;
        RECT 418.950 197.250 421.050 198.150 ;
        RECT 385.950 193.950 388.050 196.050 ;
        RECT 389.250 194.250 390.750 195.150 ;
        RECT 391.950 193.950 394.050 196.050 ;
        RECT 397.950 193.950 400.050 196.050 ;
        RECT 401.250 194.850 403.050 195.750 ;
        RECT 403.950 194.250 406.050 195.150 ;
        RECT 406.950 194.850 409.050 195.750 ;
        RECT 409.950 193.950 412.050 196.050 ;
        RECT 412.950 193.950 415.050 196.050 ;
        RECT 416.250 194.250 417.750 195.150 ;
        RECT 418.950 193.950 421.050 196.050 ;
        RECT 376.950 190.950 379.050 193.050 ;
        RECT 379.950 190.950 382.050 193.050 ;
        RECT 382.950 190.950 385.050 193.050 ;
        RECT 388.950 190.950 391.050 193.050 ;
        RECT 403.950 190.950 406.050 193.050 ;
        RECT 409.950 192.450 412.050 193.050 ;
        RECT 413.400 192.450 414.450 193.950 ;
        RECT 409.950 191.400 414.450 192.450 ;
        RECT 415.950 192.450 418.050 193.050 ;
        RECT 418.950 192.450 421.050 193.050 ;
        RECT 415.950 191.400 421.050 192.450 ;
        RECT 409.950 190.950 412.050 191.400 ;
        RECT 415.950 190.950 418.050 191.400 ;
        RECT 418.950 190.950 421.050 191.400 ;
        RECT 367.950 175.950 370.050 178.050 ;
        RECT 361.950 172.950 364.050 175.050 ;
        RECT 362.400 169.050 363.450 172.950 ;
        RECT 370.950 169.950 373.050 172.050 ;
        RECT 371.400 169.050 372.450 169.950 ;
        RECT 377.400 169.050 378.450 190.950 ;
        RECT 380.400 184.050 381.450 190.950 ;
        RECT 379.950 181.950 382.050 184.050 ;
        RECT 389.400 177.450 390.450 190.950 ;
        RECT 394.950 184.950 397.050 187.050 ;
        RECT 386.400 176.400 390.450 177.450 ;
        RECT 386.400 175.050 387.450 176.400 ;
        RECT 385.950 172.950 388.050 175.050 ;
        RECT 388.950 172.950 391.050 175.050 ;
        RECT 391.950 172.950 394.050 175.050 ;
        RECT 389.400 169.050 390.450 172.950 ;
        RECT 392.400 169.050 393.450 172.950 ;
        RECT 361.950 166.950 364.050 169.050 ;
        RECT 364.950 166.950 367.050 169.050 ;
        RECT 368.250 167.250 369.750 168.150 ;
        RECT 370.950 166.950 373.050 169.050 ;
        RECT 376.950 168.450 379.050 169.050 ;
        RECT 374.400 167.400 379.050 168.450 ;
        RECT 361.950 163.950 364.050 166.050 ;
        RECT 365.250 164.850 366.750 165.750 ;
        RECT 367.950 163.950 370.050 166.050 ;
        RECT 371.250 164.850 373.050 165.750 ;
        RECT 361.950 161.850 364.050 162.750 ;
        RECT 361.950 154.950 364.050 157.050 ;
        RECT 362.400 148.050 363.450 154.950 ;
        RECT 361.950 145.950 364.050 148.050 ;
        RECT 368.400 139.050 369.450 163.950 ;
        RECT 370.950 160.950 373.050 163.050 ;
        RECT 371.400 151.050 372.450 160.950 ;
        RECT 374.400 160.050 375.450 167.400 ;
        RECT 376.950 166.950 379.050 167.400 ;
        RECT 380.250 167.250 381.750 168.150 ;
        RECT 382.950 166.950 385.050 169.050 ;
        RECT 386.250 167.250 387.750 168.150 ;
        RECT 388.950 166.950 391.050 169.050 ;
        RECT 391.950 166.950 394.050 169.050 ;
        RECT 376.950 164.850 378.750 165.750 ;
        RECT 379.950 163.950 382.050 166.050 ;
        RECT 383.250 164.850 384.750 165.750 ;
        RECT 385.950 163.950 388.050 166.050 ;
        RECT 389.250 164.850 391.050 165.750 ;
        RECT 391.950 164.850 394.050 165.750 ;
        RECT 380.400 163.050 381.450 163.950 ;
        RECT 376.950 160.950 379.050 163.050 ;
        RECT 379.950 160.950 382.050 163.050 ;
        RECT 373.950 157.950 376.050 160.050 ;
        RECT 370.950 148.950 373.050 151.050 ;
        RECT 367.950 136.950 370.050 139.050 ;
        RECT 377.400 136.050 378.450 160.950 ;
        RECT 386.400 160.050 387.450 163.950 ;
        RECT 385.950 157.950 388.050 160.050 ;
        RECT 382.950 145.950 385.050 148.050 ;
        RECT 379.950 142.950 382.050 145.050 ;
        RECT 376.950 133.950 379.050 136.050 ;
        RECT 380.400 130.050 381.450 142.950 ;
        RECT 364.950 129.450 367.050 130.050 ;
        RECT 353.250 128.250 354.750 129.150 ;
        RECT 355.950 128.400 360.450 129.450 ;
        RECT 355.950 127.950 358.050 128.400 ;
        RECT 340.950 125.250 343.050 126.150 ;
        RECT 343.950 124.950 346.050 127.050 ;
        RECT 346.950 125.250 349.050 126.150 ;
        RECT 349.950 125.850 351.750 126.750 ;
        RECT 352.950 124.950 355.050 127.050 ;
        RECT 356.250 125.850 358.050 126.750 ;
        RECT 340.950 121.950 343.050 124.050 ;
        RECT 344.250 122.250 345.750 123.150 ;
        RECT 346.950 121.950 349.050 124.050 ;
        RECT 341.400 118.050 342.450 121.950 ;
        RECT 343.950 118.950 346.050 121.050 ;
        RECT 340.950 115.950 343.050 118.050 ;
        RECT 344.400 106.050 345.450 118.950 ;
        RECT 343.950 103.950 346.050 106.050 ;
        RECT 346.950 103.950 349.050 106.050 ;
        RECT 337.950 100.950 340.050 103.050 ;
        RECT 337.950 97.950 340.050 100.050 ;
        RECT 319.950 94.950 322.050 97.050 ;
        RECT 323.250 95.250 324.750 96.150 ;
        RECT 325.950 94.950 328.050 97.050 ;
        RECT 331.950 96.450 334.050 97.050 ;
        RECT 329.400 95.400 334.050 96.450 ;
        RECT 304.950 91.950 307.050 94.050 ;
        RECT 308.250 92.250 310.050 93.150 ;
        RECT 316.950 91.950 319.050 94.050 ;
        RECT 320.250 92.850 321.750 93.750 ;
        RECT 322.950 91.950 325.050 94.050 ;
        RECT 326.250 92.850 328.050 93.750 ;
        RECT 323.400 91.050 324.450 91.950 ;
        RECT 286.950 88.950 289.050 91.050 ;
        RECT 298.950 89.850 300.750 90.750 ;
        RECT 301.950 88.950 304.050 91.050 ;
        RECT 305.250 89.850 306.750 90.750 ;
        RECT 307.950 88.950 310.050 91.050 ;
        RECT 316.950 89.850 319.050 90.750 ;
        RECT 319.950 88.950 322.050 91.050 ;
        RECT 322.950 88.950 325.050 91.050 ;
        RECT 287.400 58.050 288.450 88.950 ;
        RECT 298.950 85.950 301.050 88.050 ;
        RECT 301.950 86.850 304.050 87.750 ;
        RECT 292.950 59.250 295.050 60.150 ;
        RECT 259.950 55.950 262.050 58.050 ;
        RECT 263.250 56.250 264.750 57.150 ;
        RECT 265.950 55.950 268.050 58.050 ;
        RECT 268.950 55.950 271.050 58.050 ;
        RECT 280.950 55.950 283.050 58.050 ;
        RECT 286.950 55.950 289.050 58.050 ;
        RECT 290.250 56.250 291.750 57.150 ;
        RECT 292.950 55.950 295.050 58.050 ;
        RECT 296.250 56.250 298.050 57.150 ;
        RECT 259.950 53.850 261.750 54.750 ;
        RECT 262.950 52.950 265.050 55.050 ;
        RECT 266.250 53.850 268.050 54.750 ;
        RECT 253.950 40.950 256.050 43.050 ;
        RECT 250.950 37.950 253.050 40.050 ;
        RECT 251.400 28.050 252.450 37.950 ;
        RECT 263.400 34.050 264.450 52.950 ;
        RECT 269.400 51.450 270.450 55.950 ;
        RECT 271.950 53.250 274.050 54.150 ;
        RECT 277.950 53.250 280.050 54.150 ;
        RECT 286.950 53.850 288.750 54.750 ;
        RECT 289.950 52.950 292.050 55.050 ;
        RECT 295.950 52.950 298.050 55.050 ;
        RECT 299.400 52.050 300.450 85.950 ;
        RECT 308.400 73.050 309.450 88.950 ;
        RECT 307.950 70.950 310.050 73.050 ;
        RECT 316.950 70.950 319.050 73.050 ;
        RECT 304.950 67.950 307.050 70.050 ;
        RECT 305.400 58.050 306.450 67.950 ;
        RECT 301.950 56.250 304.050 57.150 ;
        RECT 304.950 55.950 307.050 58.050 ;
        RECT 313.950 55.950 316.050 58.050 ;
        RECT 301.950 52.950 304.050 55.050 ;
        RECT 305.250 53.250 306.750 54.150 ;
        RECT 307.950 52.950 310.050 55.050 ;
        RECT 311.250 53.250 313.050 54.150 ;
        RECT 271.950 51.450 274.050 52.050 ;
        RECT 269.400 50.400 274.050 51.450 ;
        RECT 271.950 49.950 274.050 50.400 ;
        RECT 275.250 50.250 276.750 51.150 ;
        RECT 277.950 49.950 280.050 52.050 ;
        RECT 298.950 49.950 301.050 52.050 ;
        RECT 274.950 46.950 277.050 49.050 ;
        RECT 275.400 37.050 276.450 46.950 ;
        RECT 277.950 40.950 280.050 43.050 ;
        RECT 286.950 40.950 289.050 43.050 ;
        RECT 302.400 42.450 303.450 52.950 ;
        RECT 304.950 49.950 307.050 52.050 ;
        RECT 308.250 50.850 309.750 51.750 ;
        RECT 310.950 51.450 313.050 52.050 ;
        RECT 314.400 51.450 315.450 55.950 ;
        RECT 317.400 55.050 318.450 70.950 ;
        RECT 320.400 55.050 321.450 88.950 ;
        RECT 329.400 88.050 330.450 95.400 ;
        RECT 331.950 94.950 334.050 95.400 ;
        RECT 335.250 95.250 337.050 96.150 ;
        RECT 337.950 95.850 340.050 96.750 ;
        RECT 340.950 95.250 343.050 96.150 ;
        RECT 343.950 94.950 346.050 97.050 ;
        RECT 344.400 94.050 345.450 94.950 ;
        RECT 331.950 92.850 333.750 93.750 ;
        RECT 334.950 91.950 337.050 94.050 ;
        RECT 340.950 93.450 343.050 94.050 ;
        RECT 343.950 93.450 346.050 94.050 ;
        RECT 340.950 92.400 346.050 93.450 ;
        RECT 340.950 91.950 343.050 92.400 ;
        RECT 343.950 91.950 346.050 92.400 ;
        RECT 347.400 91.050 348.450 103.950 ;
        RECT 355.950 100.950 358.050 103.050 ;
        RECT 349.950 94.950 352.050 97.050 ;
        RECT 356.400 94.050 357.450 100.950 ;
        RECT 359.400 97.050 360.450 128.400 ;
        RECT 362.400 128.400 367.050 129.450 ;
        RECT 362.400 118.050 363.450 128.400 ;
        RECT 364.950 127.950 367.050 128.400 ;
        RECT 368.250 128.250 369.750 129.150 ;
        RECT 370.950 127.950 373.050 130.050 ;
        RECT 373.950 127.950 376.050 130.050 ;
        RECT 377.250 128.250 378.750 129.150 ;
        RECT 379.950 127.950 382.050 130.050 ;
        RECT 364.950 125.850 366.750 126.750 ;
        RECT 367.950 124.950 370.050 127.050 ;
        RECT 371.250 125.850 373.050 126.750 ;
        RECT 373.950 125.850 375.750 126.750 ;
        RECT 376.950 124.950 379.050 127.050 ;
        RECT 380.250 125.850 382.050 126.750 ;
        RECT 361.950 115.950 364.050 118.050 ;
        RECT 368.400 100.050 369.450 124.950 ;
        RECT 377.400 121.050 378.450 124.950 ;
        RECT 376.950 118.950 379.050 121.050 ;
        RECT 383.400 112.050 384.450 145.950 ;
        RECT 386.400 124.050 387.450 157.950 ;
        RECT 395.400 154.050 396.450 184.950 ;
        RECT 400.950 178.950 403.050 181.050 ;
        RECT 401.400 169.050 402.450 178.950 ;
        RECT 404.400 178.050 405.450 190.950 ;
        RECT 403.950 175.950 406.050 178.050 ;
        RECT 400.950 166.950 403.050 169.050 ;
        RECT 397.950 164.250 400.050 165.150 ;
        RECT 400.950 164.850 403.050 165.750 ;
        RECT 397.950 160.950 400.050 163.050 ;
        RECT 397.950 154.950 400.050 157.050 ;
        RECT 394.950 151.950 397.050 154.050 ;
        RECT 398.400 142.050 399.450 154.950 ;
        RECT 404.400 148.050 405.450 175.950 ;
        RECT 403.950 145.950 406.050 148.050 ;
        RECT 410.400 145.050 411.450 190.950 ;
        RECT 415.950 172.950 418.050 175.050 ;
        RECT 416.400 172.050 417.450 172.950 ;
        RECT 415.950 169.950 418.050 172.050 ;
        RECT 422.400 171.450 423.450 205.950 ;
        RECT 424.950 199.950 427.050 202.050 ;
        RECT 425.400 196.050 426.450 199.950 ;
        RECT 427.950 197.250 430.050 198.150 ;
        RECT 424.950 193.950 427.050 196.050 ;
        RECT 427.950 193.950 430.050 196.050 ;
        RECT 424.950 187.950 427.050 190.050 ;
        RECT 425.400 172.050 426.450 187.950 ;
        RECT 428.400 178.050 429.450 193.950 ;
        RECT 431.400 190.050 432.450 205.950 ;
        RECT 434.400 202.050 435.450 295.950 ;
        RECT 437.400 295.050 438.450 299.400 ;
        RECT 436.950 292.950 439.050 295.050 ;
        RECT 440.400 289.050 441.450 304.950 ;
        RECT 445.950 289.950 448.050 292.050 ;
        RECT 439.950 286.950 442.050 289.050 ;
        RECT 442.950 274.950 445.050 277.050 ;
        RECT 443.400 274.050 444.450 274.950 ;
        RECT 436.950 271.950 439.050 274.050 ;
        RECT 442.950 271.950 445.050 274.050 ;
        RECT 437.400 259.050 438.450 271.950 ;
        RECT 439.950 269.250 442.050 270.150 ;
        RECT 442.950 269.850 445.050 270.750 ;
        RECT 439.950 265.950 442.050 268.050 ;
        RECT 440.400 262.050 441.450 265.950 ;
        RECT 439.950 259.950 442.050 262.050 ;
        RECT 436.950 256.950 439.050 259.050 ;
        RECT 436.950 253.950 439.050 256.050 ;
        RECT 437.400 208.050 438.450 253.950 ;
        RECT 446.400 250.050 447.450 289.950 ;
        RECT 449.400 289.050 450.450 314.400 ;
        RECT 461.400 313.050 462.450 322.950 ;
        RECT 467.400 316.050 468.450 337.950 ;
        RECT 466.950 313.950 469.050 316.050 ;
        RECT 473.400 313.050 474.450 337.950 ;
        RECT 476.400 334.050 477.450 337.950 ;
        RECT 475.950 331.950 478.050 334.050 ;
        RECT 479.400 330.450 480.450 337.950 ;
        RECT 481.950 334.950 484.050 337.050 ;
        RECT 482.400 334.050 483.450 334.950 ;
        RECT 481.950 331.950 484.050 334.050 ;
        RECT 485.400 330.450 486.450 337.950 ;
        RECT 488.400 333.450 489.450 349.950 ;
        RECT 491.400 336.450 492.450 373.950 ;
        RECT 494.400 367.050 495.450 377.400 ;
        RECT 493.950 364.950 496.050 367.050 ;
        RECT 497.400 363.450 498.450 401.400 ;
        RECT 506.400 394.050 507.450 406.950 ;
        RECT 502.950 391.950 505.050 394.050 ;
        RECT 505.950 391.950 508.050 394.050 ;
        RECT 503.400 388.050 504.450 391.950 ;
        RECT 505.950 388.950 508.050 391.050 ;
        RECT 499.950 385.950 502.050 388.050 ;
        RECT 502.950 385.950 505.050 388.050 ;
        RECT 499.950 383.850 502.050 384.750 ;
        RECT 502.950 383.250 505.050 384.150 ;
        RECT 502.950 379.950 505.050 382.050 ;
        RECT 499.950 376.950 502.050 379.050 ;
        RECT 494.400 362.400 498.450 363.450 ;
        RECT 494.400 340.050 495.450 362.400 ;
        RECT 496.950 358.950 499.050 361.050 ;
        RECT 497.400 346.050 498.450 358.950 ;
        RECT 500.400 349.050 501.450 376.950 ;
        RECT 503.400 358.050 504.450 379.950 ;
        RECT 506.400 376.050 507.450 388.950 ;
        RECT 509.400 388.050 510.450 412.950 ;
        RECT 511.950 409.800 514.050 412.050 ;
        RECT 512.400 403.050 513.450 409.800 ;
        RECT 515.400 406.050 516.450 457.950 ;
        RECT 518.400 448.050 519.450 460.950 ;
        RECT 529.950 454.950 532.050 457.050 ;
        RECT 530.400 454.050 531.450 454.950 ;
        RECT 520.950 452.250 522.750 453.150 ;
        RECT 523.950 451.950 526.050 454.050 ;
        RECT 529.950 451.950 532.050 454.050 ;
        RECT 520.950 448.950 523.050 451.050 ;
        RECT 524.250 449.850 525.750 450.750 ;
        RECT 526.950 448.950 529.050 451.050 ;
        RECT 530.250 449.850 532.050 450.750 ;
        RECT 517.950 445.950 520.050 448.050 ;
        RECT 526.950 446.850 529.050 447.750 ;
        RECT 520.950 436.950 523.050 439.050 ;
        RECT 517.950 415.950 520.050 418.050 ;
        RECT 514.950 403.950 517.050 406.050 ;
        RECT 511.950 400.950 514.050 403.050 ;
        RECT 514.950 400.950 517.050 403.050 ;
        RECT 511.950 394.950 514.050 397.050 ;
        RECT 508.950 385.950 511.050 388.050 ;
        RECT 512.400 385.050 513.450 394.950 ;
        RECT 508.950 382.950 511.050 385.050 ;
        RECT 511.950 382.950 514.050 385.050 ;
        RECT 505.950 373.950 508.050 376.050 ;
        RECT 502.950 355.950 505.050 358.050 ;
        RECT 499.950 346.950 502.050 349.050 ;
        RECT 502.950 347.250 505.050 348.150 ;
        RECT 496.950 343.950 499.050 346.050 ;
        RECT 500.250 344.250 501.750 345.150 ;
        RECT 502.950 343.950 505.050 346.050 ;
        RECT 506.250 344.250 508.050 345.150 ;
        RECT 496.950 341.850 498.750 342.750 ;
        RECT 499.950 340.950 502.050 343.050 ;
        RECT 505.950 340.950 508.050 343.050 ;
        RECT 493.950 337.950 496.050 340.050 ;
        RECT 499.950 337.950 502.050 340.050 ;
        RECT 491.400 335.400 495.450 336.450 ;
        RECT 488.400 332.400 492.450 333.450 ;
        RECT 476.400 329.400 480.450 330.450 ;
        RECT 482.400 329.400 486.450 330.450 ;
        RECT 476.400 325.050 477.450 329.400 ;
        RECT 482.400 327.450 483.450 329.400 ;
        RECT 479.400 326.400 483.450 327.450 ;
        RECT 475.950 322.950 478.050 325.050 ;
        RECT 460.950 310.950 463.050 313.050 ;
        RECT 464.400 311.400 471.450 312.450 ;
        RECT 464.400 310.050 465.450 311.400 ;
        RECT 470.400 310.050 471.450 311.400 ;
        RECT 472.950 310.950 475.050 313.050 ;
        RECT 451.950 307.950 454.050 310.050 ;
        RECT 457.950 307.950 460.050 310.050 ;
        RECT 461.250 308.250 463.050 309.150 ;
        RECT 463.950 307.950 466.050 310.050 ;
        RECT 466.950 308.250 468.750 309.150 ;
        RECT 469.950 307.950 472.050 310.050 ;
        RECT 473.250 308.250 475.050 309.150 ;
        RECT 451.950 305.850 453.750 306.750 ;
        RECT 454.950 304.950 457.050 307.050 ;
        RECT 458.250 305.850 459.750 306.750 ;
        RECT 460.950 304.950 463.050 307.050 ;
        RECT 466.950 304.950 469.050 307.050 ;
        RECT 470.250 305.850 471.750 306.750 ;
        RECT 472.950 304.950 475.050 307.050 ;
        RECT 454.950 302.850 457.050 303.750 ;
        RECT 448.950 286.950 451.050 289.050 ;
        RECT 451.950 286.950 454.050 289.050 ;
        RECT 452.400 274.050 453.450 286.950 ;
        RECT 461.400 283.050 462.450 304.950 ;
        RECT 463.950 301.950 466.050 304.050 ;
        RECT 466.950 301.950 469.050 304.050 ;
        RECT 460.950 280.950 463.050 283.050 ;
        RECT 454.950 277.950 457.050 280.050 ;
        RECT 451.950 271.950 454.050 274.050 ;
        RECT 448.950 269.250 451.050 270.150 ;
        RECT 451.950 269.250 454.050 270.150 ;
        RECT 448.950 265.950 451.050 268.050 ;
        RECT 451.950 265.950 454.050 268.050 ;
        RECT 448.950 262.950 451.050 265.050 ;
        RECT 445.950 247.950 448.050 250.050 ;
        RECT 439.950 244.950 442.050 247.050 ;
        RECT 440.400 238.050 441.450 244.950 ;
        RECT 442.950 241.950 445.050 244.050 ;
        RECT 449.400 243.450 450.450 262.950 ;
        RECT 452.400 253.050 453.450 265.950 ;
        RECT 455.400 265.050 456.450 277.950 ;
        RECT 457.950 274.950 460.050 277.050 ;
        RECT 458.400 274.050 459.450 274.950 ;
        RECT 457.950 271.950 460.050 274.050 ;
        RECT 464.400 271.050 465.450 301.950 ;
        RECT 467.400 280.050 468.450 301.950 ;
        RECT 469.950 292.950 472.050 295.050 ;
        RECT 466.950 277.950 469.050 280.050 ;
        RECT 467.400 277.050 468.450 277.950 ;
        RECT 466.950 274.950 469.050 277.050 ;
        RECT 457.950 269.850 460.050 270.750 ;
        RECT 460.950 269.250 463.050 270.150 ;
        RECT 463.950 268.950 466.050 271.050 ;
        RECT 460.950 265.950 463.050 268.050 ;
        RECT 461.400 265.050 462.450 265.950 ;
        RECT 464.400 265.050 465.450 268.950 ;
        RECT 454.950 262.950 457.050 265.050 ;
        RECT 460.950 262.950 463.050 265.050 ;
        RECT 463.950 262.950 466.050 265.050 ;
        RECT 467.400 259.050 468.450 274.950 ;
        RECT 454.950 256.950 457.050 259.050 ;
        RECT 466.950 256.950 469.050 259.050 ;
        RECT 451.950 250.950 454.050 253.050 ;
        RECT 449.400 242.400 453.450 243.450 ;
        RECT 443.400 241.050 444.450 241.950 ;
        RECT 442.950 238.950 445.050 241.050 ;
        RECT 446.250 239.250 447.750 240.150 ;
        RECT 448.950 238.950 451.050 241.050 ;
        RECT 452.400 238.050 453.450 242.400 ;
        RECT 439.950 235.950 442.050 238.050 ;
        RECT 443.250 236.850 444.750 237.750 ;
        RECT 445.950 235.950 448.050 238.050 ;
        RECT 449.250 236.850 451.050 237.750 ;
        RECT 451.950 235.950 454.050 238.050 ;
        RECT 439.950 233.850 442.050 234.750 ;
        RECT 442.950 214.950 445.050 217.050 ;
        RECT 436.950 205.950 439.050 208.050 ;
        RECT 433.950 199.950 436.050 202.050 ;
        RECT 436.950 199.950 439.050 202.050 ;
        RECT 433.950 197.250 436.050 198.150 ;
        RECT 433.950 193.950 436.050 196.050 ;
        RECT 430.950 187.950 433.050 190.050 ;
        RECT 430.950 181.950 433.050 184.050 ;
        RECT 427.950 175.950 430.050 178.050 ;
        RECT 428.400 175.050 429.450 175.950 ;
        RECT 427.950 172.950 430.050 175.050 ;
        RECT 419.400 170.400 423.450 171.450 ;
        RECT 412.950 167.250 415.050 168.150 ;
        RECT 415.950 167.850 418.050 168.750 ;
        RECT 412.950 163.950 415.050 166.050 ;
        RECT 419.400 162.450 420.450 170.400 ;
        RECT 424.950 169.950 427.050 172.050 ;
        RECT 427.950 169.950 430.050 172.050 ;
        RECT 428.400 169.050 429.450 169.950 ;
        RECT 431.400 169.050 432.450 181.950 ;
        RECT 437.400 174.450 438.450 199.950 ;
        RECT 443.400 199.050 444.450 214.950 ;
        RECT 446.400 202.050 447.450 235.950 ;
        RECT 451.950 229.950 454.050 232.050 ;
        RECT 445.950 199.950 448.050 202.050 ;
        RECT 448.950 200.250 451.050 201.150 ;
        RECT 439.950 197.250 441.750 198.150 ;
        RECT 442.950 196.950 445.050 199.050 ;
        RECT 446.250 197.250 447.750 198.150 ;
        RECT 448.950 196.950 451.050 199.050 ;
        RECT 439.950 193.950 442.050 196.050 ;
        RECT 443.250 194.850 444.750 195.750 ;
        RECT 445.950 193.950 448.050 196.050 ;
        RECT 452.400 195.450 453.450 229.950 ;
        RECT 455.400 220.050 456.450 256.950 ;
        RECT 466.950 250.950 469.050 253.050 ;
        RECT 460.950 241.950 463.050 244.050 ;
        RECT 461.400 238.050 462.450 241.950 ;
        RECT 467.400 238.050 468.450 250.950 ;
        RECT 470.400 241.050 471.450 292.950 ;
        RECT 473.400 274.050 474.450 304.950 ;
        RECT 476.400 295.050 477.450 322.950 ;
        RECT 479.400 316.050 480.450 326.400 ;
        RECT 484.950 325.950 487.050 328.050 ;
        RECT 481.950 316.950 484.050 319.050 ;
        RECT 478.950 313.950 481.050 316.050 ;
        RECT 482.400 312.450 483.450 316.950 ;
        RECT 485.400 313.050 486.450 325.950 ;
        RECT 479.400 311.400 483.450 312.450 ;
        RECT 479.400 310.050 480.450 311.400 ;
        RECT 484.950 310.950 487.050 313.050 ;
        RECT 478.950 307.950 481.050 310.050 ;
        RECT 481.950 307.950 484.050 310.050 ;
        RECT 484.950 307.950 487.050 310.050 ;
        RECT 488.250 308.250 490.050 309.150 ;
        RECT 482.400 307.050 483.450 307.950 ;
        RECT 478.950 305.850 480.750 306.750 ;
        RECT 481.950 304.950 484.050 307.050 ;
        RECT 485.250 305.850 486.750 306.750 ;
        RECT 487.950 304.950 490.050 307.050 ;
        RECT 478.950 301.950 481.050 304.050 ;
        RECT 481.950 302.850 484.050 303.750 ;
        RECT 487.950 301.950 490.050 304.050 ;
        RECT 479.400 301.050 480.450 301.950 ;
        RECT 478.950 298.950 481.050 301.050 ;
        RECT 475.950 292.950 478.050 295.050 ;
        RECT 475.950 286.950 478.050 289.050 ;
        RECT 472.950 271.950 475.050 274.050 ;
        RECT 476.400 271.050 477.450 286.950 ;
        RECT 479.400 277.050 480.450 298.950 ;
        RECT 488.400 283.050 489.450 301.950 ;
        RECT 491.400 283.050 492.450 332.400 ;
        RECT 494.400 325.050 495.450 335.400 ;
        RECT 496.950 334.950 499.050 337.050 ;
        RECT 497.400 331.050 498.450 334.950 ;
        RECT 496.950 328.950 499.050 331.050 ;
        RECT 493.950 322.950 496.050 325.050 ;
        RECT 500.400 318.450 501.450 337.950 ;
        RECT 502.950 331.950 505.050 334.050 ;
        RECT 503.400 328.050 504.450 331.950 ;
        RECT 506.400 331.050 507.450 340.950 ;
        RECT 505.950 328.950 508.050 331.050 ;
        RECT 502.950 325.950 505.050 328.050 ;
        RECT 500.400 317.400 504.450 318.450 ;
        RECT 503.400 316.050 504.450 317.400 ;
        RECT 499.950 313.950 502.050 316.050 ;
        RECT 502.950 313.950 505.050 316.050 ;
        RECT 500.400 310.050 501.450 313.950 ;
        RECT 505.950 310.950 508.050 313.050 ;
        RECT 493.950 307.950 496.050 310.050 ;
        RECT 496.950 308.250 498.750 309.150 ;
        RECT 499.950 307.950 502.050 310.050 ;
        RECT 503.250 308.250 505.050 309.150 ;
        RECT 505.950 308.850 508.050 309.750 ;
        RECT 494.400 303.450 495.450 307.950 ;
        RECT 496.950 304.950 499.050 307.050 ;
        RECT 500.250 305.850 501.750 306.750 ;
        RECT 502.950 304.950 505.050 307.050 ;
        RECT 505.950 304.950 508.050 307.050 ;
        RECT 503.400 304.050 504.450 304.950 ;
        RECT 494.400 302.400 498.450 303.450 ;
        RECT 487.950 280.950 490.050 283.050 ;
        RECT 490.950 280.950 493.050 283.050 ;
        RECT 478.950 274.950 481.050 277.050 ;
        RECT 481.950 274.950 484.050 277.050 ;
        RECT 493.950 274.950 496.050 277.050 ;
        RECT 482.400 271.050 483.450 274.950 ;
        RECT 494.400 274.050 495.450 274.950 ;
        RECT 493.950 271.950 496.050 274.050 ;
        RECT 472.950 269.250 474.750 270.150 ;
        RECT 475.950 268.950 478.050 271.050 ;
        RECT 479.250 269.250 480.750 270.150 ;
        RECT 481.950 268.950 484.050 271.050 ;
        RECT 485.250 269.250 487.050 270.150 ;
        RECT 487.950 268.950 490.050 271.050 ;
        RECT 490.950 269.250 493.050 270.150 ;
        RECT 493.950 269.850 496.050 270.750 ;
        RECT 472.950 265.950 475.050 268.050 ;
        RECT 476.250 266.850 477.750 267.750 ;
        RECT 478.950 265.950 481.050 268.050 ;
        RECT 482.250 266.850 483.750 267.750 ;
        RECT 484.950 265.950 487.050 268.050 ;
        RECT 473.400 265.050 474.450 265.950 ;
        RECT 472.950 262.950 475.050 265.050 ;
        RECT 475.950 259.950 478.050 262.050 ;
        RECT 472.950 250.950 475.050 253.050 ;
        RECT 469.950 238.950 472.050 241.050 ;
        RECT 473.400 238.050 474.450 250.950 ;
        RECT 476.400 240.450 477.450 259.950 ;
        RECT 479.400 244.050 480.450 265.950 ;
        RECT 488.400 265.050 489.450 268.950 ;
        RECT 490.950 265.950 493.050 268.050 ;
        RECT 484.950 262.950 487.050 265.050 ;
        RECT 487.950 262.950 490.050 265.050 ;
        RECT 485.400 262.050 486.450 262.950 ;
        RECT 484.950 259.950 487.050 262.050 ;
        RECT 481.950 247.950 484.050 250.050 ;
        RECT 478.950 241.950 481.050 244.050 ;
        RECT 476.400 239.400 480.450 240.450 ;
        RECT 457.950 236.250 459.750 237.150 ;
        RECT 460.950 235.950 463.050 238.050 ;
        RECT 466.950 235.950 469.050 238.050 ;
        RECT 469.950 236.250 471.750 237.150 ;
        RECT 472.950 235.950 475.050 238.050 ;
        RECT 476.250 236.250 478.050 237.150 ;
        RECT 457.950 232.950 460.050 235.050 ;
        RECT 461.250 233.850 462.750 234.750 ;
        RECT 463.950 232.950 466.050 235.050 ;
        RECT 467.250 233.850 469.050 234.750 ;
        RECT 469.950 232.950 472.050 235.050 ;
        RECT 473.250 233.850 474.750 234.750 ;
        RECT 475.950 232.950 478.050 235.050 ;
        RECT 454.950 217.950 457.050 220.050 ;
        RECT 455.400 204.450 456.450 217.950 ;
        RECT 458.400 214.050 459.450 232.950 ;
        RECT 463.950 230.850 466.050 231.750 ;
        RECT 457.950 211.950 460.050 214.050 ;
        RECT 470.400 208.050 471.450 232.950 ;
        RECT 476.400 232.050 477.450 232.950 ;
        RECT 475.950 229.950 478.050 232.050 ;
        RECT 479.400 220.050 480.450 239.400 ;
        RECT 482.400 232.050 483.450 247.950 ;
        RECT 485.400 238.050 486.450 259.950 ;
        RECT 487.950 256.950 490.050 259.050 ;
        RECT 488.400 241.050 489.450 256.950 ;
        RECT 491.400 250.050 492.450 265.950 ;
        RECT 497.400 259.050 498.450 302.400 ;
        RECT 502.950 301.950 505.050 304.050 ;
        RECT 499.950 277.950 502.050 280.050 ;
        RECT 500.400 274.050 501.450 277.950 ;
        RECT 506.400 276.450 507.450 304.950 ;
        RECT 509.400 298.050 510.450 382.950 ;
        RECT 511.950 380.850 514.050 381.750 ;
        RECT 515.400 379.050 516.450 400.950 ;
        RECT 518.400 385.050 519.450 415.950 ;
        RECT 521.400 411.450 522.450 436.950 ;
        RECT 533.400 418.050 534.450 460.950 ;
        RECT 542.400 460.050 543.450 469.950 ;
        RECT 545.400 460.050 546.450 482.400 ;
        RECT 550.950 481.950 553.050 484.050 ;
        RECT 553.950 481.950 556.050 484.050 ;
        RECT 556.950 481.950 559.050 484.050 ;
        RECT 560.250 482.250 561.750 483.150 ;
        RECT 562.950 481.950 565.050 484.050 ;
        RECT 547.950 463.950 550.050 466.050 ;
        RECT 541.950 457.950 544.050 460.050 ;
        RECT 544.950 457.950 547.050 460.050 ;
        RECT 538.950 455.250 541.050 456.150 ;
        RECT 541.950 455.850 544.050 456.750 ;
        RECT 544.950 454.950 547.050 457.050 ;
        RECT 538.950 451.950 541.050 454.050 ;
        RECT 541.950 451.950 544.050 454.050 ;
        RECT 535.950 448.950 538.050 451.050 ;
        RECT 538.950 448.950 541.050 451.050 ;
        RECT 536.400 445.050 537.450 448.950 ;
        RECT 535.950 442.950 538.050 445.050 ;
        RECT 539.400 430.050 540.450 448.950 ;
        RECT 538.950 427.950 541.050 430.050 ;
        RECT 523.950 416.250 526.050 417.150 ;
        RECT 532.950 415.950 535.050 418.050 ;
        RECT 523.950 412.950 526.050 415.050 ;
        RECT 527.250 413.250 528.750 414.150 ;
        RECT 529.950 412.950 532.050 415.050 ;
        RECT 533.250 413.250 535.050 414.150 ;
        RECT 538.950 412.950 541.050 415.050 ;
        RECT 521.400 410.400 525.450 411.450 ;
        RECT 520.950 397.950 523.050 400.050 ;
        RECT 521.400 385.050 522.450 397.950 ;
        RECT 517.950 382.950 520.050 385.050 ;
        RECT 520.950 382.950 523.050 385.050 ;
        RECT 517.950 380.250 520.050 381.150 ;
        RECT 520.950 380.850 523.050 381.750 ;
        RECT 514.950 376.950 517.050 379.050 ;
        RECT 517.950 376.950 520.050 379.050 ;
        RECT 524.400 367.050 525.450 410.400 ;
        RECT 526.950 409.950 529.050 412.050 ;
        RECT 530.250 410.850 531.750 411.750 ;
        RECT 532.950 409.950 535.050 412.050 ;
        RECT 535.950 410.250 538.050 411.150 ;
        RECT 538.950 410.850 541.050 411.750 ;
        RECT 533.400 399.450 534.450 409.950 ;
        RECT 535.950 406.950 538.050 409.050 ;
        RECT 536.400 403.050 537.450 406.950 ;
        RECT 542.400 403.050 543.450 451.950 ;
        RECT 545.400 448.050 546.450 454.950 ;
        RECT 548.400 453.450 549.450 463.950 ;
        RECT 554.400 463.050 555.450 481.950 ;
        RECT 557.400 481.050 558.450 481.950 ;
        RECT 556.950 478.950 559.050 481.050 ;
        RECT 559.950 478.950 562.050 481.050 ;
        RECT 557.400 478.050 558.450 478.950 ;
        RECT 556.950 475.950 559.050 478.050 ;
        RECT 560.400 474.450 561.450 478.950 ;
        RECT 563.400 475.050 564.450 481.950 ;
        RECT 557.400 473.400 561.450 474.450 ;
        RECT 557.400 469.050 558.450 473.400 ;
        RECT 562.950 472.950 565.050 475.050 ;
        RECT 566.400 472.050 567.450 518.400 ;
        RECT 574.950 517.950 577.050 520.050 ;
        RECT 577.950 519.300 580.050 521.400 ;
        RECT 568.950 514.950 571.050 517.050 ;
        RECT 569.400 508.050 570.450 514.950 ;
        RECT 568.950 505.950 571.050 508.050 ;
        RECT 575.400 493.050 576.450 517.950 ;
        RECT 578.550 515.700 579.750 519.300 ;
        RECT 577.950 513.600 580.050 515.700 ;
        RECT 581.400 504.450 582.450 532.950 ;
        RECT 584.400 531.450 585.450 580.950 ;
        RECT 590.400 562.050 591.450 595.950 ;
        RECT 596.400 583.050 597.450 599.400 ;
        RECT 602.250 593.400 603.450 605.400 ;
        RECT 604.950 602.250 607.050 603.150 ;
        RECT 604.950 598.950 607.050 601.050 ;
        RECT 601.950 591.300 604.050 593.400 ;
        RECT 602.250 587.700 603.450 591.300 ;
        RECT 601.950 585.600 604.050 587.700 ;
        RECT 605.400 586.050 606.450 598.950 ;
        RECT 608.400 591.450 609.450 619.950 ;
        RECT 611.400 595.050 612.450 695.400 ;
        RECT 626.400 691.050 627.450 697.950 ;
        RECT 632.550 693.600 633.750 707.250 ;
        RECT 635.250 693.600 636.450 710.850 ;
        RECT 642.900 710.400 645.000 712.500 ;
        RECT 646.950 710.400 649.050 712.500 ;
        RECT 637.950 707.250 640.050 709.350 ;
        RECT 638.400 693.600 639.600 707.250 ;
        RECT 643.350 701.550 644.550 710.400 ;
        RECT 647.550 704.250 648.750 710.400 ;
        RECT 646.950 702.150 649.050 704.250 ;
        RECT 642.750 699.450 644.850 701.550 ;
        RECT 643.350 693.600 644.550 699.450 ;
        RECT 647.550 693.600 648.750 702.150 ;
        RECT 649.950 698.250 652.050 699.150 ;
        RECT 649.950 694.950 652.050 697.050 ;
        RECT 631.950 691.500 634.050 693.600 ;
        RECT 634.950 691.500 637.050 693.600 ;
        RECT 637.950 691.500 640.050 693.600 ;
        RECT 642.750 691.500 644.850 693.600 ;
        RECT 646.950 691.500 649.050 693.600 ;
        RECT 625.950 688.950 628.050 691.050 ;
        RECT 613.950 671.250 616.050 672.150 ;
        RECT 626.400 670.050 627.450 688.950 ;
        RECT 650.400 684.450 651.450 694.950 ;
        RECT 656.250 694.050 657.450 712.950 ;
        RECT 659.250 708.750 660.450 712.950 ;
        RECT 658.950 706.650 661.050 708.750 ;
        RECT 659.250 694.050 660.450 706.650 ;
        RECT 662.250 694.050 663.450 712.950 ;
        RECT 719.550 709.350 720.750 713.100 ;
        RECT 742.950 712.950 745.050 715.050 ;
        RECT 745.950 712.950 748.050 715.050 ;
        RECT 748.950 712.950 751.050 715.050 ;
        RECT 721.950 710.850 724.050 712.950 ;
        RECT 718.950 707.250 721.050 709.350 ;
        RECT 673.950 705.450 676.050 706.050 ;
        RECT 667.950 704.250 670.050 705.150 ;
        RECT 671.400 704.400 676.050 705.450 ;
        RECT 667.950 697.950 670.050 700.050 ;
        RECT 655.950 691.950 658.050 694.050 ;
        RECT 658.950 691.950 661.050 694.050 ;
        RECT 661.950 691.950 664.050 694.050 ;
        RECT 650.400 683.400 654.450 684.450 ;
        RECT 634.950 677.400 637.050 679.500 ;
        RECT 637.950 677.400 640.050 679.500 ;
        RECT 640.950 677.400 643.050 679.500 ;
        RECT 645.750 677.400 647.850 679.500 ;
        RECT 649.950 677.400 652.050 679.500 ;
        RECT 653.400 679.050 654.450 683.400 ;
        RECT 613.950 667.950 616.050 670.050 ;
        RECT 625.950 667.950 628.050 670.050 ;
        RECT 631.950 667.950 634.050 670.050 ;
        RECT 614.400 622.050 615.450 667.950 ;
        RECT 625.950 665.850 628.050 666.750 ;
        RECT 616.950 638.400 619.050 640.500 ;
        RECT 613.950 619.950 616.050 622.050 ;
        RECT 617.400 621.600 618.600 638.400 ;
        RECT 622.950 629.250 625.050 630.150 ;
        RECT 628.950 629.250 631.050 630.150 ;
        RECT 622.950 625.950 625.050 628.050 ;
        RECT 628.950 627.450 631.050 628.050 ;
        RECT 632.400 627.450 633.450 667.950 ;
        RECT 635.550 663.750 636.750 677.400 ;
        RECT 634.950 661.650 637.050 663.750 ;
        RECT 635.550 657.900 636.750 661.650 ;
        RECT 638.250 660.150 639.450 677.400 ;
        RECT 641.400 663.750 642.600 677.400 ;
        RECT 646.350 671.550 647.550 677.400 ;
        RECT 645.750 669.450 647.850 671.550 ;
        RECT 640.950 661.650 643.050 663.750 ;
        RECT 646.350 660.600 647.550 669.450 ;
        RECT 650.550 668.850 651.750 677.400 ;
        RECT 652.950 676.950 655.050 679.050 ;
        RECT 658.950 676.950 661.050 679.050 ;
        RECT 661.950 676.950 664.050 679.050 ;
        RECT 664.950 676.950 667.050 679.050 ;
        RECT 652.950 675.450 655.050 676.050 ;
        RECT 652.950 674.400 657.450 675.450 ;
        RECT 652.950 673.950 655.050 674.400 ;
        RECT 652.950 671.850 655.050 672.750 ;
        RECT 656.400 670.050 657.450 674.400 ;
        RECT 649.950 666.750 652.050 668.850 ;
        RECT 652.950 667.950 655.050 670.050 ;
        RECT 655.950 667.950 658.050 670.050 ;
        RECT 650.550 660.600 651.750 666.750 ;
        RECT 637.950 658.050 640.050 660.150 ;
        RECT 645.900 658.500 648.000 660.600 ;
        RECT 649.950 658.500 652.050 660.600 ;
        RECT 634.950 655.800 637.050 657.900 ;
        RECT 640.950 655.950 643.050 658.050 ;
        RECT 634.950 646.950 637.050 649.050 ;
        RECT 628.950 626.400 633.450 627.450 ;
        RECT 628.950 625.950 631.050 626.400 ;
        RECT 625.950 622.950 628.050 625.050 ;
        RECT 626.400 622.050 627.450 622.950 ;
        RECT 616.950 619.500 619.050 621.600 ;
        RECT 625.950 619.950 628.050 622.050 ;
        RECT 622.950 610.950 625.050 613.050 ;
        RECT 619.950 604.950 622.050 607.050 ;
        RECT 613.950 599.250 616.050 600.150 ;
        RECT 616.950 599.850 619.050 600.750 ;
        RECT 613.950 595.950 616.050 598.050 ;
        RECT 610.950 592.950 613.050 595.050 ;
        RECT 608.400 590.400 612.450 591.450 ;
        RECT 604.950 583.950 607.050 586.050 ;
        RECT 595.950 580.950 598.050 583.050 ;
        RECT 607.950 568.950 610.050 571.050 ;
        RECT 608.400 568.050 609.450 568.950 ;
        RECT 607.950 565.950 610.050 568.050 ;
        RECT 607.950 562.950 610.050 565.050 ;
        RECT 586.950 560.250 589.050 561.150 ;
        RECT 589.950 559.950 592.050 562.050 ;
        RECT 586.950 556.950 589.050 559.050 ;
        RECT 590.250 557.250 591.750 558.150 ;
        RECT 592.950 556.950 595.050 559.050 ;
        RECT 596.250 557.250 598.050 558.150 ;
        RECT 598.950 557.250 601.050 558.150 ;
        RECT 604.950 557.250 607.050 558.150 ;
        RECT 586.950 553.950 589.050 556.050 ;
        RECT 589.950 553.950 592.050 556.050 ;
        RECT 593.250 554.850 594.750 555.750 ;
        RECT 595.950 555.450 598.050 556.050 ;
        RECT 598.950 555.450 601.050 556.050 ;
        RECT 595.950 554.400 601.050 555.450 ;
        RECT 595.950 553.950 598.050 554.400 ;
        RECT 598.950 553.950 601.050 554.400 ;
        RECT 602.250 554.250 603.750 555.150 ;
        RECT 604.950 553.950 607.050 556.050 ;
        RECT 587.400 535.050 588.450 553.950 ;
        RECT 590.400 547.050 591.450 553.950 ;
        RECT 599.400 553.050 600.450 553.950 ;
        RECT 595.950 550.950 598.050 553.050 ;
        RECT 598.950 550.950 601.050 553.050 ;
        RECT 601.950 550.950 604.050 553.050 ;
        RECT 608.400 552.450 609.450 562.950 ;
        RECT 611.400 559.050 612.450 590.400 ;
        RECT 620.400 568.050 621.450 604.950 ;
        RECT 619.950 565.950 622.050 568.050 ;
        RECT 623.400 565.050 624.450 610.950 ;
        RECT 626.400 601.050 627.450 619.950 ;
        RECT 635.400 610.050 636.450 646.950 ;
        RECT 637.950 639.300 640.050 641.400 ;
        RECT 638.250 635.700 639.450 639.300 ;
        RECT 637.950 633.600 640.050 635.700 ;
        RECT 638.250 621.600 639.450 633.600 ;
        RECT 641.400 628.050 642.450 655.950 ;
        RECT 643.950 631.950 646.050 634.050 ;
        RECT 640.950 625.950 643.050 628.050 ;
        RECT 640.950 623.850 643.050 624.750 ;
        RECT 637.950 619.500 640.050 621.600 ;
        RECT 634.950 607.950 637.050 610.050 ;
        RECT 625.950 598.950 628.050 601.050 ;
        RECT 631.950 600.450 634.050 601.050 ;
        RECT 629.400 599.400 634.050 600.450 ;
        RECT 629.400 598.050 630.450 599.400 ;
        RECT 631.950 598.950 634.050 599.400 ;
        RECT 625.950 596.850 628.050 597.750 ;
        RECT 628.950 595.950 631.050 598.050 ;
        RECT 631.950 596.850 634.050 597.750 ;
        RECT 634.950 596.250 636.750 597.150 ;
        RECT 637.950 595.950 640.050 598.050 ;
        RECT 641.250 596.250 643.050 597.150 ;
        RECT 629.400 574.050 630.450 595.950 ;
        RECT 634.950 592.950 637.050 595.050 ;
        RECT 638.250 593.850 639.750 594.750 ;
        RECT 640.950 592.950 643.050 595.050 ;
        RECT 628.950 571.950 631.050 574.050 ;
        RECT 622.950 562.950 625.050 565.050 ;
        RECT 622.950 560.250 625.050 561.150 ;
        RECT 631.950 559.950 634.050 562.050 ;
        RECT 632.400 559.050 633.450 559.950 ;
        RECT 610.950 556.950 613.050 559.050 ;
        RECT 613.950 557.250 615.750 558.150 ;
        RECT 616.950 556.950 619.050 559.050 ;
        RECT 620.250 557.250 621.750 558.150 ;
        RECT 622.950 556.950 625.050 559.050 ;
        RECT 631.950 556.950 634.050 559.050 ;
        RECT 611.400 553.050 612.450 556.950 ;
        RECT 623.400 556.050 624.450 556.950 ;
        RECT 613.950 553.950 616.050 556.050 ;
        RECT 617.250 554.850 618.750 555.750 ;
        RECT 619.950 553.950 622.050 556.050 ;
        RECT 622.950 553.950 625.050 556.050 ;
        RECT 625.950 553.950 628.050 556.050 ;
        RECT 628.950 554.250 631.050 555.150 ;
        RECT 631.950 554.850 634.050 555.750 ;
        RECT 605.400 551.400 609.450 552.450 ;
        RECT 589.950 544.950 592.050 547.050 ;
        RECT 589.950 541.950 592.050 544.050 ;
        RECT 586.950 532.950 589.050 535.050 ;
        RECT 584.400 530.400 588.450 531.450 ;
        RECT 587.400 529.050 588.450 530.400 ;
        RECT 583.950 526.950 586.050 529.050 ;
        RECT 586.950 526.950 589.050 529.050 ;
        RECT 578.400 503.400 582.450 504.450 ;
        RECT 568.950 490.950 571.050 493.050 ;
        RECT 574.950 490.950 577.050 493.050 ;
        RECT 569.400 490.050 570.450 490.950 ;
        RECT 575.400 490.050 576.450 490.950 ;
        RECT 568.950 487.950 571.050 490.050 ;
        RECT 572.250 488.250 573.750 489.150 ;
        RECT 574.950 487.950 577.050 490.050 ;
        RECT 568.950 485.850 570.750 486.750 ;
        RECT 571.950 484.950 574.050 487.050 ;
        RECT 575.250 485.850 577.050 486.750 ;
        RECT 572.400 484.050 573.450 484.950 ;
        RECT 571.950 481.950 574.050 484.050 ;
        RECT 574.950 481.950 577.050 484.050 ;
        RECT 578.400 483.450 579.450 503.400 ;
        RECT 584.400 487.050 585.450 526.950 ;
        RECT 586.950 524.850 589.050 525.750 ;
        RECT 586.950 520.950 589.050 523.050 ;
        RECT 587.400 490.050 588.450 520.950 ;
        RECT 590.400 490.050 591.450 541.950 ;
        RECT 592.950 535.950 595.050 538.050 ;
        RECT 593.400 529.050 594.450 535.950 ;
        RECT 592.950 526.950 595.050 529.050 ;
        RECT 592.950 524.850 595.050 525.750 ;
        RECT 596.400 523.050 597.450 550.950 ;
        RECT 602.400 550.050 603.450 550.950 ;
        RECT 601.950 547.950 604.050 550.050 ;
        RECT 598.950 533.400 601.050 535.500 ;
        RECT 595.950 520.950 598.050 523.050 ;
        RECT 599.400 516.600 600.600 533.400 ;
        RECT 602.400 532.050 603.450 547.950 ;
        RECT 601.950 529.950 604.050 532.050 ;
        RECT 601.950 526.950 604.050 529.050 ;
        RECT 602.400 523.050 603.450 526.950 ;
        RECT 601.950 520.950 604.050 523.050 ;
        RECT 605.400 520.050 606.450 551.400 ;
        RECT 610.950 550.950 613.050 553.050 ;
        RECT 607.950 547.950 610.050 550.050 ;
        RECT 610.950 547.950 613.050 550.050 ;
        RECT 604.950 517.950 607.050 520.050 ;
        RECT 598.950 514.500 601.050 516.600 ;
        RECT 601.950 511.950 604.050 514.050 ;
        RECT 598.950 496.950 601.050 499.050 ;
        RECT 586.950 487.950 589.050 490.050 ;
        RECT 589.950 487.950 592.050 490.050 ;
        RECT 595.950 487.950 598.050 490.050 ;
        RECT 580.950 485.250 582.750 486.150 ;
        RECT 583.950 484.950 586.050 487.050 ;
        RECT 587.250 485.250 588.750 486.150 ;
        RECT 589.950 484.950 592.050 487.050 ;
        RECT 593.250 485.250 595.050 486.150 ;
        RECT 596.400 484.050 597.450 487.950 ;
        RECT 580.950 483.450 583.050 484.050 ;
        RECT 578.400 482.400 583.050 483.450 ;
        RECT 584.250 482.850 585.750 483.750 ;
        RECT 580.950 481.950 583.050 482.400 ;
        RECT 586.950 481.950 589.050 484.050 ;
        RECT 590.250 482.850 591.750 483.750 ;
        RECT 592.950 481.950 595.050 484.050 ;
        RECT 595.950 481.950 598.050 484.050 ;
        RECT 568.950 478.950 571.050 481.050 ;
        RECT 559.950 469.950 562.050 472.050 ;
        RECT 565.950 469.950 568.050 472.050 ;
        RECT 556.950 466.950 559.050 469.050 ;
        RECT 560.400 463.050 561.450 469.950 ;
        RECT 553.950 460.950 556.050 463.050 ;
        RECT 559.950 460.950 562.050 463.050 ;
        RECT 560.400 457.050 561.450 460.950 ;
        RECT 562.950 457.950 565.050 460.050 ;
        RECT 550.950 456.450 553.050 457.050 ;
        RECT 553.950 456.450 556.050 457.050 ;
        RECT 550.950 455.400 556.050 456.450 ;
        RECT 550.950 454.950 553.050 455.400 ;
        RECT 553.950 454.950 556.050 455.400 ;
        RECT 557.250 455.250 558.750 456.150 ;
        RECT 559.950 454.950 562.050 457.050 ;
        RECT 562.950 455.850 565.050 456.750 ;
        RECT 565.950 455.250 568.050 456.150 ;
        RECT 550.950 453.450 553.050 454.050 ;
        RECT 548.400 452.400 553.050 453.450 ;
        RECT 554.250 452.850 555.750 453.750 ;
        RECT 544.950 445.950 547.050 448.050 ;
        RECT 548.400 415.050 549.450 452.400 ;
        RECT 550.950 451.950 553.050 452.400 ;
        RECT 556.950 451.950 559.050 454.050 ;
        RECT 560.250 452.850 562.050 453.750 ;
        RECT 565.950 451.950 568.050 454.050 ;
        RECT 550.950 449.850 553.050 450.750 ;
        RECT 553.950 448.950 556.050 451.050 ;
        RECT 557.400 450.450 558.450 451.950 ;
        RECT 566.400 450.450 567.450 451.950 ;
        RECT 557.400 449.400 567.450 450.450 ;
        RECT 554.400 445.050 555.450 448.950 ;
        RECT 553.950 442.950 556.050 445.050 ;
        RECT 559.950 442.950 562.050 445.050 ;
        RECT 556.950 427.950 559.050 430.050 ;
        RECT 553.950 415.950 556.050 418.050 ;
        RECT 544.950 413.250 547.050 414.150 ;
        RECT 547.950 412.950 550.050 415.050 ;
        RECT 550.950 413.250 553.050 414.150 ;
        RECT 544.950 409.950 547.050 412.050 ;
        RECT 550.950 409.950 553.050 412.050 ;
        RECT 545.400 406.050 546.450 409.950 ;
        RECT 551.400 409.050 552.450 409.950 ;
        RECT 550.950 406.950 553.050 409.050 ;
        RECT 544.950 403.950 547.050 406.050 ;
        RECT 535.950 400.950 538.050 403.050 ;
        RECT 541.950 400.950 544.050 403.050 ;
        RECT 533.400 398.400 537.450 399.450 ;
        RECT 526.950 391.950 529.050 394.050 ;
        RECT 527.400 381.450 528.450 391.950 ;
        RECT 532.950 385.950 535.050 388.050 ;
        RECT 529.950 383.250 532.050 384.150 ;
        RECT 532.950 383.850 535.050 384.750 ;
        RECT 529.950 381.450 532.050 382.050 ;
        RECT 527.400 380.400 532.050 381.450 ;
        RECT 529.950 379.950 532.050 380.400 ;
        RECT 532.950 379.950 535.050 382.050 ;
        RECT 529.950 376.950 532.050 379.050 ;
        RECT 514.950 364.950 517.050 367.050 ;
        RECT 523.950 364.950 526.050 367.050 ;
        RECT 515.400 346.050 516.450 364.950 ;
        RECT 517.950 358.950 520.050 361.050 ;
        RECT 526.950 358.950 529.050 361.050 ;
        RECT 511.950 344.250 514.050 345.150 ;
        RECT 514.950 343.950 517.050 346.050 ;
        RECT 518.400 343.050 519.450 358.950 ;
        RECT 527.400 343.050 528.450 358.950 ;
        RECT 530.400 346.050 531.450 376.950 ;
        RECT 533.400 348.450 534.450 379.950 ;
        RECT 536.400 364.050 537.450 398.400 ;
        RECT 547.950 385.950 550.050 388.050 ;
        RECT 541.950 382.950 544.050 385.050 ;
        RECT 542.400 382.050 543.450 382.950 ;
        RECT 548.400 382.050 549.450 385.950 ;
        RECT 538.950 380.250 540.750 381.150 ;
        RECT 541.950 379.950 544.050 382.050 ;
        RECT 547.950 379.950 550.050 382.050 ;
        RECT 538.950 376.950 541.050 379.050 ;
        RECT 542.250 377.850 543.750 378.750 ;
        RECT 544.950 376.950 547.050 379.050 ;
        RECT 548.250 377.850 550.050 378.750 ;
        RECT 539.400 373.050 540.450 376.950 ;
        RECT 551.400 376.050 552.450 406.950 ;
        RECT 554.400 382.050 555.450 415.950 ;
        RECT 557.400 409.050 558.450 427.950 ;
        RECT 556.950 406.950 559.050 409.050 ;
        RECT 560.400 391.050 561.450 442.950 ;
        RECT 569.400 436.050 570.450 478.950 ;
        RECT 575.400 469.050 576.450 481.950 ;
        RECT 587.400 481.050 588.450 481.950 ;
        RECT 580.950 478.950 583.050 481.050 ;
        RECT 586.950 478.950 589.050 481.050 ;
        RECT 581.400 475.050 582.450 478.950 ;
        RECT 593.400 475.050 594.450 481.950 ;
        RECT 595.950 478.950 598.050 481.050 ;
        RECT 596.400 475.050 597.450 478.950 ;
        RECT 580.950 472.950 583.050 475.050 ;
        RECT 592.950 472.950 595.050 475.050 ;
        RECT 595.950 472.950 598.050 475.050 ;
        RECT 599.400 472.050 600.450 496.950 ;
        RECT 602.400 496.050 603.450 511.950 ;
        RECT 608.400 511.050 609.450 547.950 ;
        RECT 611.400 547.050 612.450 547.950 ;
        RECT 610.950 544.950 613.050 547.050 ;
        RECT 614.400 541.050 615.450 553.950 ;
        RECT 620.400 552.450 621.450 553.950 ;
        RECT 626.400 552.450 627.450 553.950 ;
        RECT 620.400 551.400 627.450 552.450 ;
        RECT 628.950 550.950 631.050 553.050 ;
        RECT 622.950 544.950 625.050 547.050 ;
        RECT 619.950 541.950 622.050 544.050 ;
        RECT 613.950 538.950 616.050 541.050 ;
        RECT 620.400 538.050 621.450 541.950 ;
        RECT 616.950 535.950 619.050 538.050 ;
        RECT 619.950 535.950 622.050 538.050 ;
        RECT 610.950 532.950 613.050 535.050 ;
        RECT 611.400 529.050 612.450 532.950 ;
        RECT 617.400 529.050 618.450 535.950 ;
        RECT 610.950 526.950 613.050 529.050 ;
        RECT 614.250 527.250 615.750 528.150 ;
        RECT 616.950 526.950 619.050 529.050 ;
        RECT 619.950 526.950 622.050 529.050 ;
        RECT 620.400 526.050 621.450 526.950 ;
        RECT 610.950 524.850 612.750 525.750 ;
        RECT 613.950 523.950 616.050 526.050 ;
        RECT 617.250 524.850 618.750 525.750 ;
        RECT 619.950 523.950 622.050 526.050 ;
        RECT 613.950 520.950 616.050 523.050 ;
        RECT 619.950 521.850 622.050 522.750 ;
        RECT 610.950 517.950 613.050 520.050 ;
        RECT 607.950 508.950 610.050 511.050 ;
        RECT 607.950 502.950 610.050 505.050 ;
        RECT 601.950 493.950 604.050 496.050 ;
        RECT 608.400 493.050 609.450 502.950 ;
        RECT 601.950 490.950 604.050 493.050 ;
        RECT 607.950 490.950 610.050 493.050 ;
        RECT 602.400 490.050 603.450 490.950 ;
        RECT 601.950 487.950 604.050 490.050 ;
        RECT 605.250 488.250 606.750 489.150 ;
        RECT 607.950 487.950 610.050 490.050 ;
        RECT 601.950 485.850 603.750 486.750 ;
        RECT 604.950 484.950 607.050 487.050 ;
        RECT 608.250 485.850 610.050 486.750 ;
        RECT 601.950 481.950 604.050 484.050 ;
        RECT 589.950 469.950 592.050 472.050 ;
        RECT 598.950 469.950 601.050 472.050 ;
        RECT 574.950 466.950 577.050 469.050 ;
        RECT 586.950 466.950 589.050 469.050 ;
        RECT 571.950 463.950 574.050 466.050 ;
        RECT 572.400 457.050 573.450 463.950 ;
        RECT 571.950 454.950 574.050 457.050 ;
        RECT 575.250 455.250 576.750 456.150 ;
        RECT 577.950 454.950 580.050 457.050 ;
        RECT 583.950 454.950 586.050 457.050 ;
        RECT 571.950 452.850 573.750 453.750 ;
        RECT 574.950 451.950 577.050 454.050 ;
        RECT 578.250 452.850 579.750 453.750 ;
        RECT 580.950 451.950 583.050 454.050 ;
        RECT 580.950 449.850 583.050 450.750 ;
        RECT 574.950 445.950 577.050 448.050 ;
        RECT 568.950 433.950 571.050 436.050 ;
        RECT 568.950 419.250 571.050 420.150 ;
        RECT 562.950 415.950 565.050 418.050 ;
        RECT 566.250 416.250 567.750 417.150 ;
        RECT 568.950 415.950 571.050 418.050 ;
        RECT 572.250 416.250 574.050 417.150 ;
        RECT 562.950 413.850 564.750 414.750 ;
        RECT 565.950 412.950 568.050 415.050 ;
        RECT 571.950 412.950 574.050 415.050 ;
        RECT 565.950 406.950 568.050 409.050 ;
        RECT 562.950 391.950 565.050 394.050 ;
        RECT 559.950 388.950 562.050 391.050 ;
        RECT 559.950 382.950 562.050 385.050 ;
        RECT 560.400 382.050 561.450 382.950 ;
        RECT 553.950 379.950 556.050 382.050 ;
        RECT 556.950 380.250 558.750 381.150 ;
        RECT 559.950 379.950 562.050 382.050 ;
        RECT 563.400 379.050 564.450 391.950 ;
        RECT 566.400 382.050 567.450 406.950 ;
        RECT 572.400 403.050 573.450 412.950 ;
        RECT 571.950 400.950 574.050 403.050 ;
        RECT 571.950 394.950 574.050 397.050 ;
        RECT 568.950 388.950 571.050 391.050 ;
        RECT 565.950 379.950 568.050 382.050 ;
        RECT 556.950 376.950 559.050 379.050 ;
        RECT 560.250 377.850 561.750 378.750 ;
        RECT 562.950 376.950 565.050 379.050 ;
        RECT 566.250 377.850 568.050 378.750 ;
        RECT 544.950 374.850 547.050 375.750 ;
        RECT 550.950 373.950 553.050 376.050 ;
        RECT 538.950 370.950 541.050 373.050 ;
        RECT 553.950 367.950 556.050 370.050 ;
        RECT 535.950 361.950 538.050 364.050 ;
        RECT 538.950 355.950 541.050 358.050 ;
        RECT 533.400 347.400 537.450 348.450 ;
        RECT 529.950 343.950 532.050 346.050 ;
        RECT 532.950 344.250 535.050 345.150 ;
        RECT 511.950 340.950 514.050 343.050 ;
        RECT 515.250 341.250 516.750 342.150 ;
        RECT 517.950 340.950 520.050 343.050 ;
        RECT 521.250 341.250 523.050 342.150 ;
        RECT 523.950 341.250 525.750 342.150 ;
        RECT 526.950 340.950 529.050 343.050 ;
        RECT 530.250 341.250 531.750 342.150 ;
        RECT 532.950 340.950 535.050 343.050 ;
        RECT 512.400 334.050 513.450 340.950 ;
        RECT 514.950 337.950 517.050 340.050 ;
        RECT 518.250 338.850 519.750 339.750 ;
        RECT 520.950 337.950 523.050 340.050 ;
        RECT 523.950 337.950 526.050 340.050 ;
        RECT 527.250 338.850 528.750 339.750 ;
        RECT 529.950 337.950 532.050 340.050 ;
        RECT 532.950 337.950 535.050 340.050 ;
        RECT 515.400 337.050 516.450 337.950 ;
        RECT 514.950 334.950 517.050 337.050 ;
        RECT 520.950 334.950 523.050 337.050 ;
        RECT 511.950 331.950 514.050 334.050 ;
        RECT 511.950 325.950 514.050 328.050 ;
        RECT 514.950 325.950 517.050 328.050 ;
        RECT 512.400 313.050 513.450 325.950 ;
        RECT 515.400 313.050 516.450 325.950 ;
        RECT 517.950 322.950 520.050 325.050 ;
        RECT 511.950 310.950 514.050 313.050 ;
        RECT 514.950 310.950 517.050 313.050 ;
        RECT 511.950 308.250 514.050 309.150 ;
        RECT 514.950 308.850 517.050 309.750 ;
        RECT 518.400 307.050 519.450 322.950 ;
        RECT 511.950 304.950 514.050 307.050 ;
        RECT 517.950 304.950 520.050 307.050 ;
        RECT 512.400 304.050 513.450 304.950 ;
        RECT 511.950 301.950 514.050 304.050 ;
        RECT 521.400 301.050 522.450 334.950 ;
        RECT 524.400 334.050 525.450 337.950 ;
        RECT 523.950 331.950 526.050 334.050 ;
        RECT 526.950 331.950 529.050 334.050 ;
        RECT 527.400 319.050 528.450 331.950 ;
        RECT 530.400 319.050 531.450 337.950 ;
        RECT 526.950 316.950 529.050 319.050 ;
        RECT 529.950 316.950 532.050 319.050 ;
        RECT 526.950 310.950 529.050 313.050 ;
        RECT 527.400 310.050 528.450 310.950 ;
        RECT 523.950 308.250 525.750 309.150 ;
        RECT 526.950 307.950 529.050 310.050 ;
        RECT 530.250 308.250 532.050 309.150 ;
        RECT 523.950 304.950 526.050 307.050 ;
        RECT 527.250 305.850 528.750 306.750 ;
        RECT 529.950 304.950 532.050 307.050 ;
        RECT 517.950 298.950 520.050 301.050 ;
        RECT 520.950 298.950 523.050 301.050 ;
        RECT 526.950 298.950 529.050 301.050 ;
        RECT 508.950 295.950 511.050 298.050 ;
        RECT 511.950 292.950 514.050 295.050 ;
        RECT 503.400 275.400 507.450 276.450 ;
        RECT 503.400 274.050 504.450 275.400 ;
        RECT 499.950 271.950 502.050 274.050 ;
        RECT 502.950 271.950 505.050 274.050 ;
        RECT 506.250 272.250 507.750 273.150 ;
        RECT 508.950 271.950 511.050 274.050 ;
        RECT 499.950 269.250 502.050 270.150 ;
        RECT 502.950 269.850 504.750 270.750 ;
        RECT 505.950 268.950 508.050 271.050 ;
        RECT 509.250 269.850 511.050 270.750 ;
        RECT 499.950 265.950 502.050 268.050 ;
        RECT 505.950 265.950 508.050 268.050 ;
        RECT 512.400 267.450 513.450 292.950 ;
        RECT 518.400 273.450 519.450 298.950 ;
        RECT 527.400 277.050 528.450 298.950 ;
        RECT 533.400 292.050 534.450 337.950 ;
        RECT 536.400 325.050 537.450 347.400 ;
        RECT 539.400 343.050 540.450 355.950 ;
        RECT 554.400 352.050 555.450 367.950 ;
        RECT 557.400 355.050 558.450 376.950 ;
        RECT 562.950 374.850 565.050 375.750 ;
        RECT 569.400 375.450 570.450 388.950 ;
        RECT 572.400 382.050 573.450 394.950 ;
        RECT 575.400 391.050 576.450 445.950 ;
        RECT 580.950 433.950 583.050 436.050 ;
        RECT 581.400 430.050 582.450 433.950 ;
        RECT 580.950 427.950 583.050 430.050 ;
        RECT 580.950 415.950 583.050 418.050 ;
        RECT 581.400 415.050 582.450 415.950 ;
        RECT 580.950 414.450 583.050 415.050 ;
        RECT 584.400 414.450 585.450 454.950 ;
        RECT 587.400 439.050 588.450 466.950 ;
        RECT 590.400 447.450 591.450 469.950 ;
        RECT 602.400 469.050 603.450 481.950 ;
        RECT 605.400 480.450 606.450 484.950 ;
        RECT 607.950 480.450 610.050 481.050 ;
        RECT 605.400 479.400 610.050 480.450 ;
        RECT 607.950 478.950 610.050 479.400 ;
        RECT 592.950 466.950 595.050 469.050 ;
        RECT 601.950 466.950 604.050 469.050 ;
        RECT 593.400 457.050 594.450 466.950 ;
        RECT 601.950 463.950 604.050 466.050 ;
        RECT 598.950 460.950 601.050 463.050 ;
        RECT 592.950 454.950 595.050 457.050 ;
        RECT 595.950 454.950 598.050 457.050 ;
        RECT 596.400 454.050 597.450 454.950 ;
        RECT 592.950 452.250 594.750 453.150 ;
        RECT 595.950 451.950 598.050 454.050 ;
        RECT 599.400 451.050 600.450 460.950 ;
        RECT 602.400 454.050 603.450 463.950 ;
        RECT 611.400 460.050 612.450 517.950 ;
        RECT 614.400 511.050 615.450 520.950 ;
        RECT 616.950 514.950 619.050 517.050 ;
        RECT 613.950 508.950 616.050 511.050 ;
        RECT 617.400 493.050 618.450 514.950 ;
        RECT 616.950 490.950 619.050 493.050 ;
        RECT 617.400 487.050 618.450 490.950 ;
        RECT 613.950 485.250 616.050 486.150 ;
        RECT 616.950 484.950 619.050 487.050 ;
        RECT 619.950 485.250 622.050 486.150 ;
        RECT 613.950 481.950 616.050 484.050 ;
        RECT 617.250 482.250 618.750 483.150 ;
        RECT 619.950 481.950 622.050 484.050 ;
        RECT 614.400 481.050 615.450 481.950 ;
        RECT 613.950 478.950 616.050 481.050 ;
        RECT 616.950 478.950 619.050 481.050 ;
        RECT 617.400 475.050 618.450 478.950 ;
        RECT 616.950 472.950 619.050 475.050 ;
        RECT 620.400 469.050 621.450 481.950 ;
        RECT 619.950 466.950 622.050 469.050 ;
        RECT 613.950 460.950 616.050 463.050 ;
        RECT 623.400 462.450 624.450 544.950 ;
        RECT 635.400 541.050 636.450 592.950 ;
        RECT 640.950 589.950 643.050 592.050 ;
        RECT 637.950 571.950 640.050 574.050 ;
        RECT 634.950 538.950 637.050 541.050 ;
        RECT 638.400 529.050 639.450 571.950 ;
        RECT 641.400 550.050 642.450 589.950 ;
        RECT 644.400 586.050 645.450 631.950 ;
        RECT 649.950 630.450 652.050 631.050 ;
        RECT 653.400 630.450 654.450 667.950 ;
        RECT 659.250 658.050 660.450 676.950 ;
        RECT 662.250 664.350 663.450 676.950 ;
        RECT 661.950 662.250 664.050 664.350 ;
        RECT 662.250 658.050 663.450 662.250 ;
        RECT 665.250 658.050 666.450 676.950 ;
        RECT 658.950 655.950 661.050 658.050 ;
        RECT 661.950 655.950 664.050 658.050 ;
        RECT 664.950 655.950 667.050 658.050 ;
        RECT 658.950 649.950 661.050 652.050 ;
        RECT 659.400 631.050 660.450 649.950 ;
        RECT 668.400 634.050 669.450 697.950 ;
        RECT 671.400 682.050 672.450 704.400 ;
        RECT 673.950 703.950 676.050 704.400 ;
        RECT 709.950 704.250 712.050 705.150 ;
        RECT 673.950 701.850 676.050 702.750 ;
        RECT 682.950 701.250 684.750 702.150 ;
        RECT 685.950 700.950 688.050 703.050 ;
        RECT 691.950 702.450 694.050 703.050 ;
        RECT 691.950 701.400 696.450 702.450 ;
        RECT 691.950 700.950 694.050 701.400 ;
        RECT 682.950 697.950 685.050 700.050 ;
        RECT 686.250 698.850 688.050 699.750 ;
        RECT 688.950 698.250 691.050 699.150 ;
        RECT 691.950 698.850 694.050 699.750 ;
        RECT 670.950 679.950 673.050 682.050 ;
        RECT 671.400 670.050 672.450 679.950 ;
        RECT 670.950 667.950 673.050 670.050 ;
        RECT 676.950 668.250 679.050 669.150 ;
        RECT 670.950 665.850 673.050 666.750 ;
        RECT 670.950 658.950 673.050 661.050 ;
        RECT 661.950 631.950 664.050 634.050 ;
        RECT 664.950 632.250 667.050 633.150 ;
        RECT 667.950 631.950 670.050 634.050 ;
        RECT 649.950 629.400 654.450 630.450 ;
        RECT 649.950 628.950 652.050 629.400 ;
        RECT 655.950 629.250 658.050 630.150 ;
        RECT 658.950 628.950 661.050 631.050 ;
        RECT 646.950 625.950 649.050 628.050 ;
        RECT 649.950 626.850 652.050 627.750 ;
        RECT 652.950 625.950 655.050 628.050 ;
        RECT 655.950 625.950 658.050 628.050 ;
        RECT 659.250 626.250 661.050 627.150 ;
        RECT 647.400 616.050 648.450 625.950 ;
        RECT 646.950 613.950 649.050 616.050 ;
        RECT 653.400 607.050 654.450 625.950 ;
        RECT 656.400 616.050 657.450 625.950 ;
        RECT 658.950 622.950 661.050 625.050 ;
        RECT 655.950 613.950 658.050 616.050 ;
        RECT 662.400 613.050 663.450 631.950 ;
        RECT 671.400 631.050 672.450 658.950 ;
        RECT 683.400 649.050 684.450 697.950 ;
        RECT 688.950 694.950 691.050 697.050 ;
        RECT 685.950 668.250 687.750 669.150 ;
        RECT 688.950 667.950 691.050 670.050 ;
        RECT 692.250 668.250 694.050 669.150 ;
        RECT 685.950 664.950 688.050 667.050 ;
        RECT 689.250 665.850 690.750 666.750 ;
        RECT 691.950 664.950 694.050 667.050 ;
        RECT 682.950 646.950 685.050 649.050 ;
        RECT 686.400 646.050 687.450 664.950 ;
        RECT 695.400 664.050 696.450 701.400 ;
        RECT 697.950 700.950 700.050 703.050 ;
        RECT 709.950 700.950 712.050 703.050 ;
        RECT 697.950 698.850 700.050 699.750 ;
        RECT 710.400 691.050 711.450 700.950 ;
        RECT 719.550 693.600 720.750 707.250 ;
        RECT 722.250 693.600 723.450 710.850 ;
        RECT 729.900 710.400 732.000 712.500 ;
        RECT 733.950 710.400 736.050 712.500 ;
        RECT 724.950 707.250 727.050 709.350 ;
        RECT 725.400 693.600 726.600 707.250 ;
        RECT 730.350 701.550 731.550 710.400 ;
        RECT 734.550 704.250 735.750 710.400 ;
        RECT 733.950 702.150 736.050 704.250 ;
        RECT 729.750 699.450 731.850 701.550 ;
        RECT 730.350 693.600 731.550 699.450 ;
        RECT 734.550 693.600 735.750 702.150 ;
        RECT 736.950 698.250 739.050 699.150 ;
        RECT 736.950 694.950 739.050 697.050 ;
        RECT 718.950 691.500 721.050 693.600 ;
        RECT 721.950 691.500 724.050 693.600 ;
        RECT 724.950 691.500 727.050 693.600 ;
        RECT 729.750 691.500 731.850 693.600 ;
        RECT 733.950 691.500 736.050 693.600 ;
        RECT 709.950 688.950 712.050 691.050 ;
        RECT 721.950 673.950 724.050 676.050 ;
        RECT 737.400 673.050 738.450 694.950 ;
        RECT 743.250 694.050 744.450 712.950 ;
        RECT 746.250 708.750 747.450 712.950 ;
        RECT 745.950 706.650 748.050 708.750 ;
        RECT 746.250 694.050 747.450 706.650 ;
        RECT 749.250 694.050 750.450 712.950 ;
        RECT 760.950 705.450 763.050 706.050 ;
        RECT 754.950 704.250 757.050 705.150 ;
        RECT 758.400 704.400 763.050 705.450 ;
        RECT 742.950 691.950 745.050 694.050 ;
        RECT 745.950 691.950 748.050 694.050 ;
        RECT 748.950 691.950 751.050 694.050 ;
        RECT 758.400 682.050 759.450 704.400 ;
        RECT 760.950 703.950 763.050 704.400 ;
        RECT 760.950 701.850 763.050 702.750 ;
        RECT 757.950 679.950 760.050 682.050 ;
        RECT 760.950 679.950 763.050 682.050 ;
        RECT 703.950 670.950 706.050 673.050 ;
        RECT 707.250 671.250 708.750 672.150 ;
        RECT 709.950 670.950 712.050 673.050 ;
        RECT 718.950 672.450 721.050 673.050 ;
        RECT 716.400 671.400 721.050 672.450 ;
        RECT 722.250 671.850 723.750 672.750 ;
        RECT 704.250 668.850 705.750 669.750 ;
        RECT 706.950 667.950 709.050 670.050 ;
        RECT 710.250 668.850 712.050 669.750 ;
        RECT 700.950 665.850 703.050 666.750 ;
        RECT 709.950 664.950 712.050 667.050 ;
        RECT 694.950 661.950 697.050 664.050 ;
        RECT 676.950 643.950 679.050 646.050 ;
        RECT 685.950 643.950 688.050 646.050 ;
        RECT 677.400 634.050 678.450 643.950 ;
        RECT 700.950 637.950 703.050 640.050 ;
        RECT 691.950 634.950 694.050 637.050 ;
        RECT 676.950 631.950 679.050 634.050 ;
        RECT 679.950 632.250 682.050 633.150 ;
        RECT 664.950 628.950 667.050 631.050 ;
        RECT 668.250 629.250 669.750 630.150 ;
        RECT 670.950 628.950 673.050 631.050 ;
        RECT 674.250 629.250 676.050 630.150 ;
        RECT 676.950 628.950 679.050 631.050 ;
        RECT 679.950 628.950 682.050 631.050 ;
        RECT 683.250 629.250 684.750 630.150 ;
        RECT 689.250 629.250 691.050 630.150 ;
        RECT 655.950 610.950 658.050 613.050 ;
        RECT 661.950 610.950 664.050 613.050 ;
        RECT 652.950 604.950 655.050 607.050 ;
        RECT 652.950 601.950 655.050 604.050 ;
        RECT 656.400 601.050 657.450 610.950 ;
        RECT 661.950 604.950 664.050 607.050 ;
        RECT 662.400 604.050 663.450 604.950 ;
        RECT 665.400 604.050 666.450 628.950 ;
        RECT 667.950 625.950 670.050 628.050 ;
        RECT 671.250 626.850 672.750 627.750 ;
        RECT 673.950 625.950 676.050 628.050 ;
        RECT 668.400 625.050 669.450 625.950 ;
        RECT 667.950 622.950 670.050 625.050 ;
        RECT 677.400 619.050 678.450 628.950 ;
        RECT 679.950 625.950 682.050 628.050 ;
        RECT 682.950 625.950 685.050 628.050 ;
        RECT 686.250 626.850 687.750 627.750 ;
        RECT 692.400 627.450 693.450 634.950 ;
        RECT 701.400 633.450 702.450 637.950 ;
        RECT 698.400 632.400 702.450 633.450 ;
        RECT 710.400 633.450 711.450 664.950 ;
        RECT 716.400 661.050 717.450 671.400 ;
        RECT 718.950 670.950 721.050 671.400 ;
        RECT 736.950 670.950 739.050 673.050 ;
        RECT 745.950 671.850 748.050 672.750 ;
        RECT 748.950 671.250 751.050 672.150 ;
        RECT 751.950 670.950 754.050 673.050 ;
        RECT 754.950 671.850 757.050 672.750 ;
        RECT 757.950 671.250 760.050 672.150 ;
        RECT 718.950 668.850 721.050 669.750 ;
        RECT 721.950 667.950 724.050 670.050 ;
        RECT 724.950 668.850 727.050 669.750 ;
        RECT 730.950 668.250 732.750 669.150 ;
        RECT 733.950 667.950 736.050 670.050 ;
        RECT 739.950 667.950 742.050 670.050 ;
        RECT 748.950 667.950 751.050 670.050 ;
        RECT 718.950 661.950 721.050 664.050 ;
        RECT 715.950 658.950 718.050 661.050 ;
        RECT 715.950 643.950 718.050 646.050 ;
        RECT 716.400 634.050 717.450 643.950 ;
        RECT 710.400 632.400 714.450 633.450 ;
        RECT 698.400 631.050 699.450 632.400 ;
        RECT 713.400 631.050 714.450 632.400 ;
        RECT 715.950 631.950 718.050 634.050 ;
        RECT 694.950 629.250 696.750 630.150 ;
        RECT 697.950 628.950 700.050 631.050 ;
        RECT 701.250 629.250 702.750 630.150 ;
        RECT 703.950 628.950 706.050 631.050 ;
        RECT 707.250 629.250 709.050 630.150 ;
        RECT 712.950 628.950 715.050 631.050 ;
        RECT 694.950 627.450 697.050 628.050 ;
        RECT 692.400 626.400 697.050 627.450 ;
        RECT 698.250 626.850 699.750 627.750 ;
        RECT 694.950 625.950 697.050 626.400 ;
        RECT 700.950 625.950 703.050 628.050 ;
        RECT 704.250 626.850 705.750 627.750 ;
        RECT 706.950 625.950 709.050 628.050 ;
        RECT 709.950 626.250 712.050 627.150 ;
        RECT 712.950 626.850 715.050 627.750 ;
        RECT 680.400 625.050 681.450 625.950 ;
        RECT 679.950 622.950 682.050 625.050 ;
        RECT 685.950 622.950 688.050 625.050 ;
        RECT 667.950 616.950 670.050 619.050 ;
        RECT 676.950 616.950 679.050 619.050 ;
        RECT 682.950 616.950 685.050 619.050 ;
        RECT 661.950 601.950 664.050 604.050 ;
        RECT 664.950 601.950 667.050 604.050 ;
        RECT 668.400 601.050 669.450 616.950 ;
        RECT 670.950 607.950 673.050 610.050 ;
        RECT 649.950 598.950 652.050 601.050 ;
        RECT 653.250 599.850 654.750 600.750 ;
        RECT 655.950 598.950 658.050 601.050 ;
        RECT 658.950 599.250 661.050 600.150 ;
        RECT 661.950 599.850 664.050 600.750 ;
        RECT 664.950 599.250 666.750 600.150 ;
        RECT 667.950 598.950 670.050 601.050 ;
        RECT 649.950 596.850 652.050 597.750 ;
        RECT 652.950 595.950 655.050 598.050 ;
        RECT 655.950 596.850 658.050 597.750 ;
        RECT 658.950 595.950 661.050 598.050 ;
        RECT 661.950 595.950 664.050 598.050 ;
        RECT 664.950 595.950 667.050 598.050 ;
        RECT 668.250 596.850 670.050 597.750 ;
        RECT 643.950 583.950 646.050 586.050 ;
        RECT 646.950 562.950 649.050 565.050 ;
        RECT 649.950 562.950 652.050 565.050 ;
        RECT 647.400 559.050 648.450 562.950 ;
        RECT 650.400 559.050 651.450 562.950 ;
        RECT 653.400 562.050 654.450 595.950 ;
        RECT 659.400 592.050 660.450 595.950 ;
        RECT 662.400 592.050 663.450 595.950 ;
        RECT 667.950 592.950 670.050 595.050 ;
        RECT 658.950 589.950 661.050 592.050 ;
        RECT 661.950 589.950 664.050 592.050 ;
        RECT 658.950 583.950 661.050 586.050 ;
        RECT 659.400 565.050 660.450 583.950 ;
        RECT 658.950 562.950 661.050 565.050 ;
        RECT 652.950 559.950 655.050 562.050 ;
        RECT 656.250 560.250 657.750 561.150 ;
        RECT 658.950 559.950 661.050 562.050 ;
        RECT 668.400 559.050 669.450 592.950 ;
        RECT 671.400 562.050 672.450 607.950 ;
        RECT 673.950 604.950 676.050 607.050 ;
        RECT 674.400 601.050 675.450 604.950 ;
        RECT 673.950 598.950 676.050 601.050 ;
        RECT 677.250 599.250 678.750 600.150 ;
        RECT 679.950 598.950 682.050 601.050 ;
        RECT 683.400 598.050 684.450 616.950 ;
        RECT 673.950 596.850 675.750 597.750 ;
        RECT 676.950 595.950 679.050 598.050 ;
        RECT 680.250 596.850 681.750 597.750 ;
        RECT 682.950 595.950 685.050 598.050 ;
        RECT 673.950 580.950 676.050 583.050 ;
        RECT 670.950 559.950 673.050 562.050 ;
        RECT 643.950 556.950 646.050 559.050 ;
        RECT 646.950 556.950 649.050 559.050 ;
        RECT 649.950 556.950 652.050 559.050 ;
        RECT 652.950 557.850 654.750 558.750 ;
        RECT 655.950 556.950 658.050 559.050 ;
        RECT 659.250 557.850 661.050 558.750 ;
        RECT 661.950 556.950 664.050 559.050 ;
        RECT 664.950 557.250 667.050 558.150 ;
        RECT 667.950 556.950 670.050 559.050 ;
        RECT 670.950 557.250 673.050 558.150 ;
        RECT 643.950 554.850 646.050 555.750 ;
        RECT 646.950 554.250 649.050 555.150 ;
        RECT 649.950 553.950 652.050 556.050 ;
        RECT 646.950 552.450 649.050 553.050 ;
        RECT 650.400 552.450 651.450 553.950 ;
        RECT 646.950 551.400 651.450 552.450 ;
        RECT 646.950 550.950 649.050 551.400 ;
        RECT 652.950 550.950 655.050 553.050 ;
        RECT 640.950 547.950 643.050 550.050 ;
        RECT 653.400 547.050 654.450 550.950 ;
        RECT 652.950 544.950 655.050 547.050 ;
        RECT 628.950 526.950 631.050 529.050 ;
        RECT 634.950 526.950 637.050 529.050 ;
        RECT 637.950 526.950 640.050 529.050 ;
        RECT 643.950 526.950 646.050 529.050 ;
        RECT 629.400 526.050 630.450 526.950 ;
        RECT 635.400 526.050 636.450 526.950 ;
        RECT 625.950 524.250 627.750 525.150 ;
        RECT 628.950 523.950 631.050 526.050 ;
        RECT 632.250 524.250 634.050 525.150 ;
        RECT 634.950 523.950 637.050 526.050 ;
        RECT 637.950 524.850 640.050 525.750 ;
        RECT 643.950 524.850 646.050 525.750 ;
        RECT 649.950 523.950 652.050 526.050 ;
        RECT 652.950 524.250 654.750 525.150 ;
        RECT 655.950 523.950 658.050 526.050 ;
        RECT 659.250 524.250 661.050 525.150 ;
        RECT 625.950 520.950 628.050 523.050 ;
        RECT 629.250 521.850 630.750 522.750 ;
        RECT 631.950 522.450 634.050 523.050 ;
        RECT 635.400 522.450 636.450 523.950 ;
        RECT 631.950 521.400 636.450 522.450 ;
        RECT 631.950 520.950 634.050 521.400 ;
        RECT 626.400 520.050 627.450 520.950 ;
        RECT 625.950 517.950 628.050 520.050 ;
        RECT 626.400 517.050 627.450 517.950 ;
        RECT 625.950 514.950 628.050 517.050 ;
        RECT 625.950 496.950 628.050 499.050 ;
        RECT 620.400 461.400 624.450 462.450 ;
        RECT 614.400 460.050 615.450 460.950 ;
        RECT 607.950 457.950 610.050 460.050 ;
        RECT 610.950 457.950 613.050 460.050 ;
        RECT 613.950 457.950 616.050 460.050 ;
        RECT 608.400 457.050 609.450 457.950 ;
        RECT 604.950 454.950 607.050 457.050 ;
        RECT 607.950 454.950 610.050 457.050 ;
        RECT 611.250 455.250 613.050 456.150 ;
        RECT 613.950 455.850 616.050 456.750 ;
        RECT 616.950 455.250 619.050 456.150 ;
        RECT 601.950 451.950 604.050 454.050 ;
        RECT 592.950 448.950 595.050 451.050 ;
        RECT 596.250 449.850 597.750 450.750 ;
        RECT 598.950 448.950 601.050 451.050 ;
        RECT 602.250 449.850 604.050 450.750 ;
        RECT 605.400 448.050 606.450 454.950 ;
        RECT 607.950 452.850 609.750 453.750 ;
        RECT 610.950 451.950 613.050 454.050 ;
        RECT 613.950 451.950 616.050 454.050 ;
        RECT 616.950 451.950 619.050 454.050 ;
        RECT 607.950 448.950 610.050 451.050 ;
        RECT 590.400 446.400 594.450 447.450 ;
        RECT 598.950 446.850 601.050 447.750 ;
        RECT 586.950 436.950 589.050 439.050 ;
        RECT 593.400 427.050 594.450 446.400 ;
        RECT 604.950 445.950 607.050 448.050 ;
        RECT 608.400 445.050 609.450 448.950 ;
        RECT 607.950 442.950 610.050 445.050 ;
        RECT 607.950 436.950 610.050 439.050 ;
        RECT 589.950 424.950 592.050 427.050 ;
        RECT 592.950 424.950 595.050 427.050 ;
        RECT 590.400 421.050 591.450 424.950 ;
        RECT 589.950 418.950 592.050 421.050 ;
        RECT 577.950 413.250 579.750 414.150 ;
        RECT 580.950 413.400 585.450 414.450 ;
        RECT 580.950 412.950 583.050 413.400 ;
        RECT 586.950 412.950 589.050 415.050 ;
        RECT 577.950 409.950 580.050 412.050 ;
        RECT 581.250 410.850 583.050 411.750 ;
        RECT 583.950 410.250 586.050 411.150 ;
        RECT 586.950 410.850 589.050 411.750 ;
        RECT 578.400 406.050 579.450 409.950 ;
        RECT 583.950 406.950 586.050 409.050 ;
        RECT 584.400 406.050 585.450 406.950 ;
        RECT 577.950 403.950 580.050 406.050 ;
        RECT 583.950 403.950 586.050 406.050 ;
        RECT 584.400 403.050 585.450 403.950 ;
        RECT 583.950 400.950 586.050 403.050 ;
        RECT 580.950 391.950 583.050 394.050 ;
        RECT 586.950 391.950 589.050 394.050 ;
        RECT 574.950 388.950 577.050 391.050 ;
        RECT 581.400 385.050 582.450 391.950 ;
        RECT 583.950 388.950 586.050 391.050 ;
        RECT 574.950 382.950 577.050 385.050 ;
        RECT 578.250 383.250 579.750 384.150 ;
        RECT 580.950 382.950 583.050 385.050 ;
        RECT 571.950 379.950 574.050 382.050 ;
        RECT 575.250 380.850 576.750 381.750 ;
        RECT 577.950 379.950 580.050 382.050 ;
        RECT 581.250 380.850 583.050 381.750 ;
        RECT 571.950 377.850 574.050 378.750 ;
        RECT 569.400 374.400 573.450 375.450 ;
        RECT 568.950 370.950 571.050 373.050 ;
        RECT 556.950 352.950 559.050 355.050 ;
        RECT 562.950 352.950 565.050 355.050 ;
        RECT 557.400 352.050 558.450 352.950 ;
        RECT 550.950 349.950 553.050 352.050 ;
        RECT 553.950 349.950 556.050 352.050 ;
        RECT 556.950 349.950 559.050 352.050 ;
        RECT 551.400 349.050 552.450 349.950 ;
        RECT 544.950 346.950 547.050 349.050 ;
        RECT 550.950 346.950 553.050 349.050 ;
        RECT 557.400 348.450 558.450 349.950 ;
        RECT 554.400 347.400 558.450 348.450 ;
        RECT 545.400 346.050 546.450 346.950 ;
        RECT 544.950 343.950 547.050 346.050 ;
        RECT 545.400 343.050 546.450 343.950 ;
        RECT 551.400 343.050 552.450 346.950 ;
        RECT 538.950 340.950 541.050 343.050 ;
        RECT 544.950 340.950 547.050 343.050 ;
        RECT 548.250 341.250 550.050 342.150 ;
        RECT 550.950 340.950 553.050 343.050 ;
        RECT 554.400 342.450 555.450 347.400 ;
        RECT 556.950 344.250 559.050 345.150 ;
        RECT 563.400 343.050 564.450 352.950 ;
        RECT 556.950 342.450 559.050 343.050 ;
        RECT 554.400 341.400 559.050 342.450 ;
        RECT 556.950 340.950 559.050 341.400 ;
        RECT 560.250 341.250 561.750 342.150 ;
        RECT 562.950 340.950 565.050 343.050 ;
        RECT 566.250 341.250 568.050 342.150 ;
        RECT 538.950 338.850 541.050 339.750 ;
        RECT 541.950 338.250 544.050 339.150 ;
        RECT 544.950 338.850 546.750 339.750 ;
        RECT 547.950 337.950 550.050 340.050 ;
        RECT 553.950 337.950 556.050 340.050 ;
        RECT 559.950 337.950 562.050 340.050 ;
        RECT 563.250 338.850 564.750 339.750 ;
        RECT 565.950 337.950 568.050 340.050 ;
        RECT 541.950 334.950 544.050 337.050 ;
        RECT 542.400 331.050 543.450 334.950 ;
        RECT 541.950 328.950 544.050 331.050 ;
        RECT 544.950 328.950 547.050 331.050 ;
        RECT 535.950 322.950 538.050 325.050 ;
        RECT 535.950 319.950 538.050 322.050 ;
        RECT 541.950 319.950 544.050 322.050 ;
        RECT 536.400 313.050 537.450 319.950 ;
        RECT 542.400 316.050 543.450 319.950 ;
        RECT 545.400 319.050 546.450 328.950 ;
        RECT 548.400 319.050 549.450 337.950 ;
        RECT 544.950 316.950 547.050 319.050 ;
        RECT 547.950 316.950 550.050 319.050 ;
        RECT 541.950 313.950 544.050 316.050 ;
        RECT 547.950 313.950 550.050 316.050 ;
        RECT 535.950 310.950 538.050 313.050 ;
        RECT 539.250 311.250 541.050 312.150 ;
        RECT 541.950 311.850 544.050 312.750 ;
        RECT 544.950 311.250 547.050 312.150 ;
        RECT 535.950 308.850 537.750 309.750 ;
        RECT 538.950 307.950 541.050 310.050 ;
        RECT 544.950 307.950 547.050 310.050 ;
        RECT 539.400 307.050 540.450 307.950 ;
        RECT 538.950 304.950 541.050 307.050 ;
        RECT 545.400 301.050 546.450 307.950 ;
        RECT 548.400 307.050 549.450 313.950 ;
        RECT 554.400 310.050 555.450 337.950 ;
        RECT 560.400 337.050 561.450 337.950 ;
        RECT 559.950 334.950 562.050 337.050 ;
        RECT 569.400 334.050 570.450 370.950 ;
        RECT 572.400 358.050 573.450 374.400 ;
        RECT 577.950 367.950 580.050 370.050 ;
        RECT 571.950 355.950 574.050 358.050 ;
        RECT 571.950 352.950 574.050 355.050 ;
        RECT 572.400 340.050 573.450 352.950 ;
        RECT 574.950 343.950 577.050 346.050 ;
        RECT 575.400 342.900 576.450 343.950 ;
        RECT 574.950 340.800 577.050 342.900 ;
        RECT 571.950 337.950 574.050 340.050 ;
        RECT 574.950 338.700 577.050 339.600 ;
        RECT 568.950 331.950 571.050 334.050 ;
        RECT 572.400 331.050 573.450 337.950 ;
        RECT 578.400 337.050 579.450 367.950 ;
        RECT 584.400 346.050 585.450 388.950 ;
        RECT 587.400 385.050 588.450 391.950 ;
        RECT 590.400 391.050 591.450 418.950 ;
        RECT 592.950 416.250 595.050 417.150 ;
        RECT 608.400 415.050 609.450 436.950 ;
        RECT 614.400 424.050 615.450 451.950 ;
        RECT 617.400 448.050 618.450 451.950 ;
        RECT 620.400 451.050 621.450 461.400 ;
        RECT 626.400 460.050 627.450 496.950 ;
        RECT 628.950 487.950 631.050 490.050 ;
        RECT 646.950 488.250 649.050 489.150 ;
        RECT 629.400 487.050 630.450 487.950 ;
        RECT 628.950 484.950 631.050 487.050 ;
        RECT 634.950 484.950 637.050 487.050 ;
        RECT 637.950 485.250 639.750 486.150 ;
        RECT 640.950 484.950 643.050 487.050 ;
        RECT 646.950 486.450 649.050 487.050 ;
        RECT 650.400 486.450 651.450 523.950 ;
        RECT 652.950 520.950 655.050 523.050 ;
        RECT 656.250 521.850 657.750 522.750 ;
        RECT 658.950 520.950 661.050 523.050 ;
        RECT 653.400 520.050 654.450 520.950 ;
        RECT 652.950 517.950 655.050 520.050 ;
        RECT 652.950 508.950 655.050 511.050 ;
        RECT 644.250 485.250 645.750 486.150 ;
        RECT 646.950 485.400 651.450 486.450 ;
        RECT 646.950 484.950 649.050 485.400 ;
        RECT 628.950 482.850 631.050 483.750 ;
        RECT 631.950 482.250 634.050 483.150 ;
        RECT 631.950 478.950 634.050 481.050 ;
        RECT 628.950 472.950 631.050 475.050 ;
        RECT 629.400 466.050 630.450 472.950 ;
        RECT 635.400 469.050 636.450 484.950 ;
        RECT 637.950 481.950 640.050 484.050 ;
        RECT 641.250 482.850 642.750 483.750 ;
        RECT 643.950 481.950 646.050 484.050 ;
        RECT 644.400 472.050 645.450 481.950 ;
        RECT 650.400 481.050 651.450 485.400 ;
        RECT 649.950 478.950 652.050 481.050 ;
        RECT 653.400 472.050 654.450 508.950 ;
        RECT 659.400 490.050 660.450 520.950 ;
        RECT 662.400 520.050 663.450 556.950 ;
        RECT 664.950 553.950 667.050 556.050 ;
        RECT 668.250 554.250 669.750 555.150 ;
        RECT 670.950 553.950 673.050 556.050 ;
        RECT 664.950 550.950 667.050 553.050 ;
        RECT 667.950 550.950 670.050 553.050 ;
        RECT 665.400 529.050 666.450 550.950 ;
        RECT 668.400 547.050 669.450 550.950 ;
        RECT 671.400 550.050 672.450 553.950 ;
        RECT 670.950 547.950 673.050 550.050 ;
        RECT 667.950 544.950 670.050 547.050 ;
        RECT 664.950 526.950 667.050 529.050 ;
        RECT 674.400 526.050 675.450 580.950 ;
        RECT 677.400 577.050 678.450 595.950 ;
        RECT 682.950 593.850 685.050 594.750 ;
        RECT 676.950 574.950 679.050 577.050 ;
        RECT 686.400 568.050 687.450 622.950 ;
        RECT 695.400 613.050 696.450 625.950 ;
        RECT 701.400 616.050 702.450 625.950 ;
        RECT 707.400 616.050 708.450 625.950 ;
        RECT 709.950 622.950 712.050 625.050 ;
        RECT 700.950 613.950 703.050 616.050 ;
        RECT 706.950 613.950 709.050 616.050 ;
        RECT 694.950 610.950 697.050 613.050 ;
        RECT 700.950 610.950 703.050 613.050 ;
        RECT 701.400 604.050 702.450 610.950 ;
        RECT 710.400 610.050 711.450 622.950 ;
        RECT 716.400 619.050 717.450 631.950 ;
        RECT 715.950 616.950 718.050 619.050 ;
        RECT 709.950 607.950 712.050 610.050 ;
        RECT 688.950 601.950 691.050 604.050 ;
        RECT 700.950 601.950 703.050 604.050 ;
        RECT 689.400 595.050 690.450 601.950 ;
        RECT 716.400 601.050 717.450 616.950 ;
        RECT 691.950 599.250 694.050 600.150 ;
        RECT 694.950 599.850 697.050 600.750 ;
        RECT 701.250 599.850 702.750 600.750 ;
        RECT 703.950 598.950 706.050 601.050 ;
        RECT 709.950 599.850 712.050 600.750 ;
        RECT 712.950 599.250 715.050 600.150 ;
        RECT 715.950 598.950 718.050 601.050 ;
        RECT 691.950 595.950 694.050 598.050 ;
        RECT 697.950 596.850 700.050 597.750 ;
        RECT 703.950 596.850 706.050 597.750 ;
        RECT 706.950 595.950 709.050 598.050 ;
        RECT 712.950 595.950 715.050 598.050 ;
        RECT 688.950 592.950 691.050 595.050 ;
        RECT 692.400 570.450 693.450 595.950 ;
        RECT 697.950 592.950 700.050 595.050 ;
        RECT 698.400 571.050 699.450 592.950 ;
        RECT 689.400 569.400 693.450 570.450 ;
        RECT 685.950 565.950 688.050 568.050 ;
        RECT 689.400 561.450 690.450 569.400 ;
        RECT 697.950 568.950 700.050 571.050 ;
        RECT 691.950 565.950 694.050 568.050 ;
        RECT 686.400 560.400 690.450 561.450 ;
        RECT 686.400 559.050 687.450 560.400 ;
        RECT 676.950 557.250 678.750 558.150 ;
        RECT 679.950 556.950 682.050 559.050 ;
        RECT 683.250 557.250 684.750 558.150 ;
        RECT 685.950 556.950 688.050 559.050 ;
        RECT 689.250 557.250 691.050 558.150 ;
        RECT 676.950 553.950 679.050 556.050 ;
        RECT 680.250 554.850 681.750 555.750 ;
        RECT 682.950 553.950 685.050 556.050 ;
        RECT 686.250 554.850 687.750 555.750 ;
        RECT 688.950 553.950 691.050 556.050 ;
        RECT 677.400 544.050 678.450 553.950 ;
        RECT 683.400 552.450 684.450 553.950 ;
        RECT 692.400 553.050 693.450 565.950 ;
        RECT 698.400 559.050 699.450 568.950 ;
        RECT 707.400 568.050 708.450 595.950 ;
        RECT 709.950 586.950 712.050 589.050 ;
        RECT 700.950 565.950 703.050 568.050 ;
        RECT 706.950 565.950 709.050 568.050 ;
        RECT 701.400 562.050 702.450 565.950 ;
        RECT 710.400 564.450 711.450 586.950 ;
        RECT 713.400 568.050 714.450 595.950 ;
        RECT 712.950 565.950 715.050 568.050 ;
        RECT 719.400 565.050 720.450 661.950 ;
        RECT 722.400 655.050 723.450 667.950 ;
        RECT 727.950 664.950 730.050 667.050 ;
        RECT 730.950 664.950 733.050 667.050 ;
        RECT 734.250 665.850 735.750 666.750 ;
        RECT 736.950 664.950 739.050 667.050 ;
        RECT 740.250 665.850 742.050 666.750 ;
        RECT 742.950 664.950 745.050 667.050 ;
        RECT 721.950 652.950 724.050 655.050 ;
        RECT 724.950 637.950 727.050 640.050 ;
        RECT 725.400 637.050 726.450 637.950 ;
        RECT 724.950 634.950 727.050 637.050 ;
        RECT 725.400 631.050 726.450 634.950 ;
        RECT 728.400 634.050 729.450 664.950 ;
        RECT 731.400 652.050 732.450 664.950 ;
        RECT 736.950 662.850 739.050 663.750 ;
        RECT 730.950 649.950 733.050 652.050 ;
        RECT 736.950 646.950 739.050 649.050 ;
        RECT 727.950 631.950 730.050 634.050 ;
        RECT 721.950 629.250 723.750 630.150 ;
        RECT 724.950 628.950 727.050 631.050 ;
        RECT 728.250 629.250 729.750 630.150 ;
        RECT 730.950 628.950 733.050 631.050 ;
        RECT 734.250 629.250 736.050 630.150 ;
        RECT 721.950 625.950 724.050 628.050 ;
        RECT 725.250 626.850 726.750 627.750 ;
        RECT 727.950 625.950 730.050 628.050 ;
        RECT 731.250 626.850 732.750 627.750 ;
        RECT 733.950 625.950 736.050 628.050 ;
        RECT 724.950 622.950 727.050 625.050 ;
        RECT 725.400 616.050 726.450 622.950 ;
        RECT 724.950 613.950 727.050 616.050 ;
        RECT 725.400 604.050 726.450 613.950 ;
        RECT 728.400 604.050 729.450 625.950 ;
        RECT 737.400 607.050 738.450 646.950 ;
        RECT 743.400 643.050 744.450 664.950 ;
        RECT 749.400 646.050 750.450 667.950 ;
        RECT 748.950 643.950 751.050 646.050 ;
        RECT 742.950 640.950 745.050 643.050 ;
        RECT 752.400 636.450 753.450 670.950 ;
        RECT 757.950 669.450 760.050 670.050 ;
        RECT 761.400 669.450 762.450 679.950 ;
        RECT 757.950 668.400 762.450 669.450 ;
        RECT 757.950 667.950 760.050 668.400 ;
        RECT 766.950 667.950 769.050 670.050 ;
        RECT 749.400 635.400 753.450 636.450 ;
        RECT 742.950 628.950 745.050 631.050 ;
        RECT 745.950 628.950 748.050 631.050 ;
        RECT 739.950 626.250 742.050 627.150 ;
        RECT 742.950 626.850 745.050 627.750 ;
        RECT 739.950 622.950 742.050 625.050 ;
        RECT 740.400 622.050 741.450 622.950 ;
        RECT 739.950 619.950 742.050 622.050 ;
        RECT 730.950 604.950 733.050 607.050 ;
        RECT 736.950 604.950 739.050 607.050 ;
        RECT 724.950 601.950 727.050 604.050 ;
        RECT 727.950 601.950 730.050 604.050 ;
        RECT 725.250 599.850 726.750 600.750 ;
        RECT 727.950 598.950 730.050 601.050 ;
        RECT 721.950 596.850 724.050 597.750 ;
        RECT 724.950 595.950 727.050 598.050 ;
        RECT 727.950 596.850 730.050 597.750 ;
        RECT 707.400 563.400 711.450 564.450 ;
        RECT 700.950 559.950 703.050 562.050 ;
        RECT 703.950 560.250 706.050 561.150 ;
        RECT 694.950 557.250 696.750 558.150 ;
        RECT 697.950 556.950 700.050 559.050 ;
        RECT 701.250 557.250 702.750 558.150 ;
        RECT 703.950 556.950 706.050 559.050 ;
        RECT 704.400 556.050 705.450 556.950 ;
        RECT 694.950 553.950 697.050 556.050 ;
        RECT 698.250 554.850 699.750 555.750 ;
        RECT 700.950 553.950 703.050 556.050 ;
        RECT 703.950 553.950 706.050 556.050 ;
        RECT 685.950 552.450 688.050 553.050 ;
        RECT 683.400 551.400 688.050 552.450 ;
        RECT 685.950 550.950 688.050 551.400 ;
        RECT 691.950 550.950 694.050 553.050 ;
        RECT 695.400 550.050 696.450 553.950 ;
        RECT 697.950 550.950 700.050 553.050 ;
        RECT 682.950 547.950 685.050 550.050 ;
        RECT 694.950 547.950 697.050 550.050 ;
        RECT 676.950 541.950 679.050 544.050 ;
        RECT 664.950 524.250 666.750 525.150 ;
        RECT 667.950 523.950 670.050 526.050 ;
        RECT 671.250 524.250 673.050 525.150 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 664.950 520.950 667.050 523.050 ;
        RECT 668.250 521.850 669.750 522.750 ;
        RECT 670.950 520.950 673.050 523.050 ;
        RECT 661.950 517.950 664.050 520.050 ;
        RECT 662.400 496.050 663.450 517.950 ;
        RECT 665.400 517.050 666.450 520.950 ;
        RECT 664.950 514.950 667.050 517.050 ;
        RECT 671.400 511.050 672.450 520.950 ;
        RECT 670.950 508.950 673.050 511.050 ;
        RECT 677.400 502.050 678.450 541.950 ;
        RECT 679.950 527.250 682.050 528.150 ;
        RECT 679.950 523.950 682.050 526.050 ;
        RECT 679.950 520.950 682.050 523.050 ;
        RECT 676.950 499.950 679.050 502.050 ;
        RECT 661.950 493.950 664.050 496.050 ;
        RECT 658.950 487.950 661.050 490.050 ;
        RECT 655.950 485.250 657.750 486.150 ;
        RECT 658.950 484.950 661.050 487.050 ;
        RECT 662.250 485.250 663.750 486.150 ;
        RECT 664.950 484.950 667.050 487.050 ;
        RECT 668.250 485.250 670.050 486.150 ;
        RECT 670.950 485.250 673.050 486.150 ;
        RECT 676.950 485.250 679.050 486.150 ;
        RECT 655.950 481.950 658.050 484.050 ;
        RECT 659.250 482.850 660.750 483.750 ;
        RECT 661.950 481.950 664.050 484.050 ;
        RECT 665.250 482.850 666.750 483.750 ;
        RECT 667.950 483.450 670.050 484.050 ;
        RECT 670.950 483.450 673.050 484.050 ;
        RECT 667.950 482.400 673.050 483.450 ;
        RECT 667.950 481.950 670.050 482.400 ;
        RECT 670.950 481.950 673.050 482.400 ;
        RECT 674.250 482.250 675.750 483.150 ;
        RECT 676.950 481.950 679.050 484.050 ;
        RECT 656.400 481.050 657.450 481.950 ;
        RECT 655.950 478.950 658.050 481.050 ;
        RECT 658.950 478.950 661.050 481.050 ;
        RECT 643.950 469.950 646.050 472.050 ;
        RECT 652.950 469.950 655.050 472.050 ;
        RECT 634.950 466.950 637.050 469.050 ;
        RECT 628.950 463.950 631.050 466.050 ;
        RECT 643.950 463.950 646.050 466.050 ;
        RECT 622.950 457.950 625.050 460.050 ;
        RECT 625.950 457.950 628.050 460.050 ;
        RECT 637.950 457.950 640.050 460.050 ;
        RECT 623.400 457.050 624.450 457.950 ;
        RECT 622.950 454.950 625.050 457.050 ;
        RECT 626.250 455.250 627.750 456.150 ;
        RECT 628.950 454.950 631.050 457.050 ;
        RECT 632.250 455.250 633.750 456.150 ;
        RECT 634.950 454.950 637.050 457.050 ;
        RECT 622.950 452.850 624.750 453.750 ;
        RECT 625.950 451.950 628.050 454.050 ;
        RECT 629.250 452.850 630.750 453.750 ;
        RECT 631.950 451.950 634.050 454.050 ;
        RECT 635.250 452.850 637.050 453.750 ;
        RECT 626.400 451.050 627.450 451.950 ;
        RECT 619.950 448.950 622.050 451.050 ;
        RECT 625.950 448.950 628.050 451.050 ;
        RECT 616.950 445.950 619.050 448.050 ;
        RECT 619.950 442.950 622.050 445.050 ;
        RECT 620.400 436.050 621.450 442.950 ;
        RECT 619.950 433.950 622.050 436.050 ;
        RECT 622.950 433.950 625.050 436.050 ;
        RECT 613.950 421.950 616.050 424.050 ;
        RECT 616.950 421.950 619.050 424.050 ;
        RECT 613.950 416.250 616.050 417.150 ;
        RECT 617.400 415.050 618.450 421.950 ;
        RECT 623.400 418.050 624.450 433.950 ;
        RECT 626.400 421.050 627.450 448.950 ;
        RECT 632.400 433.050 633.450 451.950 ;
        RECT 631.950 430.950 634.050 433.050 ;
        RECT 638.400 432.450 639.450 457.950 ;
        RECT 644.400 454.050 645.450 463.950 ;
        RECT 659.400 460.050 660.450 478.950 ;
        RECT 662.400 475.050 663.450 481.950 ;
        RECT 668.400 475.050 669.450 481.950 ;
        RECT 673.950 478.950 676.050 481.050 ;
        RECT 676.950 478.950 679.050 481.050 ;
        RECT 661.950 472.950 664.050 475.050 ;
        RECT 667.950 472.950 670.050 475.050 ;
        RECT 674.400 474.450 675.450 478.950 ;
        RECT 671.400 473.400 675.450 474.450 ;
        RECT 649.950 459.450 652.050 460.050 ;
        RECT 647.400 458.400 652.050 459.450 ;
        RECT 647.400 457.050 648.450 458.400 ;
        RECT 649.950 457.950 652.050 458.400 ;
        RECT 658.950 457.950 661.050 460.050 ;
        RECT 664.950 457.950 667.050 460.050 ;
        RECT 665.400 457.050 666.450 457.950 ;
        RECT 646.950 454.950 649.050 457.050 ;
        RECT 649.950 455.850 652.050 456.750 ;
        RECT 658.950 456.450 661.050 457.050 ;
        RECT 652.950 455.250 655.050 456.150 ;
        RECT 656.400 455.400 661.050 456.450 ;
        RECT 640.950 452.250 642.750 453.150 ;
        RECT 643.950 451.950 646.050 454.050 ;
        RECT 647.250 452.250 649.050 453.150 ;
        RECT 649.950 451.950 652.050 454.050 ;
        RECT 652.950 453.450 655.050 454.050 ;
        RECT 656.400 453.450 657.450 455.400 ;
        RECT 658.950 454.950 661.050 455.400 ;
        RECT 662.250 455.250 663.750 456.150 ;
        RECT 664.950 454.950 667.050 457.050 ;
        RECT 668.400 454.050 669.450 472.950 ;
        RECT 671.400 469.050 672.450 473.400 ;
        RECT 673.950 469.950 676.050 472.050 ;
        RECT 670.950 466.950 673.050 469.050 ;
        RECT 670.950 454.950 673.050 457.050 ;
        RECT 652.950 452.400 657.450 453.450 ;
        RECT 658.950 452.850 660.750 453.750 ;
        RECT 652.950 451.950 655.050 452.400 ;
        RECT 661.950 451.950 664.050 454.050 ;
        RECT 665.250 452.850 666.750 453.750 ;
        RECT 667.950 451.950 670.050 454.050 ;
        RECT 640.950 448.950 643.050 451.050 ;
        RECT 644.250 449.850 645.750 450.750 ;
        RECT 646.950 448.950 649.050 451.050 ;
        RECT 647.400 445.050 648.450 448.950 ;
        RECT 646.950 442.950 649.050 445.050 ;
        RECT 650.400 436.050 651.450 451.950 ;
        RECT 662.400 442.050 663.450 451.950 ;
        RECT 664.950 448.950 667.050 451.050 ;
        RECT 667.950 449.850 670.050 450.750 ;
        RECT 665.400 442.050 666.450 448.950 ;
        RECT 671.400 447.450 672.450 454.950 ;
        RECT 674.400 451.050 675.450 469.950 ;
        RECT 677.400 463.050 678.450 478.950 ;
        RECT 680.400 475.050 681.450 520.950 ;
        RECT 683.400 493.050 684.450 547.950 ;
        RECT 691.950 544.950 694.050 547.050 ;
        RECT 682.950 490.950 685.050 493.050 ;
        RECT 688.950 490.950 691.050 493.050 ;
        RECT 689.400 490.050 690.450 490.950 ;
        RECT 682.950 487.950 685.050 490.050 ;
        RECT 686.250 488.250 687.750 489.150 ;
        RECT 688.950 487.950 691.050 490.050 ;
        RECT 682.950 485.850 684.750 486.750 ;
        RECT 685.950 484.950 688.050 487.050 ;
        RECT 689.250 485.850 691.050 486.750 ;
        RECT 692.400 483.450 693.450 544.950 ;
        RECT 694.950 538.950 697.050 541.050 ;
        RECT 695.400 529.050 696.450 538.950 ;
        RECT 698.400 538.050 699.450 550.950 ;
        RECT 697.950 535.950 700.050 538.050 ;
        RECT 697.950 532.950 700.050 535.050 ;
        RECT 694.950 526.950 697.050 529.050 ;
        RECT 698.400 492.450 699.450 532.950 ;
        RECT 703.950 529.950 706.050 532.050 ;
        RECT 700.950 527.250 703.050 528.150 ;
        RECT 704.400 520.050 705.450 529.950 ;
        RECT 703.950 517.950 706.050 520.050 ;
        RECT 695.400 491.400 699.450 492.450 ;
        RECT 695.400 487.050 696.450 491.400 ;
        RECT 707.400 490.050 708.450 563.400 ;
        RECT 712.950 563.250 715.050 564.150 ;
        RECT 718.950 562.950 721.050 565.050 ;
        RECT 709.950 560.250 711.750 561.150 ;
        RECT 712.950 559.950 715.050 562.050 ;
        RECT 716.250 560.250 717.750 561.150 ;
        RECT 718.950 559.950 721.050 562.050 ;
        RECT 725.400 561.450 726.450 595.950 ;
        RECT 731.400 583.050 732.450 604.950 ;
        RECT 739.950 601.950 742.050 604.050 ;
        RECT 740.400 601.050 741.450 601.950 ;
        RECT 733.950 598.950 736.050 601.050 ;
        RECT 737.250 599.250 738.750 600.150 ;
        RECT 739.950 598.950 742.050 601.050 ;
        RECT 746.400 598.050 747.450 628.950 ;
        RECT 749.400 604.050 750.450 635.400 ;
        RECT 751.950 632.250 754.050 633.150 ;
        RECT 751.950 628.950 754.050 631.050 ;
        RECT 755.250 629.250 756.750 630.150 ;
        RECT 757.950 628.950 760.050 631.050 ;
        RECT 761.250 629.250 763.050 630.150 ;
        RECT 754.950 625.950 757.050 628.050 ;
        RECT 758.250 626.850 759.750 627.750 ;
        RECT 760.950 627.450 763.050 628.050 ;
        RECT 760.950 626.400 765.450 627.450 ;
        RECT 760.950 625.950 763.050 626.400 ;
        RECT 755.400 607.050 756.450 625.950 ;
        RECT 757.950 622.950 760.050 625.050 ;
        RECT 760.950 622.950 763.050 625.050 ;
        RECT 754.950 604.950 757.050 607.050 ;
        RECT 748.950 601.950 751.050 604.050 ;
        RECT 751.950 601.950 754.050 604.050 ;
        RECT 758.400 601.050 759.450 622.950 ;
        RECT 748.950 599.250 751.050 600.150 ;
        RECT 751.950 599.850 754.050 600.750 ;
        RECT 754.950 599.250 756.750 600.150 ;
        RECT 757.950 598.950 760.050 601.050 ;
        RECT 733.950 596.850 735.750 597.750 ;
        RECT 736.950 595.950 739.050 598.050 ;
        RECT 740.250 596.850 741.750 597.750 ;
        RECT 742.950 595.950 745.050 598.050 ;
        RECT 745.950 595.950 748.050 598.050 ;
        RECT 748.950 595.950 751.050 598.050 ;
        RECT 751.950 595.950 754.050 598.050 ;
        RECT 754.950 595.950 757.050 598.050 ;
        RECT 758.250 596.850 760.050 597.750 ;
        RECT 737.400 592.050 738.450 595.950 ;
        RECT 739.950 592.950 742.050 595.050 ;
        RECT 742.950 593.850 745.050 594.750 ;
        RECT 736.950 589.950 739.050 592.050 ;
        RECT 730.950 580.950 733.050 583.050 ;
        RECT 730.950 577.950 733.050 580.050 ;
        RECT 722.400 560.400 726.450 561.450 ;
        RECT 709.950 556.950 712.050 559.050 ;
        RECT 709.950 553.950 712.050 556.050 ;
        RECT 710.400 532.050 711.450 553.950 ;
        RECT 713.400 550.050 714.450 559.950 ;
        RECT 715.950 556.950 718.050 559.050 ;
        RECT 719.250 557.850 721.050 558.750 ;
        RECT 712.950 547.950 715.050 550.050 ;
        RECT 709.950 529.950 712.050 532.050 ;
        RECT 712.950 531.450 715.050 532.050 ;
        RECT 716.400 531.450 717.450 556.950 ;
        RECT 722.400 550.050 723.450 560.400 ;
        RECT 731.400 559.050 732.450 577.950 ;
        RECT 736.950 568.950 739.050 571.050 ;
        RECT 727.950 558.450 730.050 559.050 ;
        RECT 725.400 557.400 730.050 558.450 ;
        RECT 721.950 547.950 724.050 550.050 ;
        RECT 725.400 544.050 726.450 557.400 ;
        RECT 727.950 556.950 730.050 557.400 ;
        RECT 730.950 556.950 733.050 559.050 ;
        RECT 733.950 556.950 736.050 559.050 ;
        RECT 727.950 554.850 730.050 555.750 ;
        RECT 733.950 554.850 736.050 555.750 ;
        RECT 721.950 541.950 724.050 544.050 ;
        RECT 724.950 541.950 727.050 544.050 ;
        RECT 718.950 531.450 721.050 532.050 ;
        RECT 712.950 530.400 721.050 531.450 ;
        RECT 712.950 529.950 715.050 530.400 ;
        RECT 718.950 529.950 721.050 530.400 ;
        RECT 722.400 529.050 723.450 541.950 ;
        RECT 730.950 529.950 733.050 532.050 ;
        RECT 709.950 527.250 712.050 528.150 ;
        RECT 712.950 527.850 715.050 528.750 ;
        RECT 715.950 526.950 718.050 529.050 ;
        RECT 719.250 527.850 720.750 528.750 ;
        RECT 721.950 526.950 724.050 529.050 ;
        RECT 724.950 526.950 727.050 529.050 ;
        RECT 709.950 523.950 712.050 526.050 ;
        RECT 715.950 524.850 718.050 525.750 ;
        RECT 721.950 524.850 724.050 525.750 ;
        RECT 710.400 514.050 711.450 523.950 ;
        RECT 721.950 520.950 724.050 523.050 ;
        RECT 725.400 522.450 726.450 526.950 ;
        RECT 731.400 526.050 732.450 529.950 ;
        RECT 737.400 526.050 738.450 568.950 ;
        RECT 740.400 562.050 741.450 592.950 ;
        RECT 749.400 589.050 750.450 595.950 ;
        RECT 748.950 586.950 751.050 589.050 ;
        RECT 748.950 583.950 751.050 586.050 ;
        RECT 742.950 580.950 745.050 583.050 ;
        RECT 739.950 559.950 742.050 562.050 ;
        RECT 739.950 557.250 742.050 558.150 ;
        RECT 739.950 553.950 742.050 556.050 ;
        RECT 740.400 550.050 741.450 553.950 ;
        RECT 739.950 547.950 742.050 550.050 ;
        RECT 739.950 535.950 742.050 538.050 ;
        RECT 727.950 524.250 729.750 525.150 ;
        RECT 730.950 523.950 733.050 526.050 ;
        RECT 734.250 524.250 736.050 525.150 ;
        RECT 736.950 523.950 739.050 526.050 ;
        RECT 727.950 522.450 730.050 523.050 ;
        RECT 725.400 521.400 730.050 522.450 ;
        RECT 731.250 521.850 732.750 522.750 ;
        RECT 727.950 520.950 730.050 521.400 ;
        RECT 733.950 520.950 736.050 523.050 ;
        RECT 709.950 511.950 712.050 514.050 ;
        RECT 722.400 493.050 723.450 520.950 ;
        RECT 734.400 520.050 735.450 520.950 ;
        RECT 733.950 517.950 736.050 520.050 ;
        RECT 733.950 514.950 736.050 517.050 ;
        RECT 724.950 511.950 727.050 514.050 ;
        RECT 712.950 490.950 715.050 493.050 ;
        RECT 721.950 490.950 724.050 493.050 ;
        RECT 697.950 488.250 700.050 489.150 ;
        RECT 706.950 487.950 709.050 490.050 ;
        RECT 713.400 487.050 714.450 490.950 ;
        RECT 725.400 489.450 726.450 511.950 ;
        RECT 718.950 488.250 721.050 489.150 ;
        RECT 722.400 488.400 726.450 489.450 ;
        RECT 694.950 484.950 697.050 487.050 ;
        RECT 697.950 484.950 700.050 487.050 ;
        RECT 701.250 485.250 702.750 486.150 ;
        RECT 703.950 484.950 706.050 487.050 ;
        RECT 707.250 485.250 709.050 486.150 ;
        RECT 709.950 485.250 711.750 486.150 ;
        RECT 712.950 484.950 715.050 487.050 ;
        RECT 716.250 485.250 717.750 486.150 ;
        RECT 718.950 484.950 721.050 487.050 ;
        RECT 689.400 482.400 693.450 483.450 ;
        RECT 682.950 475.950 685.050 478.050 ;
        RECT 679.950 472.950 682.050 475.050 ;
        RECT 679.950 466.950 682.050 469.050 ;
        RECT 676.950 460.950 679.050 463.050 ;
        RECT 680.400 457.050 681.450 466.950 ;
        RECT 683.400 463.050 684.450 475.950 ;
        RECT 689.400 475.050 690.450 482.400 ;
        RECT 694.950 481.950 697.050 484.050 ;
        RECT 691.950 478.950 694.050 481.050 ;
        RECT 688.950 472.950 691.050 475.050 ;
        RECT 688.950 469.950 691.050 472.050 ;
        RECT 682.950 460.950 685.050 463.050 ;
        RECT 685.950 460.950 688.050 463.050 ;
        RECT 686.400 460.050 687.450 460.950 ;
        RECT 685.950 457.950 688.050 460.050 ;
        RECT 679.950 454.950 682.050 457.050 ;
        RECT 686.400 454.050 687.450 457.950 ;
        RECT 676.950 452.250 678.750 453.150 ;
        RECT 679.950 451.950 682.050 454.050 ;
        RECT 682.950 451.950 685.050 454.050 ;
        RECT 685.950 451.950 688.050 454.050 ;
        RECT 683.400 451.050 684.450 451.950 ;
        RECT 673.950 448.950 676.050 451.050 ;
        RECT 676.950 448.950 679.050 451.050 ;
        RECT 680.250 449.850 681.750 450.750 ;
        RECT 682.950 448.950 685.050 451.050 ;
        RECT 686.250 449.850 688.050 450.750 ;
        RECT 677.400 448.050 678.450 448.950 ;
        RECT 668.400 446.400 672.450 447.450 ;
        RECT 661.950 439.950 664.050 442.050 ;
        RECT 664.950 439.950 667.050 442.050 ;
        RECT 668.400 438.450 669.450 446.400 ;
        RECT 673.950 445.950 676.050 448.050 ;
        RECT 676.950 445.950 679.050 448.050 ;
        RECT 682.950 446.850 685.050 447.750 ;
        RECT 670.950 442.950 673.050 445.050 ;
        RECT 665.400 437.400 669.450 438.450 ;
        RECT 643.950 433.950 646.050 436.050 ;
        RECT 649.950 433.950 652.050 436.050 ;
        RECT 638.400 431.400 642.450 432.450 ;
        RECT 637.950 427.950 640.050 430.050 ;
        RECT 638.400 424.050 639.450 427.950 ;
        RECT 637.950 421.950 640.050 424.050 ;
        RECT 625.950 418.950 628.050 421.050 ;
        RECT 628.950 419.250 631.050 420.150 ;
        RECT 622.950 417.450 625.050 418.050 ;
        RECT 620.400 416.400 625.050 417.450 ;
        RECT 592.950 412.950 595.050 415.050 ;
        RECT 596.250 413.250 597.750 414.150 ;
        RECT 598.950 412.950 601.050 415.050 ;
        RECT 602.250 413.250 604.050 414.150 ;
        RECT 604.950 413.250 606.750 414.150 ;
        RECT 607.950 412.950 610.050 415.050 ;
        RECT 613.950 414.450 616.050 415.050 ;
        RECT 616.950 414.450 619.050 415.050 ;
        RECT 611.250 413.250 612.750 414.150 ;
        RECT 613.950 413.400 619.050 414.450 ;
        RECT 613.950 412.950 616.050 413.400 ;
        RECT 616.950 412.950 619.050 413.400 ;
        RECT 593.400 412.050 594.450 412.950 ;
        RECT 592.950 409.950 595.050 412.050 ;
        RECT 595.950 409.950 598.050 412.050 ;
        RECT 599.250 410.850 600.750 411.750 ;
        RECT 601.950 409.950 604.050 412.050 ;
        RECT 604.950 409.950 607.050 412.050 ;
        RECT 608.250 410.850 609.750 411.750 ;
        RECT 610.950 409.950 613.050 412.050 ;
        RECT 616.950 409.950 619.050 412.050 ;
        RECT 593.400 408.450 594.450 409.950 ;
        RECT 605.400 408.450 606.450 409.950 ;
        RECT 593.400 407.400 606.450 408.450 ;
        RECT 598.950 394.950 601.050 397.050 ;
        RECT 589.950 388.950 592.050 391.050 ;
        RECT 592.950 385.950 595.050 388.050 ;
        RECT 599.400 387.450 600.450 394.950 ;
        RECT 604.950 388.950 607.050 391.050 ;
        RECT 601.950 387.450 604.050 388.050 ;
        RECT 599.400 386.400 604.050 387.450 ;
        RECT 605.400 387.450 606.450 388.950 ;
        RECT 605.400 386.400 609.450 387.450 ;
        RECT 593.400 385.050 594.450 385.950 ;
        RECT 599.400 385.050 600.450 386.400 ;
        RECT 601.950 385.950 604.050 386.400 ;
        RECT 586.950 382.950 589.050 385.050 ;
        RECT 590.250 383.250 591.750 384.150 ;
        RECT 592.950 382.950 595.050 385.050 ;
        RECT 598.950 382.950 601.050 385.050 ;
        RECT 601.950 383.850 604.050 384.750 ;
        RECT 604.950 383.250 607.050 384.150 ;
        RECT 586.950 380.850 588.750 381.750 ;
        RECT 589.950 379.950 592.050 382.050 ;
        RECT 593.250 380.850 594.750 381.750 ;
        RECT 595.950 379.950 598.050 382.050 ;
        RECT 590.400 364.050 591.450 379.950 ;
        RECT 595.950 377.850 598.050 378.750 ;
        RECT 589.950 361.950 592.050 364.050 ;
        RECT 595.950 355.950 598.050 358.050 ;
        RECT 592.950 352.950 595.050 355.050 ;
        RECT 586.950 349.950 589.050 352.050 ;
        RECT 583.950 343.950 586.050 346.050 ;
        RECT 580.950 341.100 582.750 342.000 ;
        RECT 583.950 340.800 586.050 343.050 ;
        RECT 580.950 337.800 583.050 340.050 ;
        RECT 584.250 338.700 586.050 339.600 ;
        RECT 587.400 339.450 588.450 349.950 ;
        RECT 589.950 341.100 592.050 342.000 ;
        RECT 589.950 339.450 592.050 339.900 ;
        RECT 587.400 338.400 592.050 339.450 ;
        RECT 577.950 334.950 580.050 337.050 ;
        RECT 583.950 334.950 586.050 337.050 ;
        RECT 589.950 334.950 592.050 338.400 ;
        RECT 559.950 328.950 562.050 331.050 ;
        RECT 562.950 328.950 565.050 331.050 ;
        RECT 568.950 328.950 571.050 331.050 ;
        RECT 571.950 328.950 574.050 331.050 ;
        RECT 560.400 325.050 561.450 328.950 ;
        RECT 556.950 322.950 559.050 325.050 ;
        RECT 559.950 322.950 562.050 325.050 ;
        RECT 557.400 312.450 558.450 322.950 ;
        RECT 563.400 322.050 564.450 328.950 ;
        RECT 569.400 327.450 570.450 328.950 ;
        RECT 584.400 327.450 585.450 334.950 ;
        RECT 569.400 326.400 573.450 327.450 ;
        RECT 565.950 322.950 568.050 325.050 ;
        RECT 562.950 319.950 565.050 322.050 ;
        RECT 557.400 311.400 561.450 312.450 ;
        RECT 550.950 308.250 552.750 309.150 ;
        RECT 553.950 307.950 556.050 310.050 ;
        RECT 557.250 308.250 559.050 309.150 ;
        RECT 547.950 304.950 550.050 307.050 ;
        RECT 550.950 304.950 553.050 307.050 ;
        RECT 554.250 305.850 555.750 306.750 ;
        RECT 556.950 304.950 559.050 307.050 ;
        RECT 553.950 301.950 556.050 304.050 ;
        RECT 544.950 298.950 547.050 301.050 ;
        RECT 535.950 292.950 538.050 295.050 ;
        RECT 532.950 289.950 535.050 292.050 ;
        RECT 526.950 274.950 529.050 277.050 ;
        RECT 536.400 274.050 537.450 292.950 ;
        RECT 541.950 286.950 544.050 289.050 ;
        RECT 542.400 283.050 543.450 286.950 ;
        RECT 538.950 280.950 541.050 283.050 ;
        RECT 541.950 280.950 544.050 283.050 ;
        RECT 520.950 273.450 523.050 274.050 ;
        RECT 529.950 273.450 532.050 274.050 ;
        RECT 518.400 272.400 523.050 273.450 ;
        RECT 520.950 271.950 523.050 272.400 ;
        RECT 523.950 272.250 526.050 273.150 ;
        RECT 527.400 272.400 532.050 273.450 ;
        RECT 514.950 269.250 516.750 270.150 ;
        RECT 517.950 268.950 520.050 271.050 ;
        RECT 521.250 269.250 522.750 270.150 ;
        RECT 523.950 268.950 526.050 271.050 ;
        RECT 514.950 267.450 517.050 268.050 ;
        RECT 512.400 266.400 517.050 267.450 ;
        RECT 518.250 266.850 519.750 267.750 ;
        RECT 520.950 267.450 523.050 268.050 ;
        RECT 523.950 267.450 526.050 268.050 ;
        RECT 514.950 265.950 517.050 266.400 ;
        RECT 520.950 266.400 526.050 267.450 ;
        RECT 520.950 265.950 523.050 266.400 ;
        RECT 523.950 265.950 526.050 266.400 ;
        RECT 500.400 265.050 501.450 265.950 ;
        RECT 499.950 262.950 502.050 265.050 ;
        RECT 496.950 256.950 499.050 259.050 ;
        RECT 490.950 247.950 493.050 250.050 ;
        RECT 496.950 247.950 499.050 250.050 ;
        RECT 490.950 243.450 493.050 244.050 ;
        RECT 493.950 243.450 496.050 244.050 ;
        RECT 490.950 242.400 496.050 243.450 ;
        RECT 490.950 241.950 493.050 242.400 ;
        RECT 493.950 241.950 496.050 242.400 ;
        RECT 487.950 238.950 490.050 241.050 ;
        RECT 491.250 239.250 492.750 240.150 ;
        RECT 493.950 238.950 496.050 241.050 ;
        RECT 484.950 235.950 487.050 238.050 ;
        RECT 488.250 236.850 489.750 237.750 ;
        RECT 490.950 235.950 493.050 238.050 ;
        RECT 494.250 236.850 496.050 237.750 ;
        RECT 484.950 233.850 487.050 234.750 ;
        RECT 481.950 229.950 484.050 232.050 ;
        RECT 478.950 217.950 481.050 220.050 ;
        RECT 475.950 208.950 478.050 211.050 ;
        RECT 463.950 205.950 466.050 208.050 ;
        RECT 469.950 205.950 472.050 208.050 ;
        RECT 455.400 203.400 459.450 204.450 ;
        RECT 458.400 202.050 459.450 203.400 ;
        RECT 464.400 202.050 465.450 205.950 ;
        RECT 469.950 203.250 472.050 204.150 ;
        RECT 476.400 202.050 477.450 208.950 ;
        RECT 479.400 202.050 480.450 217.950 ;
        RECT 482.400 217.050 483.450 229.950 ;
        RECT 484.950 220.950 487.050 223.050 ;
        RECT 481.950 214.950 484.050 217.050 ;
        RECT 485.400 205.050 486.450 220.950 ;
        RECT 491.400 208.050 492.450 235.950 ;
        RECT 493.950 232.950 496.050 235.050 ;
        RECT 497.400 234.450 498.450 247.950 ;
        RECT 506.400 241.050 507.450 265.950 ;
        RECT 515.400 264.450 516.450 265.950 ;
        RECT 520.950 264.450 523.050 265.050 ;
        RECT 515.400 263.400 523.050 264.450 ;
        RECT 520.950 262.950 523.050 263.400 ;
        RECT 527.400 262.050 528.450 272.400 ;
        RECT 529.950 271.950 532.050 272.400 ;
        RECT 533.250 272.250 534.750 273.150 ;
        RECT 535.950 271.950 538.050 274.050 ;
        RECT 529.950 269.850 531.750 270.750 ;
        RECT 532.950 268.950 535.050 271.050 ;
        RECT 536.250 269.850 538.050 270.750 ;
        RECT 533.400 268.050 534.450 268.950 ;
        RECT 529.950 265.950 532.050 268.050 ;
        RECT 532.950 265.950 535.050 268.050 ;
        RECT 514.950 259.950 517.050 262.050 ;
        RECT 526.950 259.950 529.050 262.050 ;
        RECT 508.950 250.950 511.050 253.050 ;
        RECT 509.400 244.050 510.450 250.950 ;
        RECT 508.950 241.950 511.050 244.050 ;
        RECT 515.400 243.450 516.450 259.950 ;
        RECT 530.400 253.050 531.450 265.950 ;
        RECT 539.400 262.050 540.450 280.950 ;
        RECT 544.950 274.950 547.050 277.050 ;
        RECT 545.400 271.050 546.450 274.950 ;
        RECT 550.950 272.250 553.050 273.150 ;
        RECT 541.950 269.250 543.750 270.150 ;
        RECT 544.950 268.950 547.050 271.050 ;
        RECT 550.950 270.450 553.050 271.050 ;
        RECT 554.400 270.450 555.450 301.950 ;
        RECT 557.400 295.050 558.450 304.950 ;
        RECT 556.950 292.950 559.050 295.050 ;
        RECT 560.400 271.050 561.450 311.400 ;
        RECT 566.400 310.050 567.450 322.950 ;
        RECT 568.950 319.950 571.050 322.050 ;
        RECT 569.400 310.050 570.450 319.950 ;
        RECT 572.400 310.050 573.450 326.400 ;
        RECT 581.400 326.400 585.450 327.450 ;
        RECT 581.400 324.450 582.450 326.400 ;
        RECT 578.400 323.400 582.450 324.450 ;
        RECT 578.400 322.050 579.450 323.400 ;
        RECT 583.950 322.950 586.050 325.050 ;
        RECT 577.950 319.950 580.050 322.050 ;
        RECT 580.950 319.950 583.050 322.050 ;
        RECT 574.950 313.950 577.050 316.050 ;
        RECT 574.950 311.850 577.050 312.750 ;
        RECT 577.950 311.250 580.050 312.150 ;
        RECT 562.950 308.250 564.750 309.150 ;
        RECT 565.950 307.950 568.050 310.050 ;
        RECT 568.950 307.950 571.050 310.050 ;
        RECT 571.950 309.450 574.050 310.050 ;
        RECT 571.950 308.400 576.450 309.450 ;
        RECT 571.950 307.950 574.050 308.400 ;
        RECT 562.950 304.950 565.050 307.050 ;
        RECT 566.250 305.850 567.750 306.750 ;
        RECT 568.950 304.950 571.050 307.050 ;
        RECT 572.250 305.850 574.050 306.750 ;
        RECT 565.950 301.950 568.050 304.050 ;
        RECT 568.950 302.850 571.050 303.750 ;
        RECT 566.400 274.050 567.450 301.950 ;
        RECT 575.400 298.050 576.450 308.400 ;
        RECT 577.950 307.950 580.050 310.050 ;
        RECT 581.400 306.450 582.450 319.950 ;
        RECT 584.400 316.050 585.450 322.950 ;
        RECT 593.400 322.050 594.450 352.950 ;
        RECT 596.400 343.050 597.450 355.950 ;
        RECT 599.400 352.050 600.450 382.950 ;
        RECT 604.950 379.950 607.050 382.050 ;
        RECT 604.950 370.950 607.050 373.050 ;
        RECT 605.400 367.050 606.450 370.950 ;
        RECT 601.950 364.950 604.050 367.050 ;
        RECT 604.950 364.950 607.050 367.050 ;
        RECT 598.950 349.950 601.050 352.050 ;
        RECT 595.950 340.950 598.050 343.050 ;
        RECT 598.950 340.950 601.050 343.050 ;
        RECT 595.950 338.250 598.050 339.150 ;
        RECT 598.950 338.850 601.050 339.750 ;
        RECT 595.950 334.950 598.050 337.050 ;
        RECT 598.950 334.950 601.050 337.050 ;
        RECT 595.950 333.450 598.050 334.050 ;
        RECT 599.400 333.450 600.450 334.950 ;
        RECT 595.950 332.400 600.450 333.450 ;
        RECT 595.950 331.950 598.050 332.400 ;
        RECT 602.400 325.050 603.450 364.950 ;
        RECT 608.400 361.050 609.450 386.400 ;
        RECT 604.950 358.950 607.050 361.050 ;
        RECT 607.950 358.950 610.050 361.050 ;
        RECT 605.400 339.450 606.450 358.950 ;
        RECT 611.400 358.050 612.450 409.950 ;
        RECT 613.950 406.950 616.050 409.050 ;
        RECT 614.400 394.050 615.450 406.950 ;
        RECT 617.400 400.050 618.450 409.950 ;
        RECT 620.400 406.050 621.450 416.400 ;
        RECT 622.950 415.950 625.050 416.400 ;
        RECT 626.250 416.250 627.750 417.150 ;
        RECT 628.950 415.950 631.050 418.050 ;
        RECT 632.250 416.250 634.050 417.150 ;
        RECT 622.950 413.850 624.750 414.750 ;
        RECT 625.950 412.950 628.050 415.050 ;
        RECT 622.950 406.950 625.050 409.050 ;
        RECT 619.950 403.950 622.050 406.050 ;
        RECT 616.950 397.950 619.050 400.050 ;
        RECT 623.400 397.050 624.450 406.950 ;
        RECT 629.400 406.050 630.450 415.950 ;
        RECT 638.400 415.050 639.450 421.950 ;
        RECT 641.400 418.050 642.450 431.400 ;
        RECT 644.400 418.050 645.450 433.950 ;
        RECT 646.950 430.950 649.050 433.050 ;
        RECT 647.400 418.050 648.450 430.950 ;
        RECT 640.950 415.950 643.050 418.050 ;
        RECT 643.950 415.950 646.050 418.050 ;
        RECT 646.950 415.950 649.050 418.050 ;
        RECT 652.950 415.950 655.050 418.050 ;
        RECT 641.400 415.050 642.450 415.950 ;
        RECT 653.400 415.050 654.450 415.950 ;
        RECT 631.950 414.450 634.050 415.050 ;
        RECT 634.950 414.450 637.050 415.050 ;
        RECT 631.950 413.400 637.050 414.450 ;
        RECT 631.950 412.950 634.050 413.400 ;
        RECT 634.950 412.950 637.050 413.400 ;
        RECT 637.950 412.950 640.050 415.050 ;
        RECT 640.950 412.950 643.050 415.050 ;
        RECT 644.250 413.250 646.050 414.150 ;
        RECT 646.950 412.950 649.050 415.050 ;
        RECT 649.950 413.250 651.750 414.150 ;
        RECT 652.950 412.950 655.050 415.050 ;
        RECT 656.250 413.250 657.750 414.150 ;
        RECT 658.950 412.950 661.050 415.050 ;
        RECT 662.250 413.250 664.050 414.150 ;
        RECT 628.950 403.950 631.050 406.050 ;
        RECT 632.400 403.050 633.450 412.950 ;
        RECT 634.950 410.850 637.050 411.750 ;
        RECT 637.950 410.250 640.050 411.150 ;
        RECT 640.950 410.850 642.750 411.750 ;
        RECT 643.950 409.950 646.050 412.050 ;
        RECT 637.950 406.950 640.050 409.050 ;
        RECT 638.400 406.050 639.450 406.950 ;
        RECT 637.950 403.950 640.050 406.050 ;
        RECT 631.950 400.950 634.050 403.050 ;
        RECT 622.950 394.950 625.050 397.050 ;
        RECT 613.950 391.950 616.050 394.050 ;
        RECT 637.950 391.950 640.050 394.050 ;
        RECT 616.950 385.950 619.050 388.050 ;
        RECT 631.950 385.950 634.050 388.050 ;
        RECT 617.400 382.050 618.450 385.950 ;
        RECT 622.950 382.950 625.050 385.050 ;
        RECT 623.400 382.050 624.450 382.950 ;
        RECT 632.400 382.050 633.450 385.950 ;
        RECT 613.950 380.250 615.750 381.150 ;
        RECT 616.950 379.950 619.050 382.050 ;
        RECT 622.950 379.950 625.050 382.050 ;
        RECT 625.950 379.950 628.050 382.050 ;
        RECT 631.950 379.950 634.050 382.050 ;
        RECT 635.250 380.250 637.050 381.150 ;
        RECT 613.950 376.950 616.050 379.050 ;
        RECT 617.250 377.850 618.750 378.750 ;
        RECT 619.950 376.950 622.050 379.050 ;
        RECT 623.250 377.850 625.050 378.750 ;
        RECT 625.950 377.850 627.750 378.750 ;
        RECT 628.950 376.950 631.050 379.050 ;
        RECT 632.250 377.850 633.750 378.750 ;
        RECT 634.950 376.950 637.050 379.050 ;
        RECT 613.950 373.950 616.050 376.050 ;
        RECT 619.950 374.850 622.050 375.750 ;
        RECT 628.950 374.850 631.050 375.750 ;
        RECT 610.950 355.950 613.050 358.050 ;
        RECT 610.950 343.950 613.050 346.050 ;
        RECT 611.400 343.050 612.450 343.950 ;
        RECT 614.400 343.050 615.450 373.950 ;
        RECT 631.950 367.950 634.050 370.050 ;
        RECT 632.400 361.050 633.450 367.950 ;
        RECT 619.950 358.950 622.050 361.050 ;
        RECT 631.950 358.950 634.050 361.050 ;
        RECT 607.950 341.250 609.750 342.150 ;
        RECT 610.950 340.950 613.050 343.050 ;
        RECT 613.950 340.950 616.050 343.050 ;
        RECT 616.950 340.950 619.050 343.050 ;
        RECT 607.950 339.450 610.050 340.050 ;
        RECT 605.400 338.400 610.050 339.450 ;
        RECT 611.250 338.850 613.050 339.750 ;
        RECT 607.950 337.950 610.050 338.400 ;
        RECT 613.950 338.250 616.050 339.150 ;
        RECT 616.950 338.850 619.050 339.750 ;
        RECT 610.950 334.950 613.050 337.050 ;
        RECT 613.950 334.950 616.050 337.050 ;
        RECT 601.950 322.950 604.050 325.050 ;
        RECT 592.950 319.950 595.050 322.050 ;
        RECT 583.950 313.950 586.050 316.050 ;
        RECT 601.950 313.950 604.050 316.050 ;
        RECT 607.950 313.950 610.050 316.050 ;
        RECT 602.400 313.050 603.450 313.950 ;
        RECT 608.400 313.050 609.450 313.950 ;
        RECT 611.400 313.050 612.450 334.950 ;
        RECT 620.400 334.050 621.450 358.950 ;
        RECT 635.400 354.450 636.450 376.950 ;
        RECT 638.400 354.450 639.450 391.950 ;
        RECT 640.950 385.950 643.050 388.050 ;
        RECT 641.400 370.050 642.450 385.950 ;
        RECT 644.400 384.450 645.450 409.950 ;
        RECT 647.400 388.050 648.450 412.950 ;
        RECT 649.950 409.950 652.050 412.050 ;
        RECT 653.250 410.850 654.750 411.750 ;
        RECT 655.950 409.950 658.050 412.050 ;
        RECT 659.250 410.850 660.750 411.750 ;
        RECT 661.950 409.950 664.050 412.050 ;
        RECT 649.950 406.950 652.050 409.050 ;
        RECT 655.950 406.950 658.050 409.050 ;
        RECT 646.950 385.950 649.050 388.050 ;
        RECT 650.400 385.050 651.450 406.950 ;
        RECT 652.950 385.950 655.050 388.050 ;
        RECT 653.400 385.050 654.450 385.950 ;
        RECT 644.400 383.400 648.450 384.450 ;
        RECT 647.400 382.050 648.450 383.400 ;
        RECT 649.950 382.950 652.050 385.050 ;
        RECT 652.950 382.950 655.050 385.050 ;
        RECT 643.950 380.250 645.750 381.150 ;
        RECT 646.950 379.950 649.050 382.050 ;
        RECT 649.950 379.950 652.050 382.050 ;
        RECT 652.950 381.450 655.050 382.050 ;
        RECT 656.400 381.450 657.450 406.950 ;
        RECT 658.950 400.950 661.050 403.050 ;
        RECT 659.400 388.050 660.450 400.950 ;
        RECT 661.950 397.950 664.050 400.050 ;
        RECT 662.400 388.050 663.450 397.950 ;
        RECT 665.400 388.050 666.450 437.400 ;
        RECT 667.950 421.950 670.050 424.050 ;
        RECT 668.400 406.050 669.450 421.950 ;
        RECT 671.400 418.050 672.450 442.950 ;
        RECT 674.400 421.050 675.450 445.950 ;
        RECT 682.950 444.450 685.050 445.050 ;
        RECT 685.950 444.450 688.050 445.050 ;
        RECT 682.950 443.400 688.050 444.450 ;
        RECT 682.950 442.950 685.050 443.400 ;
        RECT 685.950 442.950 688.050 443.400 ;
        RECT 689.400 442.050 690.450 469.950 ;
        RECT 692.400 454.050 693.450 478.950 ;
        RECT 695.400 460.050 696.450 481.950 ;
        RECT 698.400 481.050 699.450 484.950 ;
        RECT 700.950 481.950 703.050 484.050 ;
        RECT 704.250 482.850 705.750 483.750 ;
        RECT 706.950 481.950 709.050 484.050 ;
        RECT 709.950 481.950 712.050 484.050 ;
        RECT 713.250 482.850 714.750 483.750 ;
        RECT 715.950 481.950 718.050 484.050 ;
        RECT 697.950 478.950 700.050 481.050 ;
        RECT 698.400 460.050 699.450 478.950 ;
        RECT 701.400 478.050 702.450 481.950 ;
        RECT 707.400 478.050 708.450 481.950 ;
        RECT 710.400 481.050 711.450 481.950 ;
        RECT 709.950 478.950 712.050 481.050 ;
        RECT 700.950 475.950 703.050 478.050 ;
        RECT 706.950 475.950 709.050 478.050 ;
        RECT 715.950 475.950 718.050 478.050 ;
        RECT 712.950 472.950 715.050 475.050 ;
        RECT 709.950 466.950 712.050 469.050 ;
        RECT 703.950 460.950 706.050 463.050 ;
        RECT 704.400 460.050 705.450 460.950 ;
        RECT 710.400 460.050 711.450 466.950 ;
        RECT 694.950 457.950 697.050 460.050 ;
        RECT 697.950 457.950 700.050 460.050 ;
        RECT 703.950 457.950 706.050 460.050 ;
        RECT 709.950 457.950 712.050 460.050 ;
        RECT 694.950 455.250 697.050 456.150 ;
        RECT 697.950 455.850 700.050 456.750 ;
        RECT 700.950 455.250 703.050 456.150 ;
        RECT 703.950 455.850 706.050 456.750 ;
        RECT 706.950 455.250 708.750 456.150 ;
        RECT 709.950 454.950 712.050 457.050 ;
        RECT 691.950 451.950 694.050 454.050 ;
        RECT 694.950 451.950 697.050 454.050 ;
        RECT 697.950 451.950 700.050 454.050 ;
        RECT 700.950 451.950 703.050 454.050 ;
        RECT 703.950 451.950 706.050 454.050 ;
        RECT 706.950 451.950 709.050 454.050 ;
        RECT 710.250 452.850 712.050 453.750 ;
        RECT 691.950 448.950 694.050 451.050 ;
        RECT 688.950 439.950 691.050 442.050 ;
        RECT 682.950 436.950 685.050 439.050 ;
        RECT 688.950 436.950 691.050 439.050 ;
        RECT 676.950 433.950 679.050 436.050 ;
        RECT 673.950 418.950 676.050 421.050 ;
        RECT 677.400 418.050 678.450 433.950 ;
        RECT 679.950 424.950 682.050 427.050 ;
        RECT 670.950 415.950 673.050 418.050 ;
        RECT 674.250 416.250 675.750 417.150 ;
        RECT 676.950 415.950 679.050 418.050 ;
        RECT 670.950 413.850 672.750 414.750 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 677.250 413.850 679.050 414.750 ;
        RECT 670.950 409.950 673.050 412.050 ;
        RECT 667.950 403.950 670.050 406.050 ;
        RECT 667.950 397.950 670.050 400.050 ;
        RECT 658.950 385.950 661.050 388.050 ;
        RECT 661.950 385.950 664.050 388.050 ;
        RECT 664.950 385.950 667.050 388.050 ;
        RECT 658.950 383.250 661.050 384.150 ;
        RECT 661.950 383.850 664.050 384.750 ;
        RECT 664.950 382.950 667.050 385.050 ;
        RECT 652.950 380.400 657.450 381.450 ;
        RECT 652.950 379.950 655.050 380.400 ;
        RECT 650.400 379.050 651.450 379.950 ;
        RECT 643.950 376.950 646.050 379.050 ;
        RECT 647.250 377.850 648.750 378.750 ;
        RECT 649.950 376.950 652.050 379.050 ;
        RECT 653.250 377.850 655.050 378.750 ;
        RECT 644.400 373.050 645.450 376.950 ;
        RECT 646.950 373.950 649.050 376.050 ;
        RECT 649.950 374.850 652.050 375.750 ;
        RECT 652.950 373.950 655.050 376.050 ;
        RECT 643.950 370.950 646.050 373.050 ;
        RECT 640.950 367.950 643.050 370.050 ;
        RECT 640.950 361.950 643.050 364.050 ;
        RECT 635.400 353.400 639.450 354.450 ;
        RECT 634.950 349.950 637.050 352.050 ;
        RECT 625.950 347.250 628.050 348.150 ;
        RECT 631.950 346.950 634.050 349.050 ;
        RECT 632.400 346.050 633.450 346.950 ;
        RECT 622.950 344.250 624.750 345.150 ;
        RECT 625.950 343.950 628.050 346.050 ;
        RECT 629.250 344.250 630.750 345.150 ;
        RECT 631.950 343.950 634.050 346.050 ;
        RECT 622.950 340.950 625.050 343.050 ;
        RECT 628.950 340.950 631.050 343.050 ;
        RECT 632.250 341.850 634.050 342.750 ;
        RECT 623.400 337.050 624.450 340.950 ;
        RECT 622.950 334.950 625.050 337.050 ;
        RECT 613.950 331.950 616.050 334.050 ;
        RECT 619.950 331.950 622.050 334.050 ;
        RECT 583.950 310.950 586.050 313.050 ;
        RECT 589.950 310.950 592.050 313.050 ;
        RECT 595.950 312.450 598.050 313.050 ;
        RECT 593.250 311.250 594.750 312.150 ;
        RECT 595.950 311.400 600.450 312.450 ;
        RECT 595.950 310.950 598.050 311.400 ;
        RECT 578.400 305.400 582.450 306.450 ;
        RECT 571.950 295.950 574.050 298.050 ;
        RECT 574.950 295.950 577.050 298.050 ;
        RECT 565.950 271.950 568.050 274.050 ;
        RECT 548.250 269.250 549.750 270.150 ;
        RECT 550.950 269.400 555.450 270.450 ;
        RECT 550.950 268.950 553.050 269.400 ;
        RECT 556.950 269.250 559.050 270.150 ;
        RECT 559.950 268.950 562.050 271.050 ;
        RECT 562.950 269.250 565.050 270.150 ;
        RECT 565.950 268.950 568.050 271.050 ;
        RECT 568.950 269.250 571.050 270.150 ;
        RECT 541.950 265.950 544.050 268.050 ;
        RECT 545.250 266.850 546.750 267.750 ;
        RECT 547.950 265.950 550.050 268.050 ;
        RECT 553.950 265.950 556.050 268.050 ;
        RECT 556.950 265.950 559.050 268.050 ;
        RECT 560.250 266.250 561.750 267.150 ;
        RECT 562.950 265.950 565.050 268.050 ;
        RECT 532.950 259.950 535.050 262.050 ;
        RECT 538.950 259.950 541.050 262.050 ;
        RECT 529.950 250.950 532.050 253.050 ;
        RECT 515.400 242.400 519.450 243.450 ;
        RECT 518.400 241.050 519.450 242.400 ;
        RECT 529.950 241.950 532.050 244.050 ;
        RECT 530.400 241.050 531.450 241.950 ;
        RECT 505.950 238.950 508.050 241.050 ;
        RECT 508.950 239.850 511.050 240.750 ;
        RECT 511.950 239.250 514.050 240.150 ;
        RECT 514.950 238.950 517.050 241.050 ;
        RECT 517.950 238.950 520.050 241.050 ;
        RECT 521.250 239.250 522.750 240.150 ;
        RECT 523.950 238.950 526.050 241.050 ;
        RECT 527.250 239.250 528.750 240.150 ;
        RECT 529.950 238.950 532.050 241.050 ;
        RECT 499.950 236.250 501.750 237.150 ;
        RECT 502.950 235.950 505.050 238.050 ;
        RECT 506.250 236.250 508.050 237.150 ;
        RECT 511.950 235.950 514.050 238.050 ;
        RECT 499.950 234.450 502.050 235.050 ;
        RECT 497.400 233.400 502.050 234.450 ;
        RECT 503.250 233.850 504.750 234.750 ;
        RECT 494.400 208.050 495.450 232.950 ;
        RECT 490.950 205.950 493.050 208.050 ;
        RECT 493.950 205.950 496.050 208.050 ;
        RECT 484.950 202.950 487.050 205.050 ;
        RECT 457.950 199.950 460.050 202.050 ;
        RECT 461.250 200.250 462.750 201.150 ;
        RECT 463.950 199.950 466.050 202.050 ;
        RECT 466.950 200.250 468.750 201.150 ;
        RECT 469.950 199.950 472.050 202.050 ;
        RECT 473.250 200.250 474.750 201.150 ;
        RECT 475.950 199.950 478.050 202.050 ;
        RECT 478.950 199.950 481.050 202.050 ;
        RECT 457.950 197.850 459.750 198.750 ;
        RECT 460.950 196.950 463.050 199.050 ;
        RECT 464.250 197.850 466.050 198.750 ;
        RECT 466.950 196.950 469.050 199.050 ;
        RECT 449.400 194.400 453.450 195.450 ;
        RECT 434.400 173.400 438.450 174.450 ;
        RECT 421.950 166.950 424.050 169.050 ;
        RECT 425.250 167.250 426.750 168.150 ;
        RECT 427.950 166.950 430.050 169.050 ;
        RECT 430.950 166.950 433.050 169.050 ;
        RECT 421.950 164.850 423.750 165.750 ;
        RECT 424.950 163.950 427.050 166.050 ;
        RECT 428.250 164.850 429.750 165.750 ;
        RECT 430.950 163.950 433.050 166.050 ;
        RECT 419.400 161.400 423.450 162.450 ;
        RECT 430.950 161.850 433.050 162.750 ;
        RECT 409.950 142.950 412.050 145.050 ;
        RECT 415.950 142.950 418.050 145.050 ;
        RECT 391.950 139.950 394.050 142.050 ;
        RECT 397.950 139.950 400.050 142.050 ;
        RECT 392.400 130.050 393.450 139.950 ;
        RECT 397.950 133.950 400.050 136.050 ;
        RECT 412.950 133.950 415.050 136.050 ;
        RECT 391.950 127.950 394.050 130.050 ;
        RECT 392.400 127.050 393.450 127.950 ;
        RECT 398.400 127.050 399.450 133.950 ;
        RECT 403.950 131.250 406.050 132.150 ;
        RECT 400.950 128.250 402.750 129.150 ;
        RECT 403.950 127.950 406.050 130.050 ;
        RECT 407.250 128.250 408.750 129.150 ;
        RECT 409.950 127.950 412.050 130.050 ;
        RECT 413.400 127.050 414.450 133.950 ;
        RECT 388.950 125.250 390.750 126.150 ;
        RECT 391.950 124.950 394.050 127.050 ;
        RECT 397.950 124.950 400.050 127.050 ;
        RECT 400.950 124.950 403.050 127.050 ;
        RECT 406.950 124.950 409.050 127.050 ;
        RECT 410.250 125.850 412.050 126.750 ;
        RECT 412.950 124.950 415.050 127.050 ;
        RECT 385.950 121.950 388.050 124.050 ;
        RECT 388.950 121.950 391.050 124.050 ;
        RECT 392.250 122.850 394.050 123.750 ;
        RECT 394.950 122.250 397.050 123.150 ;
        RECT 397.950 122.850 400.050 123.750 ;
        RECT 379.950 109.950 382.050 112.050 ;
        RECT 382.950 109.950 385.050 112.050 ;
        RECT 367.950 97.950 370.050 100.050 ;
        RECT 373.950 97.950 376.050 100.050 ;
        RECT 374.400 97.050 375.450 97.950 ;
        RECT 358.950 96.450 361.050 97.050 ;
        RECT 361.950 96.450 364.050 97.050 ;
        RECT 358.950 95.400 364.050 96.450 ;
        RECT 358.950 94.950 361.050 95.400 ;
        RECT 361.950 94.950 364.050 95.400 ;
        RECT 365.250 95.250 366.750 96.150 ;
        RECT 367.950 94.950 370.050 97.050 ;
        RECT 371.250 95.250 372.750 96.150 ;
        RECT 373.950 94.950 376.050 97.050 ;
        RECT 376.950 94.950 379.050 97.050 ;
        RECT 349.950 92.850 352.050 93.750 ;
        RECT 352.950 92.250 355.050 93.150 ;
        RECT 355.950 91.950 358.050 94.050 ;
        RECT 358.950 92.850 361.050 93.750 ;
        RECT 361.950 92.850 363.750 93.750 ;
        RECT 364.950 91.950 367.050 94.050 ;
        RECT 368.250 92.850 369.750 93.750 ;
        RECT 370.950 91.950 373.050 94.050 ;
        RECT 374.250 92.850 376.050 93.750 ;
        RECT 346.950 88.950 349.050 91.050 ;
        RECT 352.950 90.450 355.050 91.050 ;
        RECT 356.400 90.450 357.450 91.950 ;
        RECT 352.950 89.400 357.450 90.450 ;
        RECT 352.950 88.950 355.050 89.400 ;
        RECT 328.950 85.950 331.050 88.050 ;
        RECT 334.950 79.950 337.050 82.050 ;
        RECT 335.400 70.050 336.450 79.950 ;
        RECT 347.400 70.050 348.450 88.950 ;
        RECT 358.950 85.950 361.050 88.050 ;
        RECT 334.950 67.950 337.050 70.050 ;
        RECT 346.950 67.950 349.050 70.050 ;
        RECT 335.400 58.050 336.450 67.950 ;
        RECT 340.950 59.250 343.050 60.150 ;
        RECT 352.950 59.250 355.050 60.150 ;
        RECT 359.400 58.050 360.450 85.950 ;
        RECT 377.400 64.050 378.450 94.950 ;
        RECT 380.400 94.050 381.450 109.950 ;
        RECT 389.400 106.050 390.450 121.950 ;
        RECT 401.400 121.050 402.450 124.950 ;
        RECT 394.950 118.950 397.050 121.050 ;
        RECT 400.950 118.950 403.050 121.050 ;
        RECT 394.950 109.950 397.050 112.050 ;
        RECT 397.950 109.950 400.050 112.050 ;
        RECT 388.950 103.950 391.050 106.050 ;
        RECT 391.950 100.950 394.050 103.050 ;
        RECT 382.950 97.950 385.050 100.050 ;
        RECT 379.950 91.950 382.050 94.050 ;
        RECT 383.400 91.050 384.450 97.950 ;
        RECT 385.950 91.950 388.050 94.050 ;
        RECT 389.250 92.250 391.050 93.150 ;
        RECT 379.950 89.850 381.750 90.750 ;
        RECT 382.950 88.950 385.050 91.050 ;
        RECT 386.250 89.850 387.750 90.750 ;
        RECT 388.950 88.950 391.050 91.050 ;
        RECT 382.950 86.850 385.050 87.750 ;
        RECT 382.950 70.950 385.050 73.050 ;
        RECT 376.950 61.950 379.050 64.050 ;
        RECT 376.950 59.250 379.050 60.150 ;
        RECT 383.400 58.050 384.450 70.950 ;
        RECT 385.950 61.950 388.050 64.050 ;
        RECT 386.400 61.050 387.450 61.950 ;
        RECT 389.400 61.050 390.450 88.950 ;
        RECT 392.400 73.050 393.450 100.950 ;
        RECT 395.400 90.450 396.450 109.950 ;
        RECT 398.400 97.050 399.450 109.950 ;
        RECT 407.400 109.050 408.450 124.950 ;
        RECT 406.950 106.950 409.050 109.050 ;
        RECT 416.400 108.450 417.450 142.950 ;
        RECT 422.400 130.050 423.450 161.400 ;
        RECT 434.400 138.450 435.450 173.400 ;
        RECT 442.950 169.950 445.050 172.050 ;
        RECT 443.400 166.050 444.450 169.950 ;
        RECT 439.950 164.250 441.750 165.150 ;
        RECT 442.950 163.950 445.050 166.050 ;
        RECT 446.250 164.250 448.050 165.150 ;
        RECT 439.950 160.950 442.050 163.050 ;
        RECT 443.250 161.850 444.750 162.750 ;
        RECT 445.950 160.950 448.050 163.050 ;
        RECT 449.400 162.450 450.450 194.400 ;
        RECT 467.400 193.050 468.450 196.950 ;
        RECT 470.400 196.050 471.450 199.950 ;
        RECT 485.400 199.050 486.450 202.950 ;
        RECT 490.950 200.250 493.050 201.150 ;
        RECT 494.400 199.050 495.450 205.950 ;
        RECT 497.400 202.050 498.450 233.400 ;
        RECT 499.950 232.950 502.050 233.400 ;
        RECT 505.950 232.950 508.050 235.050 ;
        RECT 515.400 234.450 516.450 238.950 ;
        RECT 517.950 236.850 519.750 237.750 ;
        RECT 520.950 235.950 523.050 238.050 ;
        RECT 524.250 236.850 525.750 237.750 ;
        RECT 526.950 235.950 529.050 238.050 ;
        RECT 530.250 236.850 532.050 237.750 ;
        RECT 512.400 233.400 516.450 234.450 ;
        RECT 499.950 229.950 502.050 232.050 ;
        RECT 500.400 202.050 501.450 229.950 ;
        RECT 506.400 220.050 507.450 232.950 ;
        RECT 505.950 217.950 508.050 220.050 ;
        RECT 508.950 214.950 511.050 217.050 ;
        RECT 496.950 199.950 499.050 202.050 ;
        RECT 499.950 199.950 502.050 202.050 ;
        RECT 505.950 200.250 508.050 201.150 ;
        RECT 500.400 199.050 501.450 199.950 ;
        RECT 472.950 196.950 475.050 199.050 ;
        RECT 476.250 197.850 478.050 198.750 ;
        RECT 478.950 196.950 481.050 199.050 ;
        RECT 481.950 197.250 483.750 198.150 ;
        RECT 484.950 196.950 487.050 199.050 ;
        RECT 488.250 197.250 489.750 198.150 ;
        RECT 490.950 196.950 493.050 199.050 ;
        RECT 493.950 196.950 496.050 199.050 ;
        RECT 496.950 197.250 498.750 198.150 ;
        RECT 499.950 196.950 502.050 199.050 ;
        RECT 503.250 197.250 504.750 198.150 ;
        RECT 505.950 196.950 508.050 199.050 ;
        RECT 469.950 193.950 472.050 196.050 ;
        RECT 475.950 193.950 478.050 196.050 ;
        RECT 460.950 190.950 463.050 193.050 ;
        RECT 466.950 190.950 469.050 193.050 ;
        RECT 451.950 169.950 454.050 172.050 ;
        RECT 454.950 169.950 457.050 172.050 ;
        RECT 452.400 169.050 453.450 169.950 ;
        RECT 451.950 166.950 454.050 169.050 ;
        RECT 455.250 167.850 456.750 168.750 ;
        RECT 457.950 166.950 460.050 169.050 ;
        RECT 451.950 164.850 454.050 165.750 ;
        RECT 457.950 164.850 460.050 165.750 ;
        RECT 449.400 161.400 453.450 162.450 ;
        RECT 440.400 160.050 441.450 160.950 ;
        RECT 436.950 157.950 439.050 160.050 ;
        RECT 439.950 157.950 442.050 160.050 ;
        RECT 437.400 148.050 438.450 157.950 ;
        RECT 436.950 145.950 439.050 148.050 ;
        RECT 434.400 137.400 438.450 138.450 ;
        RECT 433.950 133.950 436.050 136.050 ;
        RECT 427.950 131.250 430.050 132.150 ;
        RECT 434.400 130.050 435.450 133.950 ;
        RECT 418.950 127.950 421.050 130.050 ;
        RECT 421.950 127.950 424.050 130.050 ;
        RECT 425.250 128.250 426.750 129.150 ;
        RECT 427.950 127.950 430.050 130.050 ;
        RECT 431.250 128.250 433.050 129.150 ;
        RECT 433.950 127.950 436.050 130.050 ;
        RECT 419.400 112.050 420.450 127.950 ;
        RECT 421.950 125.850 423.750 126.750 ;
        RECT 424.950 124.950 427.050 127.050 ;
        RECT 425.400 124.050 426.450 124.950 ;
        RECT 421.950 121.950 424.050 124.050 ;
        RECT 424.950 121.950 427.050 124.050 ;
        RECT 418.950 109.950 421.050 112.050 ;
        RECT 416.400 107.400 420.450 108.450 ;
        RECT 412.950 100.950 415.050 103.050 ;
        RECT 413.400 100.050 414.450 100.950 ;
        RECT 403.950 97.950 406.050 100.050 ;
        RECT 412.950 97.950 415.050 100.050 ;
        RECT 397.950 94.950 400.050 97.050 ;
        RECT 397.950 92.250 399.750 93.150 ;
        RECT 400.950 91.950 403.050 94.050 ;
        RECT 404.400 91.050 405.450 97.950 ;
        RECT 419.400 97.050 420.450 107.400 ;
        RECT 409.950 95.250 412.050 96.150 ;
        RECT 412.950 95.850 415.050 96.750 ;
        RECT 415.950 95.250 417.750 96.150 ;
        RECT 418.950 94.950 421.050 97.050 ;
        RECT 406.950 93.450 409.050 94.050 ;
        RECT 409.950 93.450 412.050 94.050 ;
        RECT 406.950 92.400 412.050 93.450 ;
        RECT 406.950 91.950 409.050 92.400 ;
        RECT 409.950 91.950 412.050 92.400 ;
        RECT 415.950 91.950 418.050 94.050 ;
        RECT 419.250 92.850 421.050 93.750 ;
        RECT 397.950 90.450 400.050 91.050 ;
        RECT 395.400 89.400 400.050 90.450 ;
        RECT 401.250 89.850 402.750 90.750 ;
        RECT 397.950 88.950 400.050 89.400 ;
        RECT 403.950 88.950 406.050 91.050 ;
        RECT 407.250 89.850 409.050 90.750 ;
        RECT 403.950 86.850 406.050 87.750 ;
        RECT 397.950 82.950 400.050 85.050 ;
        RECT 391.950 70.950 394.050 73.050 ;
        RECT 385.950 58.950 388.050 61.050 ;
        RECT 388.950 58.950 391.050 61.050 ;
        RECT 391.950 59.250 394.050 60.150 ;
        RECT 398.400 58.050 399.450 82.950 ;
        RECT 410.400 82.050 411.450 91.950 ;
        RECT 412.950 88.950 415.050 91.050 ;
        RECT 409.950 79.950 412.050 82.050 ;
        RECT 409.950 67.950 412.050 70.050 ;
        RECT 410.400 58.050 411.450 67.950 ;
        RECT 413.400 58.050 414.450 88.950 ;
        RECT 416.400 82.050 417.450 91.950 ;
        RECT 415.950 79.950 418.050 82.050 ;
        RECT 422.400 76.050 423.450 121.950 ;
        RECT 428.400 106.050 429.450 127.950 ;
        RECT 430.950 124.950 433.050 127.050 ;
        RECT 433.950 124.950 436.050 127.050 ;
        RECT 430.950 121.950 433.050 124.050 ;
        RECT 431.400 121.050 432.450 121.950 ;
        RECT 430.950 118.950 433.050 121.050 ;
        RECT 434.400 112.050 435.450 124.950 ;
        RECT 433.950 109.950 436.050 112.050 ;
        RECT 427.950 103.950 430.050 106.050 ;
        RECT 437.400 100.050 438.450 137.400 ;
        RECT 439.950 128.250 442.050 129.150 ;
        RECT 439.950 124.950 442.050 127.050 ;
        RECT 443.250 125.250 444.750 126.150 ;
        RECT 445.950 124.950 448.050 127.050 ;
        RECT 449.250 125.250 451.050 126.150 ;
        RECT 440.400 109.050 441.450 124.950 ;
        RECT 442.950 121.950 445.050 124.050 ;
        RECT 446.250 122.850 447.750 123.750 ;
        RECT 448.950 121.950 451.050 124.050 ;
        RECT 449.400 121.050 450.450 121.950 ;
        RECT 448.950 118.950 451.050 121.050 ;
        RECT 439.950 106.950 442.050 109.050 ;
        RECT 442.950 103.950 445.050 106.050 ;
        RECT 439.950 100.950 442.050 103.050 ;
        RECT 436.950 97.950 439.050 100.050 ;
        RECT 440.400 97.050 441.450 100.950 ;
        RECT 427.950 96.450 430.050 97.050 ;
        RECT 425.400 95.400 430.050 96.450 ;
        RECT 425.400 85.050 426.450 95.400 ;
        RECT 427.950 94.950 430.050 95.400 ;
        RECT 431.250 95.250 432.750 96.150 ;
        RECT 433.950 94.950 436.050 97.050 ;
        RECT 437.250 95.250 438.750 96.150 ;
        RECT 439.950 94.950 442.050 97.050 ;
        RECT 443.400 94.050 444.450 103.950 ;
        RECT 452.400 97.050 453.450 161.400 ;
        RECT 454.950 139.950 457.050 142.050 ;
        RECT 455.400 130.050 456.450 139.950 ;
        RECT 461.400 133.050 462.450 190.950 ;
        RECT 476.400 190.050 477.450 193.950 ;
        RECT 479.400 192.450 480.450 196.950 ;
        RECT 481.950 193.950 484.050 196.050 ;
        RECT 485.250 194.850 486.750 195.750 ;
        RECT 487.950 193.950 490.050 196.050 ;
        RECT 493.950 193.950 496.050 196.050 ;
        RECT 496.950 193.950 499.050 196.050 ;
        RECT 500.250 194.850 501.750 195.750 ;
        RECT 502.950 193.950 505.050 196.050 ;
        RECT 488.400 192.450 489.450 193.950 ;
        RECT 479.400 191.400 489.450 192.450 ;
        RECT 475.950 187.950 478.050 190.050 ;
        RECT 490.950 187.950 493.050 190.050 ;
        RECT 472.950 175.950 475.050 178.050 ;
        RECT 478.950 175.950 481.050 178.050 ;
        RECT 466.950 166.950 469.050 169.050 ;
        RECT 467.400 166.050 468.450 166.950 ;
        RECT 463.950 164.250 465.750 165.150 ;
        RECT 466.950 163.950 469.050 166.050 ;
        RECT 470.250 164.250 472.050 165.150 ;
        RECT 473.400 163.050 474.450 175.950 ;
        RECT 475.950 169.950 478.050 172.050 ;
        RECT 463.950 160.950 466.050 163.050 ;
        RECT 467.250 161.850 468.750 162.750 ;
        RECT 469.950 160.950 472.050 163.050 ;
        RECT 472.950 160.950 475.050 163.050 ;
        RECT 470.400 148.050 471.450 160.950 ;
        RECT 469.950 145.950 472.050 148.050 ;
        RECT 476.400 142.050 477.450 169.950 ;
        RECT 479.400 169.050 480.450 175.950 ;
        RECT 484.950 169.950 487.050 172.050 ;
        RECT 485.400 169.050 486.450 169.950 ;
        RECT 491.400 169.050 492.450 187.950 ;
        RECT 494.400 177.450 495.450 193.950 ;
        RECT 497.400 193.050 498.450 193.950 ;
        RECT 496.950 190.950 499.050 193.050 ;
        RECT 499.950 178.950 502.050 181.050 ;
        RECT 494.400 176.400 498.450 177.450 ;
        RECT 497.400 169.050 498.450 176.400 ;
        RECT 478.950 166.950 481.050 169.050 ;
        RECT 482.250 167.250 483.750 168.150 ;
        RECT 484.950 166.950 487.050 169.050 ;
        RECT 490.950 168.450 493.050 169.050 ;
        RECT 488.250 167.250 489.750 168.150 ;
        RECT 490.950 167.400 495.450 168.450 ;
        RECT 490.950 166.950 493.050 167.400 ;
        RECT 494.400 166.050 495.450 167.400 ;
        RECT 496.950 166.950 499.050 169.050 ;
        RECT 500.400 166.050 501.450 178.950 ;
        RECT 503.400 178.050 504.450 193.950 ;
        RECT 502.950 175.950 505.050 178.050 ;
        RECT 505.950 169.950 508.050 172.050 ;
        RECT 509.400 171.450 510.450 214.950 ;
        RECT 512.400 196.050 513.450 233.400 ;
        RECT 521.400 220.050 522.450 235.950 ;
        RECT 523.950 232.950 526.050 235.050 ;
        RECT 524.400 229.050 525.450 232.950 ;
        RECT 527.400 229.050 528.450 235.950 ;
        RECT 523.950 226.950 526.050 229.050 ;
        RECT 526.950 226.950 529.050 229.050 ;
        RECT 520.950 217.950 523.050 220.050 ;
        RECT 533.400 217.050 534.450 259.950 ;
        RECT 548.400 253.050 549.450 265.950 ;
        RECT 538.950 250.950 541.050 253.050 ;
        RECT 547.950 250.950 550.050 253.050 ;
        RECT 539.400 241.050 540.450 250.950 ;
        RECT 554.400 244.050 555.450 265.950 ;
        RECT 557.400 265.050 558.450 265.950 ;
        RECT 556.950 262.950 559.050 265.050 ;
        RECT 559.950 262.950 562.050 265.050 ;
        RECT 560.400 250.050 561.450 262.950 ;
        RECT 559.950 247.950 562.050 250.050 ;
        RECT 559.950 244.950 562.050 247.050 ;
        RECT 544.950 241.950 547.050 244.050 ;
        RECT 547.950 241.950 550.050 244.050 ;
        RECT 553.950 241.950 556.050 244.050 ;
        RECT 545.400 241.050 546.450 241.950 ;
        RECT 535.950 238.950 538.050 241.050 ;
        RECT 538.950 238.950 541.050 241.050 ;
        RECT 542.250 239.250 543.750 240.150 ;
        RECT 544.950 238.950 547.050 241.050 ;
        RECT 532.950 214.950 535.050 217.050 ;
        RECT 536.400 211.050 537.450 238.950 ;
        RECT 548.400 238.050 549.450 241.950 ;
        RECT 553.950 238.950 556.050 241.050 ;
        RECT 556.950 238.950 559.050 241.050 ;
        RECT 554.400 238.050 555.450 238.950 ;
        RECT 538.950 236.850 540.750 237.750 ;
        RECT 541.950 235.950 544.050 238.050 ;
        RECT 545.250 236.850 546.750 237.750 ;
        RECT 547.950 235.950 550.050 238.050 ;
        RECT 553.950 235.950 556.050 238.050 ;
        RECT 538.950 223.950 541.050 226.050 ;
        RECT 520.950 208.950 523.050 211.050 ;
        RECT 535.950 208.950 538.050 211.050 ;
        RECT 517.950 199.950 520.050 202.050 ;
        RECT 518.400 199.050 519.450 199.950 ;
        RECT 517.950 196.950 520.050 199.050 ;
        RECT 511.950 193.950 514.050 196.050 ;
        RECT 514.950 194.250 517.050 195.150 ;
        RECT 517.950 194.850 520.050 195.750 ;
        RECT 514.950 190.950 517.050 193.050 ;
        RECT 517.950 178.950 520.050 181.050 ;
        RECT 511.950 171.450 514.050 172.050 ;
        RECT 509.400 170.400 514.050 171.450 ;
        RECT 478.950 164.850 480.750 165.750 ;
        RECT 481.950 163.950 484.050 166.050 ;
        RECT 485.250 164.850 486.750 165.750 ;
        RECT 487.950 163.950 490.050 166.050 ;
        RECT 491.250 164.850 493.050 165.750 ;
        RECT 493.950 163.950 496.050 166.050 ;
        RECT 499.950 163.950 502.050 166.050 ;
        RECT 503.250 164.250 505.050 165.150 ;
        RECT 482.400 160.050 483.450 163.950 ;
        RECT 488.400 163.050 489.450 163.950 ;
        RECT 487.950 160.950 490.050 163.050 ;
        RECT 493.950 161.850 495.750 162.750 ;
        RECT 496.950 160.950 499.050 163.050 ;
        RECT 500.250 161.850 501.750 162.750 ;
        RECT 502.950 160.950 505.050 163.050 ;
        RECT 481.950 157.950 484.050 160.050 ;
        RECT 488.400 148.050 489.450 160.950 ;
        RECT 496.950 158.850 499.050 159.750 ;
        RECT 490.950 151.950 493.050 154.050 ;
        RECT 491.400 148.050 492.450 151.950 ;
        RECT 493.950 148.950 496.050 151.050 ;
        RECT 499.950 148.950 502.050 151.050 ;
        RECT 487.950 145.950 490.050 148.050 ;
        RECT 490.950 145.950 493.050 148.050 ;
        RECT 475.950 139.950 478.050 142.050 ;
        RECT 460.950 130.950 463.050 133.050 ;
        RECT 454.950 127.950 457.050 130.050 ;
        RECT 476.400 127.050 477.450 139.950 ;
        RECT 487.950 130.950 490.050 133.050 ;
        RECT 488.400 130.050 489.450 130.950 ;
        RECT 494.400 130.050 495.450 148.950 ;
        RECT 500.400 130.050 501.450 148.950 ;
        RECT 503.400 136.050 504.450 160.950 ;
        RECT 506.400 142.050 507.450 169.950 ;
        RECT 505.950 139.950 508.050 142.050 ;
        RECT 502.950 133.950 505.050 136.050 ;
        RECT 487.950 127.950 490.050 130.050 ;
        RECT 491.250 128.250 492.750 129.150 ;
        RECT 493.950 127.950 496.050 130.050 ;
        RECT 499.950 127.950 502.050 130.050 ;
        RECT 503.400 129.450 504.450 133.950 ;
        RECT 509.400 133.050 510.450 170.400 ;
        RECT 511.950 169.950 514.050 170.400 ;
        RECT 511.950 167.850 514.050 168.750 ;
        RECT 514.950 167.250 517.050 168.150 ;
        RECT 514.950 163.950 517.050 166.050 ;
        RECT 508.950 130.950 511.050 133.050 ;
        RECT 515.400 130.050 516.450 163.950 ;
        RECT 518.400 160.050 519.450 178.950 ;
        RECT 517.950 157.950 520.050 160.050 ;
        RECT 521.400 142.050 522.450 208.950 ;
        RECT 539.400 205.050 540.450 223.950 ;
        RECT 542.400 223.050 543.450 235.950 ;
        RECT 557.400 235.050 558.450 238.950 ;
        RECT 560.400 238.050 561.450 244.950 ;
        RECT 563.400 241.050 564.450 265.950 ;
        RECT 566.400 241.050 567.450 268.950 ;
        RECT 568.950 267.450 571.050 268.050 ;
        RECT 572.400 267.450 573.450 295.950 ;
        RECT 574.950 289.950 577.050 292.050 ;
        RECT 575.400 279.450 576.450 289.950 ;
        RECT 578.400 289.050 579.450 305.400 ;
        RECT 580.950 301.950 583.050 304.050 ;
        RECT 581.400 301.050 582.450 301.950 ;
        RECT 580.950 298.950 583.050 301.050 ;
        RECT 584.400 292.050 585.450 310.950 ;
        RECT 586.950 307.950 589.050 310.050 ;
        RECT 590.250 308.850 591.750 309.750 ;
        RECT 592.950 307.950 595.050 310.050 ;
        RECT 596.250 308.850 598.050 309.750 ;
        RECT 586.950 305.850 589.050 306.750 ;
        RECT 589.950 304.950 592.050 307.050 ;
        RECT 592.950 304.950 595.050 307.050 ;
        RECT 586.950 301.950 589.050 304.050 ;
        RECT 583.950 289.950 586.050 292.050 ;
        RECT 577.950 286.950 580.050 289.050 ;
        RECT 575.400 278.400 579.450 279.450 ;
        RECT 574.950 269.250 577.050 270.150 ;
        RECT 568.950 266.400 573.450 267.450 ;
        RECT 568.950 265.950 571.050 266.400 ;
        RECT 574.950 265.950 577.050 268.050 ;
        RECT 568.950 262.950 571.050 265.050 ;
        RECT 562.950 238.950 565.050 241.050 ;
        RECT 565.950 238.950 568.050 241.050 ;
        RECT 569.400 238.050 570.450 262.950 ;
        RECT 575.400 262.050 576.450 265.950 ;
        RECT 571.950 259.950 574.050 262.050 ;
        RECT 574.950 259.950 577.050 262.050 ;
        RECT 572.400 238.050 573.450 259.950 ;
        RECT 578.400 241.050 579.450 278.400 ;
        RECT 580.950 277.950 583.050 280.050 ;
        RECT 581.400 244.050 582.450 277.950 ;
        RECT 583.950 274.950 586.050 277.050 ;
        RECT 587.400 276.450 588.450 301.950 ;
        RECT 590.400 286.050 591.450 304.950 ;
        RECT 593.400 298.050 594.450 304.950 ;
        RECT 599.400 298.050 600.450 311.400 ;
        RECT 601.950 310.950 604.050 313.050 ;
        RECT 605.250 311.250 606.750 312.150 ;
        RECT 607.950 310.950 610.050 313.050 ;
        RECT 610.950 310.950 613.050 313.050 ;
        RECT 601.950 308.850 603.750 309.750 ;
        RECT 604.950 307.950 607.050 310.050 ;
        RECT 608.250 308.850 609.750 309.750 ;
        RECT 610.950 307.950 613.050 310.050 ;
        RECT 605.400 298.050 606.450 307.950 ;
        RECT 610.950 305.850 613.050 306.750 ;
        RECT 592.950 295.950 595.050 298.050 ;
        RECT 598.950 295.950 601.050 298.050 ;
        RECT 604.950 295.950 607.050 298.050 ;
        RECT 610.950 289.950 613.050 292.050 ;
        RECT 589.950 283.950 592.050 286.050 ;
        RECT 601.950 277.950 604.050 280.050 ;
        RECT 602.400 277.050 603.450 277.950 ;
        RECT 587.400 275.400 591.450 276.450 ;
        RECT 584.400 274.050 585.450 274.950 ;
        RECT 590.400 274.050 591.450 275.400 ;
        RECT 595.950 274.950 598.050 277.050 ;
        RECT 601.950 274.950 604.050 277.050 ;
        RECT 583.950 271.950 586.050 274.050 ;
        RECT 587.250 272.250 588.750 273.150 ;
        RECT 589.950 271.950 592.050 274.050 ;
        RECT 596.400 271.050 597.450 274.950 ;
        RECT 602.400 271.050 603.450 274.950 ;
        RECT 607.950 271.950 610.050 274.050 ;
        RECT 583.950 269.850 585.750 270.750 ;
        RECT 586.950 268.950 589.050 271.050 ;
        RECT 590.250 269.850 592.050 270.750 ;
        RECT 592.950 269.250 594.750 270.150 ;
        RECT 595.950 268.950 598.050 271.050 ;
        RECT 599.250 269.250 600.750 270.150 ;
        RECT 601.950 268.950 604.050 271.050 ;
        RECT 605.250 269.250 607.050 270.150 ;
        RECT 587.400 259.050 588.450 268.950 ;
        RECT 592.950 265.950 595.050 268.050 ;
        RECT 596.250 266.850 597.750 267.750 ;
        RECT 598.950 265.950 601.050 268.050 ;
        RECT 602.250 266.850 603.750 267.750 ;
        RECT 604.950 267.450 607.050 268.050 ;
        RECT 608.400 267.450 609.450 271.950 ;
        RECT 604.950 266.400 609.450 267.450 ;
        RECT 604.950 265.950 607.050 266.400 ;
        RECT 598.950 262.950 601.050 265.050 ;
        RECT 601.950 262.950 604.050 265.050 ;
        RECT 586.950 256.950 589.050 259.050 ;
        RECT 583.950 253.950 586.050 256.050 ;
        RECT 584.400 244.050 585.450 253.950 ;
        RECT 587.400 244.050 588.450 256.950 ;
        RECT 589.950 253.950 592.050 256.050 ;
        RECT 590.400 244.050 591.450 253.950 ;
        RECT 595.950 250.950 598.050 253.050 ;
        RECT 580.950 241.950 583.050 244.050 ;
        RECT 583.950 241.950 586.050 244.050 ;
        RECT 586.950 241.950 589.050 244.050 ;
        RECT 589.950 241.950 592.050 244.050 ;
        RECT 592.950 241.950 595.050 244.050 ;
        RECT 577.950 238.950 580.050 241.050 ;
        RECT 584.400 240.450 585.450 241.950 ;
        RECT 593.400 241.050 594.450 241.950 ;
        RECT 586.950 240.450 589.050 241.050 ;
        RECT 584.400 239.400 589.050 240.450 ;
        RECT 590.250 239.850 591.750 240.750 ;
        RECT 586.950 238.950 589.050 239.400 ;
        RECT 592.950 238.950 595.050 241.050 ;
        RECT 559.950 235.950 562.050 238.050 ;
        RECT 563.250 236.250 565.050 237.150 ;
        RECT 565.950 235.950 568.050 238.050 ;
        RECT 568.950 235.950 571.050 238.050 ;
        RECT 571.950 235.950 574.050 238.050 ;
        RECT 574.950 236.250 576.750 237.150 ;
        RECT 577.950 235.950 580.050 238.050 ;
        RECT 581.250 236.250 583.050 237.150 ;
        RECT 583.950 235.950 586.050 238.050 ;
        RECT 586.950 236.850 589.050 237.750 ;
        RECT 589.950 235.950 592.050 238.050 ;
        RECT 592.950 236.850 595.050 237.750 ;
        RECT 547.950 233.850 550.050 234.750 ;
        RECT 553.950 233.850 555.750 234.750 ;
        RECT 556.950 232.950 559.050 235.050 ;
        RECT 560.250 233.850 561.750 234.750 ;
        RECT 562.950 232.950 565.050 235.050 ;
        RECT 550.950 229.950 553.050 232.050 ;
        RECT 556.950 230.850 559.050 231.750 ;
        RECT 566.400 231.450 567.450 235.950 ;
        RECT 568.950 232.950 571.050 235.050 ;
        RECT 574.950 234.450 577.050 235.050 ;
        RECT 572.400 233.400 577.050 234.450 ;
        RECT 578.250 233.850 579.750 234.750 ;
        RECT 563.400 230.400 567.450 231.450 ;
        RECT 551.400 229.050 552.450 229.950 ;
        RECT 550.950 226.950 553.050 229.050 ;
        RECT 541.950 220.950 544.050 223.050 ;
        RECT 553.950 211.950 556.050 214.050 ;
        RECT 547.950 208.950 550.050 211.050 ;
        RECT 550.950 208.950 553.050 211.050 ;
        RECT 544.950 205.950 547.050 208.050 ;
        RECT 535.950 203.250 538.050 204.150 ;
        RECT 538.950 202.950 541.050 205.050 ;
        RECT 541.950 202.950 544.050 205.050 ;
        RECT 542.400 202.050 543.450 202.950 ;
        RECT 529.950 201.450 532.050 202.050 ;
        RECT 527.400 200.400 532.050 201.450 ;
        RECT 527.400 199.050 528.450 200.400 ;
        RECT 529.950 199.950 532.050 200.400 ;
        RECT 532.950 200.250 534.750 201.150 ;
        RECT 535.950 199.950 538.050 202.050 ;
        RECT 539.250 200.250 540.750 201.150 ;
        RECT 541.950 199.950 544.050 202.050 ;
        RECT 526.950 196.950 529.050 199.050 ;
        RECT 529.950 196.950 532.050 199.050 ;
        RECT 532.950 196.950 535.050 199.050 ;
        RECT 523.950 194.250 526.050 195.150 ;
        RECT 526.950 194.850 529.050 195.750 ;
        RECT 530.400 193.050 531.450 196.950 ;
        RECT 536.400 196.050 537.450 199.950 ;
        RECT 545.400 199.050 546.450 205.950 ;
        RECT 538.950 196.950 541.050 199.050 ;
        RECT 542.250 197.850 544.050 198.750 ;
        RECT 544.950 196.950 547.050 199.050 ;
        RECT 532.950 193.950 535.050 196.050 ;
        RECT 535.950 193.950 538.050 196.050 ;
        RECT 544.950 193.950 547.050 196.050 ;
        RECT 523.950 190.950 526.050 193.050 ;
        RECT 529.950 190.950 532.050 193.050 ;
        RECT 526.950 166.950 529.050 169.050 ;
        RECT 527.400 166.050 528.450 166.950 ;
        RECT 523.950 164.250 525.750 165.150 ;
        RECT 526.950 163.950 529.050 166.050 ;
        RECT 530.250 164.250 532.050 165.150 ;
        RECT 533.400 163.050 534.450 193.950 ;
        RECT 535.950 175.950 538.050 178.050 ;
        RECT 523.950 160.950 526.050 163.050 ;
        RECT 527.250 161.850 528.750 162.750 ;
        RECT 529.950 160.950 532.050 163.050 ;
        RECT 532.950 160.950 535.050 163.050 ;
        RECT 530.400 151.050 531.450 160.950 ;
        RECT 536.400 154.050 537.450 175.950 ;
        RECT 545.400 172.050 546.450 193.950 ;
        RECT 548.400 172.050 549.450 208.950 ;
        RECT 551.400 208.050 552.450 208.950 ;
        RECT 550.950 205.950 553.050 208.050 ;
        RECT 554.400 204.450 555.450 211.950 ;
        RECT 551.400 203.400 555.450 204.450 ;
        RECT 551.400 202.050 552.450 203.400 ;
        RECT 550.950 199.950 553.050 202.050 ;
        RECT 554.250 200.250 555.750 201.150 ;
        RECT 556.950 199.950 559.050 202.050 ;
        RECT 550.950 197.850 552.750 198.750 ;
        RECT 553.950 196.950 556.050 199.050 ;
        RECT 557.250 197.850 559.050 198.750 ;
        RECT 559.950 197.250 562.050 198.150 ;
        RECT 559.950 193.950 562.050 196.050 ;
        RECT 556.950 181.950 559.050 184.050 ;
        RECT 544.950 169.950 547.050 172.050 ;
        RECT 547.950 169.950 550.050 172.050 ;
        RECT 547.950 166.950 550.050 169.050 ;
        RECT 538.950 164.250 540.750 165.150 ;
        RECT 541.950 163.950 544.050 166.050 ;
        RECT 545.250 164.250 547.050 165.150 ;
        RECT 538.950 160.950 541.050 163.050 ;
        RECT 542.250 161.850 543.750 162.750 ;
        RECT 544.950 160.950 547.050 163.050 ;
        RECT 539.400 160.050 540.450 160.950 ;
        RECT 538.950 157.950 541.050 160.050 ;
        RECT 544.950 157.950 547.050 160.050 ;
        RECT 545.400 157.050 546.450 157.950 ;
        RECT 544.950 154.950 547.050 157.050 ;
        RECT 535.950 151.950 538.050 154.050 ;
        RECT 544.950 151.950 547.050 154.050 ;
        RECT 529.950 148.950 532.050 151.050 ;
        RECT 529.950 142.950 532.050 145.050 ;
        RECT 538.950 142.950 541.050 145.050 ;
        RECT 517.950 139.950 520.050 142.050 ;
        RECT 520.950 139.950 523.050 142.050 ;
        RECT 503.400 128.400 507.450 129.450 ;
        RECT 454.950 125.250 456.750 126.150 ;
        RECT 457.950 124.950 460.050 127.050 ;
        RECT 463.950 126.450 466.050 127.050 ;
        RECT 463.950 125.400 468.450 126.450 ;
        RECT 463.950 124.950 466.050 125.400 ;
        RECT 454.950 121.950 457.050 124.050 ;
        RECT 458.250 122.850 460.050 123.750 ;
        RECT 460.950 122.250 463.050 123.150 ;
        RECT 463.950 122.850 466.050 123.750 ;
        RECT 455.400 121.050 456.450 121.950 ;
        RECT 454.950 118.950 457.050 121.050 ;
        RECT 457.950 118.950 460.050 121.050 ;
        RECT 460.950 118.950 463.050 121.050 ;
        RECT 458.400 117.450 459.450 118.950 ;
        RECT 455.400 116.400 459.450 117.450 ;
        RECT 455.400 100.050 456.450 116.400 ;
        RECT 461.400 100.050 462.450 118.950 ;
        RECT 467.400 103.050 468.450 125.400 ;
        RECT 469.950 124.950 472.050 127.050 ;
        RECT 472.950 125.250 474.750 126.150 ;
        RECT 475.950 124.950 478.050 127.050 ;
        RECT 481.950 124.950 484.050 127.050 ;
        RECT 487.950 125.850 489.750 126.750 ;
        RECT 490.950 124.950 493.050 127.050 ;
        RECT 494.250 125.850 496.050 126.750 ;
        RECT 499.950 124.950 502.050 127.050 ;
        RECT 502.950 124.950 505.050 127.050 ;
        RECT 506.400 126.450 507.450 128.400 ;
        RECT 508.950 128.250 511.050 129.150 ;
        RECT 514.950 127.950 517.050 130.050 ;
        RECT 518.400 129.450 519.450 139.950 ;
        RECT 518.400 128.400 522.450 129.450 ;
        RECT 508.950 126.450 511.050 127.050 ;
        RECT 506.400 125.400 511.050 126.450 ;
        RECT 508.950 124.950 511.050 125.400 ;
        RECT 512.250 125.250 513.750 126.150 ;
        RECT 514.950 124.950 517.050 127.050 ;
        RECT 518.250 125.250 520.050 126.150 ;
        RECT 470.400 121.050 471.450 124.950 ;
        RECT 472.950 121.950 475.050 124.050 ;
        RECT 476.250 122.850 478.050 123.750 ;
        RECT 478.950 122.250 481.050 123.150 ;
        RECT 481.950 122.850 484.050 123.750 ;
        RECT 469.950 118.950 472.050 121.050 ;
        RECT 473.400 118.050 474.450 121.950 ;
        RECT 475.950 118.950 478.050 121.050 ;
        RECT 478.950 118.950 481.050 121.050 ;
        RECT 472.950 115.950 475.050 118.050 ;
        RECT 466.950 100.950 469.050 103.050 ;
        RECT 454.950 97.950 457.050 100.050 ;
        RECT 457.950 97.950 460.050 100.050 ;
        RECT 460.950 97.950 463.050 100.050 ;
        RECT 469.950 97.950 472.050 100.050 ;
        RECT 445.950 94.950 448.050 97.050 ;
        RECT 451.950 94.950 454.050 97.050 ;
        RECT 446.400 94.050 447.450 94.950 ;
        RECT 427.950 92.850 429.750 93.750 ;
        RECT 430.950 91.950 433.050 94.050 ;
        RECT 434.250 92.850 435.750 93.750 ;
        RECT 436.950 91.950 439.050 94.050 ;
        RECT 440.250 92.850 442.050 93.750 ;
        RECT 442.950 91.950 445.050 94.050 ;
        RECT 445.950 91.950 448.050 94.050 ;
        RECT 451.950 91.950 454.050 94.050 ;
        RECT 455.250 92.250 457.050 93.150 ;
        RECT 431.400 88.050 432.450 91.950 ;
        RECT 439.950 88.950 442.050 91.050 ;
        RECT 442.950 88.950 445.050 91.050 ;
        RECT 445.950 89.850 447.750 90.750 ;
        RECT 448.950 88.950 451.050 91.050 ;
        RECT 452.250 89.850 453.750 90.750 ;
        RECT 454.950 88.950 457.050 91.050 ;
        RECT 430.950 85.950 433.050 88.050 ;
        RECT 424.950 82.950 427.050 85.050 ;
        RECT 421.950 73.950 424.050 76.050 ;
        RECT 418.950 67.950 421.050 70.050 ;
        RECT 427.950 67.950 430.050 70.050 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 334.950 55.950 337.050 58.050 ;
        RECT 338.250 56.250 339.750 57.150 ;
        RECT 340.950 55.950 343.050 58.050 ;
        RECT 344.250 56.250 346.050 57.150 ;
        RECT 349.950 56.250 351.750 57.150 ;
        RECT 352.950 55.950 355.050 58.050 ;
        RECT 356.250 56.250 357.750 57.150 ;
        RECT 358.950 55.950 361.050 58.050 ;
        RECT 364.950 55.950 367.050 58.050 ;
        RECT 373.950 56.250 375.750 57.150 ;
        RECT 376.950 55.950 379.050 58.050 ;
        RECT 380.250 56.250 381.750 57.150 ;
        RECT 382.950 55.950 385.050 58.050 ;
        RECT 385.950 55.950 388.050 58.050 ;
        RECT 388.950 56.250 390.750 57.150 ;
        RECT 391.950 55.950 394.050 58.050 ;
        RECT 395.250 56.250 396.750 57.150 ;
        RECT 397.950 55.950 400.050 58.050 ;
        RECT 409.950 55.950 412.050 58.050 ;
        RECT 412.950 55.950 415.050 58.050 ;
        RECT 415.950 56.250 418.050 57.150 ;
        RECT 316.950 52.950 319.050 55.050 ;
        RECT 319.950 52.950 322.050 55.050 ;
        RECT 322.950 52.950 325.050 55.050 ;
        RECT 326.250 53.250 328.050 54.150 ;
        RECT 329.400 52.050 330.450 55.950 ;
        RECT 334.950 53.850 336.750 54.750 ;
        RECT 337.950 52.950 340.050 55.050 ;
        RECT 310.950 50.400 315.450 51.450 ;
        RECT 316.950 50.850 319.050 51.750 ;
        RECT 310.950 49.950 313.050 50.400 ;
        RECT 319.950 50.250 322.050 51.150 ;
        RECT 322.950 50.850 324.750 51.750 ;
        RECT 325.950 49.950 328.050 52.050 ;
        RECT 328.950 49.950 331.050 52.050 ;
        RECT 305.400 49.050 306.450 49.950 ;
        RECT 304.950 46.950 307.050 49.050 ;
        RECT 313.950 46.950 316.050 49.050 ;
        RECT 319.950 46.950 322.050 49.050 ;
        RECT 322.950 46.950 325.050 49.050 ;
        RECT 304.950 43.950 307.050 46.050 ;
        RECT 305.400 42.450 306.450 43.950 ;
        RECT 302.400 41.400 306.450 42.450 ;
        RECT 274.950 34.950 277.050 37.050 ;
        RECT 256.950 31.950 259.050 34.050 ;
        RECT 262.950 31.950 265.050 34.050 ;
        RECT 271.950 31.950 274.050 34.050 ;
        RECT 250.950 25.950 253.050 28.050 ;
        RECT 235.950 22.950 238.050 25.050 ;
        RECT 239.250 23.250 241.050 24.150 ;
        RECT 241.950 23.850 244.050 24.750 ;
        RECT 244.950 23.250 247.050 24.150 ;
        RECT 247.950 22.950 250.050 25.050 ;
        RECT 220.950 19.950 223.050 22.050 ;
        RECT 224.250 20.850 225.750 21.750 ;
        RECT 226.950 19.950 229.050 22.050 ;
        RECT 230.250 20.850 232.050 21.750 ;
        RECT 232.950 19.950 235.050 22.050 ;
        RECT 235.950 20.850 237.750 21.750 ;
        RECT 238.950 19.950 241.050 22.050 ;
        RECT 244.950 19.950 247.050 22.050 ;
        RECT 247.950 21.450 250.050 22.050 ;
        RECT 251.400 21.450 252.450 25.950 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 257.400 24.450 258.450 31.950 ;
        RECT 265.950 25.950 268.050 28.050 ;
        RECT 272.400 25.050 273.450 31.950 ;
        RECT 257.400 23.400 261.450 24.450 ;
        RECT 254.400 22.050 255.450 22.950 ;
        RECT 247.950 20.400 252.450 21.450 ;
        RECT 247.950 19.950 250.050 20.400 ;
        RECT 253.950 19.950 256.050 22.050 ;
        RECT 260.400 21.450 261.450 23.400 ;
        RECT 262.950 23.250 265.050 24.150 ;
        RECT 265.950 23.850 268.050 24.750 ;
        RECT 268.950 23.250 270.750 24.150 ;
        RECT 271.950 22.950 274.050 25.050 ;
        RECT 275.400 22.050 276.450 34.950 ;
        RECT 278.400 25.050 279.450 40.950 ;
        RECT 287.400 31.050 288.450 40.950 ;
        RECT 286.950 28.950 289.050 31.050 ;
        RECT 298.950 28.950 301.050 31.050 ;
        RECT 277.950 22.950 280.050 25.050 ;
        RECT 281.250 23.250 282.750 24.150 ;
        RECT 283.950 22.950 286.050 25.050 ;
        RECT 287.400 22.050 288.450 28.950 ;
        RECT 292.950 25.950 295.050 28.050 ;
        RECT 293.400 22.050 294.450 25.950 ;
        RECT 295.950 22.950 298.050 25.050 ;
        RECT 262.950 21.450 265.050 22.050 ;
        RECT 257.250 20.250 259.050 21.150 ;
        RECT 260.400 20.400 265.050 21.450 ;
        RECT 262.950 19.950 265.050 20.400 ;
        RECT 268.950 19.950 271.050 22.050 ;
        RECT 272.250 20.850 274.050 21.750 ;
        RECT 274.950 19.950 277.050 22.050 ;
        RECT 277.950 20.850 279.750 21.750 ;
        RECT 280.950 19.950 283.050 22.050 ;
        RECT 284.250 20.850 285.750 21.750 ;
        RECT 286.950 19.950 289.050 22.050 ;
        RECT 292.950 19.950 295.050 22.050 ;
        RECT 263.400 19.050 264.450 19.950 ;
        RECT 296.400 19.050 297.450 22.950 ;
        RECT 299.400 22.050 300.450 28.950 ;
        RECT 298.950 19.950 301.050 22.050 ;
        RECT 302.250 20.250 304.050 21.150 ;
        RECT 208.950 17.400 213.450 18.450 ;
        RECT 220.950 17.850 223.050 18.750 ;
        RECT 247.950 17.850 249.750 18.750 ;
        RECT 208.950 16.950 211.050 17.400 ;
        RECT 250.950 16.950 253.050 19.050 ;
        RECT 254.250 17.850 255.750 18.750 ;
        RECT 256.950 18.450 259.050 19.050 ;
        RECT 259.950 18.450 262.050 19.050 ;
        RECT 256.950 17.400 262.050 18.450 ;
        RECT 256.950 16.950 259.050 17.400 ;
        RECT 259.950 16.950 262.050 17.400 ;
        RECT 262.950 16.950 265.050 19.050 ;
        RECT 265.950 18.450 268.050 19.050 ;
        RECT 268.950 18.450 271.050 19.050 ;
        RECT 265.950 17.400 271.050 18.450 ;
        RECT 286.950 17.850 289.050 18.750 ;
        RECT 292.950 17.850 294.750 18.750 ;
        RECT 265.950 16.950 268.050 17.400 ;
        RECT 268.950 16.950 271.050 17.400 ;
        RECT 295.950 16.950 298.050 19.050 ;
        RECT 299.250 17.850 300.750 18.750 ;
        RECT 301.950 18.450 304.050 19.050 ;
        RECT 305.400 18.450 306.450 41.400 ;
        RECT 314.400 25.050 315.450 46.950 ;
        RECT 323.400 43.050 324.450 46.950 ;
        RECT 322.950 40.950 325.050 43.050 ;
        RECT 326.400 37.050 327.450 49.950 ;
        RECT 341.400 46.050 342.450 55.950 ;
        RECT 343.950 52.950 346.050 55.050 ;
        RECT 349.950 52.950 352.050 55.050 ;
        RECT 340.950 43.950 343.050 46.050 ;
        RECT 344.400 43.050 345.450 52.950 ;
        RECT 350.400 52.050 351.450 52.950 ;
        RECT 349.950 49.950 352.050 52.050 ;
        RECT 353.400 46.050 354.450 55.950 ;
        RECT 355.950 52.950 358.050 55.050 ;
        RECT 359.250 53.850 361.050 54.750 ;
        RECT 352.950 43.950 355.050 46.050 ;
        RECT 343.950 40.950 346.050 43.050 ;
        RECT 356.400 42.450 357.450 52.950 ;
        RECT 350.400 41.400 357.450 42.450 ;
        RECT 340.950 37.950 343.050 40.050 ;
        RECT 325.950 34.950 328.050 37.050 ;
        RECT 319.950 25.950 322.050 28.050 ;
        RECT 313.950 22.950 316.050 25.050 ;
        RECT 317.250 23.250 319.050 24.150 ;
        RECT 319.950 23.850 322.050 24.750 ;
        RECT 322.950 23.250 325.050 24.150 ;
        RECT 313.950 20.850 315.750 21.750 ;
        RECT 316.950 19.950 319.050 22.050 ;
        RECT 322.950 19.950 325.050 22.050 ;
        RECT 326.400 19.050 327.450 34.950 ;
        RECT 331.950 25.950 334.050 28.050 ;
        RECT 334.950 25.950 337.050 28.050 ;
        RECT 328.950 22.950 331.050 25.050 ;
        RECT 329.400 22.050 330.450 22.950 ;
        RECT 328.950 19.950 331.050 22.050 ;
        RECT 332.400 19.050 333.450 25.950 ;
        RECT 335.400 22.050 336.450 25.950 ;
        RECT 334.950 19.950 337.050 22.050 ;
        RECT 338.250 20.250 340.050 21.150 ;
        RECT 301.950 17.400 306.450 18.450 ;
        RECT 301.950 16.950 304.050 17.400 ;
        RECT 325.950 16.950 328.050 19.050 ;
        RECT 328.950 17.850 330.750 18.750 ;
        RECT 331.950 16.950 334.050 19.050 ;
        RECT 335.250 17.850 336.750 18.750 ;
        RECT 337.950 18.450 340.050 19.050 ;
        RECT 341.400 18.450 342.450 37.950 ;
        RECT 346.950 25.950 349.050 28.050 ;
        RECT 347.400 22.050 348.450 25.950 ;
        RECT 350.400 25.050 351.450 41.400 ;
        RECT 358.950 34.950 361.050 37.050 ;
        RECT 355.950 31.950 358.050 34.050 ;
        RECT 356.400 25.050 357.450 31.950 ;
        RECT 359.400 25.050 360.450 34.950 ;
        RECT 365.400 25.050 366.450 55.950 ;
        RECT 367.950 52.950 370.050 55.050 ;
        RECT 373.950 52.950 376.050 55.050 ;
        RECT 379.950 54.450 382.050 55.050 ;
        RECT 377.400 53.400 382.050 54.450 ;
        RECT 383.250 53.850 385.050 54.750 ;
        RECT 374.400 52.050 375.450 52.950 ;
        RECT 367.950 50.850 370.050 51.750 ;
        RECT 370.950 50.250 373.050 51.150 ;
        RECT 373.950 49.950 376.050 52.050 ;
        RECT 370.950 46.950 373.050 49.050 ;
        RECT 371.400 43.050 372.450 46.950 ;
        RECT 377.400 46.050 378.450 53.400 ;
        RECT 379.950 52.950 382.050 53.400 ;
        RECT 386.400 49.050 387.450 55.950 ;
        RECT 392.400 55.050 393.450 55.950 ;
        RECT 410.400 55.050 411.450 55.950 ;
        RECT 388.950 52.950 391.050 55.050 ;
        RECT 391.950 52.950 394.050 55.050 ;
        RECT 394.950 52.950 397.050 55.050 ;
        RECT 398.250 53.850 400.050 54.750 ;
        RECT 406.950 53.250 408.750 54.150 ;
        RECT 409.950 52.950 412.050 55.050 ;
        RECT 415.950 54.450 418.050 55.050 ;
        RECT 419.400 54.450 420.450 67.950 ;
        RECT 424.950 61.950 427.050 64.050 ;
        RECT 425.400 61.050 426.450 61.950 ;
        RECT 424.950 58.950 427.050 61.050 ;
        RECT 421.950 55.950 424.050 58.050 ;
        RECT 422.400 55.050 423.450 55.950 ;
        RECT 425.400 55.050 426.450 58.950 ;
        RECT 428.400 55.050 429.450 67.950 ;
        RECT 440.400 61.050 441.450 88.950 ;
        RECT 443.400 85.050 444.450 88.950 ;
        RECT 458.400 88.050 459.450 97.950 ;
        RECT 460.950 94.950 463.050 97.050 ;
        RECT 463.950 94.950 466.050 97.050 ;
        RECT 467.250 95.250 469.050 96.150 ;
        RECT 469.950 95.850 472.050 96.750 ;
        RECT 472.950 95.250 475.050 96.150 ;
        RECT 461.400 91.050 462.450 94.950 ;
        RECT 463.950 92.850 465.750 93.750 ;
        RECT 466.950 91.950 469.050 94.050 ;
        RECT 472.950 91.950 475.050 94.050 ;
        RECT 460.950 88.950 463.050 91.050 ;
        RECT 445.950 85.950 448.050 88.050 ;
        RECT 448.950 86.850 451.050 87.750 ;
        RECT 457.950 85.950 460.050 88.050 ;
        RECT 446.400 85.050 447.450 85.950 ;
        RECT 473.400 85.050 474.450 91.950 ;
        RECT 476.400 85.050 477.450 118.950 ;
        RECT 479.400 118.050 480.450 118.950 ;
        RECT 478.950 115.950 481.050 118.050 ;
        RECT 487.950 109.950 490.050 112.050 ;
        RECT 488.400 106.050 489.450 109.950 ;
        RECT 484.950 103.950 487.050 106.050 ;
        RECT 487.950 103.950 490.050 106.050 ;
        RECT 481.950 100.950 484.050 103.050 ;
        RECT 482.400 100.050 483.450 100.950 ;
        RECT 481.950 97.950 484.050 100.050 ;
        RECT 478.950 95.250 481.050 96.150 ;
        RECT 481.950 95.850 484.050 96.750 ;
        RECT 478.950 91.950 481.050 94.050 ;
        RECT 481.950 91.950 484.050 94.050 ;
        RECT 442.950 82.950 445.050 85.050 ;
        RECT 445.950 82.950 448.050 85.050 ;
        RECT 472.950 82.950 475.050 85.050 ;
        RECT 475.950 82.950 478.050 85.050 ;
        RECT 482.400 82.050 483.450 91.950 ;
        RECT 485.400 90.450 486.450 103.950 ;
        RECT 491.400 103.050 492.450 124.950 ;
        RECT 496.950 122.250 499.050 123.150 ;
        RECT 499.950 122.850 502.050 123.750 ;
        RECT 503.400 121.050 504.450 124.950 ;
        RECT 521.400 124.050 522.450 128.400 ;
        RECT 523.950 128.250 526.050 129.150 ;
        RECT 530.400 127.050 531.450 142.950 ;
        RECT 539.400 127.050 540.450 142.950 ;
        RECT 545.400 136.050 546.450 151.950 ;
        RECT 544.950 133.950 547.050 136.050 ;
        RECT 548.400 133.050 549.450 166.950 ;
        RECT 550.950 164.250 552.750 165.150 ;
        RECT 553.950 163.950 556.050 166.050 ;
        RECT 557.400 163.050 558.450 181.950 ;
        RECT 559.950 172.950 562.050 175.050 ;
        RECT 560.400 166.050 561.450 172.950 ;
        RECT 563.400 166.050 564.450 230.400 ;
        RECT 569.400 228.450 570.450 232.950 ;
        RECT 566.400 227.400 570.450 228.450 ;
        RECT 566.400 202.050 567.450 227.400 ;
        RECT 568.950 223.950 571.050 226.050 ;
        RECT 569.400 208.050 570.450 223.950 ;
        RECT 568.950 205.950 571.050 208.050 ;
        RECT 572.400 202.050 573.450 233.400 ;
        RECT 574.950 232.950 577.050 233.400 ;
        RECT 580.950 232.950 583.050 235.050 ;
        RECT 574.950 229.950 577.050 232.050 ;
        RECT 575.400 211.050 576.450 229.950 ;
        RECT 574.950 208.950 577.050 211.050 ;
        RECT 581.400 208.050 582.450 232.950 ;
        RECT 584.400 220.050 585.450 235.950 ;
        RECT 590.400 226.050 591.450 235.950 ;
        RECT 596.400 235.050 597.450 250.950 ;
        RECT 592.950 232.950 595.050 235.050 ;
        RECT 595.950 232.950 598.050 235.050 ;
        RECT 589.950 223.950 592.050 226.050 ;
        RECT 583.950 217.950 586.050 220.050 ;
        RECT 593.400 214.050 594.450 232.950 ;
        RECT 599.400 231.450 600.450 262.950 ;
        RECT 602.400 241.050 603.450 262.950 ;
        RECT 605.400 262.050 606.450 265.950 ;
        RECT 604.950 259.950 607.050 262.050 ;
        RECT 607.950 250.950 610.050 253.050 ;
        RECT 608.400 243.450 609.450 250.950 ;
        RECT 611.400 247.050 612.450 289.950 ;
        RECT 614.400 265.050 615.450 331.950 ;
        RECT 623.400 319.050 624.450 334.950 ;
        RECT 629.400 322.050 630.450 340.950 ;
        RECT 631.950 337.950 634.050 340.050 ;
        RECT 635.400 339.450 636.450 349.950 ;
        RECT 638.400 346.050 639.450 353.400 ;
        RECT 637.950 343.950 640.050 346.050 ;
        RECT 641.400 343.050 642.450 361.950 ;
        RECT 647.400 349.050 648.450 373.950 ;
        RECT 653.400 367.050 654.450 373.950 ;
        RECT 652.950 364.950 655.050 367.050 ;
        RECT 656.400 352.050 657.450 380.400 ;
        RECT 658.950 379.950 661.050 382.050 ;
        RECT 661.950 379.950 664.050 382.050 ;
        RECT 659.400 379.050 660.450 379.950 ;
        RECT 658.950 376.950 661.050 379.050 ;
        RECT 658.950 355.950 661.050 358.050 ;
        RECT 655.950 349.950 658.050 352.050 ;
        RECT 646.950 346.950 649.050 349.050 ;
        RECT 649.950 346.950 652.050 349.050 ;
        RECT 646.950 344.250 649.050 345.150 ;
        RECT 637.950 341.250 639.750 342.150 ;
        RECT 640.950 340.950 643.050 343.050 ;
        RECT 646.950 342.450 649.050 343.050 ;
        RECT 650.400 342.450 651.450 346.950 ;
        RECT 652.950 343.950 655.050 346.050 ;
        RECT 644.250 341.250 645.750 342.150 ;
        RECT 646.950 341.400 651.450 342.450 ;
        RECT 646.950 340.950 649.050 341.400 ;
        RECT 637.950 339.450 640.050 340.050 ;
        RECT 635.400 338.400 640.050 339.450 ;
        RECT 641.250 338.850 642.750 339.750 ;
        RECT 637.950 337.950 640.050 338.400 ;
        RECT 643.950 337.950 646.050 340.050 ;
        RECT 628.950 319.950 631.050 322.050 ;
        RECT 616.950 316.950 619.050 319.050 ;
        RECT 622.950 316.950 625.050 319.050 ;
        RECT 617.400 310.050 618.450 316.950 ;
        RECT 623.400 316.050 624.450 316.950 ;
        RECT 619.950 313.950 622.050 316.050 ;
        RECT 622.950 313.950 625.050 316.050 ;
        RECT 628.950 313.950 631.050 316.050 ;
        RECT 632.400 315.450 633.450 337.950 ;
        RECT 637.950 322.950 640.050 325.050 ;
        RECT 632.400 314.400 636.450 315.450 ;
        RECT 616.950 307.950 619.050 310.050 ;
        RECT 616.950 304.950 619.050 307.050 ;
        RECT 617.400 301.050 618.450 304.950 ;
        RECT 616.950 298.950 619.050 301.050 ;
        RECT 620.400 295.050 621.450 313.950 ;
        RECT 622.950 310.950 625.050 313.050 ;
        RECT 626.250 311.250 628.050 312.150 ;
        RECT 628.950 311.850 631.050 312.750 ;
        RECT 631.950 311.250 634.050 312.150 ;
        RECT 622.950 308.850 624.750 309.750 ;
        RECT 625.950 307.950 628.050 310.050 ;
        RECT 628.950 307.950 631.050 310.050 ;
        RECT 631.950 307.950 634.050 310.050 ;
        RECT 619.950 292.950 622.050 295.050 ;
        RECT 619.950 289.950 622.050 292.050 ;
        RECT 620.400 271.050 621.450 289.950 ;
        RECT 629.400 280.050 630.450 307.950 ;
        RECT 632.400 295.050 633.450 307.950 ;
        RECT 635.400 304.050 636.450 314.400 ;
        RECT 638.400 304.050 639.450 322.950 ;
        RECT 644.400 322.050 645.450 337.950 ;
        RECT 640.950 319.950 643.050 322.050 ;
        RECT 643.950 319.950 646.050 322.050 ;
        RECT 641.400 313.050 642.450 319.950 ;
        RECT 647.400 316.050 648.450 340.950 ;
        RECT 653.400 336.450 654.450 343.950 ;
        RECT 659.400 343.050 660.450 355.950 ;
        RECT 662.400 355.050 663.450 379.950 ;
        RECT 661.950 352.950 664.050 355.050 ;
        RECT 665.400 351.450 666.450 382.950 ;
        RECT 668.400 382.050 669.450 397.950 ;
        RECT 671.400 394.050 672.450 409.950 ;
        RECT 674.400 400.050 675.450 412.950 ;
        RECT 676.950 409.950 679.050 412.050 ;
        RECT 677.400 403.050 678.450 409.950 ;
        RECT 676.950 400.950 679.050 403.050 ;
        RECT 673.950 397.950 676.050 400.050 ;
        RECT 676.950 394.950 679.050 397.050 ;
        RECT 677.400 394.050 678.450 394.950 ;
        RECT 670.950 391.950 673.050 394.050 ;
        RECT 676.950 391.950 679.050 394.050 ;
        RECT 670.950 388.950 673.050 391.050 ;
        RECT 671.400 385.050 672.450 388.950 ;
        RECT 677.400 385.050 678.450 391.950 ;
        RECT 670.950 382.950 673.050 385.050 ;
        RECT 674.250 383.250 675.750 384.150 ;
        RECT 676.950 382.950 679.050 385.050 ;
        RECT 667.950 379.950 670.050 382.050 ;
        RECT 671.250 380.850 672.750 381.750 ;
        RECT 673.950 379.950 676.050 382.050 ;
        RECT 677.250 380.850 679.050 381.750 ;
        RECT 667.950 377.850 670.050 378.750 ;
        RECT 667.950 367.950 670.050 370.050 ;
        RECT 662.400 350.400 666.450 351.450 ;
        RECT 662.400 346.050 663.450 350.400 ;
        RECT 661.950 343.950 664.050 346.050 ;
        RECT 664.950 343.950 667.050 346.050 ;
        RECT 665.400 343.050 666.450 343.950 ;
        RECT 655.950 341.250 657.750 342.150 ;
        RECT 658.950 340.950 661.050 343.050 ;
        RECT 664.950 340.950 667.050 343.050 ;
        RECT 655.950 337.950 658.050 340.050 ;
        RECT 659.250 338.850 661.050 339.750 ;
        RECT 661.950 338.250 664.050 339.150 ;
        RECT 664.950 338.850 667.050 339.750 ;
        RECT 668.400 339.450 669.450 367.950 ;
        RECT 674.400 367.050 675.450 379.950 ;
        RECT 680.400 376.050 681.450 424.950 ;
        RECT 683.400 421.050 684.450 436.950 ;
        RECT 685.950 433.950 688.050 436.050 ;
        RECT 682.950 418.950 685.050 421.050 ;
        RECT 686.400 418.050 687.450 433.950 ;
        RECT 685.950 415.950 688.050 418.050 ;
        RECT 686.400 415.050 687.450 415.950 ;
        RECT 689.400 415.050 690.450 436.950 ;
        RECT 692.400 433.050 693.450 448.950 ;
        RECT 695.400 448.050 696.450 451.950 ;
        RECT 694.950 445.950 697.050 448.050 ;
        RECT 698.400 436.050 699.450 451.950 ;
        RECT 701.400 448.050 702.450 451.950 ;
        RECT 700.950 445.950 703.050 448.050 ;
        RECT 700.950 442.950 703.050 445.050 ;
        RECT 697.950 433.950 700.050 436.050 ;
        RECT 691.950 430.950 694.050 433.050 ;
        RECT 701.400 427.050 702.450 442.950 ;
        RECT 704.400 433.050 705.450 451.950 ;
        RECT 713.400 445.050 714.450 472.950 ;
        RECT 716.400 454.050 717.450 475.950 ;
        RECT 719.400 472.050 720.450 484.950 ;
        RECT 722.400 475.050 723.450 488.400 ;
        RECT 734.400 487.050 735.450 514.950 ;
        RECT 740.400 492.450 741.450 535.950 ;
        RECT 743.400 535.050 744.450 580.950 ;
        RECT 745.950 562.950 748.050 565.050 ;
        RECT 746.400 562.050 747.450 562.950 ;
        RECT 749.400 562.050 750.450 583.950 ;
        RECT 745.950 559.950 748.050 562.050 ;
        RECT 748.950 559.950 751.050 562.050 ;
        RECT 745.950 557.850 748.050 558.750 ;
        RECT 748.950 557.250 751.050 558.150 ;
        RECT 748.950 553.950 751.050 556.050 ;
        RECT 742.950 532.950 745.050 535.050 ;
        RECT 742.950 529.950 745.050 532.050 ;
        RECT 742.950 527.850 745.050 528.750 ;
        RECT 745.950 527.250 748.050 528.150 ;
        RECT 745.950 523.950 748.050 526.050 ;
        RECT 752.400 523.050 753.450 595.950 ;
        RECT 755.400 592.050 756.450 595.950 ;
        RECT 761.400 594.450 762.450 622.950 ;
        RECT 764.400 621.450 765.450 626.400 ;
        RECT 767.400 625.050 768.450 667.950 ;
        RECT 769.950 634.950 772.050 637.050 ;
        RECT 766.950 622.950 769.050 625.050 ;
        RECT 764.400 620.400 768.450 621.450 ;
        RECT 763.950 601.950 766.050 604.050 ;
        RECT 758.400 593.400 762.450 594.450 ;
        RECT 754.950 589.950 757.050 592.050 ;
        RECT 754.950 586.950 757.050 589.050 ;
        RECT 755.400 538.050 756.450 586.950 ;
        RECT 754.950 535.950 757.050 538.050 ;
        RECT 754.950 524.850 757.050 525.750 ;
        RECT 745.950 520.950 748.050 523.050 ;
        RECT 751.950 520.950 754.050 523.050 ;
        RECT 737.400 491.400 741.450 492.450 ;
        RECT 724.950 485.250 727.050 486.150 ;
        RECT 730.950 485.250 733.050 486.150 ;
        RECT 733.950 484.950 736.050 487.050 ;
        RECT 724.950 481.950 727.050 484.050 ;
        RECT 730.950 483.450 733.050 484.050 ;
        RECT 733.950 483.450 736.050 484.050 ;
        RECT 728.250 482.250 729.750 483.150 ;
        RECT 730.950 482.400 736.050 483.450 ;
        RECT 730.950 481.950 733.050 482.400 ;
        RECT 733.950 481.950 736.050 482.400 ;
        RECT 725.400 481.050 726.450 481.950 ;
        RECT 724.950 478.950 727.050 481.050 ;
        RECT 727.950 478.950 730.050 481.050 ;
        RECT 730.950 478.950 733.050 481.050 ;
        RECT 725.400 478.050 726.450 478.950 ;
        RECT 724.950 475.950 727.050 478.050 ;
        RECT 721.950 472.950 724.050 475.050 ;
        RECT 727.950 472.950 730.050 475.050 ;
        RECT 718.950 469.950 721.050 472.050 ;
        RECT 718.950 463.950 721.050 466.050 ;
        RECT 721.950 463.950 724.050 466.050 ;
        RECT 719.400 463.050 720.450 463.950 ;
        RECT 718.950 460.950 721.050 463.050 ;
        RECT 719.400 457.050 720.450 460.950 ;
        RECT 722.400 460.050 723.450 463.950 ;
        RECT 721.950 457.950 724.050 460.050 ;
        RECT 724.950 457.950 727.050 460.050 ;
        RECT 725.400 457.050 726.450 457.950 ;
        RECT 718.950 454.950 721.050 457.050 ;
        RECT 722.250 455.850 723.750 456.750 ;
        RECT 724.950 454.950 727.050 457.050 ;
        RECT 728.400 456.450 729.450 472.950 ;
        RECT 731.400 460.050 732.450 478.950 ;
        RECT 734.400 463.050 735.450 481.950 ;
        RECT 737.400 475.050 738.450 491.400 ;
        RECT 742.950 484.950 745.050 487.050 ;
        RECT 742.950 482.850 745.050 483.750 ;
        RECT 736.950 472.950 739.050 475.050 ;
        RECT 736.950 466.950 739.050 469.050 ;
        RECT 733.950 460.950 736.050 463.050 ;
        RECT 734.400 460.050 735.450 460.950 ;
        RECT 730.950 457.950 733.050 460.050 ;
        RECT 733.950 457.950 736.050 460.050 ;
        RECT 737.400 457.050 738.450 466.950 ;
        RECT 728.400 455.400 732.450 456.450 ;
        RECT 733.950 455.850 735.750 456.750 ;
        RECT 715.950 451.950 718.050 454.050 ;
        RECT 718.950 452.850 721.050 453.750 ;
        RECT 724.950 452.850 727.050 453.750 ;
        RECT 727.950 451.950 730.050 454.050 ;
        RECT 728.400 450.450 729.450 451.950 ;
        RECT 725.400 449.400 729.450 450.450 ;
        RECT 718.950 445.950 721.050 448.050 ;
        RECT 712.950 442.950 715.050 445.050 ;
        RECT 706.950 439.950 709.050 442.050 ;
        RECT 703.950 430.950 706.050 433.050 ;
        RECT 703.950 427.950 706.050 430.050 ;
        RECT 700.950 424.950 703.050 427.050 ;
        RECT 697.950 419.250 700.050 420.150 ;
        RECT 704.400 418.050 705.450 427.950 ;
        RECT 694.950 416.250 696.750 417.150 ;
        RECT 697.950 415.950 700.050 418.050 ;
        RECT 701.250 416.250 702.750 417.150 ;
        RECT 703.950 415.950 706.050 418.050 ;
        RECT 682.950 413.250 684.750 414.150 ;
        RECT 685.950 412.950 688.050 415.050 ;
        RECT 688.950 412.950 691.050 415.050 ;
        RECT 691.950 412.950 694.050 415.050 ;
        RECT 694.950 412.950 697.050 415.050 ;
        RECT 700.950 412.950 703.050 415.050 ;
        RECT 704.250 413.850 706.050 414.750 ;
        RECT 682.950 409.950 685.050 412.050 ;
        RECT 686.250 410.850 688.050 411.750 ;
        RECT 688.950 410.250 691.050 411.150 ;
        RECT 691.950 410.850 694.050 411.750 ;
        RECT 688.950 408.450 691.050 409.050 ;
        RECT 695.400 408.450 696.450 412.950 ;
        RECT 688.950 407.400 696.450 408.450 ;
        RECT 688.950 406.950 691.050 407.400 ;
        RECT 688.950 403.950 691.050 406.050 ;
        RECT 685.950 394.950 688.050 397.050 ;
        RECT 682.950 385.950 685.050 388.050 ;
        RECT 679.950 373.950 682.050 376.050 ;
        RECT 673.950 364.950 676.050 367.050 ;
        RECT 670.950 346.950 673.050 349.050 ;
        RECT 676.950 347.250 679.050 348.150 ;
        RECT 671.400 346.050 672.450 346.950 ;
        RECT 670.950 343.950 673.050 346.050 ;
        RECT 674.250 344.250 675.750 345.150 ;
        RECT 676.950 343.950 679.050 346.050 ;
        RECT 680.250 344.250 682.050 345.150 ;
        RECT 670.950 341.850 672.750 342.750 ;
        RECT 673.950 340.950 676.050 343.050 ;
        RECT 668.400 338.400 672.450 339.450 ;
        RECT 671.400 337.050 672.450 338.400 ;
        RECT 653.400 335.400 657.450 336.450 ;
        RECT 652.950 331.950 655.050 334.050 ;
        RECT 649.950 316.950 652.050 319.050 ;
        RECT 643.950 313.950 646.050 316.050 ;
        RECT 646.950 313.950 649.050 316.050 ;
        RECT 640.950 310.950 643.050 313.050 ;
        RECT 644.400 312.450 645.450 313.950 ;
        RECT 644.400 311.400 648.450 312.450 ;
        RECT 640.950 308.250 642.750 309.150 ;
        RECT 643.950 307.950 646.050 310.050 ;
        RECT 647.400 307.050 648.450 311.400 ;
        RECT 650.400 310.050 651.450 316.950 ;
        RECT 649.950 307.950 652.050 310.050 ;
        RECT 640.950 304.950 643.050 307.050 ;
        RECT 644.250 305.850 645.750 306.750 ;
        RECT 646.950 304.950 649.050 307.050 ;
        RECT 650.250 305.850 652.050 306.750 ;
        RECT 634.950 301.950 637.050 304.050 ;
        RECT 637.950 301.950 640.050 304.050 ;
        RECT 643.950 301.950 646.050 304.050 ;
        RECT 646.950 302.850 649.050 303.750 ;
        RECT 634.950 295.950 637.050 298.050 ;
        RECT 640.950 295.950 643.050 298.050 ;
        RECT 631.950 292.950 634.050 295.050 ;
        RECT 628.950 277.950 631.050 280.050 ;
        RECT 631.950 274.950 634.050 277.050 ;
        RECT 632.400 274.050 633.450 274.950 ;
        RECT 625.950 271.950 628.050 274.050 ;
        RECT 629.250 272.250 630.750 273.150 ;
        RECT 631.950 271.950 634.050 274.050 ;
        RECT 616.950 269.250 619.050 270.150 ;
        RECT 619.950 268.950 622.050 271.050 ;
        RECT 622.950 269.250 625.050 270.150 ;
        RECT 625.950 269.850 627.750 270.750 ;
        RECT 628.950 268.950 631.050 271.050 ;
        RECT 632.250 269.850 634.050 270.750 ;
        RECT 616.950 265.950 619.050 268.050 ;
        RECT 620.250 266.250 621.750 267.150 ;
        RECT 622.950 265.950 625.050 268.050 ;
        RECT 625.950 265.950 628.050 268.050 ;
        RECT 613.950 262.950 616.050 265.050 ;
        RECT 617.400 259.050 618.450 265.950 ;
        RECT 619.950 262.950 622.050 265.050 ;
        RECT 623.400 262.050 624.450 265.950 ;
        RECT 619.950 259.950 622.050 262.050 ;
        RECT 622.950 259.950 625.050 262.050 ;
        RECT 616.950 256.950 619.050 259.050 ;
        RECT 620.400 256.050 621.450 259.950 ;
        RECT 616.950 253.950 619.050 256.050 ;
        RECT 619.950 253.950 622.050 256.050 ;
        RECT 613.950 247.950 616.050 250.050 ;
        RECT 610.950 244.950 613.050 247.050 ;
        RECT 610.950 243.450 613.050 244.050 ;
        RECT 608.400 242.400 613.050 243.450 ;
        RECT 610.950 241.950 613.050 242.400 ;
        RECT 614.400 241.050 615.450 247.950 ;
        RECT 601.950 238.950 604.050 241.050 ;
        RECT 610.950 239.850 612.750 240.750 ;
        RECT 613.950 238.950 616.050 241.050 ;
        RECT 601.950 236.250 603.750 237.150 ;
        RECT 604.950 235.950 607.050 238.050 ;
        RECT 608.250 236.250 610.050 237.150 ;
        RECT 610.950 235.950 613.050 238.050 ;
        RECT 613.950 236.850 616.050 237.750 ;
        RECT 601.950 232.950 604.050 235.050 ;
        RECT 605.250 233.850 606.750 234.750 ;
        RECT 607.950 232.950 610.050 235.050 ;
        RECT 599.400 230.400 603.450 231.450 ;
        RECT 595.950 226.950 598.050 229.050 ;
        RECT 596.400 223.050 597.450 226.950 ;
        RECT 595.950 220.950 598.050 223.050 ;
        RECT 592.950 211.950 595.050 214.050 ;
        RECT 592.950 208.950 595.050 211.050 ;
        RECT 598.950 208.950 601.050 211.050 ;
        RECT 580.950 205.950 583.050 208.050 ;
        RECT 589.950 202.950 592.050 205.050 ;
        RECT 565.950 199.950 568.050 202.050 ;
        RECT 571.950 199.950 574.050 202.050 ;
        RECT 577.950 199.950 580.050 202.050 ;
        RECT 583.950 199.950 586.050 202.050 ;
        RECT 565.950 197.850 568.050 198.750 ;
        RECT 568.950 197.250 571.050 198.150 ;
        RECT 568.950 193.950 571.050 196.050 ;
        RECT 569.400 187.050 570.450 193.950 ;
        RECT 568.950 184.950 571.050 187.050 ;
        RECT 572.400 181.050 573.450 199.950 ;
        RECT 578.400 199.050 579.450 199.950 ;
        RECT 584.400 199.050 585.450 199.950 ;
        RECT 574.950 197.250 576.750 198.150 ;
        RECT 577.950 196.950 580.050 199.050 ;
        RECT 581.250 197.250 582.750 198.150 ;
        RECT 583.950 196.950 586.050 199.050 ;
        RECT 587.250 197.250 589.050 198.150 ;
        RECT 574.950 193.950 577.050 196.050 ;
        RECT 578.250 194.850 579.750 195.750 ;
        RECT 580.950 193.950 583.050 196.050 ;
        RECT 584.250 194.850 585.750 195.750 ;
        RECT 586.950 193.950 589.050 196.050 ;
        RECT 575.400 190.050 576.450 193.950 ;
        RECT 581.400 193.050 582.450 193.950 ;
        RECT 580.950 190.950 583.050 193.050 ;
        RECT 586.950 190.950 589.050 193.050 ;
        RECT 574.950 187.950 577.050 190.050 ;
        RECT 571.950 178.950 574.050 181.050 ;
        RECT 565.950 175.950 568.050 178.050 ;
        RECT 559.950 163.950 562.050 166.050 ;
        RECT 562.950 163.950 565.050 166.050 ;
        RECT 550.950 160.950 553.050 163.050 ;
        RECT 554.250 161.850 555.750 162.750 ;
        RECT 556.950 160.950 559.050 163.050 ;
        RECT 560.250 161.850 562.050 162.750 ;
        RECT 551.400 157.050 552.450 160.950 ;
        RECT 556.950 158.850 559.050 159.750 ;
        RECT 550.950 154.950 553.050 157.050 ;
        RECT 566.400 151.050 567.450 175.950 ;
        RECT 571.950 166.950 574.050 169.050 ;
        RECT 577.950 168.450 580.050 169.050 ;
        RECT 581.400 168.450 582.450 190.950 ;
        RECT 587.400 178.050 588.450 190.950 ;
        RECT 590.400 181.050 591.450 202.950 ;
        RECT 593.400 195.450 594.450 208.950 ;
        RECT 599.400 208.050 600.450 208.950 ;
        RECT 598.950 205.950 601.050 208.050 ;
        RECT 595.950 202.950 598.050 205.050 ;
        RECT 596.400 202.050 597.450 202.950 ;
        RECT 595.950 199.950 598.050 202.050 ;
        RECT 595.950 197.250 598.050 198.150 ;
        RECT 599.400 196.050 600.450 205.950 ;
        RECT 602.400 202.050 603.450 230.400 ;
        RECT 611.400 229.050 612.450 235.950 ;
        RECT 610.950 226.950 613.050 229.050 ;
        RECT 610.950 214.950 613.050 217.050 ;
        RECT 604.950 211.950 607.050 214.050 ;
        RECT 605.400 202.050 606.450 211.950 ;
        RECT 607.950 202.950 610.050 205.050 ;
        RECT 601.950 199.950 604.050 202.050 ;
        RECT 604.950 199.950 607.050 202.050 ;
        RECT 601.950 197.850 604.050 198.750 ;
        RECT 604.950 197.250 607.050 198.150 ;
        RECT 595.950 195.450 598.050 196.050 ;
        RECT 593.400 194.400 598.050 195.450 ;
        RECT 593.400 190.050 594.450 194.400 ;
        RECT 595.950 193.950 598.050 194.400 ;
        RECT 598.950 193.950 601.050 196.050 ;
        RECT 604.950 193.950 607.050 196.050 ;
        RECT 605.400 190.050 606.450 193.950 ;
        RECT 592.950 187.950 595.050 190.050 ;
        RECT 604.950 187.950 607.050 190.050 ;
        RECT 601.950 181.950 604.050 184.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 586.950 175.950 589.050 178.050 ;
        RECT 589.950 175.950 592.050 178.050 ;
        RECT 598.950 175.950 601.050 178.050 ;
        RECT 575.250 167.250 576.750 168.150 ;
        RECT 577.950 167.400 582.450 168.450 ;
        RECT 577.950 166.950 580.050 167.400 ;
        RECT 568.950 163.950 571.050 166.050 ;
        RECT 572.250 164.850 573.750 165.750 ;
        RECT 574.950 163.950 577.050 166.050 ;
        RECT 578.250 164.850 580.050 165.750 ;
        RECT 580.950 163.950 583.050 166.050 ;
        RECT 583.950 164.250 585.750 165.150 ;
        RECT 586.950 163.950 589.050 166.050 ;
        RECT 575.400 163.050 576.450 163.950 ;
        RECT 568.950 161.850 571.050 162.750 ;
        RECT 574.950 160.950 577.050 163.050 ;
        RECT 568.950 154.950 571.050 157.050 ;
        RECT 565.950 148.950 568.050 151.050 ;
        RECT 569.400 136.050 570.450 154.950 ;
        RECT 562.950 133.950 565.050 136.050 ;
        RECT 568.950 133.950 571.050 136.050 ;
        RECT 547.950 130.950 550.050 133.050 ;
        RECT 553.950 131.250 556.050 132.150 ;
        RECT 544.950 128.250 547.050 129.150 ;
        RECT 523.950 124.950 526.050 127.050 ;
        RECT 527.250 125.250 528.750 126.150 ;
        RECT 529.950 124.950 532.050 127.050 ;
        RECT 533.250 125.250 535.050 126.150 ;
        RECT 535.950 125.250 537.750 126.150 ;
        RECT 538.950 124.950 541.050 127.050 ;
        RECT 544.950 126.450 547.050 127.050 ;
        RECT 548.400 126.450 549.450 130.950 ;
        RECT 550.950 128.250 552.750 129.150 ;
        RECT 553.950 127.950 556.050 130.050 ;
        RECT 557.250 128.250 558.750 129.150 ;
        RECT 559.950 127.950 562.050 130.050 ;
        RECT 542.250 125.250 543.750 126.150 ;
        RECT 544.950 125.400 549.450 126.450 ;
        RECT 544.950 124.950 547.050 125.400 ;
        RECT 550.950 124.950 553.050 127.050 ;
        RECT 511.950 121.950 514.050 124.050 ;
        RECT 515.250 122.850 516.750 123.750 ;
        RECT 517.950 123.450 520.050 124.050 ;
        RECT 520.950 123.450 523.050 124.050 ;
        RECT 517.950 122.400 523.050 123.450 ;
        RECT 517.950 121.950 520.050 122.400 ;
        RECT 520.950 121.950 523.050 122.400 ;
        RECT 496.950 118.950 499.050 121.050 ;
        RECT 502.950 118.950 505.050 121.050 ;
        RECT 512.400 115.050 513.450 121.950 ;
        RECT 524.400 118.050 525.450 124.950 ;
        RECT 551.400 124.050 552.450 124.950 ;
        RECT 526.950 121.950 529.050 124.050 ;
        RECT 530.250 122.850 531.750 123.750 ;
        RECT 532.950 121.950 535.050 124.050 ;
        RECT 535.950 121.950 538.050 124.050 ;
        RECT 539.250 122.850 540.750 123.750 ;
        RECT 541.950 121.950 544.050 124.050 ;
        RECT 544.950 121.950 547.050 124.050 ;
        RECT 547.950 121.950 550.050 124.050 ;
        RECT 550.950 121.950 553.050 124.050 ;
        RECT 523.950 115.950 526.050 118.050 ;
        RECT 511.950 112.950 514.050 115.050 ;
        RECT 527.400 112.050 528.450 121.950 ;
        RECT 542.400 115.050 543.450 121.950 ;
        RECT 541.950 112.950 544.050 115.050 ;
        RECT 526.950 109.950 529.050 112.050 ;
        RECT 490.950 100.950 493.050 103.050 ;
        RECT 502.950 100.950 505.050 103.050 ;
        RECT 514.950 100.950 517.050 103.050 ;
        RECT 490.950 97.950 493.050 100.050 ;
        RECT 491.400 94.050 492.450 97.950 ;
        RECT 487.950 92.250 489.750 93.150 ;
        RECT 490.950 91.950 493.050 94.050 ;
        RECT 496.950 93.450 499.050 94.050 ;
        RECT 496.950 92.400 501.450 93.450 ;
        RECT 496.950 91.950 499.050 92.400 ;
        RECT 487.950 90.450 490.050 91.050 ;
        RECT 485.400 89.400 490.050 90.450 ;
        RECT 491.250 89.850 492.750 90.750 ;
        RECT 487.950 88.950 490.050 89.400 ;
        RECT 493.950 88.950 496.050 91.050 ;
        RECT 497.250 89.850 499.050 90.750 ;
        RECT 493.950 86.850 496.050 87.750 ;
        RECT 500.400 85.050 501.450 92.400 ;
        RECT 499.950 82.950 502.050 85.050 ;
        RECT 481.950 79.950 484.050 82.050 ;
        RECT 460.950 76.950 463.050 79.050 ;
        RECT 439.950 58.950 442.050 61.050 ;
        RECT 454.950 59.250 457.050 60.150 ;
        RECT 461.400 58.050 462.450 76.950 ;
        RECT 463.950 70.950 466.050 73.050 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 445.950 56.250 448.050 57.150 ;
        RECT 451.950 56.250 453.750 57.150 ;
        RECT 454.950 55.950 457.050 58.050 ;
        RECT 458.250 56.250 459.750 57.150 ;
        RECT 460.950 55.950 463.050 58.050 ;
        RECT 413.250 53.250 414.750 54.150 ;
        RECT 415.950 53.400 420.450 54.450 ;
        RECT 415.950 52.950 418.050 53.400 ;
        RECT 421.950 52.950 424.050 55.050 ;
        RECT 424.950 52.950 427.050 55.050 ;
        RECT 427.950 52.950 430.050 55.050 ;
        RECT 431.250 53.250 433.050 54.150 ;
        RECT 379.950 46.950 382.050 49.050 ;
        RECT 385.950 46.950 388.050 49.050 ;
        RECT 376.950 43.950 379.050 46.050 ;
        RECT 370.950 40.950 373.050 43.050 ;
        RECT 371.400 37.050 372.450 40.950 ;
        RECT 377.400 40.050 378.450 43.950 ;
        RECT 376.950 37.950 379.050 40.050 ;
        RECT 370.950 34.950 373.050 37.050 ;
        RECT 367.950 28.950 370.050 31.050 ;
        RECT 349.950 22.950 352.050 25.050 ;
        RECT 353.250 23.250 354.750 24.150 ;
        RECT 355.950 22.950 358.050 25.050 ;
        RECT 358.950 22.950 361.050 25.050 ;
        RECT 362.250 23.250 363.750 24.150 ;
        RECT 364.950 22.950 367.050 25.050 ;
        RECT 368.400 22.050 369.450 28.950 ;
        RECT 373.950 25.950 376.050 28.050 ;
        RECT 374.400 24.450 375.450 25.950 ;
        RECT 376.950 24.450 379.050 25.200 ;
        RECT 374.400 23.400 379.050 24.450 ;
        RECT 376.950 23.100 379.050 23.400 ;
        RECT 346.950 19.950 349.050 22.050 ;
        RECT 350.250 20.850 351.750 21.750 ;
        RECT 352.950 19.950 355.050 22.050 ;
        RECT 356.250 20.850 358.050 21.750 ;
        RECT 358.950 20.850 360.750 21.750 ;
        RECT 361.950 19.950 364.050 22.050 ;
        RECT 365.250 20.850 366.750 21.750 ;
        RECT 367.950 19.950 370.050 22.050 ;
        RECT 376.950 21.000 379.050 21.900 ;
        RECT 380.400 21.450 381.450 46.950 ;
        RECT 389.400 37.050 390.450 52.950 ;
        RECT 391.950 49.950 394.050 52.050 ;
        RECT 392.400 49.050 393.450 49.950 ;
        RECT 391.950 46.950 394.050 49.050 ;
        RECT 395.400 46.050 396.450 52.950 ;
        RECT 406.950 49.950 409.050 52.050 ;
        RECT 410.250 50.850 411.750 51.750 ;
        RECT 412.950 49.950 415.050 52.050 ;
        RECT 421.950 50.850 424.050 51.750 ;
        RECT 424.950 50.250 427.050 51.150 ;
        RECT 427.950 50.850 429.750 51.750 ;
        RECT 430.950 49.950 433.050 52.050 ;
        RECT 394.950 43.950 397.050 46.050 ;
        RECT 391.950 37.950 394.050 40.050 ;
        RECT 388.950 34.950 391.050 37.050 ;
        RECT 392.400 27.450 393.450 37.950 ;
        RECT 389.400 26.400 393.450 27.450 ;
        RECT 403.950 27.450 406.050 28.050 ;
        RECT 407.400 27.450 408.450 49.950 ;
        RECT 413.400 46.050 414.450 49.950 ;
        RECT 424.950 46.950 427.050 49.050 ;
        RECT 412.950 43.950 415.050 46.050 ;
        RECT 434.400 40.050 435.450 55.950 ;
        RECT 455.400 55.050 456.450 55.950 ;
        RECT 436.950 53.250 438.750 54.150 ;
        RECT 439.950 52.950 442.050 55.050 ;
        RECT 443.250 53.250 444.750 54.150 ;
        RECT 445.950 52.950 448.050 55.050 ;
        RECT 451.950 52.950 454.050 55.050 ;
        RECT 454.950 52.950 457.050 55.050 ;
        RECT 457.950 52.950 460.050 55.050 ;
        RECT 461.250 53.850 463.050 54.750 ;
        RECT 436.950 49.950 439.050 52.050 ;
        RECT 440.250 50.850 441.750 51.750 ;
        RECT 442.950 49.950 445.050 52.050 ;
        RECT 448.950 49.950 451.050 52.050 ;
        RECT 437.400 49.050 438.450 49.950 ;
        RECT 436.950 46.950 439.050 49.050 ;
        RECT 439.950 40.950 442.050 43.050 ;
        RECT 412.950 37.950 415.050 40.050 ;
        RECT 433.950 37.950 436.050 40.050 ;
        RECT 413.400 34.050 414.450 37.950 ;
        RECT 412.950 31.950 415.050 34.050 ;
        RECT 403.950 26.400 408.450 27.450 ;
        RECT 385.950 24.450 388.050 25.200 ;
        RECT 389.400 24.450 390.450 26.400 ;
        RECT 403.950 25.950 406.050 26.400 ;
        RECT 409.950 25.950 412.050 28.050 ;
        RECT 404.400 25.050 405.450 25.950 ;
        RECT 410.400 25.050 411.450 25.950 ;
        RECT 382.950 23.400 384.750 24.300 ;
        RECT 385.950 23.400 390.450 24.450 ;
        RECT 391.950 23.400 394.050 24.300 ;
        RECT 385.950 23.100 388.050 23.400 ;
        RECT 403.950 22.950 406.050 25.050 ;
        RECT 407.250 23.250 408.750 24.150 ;
        RECT 409.950 22.950 412.050 25.050 ;
        RECT 382.950 21.450 385.050 22.200 ;
        RECT 380.400 20.400 385.050 21.450 ;
        RECT 386.250 21.000 388.050 21.900 ;
        RECT 382.950 20.100 385.050 20.400 ;
        RECT 353.400 19.050 354.450 19.950 ;
        RECT 383.400 19.050 384.450 20.100 ;
        RECT 391.950 19.950 394.050 22.200 ;
        RECT 413.400 22.050 414.450 31.950 ;
        RECT 430.950 25.950 433.050 28.050 ;
        RECT 440.400 25.050 441.450 40.950 ;
        RECT 443.400 31.050 444.450 49.950 ;
        RECT 449.400 34.050 450.450 49.950 ;
        RECT 448.950 31.950 451.050 34.050 ;
        RECT 442.950 28.950 445.050 31.050 ;
        RECT 452.400 28.050 453.450 52.950 ;
        RECT 451.950 25.950 454.050 28.050 ;
        RECT 424.950 22.950 427.050 25.050 ;
        RECT 428.250 23.250 430.050 24.150 ;
        RECT 430.950 23.850 433.050 24.750 ;
        RECT 439.950 24.450 442.050 25.050 ;
        RECT 433.950 23.250 436.050 24.150 ;
        RECT 437.400 23.400 442.050 24.450 ;
        RECT 403.950 20.850 405.750 21.750 ;
        RECT 406.950 19.950 409.050 22.050 ;
        RECT 410.250 20.850 411.750 21.750 ;
        RECT 412.950 19.950 415.050 22.050 ;
        RECT 424.950 20.850 426.750 21.750 ;
        RECT 427.950 19.950 430.050 22.050 ;
        RECT 433.950 21.450 436.050 22.050 ;
        RECT 437.400 21.450 438.450 23.400 ;
        RECT 439.950 22.950 442.050 23.400 ;
        RECT 448.950 22.950 451.050 25.050 ;
        RECT 452.400 22.050 453.450 25.950 ;
        RECT 455.400 24.450 456.450 52.950 ;
        RECT 458.400 43.050 459.450 52.950 ;
        RECT 464.400 52.050 465.450 70.950 ;
        RECT 466.950 67.950 469.050 70.050 ;
        RECT 467.400 55.050 468.450 67.950 ;
        RECT 481.950 61.950 484.050 64.050 ;
        RECT 475.950 59.250 478.050 60.150 ;
        RECT 482.400 58.050 483.450 61.950 ;
        RECT 487.950 59.250 490.050 60.150 ;
        RECT 503.400 58.050 504.450 100.950 ;
        RECT 505.950 97.950 508.050 100.050 ;
        RECT 506.400 94.050 507.450 97.950 ;
        RECT 515.400 97.050 516.450 100.950 ;
        RECT 517.950 97.950 520.050 100.050 ;
        RECT 526.950 97.950 529.050 100.050 ;
        RECT 541.950 97.950 544.050 100.050 ;
        RECT 545.400 99.450 546.450 121.950 ;
        RECT 548.400 103.050 549.450 121.950 ;
        RECT 551.400 121.050 552.450 121.950 ;
        RECT 554.400 121.050 555.450 127.950 ;
        RECT 563.400 127.050 564.450 133.950 ;
        RECT 571.950 131.250 574.050 132.150 ;
        RECT 565.950 127.950 568.050 130.050 ;
        RECT 568.950 128.250 570.750 129.150 ;
        RECT 571.950 127.950 574.050 130.050 ;
        RECT 575.250 128.250 576.750 129.150 ;
        RECT 577.950 127.950 580.050 130.050 ;
        RECT 556.950 124.950 559.050 127.050 ;
        RECT 560.250 125.850 562.050 126.750 ;
        RECT 562.950 124.950 565.050 127.050 ;
        RECT 550.950 118.950 553.050 121.050 ;
        RECT 553.950 118.950 556.050 121.050 ;
        RECT 554.400 118.050 555.450 118.950 ;
        RECT 566.400 118.050 567.450 127.950 ;
        RECT 568.950 124.950 571.050 127.050 ;
        RECT 569.400 124.050 570.450 124.950 ;
        RECT 568.950 121.950 571.050 124.050 ;
        RECT 553.950 115.950 556.050 118.050 ;
        RECT 565.950 115.950 568.050 118.050 ;
        RECT 550.950 103.950 553.050 106.050 ;
        RECT 547.950 100.950 550.050 103.050 ;
        RECT 545.400 98.400 549.450 99.450 ;
        RECT 508.950 94.950 511.050 97.050 ;
        RECT 512.250 95.250 513.750 96.150 ;
        RECT 514.950 94.950 517.050 97.050 ;
        RECT 505.950 91.950 508.050 94.050 ;
        RECT 509.250 92.850 510.750 93.750 ;
        RECT 511.950 91.950 514.050 94.050 ;
        RECT 515.250 92.850 517.050 93.750 ;
        RECT 505.950 89.850 508.050 90.750 ;
        RECT 514.950 88.950 517.050 91.050 ;
        RECT 518.400 90.450 519.450 97.950 ;
        RECT 520.950 92.250 522.750 93.150 ;
        RECT 523.950 91.950 526.050 94.050 ;
        RECT 527.400 91.050 528.450 97.950 ;
        RECT 535.950 94.950 538.050 97.050 ;
        RECT 539.250 95.250 541.050 96.150 ;
        RECT 541.950 95.850 544.050 96.750 ;
        RECT 544.950 95.250 547.050 96.150 ;
        RECT 529.950 93.450 532.050 94.050 ;
        RECT 529.950 92.400 534.450 93.450 ;
        RECT 535.950 92.850 537.750 93.750 ;
        RECT 529.950 91.950 532.050 92.400 ;
        RECT 533.400 91.050 534.450 92.400 ;
        RECT 538.950 91.950 541.050 94.050 ;
        RECT 544.950 91.950 547.050 94.050 ;
        RECT 520.950 90.450 523.050 91.050 ;
        RECT 518.400 89.400 523.050 90.450 ;
        RECT 524.250 89.850 525.750 90.750 ;
        RECT 520.950 88.950 523.050 89.400 ;
        RECT 526.950 88.950 529.050 91.050 ;
        RECT 530.250 89.850 532.050 90.750 ;
        RECT 532.950 88.950 535.050 91.050 ;
        RECT 515.400 79.050 516.450 88.950 ;
        RECT 526.950 86.850 529.050 87.750 ;
        RECT 514.950 76.950 517.050 79.050 ;
        RECT 517.950 59.250 520.050 60.150 ;
        RECT 533.400 58.050 534.450 88.950 ;
        RECT 539.400 67.050 540.450 91.950 ;
        RECT 545.400 91.050 546.450 91.950 ;
        RECT 544.950 88.950 547.050 91.050 ;
        RECT 544.950 85.950 547.050 88.050 ;
        RECT 541.950 76.950 544.050 79.050 ;
        RECT 538.950 64.950 541.050 67.050 ;
        RECT 469.950 55.950 472.050 58.050 ;
        RECT 473.250 56.250 474.750 57.150 ;
        RECT 475.950 55.950 478.050 58.050 ;
        RECT 479.250 56.250 481.050 57.150 ;
        RECT 481.950 55.950 484.050 58.050 ;
        RECT 484.950 56.250 486.750 57.150 ;
        RECT 487.950 55.950 490.050 58.050 ;
        RECT 491.250 56.250 492.750 57.150 ;
        RECT 493.950 55.950 496.050 58.050 ;
        RECT 496.950 55.950 499.050 58.050 ;
        RECT 499.950 55.950 502.050 58.050 ;
        RECT 502.950 55.950 505.050 58.050 ;
        RECT 511.950 55.950 514.050 58.050 ;
        RECT 514.950 56.250 516.750 57.150 ;
        RECT 517.950 55.950 520.050 58.050 ;
        RECT 521.250 56.250 522.750 57.150 ;
        RECT 523.950 55.950 526.050 58.050 ;
        RECT 532.950 55.950 535.050 58.050 ;
        RECT 538.950 56.250 541.050 57.150 ;
        RECT 466.950 52.950 469.050 55.050 ;
        RECT 469.950 53.850 471.750 54.750 ;
        RECT 472.950 52.950 475.050 55.050 ;
        RECT 478.950 52.950 481.050 55.050 ;
        RECT 484.950 52.950 487.050 55.050 ;
        RECT 490.950 52.950 493.050 55.050 ;
        RECT 494.250 53.850 496.050 54.750 ;
        RECT 463.950 49.950 466.050 52.050 ;
        RECT 475.950 51.450 478.050 52.050 ;
        RECT 473.400 50.400 478.050 51.450 ;
        RECT 473.400 46.050 474.450 50.400 ;
        RECT 475.950 49.950 478.050 50.400 ;
        RECT 475.950 46.950 478.050 49.050 ;
        RECT 476.400 46.050 477.450 46.950 ;
        RECT 472.950 43.950 475.050 46.050 ;
        RECT 475.950 43.950 478.050 46.050 ;
        RECT 457.950 40.950 460.050 43.050 ;
        RECT 463.950 40.950 466.050 43.050 ;
        RECT 464.400 25.050 465.450 40.950 ;
        RECT 469.950 25.950 472.050 28.050 ;
        RECT 470.400 25.050 471.450 25.950 ;
        RECT 457.950 24.450 460.050 25.050 ;
        RECT 455.400 23.400 460.050 24.450 ;
        RECT 457.950 22.950 460.050 23.400 ;
        RECT 461.250 23.250 462.750 24.150 ;
        RECT 463.950 22.950 466.050 25.050 ;
        RECT 467.250 23.250 468.750 24.150 ;
        RECT 469.950 22.950 472.050 25.050 ;
        RECT 476.400 22.050 477.450 43.950 ;
        RECT 479.400 40.050 480.450 52.950 ;
        RECT 485.400 40.050 486.450 52.950 ;
        RECT 491.400 52.050 492.450 52.950 ;
        RECT 497.400 52.050 498.450 55.950 ;
        RECT 500.400 55.050 501.450 55.950 ;
        RECT 499.950 52.950 502.050 55.050 ;
        RECT 505.950 52.950 508.050 55.050 ;
        RECT 509.250 53.250 511.050 54.150 ;
        RECT 487.950 49.950 490.050 52.050 ;
        RECT 490.950 49.950 493.050 52.050 ;
        RECT 496.950 49.950 499.050 52.050 ;
        RECT 499.950 50.850 502.050 51.750 ;
        RECT 502.950 50.250 505.050 51.150 ;
        RECT 505.950 50.850 507.750 51.750 ;
        RECT 508.950 49.950 511.050 52.050 ;
        RECT 488.400 49.050 489.450 49.950 ;
        RECT 487.950 46.950 490.050 49.050 ;
        RECT 502.950 46.950 505.050 49.050 ;
        RECT 509.400 40.050 510.450 49.950 ;
        RECT 478.950 37.950 481.050 40.050 ;
        RECT 484.950 37.950 487.050 40.050 ;
        RECT 508.950 37.950 511.050 40.050 ;
        RECT 512.400 34.050 513.450 55.950 ;
        RECT 514.950 52.950 517.050 55.050 ;
        RECT 515.400 46.050 516.450 52.950 ;
        RECT 518.400 49.050 519.450 55.950 ;
        RECT 520.950 52.950 523.050 55.050 ;
        RECT 524.250 53.850 526.050 54.750 ;
        RECT 526.950 52.950 529.050 55.050 ;
        RECT 529.950 53.250 531.750 54.150 ;
        RECT 532.950 52.950 535.050 55.050 ;
        RECT 536.250 53.250 537.750 54.150 ;
        RECT 538.950 52.950 541.050 55.050 ;
        RECT 521.400 52.050 522.450 52.950 ;
        RECT 520.950 49.950 523.050 52.050 ;
        RECT 517.950 46.950 520.050 49.050 ;
        RECT 514.950 43.950 517.050 46.050 ;
        RECT 527.400 40.050 528.450 52.950 ;
        RECT 542.400 52.050 543.450 76.950 ;
        RECT 545.400 64.050 546.450 85.950 ;
        RECT 548.400 64.050 549.450 98.400 ;
        RECT 551.400 97.050 552.450 103.950 ;
        RECT 572.400 100.050 573.450 127.950 ;
        RECT 581.400 127.050 582.450 163.950 ;
        RECT 590.400 163.050 591.450 175.950 ;
        RECT 592.950 172.950 595.050 175.050 ;
        RECT 593.400 166.050 594.450 172.950 ;
        RECT 599.400 172.050 600.450 175.950 ;
        RECT 602.400 172.050 603.450 181.950 ;
        RECT 598.950 169.950 601.050 172.050 ;
        RECT 601.950 169.950 604.050 172.050 ;
        RECT 595.950 167.250 598.050 168.150 ;
        RECT 598.950 167.850 601.050 168.750 ;
        RECT 601.950 167.250 603.750 168.150 ;
        RECT 604.950 166.950 607.050 169.050 ;
        RECT 608.400 166.050 609.450 202.950 ;
        RECT 611.400 202.050 612.450 214.950 ;
        RECT 613.950 202.950 616.050 205.050 ;
        RECT 610.950 199.950 613.050 202.050 ;
        RECT 614.400 201.450 615.450 202.950 ;
        RECT 617.400 201.450 618.450 253.950 ;
        RECT 626.400 250.050 627.450 265.950 ;
        RECT 629.400 262.050 630.450 268.950 ;
        RECT 635.400 267.450 636.450 295.950 ;
        RECT 637.950 292.950 640.050 295.050 ;
        RECT 632.400 266.400 636.450 267.450 ;
        RECT 628.950 259.950 631.050 262.050 ;
        RECT 628.950 256.950 631.050 259.050 ;
        RECT 619.950 247.950 622.050 250.050 ;
        RECT 625.950 247.950 628.050 250.050 ;
        RECT 620.400 244.050 621.450 247.950 ;
        RECT 622.950 244.950 625.050 247.050 ;
        RECT 619.950 241.950 622.050 244.050 ;
        RECT 619.950 239.250 622.050 240.150 ;
        RECT 619.950 235.950 622.050 238.050 ;
        RECT 619.950 232.950 622.050 235.050 ;
        RECT 620.400 205.050 621.450 232.950 ;
        RECT 619.950 202.950 622.050 205.050 ;
        RECT 614.400 200.400 618.450 201.450 ;
        RECT 614.400 199.050 615.450 200.400 ;
        RECT 619.950 200.250 622.050 201.150 ;
        RECT 610.950 197.250 612.750 198.150 ;
        RECT 613.950 196.950 616.050 199.050 ;
        RECT 617.250 197.250 618.750 198.150 ;
        RECT 619.950 196.950 622.050 199.050 ;
        RECT 610.950 193.950 613.050 196.050 ;
        RECT 614.250 194.850 615.750 195.750 ;
        RECT 616.950 193.950 619.050 196.050 ;
        RECT 611.400 193.050 612.450 193.950 ;
        RECT 610.950 190.950 613.050 193.050 ;
        RECT 611.400 169.050 612.450 190.950 ;
        RECT 617.400 184.050 618.450 193.950 ;
        RECT 616.950 181.950 619.050 184.050 ;
        RECT 620.400 178.050 621.450 196.950 ;
        RECT 619.950 175.950 622.050 178.050 ;
        RECT 616.950 172.950 619.050 175.050 ;
        RECT 617.400 169.050 618.450 172.950 ;
        RECT 619.950 169.950 622.050 172.050 ;
        RECT 610.950 166.950 613.050 169.050 ;
        RECT 614.250 167.250 615.750 168.150 ;
        RECT 616.950 166.950 619.050 169.050 ;
        RECT 620.400 166.050 621.450 169.950 ;
        RECT 592.950 165.450 595.050 166.050 ;
        RECT 595.950 165.450 598.050 166.050 ;
        RECT 592.950 164.400 598.050 165.450 ;
        RECT 592.950 163.950 595.050 164.400 ;
        RECT 595.950 163.950 598.050 164.400 ;
        RECT 598.950 163.950 601.050 166.050 ;
        RECT 601.950 163.950 604.050 166.050 ;
        RECT 605.250 164.850 607.050 165.750 ;
        RECT 607.950 163.950 610.050 166.050 ;
        RECT 610.950 164.850 612.750 165.750 ;
        RECT 613.950 163.950 616.050 166.050 ;
        RECT 617.250 164.850 618.750 165.750 ;
        RECT 619.950 163.950 622.050 166.050 ;
        RECT 583.950 160.950 586.050 163.050 ;
        RECT 587.250 161.850 588.750 162.750 ;
        RECT 589.950 160.950 592.050 163.050 ;
        RECT 593.250 161.850 595.050 162.750 ;
        RECT 584.400 145.050 585.450 160.950 ;
        RECT 589.950 158.850 592.050 159.750 ;
        RECT 592.950 154.950 595.050 157.050 ;
        RECT 595.950 154.950 598.050 157.050 ;
        RECT 583.950 142.950 586.050 145.050 ;
        RECT 583.950 139.950 586.050 142.050 ;
        RECT 589.950 139.950 592.050 142.050 ;
        RECT 574.950 124.950 577.050 127.050 ;
        RECT 578.250 125.850 580.050 126.750 ;
        RECT 580.950 124.950 583.050 127.050 ;
        RECT 584.400 123.450 585.450 139.950 ;
        RECT 590.400 136.050 591.450 139.950 ;
        RECT 593.400 136.050 594.450 154.950 ;
        RECT 596.400 145.050 597.450 154.950 ;
        RECT 599.400 151.050 600.450 163.950 ;
        RECT 613.950 160.950 616.050 163.050 ;
        RECT 616.950 160.950 619.050 163.050 ;
        RECT 619.950 161.850 622.050 162.750 ;
        RECT 598.950 148.950 601.050 151.050 ;
        RECT 607.950 148.950 610.050 151.050 ;
        RECT 595.950 142.950 598.050 145.050 ;
        RECT 589.950 133.950 592.050 136.050 ;
        RECT 592.950 133.950 595.050 136.050 ;
        RECT 589.950 127.950 592.050 130.050 ;
        RECT 590.400 127.050 591.450 127.950 ;
        RECT 596.400 127.050 597.450 142.950 ;
        RECT 608.400 133.050 609.450 148.950 ;
        RECT 614.400 148.050 615.450 160.950 ;
        RECT 613.950 145.950 616.050 148.050 ;
        RECT 613.950 139.950 616.050 142.050 ;
        RECT 604.950 131.250 607.050 132.150 ;
        RECT 607.950 130.950 610.050 133.050 ;
        RECT 601.950 128.250 603.750 129.150 ;
        RECT 604.950 127.950 607.050 130.050 ;
        RECT 608.250 128.250 609.750 129.150 ;
        RECT 610.950 127.950 613.050 130.050 ;
        RECT 586.950 125.250 588.750 126.150 ;
        RECT 589.950 124.950 592.050 127.050 ;
        RECT 593.250 125.250 594.750 126.150 ;
        RECT 595.950 124.950 598.050 127.050 ;
        RECT 599.250 125.250 601.050 126.150 ;
        RECT 601.950 124.950 604.050 127.050 ;
        RECT 581.400 122.400 585.450 123.450 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 556.950 97.950 559.050 100.050 ;
        RECT 565.950 97.950 568.050 100.050 ;
        RECT 571.950 97.950 574.050 100.050 ;
        RECT 550.950 94.950 553.050 97.050 ;
        RECT 554.250 95.250 556.050 96.150 ;
        RECT 556.950 95.850 559.050 96.750 ;
        RECT 559.950 95.250 562.050 96.150 ;
        RECT 562.950 94.950 565.050 97.050 ;
        RECT 563.400 94.050 564.450 94.950 ;
        RECT 550.950 92.850 552.750 93.750 ;
        RECT 553.950 91.950 556.050 94.050 ;
        RECT 559.950 91.950 562.050 94.050 ;
        RECT 562.950 91.950 565.050 94.050 ;
        RECT 544.950 61.950 547.050 64.050 ;
        RECT 547.950 61.950 550.050 64.050 ;
        RECT 547.950 59.250 550.050 60.150 ;
        RECT 560.400 58.050 561.450 91.950 ;
        RECT 566.400 91.050 567.450 97.950 ;
        RECT 568.950 91.950 571.050 94.050 ;
        RECT 572.250 92.250 574.050 93.150 ;
        RECT 562.950 89.850 564.750 90.750 ;
        RECT 565.950 88.950 568.050 91.050 ;
        RECT 569.250 89.850 570.750 90.750 ;
        RECT 571.950 88.950 574.050 91.050 ;
        RECT 562.950 85.950 565.050 88.050 ;
        RECT 565.950 86.850 568.050 87.750 ;
        RECT 563.400 58.050 564.450 85.950 ;
        RECT 572.400 76.050 573.450 88.950 ;
        RECT 571.950 73.950 574.050 76.050 ;
        RECT 571.950 64.950 574.050 67.050 ;
        RECT 544.950 56.250 546.750 57.150 ;
        RECT 547.950 55.950 550.050 58.050 ;
        RECT 551.250 56.250 552.750 57.150 ;
        RECT 553.950 55.950 556.050 58.050 ;
        RECT 559.950 55.950 562.050 58.050 ;
        RECT 562.950 55.950 565.050 58.050 ;
        RECT 568.950 56.250 571.050 57.150 ;
        RECT 544.950 52.950 547.050 55.050 ;
        RECT 548.400 52.050 549.450 55.950 ;
        RECT 550.950 52.950 553.050 55.050 ;
        RECT 554.250 53.850 556.050 54.750 ;
        RECT 556.950 52.950 559.050 55.050 ;
        RECT 559.950 53.250 561.750 54.150 ;
        RECT 562.950 52.950 565.050 55.050 ;
        RECT 568.950 54.450 571.050 55.050 ;
        RECT 572.400 54.450 573.450 64.950 ;
        RECT 566.250 53.250 567.750 54.150 ;
        RECT 568.950 53.400 573.450 54.450 ;
        RECT 568.950 52.950 571.050 53.400 ;
        RECT 529.950 49.950 532.050 52.050 ;
        RECT 533.250 50.850 534.750 51.750 ;
        RECT 535.950 51.450 538.050 52.050 ;
        RECT 538.950 51.450 541.050 52.050 ;
        RECT 535.950 50.400 541.050 51.450 ;
        RECT 535.950 49.950 538.050 50.400 ;
        RECT 538.950 49.950 541.050 50.400 ;
        RECT 541.950 49.950 544.050 52.050 ;
        RECT 547.950 49.950 550.050 52.050 ;
        RECT 530.400 46.050 531.450 49.950 ;
        RECT 551.400 49.050 552.450 52.950 ;
        RECT 550.950 46.950 553.050 49.050 ;
        RECT 529.950 43.950 532.050 46.050 ;
        RECT 530.400 43.050 531.450 43.950 ;
        RECT 551.400 43.050 552.450 46.950 ;
        RECT 529.950 40.950 532.050 43.050 ;
        RECT 550.950 40.950 553.050 43.050 ;
        RECT 557.400 40.050 558.450 52.950 ;
        RECT 559.950 49.950 562.050 52.050 ;
        RECT 563.250 50.850 564.750 51.750 ;
        RECT 565.950 49.950 568.050 52.050 ;
        RECT 560.400 46.050 561.450 49.950 ;
        RECT 562.950 46.950 565.050 49.050 ;
        RECT 559.950 43.950 562.050 46.050 ;
        RECT 526.950 37.950 529.050 40.050 ;
        RECT 556.950 37.950 559.050 40.050 ;
        RECT 535.950 34.950 538.050 37.050 ;
        RECT 487.950 31.950 490.050 34.050 ;
        RECT 511.950 31.950 514.050 34.050 ;
        RECT 529.950 31.950 532.050 34.050 ;
        RECT 481.950 25.950 484.050 28.050 ;
        RECT 433.950 20.400 438.450 21.450 ;
        RECT 439.950 20.850 442.050 21.750 ;
        RECT 433.950 19.950 436.050 20.400 ;
        RECT 442.950 20.250 445.050 21.150 ;
        RECT 448.950 20.850 451.050 21.750 ;
        RECT 451.950 19.950 454.050 22.050 ;
        RECT 457.950 20.850 459.750 21.750 ;
        RECT 460.950 19.950 463.050 22.050 ;
        RECT 464.250 20.850 465.750 21.750 ;
        RECT 466.950 19.950 469.050 22.050 ;
        RECT 470.250 20.850 472.050 21.750 ;
        RECT 472.950 20.250 474.750 21.150 ;
        RECT 475.950 19.950 478.050 22.050 ;
        RECT 479.250 20.250 481.050 21.150 ;
        RECT 407.400 19.050 408.450 19.950 ;
        RECT 467.400 19.050 468.450 19.950 ;
        RECT 482.400 19.050 483.450 25.950 ;
        RECT 488.400 22.050 489.450 31.950 ;
        RECT 508.950 28.950 511.050 31.050 ;
        RECT 526.950 28.950 529.050 31.050 ;
        RECT 496.950 25.950 499.050 28.050 ;
        RECT 497.400 25.050 498.450 25.950 ;
        RECT 490.950 22.950 493.050 25.050 ;
        RECT 494.250 23.250 495.750 24.150 ;
        RECT 496.950 22.950 499.050 25.050 ;
        RECT 502.950 22.950 505.050 25.050 ;
        RECT 487.950 19.950 490.050 22.050 ;
        RECT 491.250 20.850 492.750 21.750 ;
        RECT 493.950 19.950 496.050 22.050 ;
        RECT 497.250 20.850 499.050 21.750 ;
        RECT 502.950 20.850 505.050 21.750 ;
        RECT 505.950 20.250 508.050 21.150 ;
        RECT 337.950 17.400 342.450 18.450 ;
        RECT 346.950 17.850 349.050 18.750 ;
        RECT 337.950 16.950 340.050 17.400 ;
        RECT 352.950 16.950 355.050 19.050 ;
        RECT 367.950 17.850 370.050 18.750 ;
        RECT 382.950 16.950 385.050 19.050 ;
        RECT 406.950 16.950 409.050 19.050 ;
        RECT 412.950 17.850 415.050 18.750 ;
        RECT 442.950 16.950 445.050 19.050 ;
        RECT 466.950 16.950 469.050 19.050 ;
        RECT 472.950 16.950 475.050 19.050 ;
        RECT 476.250 17.850 477.750 18.750 ;
        RECT 478.950 16.950 481.050 19.050 ;
        RECT 481.950 16.950 484.050 19.050 ;
        RECT 487.950 17.850 490.050 18.750 ;
        RECT 505.950 18.450 508.050 19.050 ;
        RECT 509.400 18.450 510.450 28.950 ;
        RECT 517.950 25.950 520.050 28.050 ;
        RECT 523.950 25.950 526.050 28.050 ;
        RECT 511.950 22.950 514.050 25.050 ;
        RECT 518.400 22.050 519.450 25.950 ;
        RECT 527.400 25.050 528.450 28.950 ;
        RECT 530.400 25.050 531.450 31.950 ;
        RECT 536.400 25.050 537.450 34.950 ;
        RECT 547.950 31.950 550.050 34.050 ;
        RECT 548.400 28.050 549.450 31.950 ;
        RECT 538.950 25.950 541.050 28.050 ;
        RECT 547.950 25.950 550.050 28.050 ;
        RECT 559.950 25.950 562.050 28.050 ;
        RECT 520.950 22.950 523.050 25.050 ;
        RECT 524.250 23.850 525.750 24.750 ;
        RECT 526.950 22.950 529.050 25.050 ;
        RECT 529.950 22.950 532.050 25.050 ;
        RECT 533.250 23.250 534.750 24.150 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 539.400 22.050 540.450 25.950 ;
        RECT 547.950 23.850 550.050 24.750 ;
        RECT 560.400 24.450 561.450 25.950 ;
        RECT 563.400 24.450 564.450 46.950 ;
        RECT 569.400 37.050 570.450 52.950 ;
        RECT 575.400 52.050 576.450 100.950 ;
        RECT 581.400 100.050 582.450 122.400 ;
        RECT 586.950 121.950 589.050 124.050 ;
        RECT 590.250 122.850 591.750 123.750 ;
        RECT 592.950 121.950 595.050 124.050 ;
        RECT 596.250 122.850 597.750 123.750 ;
        RECT 598.950 121.950 601.050 124.050 ;
        RECT 601.950 121.950 604.050 124.050 ;
        RECT 583.950 118.950 586.050 121.050 ;
        RECT 577.950 97.950 580.050 100.050 ;
        RECT 580.950 97.950 583.050 100.050 ;
        RECT 577.950 95.850 580.050 96.750 ;
        RECT 580.950 95.250 583.050 96.150 ;
        RECT 580.950 93.450 583.050 94.050 ;
        RECT 584.400 93.450 585.450 118.950 ;
        RECT 587.400 112.050 588.450 121.950 ;
        RECT 586.950 109.950 589.050 112.050 ;
        RECT 593.400 103.050 594.450 121.950 ;
        RECT 592.950 100.950 595.050 103.050 ;
        RECT 589.950 99.450 592.050 100.050 ;
        RECT 580.950 92.400 585.450 93.450 ;
        RECT 587.400 98.400 592.050 99.450 ;
        RECT 580.950 91.950 583.050 92.400 ;
        RECT 587.400 85.050 588.450 98.400 ;
        RECT 589.950 97.950 592.050 98.400 ;
        RECT 598.950 97.950 601.050 100.050 ;
        RECT 589.950 95.850 592.050 96.750 ;
        RECT 592.950 95.250 595.050 96.150 ;
        RECT 595.950 94.950 598.050 97.050 ;
        RECT 592.950 91.950 595.050 94.050 ;
        RECT 596.400 91.050 597.450 94.950 ;
        RECT 595.950 88.950 598.050 91.050 ;
        RECT 599.400 88.050 600.450 97.950 ;
        RECT 598.950 85.950 601.050 88.050 ;
        RECT 586.950 82.950 589.050 85.050 ;
        RECT 587.400 67.050 588.450 82.950 ;
        RECT 586.950 64.950 589.050 67.050 ;
        RECT 583.950 61.950 586.050 64.050 ;
        RECT 584.400 61.050 585.450 61.950 ;
        RECT 583.950 58.950 586.050 61.050 ;
        RECT 586.950 58.950 589.050 61.050 ;
        RECT 584.400 58.050 585.450 58.950 ;
        RECT 577.950 55.950 580.050 58.050 ;
        RECT 581.250 56.250 582.750 57.150 ;
        RECT 583.950 55.950 586.050 58.050 ;
        RECT 577.950 53.850 579.750 54.750 ;
        RECT 580.950 52.950 583.050 55.050 ;
        RECT 584.250 53.850 586.050 54.750 ;
        RECT 571.950 49.950 574.050 52.050 ;
        RECT 574.950 49.950 577.050 52.050 ;
        RECT 572.400 46.050 573.450 49.950 ;
        RECT 581.400 49.050 582.450 52.950 ;
        RECT 587.400 51.450 588.450 58.950 ;
        RECT 589.950 53.250 592.050 54.150 ;
        RECT 595.950 53.250 598.050 54.150 ;
        RECT 589.950 51.450 592.050 52.050 ;
        RECT 587.400 50.400 592.050 51.450 ;
        RECT 589.950 49.950 592.050 50.400 ;
        RECT 593.250 50.250 594.750 51.150 ;
        RECT 595.950 49.950 598.050 52.050 ;
        RECT 596.400 49.050 597.450 49.950 ;
        RECT 580.950 46.950 583.050 49.050 ;
        RECT 586.950 46.950 589.050 49.050 ;
        RECT 592.950 46.950 595.050 49.050 ;
        RECT 595.950 46.950 598.050 49.050 ;
        RECT 571.950 43.950 574.050 46.050 ;
        RECT 580.950 43.950 583.050 46.050 ;
        RECT 568.950 34.950 571.050 37.050 ;
        RECT 581.400 31.050 582.450 43.950 ;
        RECT 580.950 28.950 583.050 31.050 ;
        RECT 581.400 25.050 582.450 28.950 ;
        RECT 583.950 27.450 586.050 28.050 ;
        RECT 587.400 27.450 588.450 46.950 ;
        RECT 593.400 46.050 594.450 46.950 ;
        RECT 602.400 46.050 603.450 121.950 ;
        RECT 605.400 112.050 606.450 127.950 ;
        RECT 607.950 124.950 610.050 127.050 ;
        RECT 611.250 125.850 613.050 126.750 ;
        RECT 608.400 121.050 609.450 124.950 ;
        RECT 610.950 121.950 613.050 124.050 ;
        RECT 607.950 118.950 610.050 121.050 ;
        RECT 604.950 109.950 607.050 112.050 ;
        RECT 611.400 106.050 612.450 121.950 ;
        RECT 610.950 103.950 613.050 106.050 ;
        RECT 614.400 99.450 615.450 139.950 ;
        RECT 617.400 133.050 618.450 160.950 ;
        RECT 623.400 133.050 624.450 244.950 ;
        RECT 625.950 241.950 628.050 244.050 ;
        RECT 626.400 208.050 627.450 241.950 ;
        RECT 629.400 232.050 630.450 256.950 ;
        RECT 632.400 241.050 633.450 266.400 ;
        RECT 638.400 250.050 639.450 292.950 ;
        RECT 641.400 262.050 642.450 295.950 ;
        RECT 644.400 292.050 645.450 301.950 ;
        RECT 643.950 289.950 646.050 292.050 ;
        RECT 653.400 289.050 654.450 331.950 ;
        RECT 656.400 313.050 657.450 335.400 ;
        RECT 661.950 334.950 664.050 337.050 ;
        RECT 667.950 334.950 670.050 337.050 ;
        RECT 670.950 334.950 673.050 337.050 ;
        RECT 658.950 322.950 661.050 325.050 ;
        RECT 655.950 310.950 658.050 313.050 ;
        RECT 659.400 310.050 660.450 322.950 ;
        RECT 668.400 316.050 669.450 334.950 ;
        RECT 677.400 334.050 678.450 343.950 ;
        RECT 679.950 340.950 682.050 343.050 ;
        RECT 680.400 340.050 681.450 340.950 ;
        RECT 679.950 337.950 682.050 340.050 ;
        RECT 676.950 331.950 679.050 334.050 ;
        RECT 670.950 328.950 673.050 331.050 ;
        RECT 664.950 313.950 667.050 316.050 ;
        RECT 667.950 313.950 670.050 316.050 ;
        RECT 661.950 310.950 664.050 313.050 ;
        RECT 655.950 308.250 657.750 309.150 ;
        RECT 658.950 307.950 661.050 310.050 ;
        RECT 662.400 307.050 663.450 310.950 ;
        RECT 665.400 310.050 666.450 313.950 ;
        RECT 671.400 313.050 672.450 328.950 ;
        RECT 676.950 313.950 679.050 316.050 ;
        RECT 667.950 310.950 670.050 313.050 ;
        RECT 670.950 310.950 673.050 313.050 ;
        RECT 674.250 311.250 676.050 312.150 ;
        RECT 676.950 311.850 679.050 312.750 ;
        RECT 679.950 311.250 682.050 312.150 ;
        RECT 664.950 307.950 667.050 310.050 ;
        RECT 655.950 304.950 658.050 307.050 ;
        RECT 659.250 305.850 660.750 306.750 ;
        RECT 661.950 304.950 664.050 307.050 ;
        RECT 665.250 305.850 667.050 306.750 ;
        RECT 661.950 302.850 664.050 303.750 ;
        RECT 664.950 298.950 667.050 301.050 ;
        RECT 646.950 286.950 649.050 289.050 ;
        RECT 652.950 286.950 655.050 289.050 ;
        RECT 643.950 283.950 646.050 286.050 ;
        RECT 644.400 283.050 645.450 283.950 ;
        RECT 643.950 280.950 646.050 283.050 ;
        RECT 644.400 274.050 645.450 280.950 ;
        RECT 647.400 276.450 648.450 286.950 ;
        RECT 665.400 286.050 666.450 298.950 ;
        RECT 664.950 283.950 667.050 286.050 ;
        RECT 655.950 280.950 658.050 283.050 ;
        RECT 652.950 277.950 655.050 280.050 ;
        RECT 647.400 275.400 651.450 276.450 ;
        RECT 650.400 274.050 651.450 275.400 ;
        RECT 653.400 274.050 654.450 277.950 ;
        RECT 643.950 271.950 646.050 274.050 ;
        RECT 647.250 272.250 648.750 273.150 ;
        RECT 649.950 271.950 652.050 274.050 ;
        RECT 652.950 271.950 655.050 274.050 ;
        RECT 656.400 271.050 657.450 280.950 ;
        RECT 668.400 279.450 669.450 310.950 ;
        RECT 670.950 308.850 672.750 309.750 ;
        RECT 673.950 307.950 676.050 310.050 ;
        RECT 679.950 307.950 682.050 310.050 ;
        RECT 680.400 307.050 681.450 307.950 ;
        RECT 670.950 304.950 673.050 307.050 ;
        RECT 679.950 304.950 682.050 307.050 ;
        RECT 671.400 301.050 672.450 304.950 ;
        RECT 676.950 301.950 679.050 304.050 ;
        RECT 670.950 298.950 673.050 301.050 ;
        RECT 673.950 286.950 676.050 289.050 ;
        RECT 665.400 278.400 669.450 279.450 ;
        RECT 661.950 272.250 664.050 273.150 ;
        RECT 643.950 269.850 645.750 270.750 ;
        RECT 646.950 268.950 649.050 271.050 ;
        RECT 650.250 269.850 652.050 270.750 ;
        RECT 652.950 269.250 654.750 270.150 ;
        RECT 655.950 268.950 658.050 271.050 ;
        RECT 659.250 269.250 660.750 270.150 ;
        RECT 661.950 268.950 664.050 271.050 ;
        RECT 643.950 265.950 646.050 268.050 ;
        RECT 640.950 259.950 643.050 262.050 ;
        RECT 644.400 259.050 645.450 265.950 ;
        RECT 647.400 265.050 648.450 268.950 ;
        RECT 649.950 265.950 652.050 268.050 ;
        RECT 652.950 265.950 655.050 268.050 ;
        RECT 656.250 266.850 657.750 267.750 ;
        RECT 658.950 265.950 661.050 268.050 ;
        RECT 661.950 265.950 664.050 268.050 ;
        RECT 646.950 262.950 649.050 265.050 ;
        RECT 643.950 256.950 646.050 259.050 ;
        RECT 637.950 247.950 640.050 250.050 ;
        RECT 637.950 244.950 640.050 247.050 ;
        RECT 643.950 244.950 646.050 247.050 ;
        RECT 638.400 244.050 639.450 244.950 ;
        RECT 637.950 241.950 640.050 244.050 ;
        RECT 631.950 238.950 634.050 241.050 ;
        RECT 635.250 239.250 637.050 240.150 ;
        RECT 637.950 239.850 640.050 240.750 ;
        RECT 640.950 239.250 643.050 240.150 ;
        RECT 631.950 236.850 633.750 237.750 ;
        RECT 634.950 235.950 637.050 238.050 ;
        RECT 640.950 235.950 643.050 238.050 ;
        RECT 628.950 229.950 631.050 232.050 ;
        RECT 631.950 226.950 634.050 229.050 ;
        RECT 632.400 210.450 633.450 226.950 ;
        RECT 635.400 226.050 636.450 235.950 ;
        RECT 637.950 229.950 640.050 232.050 ;
        RECT 634.950 223.950 637.050 226.050 ;
        RECT 638.400 223.050 639.450 229.950 ;
        RECT 641.400 223.050 642.450 235.950 ;
        RECT 637.950 220.950 640.050 223.050 ;
        RECT 640.950 220.950 643.050 223.050 ;
        RECT 632.400 209.400 636.450 210.450 ;
        RECT 625.950 205.950 628.050 208.050 ;
        RECT 631.950 205.950 634.050 208.050 ;
        RECT 628.950 196.950 631.050 199.050 ;
        RECT 625.950 194.250 628.050 195.150 ;
        RECT 628.950 194.850 631.050 195.750 ;
        RECT 632.400 195.450 633.450 205.950 ;
        RECT 635.400 205.050 636.450 209.400 ;
        RECT 638.400 205.050 639.450 220.950 ;
        RECT 640.950 208.950 643.050 211.050 ;
        RECT 634.950 202.950 637.050 205.050 ;
        RECT 637.950 202.950 640.050 205.050 ;
        RECT 641.400 204.450 642.450 208.950 ;
        RECT 644.400 208.050 645.450 244.950 ;
        RECT 650.400 244.050 651.450 265.950 ;
        RECT 653.400 256.050 654.450 265.950 ;
        RECT 652.950 253.950 655.050 256.050 ;
        RECT 659.400 255.450 660.450 265.950 ;
        RECT 662.400 262.050 663.450 265.950 ;
        RECT 661.950 259.950 664.050 262.050 ;
        RECT 656.400 254.400 660.450 255.450 ;
        RECT 656.400 244.050 657.450 254.400 ;
        RECT 658.950 250.950 661.050 253.050 ;
        RECT 649.950 241.950 652.050 244.050 ;
        RECT 655.950 241.950 658.050 244.050 ;
        RECT 655.950 238.950 658.050 241.050 ;
        RECT 646.950 236.250 648.750 237.150 ;
        RECT 649.950 235.950 652.050 238.050 ;
        RECT 653.250 236.250 655.050 237.150 ;
        RECT 655.950 236.850 658.050 237.750 ;
        RECT 646.950 232.950 649.050 235.050 ;
        RECT 650.250 233.850 651.750 234.750 ;
        RECT 652.950 232.950 655.050 235.050 ;
        RECT 659.400 234.450 660.450 250.950 ;
        RECT 665.400 249.450 666.450 278.400 ;
        RECT 667.950 274.950 670.050 277.050 ;
        RECT 668.400 274.050 669.450 274.950 ;
        RECT 667.950 271.950 670.050 274.050 ;
        RECT 670.950 268.950 673.050 271.050 ;
        RECT 667.950 266.250 670.050 267.150 ;
        RECT 670.950 266.850 673.050 267.750 ;
        RECT 667.950 262.950 670.050 265.050 ;
        RECT 670.950 262.950 673.050 265.050 ;
        RECT 671.400 259.050 672.450 262.950 ;
        RECT 670.950 256.950 673.050 259.050 ;
        RECT 671.400 253.050 672.450 256.950 ;
        RECT 674.400 253.050 675.450 286.950 ;
        RECT 670.950 250.950 673.050 253.050 ;
        RECT 673.950 250.950 676.050 253.050 ;
        RECT 662.400 248.400 666.450 249.450 ;
        RECT 662.400 241.050 663.450 248.400 ;
        RECT 677.400 247.050 678.450 301.950 ;
        RECT 680.400 295.050 681.450 304.950 ;
        RECT 683.400 298.050 684.450 385.950 ;
        RECT 686.400 385.050 687.450 394.950 ;
        RECT 689.400 388.050 690.450 403.950 ;
        RECT 695.400 391.050 696.450 407.400 ;
        RECT 697.950 406.950 700.050 409.050 ;
        RECT 698.400 402.450 699.450 406.950 ;
        RECT 701.400 406.050 702.450 412.950 ;
        RECT 703.950 406.950 706.050 409.050 ;
        RECT 700.950 403.950 703.050 406.050 ;
        RECT 698.400 401.400 702.450 402.450 ;
        RECT 697.950 394.950 700.050 397.050 ;
        RECT 694.950 388.950 697.050 391.050 ;
        RECT 688.950 385.950 691.050 388.050 ;
        RECT 691.950 385.950 694.050 388.050 ;
        RECT 685.950 382.950 688.050 385.050 ;
        RECT 689.250 383.250 691.050 384.150 ;
        RECT 691.950 383.850 694.050 384.750 ;
        RECT 694.950 383.250 697.050 384.150 ;
        RECT 685.950 380.850 687.750 381.750 ;
        RECT 688.950 379.950 691.050 382.050 ;
        RECT 694.950 379.950 697.050 382.050 ;
        RECT 685.950 373.950 688.050 376.050 ;
        RECT 686.400 331.050 687.450 373.950 ;
        RECT 689.400 367.050 690.450 379.950 ;
        RECT 695.400 379.050 696.450 379.950 ;
        RECT 691.950 376.950 694.050 379.050 ;
        RECT 694.950 376.950 697.050 379.050 ;
        RECT 692.400 370.050 693.450 376.950 ;
        RECT 695.400 376.050 696.450 376.950 ;
        RECT 694.950 373.950 697.050 376.050 ;
        RECT 691.950 367.950 694.050 370.050 ;
        RECT 688.950 364.950 691.050 367.050 ;
        RECT 698.400 349.050 699.450 394.950 ;
        RECT 701.400 391.050 702.450 401.400 ;
        RECT 700.950 388.950 703.050 391.050 ;
        RECT 704.400 387.450 705.450 406.950 ;
        RECT 707.400 406.050 708.450 439.950 ;
        RECT 719.400 439.050 720.450 445.950 ;
        RECT 718.950 436.950 721.050 439.050 ;
        RECT 712.950 433.950 715.050 436.050 ;
        RECT 713.400 417.450 714.450 433.950 ;
        RECT 715.950 430.950 718.050 433.050 ;
        RECT 716.400 418.050 717.450 430.950 ;
        RECT 718.950 424.950 721.050 427.050 ;
        RECT 721.950 424.950 724.050 427.050 ;
        RECT 710.400 416.400 714.450 417.450 ;
        RECT 706.950 403.950 709.050 406.050 ;
        RECT 710.400 396.450 711.450 416.400 ;
        RECT 715.950 415.950 718.050 418.050 ;
        RECT 716.400 415.050 717.450 415.950 ;
        RECT 719.400 415.050 720.450 424.950 ;
        RECT 722.400 415.050 723.450 424.950 ;
        RECT 725.400 421.050 726.450 449.400 ;
        RECT 727.950 445.950 730.050 448.050 ;
        RECT 728.400 433.050 729.450 445.950 ;
        RECT 731.400 439.050 732.450 455.400 ;
        RECT 736.950 454.950 739.050 457.050 ;
        RECT 742.950 455.250 745.050 456.150 ;
        RECT 733.950 451.950 736.050 454.050 ;
        RECT 736.950 452.850 739.050 453.750 ;
        RECT 742.950 451.950 745.050 454.050 ;
        RECT 730.950 436.950 733.050 439.050 ;
        RECT 734.400 436.050 735.450 451.950 ;
        RECT 733.950 433.950 736.050 436.050 ;
        RECT 739.950 433.950 742.050 436.050 ;
        RECT 727.950 430.950 730.050 433.050 ;
        RECT 733.950 421.950 736.050 424.050 ;
        RECT 724.950 418.950 727.050 421.050 ;
        RECT 727.950 419.250 730.050 420.150 ;
        RECT 734.400 418.050 735.450 421.950 ;
        RECT 740.400 421.050 741.450 433.950 ;
        RECT 743.400 424.050 744.450 451.950 ;
        RECT 742.950 421.950 745.050 424.050 ;
        RECT 746.400 421.050 747.450 520.950 ;
        RECT 751.950 517.950 754.050 520.050 ;
        RECT 752.400 487.050 753.450 517.950 ;
        RECT 758.400 514.050 759.450 593.400 ;
        RECT 760.950 589.950 763.050 592.050 ;
        RECT 761.400 586.050 762.450 589.950 ;
        RECT 760.950 583.950 763.050 586.050 ;
        RECT 760.950 574.950 763.050 577.050 ;
        RECT 761.400 529.050 762.450 574.950 ;
        RECT 760.950 526.950 763.050 529.050 ;
        RECT 760.950 524.850 763.050 525.750 ;
        RECT 764.400 517.050 765.450 601.950 ;
        RECT 767.400 547.050 768.450 620.400 ;
        RECT 770.400 613.050 771.450 634.950 ;
        RECT 769.950 610.950 772.050 613.050 ;
        RECT 769.950 604.950 772.050 607.050 ;
        RECT 770.400 589.050 771.450 604.950 ;
        RECT 769.950 586.950 772.050 589.050 ;
        RECT 769.950 583.950 772.050 586.050 ;
        RECT 766.950 544.950 769.050 547.050 ;
        RECT 770.400 520.050 771.450 583.950 ;
        RECT 769.950 517.950 772.050 520.050 ;
        RECT 763.950 514.950 766.050 517.050 ;
        RECT 757.950 511.950 760.050 514.050 ;
        RECT 769.950 496.950 772.050 499.050 ;
        RECT 766.950 490.950 769.050 493.050 ;
        RECT 760.950 489.450 763.050 490.050 ;
        RECT 758.400 488.400 763.050 489.450 ;
        RECT 748.950 485.250 751.050 486.150 ;
        RECT 751.950 484.950 754.050 487.050 ;
        RECT 754.950 485.250 757.050 486.150 ;
        RECT 758.400 484.050 759.450 488.400 ;
        RECT 760.950 487.950 763.050 488.400 ;
        RECT 760.950 485.850 763.050 486.750 ;
        RECT 763.950 485.250 766.050 486.150 ;
        RECT 748.950 481.950 751.050 484.050 ;
        RECT 752.250 482.250 754.050 483.150 ;
        RECT 754.950 481.950 757.050 484.050 ;
        RECT 757.950 481.950 760.050 484.050 ;
        RECT 760.950 481.950 763.050 484.050 ;
        RECT 763.950 483.450 766.050 484.050 ;
        RECT 767.400 483.450 768.450 490.950 ;
        RECT 763.950 482.400 768.450 483.450 ;
        RECT 763.950 481.950 766.050 482.400 ;
        RECT 751.950 478.950 754.050 481.050 ;
        RECT 752.400 478.050 753.450 478.950 ;
        RECT 755.400 478.050 756.450 481.950 ;
        RECT 751.950 475.950 754.050 478.050 ;
        RECT 754.950 475.950 757.050 478.050 ;
        RECT 757.950 472.950 760.050 475.050 ;
        RECT 748.950 454.950 751.050 457.050 ;
        RECT 752.250 455.250 753.750 456.150 ;
        RECT 754.950 454.950 757.050 457.050 ;
        RECT 758.400 456.450 759.450 472.950 ;
        RECT 761.400 460.050 762.450 481.950 ;
        RECT 766.950 478.950 769.050 481.050 ;
        RECT 763.950 463.950 766.050 466.050 ;
        RECT 760.950 457.950 763.050 460.050 ;
        RECT 758.400 455.400 762.450 456.450 ;
        RECT 748.950 452.850 750.750 453.750 ;
        RECT 751.950 451.950 754.050 454.050 ;
        RECT 755.250 452.850 756.750 453.750 ;
        RECT 757.950 451.950 760.050 454.050 ;
        RECT 748.950 448.950 751.050 451.050 ;
        RECT 749.400 436.050 750.450 448.950 ;
        RECT 752.400 448.050 753.450 451.950 ;
        RECT 757.950 449.850 760.050 450.750 ;
        RECT 751.950 445.950 754.050 448.050 ;
        RECT 754.950 442.950 757.050 445.050 ;
        RECT 748.950 433.950 751.050 436.050 ;
        RECT 751.950 430.950 754.050 433.050 ;
        RECT 748.950 424.950 751.050 427.050 ;
        RECT 739.950 418.950 742.050 421.050 ;
        RECT 742.950 419.250 745.050 420.150 ;
        RECT 745.950 418.950 748.050 421.050 ;
        RECT 749.400 418.050 750.450 424.950 ;
        RECT 724.950 416.250 726.750 417.150 ;
        RECT 727.950 415.950 730.050 418.050 ;
        RECT 731.250 416.250 732.750 417.150 ;
        RECT 733.950 415.950 736.050 418.050 ;
        RECT 739.950 416.250 741.750 417.150 ;
        RECT 742.950 415.950 745.050 418.050 ;
        RECT 746.250 416.250 747.750 417.150 ;
        RECT 748.950 415.950 751.050 418.050 ;
        RECT 712.950 413.250 714.750 414.150 ;
        RECT 715.950 412.950 718.050 415.050 ;
        RECT 718.950 412.950 721.050 415.050 ;
        RECT 721.950 412.950 724.050 415.050 ;
        RECT 724.950 412.950 727.050 415.050 ;
        RECT 727.950 412.950 730.050 415.050 ;
        RECT 730.950 412.950 733.050 415.050 ;
        RECT 734.250 413.850 736.050 414.750 ;
        RECT 739.950 412.950 742.050 415.050 ;
        RECT 712.950 409.950 715.050 412.050 ;
        RECT 716.250 410.850 718.050 411.750 ;
        RECT 718.950 410.250 721.050 411.150 ;
        RECT 721.950 410.850 724.050 411.750 ;
        RECT 713.400 399.450 714.450 409.950 ;
        RECT 718.950 408.450 721.050 409.050 ;
        RECT 725.400 408.450 726.450 412.950 ;
        RECT 718.950 407.400 726.450 408.450 ;
        RECT 718.950 406.950 721.050 407.400 ;
        RECT 713.400 398.400 717.450 399.450 ;
        RECT 716.400 397.050 717.450 398.400 ;
        RECT 710.400 395.400 714.450 396.450 ;
        RECT 709.950 388.950 712.050 391.050 ;
        RECT 710.400 388.050 711.450 388.950 ;
        RECT 704.400 386.400 708.450 387.450 ;
        RECT 707.400 385.050 708.450 386.400 ;
        RECT 709.950 385.950 712.050 388.050 ;
        RECT 703.950 382.950 706.050 385.050 ;
        RECT 706.950 382.950 709.050 385.050 ;
        RECT 704.400 382.050 705.450 382.950 ;
        RECT 710.400 382.050 711.450 385.950 ;
        RECT 700.950 380.250 702.750 381.150 ;
        RECT 703.950 379.950 706.050 382.050 ;
        RECT 709.950 379.950 712.050 382.050 ;
        RECT 700.950 376.950 703.050 379.050 ;
        RECT 704.250 377.850 705.750 378.750 ;
        RECT 706.950 376.950 709.050 379.050 ;
        RECT 710.250 377.850 712.050 378.750 ;
        RECT 706.950 374.850 709.050 375.750 ;
        RECT 709.950 370.950 712.050 373.050 ;
        RECT 700.950 367.950 703.050 370.050 ;
        RECT 694.950 347.250 697.050 348.150 ;
        RECT 697.950 346.950 700.050 349.050 ;
        RECT 688.950 343.950 691.050 346.050 ;
        RECT 692.250 344.250 693.750 345.150 ;
        RECT 694.950 343.950 697.050 346.050 ;
        RECT 698.250 344.250 700.050 345.150 ;
        RECT 688.950 341.850 690.750 342.750 ;
        RECT 691.950 340.950 694.050 343.050 ;
        RECT 685.950 328.950 688.050 331.050 ;
        RECT 692.400 328.050 693.450 340.950 ;
        RECT 695.400 340.050 696.450 343.950 ;
        RECT 697.950 340.950 700.050 343.050 ;
        RECT 694.950 337.950 697.050 340.050 ;
        RECT 691.950 325.950 694.050 328.050 ;
        RECT 691.950 319.950 694.050 322.050 ;
        RECT 685.950 316.950 688.050 319.050 ;
        RECT 686.400 306.450 687.450 316.950 ;
        RECT 692.400 310.050 693.450 319.950 ;
        RECT 695.400 316.050 696.450 337.950 ;
        RECT 701.400 334.050 702.450 367.950 ;
        RECT 710.400 352.050 711.450 370.950 ;
        RECT 713.400 364.050 714.450 395.400 ;
        RECT 715.950 394.950 718.050 397.050 ;
        RECT 715.950 391.950 718.050 394.050 ;
        RECT 716.400 388.050 717.450 391.950 ;
        RECT 715.950 385.950 718.050 388.050 ;
        RECT 716.400 385.050 717.450 385.950 ;
        RECT 722.400 385.050 723.450 407.400 ;
        RECT 724.950 403.950 727.050 406.050 ;
        RECT 715.950 382.950 718.050 385.050 ;
        RECT 719.250 383.250 720.750 384.150 ;
        RECT 721.950 382.950 724.050 385.050 ;
        RECT 725.400 384.450 726.450 403.950 ;
        RECT 728.400 394.050 729.450 412.950 ;
        RECT 731.400 412.050 732.450 412.950 ;
        RECT 730.950 409.950 733.050 412.050 ;
        RECT 730.950 406.950 733.050 409.050 ;
        RECT 727.950 391.950 730.050 394.050 ;
        RECT 725.400 383.400 729.450 384.450 ;
        RECT 715.950 380.850 717.750 381.750 ;
        RECT 718.950 379.950 721.050 382.050 ;
        RECT 722.250 380.850 723.750 381.750 ;
        RECT 724.950 379.950 727.050 382.050 ;
        RECT 719.400 370.050 720.450 379.950 ;
        RECT 724.950 377.850 727.050 378.750 ;
        RECT 718.950 367.950 721.050 370.050 ;
        RECT 719.400 367.050 720.450 367.950 ;
        RECT 718.950 364.950 721.050 367.050 ;
        RECT 712.950 361.950 715.050 364.050 ;
        RECT 718.950 358.950 721.050 361.050 ;
        RECT 706.950 349.950 709.050 352.050 ;
        RECT 709.950 349.950 712.050 352.050 ;
        RECT 703.950 346.950 706.050 349.050 ;
        RECT 700.950 331.950 703.050 334.050 ;
        RECT 704.400 325.050 705.450 346.950 ;
        RECT 707.400 346.050 708.450 349.950 ;
        RECT 712.950 347.250 715.050 348.150 ;
        RECT 706.950 343.950 709.050 346.050 ;
        RECT 710.250 344.250 711.750 345.150 ;
        RECT 712.950 343.950 715.050 346.050 ;
        RECT 716.250 344.250 718.050 345.150 ;
        RECT 713.400 343.050 714.450 343.950 ;
        RECT 719.400 343.050 720.450 358.950 ;
        RECT 721.950 349.950 724.050 352.050 ;
        RECT 706.950 341.850 708.750 342.750 ;
        RECT 709.950 340.950 712.050 343.050 ;
        RECT 712.950 340.950 715.050 343.050 ;
        RECT 715.950 342.450 718.050 343.050 ;
        RECT 718.950 342.450 721.050 343.050 ;
        RECT 715.950 341.400 721.050 342.450 ;
        RECT 715.950 340.950 718.050 341.400 ;
        RECT 718.950 340.950 721.050 341.400 ;
        RECT 710.400 340.050 711.450 340.950 ;
        RECT 709.950 337.950 712.050 340.050 ;
        RECT 706.950 333.450 709.050 334.050 ;
        RECT 706.950 332.400 711.450 333.450 ;
        RECT 706.950 331.950 709.050 332.400 ;
        RECT 703.950 322.950 706.050 325.050 ;
        RECT 703.950 319.950 706.050 322.050 ;
        RECT 694.950 313.950 697.050 316.050 ;
        RECT 697.950 310.950 700.050 313.050 ;
        RECT 698.400 310.050 699.450 310.950 ;
        RECT 704.400 310.050 705.450 319.950 ;
        RECT 706.950 316.950 709.050 319.050 ;
        RECT 707.400 313.050 708.450 316.950 ;
        RECT 706.950 310.950 709.050 313.050 ;
        RECT 688.950 308.250 690.750 309.150 ;
        RECT 691.950 307.950 694.050 310.050 ;
        RECT 697.950 307.950 700.050 310.050 ;
        RECT 700.950 308.250 702.750 309.150 ;
        RECT 703.950 307.950 706.050 310.050 ;
        RECT 707.250 308.250 709.050 309.150 ;
        RECT 688.950 306.450 691.050 307.050 ;
        RECT 686.400 305.400 691.050 306.450 ;
        RECT 692.250 305.850 693.750 306.750 ;
        RECT 688.950 304.950 691.050 305.400 ;
        RECT 694.950 304.950 697.050 307.050 ;
        RECT 698.250 305.850 700.050 306.750 ;
        RECT 700.950 304.950 703.050 307.050 ;
        RECT 704.250 305.850 705.750 306.750 ;
        RECT 706.950 304.950 709.050 307.050 ;
        RECT 694.950 302.850 697.050 303.750 ;
        RECT 691.950 298.950 694.050 301.050 ;
        RECT 682.950 295.950 685.050 298.050 ;
        RECT 679.950 292.950 682.050 295.050 ;
        RECT 688.950 277.950 691.050 280.050 ;
        RECT 682.950 271.950 685.050 274.050 ;
        RECT 683.400 271.050 684.450 271.950 ;
        RECT 689.400 271.050 690.450 277.950 ;
        RECT 692.400 277.050 693.450 298.950 ;
        RECT 694.950 277.950 697.050 280.050 ;
        RECT 691.950 274.950 694.050 277.050 ;
        RECT 691.950 271.950 694.050 274.050 ;
        RECT 679.950 269.250 681.750 270.150 ;
        RECT 682.950 268.950 685.050 271.050 ;
        RECT 688.950 268.950 691.050 271.050 ;
        RECT 679.950 265.950 682.050 268.050 ;
        RECT 683.250 266.850 685.050 267.750 ;
        RECT 685.950 266.250 688.050 267.150 ;
        RECT 688.950 266.850 691.050 267.750 ;
        RECT 665.400 245.400 675.450 246.450 ;
        RECT 665.400 241.050 666.450 245.400 ;
        RECT 674.400 244.050 675.450 245.400 ;
        RECT 676.950 244.950 679.050 247.050 ;
        RECT 667.950 241.950 670.050 244.050 ;
        RECT 670.950 241.950 673.050 244.050 ;
        RECT 673.950 241.950 676.050 244.050 ;
        RECT 680.400 243.450 681.450 265.950 ;
        RECT 685.950 262.950 688.050 265.050 ;
        RECT 692.400 264.450 693.450 271.950 ;
        RECT 695.400 271.050 696.450 277.950 ;
        RECT 701.400 277.050 702.450 304.950 ;
        RECT 707.400 295.050 708.450 304.950 ;
        RECT 710.400 295.050 711.450 332.400 ;
        RECT 718.950 322.950 721.050 325.050 ;
        RECT 715.950 313.950 718.050 316.050 ;
        RECT 716.400 312.450 717.450 313.950 ;
        RECT 713.400 311.400 717.450 312.450 ;
        RECT 713.400 303.450 714.450 311.400 ;
        RECT 719.400 310.050 720.450 322.950 ;
        RECT 722.400 319.050 723.450 349.950 ;
        RECT 728.400 345.450 729.450 383.400 ;
        RECT 731.400 349.050 732.450 406.950 ;
        RECT 733.950 400.950 736.050 403.050 ;
        RECT 734.400 391.050 735.450 400.950 ;
        RECT 740.400 400.050 741.450 412.950 ;
        RECT 743.400 403.050 744.450 415.950 ;
        RECT 745.950 412.950 748.050 415.050 ;
        RECT 749.250 413.850 751.050 414.750 ;
        RECT 748.950 409.950 751.050 412.050 ;
        RECT 742.950 400.950 745.050 403.050 ;
        RECT 739.950 397.950 742.050 400.050 ;
        RECT 733.950 388.950 736.050 391.050 ;
        RECT 736.950 388.950 739.050 391.050 ;
        RECT 737.400 388.050 738.450 388.950 ;
        RECT 736.950 385.950 739.050 388.050 ;
        RECT 740.400 385.050 741.450 397.950 ;
        RECT 745.950 391.950 748.050 394.050 ;
        RECT 746.400 385.050 747.450 391.950 ;
        RECT 749.400 385.050 750.450 409.950 ;
        RECT 752.400 400.050 753.450 430.950 ;
        RECT 751.950 397.950 754.050 400.050 ;
        RECT 751.950 385.950 754.050 388.050 ;
        RECT 733.950 383.250 736.050 384.150 ;
        RECT 736.950 383.850 739.050 384.750 ;
        RECT 739.950 382.950 742.050 385.050 ;
        RECT 743.250 383.250 744.750 384.150 ;
        RECT 745.950 382.950 748.050 385.050 ;
        RECT 748.950 382.950 751.050 385.050 ;
        RECT 752.400 382.050 753.450 385.950 ;
        RECT 733.950 379.950 736.050 382.050 ;
        RECT 736.950 379.950 739.050 382.050 ;
        RECT 739.950 380.850 741.750 381.750 ;
        RECT 742.950 379.950 745.050 382.050 ;
        RECT 746.250 380.850 747.750 381.750 ;
        RECT 748.950 381.450 751.050 382.050 ;
        RECT 751.950 381.450 754.050 382.050 ;
        RECT 748.950 380.400 754.050 381.450 ;
        RECT 748.950 379.950 751.050 380.400 ;
        RECT 751.950 379.950 754.050 380.400 ;
        RECT 734.400 379.050 735.450 379.950 ;
        RECT 733.950 376.950 736.050 379.050 ;
        RECT 733.950 373.950 736.050 376.050 ;
        RECT 730.950 346.950 733.050 349.050 ;
        RECT 734.400 346.050 735.450 373.950 ;
        RECT 737.400 373.050 738.450 379.950 ;
        RECT 743.400 379.050 744.450 379.950 ;
        RECT 739.950 376.950 742.050 379.050 ;
        RECT 742.950 376.950 745.050 379.050 ;
        RECT 748.950 377.850 751.050 378.750 ;
        RECT 736.950 370.950 739.050 373.050 ;
        RECT 740.400 346.050 741.450 376.950 ;
        RECT 748.950 361.950 751.050 364.050 ;
        RECT 724.950 344.250 727.050 345.150 ;
        RECT 728.400 344.400 732.450 345.450 ;
        RECT 731.400 343.050 732.450 344.400 ;
        RECT 733.950 343.950 736.050 346.050 ;
        RECT 739.950 343.950 742.050 346.050 ;
        RECT 745.950 344.250 748.050 345.150 ;
        RECT 724.950 340.950 727.050 343.050 ;
        RECT 728.250 341.250 729.750 342.150 ;
        RECT 730.950 340.950 733.050 343.050 ;
        RECT 734.250 341.250 736.050 342.150 ;
        RECT 736.950 341.250 738.750 342.150 ;
        RECT 739.950 340.950 742.050 343.050 ;
        RECT 743.250 341.250 744.750 342.150 ;
        RECT 745.950 340.950 748.050 343.050 ;
        RECT 727.950 337.950 730.050 340.050 ;
        RECT 731.250 338.850 732.750 339.750 ;
        RECT 733.950 339.450 736.050 340.050 ;
        RECT 736.950 339.450 739.050 340.050 ;
        RECT 733.950 338.400 739.050 339.450 ;
        RECT 740.250 338.850 741.750 339.750 ;
        RECT 733.950 337.950 736.050 338.400 ;
        RECT 736.950 337.950 739.050 338.400 ;
        RECT 742.950 337.950 745.050 340.050 ;
        RECT 728.400 334.050 729.450 337.950 ;
        RECT 727.950 331.950 730.050 334.050 ;
        RECT 721.950 316.950 724.050 319.050 ;
        RECT 724.950 313.950 727.050 316.050 ;
        RECT 730.950 313.950 733.050 316.050 ;
        RECT 725.400 310.050 726.450 313.950 ;
        RECT 737.400 313.050 738.450 337.950 ;
        RECT 743.400 337.050 744.450 337.950 ;
        RECT 742.950 334.950 745.050 337.050 ;
        RECT 742.950 328.950 745.050 331.050 ;
        RECT 739.950 313.950 742.050 316.050 ;
        RECT 727.950 311.250 730.050 312.150 ;
        RECT 730.950 311.850 733.050 312.750 ;
        RECT 733.950 311.250 735.750 312.150 ;
        RECT 736.950 310.950 739.050 313.050 ;
        RECT 740.400 310.050 741.450 313.950 ;
        RECT 715.950 308.250 717.750 309.150 ;
        RECT 718.950 307.950 721.050 310.050 ;
        RECT 721.950 307.950 724.050 310.050 ;
        RECT 724.950 307.950 727.050 310.050 ;
        RECT 727.950 307.950 730.050 310.050 ;
        RECT 733.950 307.950 736.050 310.050 ;
        RECT 737.250 308.850 739.050 309.750 ;
        RECT 739.950 307.950 742.050 310.050 ;
        RECT 722.400 307.050 723.450 307.950 ;
        RECT 715.950 304.950 718.050 307.050 ;
        RECT 719.250 305.850 720.750 306.750 ;
        RECT 721.950 304.950 724.050 307.050 ;
        RECT 725.250 305.850 727.050 306.750 ;
        RECT 713.400 302.400 717.450 303.450 ;
        RECT 721.950 302.850 724.050 303.750 ;
        RECT 712.950 295.950 715.050 298.050 ;
        RECT 706.950 292.950 709.050 295.050 ;
        RECT 709.950 292.950 712.050 295.050 ;
        RECT 700.950 274.950 703.050 277.050 ;
        RECT 707.400 274.050 708.450 292.950 ;
        RECT 706.950 271.950 709.050 274.050 ;
        RECT 709.950 272.250 712.050 273.150 ;
        RECT 694.950 268.950 697.050 271.050 ;
        RECT 700.950 269.250 702.750 270.150 ;
        RECT 703.950 268.950 706.050 271.050 ;
        RECT 707.250 269.250 708.750 270.150 ;
        RECT 709.950 268.950 712.050 271.050 ;
        RECT 694.950 266.850 697.050 267.750 ;
        RECT 697.950 266.250 700.050 267.150 ;
        RECT 700.950 265.950 703.050 268.050 ;
        RECT 704.250 266.850 705.750 267.750 ;
        RECT 706.950 265.950 709.050 268.050 ;
        RECT 697.950 264.450 700.050 265.050 ;
        RECT 701.400 264.450 702.450 265.950 ;
        RECT 692.400 263.400 696.450 264.450 ;
        RECT 685.950 259.950 688.050 262.050 ;
        RECT 688.950 261.450 691.050 262.050 ;
        RECT 691.950 261.450 694.050 262.050 ;
        RECT 688.950 260.400 694.050 261.450 ;
        RECT 688.950 259.950 691.050 260.400 ;
        RECT 691.950 259.950 694.050 260.400 ;
        RECT 682.950 243.450 685.050 244.050 ;
        RECT 680.400 242.400 685.050 243.450 ;
        RECT 682.950 241.950 685.050 242.400 ;
        RECT 661.950 238.950 664.050 241.050 ;
        RECT 664.950 238.950 667.050 241.050 ;
        RECT 661.950 236.250 664.050 237.150 ;
        RECT 664.950 236.850 667.050 237.750 ;
        RECT 656.400 233.400 660.450 234.450 ;
        RECT 653.400 229.050 654.450 232.950 ;
        RECT 652.950 226.950 655.050 229.050 ;
        RECT 646.950 217.950 649.050 220.050 ;
        RECT 643.950 205.950 646.050 208.050 ;
        RECT 647.400 205.050 648.450 217.950 ;
        RECT 641.400 203.400 645.450 204.450 ;
        RECT 634.950 199.950 637.050 202.050 ;
        RECT 638.250 200.250 639.750 201.150 ;
        RECT 640.950 199.950 643.050 202.050 ;
        RECT 634.950 197.850 636.750 198.750 ;
        RECT 637.950 196.950 640.050 199.050 ;
        RECT 641.250 197.850 643.050 198.750 ;
        RECT 644.400 198.450 645.450 203.400 ;
        RECT 646.950 202.950 649.050 205.050 ;
        RECT 649.950 203.250 652.050 204.150 ;
        RECT 656.400 202.050 657.450 233.400 ;
        RECT 661.950 232.950 664.050 235.050 ;
        RECT 664.950 232.950 667.050 235.050 ;
        RECT 662.400 229.050 663.450 232.950 ;
        RECT 661.950 226.950 664.050 229.050 ;
        RECT 665.400 226.050 666.450 232.950 ;
        RECT 664.950 223.950 667.050 226.050 ;
        RECT 661.950 220.950 664.050 223.050 ;
        RECT 658.950 217.950 661.050 220.050 ;
        RECT 646.950 200.250 648.750 201.150 ;
        RECT 649.950 199.950 652.050 202.050 ;
        RECT 653.250 200.250 654.750 201.150 ;
        RECT 655.950 199.950 658.050 202.050 ;
        RECT 646.950 198.450 649.050 199.050 ;
        RECT 644.400 197.400 649.050 198.450 ;
        RECT 646.950 196.950 649.050 197.400 ;
        RECT 649.950 196.950 652.050 199.050 ;
        RECT 652.950 196.950 655.050 199.050 ;
        RECT 656.250 197.850 658.050 198.750 ;
        RECT 632.400 194.400 636.450 195.450 ;
        RECT 625.950 190.950 628.050 193.050 ;
        RECT 628.950 190.950 631.050 193.050 ;
        RECT 631.950 190.950 634.050 193.050 ;
        RECT 625.950 187.950 628.050 190.050 ;
        RECT 626.400 160.050 627.450 187.950 ;
        RECT 629.400 172.050 630.450 190.950 ;
        RECT 632.400 172.050 633.450 190.950 ;
        RECT 628.950 169.950 631.050 172.050 ;
        RECT 631.950 169.950 634.050 172.050 ;
        RECT 628.950 167.250 631.050 168.150 ;
        RECT 631.950 167.850 634.050 168.750 ;
        RECT 628.950 163.950 631.050 166.050 ;
        RECT 625.950 157.950 628.050 160.050 ;
        RECT 629.400 145.050 630.450 163.950 ;
        RECT 635.400 151.050 636.450 194.400 ;
        RECT 638.400 193.050 639.450 196.950 ;
        RECT 646.950 193.950 649.050 196.050 ;
        RECT 637.950 190.950 640.050 193.050 ;
        RECT 643.950 190.950 646.050 193.050 ;
        RECT 644.400 187.050 645.450 190.950 ;
        RECT 647.400 187.050 648.450 193.950 ;
        RECT 643.950 184.950 646.050 187.050 ;
        RECT 646.950 184.950 649.050 187.050 ;
        RECT 650.400 181.050 651.450 196.950 ;
        RECT 653.400 190.050 654.450 196.950 ;
        RECT 655.950 193.950 658.050 196.050 ;
        RECT 652.950 187.950 655.050 190.050 ;
        RECT 652.950 184.950 655.050 187.050 ;
        RECT 637.950 178.950 640.050 181.050 ;
        RECT 649.950 178.950 652.050 181.050 ;
        RECT 634.950 148.950 637.050 151.050 ;
        RECT 634.950 145.950 637.050 148.050 ;
        RECT 628.950 142.950 631.050 145.050 ;
        RECT 616.950 130.950 619.050 133.050 ;
        RECT 619.950 131.250 622.050 132.150 ;
        RECT 622.950 130.950 625.050 133.050 ;
        RECT 616.950 128.250 618.750 129.150 ;
        RECT 619.950 127.950 622.050 130.050 ;
        RECT 625.950 129.450 628.050 130.050 ;
        RECT 631.950 129.450 634.050 130.050 ;
        RECT 635.400 129.450 636.450 145.950 ;
        RECT 638.400 130.050 639.450 178.950 ;
        RECT 643.950 175.950 646.050 178.050 ;
        RECT 644.400 169.050 645.450 175.950 ;
        RECT 643.950 166.950 646.050 169.050 ;
        RECT 647.250 167.250 648.750 168.150 ;
        RECT 649.950 166.950 652.050 169.050 ;
        RECT 640.950 163.950 643.050 166.050 ;
        RECT 644.250 164.850 645.750 165.750 ;
        RECT 646.950 163.950 649.050 166.050 ;
        RECT 650.250 164.850 652.050 165.750 ;
        RECT 640.950 161.850 643.050 162.750 ;
        RECT 647.400 160.050 648.450 163.950 ;
        RECT 649.950 160.950 652.050 163.050 ;
        RECT 646.950 157.950 649.050 160.050 ;
        RECT 646.950 136.950 649.050 139.050 ;
        RECT 643.950 130.950 646.050 133.050 ;
        RECT 623.250 128.250 624.750 129.150 ;
        RECT 625.950 128.400 630.450 129.450 ;
        RECT 625.950 127.950 628.050 128.400 ;
        RECT 616.950 124.950 619.050 127.050 ;
        RECT 620.400 118.050 621.450 127.950 ;
        RECT 622.950 124.950 625.050 127.050 ;
        RECT 626.250 125.850 628.050 126.750 ;
        RECT 619.950 115.950 622.050 118.050 ;
        RECT 623.400 115.050 624.450 124.950 ;
        RECT 625.950 121.950 628.050 124.050 ;
        RECT 622.950 112.950 625.050 115.050 ;
        RECT 626.400 100.050 627.450 121.950 ;
        RECT 629.400 112.050 630.450 128.400 ;
        RECT 631.950 128.400 636.450 129.450 ;
        RECT 631.950 127.950 634.050 128.400 ;
        RECT 631.950 124.950 634.050 127.050 ;
        RECT 635.400 126.450 636.450 128.400 ;
        RECT 637.950 127.950 640.050 130.050 ;
        RECT 637.950 126.450 640.050 127.050 ;
        RECT 635.400 125.400 640.050 126.450 ;
        RECT 637.950 124.950 640.050 125.400 ;
        RECT 641.250 125.250 643.050 126.150 ;
        RECT 631.950 122.850 634.050 123.750 ;
        RECT 634.950 122.250 637.050 123.150 ;
        RECT 637.950 122.850 639.750 123.750 ;
        RECT 640.950 121.950 643.050 124.050 ;
        RECT 634.950 118.950 637.050 121.050 ;
        RECT 635.400 118.050 636.450 118.950 ;
        RECT 634.950 115.950 637.050 118.050 ;
        RECT 628.950 109.950 631.050 112.050 ;
        RECT 637.950 103.950 640.050 106.050 ;
        RECT 628.950 100.950 631.050 103.050 ;
        RECT 614.400 98.400 618.450 99.450 ;
        RECT 613.950 94.950 616.050 97.050 ;
        RECT 604.950 92.250 606.750 93.150 ;
        RECT 607.950 91.950 610.050 94.050 ;
        RECT 611.250 92.250 613.050 93.150 ;
        RECT 613.950 92.850 616.050 93.750 ;
        RECT 604.950 88.950 607.050 91.050 ;
        RECT 608.250 89.850 609.750 90.750 ;
        RECT 610.950 88.950 613.050 91.050 ;
        RECT 611.400 88.050 612.450 88.950 ;
        RECT 610.950 85.950 613.050 88.050 ;
        RECT 604.950 64.950 607.050 67.050 ;
        RECT 592.950 43.950 595.050 46.050 ;
        RECT 598.950 43.950 601.050 46.050 ;
        RECT 601.950 43.950 604.050 46.050 ;
        RECT 592.950 37.950 595.050 40.050 ;
        RECT 583.950 26.400 588.450 27.450 ;
        RECT 583.950 25.950 586.050 26.400 ;
        RECT 587.400 25.050 588.450 26.400 ;
        RECT 550.950 23.250 553.050 24.150 ;
        RECT 560.400 23.400 564.450 24.450 ;
        RECT 511.950 20.850 514.050 21.750 ;
        RECT 517.950 19.950 520.050 22.050 ;
        RECT 520.950 20.850 523.050 21.750 ;
        RECT 526.950 20.850 529.050 21.750 ;
        RECT 529.950 20.850 531.750 21.750 ;
        RECT 532.950 19.950 535.050 22.050 ;
        RECT 536.250 20.850 537.750 21.750 ;
        RECT 538.950 19.950 541.050 22.050 ;
        RECT 550.950 19.950 553.050 22.050 ;
        RECT 556.950 19.950 559.050 22.050 ;
        RECT 560.400 19.050 561.450 23.400 ;
        RECT 574.950 23.250 577.050 24.150 ;
        RECT 580.950 22.950 583.050 25.050 ;
        RECT 584.250 23.850 586.050 24.750 ;
        RECT 586.950 22.950 589.050 25.050 ;
        RECT 593.400 22.050 594.450 37.950 ;
        RECT 562.950 19.950 565.050 22.050 ;
        RECT 566.250 20.250 568.050 21.150 ;
        RECT 574.950 19.950 577.050 22.050 ;
        RECT 580.950 20.850 583.050 21.750 ;
        RECT 589.950 20.250 591.750 21.150 ;
        RECT 592.950 19.950 595.050 22.050 ;
        RECT 596.250 20.250 598.050 21.150 ;
        RECT 505.950 17.400 510.450 18.450 ;
        RECT 538.950 17.850 541.050 18.750 ;
        RECT 556.950 17.850 558.750 18.750 ;
        RECT 505.950 16.950 508.050 17.400 ;
        RECT 559.950 16.950 562.050 19.050 ;
        RECT 563.250 17.850 564.750 18.750 ;
        RECT 565.950 16.950 568.050 19.050 ;
        RECT 589.950 16.950 592.050 19.050 ;
        RECT 593.250 17.850 594.750 18.750 ;
        RECT 595.950 16.950 598.050 19.050 ;
        RECT 599.400 18.450 600.450 43.950 ;
        RECT 605.400 40.050 606.450 64.950 ;
        RECT 607.950 53.250 610.050 54.150 ;
        RECT 613.950 53.250 616.050 54.150 ;
        RECT 617.400 52.050 618.450 98.400 ;
        RECT 625.950 97.950 628.050 100.050 ;
        RECT 629.400 97.050 630.450 100.950 ;
        RECT 638.400 100.050 639.450 103.950 ;
        RECT 641.400 100.050 642.450 121.950 ;
        RECT 631.950 97.950 634.050 100.050 ;
        RECT 637.950 97.950 640.050 100.050 ;
        RECT 640.950 97.950 643.050 100.050 ;
        RECT 632.400 97.050 633.450 97.950 ;
        RECT 622.950 96.450 625.050 97.050 ;
        RECT 622.950 95.400 627.450 96.450 ;
        RECT 622.950 94.950 625.050 95.400 ;
        RECT 619.950 92.250 622.050 93.150 ;
        RECT 622.950 92.850 625.050 93.750 ;
        RECT 626.400 91.050 627.450 95.400 ;
        RECT 628.950 94.950 631.050 97.050 ;
        RECT 631.950 94.950 634.050 97.050 ;
        RECT 635.250 95.250 637.050 96.150 ;
        RECT 637.950 95.850 640.050 96.750 ;
        RECT 640.950 95.250 643.050 96.150 ;
        RECT 628.950 91.950 631.050 94.050 ;
        RECT 631.950 92.850 633.750 93.750 ;
        RECT 634.950 91.950 637.050 94.050 ;
        RECT 637.950 91.950 640.050 94.050 ;
        RECT 640.950 91.950 643.050 94.050 ;
        RECT 619.950 88.950 622.050 91.050 ;
        RECT 625.950 88.950 628.050 91.050 ;
        RECT 620.400 88.050 621.450 88.950 ;
        RECT 629.400 88.050 630.450 91.950 ;
        RECT 619.950 85.950 622.050 88.050 ;
        RECT 628.950 85.950 631.050 88.050 ;
        RECT 638.400 73.050 639.450 91.950 ;
        RECT 641.400 91.050 642.450 91.950 ;
        RECT 640.950 88.950 643.050 91.050 ;
        RECT 637.950 70.950 640.050 73.050 ;
        RECT 640.950 58.950 643.050 61.050 ;
        RECT 641.400 58.050 642.450 58.950 ;
        RECT 619.950 56.250 622.050 57.150 ;
        RECT 625.950 55.950 628.050 58.050 ;
        RECT 634.950 57.450 637.050 58.050 ;
        RECT 632.400 56.400 637.050 57.450 ;
        RECT 626.400 55.050 627.450 55.950 ;
        RECT 619.950 52.950 622.050 55.050 ;
        RECT 623.250 53.250 624.750 54.150 ;
        RECT 625.950 52.950 628.050 55.050 ;
        RECT 629.250 53.250 631.050 54.150 ;
        RECT 607.950 49.950 610.050 52.050 ;
        RECT 613.950 51.450 616.050 52.050 ;
        RECT 616.950 51.450 619.050 52.050 ;
        RECT 611.250 50.250 612.750 51.150 ;
        RECT 613.950 50.400 619.050 51.450 ;
        RECT 613.950 49.950 616.050 50.400 ;
        RECT 616.950 49.950 619.050 50.400 ;
        RECT 614.400 49.050 615.450 49.950 ;
        RECT 610.950 46.950 613.050 49.050 ;
        RECT 613.950 46.950 616.050 49.050 ;
        RECT 611.400 40.050 612.450 46.950 ;
        RECT 620.400 46.050 621.450 52.950 ;
        RECT 622.950 49.950 625.050 52.050 ;
        RECT 626.250 50.850 627.750 51.750 ;
        RECT 628.950 49.950 631.050 52.050 ;
        RECT 619.950 43.950 622.050 46.050 ;
        RECT 604.950 37.950 607.050 40.050 ;
        RECT 610.950 37.950 613.050 40.050 ;
        RECT 601.950 20.250 603.750 21.150 ;
        RECT 604.950 19.950 607.050 22.050 ;
        RECT 608.250 20.250 610.050 21.150 ;
        RECT 601.950 18.450 604.050 19.050 ;
        RECT 599.400 17.400 604.050 18.450 ;
        RECT 605.250 17.850 606.750 18.750 ;
        RECT 607.950 18.450 610.050 19.050 ;
        RECT 611.400 18.450 612.450 37.950 ;
        RECT 616.950 25.950 619.050 28.050 ;
        RECT 617.400 25.050 618.450 25.950 ;
        RECT 616.950 22.950 619.050 25.050 ;
        RECT 623.400 24.450 624.450 49.950 ;
        RECT 632.400 40.050 633.450 56.400 ;
        RECT 634.950 55.950 637.050 56.400 ;
        RECT 638.250 56.250 639.750 57.150 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 634.950 53.850 636.750 54.750 ;
        RECT 637.950 52.950 640.050 55.050 ;
        RECT 641.250 53.850 643.050 54.750 ;
        RECT 631.950 37.950 634.050 40.050 ;
        RECT 638.400 28.050 639.450 52.950 ;
        RECT 631.950 25.950 634.050 28.050 ;
        RECT 637.950 25.950 640.050 28.050 ;
        RECT 620.400 23.400 624.450 24.450 ;
        RECT 617.400 22.050 618.450 22.950 ;
        RECT 613.950 20.250 615.750 21.150 ;
        RECT 616.950 19.950 619.050 22.050 ;
        RECT 620.400 19.050 621.450 23.400 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 626.400 22.050 627.450 22.950 ;
        RECT 632.400 22.050 633.450 25.950 ;
        RECT 644.400 25.050 645.450 130.950 ;
        RECT 647.400 118.050 648.450 136.950 ;
        RECT 650.400 130.050 651.450 160.950 ;
        RECT 653.400 148.050 654.450 184.950 ;
        RECT 656.400 184.050 657.450 193.950 ;
        RECT 655.950 181.950 658.050 184.050 ;
        RECT 659.400 178.050 660.450 217.950 ;
        RECT 658.950 175.950 661.050 178.050 ;
        RECT 662.400 174.450 663.450 220.950 ;
        RECT 664.950 202.950 667.050 205.050 ;
        RECT 665.400 199.050 666.450 202.950 ;
        RECT 668.400 199.050 669.450 241.950 ;
        RECT 671.400 241.050 672.450 241.950 ;
        RECT 670.950 238.950 673.050 241.050 ;
        RECT 674.250 239.250 675.750 240.150 ;
        RECT 676.950 238.950 679.050 241.050 ;
        RECT 680.250 239.250 681.750 240.150 ;
        RECT 682.950 238.950 685.050 241.050 ;
        RECT 670.950 236.850 672.750 237.750 ;
        RECT 673.950 235.950 676.050 238.050 ;
        RECT 677.250 236.850 678.750 237.750 ;
        RECT 679.950 235.950 682.050 238.050 ;
        RECT 683.250 236.850 685.050 237.750 ;
        RECT 676.950 226.950 679.050 229.050 ;
        RECT 673.950 214.950 676.050 217.050 ;
        RECT 670.950 208.950 673.050 211.050 ;
        RECT 671.400 199.050 672.450 208.950 ;
        RECT 674.400 202.050 675.450 214.950 ;
        RECT 673.950 199.950 676.050 202.050 ;
        RECT 664.950 196.950 667.050 199.050 ;
        RECT 667.950 196.950 670.050 199.050 ;
        RECT 670.950 196.950 673.050 199.050 ;
        RECT 674.250 197.250 676.050 198.150 ;
        RECT 677.400 196.050 678.450 226.950 ;
        RECT 680.400 223.050 681.450 235.950 ;
        RECT 682.950 232.950 685.050 235.050 ;
        RECT 683.400 229.050 684.450 232.950 ;
        RECT 682.950 226.950 685.050 229.050 ;
        RECT 686.400 226.050 687.450 259.950 ;
        RECT 688.950 247.950 691.050 250.050 ;
        RECT 691.950 247.950 694.050 250.050 ;
        RECT 685.950 223.950 688.050 226.050 ;
        RECT 679.950 220.950 682.050 223.050 ;
        RECT 689.400 220.050 690.450 247.950 ;
        RECT 692.400 244.050 693.450 247.950 ;
        RECT 695.400 244.050 696.450 263.400 ;
        RECT 697.950 263.400 702.450 264.450 ;
        RECT 697.950 262.950 700.050 263.400 ;
        RECT 698.400 256.050 699.450 262.950 ;
        RECT 700.950 259.950 703.050 262.050 ;
        RECT 697.950 253.950 700.050 256.050 ;
        RECT 701.400 247.050 702.450 259.950 ;
        RECT 707.400 253.050 708.450 265.950 ;
        RECT 710.400 265.050 711.450 268.950 ;
        RECT 709.950 262.950 712.050 265.050 ;
        RECT 709.950 256.950 712.050 259.050 ;
        RECT 710.400 253.050 711.450 256.950 ;
        RECT 706.950 250.950 709.050 253.050 ;
        RECT 709.950 250.950 712.050 253.050 ;
        RECT 700.950 244.950 703.050 247.050 ;
        RECT 691.950 241.950 694.050 244.050 ;
        RECT 694.950 241.950 697.050 244.050 ;
        RECT 692.400 238.050 693.450 241.950 ;
        RECT 701.400 241.050 702.450 244.950 ;
        RECT 709.950 241.950 712.050 244.050 ;
        RECT 710.400 241.050 711.450 241.950 ;
        RECT 713.400 241.050 714.450 295.950 ;
        RECT 716.400 277.050 717.450 302.400 ;
        RECT 724.950 295.950 727.050 298.050 ;
        RECT 715.950 274.950 718.050 277.050 ;
        RECT 725.400 276.450 726.450 295.950 ;
        RECT 728.400 289.050 729.450 307.950 ;
        RECT 734.400 307.050 735.450 307.950 ;
        RECT 733.950 304.950 736.050 307.050 ;
        RECT 743.400 304.050 744.450 328.950 ;
        RECT 746.400 328.050 747.450 340.950 ;
        RECT 749.400 339.450 750.450 361.950 ;
        RECT 755.400 361.050 756.450 442.950 ;
        RECT 761.400 442.050 762.450 455.400 ;
        RECT 760.950 439.950 763.050 442.050 ;
        RECT 757.950 436.950 760.050 439.050 ;
        RECT 758.400 394.050 759.450 436.950 ;
        RECT 760.950 421.950 763.050 424.050 ;
        RECT 761.400 415.050 762.450 421.950 ;
        RECT 760.950 412.950 763.050 415.050 ;
        RECT 757.950 391.950 760.050 394.050 ;
        RECT 757.950 382.950 760.050 385.050 ;
        RECT 758.400 367.050 759.450 382.950 ;
        RECT 761.400 382.050 762.450 412.950 ;
        RECT 760.950 379.950 763.050 382.050 ;
        RECT 760.950 376.950 763.050 379.050 ;
        RECT 757.950 364.950 760.050 367.050 ;
        RECT 754.950 358.950 757.050 361.050 ;
        RECT 761.400 352.050 762.450 376.950 ;
        RECT 764.400 370.050 765.450 463.950 ;
        RECT 767.400 457.050 768.450 478.950 ;
        RECT 766.950 454.950 769.050 457.050 ;
        RECT 766.950 451.950 769.050 454.050 ;
        RECT 767.400 424.050 768.450 451.950 ;
        RECT 766.950 421.950 769.050 424.050 ;
        RECT 766.950 418.950 769.050 421.050 ;
        RECT 767.400 409.050 768.450 418.950 ;
        RECT 766.950 406.950 769.050 409.050 ;
        RECT 770.400 397.050 771.450 496.950 ;
        RECT 769.950 394.950 772.050 397.050 ;
        RECT 769.950 391.950 772.050 394.050 ;
        RECT 763.950 367.950 766.050 370.050 ;
        RECT 763.950 364.950 766.050 367.050 ;
        RECT 760.950 349.950 763.050 352.050 ;
        RECT 754.950 347.250 757.050 348.150 ;
        RECT 760.950 346.950 763.050 349.050 ;
        RECT 761.400 346.050 762.450 346.950 ;
        RECT 751.950 344.250 753.750 345.150 ;
        RECT 754.950 343.950 757.050 346.050 ;
        RECT 758.250 344.250 759.750 345.150 ;
        RECT 760.950 343.950 763.050 346.050 ;
        RECT 751.950 340.950 754.050 343.050 ;
        RECT 749.400 338.400 753.450 339.450 ;
        RECT 752.400 337.050 753.450 338.400 ;
        RECT 748.950 334.950 751.050 337.050 ;
        RECT 751.950 334.950 754.050 337.050 ;
        RECT 749.400 330.450 750.450 334.950 ;
        RECT 755.400 334.050 756.450 343.950 ;
        RECT 757.950 340.950 760.050 343.050 ;
        RECT 761.250 341.850 763.050 342.750 ;
        RECT 760.950 337.950 763.050 340.050 ;
        RECT 757.950 334.950 760.050 337.050 ;
        RECT 754.950 331.950 757.050 334.050 ;
        RECT 749.400 329.400 753.450 330.450 ;
        RECT 745.950 325.950 748.050 328.050 ;
        RECT 748.950 325.950 751.050 328.050 ;
        RECT 749.400 316.050 750.450 325.950 ;
        RECT 752.400 316.050 753.450 329.400 ;
        RECT 748.950 313.950 751.050 316.050 ;
        RECT 751.950 313.950 754.050 316.050 ;
        RECT 745.950 311.250 748.050 312.150 ;
        RECT 748.950 311.850 751.050 312.750 ;
        RECT 751.950 311.250 753.750 312.150 ;
        RECT 754.950 310.950 757.050 313.050 ;
        RECT 745.950 307.950 748.050 310.050 ;
        RECT 748.950 307.950 751.050 310.050 ;
        RECT 751.950 307.950 754.050 310.050 ;
        RECT 755.250 308.850 757.050 309.750 ;
        RECT 730.950 301.950 733.050 304.050 ;
        RECT 742.950 301.950 745.050 304.050 ;
        RECT 745.950 301.950 748.050 304.050 ;
        RECT 727.950 286.950 730.050 289.050 ;
        RECT 727.950 283.950 730.050 286.050 ;
        RECT 728.400 280.050 729.450 283.950 ;
        RECT 727.950 277.950 730.050 280.050 ;
        RECT 725.400 275.400 729.450 276.450 ;
        RECT 724.950 272.250 727.050 273.150 ;
        RECT 715.950 269.250 717.750 270.150 ;
        RECT 718.950 268.950 721.050 271.050 ;
        RECT 722.250 269.250 723.750 270.150 ;
        RECT 724.950 268.950 727.050 271.050 ;
        RECT 725.400 268.050 726.450 268.950 ;
        RECT 715.950 265.950 718.050 268.050 ;
        RECT 719.250 266.850 720.750 267.750 ;
        RECT 721.950 265.950 724.050 268.050 ;
        RECT 724.950 265.950 727.050 268.050 ;
        RECT 718.950 253.950 721.050 256.050 ;
        RECT 719.400 250.050 720.450 253.950 ;
        RECT 722.400 250.050 723.450 265.950 ;
        RECT 724.950 253.950 727.050 256.050 ;
        RECT 718.950 247.950 721.050 250.050 ;
        RECT 721.950 247.950 724.050 250.050 ;
        RECT 718.950 244.950 721.050 247.050 ;
        RECT 694.950 238.950 697.050 241.050 ;
        RECT 700.950 240.450 703.050 241.050 ;
        RECT 703.950 240.450 706.050 241.050 ;
        RECT 698.250 239.250 699.750 240.150 ;
        RECT 700.950 239.400 706.050 240.450 ;
        RECT 700.950 238.950 703.050 239.400 ;
        RECT 703.950 238.950 706.050 239.400 ;
        RECT 707.250 239.250 708.750 240.150 ;
        RECT 709.950 238.950 712.050 241.050 ;
        RECT 712.950 238.950 715.050 241.050 ;
        RECT 719.400 238.050 720.450 244.950 ;
        RECT 721.950 241.950 724.050 244.050 ;
        RECT 722.400 241.050 723.450 241.950 ;
        RECT 721.950 238.950 724.050 241.050 ;
        RECT 725.400 238.050 726.450 253.950 ;
        RECT 728.400 244.050 729.450 275.400 ;
        RECT 731.400 262.050 732.450 301.950 ;
        RECT 746.400 292.050 747.450 301.950 ;
        RECT 745.950 289.950 748.050 292.050 ;
        RECT 736.950 280.950 739.050 283.050 ;
        RECT 737.400 277.050 738.450 280.950 ;
        RECT 749.400 280.050 750.450 307.950 ;
        RECT 752.400 307.050 753.450 307.950 ;
        RECT 751.950 304.950 754.050 307.050 ;
        RECT 754.950 304.950 757.050 307.050 ;
        RECT 748.950 277.950 751.050 280.050 ;
        RECT 733.950 274.950 736.050 277.050 ;
        RECT 736.950 274.950 739.050 277.050 ;
        RECT 739.950 275.250 742.050 276.150 ;
        RECT 748.950 275.250 751.050 276.150 ;
        RECT 734.400 274.050 735.450 274.950 ;
        RECT 755.400 274.050 756.450 304.950 ;
        RECT 758.400 298.050 759.450 334.950 ;
        RECT 761.400 307.050 762.450 337.950 ;
        RECT 764.400 334.050 765.450 364.950 ;
        RECT 763.950 331.950 766.050 334.050 ;
        RECT 760.950 304.950 763.050 307.050 ;
        RECT 757.950 295.950 760.050 298.050 ;
        RECT 760.950 292.950 763.050 295.050 ;
        RECT 733.950 271.950 736.050 274.050 ;
        RECT 737.250 272.250 738.750 273.150 ;
        RECT 739.950 271.950 742.050 274.050 ;
        RECT 743.250 272.250 745.050 273.150 ;
        RECT 745.950 272.250 747.750 273.150 ;
        RECT 748.950 271.950 751.050 274.050 ;
        RECT 752.250 272.250 753.750 273.150 ;
        RECT 754.950 271.950 757.050 274.050 ;
        RECT 733.950 269.850 735.750 270.750 ;
        RECT 736.950 268.950 739.050 271.050 ;
        RECT 730.950 259.950 733.050 262.050 ;
        RECT 733.950 259.950 736.050 262.050 ;
        RECT 730.950 253.950 733.050 256.050 ;
        RECT 727.950 241.950 730.050 244.050 ;
        RECT 691.950 235.950 694.050 238.050 ;
        RECT 695.250 236.850 696.750 237.750 ;
        RECT 697.950 235.950 700.050 238.050 ;
        RECT 701.250 236.850 703.050 237.750 ;
        RECT 703.950 236.850 705.750 237.750 ;
        RECT 706.950 235.950 709.050 238.050 ;
        RECT 710.250 236.850 711.750 237.750 ;
        RECT 712.950 235.950 715.050 238.050 ;
        RECT 718.950 235.950 721.050 238.050 ;
        RECT 724.950 235.950 727.050 238.050 ;
        RECT 728.250 236.250 730.050 237.150 ;
        RECT 691.950 233.850 694.050 234.750 ;
        RECT 698.400 232.050 699.450 235.950 ;
        RECT 703.950 232.950 706.050 235.050 ;
        RECT 697.950 229.950 700.050 232.050 ;
        RECT 691.950 226.950 694.050 229.050 ;
        RECT 700.950 226.950 703.050 229.050 ;
        RECT 688.950 217.950 691.050 220.050 ;
        RECT 692.400 211.050 693.450 226.950 ;
        RECT 701.400 217.050 702.450 226.950 ;
        RECT 700.950 214.950 703.050 217.050 ;
        RECT 697.950 211.950 700.050 214.050 ;
        RECT 691.950 208.950 694.050 211.050 ;
        RECT 691.950 205.950 694.050 208.050 ;
        RECT 694.950 205.950 697.050 208.050 ;
        RECT 682.950 203.250 685.050 204.150 ;
        RECT 679.950 200.250 681.750 201.150 ;
        RECT 682.950 199.950 685.050 202.050 ;
        RECT 686.250 200.250 687.750 201.150 ;
        RECT 688.950 199.950 691.050 202.050 ;
        RECT 679.950 196.950 682.050 199.050 ;
        RECT 682.950 196.950 685.050 199.050 ;
        RECT 685.950 196.950 688.050 199.050 ;
        RECT 689.250 197.850 691.050 198.750 ;
        RECT 664.950 194.850 667.050 195.750 ;
        RECT 667.950 194.250 670.050 195.150 ;
        RECT 670.950 194.850 672.750 195.750 ;
        RECT 673.950 193.950 676.050 196.050 ;
        RECT 676.950 193.950 679.050 196.050 ;
        RECT 664.950 190.950 667.050 193.050 ;
        RECT 667.950 190.950 670.050 193.050 ;
        RECT 665.400 187.050 666.450 190.950 ;
        RECT 664.950 184.950 667.050 187.050 ;
        RECT 668.400 184.050 669.450 190.950 ;
        RECT 670.950 187.950 673.050 190.050 ;
        RECT 676.950 187.950 679.050 190.050 ;
        RECT 667.950 181.950 670.050 184.050 ;
        RECT 659.400 173.400 663.450 174.450 ;
        RECT 655.950 169.950 658.050 172.050 ;
        RECT 656.400 166.050 657.450 169.950 ;
        RECT 659.400 169.050 660.450 173.400 ;
        RECT 658.950 166.950 661.050 169.050 ;
        RECT 662.250 167.250 663.750 168.150 ;
        RECT 664.950 166.950 667.050 169.050 ;
        RECT 671.400 166.050 672.450 187.950 ;
        RECT 677.400 181.050 678.450 187.950 ;
        RECT 680.400 184.050 681.450 196.950 ;
        RECT 679.950 181.950 682.050 184.050 ;
        RECT 676.950 178.950 679.050 181.050 ;
        RECT 683.400 178.050 684.450 196.950 ;
        RECT 686.400 193.050 687.450 196.950 ;
        RECT 688.950 193.950 691.050 196.050 ;
        RECT 685.950 190.950 688.050 193.050 ;
        RECT 689.400 184.050 690.450 193.950 ;
        RECT 692.400 192.450 693.450 205.950 ;
        RECT 695.400 202.050 696.450 205.950 ;
        RECT 694.950 199.950 697.050 202.050 ;
        RECT 695.400 199.050 696.450 199.950 ;
        RECT 698.400 199.050 699.450 211.950 ;
        RECT 701.400 199.050 702.450 214.950 ;
        RECT 704.400 201.450 705.450 232.950 ;
        RECT 707.400 232.050 708.450 235.950 ;
        RECT 712.950 233.850 715.050 234.750 ;
        RECT 718.950 233.850 720.750 234.750 ;
        RECT 721.950 232.950 724.050 235.050 ;
        RECT 725.250 233.850 726.750 234.750 ;
        RECT 727.950 232.950 730.050 235.050 ;
        RECT 706.950 229.950 709.050 232.050 ;
        RECT 715.950 229.950 718.050 232.050 ;
        RECT 721.950 230.850 724.050 231.750 ;
        RECT 724.950 229.950 727.050 232.050 ;
        RECT 707.400 214.050 708.450 229.950 ;
        RECT 706.950 211.950 709.050 214.050 ;
        RECT 712.950 211.950 715.050 214.050 ;
        RECT 704.400 200.400 708.450 201.450 ;
        RECT 694.950 196.950 697.050 199.050 ;
        RECT 697.950 196.950 700.050 199.050 ;
        RECT 700.950 196.950 703.050 199.050 ;
        RECT 704.250 197.250 706.050 198.150 ;
        RECT 694.950 194.850 697.050 195.750 ;
        RECT 697.950 194.250 700.050 195.150 ;
        RECT 700.950 194.850 702.750 195.750 ;
        RECT 703.950 193.950 706.050 196.050 ;
        RECT 707.400 195.450 708.450 200.400 ;
        RECT 713.400 199.050 714.450 211.950 ;
        RECT 716.400 202.050 717.450 229.950 ;
        RECT 725.400 208.050 726.450 229.950 ;
        RECT 728.400 226.050 729.450 232.950 ;
        RECT 731.400 232.050 732.450 253.950 ;
        RECT 734.400 249.450 735.450 259.950 ;
        RECT 737.400 253.050 738.450 268.950 ;
        RECT 740.400 268.050 741.450 271.950 ;
        RECT 742.950 270.450 745.050 271.050 ;
        RECT 745.950 270.450 748.050 271.050 ;
        RECT 742.950 269.400 748.050 270.450 ;
        RECT 742.950 268.950 745.050 269.400 ;
        RECT 745.950 268.950 748.050 269.400 ;
        RECT 739.950 265.950 742.050 268.050 ;
        RECT 746.400 265.050 747.450 268.950 ;
        RECT 749.400 268.050 750.450 271.950 ;
        RECT 751.950 268.950 754.050 271.050 ;
        RECT 755.250 269.850 757.050 270.750 ;
        RECT 748.950 265.950 751.050 268.050 ;
        RECT 754.950 265.950 757.050 268.050 ;
        RECT 745.950 262.950 748.050 265.050 ;
        RECT 751.950 259.950 754.050 262.050 ;
        RECT 736.950 250.950 739.050 253.050 ;
        RECT 734.400 248.400 738.450 249.450 ;
        RECT 733.950 244.950 736.050 247.050 ;
        RECT 734.400 241.050 735.450 244.950 ;
        RECT 737.400 244.050 738.450 248.400 ;
        RECT 736.950 241.950 739.050 244.050 ;
        RECT 733.950 238.950 736.050 241.050 ;
        RECT 739.950 238.950 742.050 241.050 ;
        RECT 745.950 240.450 748.050 241.050 ;
        RECT 748.950 240.450 751.050 241.050 ;
        RECT 745.950 239.400 751.050 240.450 ;
        RECT 745.950 238.950 748.050 239.400 ;
        RECT 748.950 238.950 751.050 239.400 ;
        RECT 730.950 229.950 733.050 232.050 ;
        RECT 734.400 231.450 735.450 238.950 ;
        RECT 736.950 235.950 739.050 238.050 ;
        RECT 740.400 235.050 741.450 238.950 ;
        RECT 742.950 235.950 745.050 238.050 ;
        RECT 746.250 236.250 748.050 237.150 ;
        RECT 748.950 235.950 751.050 238.050 ;
        RECT 736.950 233.850 738.750 234.750 ;
        RECT 739.950 232.950 742.050 235.050 ;
        RECT 743.250 233.850 744.750 234.750 ;
        RECT 745.950 232.950 748.050 235.050 ;
        RECT 734.400 230.400 738.450 231.450 ;
        RECT 739.950 230.850 742.050 231.750 ;
        RECT 733.950 226.950 736.050 229.050 ;
        RECT 737.400 228.450 738.450 230.400 ;
        RECT 742.950 229.950 745.050 232.050 ;
        RECT 737.400 227.400 741.450 228.450 ;
        RECT 727.950 223.950 730.050 226.050 ;
        RECT 734.400 213.450 735.450 226.950 ;
        RECT 731.400 212.400 735.450 213.450 ;
        RECT 721.950 205.950 724.050 208.050 ;
        RECT 724.950 205.950 727.050 208.050 ;
        RECT 715.950 199.950 718.050 202.050 ;
        RECT 718.950 200.250 721.050 201.150 ;
        RECT 709.950 197.250 711.750 198.150 ;
        RECT 712.950 196.950 715.050 199.050 ;
        RECT 716.250 197.250 717.750 198.150 ;
        RECT 718.950 196.950 721.050 199.050 ;
        RECT 719.400 196.050 720.450 196.950 ;
        RECT 709.950 195.450 712.050 196.050 ;
        RECT 707.400 194.400 712.050 195.450 ;
        RECT 713.250 194.850 714.750 195.750 ;
        RECT 709.950 193.950 712.050 194.400 ;
        RECT 715.950 193.950 718.050 196.050 ;
        RECT 718.950 193.950 721.050 196.050 ;
        RECT 692.400 191.400 696.450 192.450 ;
        RECT 685.950 181.950 688.050 184.050 ;
        RECT 688.950 181.950 691.050 184.050 ;
        RECT 682.950 175.950 685.050 178.050 ;
        RECT 676.950 172.950 679.050 175.050 ;
        RECT 682.950 172.950 685.050 175.050 ;
        RECT 673.950 169.950 676.050 172.050 ;
        RECT 655.950 163.950 658.050 166.050 ;
        RECT 659.250 164.850 660.750 165.750 ;
        RECT 661.950 163.950 664.050 166.050 ;
        RECT 665.250 164.850 667.050 165.750 ;
        RECT 670.950 165.450 673.050 166.050 ;
        RECT 668.400 164.400 673.050 165.450 ;
        RECT 655.950 161.850 658.050 162.750 ;
        RECT 658.950 160.950 661.050 163.050 ;
        RECT 652.950 145.950 655.050 148.050 ;
        RECT 649.950 127.950 652.050 130.050 ;
        RECT 659.400 127.050 660.450 160.950 ;
        RECT 662.400 160.050 663.450 163.950 ;
        RECT 664.950 160.950 667.050 163.050 ;
        RECT 661.950 157.950 664.050 160.050 ;
        RECT 665.400 157.050 666.450 160.950 ;
        RECT 668.400 157.050 669.450 164.400 ;
        RECT 670.950 163.950 673.050 164.400 ;
        RECT 674.400 163.050 675.450 169.950 ;
        RECT 677.400 166.050 678.450 172.950 ;
        RECT 676.950 163.950 679.050 166.050 ;
        RECT 680.250 164.250 682.050 165.150 ;
        RECT 670.950 161.850 672.750 162.750 ;
        RECT 673.950 160.950 676.050 163.050 ;
        RECT 677.250 161.850 678.750 162.750 ;
        RECT 679.950 162.450 682.050 163.050 ;
        RECT 683.400 162.450 684.450 172.950 ;
        RECT 679.950 161.400 684.450 162.450 ;
        RECT 679.950 160.950 682.050 161.400 ;
        RECT 673.950 158.850 676.050 159.750 ;
        RECT 664.950 154.950 667.050 157.050 ;
        RECT 667.950 154.950 670.050 157.050 ;
        RECT 670.950 151.950 673.050 154.050 ;
        RECT 673.950 151.950 676.050 154.050 ;
        RECT 661.950 142.950 664.050 145.050 ;
        RECT 662.400 127.050 663.450 142.950 ;
        RECT 671.400 133.050 672.450 151.950 ;
        RECT 667.950 131.250 670.050 132.150 ;
        RECT 670.950 130.950 673.050 133.050 ;
        RECT 674.400 130.050 675.450 151.950 ;
        RECT 682.950 148.950 685.050 151.050 ;
        RECT 676.950 145.950 679.050 148.050 ;
        RECT 677.400 132.450 678.450 145.950 ;
        RECT 679.950 139.950 682.050 142.050 ;
        RECT 680.400 136.050 681.450 139.950 ;
        RECT 679.950 133.950 682.050 136.050 ;
        RECT 677.400 131.400 681.450 132.450 ;
        RECT 664.950 128.250 666.750 129.150 ;
        RECT 667.950 127.950 670.050 130.050 ;
        RECT 671.250 128.250 672.750 129.150 ;
        RECT 673.950 127.950 676.050 130.050 ;
        RECT 676.950 127.950 679.050 130.050 ;
        RECT 649.950 124.950 652.050 127.050 ;
        RECT 652.950 125.250 654.750 126.150 ;
        RECT 655.950 124.950 658.050 127.050 ;
        RECT 658.950 124.950 661.050 127.050 ;
        RECT 661.950 126.450 664.050 127.050 ;
        RECT 664.950 126.450 667.050 127.050 ;
        RECT 661.950 125.400 667.050 126.450 ;
        RECT 661.950 124.950 664.050 125.400 ;
        RECT 664.950 124.950 667.050 125.400 ;
        RECT 646.950 115.950 649.050 118.050 ;
        RECT 650.400 115.050 651.450 124.950 ;
        RECT 652.950 121.950 655.050 124.050 ;
        RECT 656.250 122.850 658.050 123.750 ;
        RECT 658.950 122.250 661.050 123.150 ;
        RECT 661.950 122.850 664.050 123.750 ;
        RECT 649.950 112.950 652.050 115.050 ;
        RECT 646.950 109.950 649.050 112.050 ;
        RECT 647.400 94.050 648.450 109.950 ;
        RECT 653.400 109.050 654.450 121.950 ;
        RECT 668.400 121.050 669.450 127.950 ;
        RECT 670.950 124.950 673.050 127.050 ;
        RECT 674.250 125.850 676.050 126.750 ;
        RECT 677.400 124.050 678.450 127.950 ;
        RECT 676.950 121.950 679.050 124.050 ;
        RECT 658.950 118.950 661.050 121.050 ;
        RECT 667.950 118.950 670.050 121.050 ;
        RECT 680.400 109.050 681.450 131.400 ;
        RECT 683.400 130.050 684.450 148.950 ;
        RECT 686.400 139.050 687.450 181.950 ;
        RECT 695.400 172.050 696.450 191.400 ;
        RECT 697.950 190.950 700.050 193.050 ;
        RECT 698.400 187.050 699.450 190.950 ;
        RECT 697.950 184.950 700.050 187.050 ;
        RECT 698.400 181.050 699.450 184.950 ;
        RECT 697.950 178.950 700.050 181.050 ;
        RECT 704.400 180.450 705.450 193.950 ;
        RECT 712.950 190.950 715.050 193.050 ;
        RECT 713.400 187.050 714.450 190.950 ;
        RECT 706.950 184.950 709.050 187.050 ;
        RECT 712.950 184.950 715.050 187.050 ;
        RECT 701.400 179.400 705.450 180.450 ;
        RECT 691.950 169.950 694.050 172.050 ;
        RECT 694.950 169.950 697.050 172.050 ;
        RECT 697.950 169.950 700.050 172.050 ;
        RECT 698.400 169.050 699.450 169.950 ;
        RECT 688.950 167.250 691.050 168.150 ;
        RECT 691.950 167.850 694.050 168.750 ;
        RECT 694.950 167.250 696.750 168.150 ;
        RECT 697.950 166.950 700.050 169.050 ;
        RECT 688.950 163.950 691.050 166.050 ;
        RECT 691.950 163.950 694.050 166.050 ;
        RECT 694.950 163.950 697.050 166.050 ;
        RECT 698.250 164.850 700.050 165.750 ;
        RECT 692.400 154.050 693.450 163.950 ;
        RECT 695.400 157.050 696.450 163.950 ;
        RECT 697.950 157.950 700.050 160.050 ;
        RECT 694.950 154.950 697.050 157.050 ;
        RECT 691.950 151.950 694.050 154.050 ;
        RECT 685.950 136.950 688.050 139.050 ;
        RECT 688.950 131.250 691.050 132.150 ;
        RECT 698.400 130.050 699.450 157.950 ;
        RECT 701.400 133.050 702.450 179.400 ;
        RECT 703.950 175.950 706.050 178.050 ;
        RECT 704.400 169.050 705.450 175.950 ;
        RECT 707.400 172.050 708.450 184.950 ;
        RECT 712.950 172.950 715.050 175.050 ;
        RECT 706.950 169.950 709.050 172.050 ;
        RECT 703.950 166.950 706.050 169.050 ;
        RECT 707.250 167.250 708.750 168.150 ;
        RECT 709.950 166.950 712.050 169.050 ;
        RECT 713.400 166.050 714.450 172.950 ;
        RECT 703.950 164.850 705.750 165.750 ;
        RECT 706.950 163.950 709.050 166.050 ;
        RECT 710.250 164.850 711.750 165.750 ;
        RECT 712.950 163.950 715.050 166.050 ;
        RECT 712.950 161.850 715.050 162.750 ;
        RECT 700.950 130.950 703.050 133.050 ;
        RECT 706.950 130.950 709.050 133.050 ;
        RECT 682.950 127.950 685.050 130.050 ;
        RECT 686.250 128.250 687.750 129.150 ;
        RECT 688.950 127.950 691.050 130.050 ;
        RECT 692.250 128.250 694.050 129.150 ;
        RECT 697.950 127.950 700.050 130.050 ;
        RECT 703.950 128.250 706.050 129.150 ;
        RECT 682.950 125.850 684.750 126.750 ;
        RECT 685.950 124.950 688.050 127.050 ;
        RECT 689.400 121.050 690.450 127.950 ;
        RECT 698.400 127.050 699.450 127.950 ;
        RECT 691.950 124.950 694.050 127.050 ;
        RECT 694.950 125.250 696.750 126.150 ;
        RECT 697.950 124.950 700.050 127.050 ;
        RECT 701.250 125.250 702.750 126.150 ;
        RECT 703.950 124.950 706.050 127.050 ;
        RECT 692.400 124.050 693.450 124.950 ;
        RECT 704.400 124.050 705.450 124.950 ;
        RECT 691.950 121.950 694.050 124.050 ;
        RECT 694.950 121.950 697.050 124.050 ;
        RECT 698.250 122.850 699.750 123.750 ;
        RECT 700.950 121.950 703.050 124.050 ;
        RECT 703.950 121.950 706.050 124.050 ;
        RECT 688.950 118.950 691.050 121.050 ;
        RECT 701.400 118.050 702.450 121.950 ;
        RECT 700.950 115.950 703.050 118.050 ;
        RECT 694.950 109.950 697.050 112.050 ;
        RECT 652.950 106.950 655.050 109.050 ;
        RECT 679.950 106.950 682.050 109.050 ;
        RECT 661.950 100.950 664.050 103.050 ;
        RECT 676.950 100.950 679.050 103.050 ;
        RECT 682.950 100.950 685.050 103.050 ;
        RECT 655.950 99.450 658.050 100.050 ;
        RECT 650.400 98.400 658.050 99.450 ;
        RECT 650.400 97.050 651.450 98.400 ;
        RECT 655.950 97.950 658.050 98.400 ;
        RECT 662.400 97.050 663.450 100.950 ;
        RECT 667.950 97.950 670.050 100.050 ;
        RECT 673.950 97.950 676.050 100.050 ;
        RECT 668.400 97.050 669.450 97.950 ;
        RECT 649.950 94.950 652.050 97.050 ;
        RECT 655.950 96.450 658.050 97.050 ;
        RECT 653.250 95.250 654.750 96.150 ;
        RECT 655.950 95.400 660.450 96.450 ;
        RECT 655.950 94.950 658.050 95.400 ;
        RECT 646.950 91.950 649.050 94.050 ;
        RECT 650.250 92.850 651.750 93.750 ;
        RECT 652.950 91.950 655.050 94.050 ;
        RECT 656.250 92.850 658.050 93.750 ;
        RECT 646.950 89.850 649.050 90.750 ;
        RECT 659.400 88.050 660.450 95.400 ;
        RECT 661.950 94.950 664.050 97.050 ;
        RECT 665.250 95.250 666.750 96.150 ;
        RECT 667.950 94.950 670.050 97.050 ;
        RECT 661.950 92.850 663.750 93.750 ;
        RECT 664.950 91.950 667.050 94.050 ;
        RECT 668.250 92.850 669.750 93.750 ;
        RECT 670.950 91.950 673.050 94.050 ;
        RECT 670.950 89.850 673.050 90.750 ;
        RECT 658.950 85.950 661.050 88.050 ;
        RECT 658.950 82.950 661.050 85.050 ;
        RECT 659.400 70.050 660.450 82.950 ;
        RECT 658.950 67.950 661.050 70.050 ;
        RECT 649.950 58.950 652.050 61.050 ;
        RECT 650.400 55.050 651.450 58.950 ;
        RECT 674.400 58.050 675.450 97.950 ;
        RECT 677.400 97.050 678.450 100.950 ;
        RECT 683.400 97.050 684.450 100.950 ;
        RECT 676.950 94.950 679.050 97.050 ;
        RECT 680.250 95.250 681.750 96.150 ;
        RECT 682.950 94.950 685.050 97.050 ;
        RECT 695.400 94.050 696.450 109.950 ;
        RECT 703.950 106.950 706.050 109.050 ;
        RECT 697.950 103.950 700.050 106.050 ;
        RECT 698.400 94.050 699.450 103.950 ;
        RECT 676.950 92.850 678.750 93.750 ;
        RECT 679.950 91.950 682.050 94.050 ;
        RECT 683.250 92.850 684.750 93.750 ;
        RECT 685.950 93.450 688.050 94.050 ;
        RECT 691.950 93.450 694.050 94.050 ;
        RECT 685.950 92.400 694.050 93.450 ;
        RECT 685.950 91.950 688.050 92.400 ;
        RECT 685.950 89.850 688.050 90.750 ;
        RECT 689.400 88.050 690.450 92.400 ;
        RECT 691.950 91.950 694.050 92.400 ;
        RECT 694.950 91.950 697.050 94.050 ;
        RECT 697.950 91.950 700.050 94.050 ;
        RECT 701.250 92.250 703.050 93.150 ;
        RECT 695.400 91.050 696.450 91.950 ;
        RECT 691.950 89.850 693.750 90.750 ;
        RECT 694.950 88.950 697.050 91.050 ;
        RECT 698.250 89.850 699.750 90.750 ;
        RECT 700.950 88.950 703.050 91.050 ;
        RECT 688.950 85.950 691.050 88.050 ;
        RECT 694.950 86.850 697.050 87.750 ;
        RECT 701.400 73.050 702.450 88.950 ;
        RECT 704.400 85.050 705.450 106.950 ;
        RECT 703.950 82.950 706.050 85.050 ;
        RECT 694.950 70.950 697.050 73.050 ;
        RECT 700.950 70.950 703.050 73.050 ;
        RECT 691.950 58.950 694.050 61.050 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 664.950 56.250 667.050 57.150 ;
        RECT 673.950 55.950 676.050 58.050 ;
        RECT 659.400 55.050 660.450 55.950 ;
        RECT 692.400 55.050 693.450 58.950 ;
        RECT 695.400 55.050 696.450 70.950 ;
        RECT 707.400 61.050 708.450 130.950 ;
        RECT 716.400 130.050 717.450 193.950 ;
        RECT 722.400 193.050 723.450 205.950 ;
        RECT 731.400 205.050 732.450 212.400 ;
        RECT 736.950 211.950 739.050 214.050 ;
        RECT 733.950 208.950 736.050 211.050 ;
        RECT 727.950 203.250 730.050 204.150 ;
        RECT 730.950 202.950 733.050 205.050 ;
        RECT 734.400 202.050 735.450 208.950 ;
        RECT 724.950 200.250 726.750 201.150 ;
        RECT 727.950 199.950 730.050 202.050 ;
        RECT 731.250 200.250 732.750 201.150 ;
        RECT 733.950 199.950 736.050 202.050 ;
        RECT 724.950 196.950 727.050 199.050 ;
        RECT 721.950 190.950 724.050 193.050 ;
        RECT 721.950 187.950 724.050 190.050 ;
        RECT 722.400 172.050 723.450 187.950 ;
        RECT 725.400 178.050 726.450 196.950 ;
        RECT 724.950 175.950 727.050 178.050 ;
        RECT 728.400 175.050 729.450 199.950 ;
        RECT 730.950 196.950 733.050 199.050 ;
        RECT 734.250 197.850 736.050 198.750 ;
        RECT 731.400 193.050 732.450 196.950 ;
        RECT 733.950 193.950 736.050 196.050 ;
        RECT 730.950 190.950 733.050 193.050 ;
        RECT 730.950 187.950 733.050 190.050 ;
        RECT 731.400 178.050 732.450 187.950 ;
        RECT 730.950 175.950 733.050 178.050 ;
        RECT 727.950 172.950 730.050 175.050 ;
        RECT 721.950 169.950 724.050 172.050 ;
        RECT 730.950 171.450 733.050 172.050 ;
        RECT 734.400 171.450 735.450 193.950 ;
        RECT 730.950 170.400 735.450 171.450 ;
        RECT 737.400 171.450 738.450 211.950 ;
        RECT 740.400 205.050 741.450 227.400 ;
        RECT 743.400 208.050 744.450 229.950 ;
        RECT 746.400 223.050 747.450 232.950 ;
        RECT 749.400 232.050 750.450 235.950 ;
        RECT 748.950 229.950 751.050 232.050 ;
        RECT 748.950 226.950 751.050 229.050 ;
        RECT 745.950 220.950 748.050 223.050 ;
        RECT 745.950 217.950 748.050 220.050 ;
        RECT 746.400 211.050 747.450 217.950 ;
        RECT 749.400 217.050 750.450 226.950 ;
        RECT 752.400 220.050 753.450 259.950 ;
        RECT 751.950 217.950 754.050 220.050 ;
        RECT 748.950 214.950 751.050 217.050 ;
        RECT 755.400 216.450 756.450 265.950 ;
        RECT 761.400 259.050 762.450 292.950 ;
        RECT 764.400 288.450 765.450 331.950 ;
        RECT 764.400 287.400 768.450 288.450 ;
        RECT 763.950 274.950 766.050 277.050 ;
        RECT 764.400 265.050 765.450 274.950 ;
        RECT 763.950 262.950 766.050 265.050 ;
        RECT 763.950 259.950 766.050 262.050 ;
        RECT 760.950 256.950 763.050 259.050 ;
        RECT 760.950 241.950 763.050 244.050 ;
        RECT 761.400 241.050 762.450 241.950 ;
        RECT 760.950 238.950 763.050 241.050 ;
        RECT 761.400 238.050 762.450 238.950 ;
        RECT 764.400 238.050 765.450 259.950 ;
        RECT 767.400 250.050 768.450 287.400 ;
        RECT 770.400 268.050 771.450 391.950 ;
        RECT 769.950 265.950 772.050 268.050 ;
        RECT 769.950 256.950 772.050 259.050 ;
        RECT 766.950 247.950 769.050 250.050 ;
        RECT 757.950 236.250 759.750 237.150 ;
        RECT 760.950 235.950 763.050 238.050 ;
        RECT 763.950 235.950 766.050 238.050 ;
        RECT 766.950 235.950 769.050 238.050 ;
        RECT 764.400 235.050 765.450 235.950 ;
        RECT 757.950 232.950 760.050 235.050 ;
        RECT 761.250 233.850 762.750 234.750 ;
        RECT 763.950 232.950 766.050 235.050 ;
        RECT 767.250 233.850 769.050 234.750 ;
        RECT 760.950 229.950 763.050 232.050 ;
        RECT 763.950 230.850 766.050 231.750 ;
        RECT 766.950 229.950 769.050 232.050 ;
        RECT 757.950 226.950 760.050 229.050 ;
        RECT 758.400 226.050 759.450 226.950 ;
        RECT 757.950 223.950 760.050 226.050 ;
        RECT 752.400 215.400 756.450 216.450 ;
        RECT 748.950 211.950 751.050 214.050 ;
        RECT 745.950 208.950 748.050 211.050 ;
        RECT 742.950 205.950 745.050 208.050 ;
        RECT 746.400 205.050 747.450 208.950 ;
        RECT 739.950 202.950 742.050 205.050 ;
        RECT 742.950 203.250 745.050 204.150 ;
        RECT 745.950 202.950 748.050 205.050 ;
        RECT 749.400 202.050 750.450 211.950 ;
        RECT 739.950 200.250 741.750 201.150 ;
        RECT 742.950 199.950 745.050 202.050 ;
        RECT 746.250 200.250 747.750 201.150 ;
        RECT 748.950 199.950 751.050 202.050 ;
        RECT 743.400 199.050 744.450 199.950 ;
        RECT 739.950 196.950 742.050 199.050 ;
        RECT 742.950 196.950 745.050 199.050 ;
        RECT 745.950 196.950 748.050 199.050 ;
        RECT 749.250 197.850 751.050 198.750 ;
        RECT 740.400 175.050 741.450 196.950 ;
        RECT 742.950 190.950 745.050 193.050 ;
        RECT 739.950 172.950 742.050 175.050 ;
        RECT 737.400 170.400 741.450 171.450 ;
        RECT 730.950 169.950 733.050 170.400 ;
        RECT 721.950 166.950 724.050 169.050 ;
        RECT 724.950 166.950 727.050 169.050 ;
        RECT 728.250 167.250 730.050 168.150 ;
        RECT 730.950 167.850 733.050 168.750 ;
        RECT 733.950 167.250 736.050 168.150 ;
        RECT 736.950 166.950 739.050 169.050 ;
        RECT 722.400 133.050 723.450 166.950 ;
        RECT 724.950 164.850 726.750 165.750 ;
        RECT 727.950 163.950 730.050 166.050 ;
        RECT 730.950 163.950 733.050 166.050 ;
        RECT 733.950 163.950 736.050 166.050 ;
        RECT 728.400 160.050 729.450 163.950 ;
        RECT 727.950 157.950 730.050 160.050 ;
        RECT 731.400 136.050 732.450 163.950 ;
        RECT 734.400 163.050 735.450 163.950 ;
        RECT 733.950 160.950 736.050 163.050 ;
        RECT 737.400 139.050 738.450 166.950 ;
        RECT 736.950 136.950 739.050 139.050 ;
        RECT 730.950 133.950 733.050 136.050 ;
        RECT 721.950 130.950 724.050 133.050 ;
        RECT 727.950 131.250 730.050 132.150 ;
        RECT 709.950 127.950 712.050 130.050 ;
        RECT 715.950 127.950 718.050 130.050 ;
        RECT 724.950 128.250 726.750 129.150 ;
        RECT 727.950 127.950 730.050 130.050 ;
        RECT 733.950 129.450 736.050 130.050 ;
        RECT 731.250 128.250 732.750 129.150 ;
        RECT 733.950 128.400 738.450 129.450 ;
        RECT 733.950 127.950 736.050 128.400 ;
        RECT 710.400 123.450 711.450 127.950 ;
        RECT 716.400 127.050 717.450 127.950 ;
        RECT 728.400 127.050 729.450 127.950 ;
        RECT 712.950 125.250 714.750 126.150 ;
        RECT 715.950 124.950 718.050 127.050 ;
        RECT 721.950 124.950 724.050 127.050 ;
        RECT 724.950 124.950 727.050 127.050 ;
        RECT 727.950 124.950 730.050 127.050 ;
        RECT 730.950 124.950 733.050 127.050 ;
        RECT 734.250 125.850 736.050 126.750 ;
        RECT 712.950 123.450 715.050 124.050 ;
        RECT 710.400 122.400 715.050 123.450 ;
        RECT 716.250 122.850 718.050 123.750 ;
        RECT 712.950 121.950 715.050 122.400 ;
        RECT 718.950 122.250 721.050 123.150 ;
        RECT 721.950 122.850 724.050 123.750 ;
        RECT 725.400 121.050 726.450 124.950 ;
        RECT 718.950 118.950 721.050 121.050 ;
        RECT 724.950 118.950 727.050 121.050 ;
        RECT 712.950 103.950 715.050 106.050 ;
        RECT 709.950 91.950 712.050 94.050 ;
        RECT 713.400 91.050 714.450 103.950 ;
        RECT 715.950 94.950 718.050 97.050 ;
        RECT 721.950 94.950 724.050 97.050 ;
        RECT 716.400 94.050 717.450 94.950 ;
        RECT 715.950 91.950 718.050 94.050 ;
        RECT 719.250 92.250 721.050 93.150 ;
        RECT 709.950 89.850 711.750 90.750 ;
        RECT 712.950 88.950 715.050 91.050 ;
        RECT 716.250 89.850 717.750 90.750 ;
        RECT 718.950 88.950 721.050 91.050 ;
        RECT 712.950 86.850 715.050 87.750 ;
        RECT 715.950 85.950 718.050 88.050 ;
        RECT 703.950 59.250 706.050 60.150 ;
        RECT 706.950 58.950 709.050 61.050 ;
        RECT 697.950 55.950 700.050 58.050 ;
        RECT 700.950 56.250 702.750 57.150 ;
        RECT 703.950 55.950 706.050 58.050 ;
        RECT 709.950 57.450 712.050 58.050 ;
        RECT 707.250 56.250 708.750 57.150 ;
        RECT 709.950 56.400 714.450 57.450 ;
        RECT 709.950 55.950 712.050 56.400 ;
        RECT 698.400 55.050 699.450 55.950 ;
        RECT 649.950 52.950 652.050 55.050 ;
        RECT 655.950 53.250 657.750 54.150 ;
        RECT 658.950 52.950 661.050 55.050 ;
        RECT 662.250 53.250 663.750 54.150 ;
        RECT 664.950 52.950 667.050 55.050 ;
        RECT 673.950 53.250 675.750 54.150 ;
        RECT 676.950 52.950 679.050 55.050 ;
        RECT 682.950 52.950 685.050 55.050 ;
        RECT 688.950 53.250 690.750 54.150 ;
        RECT 691.950 52.950 694.050 55.050 ;
        RECT 694.950 52.950 697.050 55.050 ;
        RECT 697.950 52.950 700.050 55.050 ;
        RECT 700.950 52.950 703.050 55.050 ;
        RECT 706.950 52.950 709.050 55.050 ;
        RECT 710.250 53.850 712.050 54.750 ;
        RECT 646.950 50.250 649.050 51.150 ;
        RECT 649.950 50.850 652.050 51.750 ;
        RECT 655.950 49.950 658.050 52.050 ;
        RECT 659.250 50.850 660.750 51.750 ;
        RECT 661.950 49.950 664.050 52.050 ;
        RECT 673.950 49.950 676.050 52.050 ;
        RECT 677.250 50.850 679.050 51.750 ;
        RECT 679.950 50.250 682.050 51.150 ;
        RECT 682.950 50.850 685.050 51.750 ;
        RECT 688.950 49.950 691.050 52.050 ;
        RECT 692.250 50.850 694.050 51.750 ;
        RECT 694.950 50.250 697.050 51.150 ;
        RECT 697.950 50.850 700.050 51.750 ;
        RECT 646.950 46.950 649.050 49.050 ;
        RECT 649.950 46.950 652.050 49.050 ;
        RECT 647.400 46.050 648.450 46.950 ;
        RECT 646.950 43.950 649.050 46.050 ;
        RECT 643.950 22.950 646.050 25.050 ;
        RECT 650.400 22.050 651.450 46.950 ;
        RECT 662.400 31.050 663.450 49.950 ;
        RECT 674.400 43.050 675.450 49.950 ;
        RECT 679.950 46.950 682.050 49.050 ;
        RECT 680.400 46.050 681.450 46.950 ;
        RECT 679.950 43.950 682.050 46.050 ;
        RECT 673.950 40.950 676.050 43.050 ;
        RECT 661.950 28.950 664.050 31.050 ;
        RECT 685.950 28.950 688.050 31.050 ;
        RECT 622.950 19.950 625.050 22.050 ;
        RECT 625.950 19.950 628.050 22.050 ;
        RECT 631.950 19.950 634.050 22.050 ;
        RECT 635.250 20.250 637.050 21.150 ;
        RECT 640.950 20.250 642.750 21.150 ;
        RECT 643.950 19.950 646.050 22.050 ;
        RECT 647.250 20.250 649.050 21.150 ;
        RECT 649.950 19.950 652.050 22.050 ;
        RECT 658.950 21.450 661.050 22.050 ;
        RECT 662.400 21.450 663.450 28.950 ;
        RECT 670.950 25.950 673.050 28.050 ;
        RECT 670.950 23.850 673.050 24.750 ;
        RECT 673.950 23.250 676.050 24.150 ;
        RECT 682.950 22.950 685.050 25.050 ;
        RECT 683.400 22.050 684.450 22.950 ;
        RECT 655.950 20.250 657.750 21.150 ;
        RECT 658.950 20.400 663.450 21.450 ;
        RECT 658.950 19.950 661.050 20.400 ;
        RECT 664.950 19.950 667.050 22.050 ;
        RECT 673.950 19.950 676.050 22.050 ;
        RECT 682.950 19.950 685.050 22.050 ;
        RECT 686.400 21.450 687.450 28.950 ;
        RECT 689.400 28.050 690.450 49.950 ;
        RECT 701.400 49.050 702.450 52.950 ;
        RECT 713.400 52.050 714.450 56.400 ;
        RECT 712.950 49.950 715.050 52.050 ;
        RECT 694.950 46.950 697.050 49.050 ;
        RECT 700.950 46.950 703.050 49.050 ;
        RECT 716.400 43.050 717.450 85.950 ;
        RECT 722.400 60.450 723.450 94.950 ;
        RECT 725.400 61.050 726.450 118.950 ;
        RECT 728.400 100.050 729.450 124.950 ;
        RECT 737.400 124.050 738.450 128.400 ;
        RECT 740.400 124.050 741.450 170.400 ;
        RECT 743.400 169.050 744.450 190.950 ;
        RECT 746.400 190.050 747.450 196.950 ;
        RECT 748.950 193.950 751.050 196.050 ;
        RECT 745.950 187.950 748.050 190.050 ;
        RECT 746.400 181.050 747.450 187.950 ;
        RECT 745.950 178.950 748.050 181.050 ;
        RECT 749.400 174.450 750.450 193.950 ;
        RECT 752.400 181.050 753.450 215.400 ;
        RECT 754.950 205.950 757.050 208.050 ;
        RECT 755.400 193.050 756.450 205.950 ;
        RECT 758.400 204.450 759.450 223.950 ;
        RECT 761.400 214.050 762.450 229.950 ;
        RECT 763.950 214.950 766.050 217.050 ;
        RECT 760.950 211.950 763.050 214.050 ;
        RECT 764.400 205.050 765.450 214.950 ;
        RECT 758.400 203.400 762.450 204.450 ;
        RECT 761.400 201.450 762.450 203.400 ;
        RECT 763.950 202.950 766.050 205.050 ;
        RECT 767.400 202.050 768.450 229.950 ;
        RECT 770.400 226.050 771.450 256.950 ;
        RECT 769.950 223.950 772.050 226.050 ;
        RECT 769.950 211.950 772.050 214.050 ;
        RECT 757.950 200.250 760.050 201.150 ;
        RECT 761.400 200.400 765.450 201.450 ;
        RECT 764.400 199.050 765.450 200.400 ;
        RECT 766.950 199.950 769.050 202.050 ;
        RECT 757.950 196.950 760.050 199.050 ;
        RECT 761.250 197.250 762.750 198.150 ;
        RECT 763.950 196.950 766.050 199.050 ;
        RECT 767.250 197.250 769.050 198.150 ;
        RECT 754.950 190.950 757.050 193.050 ;
        RECT 758.400 190.050 759.450 196.950 ;
        RECT 760.950 193.950 763.050 196.050 ;
        RECT 764.250 194.850 765.750 195.750 ;
        RECT 766.950 193.950 769.050 196.050 ;
        RECT 761.400 192.450 762.450 193.950 ;
        RECT 761.400 191.400 765.450 192.450 ;
        RECT 757.950 187.950 760.050 190.050 ;
        RECT 760.950 187.950 763.050 190.050 ;
        RECT 761.400 183.450 762.450 187.950 ;
        RECT 764.400 184.050 765.450 191.400 ;
        RECT 767.400 187.050 768.450 193.950 ;
        RECT 766.950 184.950 769.050 187.050 ;
        RECT 758.400 182.400 762.450 183.450 ;
        RECT 751.950 178.950 754.050 181.050 ;
        RECT 754.950 175.950 757.050 178.050 ;
        RECT 749.400 173.400 753.450 174.450 ;
        RECT 748.950 169.950 751.050 172.050 ;
        RECT 742.950 166.950 745.050 169.050 ;
        RECT 742.950 164.250 744.750 165.150 ;
        RECT 745.950 163.950 748.050 166.050 ;
        RECT 749.400 163.050 750.450 169.950 ;
        RECT 752.400 166.050 753.450 173.400 ;
        RECT 751.950 163.950 754.050 166.050 ;
        RECT 755.400 163.050 756.450 175.950 ;
        RECT 742.950 160.950 745.050 163.050 ;
        RECT 746.250 161.850 747.750 162.750 ;
        RECT 748.950 160.950 751.050 163.050 ;
        RECT 752.250 161.850 754.050 162.750 ;
        RECT 754.950 160.950 757.050 163.050 ;
        RECT 748.950 158.850 751.050 159.750 ;
        RECT 758.400 154.050 759.450 182.400 ;
        RECT 763.950 181.950 766.050 184.050 ;
        RECT 766.950 181.950 769.050 184.050 ;
        RECT 760.950 178.950 763.050 181.050 ;
        RECT 748.950 151.950 751.050 154.050 ;
        RECT 757.950 151.950 760.050 154.050 ;
        RECT 742.950 130.950 745.050 133.050 ;
        RECT 736.950 121.950 739.050 124.050 ;
        RECT 739.950 121.950 742.050 124.050 ;
        RECT 727.950 97.950 730.050 100.050 ;
        RECT 733.950 97.950 736.050 100.050 ;
        RECT 739.950 97.950 742.050 100.050 ;
        RECT 740.400 97.050 741.450 97.950 ;
        RECT 727.950 94.950 730.050 97.050 ;
        RECT 731.250 95.250 733.050 96.150 ;
        RECT 733.950 95.850 736.050 96.750 ;
        RECT 736.950 95.250 739.050 96.150 ;
        RECT 739.950 94.950 742.050 97.050 ;
        RECT 740.400 94.050 741.450 94.950 ;
        RECT 727.950 92.850 729.750 93.750 ;
        RECT 730.950 91.950 733.050 94.050 ;
        RECT 736.950 91.950 739.050 94.050 ;
        RECT 739.950 91.950 742.050 94.050 ;
        RECT 731.400 91.050 732.450 91.950 ;
        RECT 743.400 91.050 744.450 130.950 ;
        RECT 749.400 127.050 750.450 151.950 ;
        RECT 757.950 145.950 760.050 148.050 ;
        RECT 754.950 136.950 757.050 139.050 ;
        RECT 755.400 127.050 756.450 136.950 ;
        RECT 745.950 125.250 747.750 126.150 ;
        RECT 748.950 124.950 751.050 127.050 ;
        RECT 754.950 124.950 757.050 127.050 ;
        RECT 745.950 121.950 748.050 124.050 ;
        RECT 749.250 122.850 751.050 123.750 ;
        RECT 751.950 122.250 754.050 123.150 ;
        RECT 754.950 122.850 757.050 123.750 ;
        RECT 758.400 121.050 759.450 145.950 ;
        RECT 751.950 118.950 754.050 121.050 ;
        RECT 757.950 118.950 760.050 121.050 ;
        RECT 751.950 112.950 754.050 115.050 ;
        RECT 745.950 100.950 748.050 103.050 ;
        RECT 746.400 94.050 747.450 100.950 ;
        RECT 745.950 91.950 748.050 94.050 ;
        RECT 749.250 92.250 751.050 93.150 ;
        RECT 730.950 88.950 733.050 91.050 ;
        RECT 739.950 89.850 741.750 90.750 ;
        RECT 742.950 88.950 745.050 91.050 ;
        RECT 746.250 89.850 747.750 90.750 ;
        RECT 748.950 88.950 751.050 91.050 ;
        RECT 742.950 86.850 745.050 87.750 ;
        RECT 749.400 87.450 750.450 88.950 ;
        RECT 746.400 86.400 750.450 87.450 ;
        RECT 746.400 61.050 747.450 86.400 ;
        RECT 748.950 82.950 751.050 85.050 ;
        RECT 719.400 59.400 723.450 60.450 ;
        RECT 715.950 40.950 718.050 43.050 ;
        RECT 715.950 34.950 718.050 37.050 ;
        RECT 709.950 28.950 712.050 31.050 ;
        RECT 688.950 25.950 691.050 28.050 ;
        RECT 710.400 25.050 711.450 28.950 ;
        RECT 716.400 25.050 717.450 34.950 ;
        RECT 719.400 25.050 720.450 59.400 ;
        RECT 724.950 58.950 727.050 61.050 ;
        RECT 727.950 59.250 730.050 60.150 ;
        RECT 736.950 59.250 739.050 60.150 ;
        RECT 745.950 58.950 748.050 61.050 ;
        RECT 721.950 55.950 724.050 58.050 ;
        RECT 725.250 56.250 726.750 57.150 ;
        RECT 727.950 55.950 730.050 58.050 ;
        RECT 731.250 56.250 733.050 57.150 ;
        RECT 733.950 56.250 735.750 57.150 ;
        RECT 736.950 55.950 739.050 58.050 ;
        RECT 740.250 56.250 741.750 57.150 ;
        RECT 742.950 55.950 745.050 58.050 ;
        RECT 721.950 53.850 723.750 54.750 ;
        RECT 724.950 52.950 727.050 55.050 ;
        RECT 700.950 22.950 703.050 25.050 ;
        RECT 709.950 22.950 712.050 25.050 ;
        RECT 713.250 23.250 714.750 24.150 ;
        RECT 715.950 22.950 718.050 25.050 ;
        RECT 718.950 22.950 721.050 25.050 ;
        RECT 701.400 22.050 702.450 22.950 ;
        RECT 725.400 22.050 726.450 52.950 ;
        RECT 728.400 52.050 729.450 55.950 ;
        RECT 730.950 52.950 733.050 55.050 ;
        RECT 733.950 52.950 736.050 55.050 ;
        RECT 727.950 49.950 730.050 52.050 ;
        RECT 731.400 46.050 732.450 52.950 ;
        RECT 730.950 43.950 733.050 46.050 ;
        RECT 730.950 40.950 733.050 43.050 ;
        RECT 727.950 28.950 730.050 31.050 ;
        RECT 728.400 22.050 729.450 28.950 ;
        RECT 731.400 25.050 732.450 40.950 ;
        RECT 734.400 31.050 735.450 52.950 ;
        RECT 737.400 52.050 738.450 55.950 ;
        RECT 749.400 55.050 750.450 82.950 ;
        RECT 752.400 55.050 753.450 112.950 ;
        RECT 761.400 58.050 762.450 178.950 ;
        RECT 764.400 166.050 765.450 181.950 ;
        RECT 763.950 163.950 766.050 166.050 ;
        RECT 767.400 160.050 768.450 181.950 ;
        RECT 766.950 157.950 769.050 160.050 ;
        RECT 770.400 148.050 771.450 211.950 ;
        RECT 769.950 145.950 772.050 148.050 ;
        RECT 763.950 133.950 766.050 136.050 ;
        RECT 760.950 55.950 763.050 58.050 ;
        RECT 739.950 52.950 742.050 55.050 ;
        RECT 743.250 53.850 745.050 54.750 ;
        RECT 748.950 54.450 751.050 55.050 ;
        RECT 746.400 53.400 751.050 54.450 ;
        RECT 736.950 49.950 739.050 52.050 ;
        RECT 733.950 28.950 736.050 31.050 ;
        RECT 746.400 25.050 747.450 53.400 ;
        RECT 748.950 52.950 751.050 53.400 ;
        RECT 751.950 52.950 754.050 55.050 ;
        RECT 754.950 52.950 757.050 55.050 ;
        RECT 758.250 53.250 760.050 54.150 ;
        RECT 748.950 50.850 751.050 51.750 ;
        RECT 751.950 50.250 754.050 51.150 ;
        RECT 754.950 50.850 756.750 51.750 ;
        RECT 757.950 49.950 760.050 52.050 ;
        RECT 761.400 49.050 762.450 55.950 ;
        RECT 764.400 55.050 765.450 133.950 ;
        RECT 763.950 52.950 766.050 55.050 ;
        RECT 751.950 46.950 754.050 49.050 ;
        RECT 760.950 46.950 763.050 49.050 ;
        RECT 748.950 43.950 751.050 46.050 ;
        RECT 730.950 22.950 733.050 25.050 ;
        RECT 734.250 23.250 735.750 24.150 ;
        RECT 736.950 22.950 739.050 25.050 ;
        RECT 739.950 22.950 742.050 25.050 ;
        RECT 743.250 23.250 744.750 24.150 ;
        RECT 745.950 22.950 748.050 25.050 ;
        RECT 749.400 22.050 750.450 43.950 ;
        RECT 688.950 21.450 691.050 22.050 ;
        RECT 686.400 20.400 691.050 21.450 ;
        RECT 688.950 19.950 691.050 20.400 ;
        RECT 692.250 20.250 694.050 21.150 ;
        RECT 697.950 20.250 699.750 21.150 ;
        RECT 700.950 19.950 703.050 22.050 ;
        RECT 704.250 20.250 706.050 21.150 ;
        RECT 709.950 20.850 711.750 21.750 ;
        RECT 712.950 19.950 715.050 22.050 ;
        RECT 716.250 20.850 717.750 21.750 ;
        RECT 718.950 19.950 721.050 22.050 ;
        RECT 724.950 19.950 727.050 22.050 ;
        RECT 727.950 19.950 730.050 22.050 ;
        RECT 731.250 20.850 732.750 21.750 ;
        RECT 733.950 19.950 736.050 22.050 ;
        RECT 737.250 20.850 739.050 21.750 ;
        RECT 739.950 20.850 741.750 21.750 ;
        RECT 742.950 19.950 745.050 22.050 ;
        RECT 746.250 20.850 747.750 21.750 ;
        RECT 748.950 19.950 751.050 22.050 ;
        RECT 601.950 16.950 604.050 17.400 ;
        RECT 607.950 17.400 612.450 18.450 ;
        RECT 607.950 16.950 610.050 17.400 ;
        RECT 613.950 16.950 616.050 19.050 ;
        RECT 617.250 17.850 618.750 18.750 ;
        RECT 619.950 16.950 622.050 19.050 ;
        RECT 623.250 17.850 625.050 18.750 ;
        RECT 625.950 17.850 627.750 18.750 ;
        RECT 628.950 16.950 631.050 19.050 ;
        RECT 632.250 17.850 633.750 18.750 ;
        RECT 634.950 18.450 637.050 19.050 ;
        RECT 640.950 18.450 643.050 19.050 ;
        RECT 634.950 17.400 643.050 18.450 ;
        RECT 644.250 17.850 645.750 18.750 ;
        RECT 634.950 16.950 637.050 17.400 ;
        RECT 640.950 16.950 643.050 17.400 ;
        RECT 646.950 16.950 649.050 19.050 ;
        RECT 655.950 16.950 658.050 19.050 ;
        RECT 659.250 17.850 660.750 18.750 ;
        RECT 661.950 16.950 664.050 19.050 ;
        RECT 665.250 17.850 667.050 18.750 ;
        RECT 682.950 17.850 684.750 18.750 ;
        RECT 685.950 16.950 688.050 19.050 ;
        RECT 689.250 17.850 690.750 18.750 ;
        RECT 691.950 16.950 694.050 19.050 ;
        RECT 697.950 16.950 700.050 19.050 ;
        RECT 701.250 17.850 702.750 18.750 ;
        RECT 703.950 16.950 706.050 19.050 ;
        RECT 718.950 17.850 721.050 18.750 ;
        RECT 727.950 17.850 730.050 18.750 ;
        RECT 748.950 17.850 751.050 18.750 ;
        RECT 590.400 16.050 591.450 16.950 ;
        RECT 614.400 16.050 615.450 16.950 ;
        RECT 647.400 16.050 648.450 16.950 ;
        RECT 187.950 14.850 190.050 15.750 ;
        RECT 202.950 14.850 205.050 15.750 ;
        RECT 250.950 14.850 253.050 15.750 ;
        RECT 295.950 14.850 298.050 15.750 ;
        RECT 331.950 14.850 334.050 15.750 ;
        RECT 559.950 14.850 562.050 15.750 ;
        RECT 589.950 13.950 592.050 16.050 ;
        RECT 613.950 13.950 616.050 16.050 ;
        RECT 619.950 14.850 622.050 15.750 ;
        RECT 628.950 14.850 631.050 15.750 ;
        RECT 646.950 13.950 649.050 16.050 ;
        RECT 652.950 15.450 655.050 16.050 ;
        RECT 656.400 15.450 657.450 16.950 ;
        RECT 652.950 14.400 657.450 15.450 ;
        RECT 661.950 14.850 664.050 15.750 ;
        RECT 685.950 14.850 688.050 15.750 ;
        RECT 652.950 13.950 655.050 14.400 ;
        RECT 614.400 13.050 615.450 13.950 ;
        RECT 698.400 13.050 699.450 16.950 ;
        RECT 106.950 10.950 109.050 13.050 ;
        RECT 145.950 10.950 148.050 13.050 ;
        RECT 613.950 10.950 616.050 13.050 ;
        RECT 697.950 10.950 700.050 13.050 ;
      LAYER metal3 ;
        RECT 103.950 714.600 106.050 715.050 ;
        RECT 115.950 714.600 118.050 715.050 ;
        RECT 370.950 714.600 373.050 715.050 ;
        RECT 103.950 713.400 373.050 714.600 ;
        RECT 103.950 712.950 106.050 713.400 ;
        RECT 115.950 712.950 118.050 713.400 ;
        RECT 370.950 712.950 373.050 713.400 ;
        RECT 238.950 711.600 241.050 712.050 ;
        RECT 358.950 711.600 361.050 712.050 ;
        RECT 238.950 710.400 361.050 711.600 ;
        RECT 238.950 709.950 241.050 710.400 ;
        RECT 358.950 709.950 361.050 710.400 ;
        RECT 31.950 708.600 34.050 709.050 ;
        RECT 109.950 708.600 112.050 709.050 ;
        RECT 148.950 708.600 151.050 709.050 ;
        RECT 217.950 708.600 220.050 709.050 ;
        RECT 277.950 708.600 280.050 709.050 ;
        RECT 298.950 708.600 301.050 709.050 ;
        RECT 31.950 707.400 301.050 708.600 ;
        RECT 31.950 706.950 34.050 707.400 ;
        RECT 109.950 706.950 112.050 707.400 ;
        RECT 148.950 706.950 151.050 707.400 ;
        RECT 217.950 706.950 220.050 707.400 ;
        RECT 277.950 706.950 280.050 707.400 ;
        RECT 298.950 706.950 301.050 707.400 ;
        RECT 307.950 708.600 310.050 709.050 ;
        RECT 328.950 708.600 331.050 709.050 ;
        RECT 307.950 707.400 331.050 708.600 ;
        RECT 307.950 706.950 310.050 707.400 ;
        RECT 328.950 706.950 331.050 707.400 ;
        RECT 166.950 705.600 169.050 706.050 ;
        RECT 187.950 705.600 190.050 706.050 ;
        RECT 166.950 704.400 190.050 705.600 ;
        RECT 166.950 703.950 169.050 704.400 ;
        RECT 187.950 703.950 190.050 704.400 ;
        RECT 196.950 705.600 199.050 706.050 ;
        RECT 262.950 705.600 265.050 706.050 ;
        RECT 334.950 705.600 337.050 706.050 ;
        RECT 382.950 705.600 385.050 706.050 ;
        RECT 196.950 704.400 265.050 705.600 ;
        RECT 196.950 703.950 199.050 704.400 ;
        RECT 262.950 703.950 265.050 704.400 ;
        RECT 305.400 704.400 337.050 705.600 ;
        RECT 25.950 702.600 28.050 703.050 ;
        RECT 40.950 702.600 43.050 703.050 ;
        RECT 25.950 701.400 43.050 702.600 ;
        RECT 25.950 700.950 28.050 701.400 ;
        RECT 40.950 700.950 43.050 701.400 ;
        RECT 46.950 702.600 49.050 703.050 ;
        RECT 52.950 702.600 55.050 703.050 ;
        RECT 73.950 702.600 76.050 703.050 ;
        RECT 46.950 701.400 76.050 702.600 ;
        RECT 46.950 700.950 49.050 701.400 ;
        RECT 52.950 700.950 55.050 701.400 ;
        RECT 73.950 700.950 76.050 701.400 ;
        RECT 79.950 702.600 82.050 703.050 ;
        RECT 85.950 702.600 88.050 703.050 ;
        RECT 79.950 701.400 88.050 702.600 ;
        RECT 79.950 700.950 82.050 701.400 ;
        RECT 85.950 700.950 88.050 701.400 ;
        RECT 97.950 702.600 100.050 703.050 ;
        RECT 109.950 702.600 112.050 703.050 ;
        RECT 97.950 701.400 112.050 702.600 ;
        RECT 97.950 700.950 100.050 701.400 ;
        RECT 109.950 700.950 112.050 701.400 ;
        RECT 112.950 702.600 115.050 703.050 ;
        RECT 142.950 702.600 145.050 703.050 ;
        RECT 112.950 701.400 145.050 702.600 ;
        RECT 112.950 700.950 115.050 701.400 ;
        RECT 13.950 699.600 16.050 700.050 ;
        RECT 25.950 699.600 28.050 700.050 ;
        RECT 13.950 698.400 28.050 699.600 ;
        RECT 13.950 697.950 16.050 698.400 ;
        RECT 25.950 697.950 28.050 698.400 ;
        RECT 58.950 699.600 61.050 700.050 ;
        RECT 70.950 699.600 73.050 700.050 ;
        RECT 58.950 698.400 73.050 699.600 ;
        RECT 74.400 699.600 75.600 700.950 ;
        RECT 125.400 700.050 126.600 701.400 ;
        RECT 142.950 700.950 145.050 701.400 ;
        RECT 178.950 700.950 181.050 703.050 ;
        RECT 199.950 702.600 202.050 703.050 ;
        RECT 214.950 702.600 217.050 703.050 ;
        RECT 229.950 702.600 232.050 703.050 ;
        RECT 199.950 701.400 217.050 702.600 ;
        RECT 199.950 700.950 202.050 701.400 ;
        RECT 214.950 700.950 217.050 701.400 ;
        RECT 221.400 701.400 232.050 702.600 ;
        RECT 82.950 699.600 85.050 700.050 ;
        RECT 94.950 699.600 97.050 700.050 ;
        RECT 100.950 699.600 103.050 700.050 ;
        RECT 74.400 698.400 85.050 699.600 ;
        RECT 58.950 697.950 61.050 698.400 ;
        RECT 70.950 697.950 73.050 698.400 ;
        RECT 82.950 697.950 85.050 698.400 ;
        RECT 86.400 698.400 97.050 699.600 ;
        RECT 4.950 696.600 7.050 697.050 ;
        RECT 28.950 696.600 31.050 697.050 ;
        RECT 4.950 695.400 31.050 696.600 ;
        RECT 4.950 694.950 7.050 695.400 ;
        RECT 28.950 694.950 31.050 695.400 ;
        RECT 34.950 696.600 37.050 697.050 ;
        RECT 86.400 696.600 87.600 698.400 ;
        RECT 94.950 697.950 97.050 698.400 ;
        RECT 98.400 698.400 103.050 699.600 ;
        RECT 34.950 695.400 87.600 696.600 ;
        RECT 91.950 696.600 94.050 697.050 ;
        RECT 98.400 696.600 99.600 698.400 ;
        RECT 100.950 697.950 103.050 698.400 ;
        RECT 124.950 697.950 127.050 700.050 ;
        RECT 133.950 699.600 136.050 700.050 ;
        RECT 145.950 699.600 148.050 700.050 ;
        RECT 133.950 698.400 148.050 699.600 ;
        RECT 133.950 697.950 136.050 698.400 ;
        RECT 145.950 697.950 148.050 698.400 ;
        RECT 151.950 699.600 154.050 700.050 ;
        RECT 160.950 699.600 163.050 700.050 ;
        RECT 179.400 699.600 180.600 700.950 ;
        RECT 221.400 700.050 222.600 701.400 ;
        RECT 229.950 700.950 232.050 701.400 ;
        RECT 247.950 702.600 250.050 703.050 ;
        RECT 247.950 701.400 279.600 702.600 ;
        RECT 247.950 700.950 250.050 701.400 ;
        RECT 260.400 700.050 261.600 701.400 ;
        RECT 184.950 699.600 187.050 700.050 ;
        RECT 151.950 698.400 187.050 699.600 ;
        RECT 151.950 697.950 154.050 698.400 ;
        RECT 160.950 697.950 163.050 698.400 ;
        RECT 184.950 697.950 187.050 698.400 ;
        RECT 193.950 699.600 196.050 700.050 ;
        RECT 202.950 699.600 205.050 700.050 ;
        RECT 217.950 699.600 220.050 700.050 ;
        RECT 193.950 698.400 220.050 699.600 ;
        RECT 193.950 697.950 196.050 698.400 ;
        RECT 202.950 697.950 205.050 698.400 ;
        RECT 217.950 697.950 220.050 698.400 ;
        RECT 220.950 697.950 223.050 700.050 ;
        RECT 244.950 699.600 247.050 700.050 ;
        RECT 224.400 698.400 247.050 699.600 ;
        RECT 91.950 695.400 99.600 696.600 ;
        RECT 100.950 696.600 103.050 697.050 ;
        RECT 106.950 696.600 109.050 697.050 ;
        RECT 151.950 696.600 154.050 697.050 ;
        RECT 100.950 695.400 154.050 696.600 ;
        RECT 34.950 694.950 37.050 695.400 ;
        RECT 91.950 694.950 94.050 695.400 ;
        RECT 100.950 694.950 103.050 695.400 ;
        RECT 106.950 694.950 109.050 695.400 ;
        RECT 151.950 694.950 154.050 695.400 ;
        RECT 181.950 696.600 184.050 697.050 ;
        RECT 190.950 696.600 193.050 697.050 ;
        RECT 181.950 695.400 193.050 696.600 ;
        RECT 181.950 694.950 184.050 695.400 ;
        RECT 190.950 694.950 193.050 695.400 ;
        RECT 211.950 696.600 214.050 697.050 ;
        RECT 224.400 696.600 225.600 698.400 ;
        RECT 244.950 697.950 247.050 698.400 ;
        RECT 259.950 697.950 262.050 700.050 ;
        RECT 265.950 699.600 268.050 700.050 ;
        RECT 274.950 699.600 277.050 700.050 ;
        RECT 265.950 698.400 277.050 699.600 ;
        RECT 278.400 699.600 279.600 701.400 ;
        RECT 280.950 699.600 283.050 700.050 ;
        RECT 278.400 698.400 283.050 699.600 ;
        RECT 265.950 697.950 268.050 698.400 ;
        RECT 274.950 697.950 277.050 698.400 ;
        RECT 280.950 697.950 283.050 698.400 ;
        RECT 305.400 697.050 306.600 704.400 ;
        RECT 334.950 703.950 337.050 704.400 ;
        RECT 368.400 704.400 385.050 705.600 ;
        RECT 313.950 700.950 316.050 703.050 ;
        RECT 319.950 700.950 322.050 703.050 ;
        RECT 325.950 702.600 328.050 703.050 ;
        RECT 337.950 702.600 340.050 703.050 ;
        RECT 325.950 701.400 340.050 702.600 ;
        RECT 325.950 700.950 328.050 701.400 ;
        RECT 337.950 700.950 340.050 701.400 ;
        RECT 349.950 702.600 352.050 703.050 ;
        RECT 364.950 702.600 367.050 703.050 ;
        RECT 349.950 701.400 367.050 702.600 ;
        RECT 349.950 700.950 352.050 701.400 ;
        RECT 364.950 700.950 367.050 701.400 ;
        RECT 314.400 699.600 315.600 700.950 ;
        RECT 316.950 699.600 319.050 700.050 ;
        RECT 314.400 698.400 319.050 699.600 ;
        RECT 316.950 697.950 319.050 698.400 ;
        RECT 211.950 695.400 225.600 696.600 ;
        RECT 232.950 696.600 235.050 697.050 ;
        RECT 256.950 696.600 259.050 697.050 ;
        RECT 232.950 695.400 259.050 696.600 ;
        RECT 211.950 694.950 214.050 695.400 ;
        RECT 232.950 694.950 235.050 695.400 ;
        RECT 256.950 694.950 259.050 695.400 ;
        RECT 262.950 696.600 265.050 697.050 ;
        RECT 292.950 696.600 295.050 697.050 ;
        RECT 262.950 695.400 295.050 696.600 ;
        RECT 262.950 694.950 265.050 695.400 ;
        RECT 292.950 694.950 295.050 695.400 ;
        RECT 304.950 694.950 307.050 697.050 ;
        RECT 310.950 696.600 313.050 697.050 ;
        RECT 320.400 696.600 321.600 700.950 ;
        RECT 368.400 700.050 369.600 704.400 ;
        RECT 382.950 703.950 385.050 704.400 ;
        RECT 400.950 705.600 403.050 706.050 ;
        RECT 523.950 705.600 526.050 706.050 ;
        RECT 538.950 705.600 541.050 706.050 ;
        RECT 544.950 705.600 547.050 706.050 ;
        RECT 400.950 704.400 547.050 705.600 ;
        RECT 400.950 703.950 403.050 704.400 ;
        RECT 523.950 703.950 526.050 704.400 ;
        RECT 538.950 703.950 541.050 704.400 ;
        RECT 544.950 703.950 547.050 704.400 ;
        RECT 370.950 702.600 373.050 703.050 ;
        RECT 376.950 702.600 379.050 703.050 ;
        RECT 370.950 701.400 379.050 702.600 ;
        RECT 370.950 700.950 373.050 701.400 ;
        RECT 376.950 700.950 379.050 701.400 ;
        RECT 388.950 702.600 391.050 703.050 ;
        RECT 397.950 702.600 400.050 703.050 ;
        RECT 388.950 701.400 400.050 702.600 ;
        RECT 388.950 700.950 391.050 701.400 ;
        RECT 397.950 700.950 400.050 701.400 ;
        RECT 478.950 702.600 481.050 703.050 ;
        RECT 484.950 702.600 487.050 703.050 ;
        RECT 478.950 701.400 487.050 702.600 ;
        RECT 478.950 700.950 481.050 701.400 ;
        RECT 484.950 700.950 487.050 701.400 ;
        RECT 493.950 702.600 496.050 703.050 ;
        RECT 514.950 702.600 517.050 703.050 ;
        RECT 529.950 702.600 532.050 703.050 ;
        RECT 493.950 701.400 532.050 702.600 ;
        RECT 493.950 700.950 496.050 701.400 ;
        RECT 514.950 700.950 517.050 701.400 ;
        RECT 529.950 700.950 532.050 701.400 ;
        RECT 571.950 702.600 574.050 703.050 ;
        RECT 685.950 702.600 688.050 703.050 ;
        RECT 697.950 702.600 700.050 703.050 ;
        RECT 571.950 701.400 688.050 702.600 ;
        RECT 571.950 700.950 574.050 701.400 ;
        RECT 685.950 700.950 688.050 701.400 ;
        RECT 689.400 701.400 700.050 702.600 ;
        RECT 322.950 699.600 325.050 700.050 ;
        RECT 328.950 699.600 331.050 700.050 ;
        RECT 322.950 698.400 331.050 699.600 ;
        RECT 322.950 697.950 325.050 698.400 ;
        RECT 328.950 697.950 331.050 698.400 ;
        RECT 334.950 699.600 337.050 700.050 ;
        RECT 349.950 699.600 352.050 700.050 ;
        RECT 334.950 698.400 352.050 699.600 ;
        RECT 334.950 697.950 337.050 698.400 ;
        RECT 349.950 697.950 352.050 698.400 ;
        RECT 367.950 697.950 370.050 700.050 ;
        RECT 373.950 699.600 376.050 700.050 ;
        RECT 424.950 699.600 427.050 700.050 ;
        RECT 373.950 698.400 427.050 699.600 ;
        RECT 373.950 697.950 376.050 698.400 ;
        RECT 424.950 697.950 427.050 698.400 ;
        RECT 442.950 699.600 445.050 700.050 ;
        RECT 460.950 699.600 463.050 700.050 ;
        RECT 478.950 699.600 481.050 700.050 ;
        RECT 442.950 698.400 481.050 699.600 ;
        RECT 442.950 697.950 445.050 698.400 ;
        RECT 460.950 697.950 463.050 698.400 ;
        RECT 478.950 697.950 481.050 698.400 ;
        RECT 520.950 699.600 523.050 700.050 ;
        RECT 535.950 699.600 538.050 700.050 ;
        RECT 520.950 698.400 538.050 699.600 ;
        RECT 520.950 697.950 523.050 698.400 ;
        RECT 535.950 697.950 538.050 698.400 ;
        RECT 556.950 699.600 559.050 700.050 ;
        RECT 604.950 699.600 607.050 700.050 ;
        RECT 622.950 699.600 625.050 700.050 ;
        RECT 625.950 699.600 628.050 700.050 ;
        RECT 556.950 698.400 628.050 699.600 ;
        RECT 556.950 697.950 559.050 698.400 ;
        RECT 310.950 695.400 321.600 696.600 ;
        RECT 349.950 696.600 352.050 697.050 ;
        RECT 355.950 696.600 358.050 697.050 ;
        RECT 374.400 696.600 375.600 697.950 ;
        RECT 581.400 697.050 582.600 698.400 ;
        RECT 604.950 697.950 607.050 698.400 ;
        RECT 622.950 697.950 625.050 698.400 ;
        RECT 625.950 697.950 628.050 698.400 ;
        RECT 667.950 699.600 670.050 700.050 ;
        RECT 689.400 699.600 690.600 701.400 ;
        RECT 697.950 700.950 700.050 701.400 ;
        RECT 667.950 698.400 690.600 699.600 ;
        RECT 667.950 697.950 670.050 698.400 ;
        RECT 349.950 695.400 375.600 696.600 ;
        RECT 517.950 696.600 520.050 697.050 ;
        RECT 562.950 696.600 565.050 697.050 ;
        RECT 517.950 695.400 565.050 696.600 ;
        RECT 310.950 694.950 313.050 695.400 ;
        RECT 349.950 694.950 352.050 695.400 ;
        RECT 355.950 694.950 358.050 695.400 ;
        RECT 517.950 694.950 520.050 695.400 ;
        RECT 562.950 694.950 565.050 695.400 ;
        RECT 580.950 694.950 583.050 697.050 ;
        RECT 586.950 696.600 589.050 697.050 ;
        RECT 688.950 696.600 691.050 697.050 ;
        RECT 586.950 695.400 691.050 696.600 ;
        RECT 586.950 694.950 589.050 695.400 ;
        RECT 688.950 694.950 691.050 695.400 ;
        RECT 88.950 693.600 91.050 694.050 ;
        RECT 115.950 693.600 118.050 694.050 ;
        RECT 88.950 692.400 118.050 693.600 ;
        RECT 88.950 691.950 91.050 692.400 ;
        RECT 115.950 691.950 118.050 692.400 ;
        RECT 166.950 693.600 169.050 694.050 ;
        RECT 169.950 693.600 172.050 694.050 ;
        RECT 175.950 693.600 178.050 694.050 ;
        RECT 166.950 692.400 178.050 693.600 ;
        RECT 166.950 691.950 169.050 692.400 ;
        RECT 169.950 691.950 172.050 692.400 ;
        RECT 175.950 691.950 178.050 692.400 ;
        RECT 193.950 693.600 196.050 694.050 ;
        RECT 223.950 693.600 226.050 694.050 ;
        RECT 241.950 693.600 244.050 694.050 ;
        RECT 193.950 692.400 244.050 693.600 ;
        RECT 193.950 691.950 196.050 692.400 ;
        RECT 223.950 691.950 226.050 692.400 ;
        RECT 241.950 691.950 244.050 692.400 ;
        RECT 295.950 693.600 298.050 694.050 ;
        RECT 298.950 693.600 301.050 694.050 ;
        RECT 325.950 693.600 328.050 694.050 ;
        RECT 295.950 692.400 328.050 693.600 ;
        RECT 295.950 691.950 298.050 692.400 ;
        RECT 298.950 691.950 301.050 692.400 ;
        RECT 325.950 691.950 328.050 692.400 ;
        RECT 415.950 693.600 418.050 694.050 ;
        RECT 421.950 693.600 424.050 694.050 ;
        RECT 511.950 693.600 514.050 694.050 ;
        RECT 415.950 692.400 514.050 693.600 ;
        RECT 415.950 691.950 418.050 692.400 ;
        RECT 421.950 691.950 424.050 692.400 ;
        RECT 511.950 691.950 514.050 692.400 ;
        RECT 79.950 690.600 82.050 691.050 ;
        RECT 91.950 690.600 94.050 691.050 ;
        RECT 79.950 689.400 94.050 690.600 ;
        RECT 79.950 688.950 82.050 689.400 ;
        RECT 91.950 688.950 94.050 689.400 ;
        RECT 112.950 690.600 115.050 691.050 ;
        RECT 118.950 690.600 121.050 691.050 ;
        RECT 112.950 689.400 121.050 690.600 ;
        RECT 112.950 688.950 115.050 689.400 ;
        RECT 118.950 688.950 121.050 689.400 ;
        RECT 154.950 690.600 157.050 691.050 ;
        RECT 220.950 690.600 223.050 691.050 ;
        RECT 154.950 689.400 223.050 690.600 ;
        RECT 154.950 688.950 157.050 689.400 ;
        RECT 220.950 688.950 223.050 689.400 ;
        RECT 355.950 690.600 358.050 691.050 ;
        RECT 373.950 690.600 376.050 691.050 ;
        RECT 355.950 689.400 376.050 690.600 ;
        RECT 355.950 688.950 358.050 689.400 ;
        RECT 373.950 688.950 376.050 689.400 ;
        RECT 376.950 690.600 379.050 691.050 ;
        RECT 391.950 690.600 394.050 691.050 ;
        RECT 565.950 690.600 568.050 691.050 ;
        RECT 376.950 689.400 568.050 690.600 ;
        RECT 376.950 688.950 379.050 689.400 ;
        RECT 391.950 688.950 394.050 689.400 ;
        RECT 565.950 688.950 568.050 689.400 ;
        RECT 625.950 690.600 628.050 691.050 ;
        RECT 709.950 690.600 712.050 691.050 ;
        RECT 625.950 689.400 712.050 690.600 ;
        RECT 625.950 688.950 628.050 689.400 ;
        RECT 709.950 688.950 712.050 689.400 ;
        RECT 19.950 687.600 22.050 688.050 ;
        RECT 49.950 687.600 52.050 688.050 ;
        RECT 67.950 687.600 70.050 688.050 ;
        RECT 385.950 687.600 388.050 688.050 ;
        RECT 19.950 686.400 388.050 687.600 ;
        RECT 19.950 685.950 22.050 686.400 ;
        RECT 49.950 685.950 52.050 686.400 ;
        RECT 67.950 685.950 70.050 686.400 ;
        RECT 385.950 685.950 388.050 686.400 ;
        RECT 139.950 684.600 142.050 685.050 ;
        RECT 148.950 684.600 151.050 685.050 ;
        RECT 139.950 683.400 151.050 684.600 ;
        RECT 139.950 682.950 142.050 683.400 ;
        RECT 148.950 682.950 151.050 683.400 ;
        RECT 223.950 684.600 226.050 685.050 ;
        RECT 271.950 684.600 274.050 685.050 ;
        RECT 289.950 684.600 292.050 685.050 ;
        RECT 310.950 684.600 313.050 685.050 ;
        RECT 436.950 684.600 439.050 685.050 ;
        RECT 223.950 683.400 439.050 684.600 ;
        RECT 223.950 682.950 226.050 683.400 ;
        RECT 271.950 682.950 274.050 683.400 ;
        RECT 289.950 682.950 292.050 683.400 ;
        RECT 310.950 682.950 313.050 683.400 ;
        RECT 436.950 682.950 439.050 683.400 ;
        RECT 19.950 681.600 22.050 682.050 ;
        RECT 55.950 681.600 58.050 682.050 ;
        RECT 88.950 681.600 91.050 682.050 ;
        RECT 118.950 681.600 121.050 682.050 ;
        RECT 19.950 680.400 121.050 681.600 ;
        RECT 19.950 679.950 22.050 680.400 ;
        RECT 55.950 679.950 58.050 680.400 ;
        RECT 88.950 679.950 91.050 680.400 ;
        RECT 118.950 679.950 121.050 680.400 ;
        RECT 145.950 681.600 148.050 682.050 ;
        RECT 163.950 681.600 166.050 682.050 ;
        RECT 145.950 680.400 166.050 681.600 ;
        RECT 145.950 679.950 148.050 680.400 ;
        RECT 163.950 679.950 166.050 680.400 ;
        RECT 166.950 681.600 169.050 682.050 ;
        RECT 187.950 681.600 190.050 682.050 ;
        RECT 208.950 681.600 211.050 682.050 ;
        RECT 298.950 681.600 301.050 682.050 ;
        RECT 166.950 680.400 301.050 681.600 ;
        RECT 166.950 679.950 169.050 680.400 ;
        RECT 187.950 679.950 190.050 680.400 ;
        RECT 208.950 679.950 211.050 680.400 ;
        RECT 298.950 679.950 301.050 680.400 ;
        RECT 301.950 681.600 304.050 682.050 ;
        RECT 340.950 681.600 343.050 682.050 ;
        RECT 301.950 680.400 343.050 681.600 ;
        RECT 301.950 679.950 304.050 680.400 ;
        RECT 340.950 679.950 343.050 680.400 ;
        RECT 670.950 681.600 673.050 682.050 ;
        RECT 757.950 681.600 760.050 682.050 ;
        RECT 760.950 681.600 763.050 682.050 ;
        RECT 670.950 680.400 763.050 681.600 ;
        RECT 670.950 679.950 673.050 680.400 ;
        RECT 757.950 679.950 760.050 680.400 ;
        RECT 760.950 679.950 763.050 680.400 ;
        RECT 28.950 678.600 31.050 679.050 ;
        RECT 85.950 678.600 88.050 679.050 ;
        RECT 28.950 677.400 88.050 678.600 ;
        RECT 28.950 676.950 31.050 677.400 ;
        RECT 85.950 676.950 88.050 677.400 ;
        RECT 100.950 678.600 103.050 679.050 ;
        RECT 109.950 678.600 112.050 679.050 ;
        RECT 115.950 678.600 118.050 679.050 ;
        RECT 172.950 678.600 175.050 679.050 ;
        RECT 100.950 677.400 175.050 678.600 ;
        RECT 100.950 676.950 103.050 677.400 ;
        RECT 109.950 676.950 112.050 677.400 ;
        RECT 115.950 676.950 118.050 677.400 ;
        RECT 172.950 676.950 175.050 677.400 ;
        RECT 175.950 678.600 178.050 679.050 ;
        RECT 205.950 678.600 208.050 679.050 ;
        RECT 175.950 677.400 208.050 678.600 ;
        RECT 175.950 676.950 178.050 677.400 ;
        RECT 205.950 676.950 208.050 677.400 ;
        RECT 274.950 678.600 277.050 679.050 ;
        RECT 316.950 678.600 319.050 679.050 ;
        RECT 274.950 677.400 319.050 678.600 ;
        RECT 274.950 676.950 277.050 677.400 ;
        RECT 316.950 676.950 319.050 677.400 ;
        RECT 352.950 678.600 355.050 679.050 ;
        RECT 406.950 678.600 409.050 679.050 ;
        RECT 352.950 677.400 409.050 678.600 ;
        RECT 352.950 676.950 355.050 677.400 ;
        RECT 406.950 676.950 409.050 677.400 ;
        RECT 484.950 678.600 487.050 679.050 ;
        RECT 505.950 678.600 508.050 679.050 ;
        RECT 484.950 677.400 508.050 678.600 ;
        RECT 484.950 676.950 487.050 677.400 ;
        RECT 505.950 676.950 508.050 677.400 ;
        RECT 652.950 676.950 655.050 679.050 ;
        RECT 7.950 675.600 10.050 676.050 ;
        RECT 16.950 675.600 19.050 676.050 ;
        RECT 7.950 674.400 19.050 675.600 ;
        RECT 7.950 673.950 10.050 674.400 ;
        RECT 16.950 673.950 19.050 674.400 ;
        RECT 76.950 675.600 79.050 676.050 ;
        RECT 124.950 675.600 127.050 676.050 ;
        RECT 142.950 675.600 145.050 676.050 ;
        RECT 184.950 675.600 187.050 676.050 ;
        RECT 196.950 675.600 199.050 676.050 ;
        RECT 76.950 674.400 199.050 675.600 ;
        RECT 76.950 673.950 79.050 674.400 ;
        RECT 124.950 673.950 127.050 674.400 ;
        RECT 142.950 673.950 145.050 674.400 ;
        RECT 184.950 673.950 187.050 674.400 ;
        RECT 196.950 673.950 199.050 674.400 ;
        RECT 199.950 675.600 202.050 676.050 ;
        RECT 226.950 675.600 229.050 676.050 ;
        RECT 238.950 675.600 241.050 676.050 ;
        RECT 244.950 675.600 247.050 676.050 ;
        RECT 199.950 674.400 237.600 675.600 ;
        RECT 199.950 673.950 202.050 674.400 ;
        RECT 226.950 673.950 229.050 674.400 ;
        RECT 10.950 670.950 13.050 673.050 ;
        RECT 13.950 672.600 16.050 673.050 ;
        RECT 22.950 672.600 25.050 673.050 ;
        RECT 13.950 671.400 25.050 672.600 ;
        RECT 13.950 670.950 16.050 671.400 ;
        RECT 22.950 670.950 25.050 671.400 ;
        RECT 73.950 672.600 76.050 673.050 ;
        RECT 91.950 672.600 94.050 673.050 ;
        RECT 73.950 671.400 94.050 672.600 ;
        RECT 73.950 670.950 76.050 671.400 ;
        RECT 91.950 670.950 94.050 671.400 ;
        RECT 97.950 672.600 100.050 673.050 ;
        RECT 106.950 672.600 109.050 673.050 ;
        RECT 112.950 672.600 115.050 673.050 ;
        RECT 97.950 671.400 115.050 672.600 ;
        RECT 97.950 670.950 100.050 671.400 ;
        RECT 106.950 670.950 109.050 671.400 ;
        RECT 112.950 670.950 115.050 671.400 ;
        RECT 115.950 672.600 118.050 673.050 ;
        RECT 115.950 671.400 123.600 672.600 ;
        RECT 115.950 670.950 118.050 671.400 ;
        RECT 11.400 667.050 12.600 670.950 ;
        RECT 122.400 670.050 123.600 671.400 ;
        RECT 127.950 670.950 130.050 673.050 ;
        RECT 145.950 672.600 148.050 673.050 ;
        RECT 145.950 671.400 153.600 672.600 ;
        RECT 145.950 670.950 148.050 671.400 ;
        RECT 34.950 669.600 37.050 670.050 ;
        RECT 40.950 669.600 43.050 670.050 ;
        RECT 34.950 668.400 43.050 669.600 ;
        RECT 34.950 667.950 37.050 668.400 ;
        RECT 40.950 667.950 43.050 668.400 ;
        RECT 49.950 667.950 52.050 670.050 ;
        RECT 64.950 667.950 67.050 670.050 ;
        RECT 70.950 669.600 73.050 670.050 ;
        RECT 79.950 669.600 82.050 670.050 ;
        RECT 70.950 668.400 82.050 669.600 ;
        RECT 70.950 667.950 73.050 668.400 ;
        RECT 79.950 667.950 82.050 668.400 ;
        RECT 94.950 669.600 97.050 670.050 ;
        RECT 121.950 669.600 124.050 670.050 ;
        RECT 94.950 668.400 124.050 669.600 ;
        RECT 94.950 667.950 97.050 668.400 ;
        RECT 121.950 667.950 124.050 668.400 ;
        RECT 10.950 664.950 13.050 667.050 ;
        RECT 16.950 666.600 19.050 667.050 ;
        RECT 31.950 666.600 34.050 667.050 ;
        RECT 16.950 665.400 34.050 666.600 ;
        RECT 16.950 664.950 19.050 665.400 ;
        RECT 31.950 664.950 34.050 665.400 ;
        RECT 37.950 666.600 40.050 667.050 ;
        RECT 46.950 666.600 49.050 667.050 ;
        RECT 37.950 665.400 49.050 666.600 ;
        RECT 50.400 666.600 51.600 667.950 ;
        RECT 61.950 666.600 64.050 667.050 ;
        RECT 50.400 665.400 64.050 666.600 ;
        RECT 37.950 664.950 40.050 665.400 ;
        RECT 46.950 664.950 49.050 665.400 ;
        RECT 61.950 664.950 64.050 665.400 ;
        RECT 65.400 664.050 66.600 667.950 ;
        RECT 128.400 667.050 129.600 670.950 ;
        RECT 152.400 670.050 153.600 671.400 ;
        RECT 160.950 670.950 163.050 673.050 ;
        RECT 172.950 672.600 175.050 673.050 ;
        RECT 178.950 672.600 181.050 673.050 ;
        RECT 190.950 672.600 193.050 673.050 ;
        RECT 199.950 672.600 202.050 673.050 ;
        RECT 172.950 671.400 193.050 672.600 ;
        RECT 172.950 670.950 175.050 671.400 ;
        RECT 178.950 670.950 181.050 671.400 ;
        RECT 190.950 670.950 193.050 671.400 ;
        RECT 194.400 671.400 202.050 672.600 ;
        RECT 130.950 669.600 133.050 670.050 ;
        RECT 136.950 669.600 139.050 670.050 ;
        RECT 130.950 668.400 139.050 669.600 ;
        RECT 130.950 667.950 133.050 668.400 ;
        RECT 136.950 667.950 139.050 668.400 ;
        RECT 145.950 667.950 148.050 670.050 ;
        RECT 151.950 667.950 154.050 670.050 ;
        RECT 161.400 669.600 162.600 670.950 ;
        RECT 175.950 669.600 178.050 670.050 ;
        RECT 194.400 669.600 195.600 671.400 ;
        RECT 199.950 670.950 202.050 671.400 ;
        RECT 211.950 672.600 214.050 673.050 ;
        RECT 232.950 672.600 235.050 673.050 ;
        RECT 211.950 671.400 235.050 672.600 ;
        RECT 236.400 672.600 237.600 674.400 ;
        RECT 238.950 674.400 247.050 675.600 ;
        RECT 238.950 673.950 241.050 674.400 ;
        RECT 244.950 673.950 247.050 674.400 ;
        RECT 253.950 675.600 256.050 676.050 ;
        RECT 262.950 675.600 265.050 676.050 ;
        RECT 253.950 674.400 265.050 675.600 ;
        RECT 253.950 673.950 256.050 674.400 ;
        RECT 262.950 673.950 265.050 674.400 ;
        RECT 319.950 675.600 322.050 676.050 ;
        RECT 346.950 675.600 349.050 676.050 ;
        RECT 373.950 675.600 376.050 676.050 ;
        RECT 382.950 675.600 385.050 676.050 ;
        RECT 319.950 674.400 349.050 675.600 ;
        RECT 319.950 673.950 322.050 674.400 ;
        RECT 346.950 673.950 349.050 674.400 ;
        RECT 359.400 674.400 385.050 675.600 ;
        RECT 283.950 672.600 286.050 673.050 ;
        RECT 236.400 671.400 286.050 672.600 ;
        RECT 211.950 670.950 214.050 671.400 ;
        RECT 232.950 670.950 235.050 671.400 ;
        RECT 283.950 670.950 286.050 671.400 ;
        RECT 289.950 672.600 292.050 673.050 ;
        RECT 301.950 672.600 304.050 673.050 ;
        RECT 289.950 671.400 304.050 672.600 ;
        RECT 289.950 670.950 292.050 671.400 ;
        RECT 301.950 670.950 304.050 671.400 ;
        RECT 310.950 672.600 313.050 673.050 ;
        RECT 331.950 672.600 334.050 673.050 ;
        RECT 352.950 672.600 355.050 673.050 ;
        RECT 310.950 671.400 334.050 672.600 ;
        RECT 310.950 670.950 313.050 671.400 ;
        RECT 331.950 670.950 334.050 671.400 ;
        RECT 344.400 671.400 355.050 672.600 ;
        RECT 344.400 670.050 345.600 671.400 ;
        RECT 352.950 670.950 355.050 671.400 ;
        RECT 359.400 670.050 360.600 674.400 ;
        RECT 373.950 673.950 376.050 674.400 ;
        RECT 382.950 673.950 385.050 674.400 ;
        RECT 430.950 675.600 433.050 676.050 ;
        RECT 451.950 675.600 454.050 676.050 ;
        RECT 430.950 674.400 454.050 675.600 ;
        RECT 430.950 673.950 433.050 674.400 ;
        RECT 451.950 673.950 454.050 674.400 ;
        RECT 361.950 670.950 364.050 673.050 ;
        RECT 499.950 672.600 502.050 673.050 ;
        RECT 488.400 671.400 502.050 672.600 ;
        RECT 161.400 668.400 195.600 669.600 ;
        RECT 205.950 669.600 208.050 670.050 ;
        RECT 214.950 669.600 217.050 670.050 ;
        RECT 235.950 669.600 238.050 670.050 ;
        RECT 256.950 669.600 259.050 670.050 ;
        RECT 205.950 668.400 234.600 669.600 ;
        RECT 175.950 667.950 178.050 668.400 ;
        RECT 205.950 667.950 208.050 668.400 ;
        RECT 214.950 667.950 217.050 668.400 ;
        RECT 85.950 666.600 88.050 667.050 ;
        RECT 109.950 666.600 112.050 667.050 ;
        RECT 85.950 665.400 112.050 666.600 ;
        RECT 85.950 664.950 88.050 665.400 ;
        RECT 109.950 664.950 112.050 665.400 ;
        RECT 127.950 664.950 130.050 667.050 ;
        RECT 133.950 666.600 136.050 667.050 ;
        RECT 139.950 666.600 142.050 667.050 ;
        RECT 133.950 665.400 142.050 666.600 ;
        RECT 146.400 666.600 147.600 667.950 ;
        RECT 172.950 666.600 175.050 667.050 ;
        RECT 146.400 665.400 175.050 666.600 ;
        RECT 133.950 664.950 136.050 665.400 ;
        RECT 139.950 664.950 142.050 665.400 ;
        RECT 172.950 664.950 175.050 665.400 ;
        RECT 181.950 666.600 184.050 667.050 ;
        RECT 187.950 666.600 190.050 667.050 ;
        RECT 196.950 666.600 199.050 667.050 ;
        RECT 181.950 665.400 199.050 666.600 ;
        RECT 181.950 664.950 184.050 665.400 ;
        RECT 187.950 664.950 190.050 665.400 ;
        RECT 196.950 664.950 199.050 665.400 ;
        RECT 202.950 666.600 205.050 667.050 ;
        RECT 220.950 666.600 223.050 667.050 ;
        RECT 202.950 665.400 223.050 666.600 ;
        RECT 233.400 666.600 234.600 668.400 ;
        RECT 235.950 668.400 259.050 669.600 ;
        RECT 235.950 667.950 238.050 668.400 ;
        RECT 256.950 667.950 259.050 668.400 ;
        RECT 259.950 669.600 262.050 670.050 ;
        RECT 268.950 669.600 271.050 670.050 ;
        RECT 280.950 669.600 283.050 670.050 ;
        RECT 259.950 668.400 283.050 669.600 ;
        RECT 259.950 667.950 262.050 668.400 ;
        RECT 268.950 667.950 271.050 668.400 ;
        RECT 280.950 667.950 283.050 668.400 ;
        RECT 286.950 669.600 289.050 670.050 ;
        RECT 295.950 669.600 298.050 670.050 ;
        RECT 286.950 668.400 298.050 669.600 ;
        RECT 286.950 667.950 289.050 668.400 ;
        RECT 295.950 667.950 298.050 668.400 ;
        RECT 325.950 669.600 328.050 670.050 ;
        RECT 337.950 669.600 340.050 670.050 ;
        RECT 325.950 668.400 340.050 669.600 ;
        RECT 325.950 667.950 328.050 668.400 ;
        RECT 337.950 667.950 340.050 668.400 ;
        RECT 343.950 667.950 346.050 670.050 ;
        RECT 352.950 669.600 355.050 670.050 ;
        RECT 347.400 668.400 355.050 669.600 ;
        RECT 347.400 667.050 348.600 668.400 ;
        RECT 352.950 667.950 355.050 668.400 ;
        RECT 358.950 667.950 361.050 670.050 ;
        RECT 256.950 666.600 259.050 667.050 ;
        RECT 233.400 665.400 259.050 666.600 ;
        RECT 202.950 664.950 205.050 665.400 ;
        RECT 220.950 664.950 223.050 665.400 ;
        RECT 256.950 664.950 259.050 665.400 ;
        RECT 298.950 666.600 301.050 667.050 ;
        RECT 313.950 666.600 316.050 667.050 ;
        RECT 298.950 665.400 316.050 666.600 ;
        RECT 298.950 664.950 301.050 665.400 ;
        RECT 313.950 664.950 316.050 665.400 ;
        RECT 319.950 666.600 322.050 667.050 ;
        RECT 328.950 666.600 331.050 667.050 ;
        RECT 319.950 665.400 331.050 666.600 ;
        RECT 319.950 664.950 322.050 665.400 ;
        RECT 328.950 664.950 331.050 665.400 ;
        RECT 331.950 666.600 334.050 667.050 ;
        RECT 343.950 666.600 346.050 667.050 ;
        RECT 331.950 665.400 346.050 666.600 ;
        RECT 331.950 664.950 334.050 665.400 ;
        RECT 343.950 664.950 346.050 665.400 ;
        RECT 346.950 664.950 349.050 667.050 ;
        RECT 362.400 666.600 363.600 670.950 ;
        RECT 388.950 669.600 391.050 670.050 ;
        RECT 394.950 669.600 397.050 670.050 ;
        RECT 388.950 668.400 397.050 669.600 ;
        RECT 388.950 667.950 391.050 668.400 ;
        RECT 394.950 667.950 397.050 668.400 ;
        RECT 418.950 669.600 421.050 670.050 ;
        RECT 463.950 669.600 466.050 670.050 ;
        RECT 488.400 669.600 489.600 671.400 ;
        RECT 499.950 670.950 502.050 671.400 ;
        RECT 541.950 672.600 544.050 673.050 ;
        RECT 574.950 672.600 577.050 673.050 ;
        RECT 541.950 671.400 577.050 672.600 ;
        RECT 541.950 670.950 544.050 671.400 ;
        RECT 574.950 670.950 577.050 671.400 ;
        RECT 653.400 670.050 654.600 676.950 ;
        RECT 721.950 675.600 724.050 676.050 ;
        RECT 707.400 674.400 724.050 675.600 ;
        RECT 703.950 672.600 706.050 673.050 ;
        RECT 692.400 671.400 706.050 672.600 ;
        RECT 418.950 668.400 489.600 669.600 ;
        RECT 493.950 669.600 496.050 670.050 ;
        RECT 502.950 669.600 505.050 670.050 ;
        RECT 493.950 668.400 505.050 669.600 ;
        RECT 418.950 667.950 421.050 668.400 ;
        RECT 463.950 667.950 466.050 668.400 ;
        RECT 493.950 667.950 496.050 668.400 ;
        RECT 502.950 667.950 505.050 668.400 ;
        RECT 508.950 669.600 511.050 670.050 ;
        RECT 517.950 669.600 520.050 670.050 ;
        RECT 508.950 668.400 520.050 669.600 ;
        RECT 508.950 667.950 511.050 668.400 ;
        RECT 517.950 667.950 520.050 668.400 ;
        RECT 544.950 669.600 547.050 670.050 ;
        RECT 556.950 669.600 559.050 670.050 ;
        RECT 544.950 668.400 559.050 669.600 ;
        RECT 544.950 667.950 547.050 668.400 ;
        RECT 556.950 667.950 559.050 668.400 ;
        RECT 604.950 667.950 607.050 670.050 ;
        RECT 625.950 669.600 628.050 670.050 ;
        RECT 631.950 669.600 634.050 670.050 ;
        RECT 625.950 668.400 634.050 669.600 ;
        RECT 625.950 667.950 628.050 668.400 ;
        RECT 631.950 667.950 634.050 668.400 ;
        RECT 652.950 667.950 655.050 670.050 ;
        RECT 655.950 669.600 658.050 670.050 ;
        RECT 688.950 669.600 691.050 670.050 ;
        RECT 655.950 668.400 691.050 669.600 ;
        RECT 655.950 667.950 658.050 668.400 ;
        RECT 688.950 667.950 691.050 668.400 ;
        RECT 364.950 666.600 367.050 667.050 ;
        RECT 362.400 665.400 367.050 666.600 ;
        RECT 364.950 664.950 367.050 665.400 ;
        RECT 427.950 666.600 430.050 667.050 ;
        RECT 457.950 666.600 460.050 667.050 ;
        RECT 427.950 665.400 460.050 666.600 ;
        RECT 427.950 664.950 430.050 665.400 ;
        RECT 457.950 664.950 460.050 665.400 ;
        RECT 520.950 666.600 523.050 667.050 ;
        RECT 538.950 666.600 541.050 667.050 ;
        RECT 553.950 666.600 556.050 667.050 ;
        RECT 520.950 665.400 556.050 666.600 ;
        RECT 520.950 664.950 523.050 665.400 ;
        RECT 538.950 664.950 541.050 665.400 ;
        RECT 553.950 664.950 556.050 665.400 ;
        RECT 559.950 666.600 562.050 667.050 ;
        RECT 592.950 666.600 595.050 667.050 ;
        RECT 559.950 665.400 595.050 666.600 ;
        RECT 559.950 664.950 562.050 665.400 ;
        RECT 592.950 664.950 595.050 665.400 ;
        RECT 605.400 664.050 606.600 667.950 ;
        RECT 692.400 667.050 693.600 671.400 ;
        RECT 703.950 670.950 706.050 671.400 ;
        RECT 707.400 670.050 708.600 674.400 ;
        RECT 721.950 673.950 724.050 674.400 ;
        RECT 709.950 670.950 712.050 673.050 ;
        RECT 736.950 672.600 739.050 673.050 ;
        RECT 751.950 672.600 754.050 673.050 ;
        RECT 736.950 671.400 754.050 672.600 ;
        RECT 736.950 670.950 739.050 671.400 ;
        RECT 751.950 670.950 754.050 671.400 ;
        RECT 706.950 667.950 709.050 670.050 ;
        RECT 710.400 667.050 711.600 670.950 ;
        RECT 721.950 669.600 724.050 670.050 ;
        RECT 733.950 669.600 736.050 670.050 ;
        RECT 721.950 668.400 736.050 669.600 ;
        RECT 721.950 667.950 724.050 668.400 ;
        RECT 733.950 667.950 736.050 668.400 ;
        RECT 739.950 669.600 742.050 670.050 ;
        RECT 766.950 669.600 769.050 670.050 ;
        RECT 739.950 668.400 769.050 669.600 ;
        RECT 739.950 667.950 742.050 668.400 ;
        RECT 766.950 667.950 769.050 668.400 ;
        RECT 691.950 664.950 694.050 667.050 ;
        RECT 709.950 666.600 712.050 667.050 ;
        RECT 727.950 666.600 730.050 667.050 ;
        RECT 709.950 665.400 730.050 666.600 ;
        RECT 709.950 664.950 712.050 665.400 ;
        RECT 727.950 664.950 730.050 665.400 ;
        RECT 736.950 666.600 739.050 667.050 ;
        RECT 742.950 666.600 745.050 667.050 ;
        RECT 736.950 665.400 745.050 666.600 ;
        RECT 736.950 664.950 739.050 665.400 ;
        RECT 742.950 664.950 745.050 665.400 ;
        RECT 4.950 663.600 7.050 664.050 ;
        RECT 7.950 663.600 10.050 664.050 ;
        RECT 13.950 663.600 16.050 664.050 ;
        RECT 4.950 662.400 16.050 663.600 ;
        RECT 4.950 661.950 7.050 662.400 ;
        RECT 7.950 661.950 10.050 662.400 ;
        RECT 13.950 661.950 16.050 662.400 ;
        RECT 64.950 661.950 67.050 664.050 ;
        RECT 112.950 663.600 115.050 664.050 ;
        RECT 232.950 663.600 235.050 664.050 ;
        RECT 112.950 662.400 235.050 663.600 ;
        RECT 112.950 661.950 115.050 662.400 ;
        RECT 232.950 661.950 235.050 662.400 ;
        RECT 271.950 663.600 274.050 664.050 ;
        RECT 286.950 663.600 289.050 664.050 ;
        RECT 271.950 662.400 289.050 663.600 ;
        RECT 271.950 661.950 274.050 662.400 ;
        RECT 286.950 661.950 289.050 662.400 ;
        RECT 397.950 663.600 400.050 664.050 ;
        RECT 466.950 663.600 469.050 664.050 ;
        RECT 514.950 663.600 517.050 664.050 ;
        RECT 397.950 662.400 517.050 663.600 ;
        RECT 397.950 661.950 400.050 662.400 ;
        RECT 466.950 661.950 469.050 662.400 ;
        RECT 514.950 661.950 517.050 662.400 ;
        RECT 604.950 661.950 607.050 664.050 ;
        RECT 694.950 663.600 697.050 664.050 ;
        RECT 718.950 663.600 721.050 664.050 ;
        RECT 694.950 662.400 721.050 663.600 ;
        RECT 694.950 661.950 697.050 662.400 ;
        RECT 718.950 661.950 721.050 662.400 ;
        RECT 61.950 660.600 64.050 661.050 ;
        RECT 136.950 660.600 139.050 661.050 ;
        RECT 61.950 659.400 139.050 660.600 ;
        RECT 61.950 658.950 64.050 659.400 ;
        RECT 136.950 658.950 139.050 659.400 ;
        RECT 208.950 660.600 211.050 661.050 ;
        RECT 229.950 660.600 232.050 661.050 ;
        RECT 208.950 659.400 232.050 660.600 ;
        RECT 208.950 658.950 211.050 659.400 ;
        RECT 229.950 658.950 232.050 659.400 ;
        RECT 244.950 660.600 247.050 661.050 ;
        RECT 250.950 660.600 253.050 661.050 ;
        RECT 244.950 659.400 253.050 660.600 ;
        RECT 244.950 658.950 247.050 659.400 ;
        RECT 250.950 658.950 253.050 659.400 ;
        RECT 262.950 660.600 265.050 661.050 ;
        RECT 307.950 660.600 310.050 661.050 ;
        RECT 346.950 660.600 349.050 661.050 ;
        RECT 262.950 659.400 310.050 660.600 ;
        RECT 262.950 658.950 265.050 659.400 ;
        RECT 307.950 658.950 310.050 659.400 ;
        RECT 326.400 659.400 349.050 660.600 ;
        RECT 25.950 657.600 28.050 658.050 ;
        RECT 82.950 657.600 85.050 658.050 ;
        RECT 211.950 657.600 214.050 658.050 ;
        RECT 25.950 656.400 214.050 657.600 ;
        RECT 25.950 655.950 28.050 656.400 ;
        RECT 82.950 655.950 85.050 656.400 ;
        RECT 211.950 655.950 214.050 656.400 ;
        RECT 217.950 657.600 220.050 658.050 ;
        RECT 274.950 657.600 277.050 658.050 ;
        RECT 292.950 657.600 295.050 658.050 ;
        RECT 326.400 657.600 327.600 659.400 ;
        RECT 346.950 658.950 349.050 659.400 ;
        RECT 433.950 660.600 436.050 661.050 ;
        RECT 475.950 660.600 478.050 661.050 ;
        RECT 433.950 659.400 478.050 660.600 ;
        RECT 433.950 658.950 436.050 659.400 ;
        RECT 475.950 658.950 478.050 659.400 ;
        RECT 508.950 660.600 511.050 661.050 ;
        RECT 523.950 660.600 526.050 661.050 ;
        RECT 508.950 659.400 526.050 660.600 ;
        RECT 508.950 658.950 511.050 659.400 ;
        RECT 523.950 658.950 526.050 659.400 ;
        RECT 670.950 660.600 673.050 661.050 ;
        RECT 715.950 660.600 718.050 661.050 ;
        RECT 670.950 659.400 718.050 660.600 ;
        RECT 670.950 658.950 673.050 659.400 ;
        RECT 715.950 658.950 718.050 659.400 ;
        RECT 217.950 656.400 327.600 657.600 ;
        RECT 328.950 657.600 331.050 658.050 ;
        RECT 382.950 657.600 385.050 658.050 ;
        RECT 328.950 656.400 385.050 657.600 ;
        RECT 217.950 655.950 220.050 656.400 ;
        RECT 274.950 655.950 277.050 656.400 ;
        RECT 292.950 655.950 295.050 656.400 ;
        RECT 328.950 655.950 331.050 656.400 ;
        RECT 382.950 655.950 385.050 656.400 ;
        RECT 439.950 657.600 442.050 658.050 ;
        RECT 592.950 657.600 595.050 658.050 ;
        RECT 439.950 656.400 595.050 657.600 ;
        RECT 439.950 655.950 442.050 656.400 ;
        RECT 592.950 655.950 595.050 656.400 ;
        RECT 607.950 657.600 610.050 658.050 ;
        RECT 640.950 657.600 643.050 658.050 ;
        RECT 607.950 656.400 643.050 657.600 ;
        RECT 607.950 655.950 610.050 656.400 ;
        RECT 640.950 655.950 643.050 656.400 ;
        RECT 169.950 654.600 172.050 655.050 ;
        RECT 262.950 654.600 265.050 655.050 ;
        RECT 169.950 653.400 265.050 654.600 ;
        RECT 169.950 652.950 172.050 653.400 ;
        RECT 262.950 652.950 265.050 653.400 ;
        RECT 268.950 654.600 271.050 655.050 ;
        RECT 304.950 654.600 307.050 655.050 ;
        RECT 721.950 654.600 724.050 655.050 ;
        RECT 268.950 653.400 307.050 654.600 ;
        RECT 268.950 652.950 271.050 653.400 ;
        RECT 304.950 652.950 307.050 653.400 ;
        RECT 656.400 653.400 724.050 654.600 ;
        RECT 436.950 651.600 439.050 652.050 ;
        RECT 656.400 651.600 657.600 653.400 ;
        RECT 721.950 652.950 724.050 653.400 ;
        RECT 436.950 650.400 657.600 651.600 ;
        RECT 658.950 651.600 661.050 652.050 ;
        RECT 730.950 651.600 733.050 652.050 ;
        RECT 658.950 650.400 733.050 651.600 ;
        RECT 436.950 649.950 439.050 650.400 ;
        RECT 658.950 649.950 661.050 650.400 ;
        RECT 730.950 649.950 733.050 650.400 ;
        RECT 322.950 648.600 325.050 649.050 ;
        RECT 397.950 648.600 400.050 649.050 ;
        RECT 322.950 647.400 400.050 648.600 ;
        RECT 322.950 646.950 325.050 647.400 ;
        RECT 397.950 646.950 400.050 647.400 ;
        RECT 406.950 648.600 409.050 649.050 ;
        RECT 559.950 648.600 562.050 649.050 ;
        RECT 634.950 648.600 637.050 649.050 ;
        RECT 406.950 647.400 637.050 648.600 ;
        RECT 406.950 646.950 409.050 647.400 ;
        RECT 559.950 646.950 562.050 647.400 ;
        RECT 634.950 646.950 637.050 647.400 ;
        RECT 682.950 648.600 685.050 649.050 ;
        RECT 736.950 648.600 739.050 649.050 ;
        RECT 682.950 647.400 739.050 648.600 ;
        RECT 682.950 646.950 685.050 647.400 ;
        RECT 736.950 646.950 739.050 647.400 ;
        RECT 235.950 645.600 238.050 646.050 ;
        RECT 241.950 645.600 244.050 646.050 ;
        RECT 235.950 644.400 244.050 645.600 ;
        RECT 235.950 643.950 238.050 644.400 ;
        RECT 241.950 643.950 244.050 644.400 ;
        RECT 676.950 645.600 679.050 646.050 ;
        RECT 685.950 645.600 688.050 646.050 ;
        RECT 676.950 644.400 688.050 645.600 ;
        RECT 676.950 643.950 679.050 644.400 ;
        RECT 685.950 643.950 688.050 644.400 ;
        RECT 715.950 645.600 718.050 646.050 ;
        RECT 748.950 645.600 751.050 646.050 ;
        RECT 715.950 644.400 751.050 645.600 ;
        RECT 715.950 643.950 718.050 644.400 ;
        RECT 748.950 643.950 751.050 644.400 ;
        RECT 169.950 642.600 172.050 643.050 ;
        RECT 361.950 642.600 364.050 643.050 ;
        RECT 169.950 641.400 364.050 642.600 ;
        RECT 169.950 640.950 172.050 641.400 ;
        RECT 361.950 640.950 364.050 641.400 ;
        RECT 364.950 642.600 367.050 643.050 ;
        RECT 517.950 642.600 520.050 643.050 ;
        RECT 364.950 641.400 520.050 642.600 ;
        RECT 364.950 640.950 367.050 641.400 ;
        RECT 517.950 640.950 520.050 641.400 ;
        RECT 556.950 642.600 559.050 643.050 ;
        RECT 742.950 642.600 745.050 643.050 ;
        RECT 556.950 641.400 745.050 642.600 ;
        RECT 556.950 640.950 559.050 641.400 ;
        RECT 742.950 640.950 745.050 641.400 ;
        RECT 37.950 639.600 40.050 640.050 ;
        RECT 58.950 639.600 61.050 640.050 ;
        RECT 37.950 638.400 61.050 639.600 ;
        RECT 37.950 637.950 40.050 638.400 ;
        RECT 58.950 637.950 61.050 638.400 ;
        RECT 82.950 639.600 85.050 640.050 ;
        RECT 139.950 639.600 142.050 640.050 ;
        RECT 202.950 639.600 205.050 640.050 ;
        RECT 82.950 638.400 205.050 639.600 ;
        RECT 82.950 637.950 85.050 638.400 ;
        RECT 139.950 637.950 142.050 638.400 ;
        RECT 202.950 637.950 205.050 638.400 ;
        RECT 205.950 639.600 208.050 640.050 ;
        RECT 229.950 639.600 232.050 640.050 ;
        RECT 268.950 639.600 271.050 640.050 ;
        RECT 205.950 638.400 271.050 639.600 ;
        RECT 205.950 637.950 208.050 638.400 ;
        RECT 229.950 637.950 232.050 638.400 ;
        RECT 268.950 637.950 271.050 638.400 ;
        RECT 457.950 639.600 460.050 640.050 ;
        RECT 487.950 639.600 490.050 640.050 ;
        RECT 457.950 638.400 490.050 639.600 ;
        RECT 457.950 637.950 460.050 638.400 ;
        RECT 487.950 637.950 490.050 638.400 ;
        RECT 700.950 639.600 703.050 640.050 ;
        RECT 724.950 639.600 727.050 640.050 ;
        RECT 700.950 638.400 727.050 639.600 ;
        RECT 700.950 637.950 703.050 638.400 ;
        RECT 724.950 637.950 727.050 638.400 ;
        RECT 40.950 636.600 43.050 637.050 ;
        RECT 106.950 636.600 109.050 637.050 ;
        RECT 40.950 635.400 109.050 636.600 ;
        RECT 40.950 634.950 43.050 635.400 ;
        RECT 106.950 634.950 109.050 635.400 ;
        RECT 121.950 636.600 124.050 637.050 ;
        RECT 142.950 636.600 145.050 637.050 ;
        RECT 121.950 635.400 145.050 636.600 ;
        RECT 121.950 634.950 124.050 635.400 ;
        RECT 142.950 634.950 145.050 635.400 ;
        RECT 172.950 636.600 175.050 637.050 ;
        RECT 181.950 636.600 184.050 637.050 ;
        RECT 172.950 635.400 184.050 636.600 ;
        RECT 172.950 634.950 175.050 635.400 ;
        RECT 181.950 634.950 184.050 635.400 ;
        RECT 211.950 636.600 214.050 637.050 ;
        RECT 223.950 636.600 226.050 637.050 ;
        RECT 211.950 635.400 226.050 636.600 ;
        RECT 211.950 634.950 214.050 635.400 ;
        RECT 223.950 634.950 226.050 635.400 ;
        RECT 253.950 636.600 256.050 637.050 ;
        RECT 274.950 636.600 277.050 637.050 ;
        RECT 253.950 635.400 277.050 636.600 ;
        RECT 253.950 634.950 256.050 635.400 ;
        RECT 274.950 634.950 277.050 635.400 ;
        RECT 289.950 636.600 292.050 637.050 ;
        RECT 325.950 636.600 328.050 637.050 ;
        RECT 289.950 635.400 328.050 636.600 ;
        RECT 289.950 634.950 292.050 635.400 ;
        RECT 325.950 634.950 328.050 635.400 ;
        RECT 361.950 636.600 364.050 637.050 ;
        RECT 415.950 636.600 418.050 637.050 ;
        RECT 466.950 636.600 469.050 637.050 ;
        RECT 361.950 635.400 469.050 636.600 ;
        RECT 361.950 634.950 364.050 635.400 ;
        RECT 415.950 634.950 418.050 635.400 ;
        RECT 466.950 634.950 469.050 635.400 ;
        RECT 511.950 636.600 514.050 637.050 ;
        RECT 538.950 636.600 541.050 637.050 ;
        RECT 511.950 635.400 541.050 636.600 ;
        RECT 511.950 634.950 514.050 635.400 ;
        RECT 538.950 634.950 541.050 635.400 ;
        RECT 598.950 636.600 601.050 637.050 ;
        RECT 691.950 636.600 694.050 637.050 ;
        RECT 598.950 635.400 694.050 636.600 ;
        RECT 598.950 634.950 601.050 635.400 ;
        RECT 691.950 634.950 694.050 635.400 ;
        RECT 724.950 636.600 727.050 637.050 ;
        RECT 769.950 636.600 772.050 637.050 ;
        RECT 724.950 635.400 772.050 636.600 ;
        RECT 724.950 634.950 727.050 635.400 ;
        RECT 769.950 634.950 772.050 635.400 ;
        RECT 10.950 633.600 13.050 634.050 ;
        RECT 16.950 633.600 19.050 634.050 ;
        RECT 19.950 633.600 22.050 634.050 ;
        RECT 10.950 632.400 22.050 633.600 ;
        RECT 10.950 631.950 13.050 632.400 ;
        RECT 16.950 631.950 19.050 632.400 ;
        RECT 19.950 631.950 22.050 632.400 ;
        RECT 37.950 633.600 40.050 634.050 ;
        RECT 43.950 633.600 46.050 634.050 ;
        RECT 55.950 633.600 58.050 634.050 ;
        RECT 91.950 633.600 94.050 634.050 ;
        RECT 37.950 632.400 42.600 633.600 ;
        RECT 37.950 631.950 40.050 632.400 ;
        RECT 41.400 631.050 42.600 632.400 ;
        RECT 43.950 632.400 94.050 633.600 ;
        RECT 43.950 631.950 46.050 632.400 ;
        RECT 55.950 631.950 58.050 632.400 ;
        RECT 91.950 631.950 94.050 632.400 ;
        RECT 133.950 633.600 136.050 634.050 ;
        RECT 154.950 633.600 157.050 634.050 ;
        RECT 217.950 633.600 220.050 634.050 ;
        RECT 133.950 632.400 157.050 633.600 ;
        RECT 133.950 631.950 136.050 632.400 ;
        RECT 154.950 631.950 157.050 632.400 ;
        RECT 173.400 632.400 220.050 633.600 ;
        RECT 173.400 631.050 174.600 632.400 ;
        RECT 217.950 631.950 220.050 632.400 ;
        RECT 229.950 633.600 232.050 634.050 ;
        RECT 325.950 633.600 328.050 634.050 ;
        RECT 346.950 633.600 349.050 634.050 ;
        RECT 229.950 632.400 237.600 633.600 ;
        RECT 229.950 631.950 232.050 632.400 ;
        RECT 7.950 630.600 10.050 631.050 ;
        RECT 5.400 629.400 10.050 630.600 ;
        RECT 5.400 628.050 6.600 629.400 ;
        RECT 7.950 628.950 10.050 629.400 ;
        RECT 40.950 628.950 43.050 631.050 ;
        RECT 43.950 630.600 46.050 631.050 ;
        RECT 61.950 630.600 64.050 631.050 ;
        RECT 67.950 630.600 70.050 631.050 ;
        RECT 79.950 630.600 82.050 631.050 ;
        RECT 85.950 630.600 88.050 631.050 ;
        RECT 43.950 629.400 66.600 630.600 ;
        RECT 43.950 628.950 46.050 629.400 ;
        RECT 61.950 628.950 64.050 629.400 ;
        RECT 4.950 627.600 7.050 628.050 ;
        RECT 13.950 627.600 16.050 628.050 ;
        RECT 4.950 626.400 16.050 627.600 ;
        RECT 4.950 625.950 7.050 626.400 ;
        RECT 13.950 625.950 16.050 626.400 ;
        RECT 28.950 627.600 31.050 628.050 ;
        RECT 46.950 627.600 49.050 628.050 ;
        RECT 28.950 626.400 49.050 627.600 ;
        RECT 65.400 627.600 66.600 629.400 ;
        RECT 67.950 629.400 75.600 630.600 ;
        RECT 67.950 628.950 70.050 629.400 ;
        RECT 65.400 626.400 72.600 627.600 ;
        RECT 28.950 625.950 31.050 626.400 ;
        RECT 46.950 625.950 49.050 626.400 ;
        RECT 71.400 625.050 72.600 626.400 ;
        RECT 10.950 624.600 13.050 625.050 ;
        RECT 16.950 624.600 19.050 625.050 ;
        RECT 10.950 623.400 19.050 624.600 ;
        RECT 10.950 622.950 13.050 623.400 ;
        RECT 16.950 622.950 19.050 623.400 ;
        RECT 70.950 622.950 73.050 625.050 ;
        RECT 34.950 621.600 37.050 622.050 ;
        RECT 74.400 621.600 75.600 629.400 ;
        RECT 79.950 629.400 88.050 630.600 ;
        RECT 79.950 628.950 82.050 629.400 ;
        RECT 85.950 628.950 88.050 629.400 ;
        RECT 100.950 630.600 103.050 631.050 ;
        RECT 115.950 630.600 118.050 631.050 ;
        RECT 100.950 629.400 118.050 630.600 ;
        RECT 100.950 628.950 103.050 629.400 ;
        RECT 115.950 628.950 118.050 629.400 ;
        RECT 136.950 630.600 139.050 631.050 ;
        RECT 148.950 630.600 151.050 631.050 ;
        RECT 136.950 629.400 151.050 630.600 ;
        RECT 136.950 628.950 139.050 629.400 ;
        RECT 148.950 628.950 151.050 629.400 ;
        RECT 163.950 628.950 166.050 631.050 ;
        RECT 172.950 628.950 175.050 631.050 ;
        RECT 178.950 630.600 181.050 631.050 ;
        RECT 196.950 630.600 199.050 631.050 ;
        RECT 178.950 629.400 199.050 630.600 ;
        RECT 178.950 628.950 181.050 629.400 ;
        RECT 196.950 628.950 199.050 629.400 ;
        RECT 199.950 630.600 202.050 631.050 ;
        RECT 211.950 630.600 214.050 631.050 ;
        RECT 199.950 629.400 214.050 630.600 ;
        RECT 199.950 628.950 202.050 629.400 ;
        RECT 211.950 628.950 214.050 629.400 ;
        RECT 91.950 627.600 94.050 628.050 ;
        RECT 97.950 627.600 100.050 628.050 ;
        RECT 91.950 626.400 100.050 627.600 ;
        RECT 116.400 627.600 117.600 628.950 ;
        RECT 124.950 627.600 127.050 628.050 ;
        RECT 116.400 626.400 127.050 627.600 ;
        RECT 164.400 627.600 165.600 628.950 ;
        RECT 236.400 628.050 237.600 632.400 ;
        RECT 325.950 632.400 349.050 633.600 ;
        RECT 325.950 631.950 328.050 632.400 ;
        RECT 346.950 631.950 349.050 632.400 ;
        RECT 361.950 633.600 364.050 634.050 ;
        RECT 370.950 633.600 373.050 634.050 ;
        RECT 361.950 632.400 373.050 633.600 ;
        RECT 361.950 631.950 364.050 632.400 ;
        RECT 370.950 631.950 373.050 632.400 ;
        RECT 376.950 633.600 379.050 634.050 ;
        RECT 391.950 633.600 394.050 634.050 ;
        RECT 427.950 633.600 430.050 634.050 ;
        RECT 376.950 632.400 430.050 633.600 ;
        RECT 376.950 631.950 379.050 632.400 ;
        RECT 391.950 631.950 394.050 632.400 ;
        RECT 427.950 631.950 430.050 632.400 ;
        RECT 460.950 633.600 463.050 634.050 ;
        RECT 472.950 633.600 475.050 634.050 ;
        RECT 502.950 633.600 505.050 634.050 ;
        RECT 460.950 632.400 505.050 633.600 ;
        RECT 460.950 631.950 463.050 632.400 ;
        RECT 472.950 631.950 475.050 632.400 ;
        RECT 502.950 631.950 505.050 632.400 ;
        RECT 532.950 633.600 535.050 634.050 ;
        RECT 550.950 633.600 553.050 634.050 ;
        RECT 553.950 633.600 556.050 634.050 ;
        RECT 532.950 632.400 556.050 633.600 ;
        RECT 532.950 631.950 535.050 632.400 ;
        RECT 550.950 631.950 553.050 632.400 ;
        RECT 553.950 631.950 556.050 632.400 ;
        RECT 559.950 631.950 562.050 634.050 ;
        RECT 565.950 633.600 568.050 634.050 ;
        RECT 643.950 633.600 646.050 634.050 ;
        RECT 565.950 632.400 646.050 633.600 ;
        RECT 565.950 631.950 568.050 632.400 ;
        RECT 643.950 631.950 646.050 632.400 ;
        RECT 661.950 633.600 664.050 634.050 ;
        RECT 667.950 633.600 670.050 634.050 ;
        RECT 715.950 633.600 718.050 634.050 ;
        RECT 661.950 632.400 670.050 633.600 ;
        RECT 661.950 631.950 664.050 632.400 ;
        RECT 667.950 631.950 670.050 632.400 ;
        RECT 680.400 632.400 718.050 633.600 ;
        RECT 238.950 630.600 241.050 631.050 ;
        RECT 247.950 630.600 250.050 631.050 ;
        RECT 238.950 629.400 250.050 630.600 ;
        RECT 238.950 628.950 241.050 629.400 ;
        RECT 247.950 628.950 250.050 629.400 ;
        RECT 262.950 628.950 265.050 631.050 ;
        RECT 307.950 630.600 310.050 631.050 ;
        RECT 316.950 630.600 319.050 631.050 ;
        RECT 373.950 630.600 376.050 631.050 ;
        RECT 385.950 630.600 388.050 631.050 ;
        RECT 307.950 629.400 330.600 630.600 ;
        RECT 307.950 628.950 310.050 629.400 ;
        RECT 316.950 628.950 319.050 629.400 ;
        RECT 172.950 627.600 175.050 628.050 ;
        RECT 199.950 627.600 202.050 628.050 ;
        RECT 164.400 626.400 175.050 627.600 ;
        RECT 91.950 625.950 94.050 626.400 ;
        RECT 97.950 625.950 100.050 626.400 ;
        RECT 124.950 625.950 127.050 626.400 ;
        RECT 172.950 625.950 175.050 626.400 ;
        RECT 176.400 626.400 202.050 627.600 ;
        RECT 88.950 624.600 91.050 625.050 ;
        RECT 94.950 624.600 97.050 625.050 ;
        RECT 112.950 624.600 115.050 625.050 ;
        RECT 88.950 623.400 115.050 624.600 ;
        RECT 88.950 622.950 91.050 623.400 ;
        RECT 94.950 622.950 97.050 623.400 ;
        RECT 112.950 622.950 115.050 623.400 ;
        RECT 130.950 624.600 133.050 625.050 ;
        RECT 136.950 624.600 139.050 625.050 ;
        RECT 176.400 624.600 177.600 626.400 ;
        RECT 199.950 625.950 202.050 626.400 ;
        RECT 235.950 625.950 238.050 628.050 ;
        RECT 241.950 627.600 244.050 628.050 ;
        RECT 263.400 627.600 264.600 628.950 ;
        RECT 286.950 627.600 289.050 628.050 ;
        RECT 241.950 626.400 258.600 627.600 ;
        RECT 263.400 626.400 289.050 627.600 ;
        RECT 241.950 625.950 244.050 626.400 ;
        RECT 130.950 623.400 177.600 624.600 ;
        RECT 181.950 624.600 184.050 625.050 ;
        RECT 184.950 624.600 187.050 625.050 ;
        RECT 193.950 624.600 196.050 625.050 ;
        RECT 181.950 623.400 196.050 624.600 ;
        RECT 130.950 622.950 133.050 623.400 ;
        RECT 136.950 622.950 139.050 623.400 ;
        RECT 181.950 622.950 184.050 623.400 ;
        RECT 184.950 622.950 187.050 623.400 ;
        RECT 193.950 622.950 196.050 623.400 ;
        RECT 196.950 624.600 199.050 625.050 ;
        RECT 220.950 624.600 223.050 625.050 ;
        RECT 196.950 623.400 223.050 624.600 ;
        RECT 196.950 622.950 199.050 623.400 ;
        RECT 220.950 622.950 223.050 623.400 ;
        RECT 229.950 624.600 232.050 625.050 ;
        RECT 253.950 624.600 256.050 625.050 ;
        RECT 229.950 623.400 256.050 624.600 ;
        RECT 257.400 624.600 258.600 626.400 ;
        RECT 286.950 625.950 289.050 626.400 ;
        RECT 298.950 627.600 301.050 628.050 ;
        RECT 304.950 627.600 307.050 628.050 ;
        RECT 298.950 626.400 307.050 627.600 ;
        RECT 329.400 627.600 330.600 629.400 ;
        RECT 373.950 629.400 388.050 630.600 ;
        RECT 373.950 628.950 376.050 629.400 ;
        RECT 385.950 628.950 388.050 629.400 ;
        RECT 454.950 630.600 457.050 631.050 ;
        RECT 469.950 630.600 472.050 631.050 ;
        RECT 454.950 629.400 472.050 630.600 ;
        RECT 454.950 628.950 457.050 629.400 ;
        RECT 469.950 628.950 472.050 629.400 ;
        RECT 535.950 630.600 538.050 631.050 ;
        RECT 544.950 630.600 547.050 631.050 ;
        RECT 535.950 629.400 547.050 630.600 ;
        RECT 535.950 628.950 538.050 629.400 ;
        RECT 544.950 628.950 547.050 629.400 ;
        RECT 340.950 627.600 343.050 628.050 ;
        RECT 329.400 626.400 343.050 627.600 ;
        RECT 298.950 625.950 301.050 626.400 ;
        RECT 304.950 625.950 307.050 626.400 ;
        RECT 340.950 625.950 343.050 626.400 ;
        RECT 394.950 627.600 397.050 628.050 ;
        RECT 421.950 627.600 424.050 628.050 ;
        RECT 394.950 626.400 424.050 627.600 ;
        RECT 394.950 625.950 397.050 626.400 ;
        RECT 421.950 625.950 424.050 626.400 ;
        RECT 433.950 627.600 436.050 628.050 ;
        RECT 457.950 627.600 460.050 628.050 ;
        RECT 433.950 626.400 460.050 627.600 ;
        RECT 433.950 625.950 436.050 626.400 ;
        RECT 457.950 625.950 460.050 626.400 ;
        RECT 466.950 627.600 469.050 628.050 ;
        RECT 481.950 627.600 484.050 628.050 ;
        RECT 511.950 627.600 514.050 628.050 ;
        RECT 466.950 626.400 514.050 627.600 ;
        RECT 466.950 625.950 469.050 626.400 ;
        RECT 481.950 625.950 484.050 626.400 ;
        RECT 511.950 625.950 514.050 626.400 ;
        RECT 520.950 627.600 523.050 628.050 ;
        RECT 529.950 627.600 532.050 628.050 ;
        RECT 520.950 626.400 532.050 627.600 ;
        RECT 560.400 627.600 561.600 631.950 ;
        RECT 680.400 631.050 681.600 632.400 ;
        RECT 715.950 631.950 718.050 632.400 ;
        RECT 727.950 631.950 730.050 634.050 ;
        RECT 562.950 630.600 565.050 631.050 ;
        RECT 571.950 630.600 574.050 631.050 ;
        RECT 562.950 629.400 574.050 630.600 ;
        RECT 562.950 628.950 565.050 629.400 ;
        RECT 571.950 628.950 574.050 629.400 ;
        RECT 577.950 628.950 580.050 631.050 ;
        RECT 592.950 630.600 595.050 631.050 ;
        RECT 581.400 629.400 595.050 630.600 ;
        RECT 578.400 627.600 579.600 628.950 ;
        RECT 581.400 628.050 582.600 629.400 ;
        RECT 592.950 628.950 595.050 629.400 ;
        RECT 598.950 628.950 601.050 631.050 ;
        RECT 658.950 630.600 661.050 631.050 ;
        RECT 653.400 629.400 661.050 630.600 ;
        RECT 560.400 626.400 579.600 627.600 ;
        RECT 520.950 625.950 523.050 626.400 ;
        RECT 529.950 625.950 532.050 626.400 ;
        RECT 262.950 624.600 265.050 625.050 ;
        RECT 325.950 624.600 328.050 625.050 ;
        RECT 257.400 623.400 328.050 624.600 ;
        RECT 229.950 622.950 232.050 623.400 ;
        RECT 253.950 622.950 256.050 623.400 ;
        RECT 262.950 622.950 265.050 623.400 ;
        RECT 325.950 622.950 328.050 623.400 ;
        RECT 328.950 624.600 331.050 625.050 ;
        RECT 343.950 624.600 346.050 625.050 ;
        RECT 328.950 623.400 346.050 624.600 ;
        RECT 328.950 622.950 331.050 623.400 ;
        RECT 343.950 622.950 346.050 623.400 ;
        RECT 427.950 624.600 430.050 625.050 ;
        RECT 442.950 624.600 445.050 625.050 ;
        RECT 427.950 623.400 445.050 624.600 ;
        RECT 427.950 622.950 430.050 623.400 ;
        RECT 442.950 622.950 445.050 623.400 ;
        RECT 499.950 624.600 502.050 625.050 ;
        RECT 547.950 624.600 550.050 625.050 ;
        RECT 499.950 623.400 550.050 624.600 ;
        RECT 578.400 624.600 579.600 626.400 ;
        RECT 580.950 625.950 583.050 628.050 ;
        RECT 589.950 627.600 592.050 628.050 ;
        RECT 599.400 627.600 600.600 628.950 ;
        RECT 653.400 628.050 654.600 629.400 ;
        RECT 658.950 628.950 661.050 629.400 ;
        RECT 670.950 630.600 673.050 631.050 ;
        RECT 676.950 630.600 679.050 631.050 ;
        RECT 670.950 629.400 679.050 630.600 ;
        RECT 670.950 628.950 673.050 629.400 ;
        RECT 676.950 628.950 679.050 629.400 ;
        RECT 679.950 628.950 682.050 631.050 ;
        RECT 703.950 628.950 706.050 631.050 ;
        RECT 728.400 630.600 729.600 631.950 ;
        RECT 722.400 629.400 729.600 630.600 ;
        RECT 589.950 626.400 600.600 627.600 ;
        RECT 601.950 627.600 604.050 628.050 ;
        RECT 622.950 627.600 625.050 628.050 ;
        RECT 601.950 626.400 625.050 627.600 ;
        RECT 589.950 625.950 592.050 626.400 ;
        RECT 601.950 625.950 604.050 626.400 ;
        RECT 622.950 625.950 625.050 626.400 ;
        RECT 640.950 627.600 643.050 628.050 ;
        RECT 646.950 627.600 649.050 628.050 ;
        RECT 640.950 626.400 649.050 627.600 ;
        RECT 640.950 625.950 643.050 626.400 ;
        RECT 646.950 625.950 649.050 626.400 ;
        RECT 652.950 625.950 655.050 628.050 ;
        RECT 673.950 627.600 676.050 628.050 ;
        RECT 682.950 627.600 685.050 628.050 ;
        RECT 673.950 626.400 685.050 627.600 ;
        RECT 673.950 625.950 676.050 626.400 ;
        RECT 682.950 625.950 685.050 626.400 ;
        RECT 625.950 624.600 628.050 625.050 ;
        RECT 578.400 623.400 628.050 624.600 ;
        RECT 499.950 622.950 502.050 623.400 ;
        RECT 547.950 622.950 550.050 623.400 ;
        RECT 625.950 622.950 628.050 623.400 ;
        RECT 658.950 624.600 661.050 625.050 ;
        RECT 667.950 624.600 670.050 625.050 ;
        RECT 658.950 623.400 670.050 624.600 ;
        RECT 658.950 622.950 661.050 623.400 ;
        RECT 667.950 622.950 670.050 623.400 ;
        RECT 679.950 624.600 682.050 625.050 ;
        RECT 685.950 624.600 688.050 625.050 ;
        RECT 679.950 623.400 688.050 624.600 ;
        RECT 679.950 622.950 682.050 623.400 ;
        RECT 685.950 622.950 688.050 623.400 ;
        RECT 34.950 620.400 75.600 621.600 ;
        RECT 103.950 621.600 106.050 622.050 ;
        RECT 109.950 621.600 112.050 622.050 ;
        RECT 160.950 621.600 163.050 622.050 ;
        RECT 103.950 620.400 163.050 621.600 ;
        RECT 34.950 619.950 37.050 620.400 ;
        RECT 103.950 619.950 106.050 620.400 ;
        RECT 109.950 619.950 112.050 620.400 ;
        RECT 160.950 619.950 163.050 620.400 ;
        RECT 166.950 621.600 169.050 622.050 ;
        RECT 175.950 621.600 178.050 622.050 ;
        RECT 166.950 620.400 178.050 621.600 ;
        RECT 166.950 619.950 169.050 620.400 ;
        RECT 175.950 619.950 178.050 620.400 ;
        RECT 190.950 621.600 193.050 622.050 ;
        RECT 202.950 621.600 205.050 622.050 ;
        RECT 190.950 620.400 205.050 621.600 ;
        RECT 190.950 619.950 193.050 620.400 ;
        RECT 202.950 619.950 205.050 620.400 ;
        RECT 232.950 621.600 235.050 622.050 ;
        RECT 250.950 621.600 253.050 622.050 ;
        RECT 232.950 620.400 253.050 621.600 ;
        RECT 232.950 619.950 235.050 620.400 ;
        RECT 250.950 619.950 253.050 620.400 ;
        RECT 256.950 621.600 259.050 622.050 ;
        RECT 265.950 621.600 268.050 622.050 ;
        RECT 256.950 620.400 268.050 621.600 ;
        RECT 256.950 619.950 259.050 620.400 ;
        RECT 265.950 619.950 268.050 620.400 ;
        RECT 274.950 621.600 277.050 622.050 ;
        RECT 298.950 621.600 301.050 622.050 ;
        RECT 274.950 620.400 301.050 621.600 ;
        RECT 274.950 619.950 277.050 620.400 ;
        RECT 298.950 619.950 301.050 620.400 ;
        RECT 319.950 621.600 322.050 622.050 ;
        RECT 382.950 621.600 385.050 622.050 ;
        RECT 403.950 621.600 406.050 622.050 ;
        RECT 319.950 620.400 406.050 621.600 ;
        RECT 319.950 619.950 322.050 620.400 ;
        RECT 382.950 619.950 385.050 620.400 ;
        RECT 403.950 619.950 406.050 620.400 ;
        RECT 607.950 621.600 610.050 622.050 ;
        RECT 613.950 621.600 616.050 622.050 ;
        RECT 607.950 620.400 616.050 621.600 ;
        RECT 607.950 619.950 610.050 620.400 ;
        RECT 613.950 619.950 616.050 620.400 ;
        RECT 625.950 621.600 628.050 622.050 ;
        RECT 704.400 621.600 705.600 628.950 ;
        RECT 722.400 628.050 723.600 629.400 ;
        RECT 730.950 628.950 733.050 631.050 ;
        RECT 742.950 630.600 745.050 631.050 ;
        RECT 734.400 629.400 745.050 630.600 ;
        RECT 721.950 625.950 724.050 628.050 ;
        RECT 724.950 624.600 727.050 625.050 ;
        RECT 731.400 624.600 732.600 628.950 ;
        RECT 734.400 628.050 735.600 629.400 ;
        RECT 742.950 628.950 745.050 629.400 ;
        RECT 745.950 630.600 748.050 631.050 ;
        RECT 751.950 630.600 754.050 631.050 ;
        RECT 745.950 629.400 754.050 630.600 ;
        RECT 745.950 628.950 748.050 629.400 ;
        RECT 751.950 628.950 754.050 629.400 ;
        RECT 757.950 628.950 760.050 631.050 ;
        RECT 733.950 625.950 736.050 628.050 ;
        RECT 758.400 625.050 759.600 628.950 ;
        RECT 724.950 623.400 732.600 624.600 ;
        RECT 724.950 622.950 727.050 623.400 ;
        RECT 757.950 622.950 760.050 625.050 ;
        RECT 760.950 624.600 763.050 625.050 ;
        RECT 766.950 624.600 769.050 625.050 ;
        RECT 760.950 623.400 769.050 624.600 ;
        RECT 760.950 622.950 763.050 623.400 ;
        RECT 766.950 622.950 769.050 623.400 ;
        RECT 739.950 621.600 742.050 622.050 ;
        RECT 625.950 620.400 742.050 621.600 ;
        RECT 625.950 619.950 628.050 620.400 ;
        RECT 739.950 619.950 742.050 620.400 ;
        RECT 145.950 618.600 148.050 619.050 ;
        RECT 151.950 618.600 154.050 619.050 ;
        RECT 145.950 617.400 154.050 618.600 ;
        RECT 145.950 616.950 148.050 617.400 ;
        RECT 151.950 616.950 154.050 617.400 ;
        RECT 172.950 618.600 175.050 619.050 ;
        RECT 208.950 618.600 211.050 619.050 ;
        RECT 172.950 617.400 211.050 618.600 ;
        RECT 172.950 616.950 175.050 617.400 ;
        RECT 208.950 616.950 211.050 617.400 ;
        RECT 211.950 618.600 214.050 619.050 ;
        RECT 214.950 618.600 217.050 619.050 ;
        RECT 238.950 618.600 241.050 619.050 ;
        RECT 259.950 618.600 262.050 619.050 ;
        RECT 352.950 618.600 355.050 619.050 ;
        RECT 211.950 617.400 355.050 618.600 ;
        RECT 211.950 616.950 214.050 617.400 ;
        RECT 214.950 616.950 217.050 617.400 ;
        RECT 238.950 616.950 241.050 617.400 ;
        RECT 259.950 616.950 262.050 617.400 ;
        RECT 352.950 616.950 355.050 617.400 ;
        RECT 409.950 618.600 412.050 619.050 ;
        RECT 538.950 618.600 541.050 619.050 ;
        RECT 409.950 617.400 541.050 618.600 ;
        RECT 409.950 616.950 412.050 617.400 ;
        RECT 538.950 616.950 541.050 617.400 ;
        RECT 577.950 618.600 580.050 619.050 ;
        RECT 586.950 618.600 589.050 619.050 ;
        RECT 577.950 617.400 589.050 618.600 ;
        RECT 577.950 616.950 580.050 617.400 ;
        RECT 586.950 616.950 589.050 617.400 ;
        RECT 667.950 618.600 670.050 619.050 ;
        RECT 676.950 618.600 679.050 619.050 ;
        RECT 667.950 617.400 679.050 618.600 ;
        RECT 667.950 616.950 670.050 617.400 ;
        RECT 676.950 616.950 679.050 617.400 ;
        RECT 682.950 618.600 685.050 619.050 ;
        RECT 715.950 618.600 718.050 619.050 ;
        RECT 682.950 617.400 718.050 618.600 ;
        RECT 682.950 616.950 685.050 617.400 ;
        RECT 715.950 616.950 718.050 617.400 ;
        RECT 61.950 615.600 64.050 616.050 ;
        RECT 241.950 615.600 244.050 616.050 ;
        RECT 61.950 614.400 244.050 615.600 ;
        RECT 61.950 613.950 64.050 614.400 ;
        RECT 241.950 613.950 244.050 614.400 ;
        RECT 244.950 615.600 247.050 616.050 ;
        RECT 322.950 615.600 325.050 616.050 ;
        RECT 244.950 614.400 325.050 615.600 ;
        RECT 244.950 613.950 247.050 614.400 ;
        RECT 322.950 613.950 325.050 614.400 ;
        RECT 325.950 615.600 328.050 616.050 ;
        RECT 430.950 615.600 433.050 616.050 ;
        RECT 325.950 614.400 433.050 615.600 ;
        RECT 325.950 613.950 328.050 614.400 ;
        RECT 430.950 613.950 433.050 614.400 ;
        RECT 505.950 615.600 508.050 616.050 ;
        RECT 514.950 615.600 517.050 616.050 ;
        RECT 505.950 614.400 517.050 615.600 ;
        RECT 505.950 613.950 508.050 614.400 ;
        RECT 514.950 613.950 517.050 614.400 ;
        RECT 517.950 615.600 520.050 616.050 ;
        RECT 562.950 615.600 565.050 616.050 ;
        RECT 646.950 615.600 649.050 616.050 ;
        RECT 517.950 614.400 649.050 615.600 ;
        RECT 517.950 613.950 520.050 614.400 ;
        RECT 562.950 613.950 565.050 614.400 ;
        RECT 646.950 613.950 649.050 614.400 ;
        RECT 655.950 615.600 658.050 616.050 ;
        RECT 700.950 615.600 703.050 616.050 ;
        RECT 655.950 614.400 703.050 615.600 ;
        RECT 655.950 613.950 658.050 614.400 ;
        RECT 700.950 613.950 703.050 614.400 ;
        RECT 706.950 615.600 709.050 616.050 ;
        RECT 724.950 615.600 727.050 616.050 ;
        RECT 706.950 614.400 727.050 615.600 ;
        RECT 706.950 613.950 709.050 614.400 ;
        RECT 724.950 613.950 727.050 614.400 ;
        RECT 169.950 612.600 172.050 613.050 ;
        RECT 196.950 612.600 199.050 613.050 ;
        RECT 169.950 611.400 199.050 612.600 ;
        RECT 169.950 610.950 172.050 611.400 ;
        RECT 196.950 610.950 199.050 611.400 ;
        RECT 199.950 612.600 202.050 613.050 ;
        RECT 361.950 612.600 364.050 613.050 ;
        RECT 199.950 611.400 364.050 612.600 ;
        RECT 199.950 610.950 202.050 611.400 ;
        RECT 361.950 610.950 364.050 611.400 ;
        RECT 373.950 612.600 376.050 613.050 ;
        RECT 466.950 612.600 469.050 613.050 ;
        RECT 373.950 611.400 469.050 612.600 ;
        RECT 373.950 610.950 376.050 611.400 ;
        RECT 466.950 610.950 469.050 611.400 ;
        RECT 514.950 612.600 517.050 613.050 ;
        RECT 583.950 612.600 586.050 613.050 ;
        RECT 622.950 612.600 625.050 613.050 ;
        RECT 514.950 611.400 625.050 612.600 ;
        RECT 514.950 610.950 517.050 611.400 ;
        RECT 583.950 610.950 586.050 611.400 ;
        RECT 622.950 610.950 625.050 611.400 ;
        RECT 655.950 612.600 658.050 613.050 ;
        RECT 661.950 612.600 664.050 613.050 ;
        RECT 655.950 611.400 664.050 612.600 ;
        RECT 655.950 610.950 658.050 611.400 ;
        RECT 661.950 610.950 664.050 611.400 ;
        RECT 694.950 612.600 697.050 613.050 ;
        RECT 700.950 612.600 703.050 613.050 ;
        RECT 769.950 612.600 772.050 613.050 ;
        RECT 694.950 611.400 699.600 612.600 ;
        RECT 694.950 610.950 697.050 611.400 ;
        RECT 94.950 609.600 97.050 610.050 ;
        RECT 106.950 609.600 109.050 610.050 ;
        RECT 115.950 609.600 118.050 610.050 ;
        RECT 94.950 608.400 118.050 609.600 ;
        RECT 94.950 607.950 97.050 608.400 ;
        RECT 106.950 607.950 109.050 608.400 ;
        RECT 115.950 607.950 118.050 608.400 ;
        RECT 208.950 609.600 211.050 610.050 ;
        RECT 250.950 609.600 253.050 610.050 ;
        RECT 208.950 608.400 253.050 609.600 ;
        RECT 208.950 607.950 211.050 608.400 ;
        RECT 250.950 607.950 253.050 608.400 ;
        RECT 253.950 609.600 256.050 610.050 ;
        RECT 274.950 609.600 277.050 610.050 ;
        RECT 253.950 608.400 277.050 609.600 ;
        RECT 253.950 607.950 256.050 608.400 ;
        RECT 274.950 607.950 277.050 608.400 ;
        RECT 301.950 609.600 304.050 610.050 ;
        RECT 322.950 609.600 325.050 610.050 ;
        RECT 331.950 609.600 334.050 610.050 ;
        RECT 301.950 608.400 334.050 609.600 ;
        RECT 301.950 607.950 304.050 608.400 ;
        RECT 322.950 607.950 325.050 608.400 ;
        RECT 331.950 607.950 334.050 608.400 ;
        RECT 364.950 609.600 367.050 610.050 ;
        RECT 406.950 609.600 409.050 610.050 ;
        RECT 442.950 609.600 445.050 610.050 ;
        RECT 364.950 608.400 445.050 609.600 ;
        RECT 364.950 607.950 367.050 608.400 ;
        RECT 406.950 607.950 409.050 608.400 ;
        RECT 442.950 607.950 445.050 608.400 ;
        RECT 574.950 609.600 577.050 610.050 ;
        RECT 586.950 609.600 589.050 610.050 ;
        RECT 574.950 608.400 589.050 609.600 ;
        RECT 574.950 607.950 577.050 608.400 ;
        RECT 586.950 607.950 589.050 608.400 ;
        RECT 634.950 609.600 637.050 610.050 ;
        RECT 670.950 609.600 673.050 610.050 ;
        RECT 634.950 608.400 673.050 609.600 ;
        RECT 698.400 609.600 699.600 611.400 ;
        RECT 700.950 611.400 772.050 612.600 ;
        RECT 700.950 610.950 703.050 611.400 ;
        RECT 769.950 610.950 772.050 611.400 ;
        RECT 709.950 609.600 712.050 610.050 ;
        RECT 698.400 608.400 712.050 609.600 ;
        RECT 634.950 607.950 637.050 608.400 ;
        RECT 670.950 607.950 673.050 608.400 ;
        RECT 709.950 607.950 712.050 608.400 ;
        RECT 13.950 606.600 16.050 607.050 ;
        RECT 64.950 606.600 67.050 607.050 ;
        RECT 88.950 606.600 91.050 607.050 ;
        RECT 259.950 606.600 262.050 607.050 ;
        RECT 13.950 605.400 262.050 606.600 ;
        RECT 13.950 604.950 16.050 605.400 ;
        RECT 64.950 604.950 67.050 605.400 ;
        RECT 88.950 604.950 91.050 605.400 ;
        RECT 259.950 604.950 262.050 605.400 ;
        RECT 286.950 606.600 289.050 607.050 ;
        RECT 328.950 606.600 331.050 607.050 ;
        RECT 286.950 605.400 331.050 606.600 ;
        RECT 286.950 604.950 289.050 605.400 ;
        RECT 328.950 604.950 331.050 605.400 ;
        RECT 493.950 606.600 496.050 607.050 ;
        RECT 550.950 606.600 553.050 607.050 ;
        RECT 493.950 605.400 553.050 606.600 ;
        RECT 493.950 604.950 496.050 605.400 ;
        RECT 550.950 604.950 553.050 605.400 ;
        RECT 553.950 606.600 556.050 607.050 ;
        RECT 583.950 606.600 586.050 607.050 ;
        RECT 553.950 605.400 586.050 606.600 ;
        RECT 553.950 604.950 556.050 605.400 ;
        RECT 583.950 604.950 586.050 605.400 ;
        RECT 619.950 606.600 622.050 607.050 ;
        RECT 652.950 606.600 655.050 607.050 ;
        RECT 619.950 605.400 655.050 606.600 ;
        RECT 619.950 604.950 622.050 605.400 ;
        RECT 652.950 604.950 655.050 605.400 ;
        RECT 661.950 606.600 664.050 607.050 ;
        RECT 673.950 606.600 676.050 607.050 ;
        RECT 661.950 605.400 676.050 606.600 ;
        RECT 661.950 604.950 664.050 605.400 ;
        RECT 673.950 604.950 676.050 605.400 ;
        RECT 730.950 606.600 733.050 607.050 ;
        RECT 736.950 606.600 739.050 607.050 ;
        RECT 730.950 605.400 739.050 606.600 ;
        RECT 730.950 604.950 733.050 605.400 ;
        RECT 736.950 604.950 739.050 605.400 ;
        RECT 754.950 606.600 757.050 607.050 ;
        RECT 769.950 606.600 772.050 607.050 ;
        RECT 754.950 605.400 772.050 606.600 ;
        RECT 754.950 604.950 757.050 605.400 ;
        RECT 769.950 604.950 772.050 605.400 ;
        RECT 28.950 603.600 31.050 604.050 ;
        RECT 40.950 603.600 43.050 604.050 ;
        RECT 28.950 602.400 43.050 603.600 ;
        RECT 28.950 601.950 31.050 602.400 ;
        RECT 40.950 601.950 43.050 602.400 ;
        RECT 52.950 603.600 55.050 604.050 ;
        RECT 67.950 603.600 70.050 604.050 ;
        RECT 52.950 602.400 70.050 603.600 ;
        RECT 52.950 601.950 55.050 602.400 ;
        RECT 67.950 601.950 70.050 602.400 ;
        RECT 169.950 601.950 172.050 604.050 ;
        RECT 181.950 603.600 184.050 604.050 ;
        RECT 187.950 603.600 190.050 604.050 ;
        RECT 181.950 602.400 190.050 603.600 ;
        RECT 181.950 601.950 184.050 602.400 ;
        RECT 187.950 601.950 190.050 602.400 ;
        RECT 217.950 603.600 220.050 604.050 ;
        RECT 256.950 603.600 259.050 604.050 ;
        RECT 295.950 603.600 298.050 604.050 ;
        RECT 217.950 602.400 298.050 603.600 ;
        RECT 217.950 601.950 220.050 602.400 ;
        RECT 256.950 601.950 259.050 602.400 ;
        RECT 295.950 601.950 298.050 602.400 ;
        RECT 310.950 603.600 313.050 604.050 ;
        RECT 319.950 603.600 322.050 604.050 ;
        RECT 310.950 602.400 322.050 603.600 ;
        RECT 310.950 601.950 313.050 602.400 ;
        RECT 319.950 601.950 322.050 602.400 ;
        RECT 328.950 603.600 331.050 604.050 ;
        RECT 343.950 603.600 346.050 604.050 ;
        RECT 328.950 602.400 346.050 603.600 ;
        RECT 328.950 601.950 331.050 602.400 ;
        RECT 343.950 601.950 346.050 602.400 ;
        RECT 346.950 603.600 349.050 604.050 ;
        RECT 355.950 603.600 358.050 604.050 ;
        RECT 346.950 602.400 358.050 603.600 ;
        RECT 346.950 601.950 349.050 602.400 ;
        RECT 355.950 601.950 358.050 602.400 ;
        RECT 463.950 603.600 466.050 604.050 ;
        RECT 472.950 603.600 475.050 604.050 ;
        RECT 463.950 602.400 475.050 603.600 ;
        RECT 463.950 601.950 466.050 602.400 ;
        RECT 472.950 601.950 475.050 602.400 ;
        RECT 526.950 603.600 529.050 604.050 ;
        RECT 535.950 603.600 538.050 604.050 ;
        RECT 526.950 602.400 538.050 603.600 ;
        RECT 526.950 601.950 529.050 602.400 ;
        RECT 535.950 601.950 538.050 602.400 ;
        RECT 550.950 603.600 553.050 604.050 ;
        RECT 553.950 603.600 556.050 604.050 ;
        RECT 592.950 603.600 595.050 604.050 ;
        RECT 652.950 603.600 655.050 604.050 ;
        RECT 661.950 603.600 664.050 604.050 ;
        RECT 550.950 602.400 595.050 603.600 ;
        RECT 550.950 601.950 553.050 602.400 ;
        RECT 553.950 601.950 556.050 602.400 ;
        RECT 592.950 601.950 595.050 602.400 ;
        RECT 641.400 602.400 664.050 603.600 ;
        RECT 10.950 600.600 13.050 601.050 ;
        RECT 19.950 600.600 22.050 601.050 ;
        RECT 10.950 599.400 22.050 600.600 ;
        RECT 10.950 598.950 13.050 599.400 ;
        RECT 19.950 598.950 22.050 599.400 ;
        RECT 31.950 598.950 34.050 601.050 ;
        RECT 37.950 600.600 40.050 601.050 ;
        RECT 49.950 600.600 52.050 601.050 ;
        RECT 64.950 600.600 67.050 601.050 ;
        RECT 37.950 599.400 67.050 600.600 ;
        RECT 37.950 598.950 40.050 599.400 ;
        RECT 49.950 598.950 52.050 599.400 ;
        RECT 64.950 598.950 67.050 599.400 ;
        RECT 70.950 600.600 73.050 601.050 ;
        RECT 82.950 600.600 85.050 601.050 ;
        RECT 70.950 599.400 85.050 600.600 ;
        RECT 70.950 598.950 73.050 599.400 ;
        RECT 82.950 598.950 85.050 599.400 ;
        RECT 7.950 597.600 10.050 598.050 ;
        RECT 22.950 597.600 25.050 598.050 ;
        RECT 7.950 596.400 25.050 597.600 ;
        RECT 7.950 595.950 10.050 596.400 ;
        RECT 22.950 595.950 25.050 596.400 ;
        RECT 25.950 597.600 28.050 598.050 ;
        RECT 32.400 597.600 33.600 598.950 ;
        RECT 170.400 598.050 171.600 601.950 ;
        RECT 202.950 600.600 205.050 601.050 ;
        RECT 217.950 600.600 220.050 601.050 ;
        RECT 173.400 599.400 205.050 600.600 ;
        RECT 25.950 596.400 33.600 597.600 ;
        RECT 55.950 597.600 58.050 598.050 ;
        RECT 88.950 597.600 91.050 598.050 ;
        RECT 55.950 596.400 91.050 597.600 ;
        RECT 25.950 595.950 28.050 596.400 ;
        RECT 55.950 595.950 58.050 596.400 ;
        RECT 88.950 595.950 91.050 596.400 ;
        RECT 100.950 597.600 103.050 598.050 ;
        RECT 106.950 597.600 109.050 598.050 ;
        RECT 100.950 596.400 109.050 597.600 ;
        RECT 100.950 595.950 103.050 596.400 ;
        RECT 106.950 595.950 109.050 596.400 ;
        RECT 169.950 595.950 172.050 598.050 ;
        RECT 22.950 594.600 25.050 595.050 ;
        RECT 34.950 594.600 37.050 595.050 ;
        RECT 22.950 593.400 37.050 594.600 ;
        RECT 22.950 592.950 25.050 593.400 ;
        RECT 34.950 592.950 37.050 593.400 ;
        RECT 58.950 594.600 61.050 595.050 ;
        RECT 67.950 594.600 70.050 595.050 ;
        RECT 58.950 593.400 70.050 594.600 ;
        RECT 58.950 592.950 61.050 593.400 ;
        RECT 67.950 592.950 70.050 593.400 ;
        RECT 85.950 594.600 88.050 595.050 ;
        RECT 97.950 594.600 100.050 595.050 ;
        RECT 85.950 593.400 100.050 594.600 ;
        RECT 85.950 592.950 88.050 593.400 ;
        RECT 97.950 592.950 100.050 593.400 ;
        RECT 109.950 594.600 112.050 595.050 ;
        RECT 163.950 594.600 166.050 595.050 ;
        RECT 109.950 593.400 166.050 594.600 ;
        RECT 109.950 592.950 112.050 593.400 ;
        RECT 163.950 592.950 166.050 593.400 ;
        RECT 166.950 594.600 169.050 595.050 ;
        RECT 173.400 594.600 174.600 599.400 ;
        RECT 202.950 598.950 205.050 599.400 ;
        RECT 206.400 599.400 220.050 600.600 ;
        RECT 206.400 598.050 207.600 599.400 ;
        RECT 217.950 598.950 220.050 599.400 ;
        RECT 223.950 600.600 226.050 601.050 ;
        RECT 232.950 600.600 235.050 601.050 ;
        RECT 223.950 599.400 235.050 600.600 ;
        RECT 223.950 598.950 226.050 599.400 ;
        RECT 232.950 598.950 235.050 599.400 ;
        RECT 235.950 598.950 238.050 601.050 ;
        RECT 265.950 600.600 268.050 601.050 ;
        RECT 248.400 599.400 268.050 600.600 ;
        RECT 187.950 597.600 190.050 598.050 ;
        RECT 199.950 597.600 202.050 598.050 ;
        RECT 187.950 596.400 202.050 597.600 ;
        RECT 187.950 595.950 190.050 596.400 ;
        RECT 199.950 595.950 202.050 596.400 ;
        RECT 205.950 595.950 208.050 598.050 ;
        RECT 220.950 597.600 223.050 598.050 ;
        RECT 236.400 597.600 237.600 598.950 ;
        RECT 248.400 598.050 249.600 599.400 ;
        RECT 265.950 598.950 268.050 599.400 ;
        RECT 274.950 600.600 277.050 601.050 ;
        RECT 283.950 600.600 286.050 601.050 ;
        RECT 274.950 599.400 286.050 600.600 ;
        RECT 274.950 598.950 277.050 599.400 ;
        RECT 283.950 598.950 286.050 599.400 ;
        RECT 289.950 600.600 292.050 601.050 ;
        RECT 304.950 600.600 307.050 601.050 ;
        RECT 373.950 600.600 376.050 601.050 ;
        RECT 289.950 599.400 376.050 600.600 ;
        RECT 289.950 598.950 292.050 599.400 ;
        RECT 304.950 598.950 307.050 599.400 ;
        RECT 373.950 598.950 376.050 599.400 ;
        RECT 394.950 600.600 397.050 601.050 ;
        RECT 427.950 600.600 430.050 601.050 ;
        RECT 394.950 599.400 430.050 600.600 ;
        RECT 394.950 598.950 397.050 599.400 ;
        RECT 427.950 598.950 430.050 599.400 ;
        RECT 433.950 600.600 436.050 601.050 ;
        RECT 463.950 600.600 466.050 601.050 ;
        RECT 472.950 600.600 475.050 601.050 ;
        RECT 487.950 600.600 490.050 601.050 ;
        RECT 433.950 599.400 466.050 600.600 ;
        RECT 433.950 598.950 436.050 599.400 ;
        RECT 463.950 598.950 466.050 599.400 ;
        RECT 467.400 599.400 475.050 600.600 ;
        RECT 220.950 596.400 246.600 597.600 ;
        RECT 220.950 595.950 223.050 596.400 ;
        RECT 245.400 595.050 246.600 596.400 ;
        RECT 247.950 595.950 250.050 598.050 ;
        RECT 283.950 597.600 286.050 598.050 ;
        RECT 292.950 597.600 295.050 598.050 ;
        RECT 283.950 596.400 295.050 597.600 ;
        RECT 283.950 595.950 286.050 596.400 ;
        RECT 166.950 593.400 174.600 594.600 ;
        RECT 190.950 594.600 193.050 595.050 ;
        RECT 196.950 594.600 199.050 595.050 ;
        RECT 208.950 594.600 211.050 595.050 ;
        RECT 190.950 593.400 211.050 594.600 ;
        RECT 166.950 592.950 169.050 593.400 ;
        RECT 190.950 592.950 193.050 593.400 ;
        RECT 196.950 592.950 199.050 593.400 ;
        RECT 208.950 592.950 211.050 593.400 ;
        RECT 229.950 594.600 232.050 595.050 ;
        RECT 241.950 594.600 244.050 595.050 ;
        RECT 229.950 593.400 244.050 594.600 ;
        RECT 229.950 592.950 232.050 593.400 ;
        RECT 241.950 592.950 244.050 593.400 ;
        RECT 244.950 592.950 247.050 595.050 ;
        RECT 262.950 594.600 265.050 595.050 ;
        RECT 268.950 594.600 271.050 595.050 ;
        RECT 262.950 593.400 271.050 594.600 ;
        RECT 262.950 592.950 265.050 593.400 ;
        RECT 268.950 592.950 271.050 593.400 ;
        RECT 271.950 594.600 274.050 595.050 ;
        RECT 280.950 594.600 283.050 595.050 ;
        RECT 271.950 593.400 283.050 594.600 ;
        RECT 271.950 592.950 274.050 593.400 ;
        RECT 280.950 592.950 283.050 593.400 ;
        RECT 214.950 591.600 217.050 592.050 ;
        RECT 262.950 591.600 265.050 592.050 ;
        RECT 214.950 590.400 265.050 591.600 ;
        RECT 290.400 591.600 291.600 596.400 ;
        RECT 292.950 595.950 295.050 596.400 ;
        RECT 316.950 597.600 319.050 598.050 ;
        RECT 325.950 597.600 328.050 598.050 ;
        RECT 316.950 596.400 328.050 597.600 ;
        RECT 316.950 595.950 319.050 596.400 ;
        RECT 325.950 595.950 328.050 596.400 ;
        RECT 334.950 597.600 337.050 598.050 ;
        RECT 352.950 597.600 355.050 598.050 ;
        RECT 334.950 596.400 355.050 597.600 ;
        RECT 334.950 595.950 337.050 596.400 ;
        RECT 352.950 595.950 355.050 596.400 ;
        RECT 358.950 597.600 361.050 598.050 ;
        RECT 367.950 597.600 370.050 598.050 ;
        RECT 358.950 596.400 370.050 597.600 ;
        RECT 358.950 595.950 361.050 596.400 ;
        RECT 367.950 595.950 370.050 596.400 ;
        RECT 370.950 597.600 373.050 598.050 ;
        RECT 409.950 597.600 412.050 598.050 ;
        RECT 370.950 596.400 412.050 597.600 ;
        RECT 370.950 595.950 373.050 596.400 ;
        RECT 409.950 595.950 412.050 596.400 ;
        RECT 451.950 597.600 454.050 598.050 ;
        RECT 463.950 597.600 466.050 598.050 ;
        RECT 451.950 596.400 466.050 597.600 ;
        RECT 451.950 595.950 454.050 596.400 ;
        RECT 463.950 595.950 466.050 596.400 ;
        RECT 292.950 594.600 295.050 595.050 ;
        RECT 400.950 594.600 403.050 595.050 ;
        RECT 292.950 593.400 403.050 594.600 ;
        RECT 467.400 594.600 468.600 599.400 ;
        RECT 472.950 598.950 475.050 599.400 ;
        RECT 476.400 599.400 490.050 600.600 ;
        RECT 469.950 597.600 472.050 598.050 ;
        RECT 476.400 597.600 477.600 599.400 ;
        RECT 487.950 598.950 490.050 599.400 ;
        RECT 493.950 600.600 496.050 601.050 ;
        RECT 523.950 600.600 526.050 601.050 ;
        RECT 493.950 599.400 526.050 600.600 ;
        RECT 493.950 598.950 496.050 599.400 ;
        RECT 523.950 598.950 526.050 599.400 ;
        RECT 529.950 600.600 532.050 601.050 ;
        RECT 559.950 600.600 562.050 601.050 ;
        RECT 529.950 599.400 562.050 600.600 ;
        RECT 529.950 598.950 532.050 599.400 ;
        RECT 559.950 598.950 562.050 599.400 ;
        RECT 469.950 596.400 477.600 597.600 ;
        RECT 517.950 597.600 520.050 598.050 ;
        RECT 526.950 597.600 529.050 598.050 ;
        RECT 517.950 596.400 529.050 597.600 ;
        RECT 469.950 595.950 472.050 596.400 ;
        RECT 517.950 595.950 520.050 596.400 ;
        RECT 526.950 595.950 529.050 596.400 ;
        RECT 583.950 597.600 586.050 598.050 ;
        RECT 589.950 597.600 592.050 598.050 ;
        RECT 613.950 597.600 616.050 598.050 ;
        RECT 583.950 596.400 616.050 597.600 ;
        RECT 583.950 595.950 586.050 596.400 ;
        RECT 589.950 595.950 592.050 596.400 ;
        RECT 613.950 595.950 616.050 596.400 ;
        RECT 628.950 597.600 631.050 598.050 ;
        RECT 637.950 597.600 640.050 598.050 ;
        RECT 628.950 596.400 640.050 597.600 ;
        RECT 628.950 595.950 631.050 596.400 ;
        RECT 637.950 595.950 640.050 596.400 ;
        RECT 641.400 595.050 642.600 602.400 ;
        RECT 652.950 601.950 655.050 602.400 ;
        RECT 661.950 601.950 664.050 602.400 ;
        RECT 664.950 603.600 667.050 604.050 ;
        RECT 688.950 603.600 691.050 604.050 ;
        RECT 664.950 602.400 691.050 603.600 ;
        RECT 664.950 601.950 667.050 602.400 ;
        RECT 688.950 601.950 691.050 602.400 ;
        RECT 727.950 603.600 730.050 604.050 ;
        RECT 739.950 603.600 742.050 604.050 ;
        RECT 748.950 603.600 751.050 604.050 ;
        RECT 727.950 602.400 738.600 603.600 ;
        RECT 727.950 601.950 730.050 602.400 ;
        RECT 649.950 598.950 652.050 601.050 ;
        RECT 655.950 600.600 658.050 601.050 ;
        RECT 667.950 600.600 670.050 601.050 ;
        RECT 655.950 599.400 660.600 600.600 ;
        RECT 655.950 598.950 658.050 599.400 ;
        RECT 650.400 597.600 651.600 598.950 ;
        RECT 652.950 597.600 655.050 598.050 ;
        RECT 650.400 596.400 655.050 597.600 ;
        RECT 652.950 595.950 655.050 596.400 ;
        RECT 478.950 594.600 481.050 595.050 ;
        RECT 467.400 593.400 481.050 594.600 ;
        RECT 292.950 592.950 295.050 593.400 ;
        RECT 400.950 592.950 403.050 593.400 ;
        RECT 478.950 592.950 481.050 593.400 ;
        RECT 505.950 594.600 508.050 595.050 ;
        RECT 511.950 594.600 514.050 595.050 ;
        RECT 505.950 593.400 514.050 594.600 ;
        RECT 505.950 592.950 508.050 593.400 ;
        RECT 511.950 592.950 514.050 593.400 ;
        RECT 514.950 594.600 517.050 595.050 ;
        RECT 532.950 594.600 535.050 595.050 ;
        RECT 514.950 593.400 535.050 594.600 ;
        RECT 514.950 592.950 517.050 593.400 ;
        RECT 532.950 592.950 535.050 593.400 ;
        RECT 610.950 594.600 613.050 595.050 ;
        RECT 634.950 594.600 637.050 595.050 ;
        RECT 610.950 593.400 637.050 594.600 ;
        RECT 610.950 592.950 613.050 593.400 ;
        RECT 634.950 592.950 637.050 593.400 ;
        RECT 640.950 592.950 643.050 595.050 ;
        RECT 659.400 594.600 660.600 599.400 ;
        RECT 662.400 599.400 670.050 600.600 ;
        RECT 662.400 598.050 663.600 599.400 ;
        RECT 667.950 598.950 670.050 599.400 ;
        RECT 679.950 600.600 682.050 601.050 ;
        RECT 703.950 600.600 706.050 601.050 ;
        RECT 715.950 600.600 718.050 601.050 ;
        RECT 727.950 600.600 730.050 601.050 ;
        RECT 733.950 600.600 736.050 601.050 ;
        RECT 679.950 599.400 702.600 600.600 ;
        RECT 679.950 598.950 682.050 599.400 ;
        RECT 661.950 595.950 664.050 598.050 ;
        RECT 664.950 597.600 667.050 598.050 ;
        RECT 676.950 597.600 679.050 598.050 ;
        RECT 664.950 596.400 679.050 597.600 ;
        RECT 701.400 597.600 702.600 599.400 ;
        RECT 703.950 599.400 736.050 600.600 ;
        RECT 703.950 598.950 706.050 599.400 ;
        RECT 715.950 598.950 718.050 599.400 ;
        RECT 727.950 598.950 730.050 599.400 ;
        RECT 733.950 598.950 736.050 599.400 ;
        RECT 706.950 597.600 709.050 598.050 ;
        RECT 701.400 596.400 709.050 597.600 ;
        RECT 664.950 595.950 667.050 596.400 ;
        RECT 676.950 595.950 679.050 596.400 ;
        RECT 706.950 595.950 709.050 596.400 ;
        RECT 724.950 597.600 727.050 598.050 ;
        RECT 737.400 597.600 738.600 602.400 ;
        RECT 739.950 602.400 751.050 603.600 ;
        RECT 739.950 601.950 742.050 602.400 ;
        RECT 748.950 601.950 751.050 602.400 ;
        RECT 751.950 603.600 754.050 604.050 ;
        RECT 763.950 603.600 766.050 604.050 ;
        RECT 751.950 602.400 766.050 603.600 ;
        RECT 751.950 601.950 754.050 602.400 ;
        RECT 763.950 601.950 766.050 602.400 ;
        RECT 757.950 600.600 760.050 601.050 ;
        RECT 755.400 599.400 760.050 600.600 ;
        RECT 724.950 596.400 738.600 597.600 ;
        RECT 724.950 595.950 727.050 596.400 ;
        RECT 742.950 595.950 745.050 598.050 ;
        RECT 745.950 597.600 748.050 598.050 ;
        RECT 751.950 597.600 754.050 598.050 ;
        RECT 745.950 596.400 754.050 597.600 ;
        RECT 745.950 595.950 748.050 596.400 ;
        RECT 751.950 595.950 754.050 596.400 ;
        RECT 667.950 594.600 670.050 595.050 ;
        RECT 659.400 593.400 670.050 594.600 ;
        RECT 667.950 592.950 670.050 593.400 ;
        RECT 688.950 594.600 691.050 595.050 ;
        RECT 697.950 594.600 700.050 595.050 ;
        RECT 688.950 593.400 700.050 594.600 ;
        RECT 688.950 592.950 691.050 593.400 ;
        RECT 697.950 592.950 700.050 593.400 ;
        RECT 739.950 594.600 742.050 595.050 ;
        RECT 743.400 594.600 744.600 595.950 ;
        RECT 755.400 594.600 756.600 599.400 ;
        RECT 757.950 598.950 760.050 599.400 ;
        RECT 739.950 593.400 744.600 594.600 ;
        RECT 752.400 593.400 756.600 594.600 ;
        RECT 739.950 592.950 742.050 593.400 ;
        RECT 295.950 591.600 298.050 592.050 ;
        RECT 290.400 590.400 298.050 591.600 ;
        RECT 214.950 589.950 217.050 590.400 ;
        RECT 262.950 589.950 265.050 590.400 ;
        RECT 295.950 589.950 298.050 590.400 ;
        RECT 301.950 591.600 304.050 592.050 ;
        RECT 319.950 591.600 322.050 592.050 ;
        RECT 301.950 590.400 322.050 591.600 ;
        RECT 301.950 589.950 304.050 590.400 ;
        RECT 319.950 589.950 322.050 590.400 ;
        RECT 331.950 591.600 334.050 592.050 ;
        RECT 343.950 591.600 346.050 592.050 ;
        RECT 331.950 590.400 346.050 591.600 ;
        RECT 331.950 589.950 334.050 590.400 ;
        RECT 343.950 589.950 346.050 590.400 ;
        RECT 349.950 591.600 352.050 592.050 ;
        RECT 412.950 591.600 415.050 592.050 ;
        RECT 349.950 590.400 415.050 591.600 ;
        RECT 349.950 589.950 352.050 590.400 ;
        RECT 412.950 589.950 415.050 590.400 ;
        RECT 532.950 591.600 535.050 592.050 ;
        RECT 556.950 591.600 559.050 592.050 ;
        RECT 532.950 590.400 559.050 591.600 ;
        RECT 532.950 589.950 535.050 590.400 ;
        RECT 556.950 589.950 559.050 590.400 ;
        RECT 640.950 591.600 643.050 592.050 ;
        RECT 658.950 591.600 661.050 592.050 ;
        RECT 640.950 590.400 661.050 591.600 ;
        RECT 640.950 589.950 643.050 590.400 ;
        RECT 658.950 589.950 661.050 590.400 ;
        RECT 661.950 591.600 664.050 592.050 ;
        RECT 736.950 591.600 739.050 592.050 ;
        RECT 661.950 590.400 739.050 591.600 ;
        RECT 661.950 589.950 664.050 590.400 ;
        RECT 736.950 589.950 739.050 590.400 ;
        RECT 19.950 588.600 22.050 589.050 ;
        RECT 109.950 588.600 112.050 589.050 ;
        RECT 19.950 587.400 112.050 588.600 ;
        RECT 19.950 586.950 22.050 587.400 ;
        RECT 109.950 586.950 112.050 587.400 ;
        RECT 235.950 588.600 238.050 589.050 ;
        RECT 247.950 588.600 250.050 589.050 ;
        RECT 235.950 587.400 250.050 588.600 ;
        RECT 235.950 586.950 238.050 587.400 ;
        RECT 247.950 586.950 250.050 587.400 ;
        RECT 322.950 588.600 325.050 589.050 ;
        RECT 325.950 588.600 328.050 589.050 ;
        RECT 361.950 588.600 364.050 589.050 ;
        RECT 322.950 587.400 364.050 588.600 ;
        RECT 322.950 586.950 325.050 587.400 ;
        RECT 325.950 586.950 328.050 587.400 ;
        RECT 361.950 586.950 364.050 587.400 ;
        RECT 367.950 588.600 370.050 589.050 ;
        RECT 406.950 588.600 409.050 589.050 ;
        RECT 367.950 587.400 409.050 588.600 ;
        RECT 367.950 586.950 370.050 587.400 ;
        RECT 406.950 586.950 409.050 587.400 ;
        RECT 415.950 588.600 418.050 589.050 ;
        RECT 448.950 588.600 451.050 589.050 ;
        RECT 490.950 588.600 493.050 589.050 ;
        RECT 415.950 587.400 493.050 588.600 ;
        RECT 415.950 586.950 418.050 587.400 ;
        RECT 448.950 586.950 451.050 587.400 ;
        RECT 490.950 586.950 493.050 587.400 ;
        RECT 523.950 588.600 526.050 589.050 ;
        RECT 556.950 588.600 559.050 589.050 ;
        RECT 523.950 587.400 559.050 588.600 ;
        RECT 523.950 586.950 526.050 587.400 ;
        RECT 556.950 586.950 559.050 587.400 ;
        RECT 709.950 588.600 712.050 589.050 ;
        RECT 748.950 588.600 751.050 589.050 ;
        RECT 709.950 587.400 751.050 588.600 ;
        RECT 752.400 588.600 753.600 593.400 ;
        RECT 754.950 591.600 757.050 592.050 ;
        RECT 760.950 591.600 763.050 592.050 ;
        RECT 754.950 590.400 763.050 591.600 ;
        RECT 754.950 589.950 757.050 590.400 ;
        RECT 760.950 589.950 763.050 590.400 ;
        RECT 754.950 588.600 757.050 589.050 ;
        RECT 769.950 588.600 772.050 589.050 ;
        RECT 752.400 587.400 757.050 588.600 ;
        RECT 709.950 586.950 712.050 587.400 ;
        RECT 748.950 586.950 751.050 587.400 ;
        RECT 754.950 586.950 757.050 587.400 ;
        RECT 758.400 587.400 772.050 588.600 ;
        RECT 79.950 585.600 82.050 586.050 ;
        RECT 163.950 585.600 166.050 586.050 ;
        RECT 79.950 584.400 166.050 585.600 ;
        RECT 79.950 583.950 82.050 584.400 ;
        RECT 163.950 583.950 166.050 584.400 ;
        RECT 256.950 585.600 259.050 586.050 ;
        RECT 286.950 585.600 289.050 586.050 ;
        RECT 256.950 584.400 289.050 585.600 ;
        RECT 256.950 583.950 259.050 584.400 ;
        RECT 286.950 583.950 289.050 584.400 ;
        RECT 604.950 585.600 607.050 586.050 ;
        RECT 643.950 585.600 646.050 586.050 ;
        RECT 658.950 585.600 661.050 586.050 ;
        RECT 604.950 584.400 661.050 585.600 ;
        RECT 604.950 583.950 607.050 584.400 ;
        RECT 643.950 583.950 646.050 584.400 ;
        RECT 658.950 583.950 661.050 584.400 ;
        RECT 748.950 585.600 751.050 586.050 ;
        RECT 758.400 585.600 759.600 587.400 ;
        RECT 769.950 586.950 772.050 587.400 ;
        RECT 748.950 584.400 759.600 585.600 ;
        RECT 760.950 585.600 763.050 586.050 ;
        RECT 769.950 585.600 772.050 586.050 ;
        RECT 760.950 584.400 772.050 585.600 ;
        RECT 748.950 583.950 751.050 584.400 ;
        RECT 760.950 583.950 763.050 584.400 ;
        RECT 769.950 583.950 772.050 584.400 ;
        RECT 16.950 582.600 19.050 583.050 ;
        RECT 166.950 582.600 169.050 583.050 ;
        RECT 16.950 581.400 169.050 582.600 ;
        RECT 16.950 580.950 19.050 581.400 ;
        RECT 166.950 580.950 169.050 581.400 ;
        RECT 169.950 582.600 172.050 583.050 ;
        RECT 187.950 582.600 190.050 583.050 ;
        RECT 169.950 581.400 190.050 582.600 ;
        RECT 169.950 580.950 172.050 581.400 ;
        RECT 187.950 580.950 190.050 581.400 ;
        RECT 190.950 582.600 193.050 583.050 ;
        RECT 256.950 582.600 259.050 583.050 ;
        RECT 190.950 581.400 259.050 582.600 ;
        RECT 190.950 580.950 193.050 581.400 ;
        RECT 256.950 580.950 259.050 581.400 ;
        RECT 259.950 582.600 262.050 583.050 ;
        RECT 355.950 582.600 358.050 583.050 ;
        RECT 259.950 581.400 358.050 582.600 ;
        RECT 259.950 580.950 262.050 581.400 ;
        RECT 355.950 580.950 358.050 581.400 ;
        RECT 406.950 582.600 409.050 583.050 ;
        RECT 421.950 582.600 424.050 583.050 ;
        RECT 454.950 582.600 457.050 583.050 ;
        RECT 514.950 582.600 517.050 583.050 ;
        RECT 406.950 581.400 517.050 582.600 ;
        RECT 406.950 580.950 409.050 581.400 ;
        RECT 421.950 580.950 424.050 581.400 ;
        RECT 454.950 580.950 457.050 581.400 ;
        RECT 514.950 580.950 517.050 581.400 ;
        RECT 568.950 582.600 571.050 583.050 ;
        RECT 580.950 582.600 583.050 583.050 ;
        RECT 568.950 581.400 583.050 582.600 ;
        RECT 568.950 580.950 571.050 581.400 ;
        RECT 580.950 580.950 583.050 581.400 ;
        RECT 583.950 582.600 586.050 583.050 ;
        RECT 595.950 582.600 598.050 583.050 ;
        RECT 673.950 582.600 676.050 583.050 ;
        RECT 583.950 581.400 676.050 582.600 ;
        RECT 583.950 580.950 586.050 581.400 ;
        RECT 595.950 580.950 598.050 581.400 ;
        RECT 673.950 580.950 676.050 581.400 ;
        RECT 730.950 582.600 733.050 583.050 ;
        RECT 742.950 582.600 745.050 583.050 ;
        RECT 730.950 581.400 745.050 582.600 ;
        RECT 730.950 580.950 733.050 581.400 ;
        RECT 742.950 580.950 745.050 581.400 ;
        RECT 118.950 579.600 121.050 580.050 ;
        RECT 184.950 579.600 187.050 580.050 ;
        RECT 118.950 578.400 187.050 579.600 ;
        RECT 118.950 577.950 121.050 578.400 ;
        RECT 184.950 577.950 187.050 578.400 ;
        RECT 346.950 579.600 349.050 580.050 ;
        RECT 520.950 579.600 523.050 580.050 ;
        RECT 346.950 578.400 523.050 579.600 ;
        RECT 346.950 577.950 349.050 578.400 ;
        RECT 520.950 577.950 523.050 578.400 ;
        RECT 547.950 579.600 550.050 580.050 ;
        RECT 730.950 579.600 733.050 580.050 ;
        RECT 547.950 578.400 733.050 579.600 ;
        RECT 547.950 577.950 550.050 578.400 ;
        RECT 730.950 577.950 733.050 578.400 ;
        RECT 88.950 576.600 91.050 577.050 ;
        RECT 106.950 576.600 109.050 577.050 ;
        RECT 88.950 575.400 109.050 576.600 ;
        RECT 88.950 574.950 91.050 575.400 ;
        RECT 106.950 574.950 109.050 575.400 ;
        RECT 154.950 576.600 157.050 577.050 ;
        RECT 190.950 576.600 193.050 577.050 ;
        RECT 154.950 575.400 193.050 576.600 ;
        RECT 154.950 574.950 157.050 575.400 ;
        RECT 190.950 574.950 193.050 575.400 ;
        RECT 232.950 576.600 235.050 577.050 ;
        RECT 253.950 576.600 256.050 577.050 ;
        RECT 232.950 575.400 256.050 576.600 ;
        RECT 232.950 574.950 235.050 575.400 ;
        RECT 253.950 574.950 256.050 575.400 ;
        RECT 262.950 576.600 265.050 577.050 ;
        RECT 274.950 576.600 277.050 577.050 ;
        RECT 262.950 575.400 277.050 576.600 ;
        RECT 262.950 574.950 265.050 575.400 ;
        RECT 274.950 574.950 277.050 575.400 ;
        RECT 277.950 576.600 280.050 577.050 ;
        RECT 283.950 576.600 286.050 577.050 ;
        RECT 277.950 575.400 286.050 576.600 ;
        RECT 277.950 574.950 280.050 575.400 ;
        RECT 283.950 574.950 286.050 575.400 ;
        RECT 304.950 576.600 307.050 577.050 ;
        RECT 454.950 576.600 457.050 577.050 ;
        RECT 304.950 575.400 457.050 576.600 ;
        RECT 304.950 574.950 307.050 575.400 ;
        RECT 454.950 574.950 457.050 575.400 ;
        RECT 493.950 576.600 496.050 577.050 ;
        RECT 502.950 576.600 505.050 577.050 ;
        RECT 493.950 575.400 505.050 576.600 ;
        RECT 493.950 574.950 496.050 575.400 ;
        RECT 502.950 574.950 505.050 575.400 ;
        RECT 676.950 576.600 679.050 577.050 ;
        RECT 760.950 576.600 763.050 577.050 ;
        RECT 676.950 575.400 763.050 576.600 ;
        RECT 676.950 574.950 679.050 575.400 ;
        RECT 760.950 574.950 763.050 575.400 ;
        RECT 139.950 573.600 142.050 574.050 ;
        RECT 169.950 573.600 172.050 574.050 ;
        RECT 139.950 572.400 172.050 573.600 ;
        RECT 139.950 571.950 142.050 572.400 ;
        RECT 169.950 571.950 172.050 572.400 ;
        RECT 178.950 573.600 181.050 574.050 ;
        RECT 310.950 573.600 313.050 574.050 ;
        RECT 178.950 572.400 313.050 573.600 ;
        RECT 178.950 571.950 181.050 572.400 ;
        RECT 310.950 571.950 313.050 572.400 ;
        RECT 352.950 573.600 355.050 574.050 ;
        RECT 379.950 573.600 382.050 574.050 ;
        RECT 547.950 573.600 550.050 574.050 ;
        RECT 352.950 572.400 550.050 573.600 ;
        RECT 352.950 571.950 355.050 572.400 ;
        RECT 379.950 571.950 382.050 572.400 ;
        RECT 547.950 571.950 550.050 572.400 ;
        RECT 556.950 573.600 559.050 574.050 ;
        RECT 628.950 573.600 631.050 574.050 ;
        RECT 637.950 573.600 640.050 574.050 ;
        RECT 556.950 572.400 640.050 573.600 ;
        RECT 556.950 571.950 559.050 572.400 ;
        RECT 628.950 571.950 631.050 572.400 ;
        RECT 637.950 571.950 640.050 572.400 ;
        RECT 79.950 570.600 82.050 571.050 ;
        RECT 88.950 570.600 91.050 571.050 ;
        RECT 79.950 569.400 91.050 570.600 ;
        RECT 79.950 568.950 82.050 569.400 ;
        RECT 88.950 568.950 91.050 569.400 ;
        RECT 106.950 570.600 109.050 571.050 ;
        RECT 193.950 570.600 196.050 571.050 ;
        RECT 373.950 570.600 376.050 571.050 ;
        RECT 106.950 569.400 376.050 570.600 ;
        RECT 106.950 568.950 109.050 569.400 ;
        RECT 193.950 568.950 196.050 569.400 ;
        RECT 373.950 568.950 376.050 569.400 ;
        RECT 607.950 568.950 610.050 571.050 ;
        RECT 697.950 570.600 700.050 571.050 ;
        RECT 736.950 570.600 739.050 571.050 ;
        RECT 697.950 569.400 739.050 570.600 ;
        RECT 697.950 568.950 700.050 569.400 ;
        RECT 736.950 568.950 739.050 569.400 ;
        RECT 46.950 567.600 49.050 568.050 ;
        RECT 61.950 567.600 64.050 568.050 ;
        RECT 46.950 566.400 64.050 567.600 ;
        RECT 46.950 565.950 49.050 566.400 ;
        RECT 61.950 565.950 64.050 566.400 ;
        RECT 151.950 567.600 154.050 568.050 ;
        RECT 154.950 567.600 157.050 568.050 ;
        RECT 166.950 567.600 169.050 568.050 ;
        RECT 151.950 566.400 169.050 567.600 ;
        RECT 151.950 565.950 154.050 566.400 ;
        RECT 154.950 565.950 157.050 566.400 ;
        RECT 166.950 565.950 169.050 566.400 ;
        RECT 169.950 567.600 172.050 568.050 ;
        RECT 196.950 567.600 199.050 568.050 ;
        RECT 169.950 566.400 199.050 567.600 ;
        RECT 169.950 565.950 172.050 566.400 ;
        RECT 196.950 565.950 199.050 566.400 ;
        RECT 241.950 567.600 244.050 568.050 ;
        RECT 265.950 567.600 268.050 568.050 ;
        RECT 292.950 567.600 295.050 568.050 ;
        RECT 241.950 566.400 295.050 567.600 ;
        RECT 241.950 565.950 244.050 566.400 ;
        RECT 265.950 565.950 268.050 566.400 ;
        RECT 292.950 565.950 295.050 566.400 ;
        RECT 295.950 567.600 298.050 568.050 ;
        RECT 346.950 567.600 349.050 568.050 ;
        RECT 295.950 566.400 349.050 567.600 ;
        RECT 295.950 565.950 298.050 566.400 ;
        RECT 346.950 565.950 349.050 566.400 ;
        RECT 370.950 567.600 373.050 568.050 ;
        RECT 436.950 567.600 439.050 568.050 ;
        RECT 370.950 566.400 439.050 567.600 ;
        RECT 608.400 567.600 609.600 568.950 ;
        RECT 619.950 567.600 622.050 568.050 ;
        RECT 608.400 566.400 622.050 567.600 ;
        RECT 370.950 565.950 373.050 566.400 ;
        RECT 436.950 565.950 439.050 566.400 ;
        RECT 619.950 565.950 622.050 566.400 ;
        RECT 685.950 567.600 688.050 568.050 ;
        RECT 691.950 567.600 694.050 568.050 ;
        RECT 685.950 566.400 694.050 567.600 ;
        RECT 685.950 565.950 688.050 566.400 ;
        RECT 691.950 565.950 694.050 566.400 ;
        RECT 700.950 567.600 703.050 568.050 ;
        RECT 712.950 567.600 715.050 568.050 ;
        RECT 700.950 566.400 715.050 567.600 ;
        RECT 700.950 565.950 703.050 566.400 ;
        RECT 712.950 565.950 715.050 566.400 ;
        RECT 58.950 564.600 61.050 565.050 ;
        RECT 76.950 564.600 79.050 565.050 ;
        RECT 91.950 564.600 94.050 565.050 ;
        RECT 58.950 563.400 66.600 564.600 ;
        RECT 58.950 562.950 61.050 563.400 ;
        RECT 52.950 561.600 55.050 562.050 ;
        RECT 65.400 561.600 66.600 563.400 ;
        RECT 76.950 563.400 94.050 564.600 ;
        RECT 76.950 562.950 79.050 563.400 ;
        RECT 91.950 562.950 94.050 563.400 ;
        RECT 124.950 564.600 127.050 565.050 ;
        RECT 181.950 564.600 184.050 565.050 ;
        RECT 124.950 563.400 184.050 564.600 ;
        RECT 124.950 562.950 127.050 563.400 ;
        RECT 181.950 562.950 184.050 563.400 ;
        RECT 190.950 564.600 193.050 565.050 ;
        RECT 508.950 564.600 511.050 565.050 ;
        RECT 190.950 563.400 511.050 564.600 ;
        RECT 190.950 562.950 193.050 563.400 ;
        RECT 508.950 562.950 511.050 563.400 ;
        RECT 571.950 564.600 574.050 565.050 ;
        RECT 607.950 564.600 610.050 565.050 ;
        RECT 571.950 563.400 610.050 564.600 ;
        RECT 571.950 562.950 574.050 563.400 ;
        RECT 607.950 562.950 610.050 563.400 ;
        RECT 622.950 564.600 625.050 565.050 ;
        RECT 646.950 564.600 649.050 565.050 ;
        RECT 622.950 563.400 649.050 564.600 ;
        RECT 622.950 562.950 625.050 563.400 ;
        RECT 646.950 562.950 649.050 563.400 ;
        RECT 649.950 564.600 652.050 565.050 ;
        RECT 718.950 564.600 721.050 565.050 ;
        RECT 745.950 564.600 748.050 565.050 ;
        RECT 649.950 563.400 660.600 564.600 ;
        RECT 649.950 562.950 652.050 563.400 ;
        RECT 659.400 562.050 660.600 563.400 ;
        RECT 698.400 563.400 721.050 564.600 ;
        RECT 124.950 561.600 127.050 562.050 ;
        RECT 52.950 560.400 63.600 561.600 ;
        RECT 65.400 560.400 127.050 561.600 ;
        RECT 52.950 559.950 55.050 560.400 ;
        RECT 25.950 558.600 28.050 559.050 ;
        RECT 34.950 558.600 37.050 559.050 ;
        RECT 25.950 557.400 37.050 558.600 ;
        RECT 25.950 556.950 28.050 557.400 ;
        RECT 34.950 556.950 37.050 557.400 ;
        RECT 58.950 556.950 61.050 559.050 ;
        RECT 62.400 558.600 63.600 560.400 ;
        RECT 124.950 559.950 127.050 560.400 ;
        RECT 127.950 561.600 130.050 562.050 ;
        RECT 148.950 561.600 151.050 562.050 ;
        RECT 127.950 560.400 151.050 561.600 ;
        RECT 127.950 559.950 130.050 560.400 ;
        RECT 148.950 559.950 151.050 560.400 ;
        RECT 163.950 561.600 166.050 562.050 ;
        RECT 214.950 561.600 217.050 562.050 ;
        RECT 229.950 561.600 232.050 562.050 ;
        RECT 163.950 560.400 180.600 561.600 ;
        RECT 163.950 559.950 166.050 560.400 ;
        RECT 70.950 558.600 73.050 559.050 ;
        RECT 79.950 558.600 82.050 559.050 ;
        RECT 62.400 557.400 66.600 558.600 ;
        RECT 19.950 555.600 22.050 556.050 ;
        RECT 31.950 555.600 34.050 556.050 ;
        RECT 19.950 554.400 34.050 555.600 ;
        RECT 35.400 555.600 36.600 556.950 ;
        RECT 49.950 555.600 52.050 556.050 ;
        RECT 35.400 554.400 52.050 555.600 ;
        RECT 59.400 555.600 60.600 556.950 ;
        RECT 61.950 555.600 64.050 556.050 ;
        RECT 59.400 554.400 64.050 555.600 ;
        RECT 65.400 555.600 66.600 557.400 ;
        RECT 70.950 557.400 82.050 558.600 ;
        RECT 70.950 556.950 73.050 557.400 ;
        RECT 79.950 556.950 82.050 557.400 ;
        RECT 82.950 558.600 85.050 559.050 ;
        RECT 88.950 558.600 91.050 559.050 ;
        RECT 109.950 558.600 112.050 559.050 ;
        RECT 82.950 557.400 87.600 558.600 ;
        RECT 82.950 556.950 85.050 557.400 ;
        RECT 67.950 555.600 70.050 556.050 ;
        RECT 65.400 554.400 70.050 555.600 ;
        RECT 86.400 555.600 87.600 557.400 ;
        RECT 88.950 557.400 112.050 558.600 ;
        RECT 88.950 556.950 91.050 557.400 ;
        RECT 109.950 556.950 112.050 557.400 ;
        RECT 115.950 558.600 118.050 559.050 ;
        RECT 121.950 558.600 124.050 559.050 ;
        RECT 115.950 557.400 124.050 558.600 ;
        RECT 115.950 556.950 118.050 557.400 ;
        RECT 121.950 556.950 124.050 557.400 ;
        RECT 118.950 555.600 121.050 556.050 ;
        RECT 125.400 555.600 126.600 559.950 ;
        RECT 179.400 559.050 180.600 560.400 ;
        RECT 214.950 560.400 232.050 561.600 ;
        RECT 214.950 559.950 217.050 560.400 ;
        RECT 229.950 559.950 232.050 560.400 ;
        RECT 238.950 559.950 241.050 562.050 ;
        RECT 244.950 559.950 247.050 562.050 ;
        RECT 256.950 561.600 259.050 562.050 ;
        RECT 268.950 561.600 271.050 562.050 ;
        RECT 304.950 561.600 307.050 562.050 ;
        RECT 256.950 560.400 307.050 561.600 ;
        RECT 256.950 559.950 259.050 560.400 ;
        RECT 268.950 559.950 271.050 560.400 ;
        RECT 304.950 559.950 307.050 560.400 ;
        RECT 310.950 561.600 313.050 562.050 ;
        RECT 322.950 561.600 325.050 562.050 ;
        RECT 352.950 561.600 355.050 562.050 ;
        RECT 310.950 560.400 318.600 561.600 ;
        RECT 310.950 559.950 313.050 560.400 ;
        RECT 133.950 558.600 136.050 559.050 ;
        RECT 139.950 558.600 142.050 559.050 ;
        RECT 133.950 557.400 142.050 558.600 ;
        RECT 133.950 556.950 136.050 557.400 ;
        RECT 139.950 556.950 142.050 557.400 ;
        RECT 148.950 556.950 151.050 559.050 ;
        RECT 160.950 556.950 163.050 559.050 ;
        RECT 166.950 558.600 169.050 559.050 ;
        RECT 166.950 557.400 171.600 558.600 ;
        RECT 166.950 556.950 169.050 557.400 ;
        RECT 86.400 554.400 96.600 555.600 ;
        RECT 19.950 553.950 22.050 554.400 ;
        RECT 31.950 553.950 34.050 554.400 ;
        RECT 49.950 553.950 52.050 554.400 ;
        RECT 61.950 553.950 64.050 554.400 ;
        RECT 67.950 553.950 70.050 554.400 ;
        RECT 22.950 552.600 25.050 553.050 ;
        RECT 40.950 552.600 43.050 553.050 ;
        RECT 22.950 551.400 43.050 552.600 ;
        RECT 22.950 550.950 25.050 551.400 ;
        RECT 40.950 550.950 43.050 551.400 ;
        RECT 46.950 552.600 49.050 553.050 ;
        RECT 55.950 552.600 58.050 553.050 ;
        RECT 46.950 551.400 58.050 552.600 ;
        RECT 46.950 550.950 49.050 551.400 ;
        RECT 55.950 550.950 58.050 551.400 ;
        RECT 79.950 552.600 82.050 553.050 ;
        RECT 91.950 552.600 94.050 553.050 ;
        RECT 79.950 551.400 94.050 552.600 ;
        RECT 95.400 552.600 96.600 554.400 ;
        RECT 118.950 554.400 126.600 555.600 ;
        RECT 130.950 555.600 133.050 556.050 ;
        RECT 142.950 555.600 145.050 556.050 ;
        RECT 130.950 554.400 145.050 555.600 ;
        RECT 149.400 555.600 150.600 556.950 ;
        RECT 157.950 555.600 160.050 556.050 ;
        RECT 149.400 554.400 160.050 555.600 ;
        RECT 118.950 553.950 121.050 554.400 ;
        RECT 130.950 553.950 133.050 554.400 ;
        RECT 142.950 553.950 145.050 554.400 ;
        RECT 157.950 553.950 160.050 554.400 ;
        RECT 139.950 552.600 142.050 553.050 ;
        RECT 151.950 552.600 154.050 553.050 ;
        RECT 95.400 551.400 129.600 552.600 ;
        RECT 79.950 550.950 82.050 551.400 ;
        RECT 91.950 550.950 94.050 551.400 ;
        RECT 28.950 549.600 31.050 550.050 ;
        RECT 88.950 549.600 91.050 550.050 ;
        RECT 124.950 549.600 127.050 550.050 ;
        RECT 28.950 548.400 127.050 549.600 ;
        RECT 128.400 549.600 129.600 551.400 ;
        RECT 139.950 551.400 154.050 552.600 ;
        RECT 161.400 552.600 162.600 556.950 ;
        RECT 170.400 556.050 171.600 557.400 ;
        RECT 172.950 556.950 175.050 559.050 ;
        RECT 178.950 556.950 181.050 559.050 ;
        RECT 190.950 558.600 193.050 559.050 ;
        RECT 217.950 558.600 220.050 559.050 ;
        RECT 226.950 558.600 229.050 559.050 ;
        RECT 190.950 557.400 195.600 558.600 ;
        RECT 190.950 556.950 193.050 557.400 ;
        RECT 169.950 553.950 172.050 556.050 ;
        RECT 169.950 552.600 172.050 553.050 ;
        RECT 161.400 551.400 172.050 552.600 ;
        RECT 139.950 550.950 142.050 551.400 ;
        RECT 151.950 550.950 154.050 551.400 ;
        RECT 169.950 550.950 172.050 551.400 ;
        RECT 139.950 549.600 142.050 550.050 ;
        RECT 145.950 549.600 148.050 550.050 ;
        RECT 128.400 548.400 148.050 549.600 ;
        RECT 28.950 547.950 31.050 548.400 ;
        RECT 88.950 547.950 91.050 548.400 ;
        RECT 124.950 547.950 127.050 548.400 ;
        RECT 139.950 547.950 142.050 548.400 ;
        RECT 145.950 547.950 148.050 548.400 ;
        RECT 163.950 549.600 166.050 550.050 ;
        RECT 173.400 549.600 174.600 556.950 ;
        RECT 194.400 556.050 195.600 557.400 ;
        RECT 217.950 557.400 229.050 558.600 ;
        RECT 217.950 556.950 220.050 557.400 ;
        RECT 226.950 556.950 229.050 557.400 ;
        RECT 239.400 556.050 240.600 559.950 ;
        RECT 178.950 555.600 181.050 556.050 ;
        RECT 190.950 555.600 193.050 556.050 ;
        RECT 178.950 554.400 193.050 555.600 ;
        RECT 178.950 553.950 181.050 554.400 ;
        RECT 190.950 553.950 193.050 554.400 ;
        RECT 193.950 553.950 196.050 556.050 ;
        RECT 196.950 555.600 199.050 556.050 ;
        RECT 229.950 555.600 232.050 556.050 ;
        RECT 196.950 554.400 232.050 555.600 ;
        RECT 196.950 553.950 199.050 554.400 ;
        RECT 229.950 553.950 232.050 554.400 ;
        RECT 238.950 553.950 241.050 556.050 ;
        RECT 245.400 555.600 246.600 559.950 ;
        RECT 274.950 556.950 277.050 559.050 ;
        RECT 280.950 558.600 283.050 559.050 ;
        RECT 286.950 558.600 289.050 559.050 ;
        RECT 280.950 557.400 306.600 558.600 ;
        RECT 280.950 556.950 283.050 557.400 ;
        RECT 286.950 556.950 289.050 557.400 ;
        RECT 262.950 555.600 265.050 556.050 ;
        RECT 245.400 554.400 265.050 555.600 ;
        RECT 275.400 555.600 276.600 556.950 ;
        RECT 305.400 556.050 306.600 557.400 ;
        RECT 289.950 555.600 292.050 556.050 ;
        RECT 275.400 554.400 292.050 555.600 ;
        RECT 262.950 553.950 265.050 554.400 ;
        RECT 289.950 553.950 292.050 554.400 ;
        RECT 304.950 553.950 307.050 556.050 ;
        RECT 310.950 555.600 313.050 556.050 ;
        RECT 317.400 555.600 318.600 560.400 ;
        RECT 322.950 560.400 355.050 561.600 ;
        RECT 322.950 559.950 325.050 560.400 ;
        RECT 352.950 559.950 355.050 560.400 ;
        RECT 361.950 561.600 364.050 562.050 ;
        RECT 394.950 561.600 397.050 562.050 ;
        RECT 361.950 560.400 397.050 561.600 ;
        RECT 361.950 559.950 364.050 560.400 ;
        RECT 394.950 559.950 397.050 560.400 ;
        RECT 409.950 561.600 412.050 562.050 ;
        RECT 433.950 561.600 436.050 562.050 ;
        RECT 445.950 561.600 448.050 562.050 ;
        RECT 409.950 560.400 414.600 561.600 ;
        RECT 409.950 559.950 412.050 560.400 ;
        RECT 370.950 558.600 373.050 559.050 ;
        RECT 338.400 557.400 373.050 558.600 ;
        RECT 310.950 554.400 318.600 555.600 ;
        RECT 319.950 555.600 322.050 556.050 ;
        RECT 338.400 555.600 339.600 557.400 ;
        RECT 370.950 556.950 373.050 557.400 ;
        RECT 373.950 556.950 376.050 559.050 ;
        RECT 376.950 558.600 379.050 559.050 ;
        RECT 376.950 557.400 381.600 558.600 ;
        RECT 376.950 556.950 379.050 557.400 ;
        RECT 319.950 554.400 339.600 555.600 ;
        RECT 340.950 555.600 343.050 556.050 ;
        RECT 349.950 555.600 352.050 556.050 ;
        RECT 340.950 554.400 352.050 555.600 ;
        RECT 374.400 555.600 375.600 556.950 ;
        RECT 380.400 555.600 381.600 557.400 ;
        RECT 385.950 556.950 388.050 559.050 ;
        RECT 391.950 558.600 394.050 559.050 ;
        RECT 403.950 558.600 406.050 559.050 ;
        RECT 409.950 558.600 412.050 559.050 ;
        RECT 391.950 557.400 396.600 558.600 ;
        RECT 391.950 556.950 394.050 557.400 ;
        RECT 382.950 555.600 385.050 556.050 ;
        RECT 374.400 554.400 378.600 555.600 ;
        RECT 380.400 554.400 385.050 555.600 ;
        RECT 386.400 555.600 387.600 556.950 ;
        RECT 391.950 555.600 394.050 556.050 ;
        RECT 386.400 554.400 394.050 555.600 ;
        RECT 395.400 555.600 396.600 557.400 ;
        RECT 403.950 557.400 412.050 558.600 ;
        RECT 403.950 556.950 406.050 557.400 ;
        RECT 409.950 556.950 412.050 557.400 ;
        RECT 400.950 555.600 403.050 556.050 ;
        RECT 395.400 554.400 403.050 555.600 ;
        RECT 413.400 555.600 414.600 560.400 ;
        RECT 433.950 560.400 448.050 561.600 ;
        RECT 433.950 559.950 436.050 560.400 ;
        RECT 445.950 559.950 448.050 560.400 ;
        RECT 454.950 561.600 457.050 562.050 ;
        RECT 481.950 561.600 484.050 562.050 ;
        RECT 454.950 560.400 484.050 561.600 ;
        RECT 454.950 559.950 457.050 560.400 ;
        RECT 481.950 559.950 484.050 560.400 ;
        RECT 589.950 559.950 592.050 562.050 ;
        RECT 631.950 561.600 634.050 562.050 ;
        RECT 652.950 561.600 655.050 562.050 ;
        RECT 631.950 560.400 655.050 561.600 ;
        RECT 631.950 559.950 634.050 560.400 ;
        RECT 652.950 559.950 655.050 560.400 ;
        RECT 658.950 559.950 661.050 562.050 ;
        RECT 670.950 561.600 673.050 562.050 ;
        RECT 698.400 561.600 699.600 563.400 ;
        RECT 718.950 562.950 721.050 563.400 ;
        RECT 737.400 563.400 748.050 564.600 ;
        RECT 662.400 560.400 673.050 561.600 ;
        RECT 439.950 558.600 442.050 559.050 ;
        RECT 451.950 558.600 454.050 559.050 ;
        RECT 439.950 557.400 454.050 558.600 ;
        RECT 439.950 556.950 442.050 557.400 ;
        RECT 451.950 556.950 454.050 557.400 ;
        RECT 535.950 558.600 538.050 559.050 ;
        RECT 586.950 558.600 589.050 559.050 ;
        RECT 535.950 557.400 589.050 558.600 ;
        RECT 535.950 556.950 538.050 557.400 ;
        RECT 586.950 556.950 589.050 557.400 ;
        RECT 424.950 555.600 427.050 556.050 ;
        RECT 430.950 555.600 433.050 556.050 ;
        RECT 413.400 554.400 433.050 555.600 ;
        RECT 310.950 553.950 313.050 554.400 ;
        RECT 319.950 553.950 322.050 554.400 ;
        RECT 340.950 553.950 343.050 554.400 ;
        RECT 349.950 553.950 352.050 554.400 ;
        RECT 184.950 552.600 187.050 553.050 ;
        RECT 199.950 552.600 202.050 553.050 ;
        RECT 223.950 552.600 226.050 553.050 ;
        RECT 373.950 552.600 376.050 553.050 ;
        RECT 184.950 551.400 202.050 552.600 ;
        RECT 184.950 550.950 187.050 551.400 ;
        RECT 199.950 550.950 202.050 551.400 ;
        RECT 203.400 551.400 226.050 552.600 ;
        RECT 175.950 549.600 178.050 550.050 ;
        RECT 203.400 549.600 204.600 551.400 ;
        RECT 223.950 550.950 226.050 551.400 ;
        RECT 365.400 551.400 376.050 552.600 ;
        RECT 377.400 552.600 378.600 554.400 ;
        RECT 382.950 553.950 385.050 554.400 ;
        RECT 391.950 553.950 394.050 554.400 ;
        RECT 400.950 553.950 403.050 554.400 ;
        RECT 424.950 553.950 427.050 554.400 ;
        RECT 430.950 553.950 433.050 554.400 ;
        RECT 436.950 555.600 439.050 556.050 ;
        RECT 469.950 555.600 472.050 556.050 ;
        RECT 436.950 554.400 472.050 555.600 ;
        RECT 436.950 553.950 439.050 554.400 ;
        RECT 469.950 553.950 472.050 554.400 ;
        RECT 481.950 555.600 484.050 556.050 ;
        RECT 487.950 555.600 490.050 556.050 ;
        RECT 481.950 554.400 490.050 555.600 ;
        RECT 481.950 553.950 484.050 554.400 ;
        RECT 487.950 553.950 490.050 554.400 ;
        RECT 529.950 555.600 532.050 556.050 ;
        RECT 535.950 555.600 538.050 556.050 ;
        RECT 529.950 554.400 538.050 555.600 ;
        RECT 529.950 553.950 532.050 554.400 ;
        RECT 535.950 553.950 538.050 554.400 ;
        RECT 562.950 555.600 565.050 556.050 ;
        RECT 568.950 555.600 571.050 556.050 ;
        RECT 562.950 554.400 571.050 555.600 ;
        RECT 562.950 553.950 565.050 554.400 ;
        RECT 568.950 553.950 571.050 554.400 ;
        RECT 586.950 555.600 589.050 556.050 ;
        RECT 590.400 555.600 591.600 559.950 ;
        RECT 662.400 559.050 663.600 560.400 ;
        RECT 670.950 559.950 673.050 560.400 ;
        RECT 683.400 560.400 699.600 561.600 ;
        RECT 700.950 561.600 703.050 562.050 ;
        RECT 712.950 561.600 715.050 562.050 ;
        RECT 700.950 560.400 715.050 561.600 ;
        RECT 592.950 558.600 595.050 559.050 ;
        RECT 610.950 558.600 613.050 559.050 ;
        RECT 616.950 558.600 619.050 559.050 ;
        RECT 592.950 557.400 606.600 558.600 ;
        RECT 592.950 556.950 595.050 557.400 ;
        RECT 605.400 556.050 606.600 557.400 ;
        RECT 610.950 557.400 619.050 558.600 ;
        RECT 610.950 556.950 613.050 557.400 ;
        RECT 616.950 556.950 619.050 557.400 ;
        RECT 622.950 558.600 625.050 559.050 ;
        RECT 643.950 558.600 646.050 559.050 ;
        RECT 622.950 557.400 646.050 558.600 ;
        RECT 622.950 556.950 625.050 557.400 ;
        RECT 643.950 556.950 646.050 557.400 ;
        RECT 646.950 558.600 649.050 559.050 ;
        RECT 655.950 558.600 658.050 559.050 ;
        RECT 646.950 557.400 658.050 558.600 ;
        RECT 646.950 556.950 649.050 557.400 ;
        RECT 655.950 556.950 658.050 557.400 ;
        RECT 661.950 556.950 664.050 559.050 ;
        RECT 667.950 558.600 670.050 559.050 ;
        RECT 665.400 557.400 670.050 558.600 ;
        RECT 665.400 556.050 666.600 557.400 ;
        RECT 667.950 556.950 670.050 557.400 ;
        RECT 679.950 556.950 682.050 559.050 ;
        RECT 586.950 554.400 591.600 555.600 ;
        RECT 604.950 555.600 607.050 556.050 ;
        RECT 622.950 555.600 625.050 556.050 ;
        RECT 604.950 554.400 625.050 555.600 ;
        RECT 586.950 553.950 589.050 554.400 ;
        RECT 604.950 553.950 607.050 554.400 ;
        RECT 622.950 553.950 625.050 554.400 ;
        RECT 625.950 555.600 628.050 556.050 ;
        RECT 649.950 555.600 652.050 556.050 ;
        RECT 664.950 555.600 667.050 556.050 ;
        RECT 625.950 554.400 648.600 555.600 ;
        RECT 625.950 553.950 628.050 554.400 ;
        RECT 415.950 552.600 418.050 553.050 ;
        RECT 377.400 551.400 418.050 552.600 ;
        RECT 163.950 548.400 178.050 549.600 ;
        RECT 163.950 547.950 166.050 548.400 ;
        RECT 175.950 547.950 178.050 548.400 ;
        RECT 179.400 548.400 204.600 549.600 ;
        RECT 208.950 549.600 211.050 550.050 ;
        RECT 241.950 549.600 244.050 550.050 ;
        RECT 208.950 548.400 244.050 549.600 ;
        RECT 118.950 546.600 121.050 547.050 ;
        RECT 121.950 546.600 124.050 547.050 ;
        RECT 127.950 546.600 130.050 547.050 ;
        RECT 118.950 545.400 130.050 546.600 ;
        RECT 118.950 544.950 121.050 545.400 ;
        RECT 121.950 544.950 124.050 545.400 ;
        RECT 127.950 544.950 130.050 545.400 ;
        RECT 130.950 546.600 133.050 547.050 ;
        RECT 136.950 546.600 139.050 547.050 ;
        RECT 130.950 545.400 139.050 546.600 ;
        RECT 130.950 544.950 133.050 545.400 ;
        RECT 136.950 544.950 139.050 545.400 ;
        RECT 148.950 546.600 151.050 547.050 ;
        RECT 160.950 546.600 163.050 547.050 ;
        RECT 148.950 545.400 163.050 546.600 ;
        RECT 148.950 544.950 151.050 545.400 ;
        RECT 160.950 544.950 163.050 545.400 ;
        RECT 166.950 546.600 169.050 547.050 ;
        RECT 179.400 546.600 180.600 548.400 ;
        RECT 208.950 547.950 211.050 548.400 ;
        RECT 241.950 547.950 244.050 548.400 ;
        RECT 244.950 549.600 247.050 550.050 ;
        RECT 253.950 549.600 256.050 550.050 ;
        RECT 244.950 548.400 256.050 549.600 ;
        RECT 244.950 547.950 247.050 548.400 ;
        RECT 253.950 547.950 256.050 548.400 ;
        RECT 265.950 549.600 268.050 550.050 ;
        RECT 274.950 549.600 277.050 550.050 ;
        RECT 265.950 548.400 277.050 549.600 ;
        RECT 265.950 547.950 268.050 548.400 ;
        RECT 274.950 547.950 277.050 548.400 ;
        RECT 280.950 549.600 283.050 550.050 ;
        RECT 349.950 549.600 352.050 550.050 ;
        RECT 365.400 549.600 366.600 551.400 ;
        RECT 373.950 550.950 376.050 551.400 ;
        RECT 415.950 550.950 418.050 551.400 ;
        RECT 427.950 552.600 430.050 553.050 ;
        RECT 439.950 552.600 442.050 553.050 ;
        RECT 427.950 551.400 442.050 552.600 ;
        RECT 427.950 550.950 430.050 551.400 ;
        RECT 439.950 550.950 442.050 551.400 ;
        RECT 475.950 552.600 478.050 553.050 ;
        RECT 493.950 552.600 496.050 553.050 ;
        RECT 475.950 551.400 496.050 552.600 ;
        RECT 475.950 550.950 478.050 551.400 ;
        RECT 493.950 550.950 496.050 551.400 ;
        RECT 517.950 552.600 520.050 553.050 ;
        RECT 556.950 552.600 559.050 553.050 ;
        RECT 517.950 551.400 559.050 552.600 ;
        RECT 517.950 550.950 520.050 551.400 ;
        RECT 556.950 550.950 559.050 551.400 ;
        RECT 565.950 552.600 568.050 553.050 ;
        RECT 574.950 552.600 577.050 553.050 ;
        RECT 565.950 551.400 577.050 552.600 ;
        RECT 565.950 550.950 568.050 551.400 ;
        RECT 574.950 550.950 577.050 551.400 ;
        RECT 580.950 552.600 583.050 553.050 ;
        RECT 595.950 552.600 598.050 553.050 ;
        RECT 580.950 551.400 598.050 552.600 ;
        RECT 580.950 550.950 583.050 551.400 ;
        RECT 595.950 550.950 598.050 551.400 ;
        RECT 598.950 552.600 601.050 553.050 ;
        RECT 610.950 552.600 613.050 553.050 ;
        RECT 628.950 552.600 631.050 553.050 ;
        RECT 598.950 551.400 631.050 552.600 ;
        RECT 647.400 552.600 648.600 554.400 ;
        RECT 649.950 554.400 667.050 555.600 ;
        RECT 649.950 553.950 652.050 554.400 ;
        RECT 664.950 553.950 667.050 554.400 ;
        RECT 680.400 552.600 681.600 556.950 ;
        RECT 647.400 551.400 681.600 552.600 ;
        RECT 598.950 550.950 601.050 551.400 ;
        RECT 610.950 550.950 613.050 551.400 ;
        RECT 628.950 550.950 631.050 551.400 ;
        RECT 683.400 550.050 684.600 560.400 ;
        RECT 700.950 559.950 703.050 560.400 ;
        RECT 712.950 559.950 715.050 560.400 ;
        RECT 718.950 561.600 721.050 562.050 ;
        RECT 737.400 561.600 738.600 563.400 ;
        RECT 745.950 562.950 748.050 563.400 ;
        RECT 718.950 560.400 738.600 561.600 ;
        RECT 718.950 559.950 721.050 560.400 ;
        RECT 739.950 559.950 742.050 562.050 ;
        RECT 748.950 561.600 751.050 562.050 ;
        RECT 748.950 560.400 753.600 561.600 ;
        RECT 748.950 559.950 751.050 560.400 ;
        RECT 685.950 558.600 688.050 559.050 ;
        RECT 709.950 558.600 712.050 559.050 ;
        RECT 685.950 557.400 712.050 558.600 ;
        RECT 685.950 556.950 688.050 557.400 ;
        RECT 709.950 556.950 712.050 557.400 ;
        RECT 715.950 558.600 718.050 559.050 ;
        RECT 730.950 558.600 733.050 559.050 ;
        RECT 715.950 557.400 733.050 558.600 ;
        RECT 715.950 556.950 718.050 557.400 ;
        RECT 730.950 556.950 733.050 557.400 ;
        RECT 733.950 556.950 736.050 559.050 ;
        RECT 688.950 555.600 691.050 556.050 ;
        RECT 700.950 555.600 703.050 556.050 ;
        RECT 688.950 554.400 703.050 555.600 ;
        RECT 688.950 553.950 691.050 554.400 ;
        RECT 700.950 553.950 703.050 554.400 ;
        RECT 709.950 555.600 712.050 556.050 ;
        RECT 734.400 555.600 735.600 556.950 ;
        RECT 709.950 554.400 735.600 555.600 ;
        RECT 740.400 555.600 741.600 559.950 ;
        RECT 748.950 555.600 751.050 556.050 ;
        RECT 740.400 554.400 751.050 555.600 ;
        RECT 709.950 553.950 712.050 554.400 ;
        RECT 748.950 553.950 751.050 554.400 ;
        RECT 685.950 552.600 688.050 553.050 ;
        RECT 691.950 552.600 694.050 553.050 ;
        RECT 685.950 551.400 694.050 552.600 ;
        RECT 685.950 550.950 688.050 551.400 ;
        RECT 691.950 550.950 694.050 551.400 ;
        RECT 697.950 552.600 700.050 553.050 ;
        RECT 752.400 552.600 753.600 560.400 ;
        RECT 697.950 551.400 753.600 552.600 ;
        RECT 697.950 550.950 700.050 551.400 ;
        RECT 280.950 548.400 366.600 549.600 ;
        RECT 367.950 549.600 370.050 550.050 ;
        RECT 373.950 549.600 376.050 550.050 ;
        RECT 367.950 548.400 376.050 549.600 ;
        RECT 280.950 547.950 283.050 548.400 ;
        RECT 349.950 547.950 352.050 548.400 ;
        RECT 367.950 547.950 370.050 548.400 ;
        RECT 373.950 547.950 376.050 548.400 ;
        RECT 391.950 549.600 394.050 550.050 ;
        RECT 436.950 549.600 439.050 550.050 ;
        RECT 601.950 549.600 604.050 550.050 ;
        RECT 391.950 548.400 604.050 549.600 ;
        RECT 391.950 547.950 394.050 548.400 ;
        RECT 436.950 547.950 439.050 548.400 ;
        RECT 601.950 547.950 604.050 548.400 ;
        RECT 607.950 549.600 610.050 550.050 ;
        RECT 640.950 549.600 643.050 550.050 ;
        RECT 670.950 549.600 673.050 550.050 ;
        RECT 607.950 548.400 673.050 549.600 ;
        RECT 607.950 547.950 610.050 548.400 ;
        RECT 640.950 547.950 643.050 548.400 ;
        RECT 670.950 547.950 673.050 548.400 ;
        RECT 682.950 547.950 685.050 550.050 ;
        RECT 694.950 549.600 697.050 550.050 ;
        RECT 712.950 549.600 715.050 550.050 ;
        RECT 694.950 548.400 715.050 549.600 ;
        RECT 694.950 547.950 697.050 548.400 ;
        RECT 712.950 547.950 715.050 548.400 ;
        RECT 721.950 549.600 724.050 550.050 ;
        RECT 739.950 549.600 742.050 550.050 ;
        RECT 721.950 548.400 742.050 549.600 ;
        RECT 721.950 547.950 724.050 548.400 ;
        RECT 739.950 547.950 742.050 548.400 ;
        RECT 166.950 545.400 180.600 546.600 ;
        RECT 403.950 546.600 406.050 547.050 ;
        RECT 418.950 546.600 421.050 547.050 ;
        RECT 403.950 545.400 421.050 546.600 ;
        RECT 166.950 544.950 169.050 545.400 ;
        RECT 403.950 544.950 406.050 545.400 ;
        RECT 418.950 544.950 421.050 545.400 ;
        RECT 445.950 546.600 448.050 547.050 ;
        RECT 469.950 546.600 472.050 547.050 ;
        RECT 502.950 546.600 505.050 547.050 ;
        RECT 445.950 545.400 505.050 546.600 ;
        RECT 445.950 544.950 448.050 545.400 ;
        RECT 469.950 544.950 472.050 545.400 ;
        RECT 502.950 544.950 505.050 545.400 ;
        RECT 508.950 546.600 511.050 547.050 ;
        RECT 529.950 546.600 532.050 547.050 ;
        RECT 508.950 545.400 532.050 546.600 ;
        RECT 508.950 544.950 511.050 545.400 ;
        RECT 529.950 544.950 532.050 545.400 ;
        RECT 565.950 546.600 568.050 547.050 ;
        RECT 589.950 546.600 592.050 547.050 ;
        RECT 565.950 545.400 592.050 546.600 ;
        RECT 565.950 544.950 568.050 545.400 ;
        RECT 589.950 544.950 592.050 545.400 ;
        RECT 610.950 546.600 613.050 547.050 ;
        RECT 622.950 546.600 625.050 547.050 ;
        RECT 610.950 545.400 625.050 546.600 ;
        RECT 610.950 544.950 613.050 545.400 ;
        RECT 622.950 544.950 625.050 545.400 ;
        RECT 652.950 546.600 655.050 547.050 ;
        RECT 667.950 546.600 670.050 547.050 ;
        RECT 652.950 545.400 670.050 546.600 ;
        RECT 652.950 544.950 655.050 545.400 ;
        RECT 667.950 544.950 670.050 545.400 ;
        RECT 691.950 546.600 694.050 547.050 ;
        RECT 766.950 546.600 769.050 547.050 ;
        RECT 691.950 545.400 769.050 546.600 ;
        RECT 691.950 544.950 694.050 545.400 ;
        RECT 766.950 544.950 769.050 545.400 ;
        RECT 10.950 543.600 13.050 544.050 ;
        RECT 280.950 543.600 283.050 544.050 ;
        RECT 10.950 542.400 283.050 543.600 ;
        RECT 10.950 541.950 13.050 542.400 ;
        RECT 280.950 541.950 283.050 542.400 ;
        RECT 316.950 543.600 319.050 544.050 ;
        RECT 358.950 543.600 361.050 544.050 ;
        RECT 316.950 542.400 361.050 543.600 ;
        RECT 316.950 541.950 319.050 542.400 ;
        RECT 358.950 541.950 361.050 542.400 ;
        RECT 367.950 543.600 370.050 544.050 ;
        RECT 379.950 543.600 382.050 544.050 ;
        RECT 367.950 542.400 382.050 543.600 ;
        RECT 367.950 541.950 370.050 542.400 ;
        RECT 379.950 541.950 382.050 542.400 ;
        RECT 388.950 543.600 391.050 544.050 ;
        RECT 394.950 543.600 397.050 544.050 ;
        RECT 388.950 542.400 397.050 543.600 ;
        RECT 388.950 541.950 391.050 542.400 ;
        RECT 394.950 541.950 397.050 542.400 ;
        RECT 397.950 543.600 400.050 544.050 ;
        RECT 412.950 543.600 415.050 544.050 ;
        RECT 397.950 542.400 415.050 543.600 ;
        RECT 397.950 541.950 400.050 542.400 ;
        RECT 412.950 541.950 415.050 542.400 ;
        RECT 526.950 543.600 529.050 544.050 ;
        RECT 562.950 543.600 565.050 544.050 ;
        RECT 526.950 542.400 565.050 543.600 ;
        RECT 526.950 541.950 529.050 542.400 ;
        RECT 562.950 541.950 565.050 542.400 ;
        RECT 568.950 543.600 571.050 544.050 ;
        RECT 577.950 543.600 580.050 544.050 ;
        RECT 568.950 542.400 580.050 543.600 ;
        RECT 568.950 541.950 571.050 542.400 ;
        RECT 577.950 541.950 580.050 542.400 ;
        RECT 589.950 543.600 592.050 544.050 ;
        RECT 619.950 543.600 622.050 544.050 ;
        RECT 589.950 542.400 622.050 543.600 ;
        RECT 589.950 541.950 592.050 542.400 ;
        RECT 619.950 541.950 622.050 542.400 ;
        RECT 676.950 543.600 679.050 544.050 ;
        RECT 721.950 543.600 724.050 544.050 ;
        RECT 724.950 543.600 727.050 544.050 ;
        RECT 676.950 542.400 727.050 543.600 ;
        RECT 676.950 541.950 679.050 542.400 ;
        RECT 721.950 541.950 724.050 542.400 ;
        RECT 724.950 541.950 727.050 542.400 ;
        RECT 85.950 540.600 88.050 541.050 ;
        RECT 211.950 540.600 214.050 541.050 ;
        RECT 85.950 539.400 214.050 540.600 ;
        RECT 85.950 538.950 88.050 539.400 ;
        RECT 211.950 538.950 214.050 539.400 ;
        RECT 229.950 540.600 232.050 541.050 ;
        RECT 361.950 540.600 364.050 541.050 ;
        RECT 229.950 539.400 364.050 540.600 ;
        RECT 229.950 538.950 232.050 539.400 ;
        RECT 361.950 538.950 364.050 539.400 ;
        RECT 370.950 540.600 373.050 541.050 ;
        RECT 388.950 540.600 391.050 541.050 ;
        RECT 370.950 539.400 391.050 540.600 ;
        RECT 370.950 538.950 373.050 539.400 ;
        RECT 388.950 538.950 391.050 539.400 ;
        RECT 391.950 540.600 394.050 541.050 ;
        RECT 400.950 540.600 403.050 541.050 ;
        RECT 391.950 539.400 403.050 540.600 ;
        RECT 391.950 538.950 394.050 539.400 ;
        RECT 400.950 538.950 403.050 539.400 ;
        RECT 427.950 540.600 430.050 541.050 ;
        RECT 613.950 540.600 616.050 541.050 ;
        RECT 634.950 540.600 637.050 541.050 ;
        RECT 694.950 540.600 697.050 541.050 ;
        RECT 427.950 539.400 697.050 540.600 ;
        RECT 427.950 538.950 430.050 539.400 ;
        RECT 613.950 538.950 616.050 539.400 ;
        RECT 634.950 538.950 637.050 539.400 ;
        RECT 694.950 538.950 697.050 539.400 ;
        RECT 97.950 537.600 100.050 538.050 ;
        RECT 151.950 537.600 154.050 538.050 ;
        RECT 205.950 537.600 208.050 538.050 ;
        RECT 226.950 537.600 229.050 538.050 ;
        RECT 97.950 536.400 229.050 537.600 ;
        RECT 97.950 535.950 100.050 536.400 ;
        RECT 151.950 535.950 154.050 536.400 ;
        RECT 205.950 535.950 208.050 536.400 ;
        RECT 226.950 535.950 229.050 536.400 ;
        RECT 235.950 537.600 238.050 538.050 ;
        RECT 277.950 537.600 280.050 538.050 ;
        RECT 235.950 536.400 280.050 537.600 ;
        RECT 235.950 535.950 238.050 536.400 ;
        RECT 277.950 535.950 280.050 536.400 ;
        RECT 313.950 537.600 316.050 538.050 ;
        RECT 334.950 537.600 337.050 538.050 ;
        RECT 313.950 536.400 337.050 537.600 ;
        RECT 313.950 535.950 316.050 536.400 ;
        RECT 334.950 535.950 337.050 536.400 ;
        RECT 337.950 537.600 340.050 538.050 ;
        RECT 526.950 537.600 529.050 538.050 ;
        RECT 337.950 536.400 529.050 537.600 ;
        RECT 337.950 535.950 340.050 536.400 ;
        RECT 526.950 535.950 529.050 536.400 ;
        RECT 574.950 537.600 577.050 538.050 ;
        RECT 592.950 537.600 595.050 538.050 ;
        RECT 616.950 537.600 619.050 538.050 ;
        RECT 574.950 536.400 585.600 537.600 ;
        RECT 574.950 535.950 577.050 536.400 ;
        RECT 37.950 534.600 40.050 535.050 ;
        RECT 43.950 534.600 46.050 535.050 ;
        RECT 58.950 534.600 61.050 535.050 ;
        RECT 73.950 534.600 76.050 535.050 ;
        RECT 37.950 533.400 76.050 534.600 ;
        RECT 37.950 532.950 40.050 533.400 ;
        RECT 43.950 532.950 46.050 533.400 ;
        RECT 58.950 532.950 61.050 533.400 ;
        RECT 73.950 532.950 76.050 533.400 ;
        RECT 154.950 534.600 157.050 535.050 ;
        RECT 202.950 534.600 205.050 535.050 ;
        RECT 208.950 534.600 211.050 535.050 ;
        RECT 154.950 533.400 159.600 534.600 ;
        RECT 154.950 532.950 157.050 533.400 ;
        RECT 22.950 531.600 25.050 532.050 ;
        RECT 28.950 531.600 31.050 532.050 ;
        RECT 49.950 531.600 52.050 532.050 ;
        RECT 85.950 531.600 88.050 532.050 ;
        RECT 100.950 531.600 103.050 532.050 ;
        RECT 130.950 531.600 133.050 532.050 ;
        RECT 22.950 530.400 52.050 531.600 ;
        RECT 22.950 529.950 25.050 530.400 ;
        RECT 28.950 529.950 31.050 530.400 ;
        RECT 49.950 529.950 52.050 530.400 ;
        RECT 83.400 530.400 99.600 531.600 ;
        RECT 52.950 526.950 55.050 529.050 ;
        RECT 64.950 528.600 67.050 529.050 ;
        RECT 79.950 528.600 82.050 529.050 ;
        RECT 64.950 527.400 82.050 528.600 ;
        RECT 64.950 526.950 67.050 527.400 ;
        RECT 79.950 526.950 82.050 527.400 ;
        RECT 43.950 525.600 46.050 526.050 ;
        RECT 49.950 525.600 52.050 526.050 ;
        RECT 43.950 524.400 52.050 525.600 ;
        RECT 43.950 523.950 46.050 524.400 ;
        RECT 49.950 523.950 52.050 524.400 ;
        RECT 53.400 522.600 54.600 526.950 ;
        RECT 83.400 526.050 84.600 530.400 ;
        RECT 85.950 529.950 88.050 530.400 ;
        RECT 85.950 528.600 88.050 529.050 ;
        RECT 91.950 528.600 94.050 529.050 ;
        RECT 85.950 527.400 94.050 528.600 ;
        RECT 85.950 526.950 88.050 527.400 ;
        RECT 91.950 526.950 94.050 527.400 ;
        RECT 94.950 526.950 97.050 529.050 ;
        RECT 55.950 525.600 58.050 526.050 ;
        RECT 61.950 525.600 64.050 526.050 ;
        RECT 67.950 525.600 70.050 526.050 ;
        RECT 76.950 525.600 79.050 526.050 ;
        RECT 55.950 524.400 64.050 525.600 ;
        RECT 55.950 523.950 58.050 524.400 ;
        RECT 61.950 523.950 64.050 524.400 ;
        RECT 65.400 524.400 70.050 525.600 ;
        RECT 55.950 522.600 58.050 523.050 ;
        RECT 53.400 521.400 58.050 522.600 ;
        RECT 55.950 520.950 58.050 521.400 ;
        RECT 58.950 522.600 61.050 523.050 ;
        RECT 65.400 522.600 66.600 524.400 ;
        RECT 67.950 523.950 70.050 524.400 ;
        RECT 71.400 524.400 79.050 525.600 ;
        RECT 71.400 523.050 72.600 524.400 ;
        RECT 76.950 523.950 79.050 524.400 ;
        RECT 82.950 523.950 85.050 526.050 ;
        RECT 91.950 523.950 94.050 526.050 ;
        RECT 58.950 521.400 66.600 522.600 ;
        RECT 58.950 520.950 61.050 521.400 ;
        RECT 70.950 520.950 73.050 523.050 ;
        RECT 73.950 522.600 76.050 523.050 ;
        RECT 92.400 522.600 93.600 523.950 ;
        RECT 73.950 521.400 93.600 522.600 ;
        RECT 95.400 522.600 96.600 526.950 ;
        RECT 98.400 526.050 99.600 530.400 ;
        RECT 100.950 530.400 133.050 531.600 ;
        RECT 100.950 529.950 103.050 530.400 ;
        RECT 130.950 529.950 133.050 530.400 ;
        RECT 151.950 529.950 154.050 532.050 ;
        RECT 154.950 529.950 157.050 532.050 ;
        RECT 142.950 528.600 145.050 529.050 ;
        RECT 125.400 527.400 145.050 528.600 ;
        RECT 97.950 523.950 100.050 526.050 ;
        RECT 106.950 523.950 109.050 526.050 ;
        RECT 112.950 525.600 115.050 526.050 ;
        RECT 121.950 525.600 124.050 526.050 ;
        RECT 112.950 524.400 124.050 525.600 ;
        RECT 112.950 523.950 115.050 524.400 ;
        RECT 121.950 523.950 124.050 524.400 ;
        RECT 103.950 522.600 106.050 523.050 ;
        RECT 95.400 521.400 106.050 522.600 ;
        RECT 107.400 522.600 108.600 523.950 ;
        RECT 112.950 522.600 115.050 523.050 ;
        RECT 107.400 521.400 115.050 522.600 ;
        RECT 73.950 520.950 76.050 521.400 ;
        RECT 103.950 520.950 106.050 521.400 ;
        RECT 112.950 520.950 115.050 521.400 ;
        RECT 118.950 522.600 121.050 523.050 ;
        RECT 125.400 522.600 126.600 527.400 ;
        RECT 142.950 526.950 145.050 527.400 ;
        RECT 152.400 526.050 153.600 529.950 ;
        RECT 130.950 525.600 133.050 526.050 ;
        RECT 133.950 525.600 136.050 526.050 ;
        RECT 145.950 525.600 148.050 526.050 ;
        RECT 130.950 524.400 148.050 525.600 ;
        RECT 130.950 523.950 133.050 524.400 ;
        RECT 133.950 523.950 136.050 524.400 ;
        RECT 145.950 523.950 148.050 524.400 ;
        RECT 151.950 523.950 154.050 526.050 ;
        RECT 118.950 521.400 126.600 522.600 ;
        RECT 139.950 522.600 142.050 523.050 ;
        RECT 155.400 522.600 156.600 529.950 ;
        RECT 158.400 525.600 159.600 533.400 ;
        RECT 202.950 533.400 211.050 534.600 ;
        RECT 202.950 532.950 205.050 533.400 ;
        RECT 208.950 532.950 211.050 533.400 ;
        RECT 241.950 534.600 244.050 535.050 ;
        RECT 250.950 534.600 253.050 535.050 ;
        RECT 241.950 533.400 253.050 534.600 ;
        RECT 241.950 532.950 244.050 533.400 ;
        RECT 250.950 532.950 253.050 533.400 ;
        RECT 280.950 534.600 283.050 535.050 ;
        RECT 301.950 534.600 304.050 535.050 ;
        RECT 280.950 533.400 304.050 534.600 ;
        RECT 280.950 532.950 283.050 533.400 ;
        RECT 301.950 532.950 304.050 533.400 ;
        RECT 310.950 534.600 313.050 535.050 ;
        RECT 319.950 534.600 322.050 535.050 ;
        RECT 310.950 533.400 322.050 534.600 ;
        RECT 310.950 532.950 313.050 533.400 ;
        RECT 319.950 532.950 322.050 533.400 ;
        RECT 322.950 534.600 325.050 535.050 ;
        RECT 349.950 534.600 352.050 535.050 ;
        RECT 322.950 533.400 352.050 534.600 ;
        RECT 322.950 532.950 325.050 533.400 ;
        RECT 349.950 532.950 352.050 533.400 ;
        RECT 379.950 534.600 382.050 535.050 ;
        RECT 406.950 534.600 409.050 535.050 ;
        RECT 379.950 533.400 409.050 534.600 ;
        RECT 379.950 532.950 382.050 533.400 ;
        RECT 406.950 532.950 409.050 533.400 ;
        RECT 424.950 534.600 427.050 535.050 ;
        RECT 460.950 534.600 463.050 535.050 ;
        RECT 424.950 533.400 463.050 534.600 ;
        RECT 424.950 532.950 427.050 533.400 ;
        RECT 460.950 532.950 463.050 533.400 ;
        RECT 478.950 534.600 481.050 535.050 ;
        RECT 514.950 534.600 517.050 535.050 ;
        RECT 520.950 534.600 523.050 535.050 ;
        RECT 550.950 534.600 553.050 535.050 ;
        RECT 580.950 534.600 583.050 535.050 ;
        RECT 478.950 533.400 583.050 534.600 ;
        RECT 478.950 532.950 481.050 533.400 ;
        RECT 514.950 532.950 517.050 533.400 ;
        RECT 520.950 532.950 523.050 533.400 ;
        RECT 550.950 532.950 553.050 533.400 ;
        RECT 580.950 532.950 583.050 533.400 ;
        RECT 160.950 531.600 163.050 532.050 ;
        RECT 199.950 531.600 202.050 532.050 ;
        RECT 160.950 530.400 202.050 531.600 ;
        RECT 160.950 529.950 163.050 530.400 ;
        RECT 199.950 529.950 202.050 530.400 ;
        RECT 202.950 531.600 205.050 532.050 ;
        RECT 202.950 530.400 213.600 531.600 ;
        RECT 202.950 529.950 205.050 530.400 ;
        RECT 172.950 528.600 175.050 529.050 ;
        RECT 187.950 528.600 190.050 529.050 ;
        RECT 167.400 527.400 175.050 528.600 ;
        RECT 167.400 526.050 168.600 527.400 ;
        RECT 172.950 526.950 175.050 527.400 ;
        RECT 176.400 527.400 190.050 528.600 ;
        RECT 163.950 525.600 166.050 526.050 ;
        RECT 158.400 524.400 166.050 525.600 ;
        RECT 163.950 523.950 166.050 524.400 ;
        RECT 166.950 523.950 169.050 526.050 ;
        RECT 169.950 525.600 172.050 526.050 ;
        RECT 176.400 525.600 177.600 527.400 ;
        RECT 187.950 526.950 190.050 527.400 ;
        RECT 169.950 524.400 177.600 525.600 ;
        RECT 169.950 523.950 172.050 524.400 ;
        RECT 139.950 521.400 156.600 522.600 ;
        RECT 212.400 522.600 213.600 530.400 ;
        RECT 214.950 529.950 217.050 532.050 ;
        RECT 220.950 531.600 223.050 532.050 ;
        RECT 238.950 531.600 241.050 532.050 ;
        RECT 295.950 531.600 298.050 532.050 ;
        RECT 220.950 530.400 231.600 531.600 ;
        RECT 220.950 529.950 223.050 530.400 ;
        RECT 215.400 526.050 216.600 529.950 ;
        RECT 230.400 526.050 231.600 530.400 ;
        RECT 238.950 530.400 298.050 531.600 ;
        RECT 238.950 529.950 241.050 530.400 ;
        RECT 295.950 529.950 298.050 530.400 ;
        RECT 304.950 531.600 307.050 532.050 ;
        RECT 325.950 531.600 328.050 532.050 ;
        RECT 304.950 530.400 328.050 531.600 ;
        RECT 304.950 529.950 307.050 530.400 ;
        RECT 325.950 529.950 328.050 530.400 ;
        RECT 328.950 531.600 331.050 532.050 ;
        RECT 340.950 531.600 343.050 532.050 ;
        RECT 346.950 531.600 349.050 532.050 ;
        RECT 328.950 530.400 349.050 531.600 ;
        RECT 328.950 529.950 331.050 530.400 ;
        RECT 340.950 529.950 343.050 530.400 ;
        RECT 346.950 529.950 349.050 530.400 ;
        RECT 364.950 531.600 367.050 532.050 ;
        RECT 376.950 531.600 379.050 532.050 ;
        RECT 364.950 530.400 379.050 531.600 ;
        RECT 364.950 529.950 367.050 530.400 ;
        RECT 376.950 529.950 379.050 530.400 ;
        RECT 388.950 531.600 391.050 532.050 ;
        RECT 397.950 531.600 400.050 532.050 ;
        RECT 388.950 530.400 400.050 531.600 ;
        RECT 388.950 529.950 391.050 530.400 ;
        RECT 397.950 529.950 400.050 530.400 ;
        RECT 400.950 531.600 403.050 532.050 ;
        RECT 430.950 531.600 433.050 532.050 ;
        RECT 400.950 530.400 433.050 531.600 ;
        RECT 400.950 529.950 403.050 530.400 ;
        RECT 430.950 529.950 433.050 530.400 ;
        RECT 442.950 531.600 445.050 532.050 ;
        RECT 448.950 531.600 451.050 532.050 ;
        RECT 442.950 530.400 451.050 531.600 ;
        RECT 442.950 529.950 445.050 530.400 ;
        RECT 448.950 529.950 451.050 530.400 ;
        RECT 502.950 531.600 505.050 532.050 ;
        RECT 523.950 531.600 526.050 532.050 ;
        RECT 502.950 530.400 526.050 531.600 ;
        RECT 502.950 529.950 505.050 530.400 ;
        RECT 523.950 529.950 526.050 530.400 ;
        RECT 553.950 529.950 556.050 532.050 ;
        RECT 562.950 531.600 565.050 532.050 ;
        RECT 562.950 530.400 576.600 531.600 ;
        RECT 562.950 529.950 565.050 530.400 ;
        RECT 241.950 528.600 244.050 529.050 ;
        RECT 233.400 527.400 244.050 528.600 ;
        RECT 214.950 523.950 217.050 526.050 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 233.400 523.050 234.600 527.400 ;
        RECT 241.950 526.950 244.050 527.400 ;
        RECT 247.950 528.600 250.050 529.050 ;
        RECT 256.950 528.600 259.050 529.050 ;
        RECT 247.950 527.400 259.050 528.600 ;
        RECT 247.950 526.950 250.050 527.400 ;
        RECT 256.950 526.950 259.050 527.400 ;
        RECT 262.950 528.600 265.050 529.050 ;
        RECT 268.950 528.600 271.050 529.050 ;
        RECT 262.950 527.400 271.050 528.600 ;
        RECT 262.950 526.950 265.050 527.400 ;
        RECT 268.950 526.950 271.050 527.400 ;
        RECT 277.950 526.950 280.050 529.050 ;
        RECT 286.950 528.600 289.050 529.050 ;
        RECT 292.950 528.600 295.050 529.050 ;
        RECT 307.950 528.600 310.050 529.050 ;
        RECT 319.950 528.600 322.050 529.050 ;
        RECT 286.950 527.400 291.600 528.600 ;
        RECT 286.950 526.950 289.050 527.400 ;
        RECT 220.950 522.600 223.050 523.050 ;
        RECT 212.400 521.400 223.050 522.600 ;
        RECT 118.950 520.950 121.050 521.400 ;
        RECT 139.950 520.950 142.050 521.400 ;
        RECT 220.950 520.950 223.050 521.400 ;
        RECT 232.950 520.950 235.050 523.050 ;
        RECT 238.950 522.600 241.050 523.050 ;
        RECT 268.950 522.600 271.050 523.050 ;
        RECT 271.950 522.600 274.050 523.050 ;
        RECT 238.950 521.400 274.050 522.600 ;
        RECT 238.950 520.950 241.050 521.400 ;
        RECT 268.950 520.950 271.050 521.400 ;
        RECT 271.950 520.950 274.050 521.400 ;
        RECT 40.950 519.600 43.050 520.050 ;
        RECT 70.950 519.600 73.050 520.050 ;
        RECT 40.950 518.400 73.050 519.600 ;
        RECT 40.950 517.950 43.050 518.400 ;
        RECT 70.950 517.950 73.050 518.400 ;
        RECT 115.950 519.600 118.050 520.050 ;
        RECT 178.950 519.600 181.050 520.050 ;
        RECT 115.950 518.400 181.050 519.600 ;
        RECT 115.950 517.950 118.050 518.400 ;
        RECT 178.950 517.950 181.050 518.400 ;
        RECT 229.950 519.600 232.050 520.050 ;
        RECT 244.950 519.600 247.050 520.050 ;
        RECT 229.950 518.400 247.050 519.600 ;
        RECT 229.950 517.950 232.050 518.400 ;
        RECT 244.950 517.950 247.050 518.400 ;
        RECT 250.950 519.600 253.050 520.050 ;
        RECT 253.950 519.600 256.050 520.050 ;
        RECT 259.950 519.600 262.050 520.050 ;
        RECT 250.950 518.400 262.050 519.600 ;
        RECT 278.400 519.600 279.600 526.950 ;
        RECT 290.400 525.600 291.600 527.400 ;
        RECT 292.950 527.400 297.600 528.600 ;
        RECT 292.950 526.950 295.050 527.400 ;
        RECT 296.400 525.600 297.600 527.400 ;
        RECT 307.950 527.400 322.050 528.600 ;
        RECT 307.950 526.950 310.050 527.400 ;
        RECT 319.950 526.950 322.050 527.400 ;
        RECT 322.950 526.950 325.050 529.050 ;
        RECT 343.950 526.950 346.050 529.050 ;
        RECT 367.950 528.600 370.050 529.050 ;
        RECT 385.950 528.600 388.050 529.050 ;
        RECT 365.400 527.400 370.050 528.600 ;
        RECT 323.400 525.600 324.600 526.950 ;
        RECT 290.400 524.400 294.600 525.600 ;
        RECT 296.400 524.400 324.600 525.600 ;
        RECT 293.400 523.050 294.600 524.400 ;
        RECT 280.950 522.600 283.050 523.050 ;
        RECT 289.950 522.600 292.050 523.050 ;
        RECT 280.950 521.400 292.050 522.600 ;
        RECT 280.950 520.950 283.050 521.400 ;
        RECT 289.950 520.950 292.050 521.400 ;
        RECT 292.950 520.950 295.050 523.050 ;
        RECT 307.950 522.600 310.050 523.050 ;
        RECT 316.950 522.600 319.050 523.050 ;
        RECT 344.400 522.600 345.600 526.950 ;
        RECT 365.400 526.050 366.600 527.400 ;
        RECT 367.950 526.950 370.050 527.400 ;
        RECT 380.400 527.400 388.050 528.600 ;
        RECT 352.950 523.950 355.050 526.050 ;
        RECT 364.950 523.950 367.050 526.050 ;
        RECT 307.950 521.400 345.600 522.600 ;
        RECT 307.950 520.950 310.050 521.400 ;
        RECT 316.950 520.950 319.050 521.400 ;
        RECT 295.950 519.600 298.050 520.050 ;
        RECT 278.400 518.400 298.050 519.600 ;
        RECT 250.950 517.950 253.050 518.400 ;
        RECT 253.950 517.950 256.050 518.400 ;
        RECT 259.950 517.950 262.050 518.400 ;
        RECT 295.950 517.950 298.050 518.400 ;
        RECT 313.950 519.600 316.050 520.050 ;
        RECT 322.950 519.600 325.050 520.050 ;
        RECT 313.950 518.400 325.050 519.600 ;
        RECT 313.950 517.950 316.050 518.400 ;
        RECT 322.950 517.950 325.050 518.400 ;
        RECT 325.950 519.600 328.050 520.050 ;
        RECT 353.400 519.600 354.600 523.950 ;
        RECT 361.950 522.600 364.050 523.050 ;
        RECT 380.400 522.600 381.600 527.400 ;
        RECT 385.950 526.950 388.050 527.400 ;
        RECT 397.950 528.600 400.050 529.050 ;
        RECT 409.950 528.600 412.050 529.050 ;
        RECT 397.950 527.400 412.050 528.600 ;
        RECT 397.950 526.950 400.050 527.400 ;
        RECT 409.950 526.950 412.050 527.400 ;
        RECT 415.950 528.600 418.050 529.050 ;
        RECT 442.950 528.600 445.050 529.050 ;
        RECT 415.950 527.400 445.050 528.600 ;
        RECT 415.950 526.950 418.050 527.400 ;
        RECT 442.950 526.950 445.050 527.400 ;
        RECT 449.400 526.050 450.600 529.950 ;
        RECT 454.950 526.950 457.050 529.050 ;
        RECT 469.950 528.600 472.050 529.050 ;
        RECT 458.400 527.400 472.050 528.600 ;
        RECT 421.950 523.950 424.050 526.050 ;
        RECT 448.950 523.950 451.050 526.050 ;
        RECT 422.400 522.600 423.600 523.950 ;
        RECT 427.950 522.600 430.050 523.050 ;
        RECT 361.950 521.400 411.600 522.600 ;
        RECT 422.400 521.400 430.050 522.600 ;
        RECT 361.950 520.950 364.050 521.400 ;
        RECT 325.950 518.400 354.600 519.600 ;
        RECT 367.950 519.600 370.050 520.050 ;
        RECT 403.950 519.600 406.050 520.050 ;
        RECT 367.950 518.400 406.050 519.600 ;
        RECT 410.400 519.600 411.600 521.400 ;
        RECT 427.950 520.950 430.050 521.400 ;
        RECT 445.950 522.600 448.050 523.050 ;
        RECT 455.400 522.600 456.600 526.950 ;
        RECT 458.400 526.050 459.600 527.400 ;
        RECT 469.950 526.950 472.050 527.400 ;
        RECT 511.950 528.600 514.050 529.050 ;
        RECT 517.950 528.600 520.050 529.050 ;
        RECT 541.950 528.600 544.050 529.050 ;
        RECT 511.950 527.400 520.050 528.600 ;
        RECT 511.950 526.950 514.050 527.400 ;
        RECT 517.950 526.950 520.050 527.400 ;
        RECT 521.400 527.400 544.050 528.600 ;
        RECT 554.400 528.600 555.600 529.950 ;
        RECT 575.400 529.050 576.600 530.400 ;
        RECT 584.400 529.050 585.600 536.400 ;
        RECT 592.950 536.400 619.050 537.600 ;
        RECT 592.950 535.950 595.050 536.400 ;
        RECT 616.950 535.950 619.050 536.400 ;
        RECT 619.950 537.600 622.050 538.050 ;
        RECT 697.950 537.600 700.050 538.050 ;
        RECT 619.950 536.400 700.050 537.600 ;
        RECT 619.950 535.950 622.050 536.400 ;
        RECT 697.950 535.950 700.050 536.400 ;
        RECT 739.950 537.600 742.050 538.050 ;
        RECT 754.950 537.600 757.050 538.050 ;
        RECT 739.950 536.400 757.050 537.600 ;
        RECT 739.950 535.950 742.050 536.400 ;
        RECT 754.950 535.950 757.050 536.400 ;
        RECT 586.950 534.600 589.050 535.050 ;
        RECT 610.950 534.600 613.050 535.050 ;
        RECT 586.950 533.400 613.050 534.600 ;
        RECT 586.950 532.950 589.050 533.400 ;
        RECT 610.950 532.950 613.050 533.400 ;
        RECT 697.950 534.600 700.050 535.050 ;
        RECT 742.950 534.600 745.050 535.050 ;
        RECT 697.950 533.400 745.050 534.600 ;
        RECT 697.950 532.950 700.050 533.400 ;
        RECT 742.950 532.950 745.050 533.400 ;
        RECT 601.950 531.600 604.050 532.050 ;
        RECT 703.950 531.600 706.050 532.050 ;
        RECT 709.950 531.600 712.050 532.050 ;
        RECT 601.950 530.400 712.050 531.600 ;
        RECT 601.950 529.950 604.050 530.400 ;
        RECT 703.950 529.950 706.050 530.400 ;
        RECT 709.950 529.950 712.050 530.400 ;
        RECT 730.950 531.600 733.050 532.050 ;
        RECT 742.950 531.600 745.050 532.050 ;
        RECT 730.950 530.400 745.050 531.600 ;
        RECT 730.950 529.950 733.050 530.400 ;
        RECT 742.950 529.950 745.050 530.400 ;
        RECT 562.950 528.600 565.050 529.050 ;
        RECT 554.400 527.400 565.050 528.600 ;
        RECT 521.400 526.050 522.600 527.400 ;
        RECT 541.950 526.950 544.050 527.400 ;
        RECT 562.950 526.950 565.050 527.400 ;
        RECT 574.950 526.950 577.050 529.050 ;
        RECT 583.950 528.600 586.050 529.050 ;
        RECT 601.950 528.600 604.050 529.050 ;
        RECT 583.950 527.400 604.050 528.600 ;
        RECT 583.950 526.950 586.050 527.400 ;
        RECT 601.950 526.950 604.050 527.400 ;
        RECT 619.950 528.600 622.050 529.050 ;
        RECT 628.950 528.600 631.050 529.050 ;
        RECT 619.950 527.400 631.050 528.600 ;
        RECT 619.950 526.950 622.050 527.400 ;
        RECT 628.950 526.950 631.050 527.400 ;
        RECT 634.950 528.600 637.050 529.050 ;
        RECT 643.950 528.600 646.050 529.050 ;
        RECT 634.950 527.400 646.050 528.600 ;
        RECT 634.950 526.950 637.050 527.400 ;
        RECT 643.950 526.950 646.050 527.400 ;
        RECT 664.950 526.950 667.050 529.050 ;
        RECT 694.950 528.600 697.050 529.050 ;
        RECT 715.950 528.600 718.050 529.050 ;
        RECT 724.950 528.600 727.050 529.050 ;
        RECT 760.950 528.600 763.050 529.050 ;
        RECT 694.950 527.400 727.050 528.600 ;
        RECT 694.950 526.950 697.050 527.400 ;
        RECT 715.950 526.950 718.050 527.400 ;
        RECT 724.950 526.950 727.050 527.400 ;
        RECT 758.400 527.400 763.050 528.600 ;
        RECT 457.950 523.950 460.050 526.050 ;
        RECT 463.950 525.600 466.050 526.050 ;
        RECT 472.950 525.600 475.050 526.050 ;
        RECT 463.950 524.400 475.050 525.600 ;
        RECT 463.950 523.950 466.050 524.400 ;
        RECT 472.950 523.950 475.050 524.400 ;
        RECT 520.950 523.950 523.050 526.050 ;
        RECT 526.950 525.600 529.050 526.050 ;
        RECT 535.950 525.600 538.050 526.050 ;
        RECT 526.950 524.400 538.050 525.600 ;
        RECT 526.950 523.950 529.050 524.400 ;
        RECT 535.950 523.950 538.050 524.400 ;
        RECT 541.950 525.600 544.050 526.050 ;
        RECT 613.950 525.600 616.050 526.050 ;
        RECT 634.950 525.600 637.050 526.050 ;
        RECT 541.950 524.400 637.050 525.600 ;
        RECT 541.950 523.950 544.050 524.400 ;
        RECT 613.950 523.950 616.050 524.400 ;
        RECT 634.950 523.950 637.050 524.400 ;
        RECT 649.950 525.600 652.050 526.050 ;
        RECT 655.950 525.600 658.050 526.050 ;
        RECT 649.950 524.400 658.050 525.600 ;
        RECT 649.950 523.950 652.050 524.400 ;
        RECT 655.950 523.950 658.050 524.400 ;
        RECT 445.950 521.400 456.600 522.600 ;
        RECT 460.950 522.600 463.050 523.050 ;
        RECT 484.950 522.600 487.050 523.050 ;
        RECT 502.950 522.600 505.050 523.050 ;
        RECT 460.950 521.400 505.050 522.600 ;
        RECT 445.950 520.950 448.050 521.400 ;
        RECT 460.950 520.950 463.050 521.400 ;
        RECT 484.950 520.950 487.050 521.400 ;
        RECT 502.950 520.950 505.050 521.400 ;
        RECT 505.950 522.600 508.050 523.050 ;
        RECT 520.950 522.600 523.050 523.050 ;
        RECT 505.950 521.400 523.050 522.600 ;
        RECT 505.950 520.950 508.050 521.400 ;
        RECT 520.950 520.950 523.050 521.400 ;
        RECT 523.950 522.600 526.050 523.050 ;
        RECT 529.950 522.600 532.050 523.050 ;
        RECT 523.950 521.400 532.050 522.600 ;
        RECT 523.950 520.950 526.050 521.400 ;
        RECT 529.950 520.950 532.050 521.400 ;
        RECT 562.950 522.600 565.050 523.050 ;
        RECT 574.950 522.600 577.050 523.050 ;
        RECT 562.950 521.400 577.050 522.600 ;
        RECT 562.950 520.950 565.050 521.400 ;
        RECT 574.950 520.950 577.050 521.400 ;
        RECT 586.950 522.600 589.050 523.050 ;
        RECT 595.950 522.600 598.050 523.050 ;
        RECT 586.950 521.400 598.050 522.600 ;
        RECT 586.950 520.950 589.050 521.400 ;
        RECT 595.950 520.950 598.050 521.400 ;
        RECT 601.950 522.600 604.050 523.050 ;
        RECT 613.950 522.600 616.050 523.050 ;
        RECT 601.950 521.400 616.050 522.600 ;
        RECT 601.950 520.950 604.050 521.400 ;
        RECT 613.950 520.950 616.050 521.400 ;
        RECT 658.950 522.600 661.050 523.050 ;
        RECT 665.400 522.600 666.600 526.950 ;
        RECT 667.950 523.950 670.050 526.050 ;
        RECT 673.950 525.600 676.050 526.050 ;
        RECT 679.950 525.600 682.050 526.050 ;
        RECT 673.950 524.400 682.050 525.600 ;
        RECT 673.950 523.950 676.050 524.400 ;
        RECT 679.950 523.950 682.050 524.400 ;
        RECT 709.950 525.600 712.050 526.050 ;
        RECT 736.950 525.600 739.050 526.050 ;
        RECT 709.950 524.400 739.050 525.600 ;
        RECT 709.950 523.950 712.050 524.400 ;
        RECT 736.950 523.950 739.050 524.400 ;
        RECT 745.950 525.600 748.050 526.050 ;
        RECT 758.400 525.600 759.600 527.400 ;
        RECT 760.950 526.950 763.050 527.400 ;
        RECT 745.950 524.400 759.600 525.600 ;
        RECT 745.950 523.950 748.050 524.400 ;
        RECT 658.950 521.400 666.600 522.600 ;
        RECT 668.400 522.600 669.600 523.950 ;
        RECT 679.950 522.600 682.050 523.050 ;
        RECT 721.950 522.600 724.050 523.050 ;
        RECT 668.400 521.400 724.050 522.600 ;
        RECT 658.950 520.950 661.050 521.400 ;
        RECT 679.950 520.950 682.050 521.400 ;
        RECT 721.950 520.950 724.050 521.400 ;
        RECT 745.950 522.600 748.050 523.050 ;
        RECT 751.950 522.600 754.050 523.050 ;
        RECT 745.950 521.400 754.050 522.600 ;
        RECT 745.950 520.950 748.050 521.400 ;
        RECT 751.950 520.950 754.050 521.400 ;
        RECT 433.950 519.600 436.050 520.050 ;
        RECT 445.950 519.600 448.050 520.050 ;
        RECT 410.400 518.400 448.050 519.600 ;
        RECT 325.950 517.950 328.050 518.400 ;
        RECT 367.950 517.950 370.050 518.400 ;
        RECT 403.950 517.950 406.050 518.400 ;
        RECT 433.950 517.950 436.050 518.400 ;
        RECT 445.950 517.950 448.050 518.400 ;
        RECT 448.950 519.600 451.050 520.050 ;
        RECT 454.950 519.600 457.050 520.050 ;
        RECT 448.950 518.400 457.050 519.600 ;
        RECT 448.950 517.950 451.050 518.400 ;
        RECT 454.950 517.950 457.050 518.400 ;
        RECT 472.950 519.600 475.050 520.050 ;
        RECT 490.950 519.600 493.050 520.050 ;
        RECT 472.950 518.400 493.050 519.600 ;
        RECT 472.950 517.950 475.050 518.400 ;
        RECT 490.950 517.950 493.050 518.400 ;
        RECT 574.950 519.600 577.050 520.050 ;
        RECT 604.950 519.600 607.050 520.050 ;
        RECT 610.950 519.600 613.050 520.050 ;
        RECT 625.950 519.600 628.050 520.050 ;
        RECT 574.950 518.400 628.050 519.600 ;
        RECT 574.950 517.950 577.050 518.400 ;
        RECT 604.950 517.950 607.050 518.400 ;
        RECT 610.950 517.950 613.050 518.400 ;
        RECT 625.950 517.950 628.050 518.400 ;
        RECT 652.950 519.600 655.050 520.050 ;
        RECT 661.950 519.600 664.050 520.050 ;
        RECT 652.950 518.400 664.050 519.600 ;
        RECT 652.950 517.950 655.050 518.400 ;
        RECT 661.950 517.950 664.050 518.400 ;
        RECT 703.950 519.600 706.050 520.050 ;
        RECT 733.950 519.600 736.050 520.050 ;
        RECT 703.950 518.400 736.050 519.600 ;
        RECT 703.950 517.950 706.050 518.400 ;
        RECT 733.950 517.950 736.050 518.400 ;
        RECT 751.950 519.600 754.050 520.050 ;
        RECT 769.950 519.600 772.050 520.050 ;
        RECT 751.950 518.400 772.050 519.600 ;
        RECT 751.950 517.950 754.050 518.400 ;
        RECT 769.950 517.950 772.050 518.400 ;
        RECT 31.950 516.600 34.050 517.050 ;
        RECT 40.950 516.600 43.050 517.050 ;
        RECT 61.950 516.600 64.050 517.050 ;
        RECT 31.950 515.400 64.050 516.600 ;
        RECT 31.950 514.950 34.050 515.400 ;
        RECT 40.950 514.950 43.050 515.400 ;
        RECT 61.950 514.950 64.050 515.400 ;
        RECT 64.950 516.600 67.050 517.050 ;
        RECT 118.950 516.600 121.050 517.050 ;
        RECT 64.950 515.400 121.050 516.600 ;
        RECT 64.950 514.950 67.050 515.400 ;
        RECT 118.950 514.950 121.050 515.400 ;
        RECT 220.950 516.600 223.050 517.050 ;
        RECT 238.950 516.600 241.050 517.050 ;
        RECT 220.950 515.400 241.050 516.600 ;
        RECT 220.950 514.950 223.050 515.400 ;
        RECT 238.950 514.950 241.050 515.400 ;
        RECT 244.950 516.600 247.050 517.050 ;
        RECT 304.950 516.600 307.050 517.050 ;
        RECT 244.950 515.400 307.050 516.600 ;
        RECT 244.950 514.950 247.050 515.400 ;
        RECT 304.950 514.950 307.050 515.400 ;
        RECT 310.950 516.600 313.050 517.050 ;
        RECT 316.950 516.600 319.050 517.050 ;
        RECT 310.950 515.400 319.050 516.600 ;
        RECT 310.950 514.950 313.050 515.400 ;
        RECT 316.950 514.950 319.050 515.400 ;
        RECT 319.950 516.600 322.050 517.050 ;
        RECT 355.950 516.600 358.050 517.050 ;
        RECT 442.950 516.600 445.050 517.050 ;
        RECT 319.950 515.400 445.050 516.600 ;
        RECT 319.950 514.950 322.050 515.400 ;
        RECT 355.950 514.950 358.050 515.400 ;
        RECT 442.950 514.950 445.050 515.400 ;
        RECT 451.950 516.600 454.050 517.050 ;
        RECT 478.950 516.600 481.050 517.050 ;
        RECT 451.950 515.400 481.050 516.600 ;
        RECT 451.950 514.950 454.050 515.400 ;
        RECT 478.950 514.950 481.050 515.400 ;
        RECT 481.950 516.600 484.050 517.050 ;
        RECT 490.950 516.600 493.050 517.050 ;
        RECT 481.950 515.400 493.050 516.600 ;
        RECT 481.950 514.950 484.050 515.400 ;
        RECT 490.950 514.950 493.050 515.400 ;
        RECT 505.950 516.600 508.050 517.050 ;
        RECT 547.950 516.600 550.050 517.050 ;
        RECT 505.950 515.400 550.050 516.600 ;
        RECT 505.950 514.950 508.050 515.400 ;
        RECT 547.950 514.950 550.050 515.400 ;
        RECT 568.950 516.600 571.050 517.050 ;
        RECT 616.950 516.600 619.050 517.050 ;
        RECT 568.950 515.400 619.050 516.600 ;
        RECT 568.950 514.950 571.050 515.400 ;
        RECT 616.950 514.950 619.050 515.400 ;
        RECT 625.950 516.600 628.050 517.050 ;
        RECT 664.950 516.600 667.050 517.050 ;
        RECT 625.950 515.400 667.050 516.600 ;
        RECT 625.950 514.950 628.050 515.400 ;
        RECT 664.950 514.950 667.050 515.400 ;
        RECT 733.950 516.600 736.050 517.050 ;
        RECT 763.950 516.600 766.050 517.050 ;
        RECT 733.950 515.400 766.050 516.600 ;
        RECT 733.950 514.950 736.050 515.400 ;
        RECT 763.950 514.950 766.050 515.400 ;
        RECT 58.950 513.600 61.050 514.050 ;
        RECT 109.950 513.600 112.050 514.050 ;
        RECT 58.950 512.400 112.050 513.600 ;
        RECT 58.950 511.950 61.050 512.400 ;
        RECT 109.950 511.950 112.050 512.400 ;
        RECT 130.950 513.600 133.050 514.050 ;
        RECT 220.950 513.600 223.050 514.050 ;
        RECT 130.950 512.400 223.050 513.600 ;
        RECT 130.950 511.950 133.050 512.400 ;
        RECT 220.950 511.950 223.050 512.400 ;
        RECT 301.950 513.600 304.050 514.050 ;
        RECT 337.950 513.600 340.050 514.050 ;
        RECT 301.950 512.400 340.050 513.600 ;
        RECT 301.950 511.950 304.050 512.400 ;
        RECT 337.950 511.950 340.050 512.400 ;
        RECT 358.950 513.600 361.050 514.050 ;
        RECT 412.950 513.600 415.050 514.050 ;
        RECT 358.950 512.400 415.050 513.600 ;
        RECT 358.950 511.950 361.050 512.400 ;
        RECT 412.950 511.950 415.050 512.400 ;
        RECT 457.950 513.600 460.050 514.050 ;
        RECT 475.950 513.600 478.050 514.050 ;
        RECT 457.950 512.400 478.050 513.600 ;
        RECT 457.950 511.950 460.050 512.400 ;
        RECT 475.950 511.950 478.050 512.400 ;
        RECT 502.950 513.600 505.050 514.050 ;
        RECT 532.950 513.600 535.050 514.050 ;
        RECT 502.950 512.400 535.050 513.600 ;
        RECT 502.950 511.950 505.050 512.400 ;
        RECT 532.950 511.950 535.050 512.400 ;
        RECT 535.950 513.600 538.050 514.050 ;
        RECT 559.950 513.600 562.050 514.050 ;
        RECT 535.950 512.400 562.050 513.600 ;
        RECT 535.950 511.950 538.050 512.400 ;
        RECT 559.950 511.950 562.050 512.400 ;
        RECT 601.950 513.600 604.050 514.050 ;
        RECT 709.950 513.600 712.050 514.050 ;
        RECT 601.950 512.400 712.050 513.600 ;
        RECT 601.950 511.950 604.050 512.400 ;
        RECT 709.950 511.950 712.050 512.400 ;
        RECT 724.950 513.600 727.050 514.050 ;
        RECT 757.950 513.600 760.050 514.050 ;
        RECT 724.950 512.400 760.050 513.600 ;
        RECT 724.950 511.950 727.050 512.400 ;
        RECT 757.950 511.950 760.050 512.400 ;
        RECT 241.950 510.600 244.050 511.050 ;
        RECT 265.950 510.600 268.050 511.050 ;
        RECT 241.950 509.400 268.050 510.600 ;
        RECT 241.950 508.950 244.050 509.400 ;
        RECT 265.950 508.950 268.050 509.400 ;
        RECT 268.950 510.600 271.050 511.050 ;
        RECT 472.950 510.600 475.050 511.050 ;
        RECT 268.950 509.400 475.050 510.600 ;
        RECT 268.950 508.950 271.050 509.400 ;
        RECT 472.950 508.950 475.050 509.400 ;
        RECT 478.950 510.600 481.050 511.050 ;
        RECT 493.950 510.600 496.050 511.050 ;
        RECT 478.950 509.400 496.050 510.600 ;
        RECT 478.950 508.950 481.050 509.400 ;
        RECT 493.950 508.950 496.050 509.400 ;
        RECT 529.950 510.600 532.050 511.050 ;
        RECT 607.950 510.600 610.050 511.050 ;
        RECT 529.950 509.400 610.050 510.600 ;
        RECT 529.950 508.950 532.050 509.400 ;
        RECT 607.950 508.950 610.050 509.400 ;
        RECT 613.950 510.600 616.050 511.050 ;
        RECT 652.950 510.600 655.050 511.050 ;
        RECT 670.950 510.600 673.050 511.050 ;
        RECT 613.950 509.400 673.050 510.600 ;
        RECT 613.950 508.950 616.050 509.400 ;
        RECT 652.950 508.950 655.050 509.400 ;
        RECT 670.950 508.950 673.050 509.400 ;
        RECT 160.950 507.600 163.050 508.050 ;
        RECT 184.950 507.600 187.050 508.050 ;
        RECT 223.950 507.600 226.050 508.050 ;
        RECT 301.950 507.600 304.050 508.050 ;
        RECT 160.950 506.400 304.050 507.600 ;
        RECT 160.950 505.950 163.050 506.400 ;
        RECT 184.950 505.950 187.050 506.400 ;
        RECT 223.950 505.950 226.050 506.400 ;
        RECT 301.950 505.950 304.050 506.400 ;
        RECT 391.950 507.600 394.050 508.050 ;
        RECT 427.950 507.600 430.050 508.050 ;
        RECT 469.950 507.600 472.050 508.050 ;
        RECT 391.950 506.400 426.600 507.600 ;
        RECT 391.950 505.950 394.050 506.400 ;
        RECT 16.950 504.600 19.050 505.050 ;
        RECT 265.950 504.600 268.050 505.050 ;
        RECT 16.950 503.400 268.050 504.600 ;
        RECT 16.950 502.950 19.050 503.400 ;
        RECT 265.950 502.950 268.050 503.400 ;
        RECT 274.950 504.600 277.050 505.050 ;
        RECT 301.950 504.600 304.050 505.050 ;
        RECT 274.950 503.400 304.050 504.600 ;
        RECT 274.950 502.950 277.050 503.400 ;
        RECT 301.950 502.950 304.050 503.400 ;
        RECT 322.950 504.600 325.050 505.050 ;
        RECT 346.950 504.600 349.050 505.050 ;
        RECT 322.950 503.400 349.050 504.600 ;
        RECT 425.400 504.600 426.600 506.400 ;
        RECT 427.950 506.400 472.050 507.600 ;
        RECT 427.950 505.950 430.050 506.400 ;
        RECT 469.950 505.950 472.050 506.400 ;
        RECT 520.950 507.600 523.050 508.050 ;
        RECT 568.950 507.600 571.050 508.050 ;
        RECT 520.950 506.400 571.050 507.600 ;
        RECT 520.950 505.950 523.050 506.400 ;
        RECT 568.950 505.950 571.050 506.400 ;
        RECT 535.950 504.600 538.050 505.050 ;
        RECT 425.400 503.400 538.050 504.600 ;
        RECT 322.950 502.950 325.050 503.400 ;
        RECT 346.950 502.950 349.050 503.400 ;
        RECT 535.950 502.950 538.050 503.400 ;
        RECT 538.950 504.600 541.050 505.050 ;
        RECT 607.950 504.600 610.050 505.050 ;
        RECT 538.950 503.400 610.050 504.600 ;
        RECT 538.950 502.950 541.050 503.400 ;
        RECT 607.950 502.950 610.050 503.400 ;
        RECT 88.950 501.600 91.050 502.050 ;
        RECT 142.950 501.600 145.050 502.050 ;
        RECT 199.950 501.600 202.050 502.050 ;
        RECT 88.950 500.400 202.050 501.600 ;
        RECT 88.950 499.950 91.050 500.400 ;
        RECT 142.950 499.950 145.050 500.400 ;
        RECT 199.950 499.950 202.050 500.400 ;
        RECT 277.950 501.600 280.050 502.050 ;
        RECT 364.950 501.600 367.050 502.050 ;
        RECT 277.950 500.400 367.050 501.600 ;
        RECT 277.950 499.950 280.050 500.400 ;
        RECT 364.950 499.950 367.050 500.400 ;
        RECT 388.950 501.600 391.050 502.050 ;
        RECT 436.950 501.600 439.050 502.050 ;
        RECT 388.950 500.400 439.050 501.600 ;
        RECT 388.950 499.950 391.050 500.400 ;
        RECT 436.950 499.950 439.050 500.400 ;
        RECT 454.950 501.600 457.050 502.050 ;
        RECT 553.950 501.600 556.050 502.050 ;
        RECT 676.950 501.600 679.050 502.050 ;
        RECT 454.950 500.400 679.050 501.600 ;
        RECT 454.950 499.950 457.050 500.400 ;
        RECT 553.950 499.950 556.050 500.400 ;
        RECT 676.950 499.950 679.050 500.400 ;
        RECT 46.950 498.600 49.050 499.050 ;
        RECT 58.950 498.600 61.050 499.050 ;
        RECT 46.950 497.400 61.050 498.600 ;
        RECT 46.950 496.950 49.050 497.400 ;
        RECT 58.950 496.950 61.050 497.400 ;
        RECT 61.950 498.600 64.050 499.050 ;
        RECT 76.950 498.600 79.050 499.050 ;
        RECT 61.950 497.400 79.050 498.600 ;
        RECT 61.950 496.950 64.050 497.400 ;
        RECT 76.950 496.950 79.050 497.400 ;
        RECT 175.950 498.600 178.050 499.050 ;
        RECT 271.950 498.600 274.050 499.050 ;
        RECT 346.950 498.600 349.050 499.050 ;
        RECT 175.950 497.400 349.050 498.600 ;
        RECT 175.950 496.950 178.050 497.400 ;
        RECT 271.950 496.950 274.050 497.400 ;
        RECT 346.950 496.950 349.050 497.400 ;
        RECT 355.950 498.600 358.050 499.050 ;
        RECT 370.950 498.600 373.050 499.050 ;
        RECT 355.950 497.400 373.050 498.600 ;
        RECT 355.950 496.950 358.050 497.400 ;
        RECT 370.950 496.950 373.050 497.400 ;
        RECT 409.950 498.600 412.050 499.050 ;
        RECT 529.950 498.600 532.050 499.050 ;
        RECT 409.950 497.400 532.050 498.600 ;
        RECT 409.950 496.950 412.050 497.400 ;
        RECT 529.950 496.950 532.050 497.400 ;
        RECT 532.950 498.600 535.050 499.050 ;
        RECT 556.950 498.600 559.050 499.050 ;
        RECT 532.950 497.400 559.050 498.600 ;
        RECT 532.950 496.950 535.050 497.400 ;
        RECT 556.950 496.950 559.050 497.400 ;
        RECT 562.950 498.600 565.050 499.050 ;
        RECT 598.950 498.600 601.050 499.050 ;
        RECT 562.950 497.400 601.050 498.600 ;
        RECT 562.950 496.950 565.050 497.400 ;
        RECT 598.950 496.950 601.050 497.400 ;
        RECT 625.950 498.600 628.050 499.050 ;
        RECT 769.950 498.600 772.050 499.050 ;
        RECT 625.950 497.400 772.050 498.600 ;
        RECT 625.950 496.950 628.050 497.400 ;
        RECT 769.950 496.950 772.050 497.400 ;
        RECT 13.950 495.600 16.050 496.050 ;
        RECT 19.950 495.600 22.050 496.050 ;
        RECT 13.950 494.400 22.050 495.600 ;
        RECT 13.950 493.950 16.050 494.400 ;
        RECT 19.950 493.950 22.050 494.400 ;
        RECT 55.950 495.600 58.050 496.050 ;
        RECT 61.950 495.600 64.050 496.050 ;
        RECT 103.950 495.600 106.050 496.050 ;
        RECT 55.950 494.400 106.050 495.600 ;
        RECT 55.950 493.950 58.050 494.400 ;
        RECT 61.950 493.950 64.050 494.400 ;
        RECT 103.950 493.950 106.050 494.400 ;
        RECT 205.950 495.600 208.050 496.050 ;
        RECT 292.950 495.600 295.050 496.050 ;
        RECT 205.950 494.400 295.050 495.600 ;
        RECT 205.950 493.950 208.050 494.400 ;
        RECT 292.950 493.950 295.050 494.400 ;
        RECT 295.950 495.600 298.050 496.050 ;
        RECT 340.950 495.600 343.050 496.050 ;
        RECT 295.950 494.400 343.050 495.600 ;
        RECT 295.950 493.950 298.050 494.400 ;
        RECT 340.950 493.950 343.050 494.400 ;
        RECT 364.950 495.600 367.050 496.050 ;
        RECT 382.950 495.600 385.050 496.050 ;
        RECT 364.950 494.400 385.050 495.600 ;
        RECT 364.950 493.950 367.050 494.400 ;
        RECT 382.950 493.950 385.050 494.400 ;
        RECT 400.950 495.600 403.050 496.050 ;
        RECT 415.950 495.600 418.050 496.050 ;
        RECT 400.950 494.400 418.050 495.600 ;
        RECT 400.950 493.950 403.050 494.400 ;
        RECT 415.950 493.950 418.050 494.400 ;
        RECT 421.950 495.600 424.050 496.050 ;
        RECT 448.950 495.600 451.050 496.050 ;
        RECT 421.950 494.400 451.050 495.600 ;
        RECT 421.950 493.950 424.050 494.400 ;
        RECT 448.950 493.950 451.050 494.400 ;
        RECT 460.950 495.600 463.050 496.050 ;
        RECT 472.950 495.600 475.050 496.050 ;
        RECT 460.950 494.400 475.050 495.600 ;
        RECT 460.950 493.950 463.050 494.400 ;
        RECT 472.950 493.950 475.050 494.400 ;
        RECT 487.950 495.600 490.050 496.050 ;
        RECT 601.950 495.600 604.050 496.050 ;
        RECT 661.950 495.600 664.050 496.050 ;
        RECT 487.950 494.400 604.050 495.600 ;
        RECT 487.950 493.950 490.050 494.400 ;
        RECT 601.950 493.950 604.050 494.400 ;
        RECT 605.400 494.400 664.050 495.600 ;
        RECT 16.950 492.600 19.050 493.050 ;
        RECT 58.950 492.600 61.050 493.050 ;
        RECT 67.950 492.600 70.050 493.050 ;
        RECT 16.950 491.400 70.050 492.600 ;
        RECT 16.950 490.950 19.050 491.400 ;
        RECT 58.950 490.950 61.050 491.400 ;
        RECT 67.950 490.950 70.050 491.400 ;
        RECT 76.950 490.950 79.050 493.050 ;
        RECT 112.950 492.600 115.050 493.050 ;
        RECT 154.950 492.600 157.050 493.050 ;
        RECT 166.950 492.600 169.050 493.050 ;
        RECT 112.950 491.400 138.600 492.600 ;
        RECT 112.950 490.950 115.050 491.400 ;
        RECT 7.950 489.600 10.050 490.050 ;
        RECT 16.950 489.600 19.050 490.050 ;
        RECT 7.950 488.400 19.050 489.600 ;
        RECT 7.950 487.950 10.050 488.400 ;
        RECT 16.950 487.950 19.050 488.400 ;
        RECT 22.950 489.600 25.050 490.050 ;
        RECT 52.950 489.600 55.050 490.050 ;
        RECT 61.950 489.600 64.050 490.050 ;
        RECT 22.950 488.400 55.050 489.600 ;
        RECT 22.950 487.950 25.050 488.400 ;
        RECT 19.950 486.600 22.050 487.050 ;
        RECT 25.950 486.600 28.050 487.050 ;
        RECT 19.950 485.400 28.050 486.600 ;
        RECT 19.950 484.950 22.050 485.400 ;
        RECT 25.950 484.950 28.050 485.400 ;
        RECT 28.950 486.600 31.050 487.050 ;
        RECT 34.950 486.600 37.050 487.050 ;
        RECT 28.950 485.400 37.050 486.600 ;
        RECT 28.950 484.950 31.050 485.400 ;
        RECT 34.950 484.950 37.050 485.400 ;
        RECT 47.400 484.050 48.600 488.400 ;
        RECT 52.950 487.950 55.050 488.400 ;
        RECT 56.400 488.400 64.050 489.600 ;
        RECT 49.950 486.600 52.050 487.050 ;
        RECT 56.400 486.600 57.600 488.400 ;
        RECT 61.950 487.950 64.050 488.400 ;
        RECT 67.950 489.600 70.050 490.050 ;
        RECT 73.950 489.600 76.050 490.050 ;
        RECT 67.950 488.400 76.050 489.600 ;
        RECT 67.950 487.950 70.050 488.400 ;
        RECT 73.950 487.950 76.050 488.400 ;
        RECT 77.400 487.050 78.600 490.950 ;
        RECT 79.950 489.600 82.050 490.050 ;
        RECT 100.950 489.600 103.050 490.050 ;
        RECT 79.950 488.400 103.050 489.600 ;
        RECT 79.950 487.950 82.050 488.400 ;
        RECT 100.950 487.950 103.050 488.400 ;
        RECT 121.950 489.600 124.050 490.050 ;
        RECT 127.950 489.600 130.050 490.050 ;
        RECT 133.950 489.600 136.050 490.050 ;
        RECT 121.950 488.400 136.050 489.600 ;
        RECT 121.950 487.950 124.050 488.400 ;
        RECT 127.950 487.950 130.050 488.400 ;
        RECT 133.950 487.950 136.050 488.400 ;
        RECT 49.950 485.400 57.600 486.600 ;
        RECT 49.950 484.950 52.050 485.400 ;
        RECT 76.950 484.950 79.050 487.050 ;
        RECT 82.950 486.600 85.050 487.050 ;
        RECT 88.950 486.600 91.050 487.050 ;
        RECT 82.950 485.400 91.050 486.600 ;
        RECT 82.950 484.950 85.050 485.400 ;
        RECT 88.950 484.950 91.050 485.400 ;
        RECT 115.950 486.600 118.050 487.050 ;
        RECT 127.950 486.600 130.050 487.050 ;
        RECT 137.400 486.600 138.600 491.400 ;
        RECT 154.950 491.400 169.050 492.600 ;
        RECT 154.950 490.950 157.050 491.400 ;
        RECT 166.950 490.950 169.050 491.400 ;
        RECT 184.950 492.600 187.050 493.050 ;
        RECT 193.950 492.600 196.050 493.050 ;
        RECT 184.950 491.400 196.050 492.600 ;
        RECT 184.950 490.950 187.050 491.400 ;
        RECT 193.950 490.950 196.050 491.400 ;
        RECT 274.950 492.600 277.050 493.050 ;
        RECT 328.950 492.600 331.050 493.050 ;
        RECT 274.950 491.400 331.050 492.600 ;
        RECT 274.950 490.950 277.050 491.400 ;
        RECT 328.950 490.950 331.050 491.400 ;
        RECT 373.950 492.600 376.050 493.050 ;
        RECT 382.950 492.600 385.050 493.050 ;
        RECT 373.950 491.400 385.050 492.600 ;
        RECT 373.950 490.950 376.050 491.400 ;
        RECT 382.950 490.950 385.050 491.400 ;
        RECT 406.950 492.600 409.050 493.050 ;
        RECT 436.950 492.600 439.050 493.050 ;
        RECT 406.950 491.400 439.050 492.600 ;
        RECT 406.950 490.950 409.050 491.400 ;
        RECT 436.950 490.950 439.050 491.400 ;
        RECT 439.950 492.600 442.050 493.050 ;
        RECT 460.950 492.600 463.050 493.050 ;
        RECT 511.950 492.600 514.050 493.050 ;
        RECT 544.950 492.600 547.050 493.050 ;
        RECT 562.950 492.600 565.050 493.050 ;
        RECT 439.950 491.400 463.050 492.600 ;
        RECT 439.950 490.950 442.050 491.400 ;
        RECT 460.950 490.950 463.050 491.400 ;
        RECT 464.400 491.400 514.050 492.600 ;
        RECT 205.950 489.600 208.050 490.050 ;
        RECT 164.400 488.400 208.050 489.600 ;
        RECT 164.400 487.050 165.600 488.400 ;
        RECT 205.950 487.950 208.050 488.400 ;
        RECT 208.950 489.600 211.050 490.050 ;
        RECT 244.950 489.600 247.050 490.050 ;
        RECT 208.950 488.400 247.050 489.600 ;
        RECT 208.950 487.950 211.050 488.400 ;
        RECT 244.950 487.950 247.050 488.400 ;
        RECT 253.950 489.600 256.050 490.050 ;
        RECT 262.950 489.600 265.050 490.050 ;
        RECT 253.950 488.400 265.050 489.600 ;
        RECT 253.950 487.950 256.050 488.400 ;
        RECT 262.950 487.950 265.050 488.400 ;
        RECT 265.950 489.600 268.050 490.050 ;
        RECT 310.950 489.600 313.050 490.050 ;
        RECT 391.950 489.600 394.050 490.050 ;
        RECT 265.950 488.400 313.050 489.600 ;
        RECT 265.950 487.950 268.050 488.400 ;
        RECT 310.950 487.950 313.050 488.400 ;
        RECT 356.400 488.400 394.050 489.600 ;
        RECT 115.950 485.400 123.600 486.600 ;
        RECT 115.950 484.950 118.050 485.400 ;
        RECT 46.950 481.950 49.050 484.050 ;
        RECT 112.950 483.600 115.050 484.050 ;
        RECT 118.950 483.600 121.050 484.050 ;
        RECT 112.950 482.400 121.050 483.600 ;
        RECT 122.400 483.600 123.600 485.400 ;
        RECT 127.950 485.400 138.600 486.600 ;
        RECT 127.950 484.950 130.050 485.400 ;
        RECT 163.950 484.950 166.050 487.050 ;
        RECT 169.950 486.600 172.050 487.050 ;
        RECT 169.950 485.400 177.600 486.600 ;
        RECT 169.950 484.950 172.050 485.400 ;
        RECT 136.950 483.600 139.050 484.050 ;
        RECT 122.400 482.400 139.050 483.600 ;
        RECT 112.950 481.950 115.050 482.400 ;
        RECT 118.950 481.950 121.050 482.400 ;
        RECT 136.950 481.950 139.050 482.400 ;
        RECT 157.950 483.600 160.050 484.050 ;
        RECT 163.950 483.600 166.050 484.050 ;
        RECT 157.950 482.400 166.050 483.600 ;
        RECT 157.950 481.950 160.050 482.400 ;
        RECT 163.950 481.950 166.050 482.400 ;
        RECT 176.400 481.050 177.600 485.400 ;
        RECT 190.950 484.950 193.050 487.050 ;
        RECT 196.950 486.600 199.050 487.050 ;
        RECT 202.950 486.600 205.050 487.050 ;
        RECT 217.950 486.600 220.050 487.050 ;
        RECT 226.950 486.600 229.050 487.050 ;
        RECT 196.950 485.400 205.050 486.600 ;
        RECT 196.950 484.950 199.050 485.400 ;
        RECT 202.950 484.950 205.050 485.400 ;
        RECT 206.400 485.400 229.050 486.600 ;
        RECT 191.400 483.600 192.600 484.950 ;
        RECT 206.400 483.600 207.600 485.400 ;
        RECT 217.950 484.950 220.050 485.400 ;
        RECT 226.950 484.950 229.050 485.400 ;
        RECT 295.950 484.950 298.050 487.050 ;
        RECT 356.400 486.600 357.600 488.400 ;
        RECT 391.950 487.950 394.050 488.400 ;
        RECT 394.950 489.600 397.050 490.050 ;
        RECT 406.950 489.600 409.050 490.050 ;
        RECT 394.950 488.400 409.050 489.600 ;
        RECT 394.950 487.950 397.050 488.400 ;
        RECT 406.950 487.950 409.050 488.400 ;
        RECT 433.950 489.600 436.050 490.050 ;
        RECT 464.400 489.600 465.600 491.400 ;
        RECT 511.950 490.950 514.050 491.400 ;
        RECT 524.400 491.400 547.050 492.600 ;
        RECT 433.950 488.400 465.600 489.600 ;
        RECT 466.950 489.600 469.050 490.050 ;
        RECT 520.950 489.600 523.050 490.050 ;
        RECT 466.950 488.400 523.050 489.600 ;
        RECT 433.950 487.950 436.050 488.400 ;
        RECT 466.950 487.950 469.050 488.400 ;
        RECT 520.950 487.950 523.050 488.400 ;
        RECT 308.400 485.400 357.600 486.600 ;
        RECT 358.950 486.600 361.050 487.050 ;
        RECT 370.950 486.600 373.050 487.050 ;
        RECT 358.950 485.400 373.050 486.600 ;
        RECT 191.400 482.400 207.600 483.600 ;
        RECT 208.950 483.600 211.050 484.050 ;
        RECT 229.950 483.600 232.050 484.050 ;
        RECT 208.950 482.400 232.050 483.600 ;
        RECT 208.950 481.950 211.050 482.400 ;
        RECT 229.950 481.950 232.050 482.400 ;
        RECT 244.950 483.600 247.050 484.050 ;
        RECT 280.950 483.600 283.050 484.050 ;
        RECT 289.950 483.600 292.050 484.050 ;
        RECT 244.950 482.400 279.600 483.600 ;
        RECT 244.950 481.950 247.050 482.400 ;
        RECT 37.950 480.600 40.050 481.050 ;
        RECT 43.950 480.600 46.050 481.050 ;
        RECT 70.950 480.600 73.050 481.050 ;
        RECT 37.950 479.400 73.050 480.600 ;
        RECT 37.950 478.950 40.050 479.400 ;
        RECT 43.950 478.950 46.050 479.400 ;
        RECT 70.950 478.950 73.050 479.400 ;
        RECT 79.950 480.600 82.050 481.050 ;
        RECT 85.950 480.600 88.050 481.050 ;
        RECT 115.950 480.600 118.050 481.050 ;
        RECT 79.950 479.400 118.050 480.600 ;
        RECT 79.950 478.950 82.050 479.400 ;
        RECT 85.950 478.950 88.050 479.400 ;
        RECT 115.950 478.950 118.050 479.400 ;
        RECT 130.950 480.600 133.050 481.050 ;
        RECT 142.950 480.600 145.050 481.050 ;
        RECT 130.950 479.400 145.050 480.600 ;
        RECT 130.950 478.950 133.050 479.400 ;
        RECT 142.950 478.950 145.050 479.400 ;
        RECT 148.950 480.600 151.050 481.050 ;
        RECT 166.950 480.600 169.050 481.050 ;
        RECT 148.950 479.400 169.050 480.600 ;
        RECT 148.950 478.950 151.050 479.400 ;
        RECT 166.950 478.950 169.050 479.400 ;
        RECT 175.950 478.950 178.050 481.050 ;
        RECT 181.950 480.600 184.050 481.050 ;
        RECT 193.950 480.600 196.050 481.050 ;
        RECT 181.950 479.400 196.050 480.600 ;
        RECT 181.950 478.950 184.050 479.400 ;
        RECT 193.950 478.950 196.050 479.400 ;
        RECT 214.950 480.600 217.050 481.050 ;
        RECT 253.950 480.600 256.050 481.050 ;
        RECT 214.950 479.400 256.050 480.600 ;
        RECT 278.400 480.600 279.600 482.400 ;
        RECT 280.950 482.400 292.050 483.600 ;
        RECT 280.950 481.950 283.050 482.400 ;
        RECT 289.950 481.950 292.050 482.400 ;
        RECT 296.400 481.050 297.600 484.950 ;
        RECT 298.950 483.600 301.050 484.050 ;
        RECT 308.400 483.600 309.600 485.400 ;
        RECT 358.950 484.950 361.050 485.400 ;
        RECT 370.950 484.950 373.050 485.400 ;
        RECT 376.950 486.600 379.050 487.050 ;
        RECT 400.950 486.600 403.050 487.050 ;
        RECT 376.950 485.400 403.050 486.600 ;
        RECT 376.950 484.950 379.050 485.400 ;
        RECT 400.950 484.950 403.050 485.400 ;
        RECT 421.950 486.600 424.050 487.050 ;
        RECT 424.950 486.600 427.050 487.050 ;
        RECT 421.950 485.400 427.050 486.600 ;
        RECT 421.950 484.950 424.050 485.400 ;
        RECT 424.950 484.950 427.050 485.400 ;
        RECT 442.950 486.600 445.050 487.050 ;
        RECT 463.950 486.600 466.050 487.050 ;
        RECT 478.950 486.600 481.050 487.050 ;
        RECT 442.950 485.400 481.050 486.600 ;
        RECT 442.950 484.950 445.050 485.400 ;
        RECT 463.950 484.950 466.050 485.400 ;
        RECT 478.950 484.950 481.050 485.400 ;
        RECT 499.950 486.600 502.050 487.050 ;
        RECT 508.950 486.600 511.050 487.050 ;
        RECT 524.400 486.600 525.600 491.400 ;
        RECT 544.950 490.950 547.050 491.400 ;
        RECT 551.400 491.400 565.050 492.600 ;
        RECT 551.400 490.050 552.600 491.400 ;
        RECT 562.950 490.950 565.050 491.400 ;
        RECT 568.950 492.600 571.050 493.050 ;
        RECT 605.400 492.600 606.600 494.400 ;
        RECT 661.950 493.950 664.050 494.400 ;
        RECT 568.950 491.400 606.600 492.600 ;
        RECT 616.950 492.600 619.050 493.050 ;
        RECT 688.950 492.600 691.050 493.050 ;
        RECT 616.950 491.400 691.050 492.600 ;
        RECT 568.950 490.950 571.050 491.400 ;
        RECT 616.950 490.950 619.050 491.400 ;
        RECT 688.950 490.950 691.050 491.400 ;
        RECT 712.950 492.600 715.050 493.050 ;
        RECT 766.950 492.600 769.050 493.050 ;
        RECT 712.950 491.400 769.050 492.600 ;
        RECT 712.950 490.950 715.050 491.400 ;
        RECT 766.950 490.950 769.050 491.400 ;
        RECT 526.950 489.600 529.050 490.050 ;
        RECT 541.950 489.600 544.050 490.050 ;
        RECT 526.950 488.400 544.050 489.600 ;
        RECT 526.950 487.950 529.050 488.400 ;
        RECT 541.950 487.950 544.050 488.400 ;
        RECT 550.950 487.950 553.050 490.050 ;
        RECT 556.950 489.600 559.050 490.050 ;
        RECT 586.950 489.600 589.050 490.050 ;
        RECT 554.400 488.400 559.050 489.600 ;
        RECT 554.400 487.050 555.600 488.400 ;
        RECT 556.950 487.950 559.050 488.400 ;
        RECT 581.400 488.400 589.050 489.600 ;
        RECT 499.950 485.400 511.050 486.600 ;
        RECT 499.950 484.950 502.050 485.400 ;
        RECT 508.950 484.950 511.050 485.400 ;
        RECT 515.400 485.400 525.600 486.600 ;
        RECT 526.950 486.600 529.050 487.050 ;
        RECT 532.950 486.600 535.050 487.050 ;
        RECT 526.950 485.400 535.050 486.600 ;
        RECT 298.950 482.400 309.600 483.600 ;
        RECT 298.950 481.950 301.050 482.400 ;
        RECT 310.950 481.950 313.050 484.050 ;
        RECT 379.950 483.600 382.050 484.050 ;
        RECT 391.950 483.600 394.050 484.050 ;
        RECT 379.950 482.400 394.050 483.600 ;
        RECT 379.950 481.950 382.050 482.400 ;
        RECT 391.950 481.950 394.050 482.400 ;
        RECT 397.950 483.600 400.050 484.050 ;
        RECT 412.950 483.600 415.050 484.050 ;
        RECT 397.950 482.400 415.050 483.600 ;
        RECT 422.400 483.600 423.600 484.950 ;
        RECT 422.400 482.400 429.600 483.600 ;
        RECT 397.950 481.950 400.050 482.400 ;
        RECT 412.950 481.950 415.050 482.400 ;
        RECT 286.950 480.600 289.050 481.050 ;
        RECT 278.400 479.400 289.050 480.600 ;
        RECT 214.950 478.950 217.050 479.400 ;
        RECT 253.950 478.950 256.050 479.400 ;
        RECT 286.950 478.950 289.050 479.400 ;
        RECT 295.950 478.950 298.050 481.050 ;
        RECT 301.950 480.600 304.050 481.050 ;
        RECT 311.400 480.600 312.600 481.950 ;
        RECT 301.950 479.400 312.600 480.600 ;
        RECT 322.950 480.600 325.050 481.050 ;
        RECT 328.950 480.600 331.050 481.050 ;
        RECT 322.950 479.400 331.050 480.600 ;
        RECT 301.950 478.950 304.050 479.400 ;
        RECT 322.950 478.950 325.050 479.400 ;
        RECT 328.950 478.950 331.050 479.400 ;
        RECT 364.950 480.600 367.050 481.050 ;
        RECT 379.950 480.600 382.050 481.050 ;
        RECT 424.950 480.600 427.050 481.050 ;
        RECT 364.950 479.400 382.050 480.600 ;
        RECT 364.950 478.950 367.050 479.400 ;
        RECT 379.950 478.950 382.050 479.400 ;
        RECT 383.400 479.400 427.050 480.600 ;
        RECT 10.950 477.600 13.050 478.050 ;
        RECT 28.950 477.600 31.050 478.050 ;
        RECT 112.950 477.600 115.050 478.050 ;
        RECT 10.950 476.400 115.050 477.600 ;
        RECT 10.950 475.950 13.050 476.400 ;
        RECT 28.950 475.950 31.050 476.400 ;
        RECT 112.950 475.950 115.050 476.400 ;
        RECT 124.950 477.600 127.050 478.050 ;
        RECT 139.950 477.600 142.050 478.050 ;
        RECT 208.950 477.600 211.050 478.050 ;
        RECT 124.950 476.400 211.050 477.600 ;
        RECT 124.950 475.950 127.050 476.400 ;
        RECT 139.950 475.950 142.050 476.400 ;
        RECT 208.950 475.950 211.050 476.400 ;
        RECT 235.950 477.600 238.050 478.050 ;
        RECT 250.950 477.600 253.050 478.050 ;
        RECT 235.950 476.400 253.050 477.600 ;
        RECT 235.950 475.950 238.050 476.400 ;
        RECT 250.950 475.950 253.050 476.400 ;
        RECT 253.950 477.600 256.050 478.050 ;
        RECT 307.950 477.600 310.050 478.050 ;
        RECT 383.400 477.600 384.600 479.400 ;
        RECT 424.950 478.950 427.050 479.400 ;
        RECT 428.400 478.050 429.600 482.400 ;
        RECT 445.950 480.600 448.050 481.050 ;
        RECT 487.950 480.600 490.050 481.050 ;
        RECT 445.950 479.400 490.050 480.600 ;
        RECT 500.400 480.600 501.600 484.950 ;
        RECT 515.400 484.050 516.600 485.400 ;
        RECT 526.950 484.950 529.050 485.400 ;
        RECT 532.950 484.950 535.050 485.400 ;
        RECT 538.950 486.600 541.050 487.050 ;
        RECT 547.950 486.600 550.050 487.050 ;
        RECT 538.950 485.400 550.050 486.600 ;
        RECT 538.950 484.950 541.050 485.400 ;
        RECT 547.950 484.950 550.050 485.400 ;
        RECT 553.950 484.950 556.050 487.050 ;
        RECT 559.950 486.600 562.050 487.050 ;
        RECT 557.400 485.400 562.050 486.600 ;
        RECT 502.950 483.600 505.050 484.050 ;
        RECT 502.950 482.400 507.600 483.600 ;
        RECT 502.950 481.950 505.050 482.400 ;
        RECT 502.950 480.600 505.050 481.050 ;
        RECT 500.400 479.400 505.050 480.600 ;
        RECT 506.400 480.600 507.600 482.400 ;
        RECT 514.950 481.950 517.050 484.050 ;
        RECT 550.950 483.600 553.050 484.050 ;
        RECT 536.400 482.400 553.050 483.600 ;
        RECT 536.400 481.050 537.600 482.400 ;
        RECT 550.950 481.950 553.050 482.400 ;
        RECT 553.950 483.600 556.050 484.050 ;
        RECT 557.400 483.600 558.600 485.400 ;
        RECT 559.950 484.950 562.050 485.400 ;
        RECT 553.950 482.400 558.600 483.600 ;
        RECT 562.950 483.600 565.050 484.050 ;
        RECT 571.950 483.600 574.050 484.050 ;
        RECT 562.950 482.400 574.050 483.600 ;
        RECT 553.950 481.950 556.050 482.400 ;
        RECT 562.950 481.950 565.050 482.400 ;
        RECT 571.950 481.950 574.050 482.400 ;
        RECT 574.950 483.600 577.050 484.050 ;
        RECT 581.400 483.600 582.600 488.400 ;
        RECT 586.950 487.950 589.050 488.400 ;
        RECT 589.950 489.600 592.050 490.050 ;
        RECT 595.950 489.600 598.050 490.050 ;
        RECT 589.950 488.400 598.050 489.600 ;
        RECT 589.950 487.950 592.050 488.400 ;
        RECT 595.950 487.950 598.050 488.400 ;
        RECT 607.950 489.600 610.050 490.050 ;
        RECT 628.950 489.600 631.050 490.050 ;
        RECT 607.950 488.400 631.050 489.600 ;
        RECT 607.950 487.950 610.050 488.400 ;
        RECT 628.950 487.950 631.050 488.400 ;
        RECT 658.950 489.600 661.050 490.050 ;
        RECT 682.950 489.600 685.050 490.050 ;
        RECT 658.950 488.400 685.050 489.600 ;
        RECT 658.950 487.950 661.050 488.400 ;
        RECT 583.950 484.950 586.050 487.050 ;
        RECT 589.950 486.600 592.050 487.050 ;
        RECT 616.950 486.600 619.050 487.050 ;
        RECT 589.950 485.400 619.050 486.600 ;
        RECT 589.950 484.950 592.050 485.400 ;
        RECT 616.950 484.950 619.050 485.400 ;
        RECT 634.950 486.600 637.050 487.050 ;
        RECT 640.950 486.600 643.050 487.050 ;
        RECT 634.950 485.400 643.050 486.600 ;
        RECT 634.950 484.950 637.050 485.400 ;
        RECT 640.950 484.950 643.050 485.400 ;
        RECT 658.950 484.950 661.050 487.050 ;
        RECT 574.950 482.400 582.600 483.600 ;
        RECT 574.950 481.950 577.050 482.400 ;
        RECT 529.950 480.600 532.050 481.050 ;
        RECT 506.400 479.400 532.050 480.600 ;
        RECT 445.950 478.950 448.050 479.400 ;
        RECT 487.950 478.950 490.050 479.400 ;
        RECT 502.950 478.950 505.050 479.400 ;
        RECT 529.950 478.950 532.050 479.400 ;
        RECT 535.950 478.950 538.050 481.050 ;
        RECT 538.950 480.600 541.050 481.050 ;
        RECT 556.950 480.600 559.050 481.050 ;
        RECT 538.950 479.400 559.050 480.600 ;
        RECT 538.950 478.950 541.050 479.400 ;
        RECT 556.950 478.950 559.050 479.400 ;
        RECT 568.950 480.600 571.050 481.050 ;
        RECT 584.400 480.600 585.600 484.950 ;
        RECT 595.950 483.600 598.050 484.050 ;
        RECT 601.950 483.600 604.050 484.050 ;
        RECT 595.950 482.400 604.050 483.600 ;
        RECT 595.950 481.950 598.050 482.400 ;
        RECT 601.950 481.950 604.050 482.400 ;
        RECT 613.950 483.600 616.050 484.050 ;
        RECT 637.950 483.600 640.050 484.050 ;
        RECT 659.400 483.600 660.600 484.950 ;
        RECT 613.950 482.400 660.600 483.600 ;
        RECT 613.950 481.950 616.050 482.400 ;
        RECT 637.950 481.950 640.050 482.400 ;
        RECT 568.950 479.400 585.600 480.600 ;
        RECT 586.950 480.600 589.050 481.050 ;
        RECT 613.950 480.600 616.050 481.050 ;
        RECT 586.950 479.400 616.050 480.600 ;
        RECT 568.950 478.950 571.050 479.400 ;
        RECT 586.950 478.950 589.050 479.400 ;
        RECT 613.950 478.950 616.050 479.400 ;
        RECT 631.950 480.600 634.050 481.050 ;
        RECT 649.950 480.600 652.050 481.050 ;
        RECT 655.950 480.600 658.050 481.050 ;
        RECT 631.950 479.400 658.050 480.600 ;
        RECT 631.950 478.950 634.050 479.400 ;
        RECT 649.950 478.950 652.050 479.400 ;
        RECT 655.950 478.950 658.050 479.400 ;
        RECT 658.950 480.600 661.050 481.050 ;
        RECT 662.400 480.600 663.600 488.400 ;
        RECT 682.950 487.950 685.050 488.400 ;
        RECT 706.950 489.600 709.050 490.050 ;
        RECT 706.950 488.400 765.600 489.600 ;
        RECT 706.950 487.950 709.050 488.400 ;
        RECT 664.950 484.950 667.050 487.050 ;
        RECT 685.950 486.600 688.050 487.050 ;
        RECT 697.950 486.600 700.050 487.050 ;
        RECT 685.950 485.400 700.050 486.600 ;
        RECT 685.950 484.950 688.050 485.400 ;
        RECT 697.950 484.950 700.050 485.400 ;
        RECT 703.950 486.600 706.050 487.050 ;
        RECT 712.950 486.600 715.050 487.050 ;
        RECT 703.950 485.400 715.050 486.600 ;
        RECT 703.950 484.950 706.050 485.400 ;
        RECT 712.950 484.950 715.050 485.400 ;
        RECT 718.950 486.600 721.050 487.050 ;
        RECT 742.950 486.600 745.050 487.050 ;
        RECT 718.950 485.400 745.050 486.600 ;
        RECT 718.950 484.950 721.050 485.400 ;
        RECT 742.950 484.950 745.050 485.400 ;
        RECT 751.950 486.600 754.050 487.050 ;
        RECT 751.950 485.400 762.600 486.600 ;
        RECT 751.950 484.950 754.050 485.400 ;
        RECT 665.400 483.600 666.600 484.950 ;
        RECT 761.400 484.050 762.600 485.400 ;
        RECT 676.950 483.600 679.050 484.050 ;
        RECT 665.400 482.400 679.050 483.600 ;
        RECT 676.950 481.950 679.050 482.400 ;
        RECT 694.950 483.600 697.050 484.050 ;
        RECT 715.950 483.600 718.050 484.050 ;
        RECT 694.950 482.400 718.050 483.600 ;
        RECT 694.950 481.950 697.050 482.400 ;
        RECT 715.950 481.950 718.050 482.400 ;
        RECT 733.950 483.600 736.050 484.050 ;
        RECT 748.950 483.600 751.050 484.050 ;
        RECT 757.950 483.600 760.050 484.050 ;
        RECT 733.950 482.400 760.050 483.600 ;
        RECT 733.950 481.950 736.050 482.400 ;
        RECT 748.950 481.950 751.050 482.400 ;
        RECT 757.950 481.950 760.050 482.400 ;
        RECT 760.950 481.950 763.050 484.050 ;
        RECT 677.400 480.600 678.600 481.950 ;
        RECT 658.950 479.400 663.600 480.600 ;
        RECT 674.400 479.400 678.600 480.600 ;
        RECT 697.950 480.600 700.050 481.050 ;
        RECT 709.950 480.600 712.050 481.050 ;
        RECT 727.950 480.600 730.050 481.050 ;
        RECT 697.950 479.400 712.050 480.600 ;
        RECT 658.950 478.950 661.050 479.400 ;
        RECT 253.950 476.400 384.600 477.600 ;
        RECT 253.950 475.950 256.050 476.400 ;
        RECT 307.950 475.950 310.050 476.400 ;
        RECT 427.950 475.950 430.050 478.050 ;
        RECT 436.950 477.600 439.050 478.050 ;
        RECT 556.950 477.600 559.050 478.050 ;
        RECT 674.400 477.600 675.600 479.400 ;
        RECT 697.950 478.950 700.050 479.400 ;
        RECT 709.950 478.950 712.050 479.400 ;
        RECT 716.400 479.400 730.050 480.600 ;
        RECT 764.400 480.600 765.600 488.400 ;
        RECT 766.950 480.600 769.050 481.050 ;
        RECT 764.400 479.400 769.050 480.600 ;
        RECT 716.400 478.050 717.600 479.400 ;
        RECT 727.950 478.950 730.050 479.400 ;
        RECT 766.950 478.950 769.050 479.400 ;
        RECT 436.950 476.400 546.600 477.600 ;
        RECT 436.950 475.950 439.050 476.400 ;
        RECT 94.950 474.600 97.050 475.050 ;
        RECT 148.950 474.600 151.050 475.050 ;
        RECT 94.950 473.400 151.050 474.600 ;
        RECT 94.950 472.950 97.050 473.400 ;
        RECT 148.950 472.950 151.050 473.400 ;
        RECT 193.950 474.600 196.050 475.050 ;
        RECT 214.950 474.600 217.050 475.050 ;
        RECT 193.950 473.400 217.050 474.600 ;
        RECT 193.950 472.950 196.050 473.400 ;
        RECT 214.950 472.950 217.050 473.400 ;
        RECT 283.950 474.600 286.050 475.050 ;
        RECT 289.950 474.600 292.050 475.050 ;
        RECT 283.950 473.400 292.050 474.600 ;
        RECT 283.950 472.950 286.050 473.400 ;
        RECT 289.950 472.950 292.050 473.400 ;
        RECT 304.950 474.600 307.050 475.050 ;
        RECT 496.950 474.600 499.050 475.050 ;
        RECT 304.950 473.400 499.050 474.600 ;
        RECT 545.400 474.600 546.600 476.400 ;
        RECT 556.950 476.400 675.600 477.600 ;
        RECT 682.950 477.600 685.050 478.050 ;
        RECT 700.950 477.600 703.050 478.050 ;
        RECT 682.950 476.400 703.050 477.600 ;
        RECT 556.950 475.950 559.050 476.400 ;
        RECT 682.950 475.950 685.050 476.400 ;
        RECT 700.950 475.950 703.050 476.400 ;
        RECT 706.950 477.600 709.050 478.050 ;
        RECT 715.950 477.600 718.050 478.050 ;
        RECT 706.950 476.400 718.050 477.600 ;
        RECT 706.950 475.950 709.050 476.400 ;
        RECT 715.950 475.950 718.050 476.400 ;
        RECT 724.950 477.600 727.050 478.050 ;
        RECT 751.950 477.600 754.050 478.050 ;
        RECT 754.950 477.600 757.050 478.050 ;
        RECT 724.950 476.400 757.050 477.600 ;
        RECT 724.950 475.950 727.050 476.400 ;
        RECT 751.950 475.950 754.050 476.400 ;
        RECT 754.950 475.950 757.050 476.400 ;
        RECT 562.950 474.600 565.050 475.050 ;
        RECT 545.400 473.400 565.050 474.600 ;
        RECT 304.950 472.950 307.050 473.400 ;
        RECT 496.950 472.950 499.050 473.400 ;
        RECT 562.950 472.950 565.050 473.400 ;
        RECT 580.950 474.600 583.050 475.050 ;
        RECT 592.950 474.600 595.050 475.050 ;
        RECT 580.950 473.400 595.050 474.600 ;
        RECT 580.950 472.950 583.050 473.400 ;
        RECT 592.950 472.950 595.050 473.400 ;
        RECT 595.950 474.600 598.050 475.050 ;
        RECT 616.950 474.600 619.050 475.050 ;
        RECT 595.950 473.400 619.050 474.600 ;
        RECT 595.950 472.950 598.050 473.400 ;
        RECT 616.950 472.950 619.050 473.400 ;
        RECT 628.950 474.600 631.050 475.050 ;
        RECT 661.950 474.600 664.050 475.050 ;
        RECT 628.950 473.400 664.050 474.600 ;
        RECT 628.950 472.950 631.050 473.400 ;
        RECT 661.950 472.950 664.050 473.400 ;
        RECT 667.950 474.600 670.050 475.050 ;
        RECT 679.950 474.600 682.050 475.050 ;
        RECT 667.950 473.400 682.050 474.600 ;
        RECT 667.950 472.950 670.050 473.400 ;
        RECT 679.950 472.950 682.050 473.400 ;
        RECT 688.950 474.600 691.050 475.050 ;
        RECT 712.950 474.600 715.050 475.050 ;
        RECT 688.950 473.400 715.050 474.600 ;
        RECT 688.950 472.950 691.050 473.400 ;
        RECT 712.950 472.950 715.050 473.400 ;
        RECT 721.950 474.600 724.050 475.050 ;
        RECT 727.950 474.600 730.050 475.050 ;
        RECT 721.950 473.400 730.050 474.600 ;
        RECT 721.950 472.950 724.050 473.400 ;
        RECT 727.950 472.950 730.050 473.400 ;
        RECT 736.950 474.600 739.050 475.050 ;
        RECT 757.950 474.600 760.050 475.050 ;
        RECT 736.950 473.400 760.050 474.600 ;
        RECT 736.950 472.950 739.050 473.400 ;
        RECT 757.950 472.950 760.050 473.400 ;
        RECT 127.950 471.600 130.050 472.050 ;
        RECT 136.950 471.600 139.050 472.050 ;
        RECT 142.950 471.600 145.050 472.050 ;
        RECT 286.950 471.600 289.050 472.050 ;
        RECT 127.950 470.400 289.050 471.600 ;
        RECT 127.950 469.950 130.050 470.400 ;
        RECT 136.950 469.950 139.050 470.400 ;
        RECT 142.950 469.950 145.050 470.400 ;
        RECT 286.950 469.950 289.050 470.400 ;
        RECT 367.950 471.600 370.050 472.050 ;
        RECT 385.950 471.600 388.050 472.050 ;
        RECT 367.950 470.400 388.050 471.600 ;
        RECT 367.950 469.950 370.050 470.400 ;
        RECT 385.950 469.950 388.050 470.400 ;
        RECT 442.950 471.600 445.050 472.050 ;
        RECT 457.950 471.600 460.050 472.050 ;
        RECT 442.950 470.400 460.050 471.600 ;
        RECT 442.950 469.950 445.050 470.400 ;
        RECT 457.950 469.950 460.050 470.400 ;
        RECT 463.950 471.600 466.050 472.050 ;
        RECT 517.950 471.600 520.050 472.050 ;
        RECT 538.950 471.600 541.050 472.050 ;
        RECT 463.950 470.400 541.050 471.600 ;
        RECT 463.950 469.950 466.050 470.400 ;
        RECT 517.950 469.950 520.050 470.400 ;
        RECT 538.950 469.950 541.050 470.400 ;
        RECT 541.950 471.600 544.050 472.050 ;
        RECT 559.950 471.600 562.050 472.050 ;
        RECT 541.950 470.400 562.050 471.600 ;
        RECT 541.950 469.950 544.050 470.400 ;
        RECT 559.950 469.950 562.050 470.400 ;
        RECT 565.950 471.600 568.050 472.050 ;
        RECT 589.950 471.600 592.050 472.050 ;
        RECT 565.950 470.400 592.050 471.600 ;
        RECT 565.950 469.950 568.050 470.400 ;
        RECT 589.950 469.950 592.050 470.400 ;
        RECT 598.950 471.600 601.050 472.050 ;
        RECT 643.950 471.600 646.050 472.050 ;
        RECT 598.950 470.400 646.050 471.600 ;
        RECT 598.950 469.950 601.050 470.400 ;
        RECT 643.950 469.950 646.050 470.400 ;
        RECT 652.950 471.600 655.050 472.050 ;
        RECT 673.950 471.600 676.050 472.050 ;
        RECT 652.950 470.400 676.050 471.600 ;
        RECT 652.950 469.950 655.050 470.400 ;
        RECT 673.950 469.950 676.050 470.400 ;
        RECT 688.950 471.600 691.050 472.050 ;
        RECT 718.950 471.600 721.050 472.050 ;
        RECT 688.950 470.400 721.050 471.600 ;
        RECT 688.950 469.950 691.050 470.400 ;
        RECT 718.950 469.950 721.050 470.400 ;
        RECT 40.950 468.600 43.050 469.050 ;
        RECT 73.950 468.600 76.050 469.050 ;
        RECT 82.950 468.600 85.050 469.050 ;
        RECT 151.950 468.600 154.050 469.050 ;
        RECT 268.950 468.600 271.050 469.050 ;
        RECT 40.950 467.400 154.050 468.600 ;
        RECT 40.950 466.950 43.050 467.400 ;
        RECT 73.950 466.950 76.050 467.400 ;
        RECT 82.950 466.950 85.050 467.400 ;
        RECT 151.950 466.950 154.050 467.400 ;
        RECT 155.400 467.400 271.050 468.600 ;
        RECT 155.400 465.600 156.600 467.400 ;
        RECT 268.950 466.950 271.050 467.400 ;
        RECT 280.950 468.600 283.050 469.050 ;
        RECT 292.950 468.600 295.050 469.050 ;
        RECT 280.950 467.400 295.050 468.600 ;
        RECT 280.950 466.950 283.050 467.400 ;
        RECT 292.950 466.950 295.050 467.400 ;
        RECT 301.950 468.600 304.050 469.050 ;
        RECT 307.950 468.600 310.050 469.050 ;
        RECT 301.950 467.400 310.050 468.600 ;
        RECT 301.950 466.950 304.050 467.400 ;
        RECT 307.950 466.950 310.050 467.400 ;
        RECT 358.950 468.600 361.050 469.050 ;
        RECT 394.950 468.600 397.050 469.050 ;
        RECT 409.950 468.600 412.050 469.050 ;
        RECT 418.950 468.600 421.050 469.050 ;
        RECT 358.950 467.400 421.050 468.600 ;
        RECT 358.950 466.950 361.050 467.400 ;
        RECT 394.950 466.950 397.050 467.400 ;
        RECT 409.950 466.950 412.050 467.400 ;
        RECT 418.950 466.950 421.050 467.400 ;
        RECT 526.950 468.600 529.050 469.050 ;
        RECT 556.950 468.600 559.050 469.050 ;
        RECT 526.950 467.400 559.050 468.600 ;
        RECT 526.950 466.950 529.050 467.400 ;
        RECT 556.950 466.950 559.050 467.400 ;
        RECT 574.950 468.600 577.050 469.050 ;
        RECT 586.950 468.600 589.050 469.050 ;
        RECT 574.950 467.400 589.050 468.600 ;
        RECT 574.950 466.950 577.050 467.400 ;
        RECT 586.950 466.950 589.050 467.400 ;
        RECT 592.950 468.600 595.050 469.050 ;
        RECT 601.950 468.600 604.050 469.050 ;
        RECT 592.950 467.400 604.050 468.600 ;
        RECT 592.950 466.950 595.050 467.400 ;
        RECT 601.950 466.950 604.050 467.400 ;
        RECT 619.950 468.600 622.050 469.050 ;
        RECT 634.950 468.600 637.050 469.050 ;
        RECT 670.950 468.600 673.050 469.050 ;
        RECT 619.950 467.400 673.050 468.600 ;
        RECT 619.950 466.950 622.050 467.400 ;
        RECT 634.950 466.950 637.050 467.400 ;
        RECT 670.950 466.950 673.050 467.400 ;
        RECT 679.950 468.600 682.050 469.050 ;
        RECT 709.950 468.600 712.050 469.050 ;
        RECT 736.950 468.600 739.050 469.050 ;
        RECT 679.950 467.400 739.050 468.600 ;
        RECT 679.950 466.950 682.050 467.400 ;
        RECT 709.950 466.950 712.050 467.400 ;
        RECT 736.950 466.950 739.050 467.400 ;
        RECT 62.400 464.400 156.600 465.600 ;
        RECT 160.950 465.600 163.050 466.050 ;
        RECT 220.950 465.600 223.050 466.050 ;
        RECT 160.950 464.400 223.050 465.600 ;
        RECT 16.950 462.600 19.050 463.050 ;
        RECT 25.950 462.600 28.050 463.050 ;
        RECT 16.950 461.400 28.050 462.600 ;
        RECT 16.950 460.950 19.050 461.400 ;
        RECT 25.950 460.950 28.050 461.400 ;
        RECT 55.950 462.600 58.050 463.050 ;
        RECT 62.400 462.600 63.600 464.400 ;
        RECT 160.950 463.950 163.050 464.400 ;
        RECT 220.950 463.950 223.050 464.400 ;
        RECT 223.950 465.600 226.050 466.050 ;
        RECT 247.950 465.600 250.050 466.050 ;
        RECT 265.950 465.600 268.050 466.050 ;
        RECT 325.950 465.600 328.050 466.050 ;
        RECT 223.950 464.400 328.050 465.600 ;
        RECT 223.950 463.950 226.050 464.400 ;
        RECT 247.950 463.950 250.050 464.400 ;
        RECT 265.950 463.950 268.050 464.400 ;
        RECT 325.950 463.950 328.050 464.400 ;
        RECT 376.950 465.600 379.050 466.050 ;
        RECT 382.950 465.600 385.050 466.050 ;
        RECT 376.950 464.400 385.050 465.600 ;
        RECT 376.950 463.950 379.050 464.400 ;
        RECT 382.950 463.950 385.050 464.400 ;
        RECT 418.950 465.600 421.050 466.050 ;
        RECT 433.950 465.600 436.050 466.050 ;
        RECT 418.950 464.400 436.050 465.600 ;
        RECT 418.950 463.950 421.050 464.400 ;
        RECT 433.950 463.950 436.050 464.400 ;
        RECT 478.950 465.600 481.050 466.050 ;
        RECT 523.950 465.600 526.050 466.050 ;
        RECT 478.950 464.400 526.050 465.600 ;
        RECT 478.950 463.950 481.050 464.400 ;
        RECT 523.950 463.950 526.050 464.400 ;
        RECT 547.950 465.600 550.050 466.050 ;
        RECT 571.950 465.600 574.050 466.050 ;
        RECT 547.950 464.400 574.050 465.600 ;
        RECT 547.950 463.950 550.050 464.400 ;
        RECT 571.950 463.950 574.050 464.400 ;
        RECT 601.950 465.600 604.050 466.050 ;
        RECT 628.950 465.600 631.050 466.050 ;
        RECT 601.950 464.400 631.050 465.600 ;
        RECT 601.950 463.950 604.050 464.400 ;
        RECT 628.950 463.950 631.050 464.400 ;
        RECT 643.950 465.600 646.050 466.050 ;
        RECT 718.950 465.600 721.050 466.050 ;
        RECT 643.950 464.400 721.050 465.600 ;
        RECT 643.950 463.950 646.050 464.400 ;
        RECT 718.950 463.950 721.050 464.400 ;
        RECT 721.950 465.600 724.050 466.050 ;
        RECT 763.950 465.600 766.050 466.050 ;
        RECT 721.950 464.400 766.050 465.600 ;
        RECT 721.950 463.950 724.050 464.400 ;
        RECT 763.950 463.950 766.050 464.400 ;
        RECT 55.950 461.400 63.600 462.600 ;
        RECT 130.950 462.600 133.050 463.050 ;
        RECT 172.950 462.600 175.050 463.050 ;
        RECT 130.950 461.400 175.050 462.600 ;
        RECT 55.950 460.950 58.050 461.400 ;
        RECT 130.950 460.950 133.050 461.400 ;
        RECT 172.950 460.950 175.050 461.400 ;
        RECT 184.950 462.600 187.050 463.050 ;
        RECT 211.950 462.600 214.050 463.050 ;
        RECT 223.950 462.600 226.050 463.050 ;
        RECT 247.950 462.600 250.050 463.050 ;
        RECT 184.950 461.400 210.600 462.600 ;
        RECT 184.950 460.950 187.050 461.400 ;
        RECT 7.950 459.600 10.050 460.050 ;
        RECT 55.950 459.600 58.050 460.050 ;
        RECT 7.950 458.400 58.050 459.600 ;
        RECT 7.950 457.950 10.050 458.400 ;
        RECT 55.950 457.950 58.050 458.400 ;
        RECT 58.950 459.600 61.050 460.050 ;
        RECT 91.950 459.600 94.050 460.050 ;
        RECT 58.950 458.400 94.050 459.600 ;
        RECT 58.950 457.950 61.050 458.400 ;
        RECT 91.950 457.950 94.050 458.400 ;
        RECT 100.950 459.600 103.050 460.050 ;
        RECT 118.950 459.600 121.050 460.050 ;
        RECT 100.950 458.400 121.050 459.600 ;
        RECT 100.950 457.950 103.050 458.400 ;
        RECT 118.950 457.950 121.050 458.400 ;
        RECT 175.950 459.600 178.050 460.050 ;
        RECT 184.950 459.600 187.050 460.050 ;
        RECT 193.950 459.600 196.050 460.050 ;
        RECT 175.950 458.400 187.050 459.600 ;
        RECT 175.950 457.950 178.050 458.400 ;
        RECT 184.950 457.950 187.050 458.400 ;
        RECT 188.400 458.400 196.050 459.600 ;
        RECT 209.400 459.600 210.600 461.400 ;
        RECT 211.950 461.400 226.050 462.600 ;
        RECT 211.950 460.950 214.050 461.400 ;
        RECT 223.950 460.950 226.050 461.400 ;
        RECT 230.400 461.400 250.050 462.600 ;
        RECT 217.950 459.600 220.050 460.050 ;
        RECT 209.400 458.400 220.050 459.600 ;
        RECT 13.950 456.600 16.050 457.050 ;
        RECT 22.950 456.600 25.050 457.050 ;
        RECT 59.400 456.600 60.600 457.950 ;
        RECT 13.950 455.400 21.600 456.600 ;
        RECT 13.950 454.950 16.050 455.400 ;
        RECT 20.400 454.050 21.600 455.400 ;
        RECT 22.950 455.400 60.600 456.600 ;
        RECT 106.950 456.600 109.050 457.050 ;
        RECT 121.950 456.600 124.050 457.050 ;
        RECT 151.950 456.600 154.050 457.050 ;
        RECT 106.950 455.400 124.050 456.600 ;
        RECT 22.950 454.950 25.050 455.400 ;
        RECT 106.950 454.950 109.050 455.400 ;
        RECT 121.950 454.950 124.050 455.400 ;
        RECT 143.400 455.400 154.050 456.600 ;
        RECT 143.400 454.050 144.600 455.400 ;
        RECT 151.950 454.950 154.050 455.400 ;
        RECT 166.950 456.600 169.050 457.050 ;
        RECT 178.950 456.600 181.050 457.050 ;
        RECT 166.950 455.400 181.050 456.600 ;
        RECT 166.950 454.950 169.050 455.400 ;
        RECT 178.950 454.950 181.050 455.400 ;
        RECT 181.950 456.600 184.050 457.050 ;
        RECT 188.400 456.600 189.600 458.400 ;
        RECT 193.950 457.950 196.050 458.400 ;
        RECT 217.950 457.950 220.050 458.400 ;
        RECT 220.950 459.600 223.050 460.050 ;
        RECT 230.400 459.600 231.600 461.400 ;
        RECT 247.950 460.950 250.050 461.400 ;
        RECT 337.950 462.600 340.050 463.050 ;
        RECT 400.950 462.600 403.050 463.050 ;
        RECT 337.950 461.400 403.050 462.600 ;
        RECT 337.950 460.950 340.050 461.400 ;
        RECT 400.950 460.950 403.050 461.400 ;
        RECT 412.950 462.600 415.050 463.050 ;
        RECT 463.950 462.600 466.050 463.050 ;
        RECT 412.950 461.400 466.050 462.600 ;
        RECT 412.950 460.950 415.050 461.400 ;
        RECT 463.950 460.950 466.050 461.400 ;
        RECT 508.950 462.600 511.050 463.050 ;
        RECT 517.950 462.600 520.050 463.050 ;
        RECT 508.950 461.400 520.050 462.600 ;
        RECT 508.950 460.950 511.050 461.400 ;
        RECT 517.950 460.950 520.050 461.400 ;
        RECT 532.950 462.600 535.050 463.050 ;
        RECT 553.950 462.600 556.050 463.050 ;
        RECT 532.950 461.400 556.050 462.600 ;
        RECT 532.950 460.950 535.050 461.400 ;
        RECT 553.950 460.950 556.050 461.400 ;
        RECT 559.950 462.600 562.050 463.050 ;
        RECT 598.950 462.600 601.050 463.050 ;
        RECT 613.950 462.600 616.050 463.050 ;
        RECT 682.950 462.600 685.050 463.050 ;
        RECT 559.950 461.400 567.600 462.600 ;
        RECT 559.950 460.950 562.050 461.400 ;
        RECT 220.950 458.400 231.600 459.600 ;
        RECT 232.950 459.600 235.050 460.050 ;
        RECT 241.950 459.600 244.050 460.050 ;
        RECT 232.950 458.400 244.050 459.600 ;
        RECT 220.950 457.950 223.050 458.400 ;
        RECT 232.950 457.950 235.050 458.400 ;
        RECT 241.950 457.950 244.050 458.400 ;
        RECT 262.950 459.600 265.050 460.050 ;
        RECT 271.950 459.600 274.050 460.050 ;
        RECT 262.950 458.400 274.050 459.600 ;
        RECT 262.950 457.950 265.050 458.400 ;
        RECT 271.950 457.950 274.050 458.400 ;
        RECT 274.950 459.600 277.050 460.050 ;
        RECT 295.950 459.600 298.050 460.050 ;
        RECT 337.950 459.600 340.050 460.050 ;
        RECT 274.950 458.400 298.050 459.600 ;
        RECT 274.950 457.950 277.050 458.400 ;
        RECT 295.950 457.950 298.050 458.400 ;
        RECT 314.400 458.400 340.050 459.600 ;
        RECT 181.950 455.400 189.600 456.600 ;
        RECT 181.950 454.950 184.050 455.400 ;
        RECT 190.950 454.950 193.050 457.050 ;
        RECT 196.950 456.600 199.050 457.050 ;
        RECT 205.950 456.600 208.050 457.050 ;
        RECT 214.950 456.600 217.050 457.050 ;
        RECT 196.950 455.400 208.050 456.600 ;
        RECT 196.950 454.950 199.050 455.400 ;
        RECT 205.950 454.950 208.050 455.400 ;
        RECT 209.400 455.400 217.050 456.600 ;
        RECT 4.950 453.600 7.050 454.050 ;
        RECT 13.950 453.600 16.050 454.050 ;
        RECT 4.950 452.400 16.050 453.600 ;
        RECT 4.950 451.950 7.050 452.400 ;
        RECT 13.950 451.950 16.050 452.400 ;
        RECT 19.950 451.950 22.050 454.050 ;
        RECT 64.950 453.600 67.050 454.050 ;
        RECT 85.950 453.600 88.050 454.050 ;
        RECT 64.950 452.400 88.050 453.600 ;
        RECT 64.950 451.950 67.050 452.400 ;
        RECT 85.950 451.950 88.050 452.400 ;
        RECT 112.950 451.950 115.050 454.050 ;
        RECT 118.950 453.600 121.050 454.050 ;
        RECT 116.400 452.400 121.050 453.600 ;
        RECT 31.950 450.600 34.050 451.050 ;
        RECT 46.950 450.600 49.050 451.050 ;
        RECT 31.950 449.400 49.050 450.600 ;
        RECT 31.950 448.950 34.050 449.400 ;
        RECT 46.950 448.950 49.050 449.400 ;
        RECT 52.950 450.600 55.050 451.050 ;
        RECT 61.950 450.600 64.050 451.050 ;
        RECT 52.950 449.400 64.050 450.600 ;
        RECT 52.950 448.950 55.050 449.400 ;
        RECT 61.950 448.950 64.050 449.400 ;
        RECT 113.400 447.600 114.600 451.950 ;
        RECT 116.400 451.050 117.600 452.400 ;
        RECT 118.950 451.950 121.050 452.400 ;
        RECT 124.950 453.600 127.050 454.050 ;
        RECT 139.950 453.600 142.050 454.050 ;
        RECT 124.950 452.400 142.050 453.600 ;
        RECT 124.950 451.950 127.050 452.400 ;
        RECT 139.950 451.950 142.050 452.400 ;
        RECT 142.950 451.950 145.050 454.050 ;
        RECT 169.950 451.950 172.050 454.050 ;
        RECT 191.400 453.600 192.600 454.950 ;
        RECT 193.950 453.600 196.050 454.050 ;
        RECT 209.400 453.600 210.600 455.400 ;
        RECT 214.950 454.950 217.050 455.400 ;
        RECT 229.950 454.950 232.050 457.050 ;
        RECT 247.950 454.950 250.050 457.050 ;
        RECT 250.950 456.600 253.050 457.050 ;
        RECT 259.950 456.600 262.050 457.050 ;
        RECT 250.950 455.400 262.050 456.600 ;
        RECT 250.950 454.950 253.050 455.400 ;
        RECT 259.950 454.950 262.050 455.400 ;
        RECT 268.950 456.600 271.050 457.050 ;
        RECT 277.950 456.600 280.050 457.050 ;
        RECT 314.400 456.600 315.600 458.400 ;
        RECT 337.950 457.950 340.050 458.400 ;
        RECT 343.950 459.600 346.050 460.050 ;
        RECT 364.950 459.600 367.050 460.050 ;
        RECT 343.950 458.400 367.050 459.600 ;
        RECT 343.950 457.950 346.050 458.400 ;
        RECT 364.950 457.950 367.050 458.400 ;
        RECT 379.950 459.600 382.050 460.050 ;
        RECT 397.950 459.600 400.050 460.050 ;
        RECT 379.950 458.400 400.050 459.600 ;
        RECT 379.950 457.950 382.050 458.400 ;
        RECT 397.950 457.950 400.050 458.400 ;
        RECT 415.950 459.600 418.050 460.050 ;
        RECT 427.950 459.600 430.050 460.050 ;
        RECT 415.950 458.400 430.050 459.600 ;
        RECT 415.950 457.950 418.050 458.400 ;
        RECT 427.950 457.950 430.050 458.400 ;
        RECT 505.950 459.600 508.050 460.050 ;
        RECT 514.950 459.600 517.050 460.050 ;
        RECT 505.950 458.400 517.050 459.600 ;
        RECT 505.950 457.950 508.050 458.400 ;
        RECT 514.950 457.950 517.050 458.400 ;
        RECT 544.950 457.950 547.050 460.050 ;
        RECT 562.950 457.950 565.050 460.050 ;
        RECT 566.400 459.600 567.600 461.400 ;
        RECT 598.950 461.400 685.050 462.600 ;
        RECT 598.950 460.950 601.050 461.400 ;
        RECT 613.950 460.950 616.050 461.400 ;
        RECT 682.950 460.950 685.050 461.400 ;
        RECT 685.950 462.600 688.050 463.050 ;
        RECT 703.950 462.600 706.050 463.050 ;
        RECT 685.950 461.400 706.050 462.600 ;
        RECT 685.950 460.950 688.050 461.400 ;
        RECT 703.950 460.950 706.050 461.400 ;
        RECT 718.950 462.600 721.050 463.050 ;
        RECT 733.950 462.600 736.050 463.050 ;
        RECT 718.950 461.400 736.050 462.600 ;
        RECT 718.950 460.950 721.050 461.400 ;
        RECT 733.950 460.950 736.050 461.400 ;
        RECT 607.950 459.600 610.050 460.050 ;
        RECT 566.400 458.400 610.050 459.600 ;
        RECT 268.950 455.400 280.050 456.600 ;
        RECT 268.950 454.950 271.050 455.400 ;
        RECT 277.950 454.950 280.050 455.400 ;
        RECT 290.400 455.400 315.600 456.600 ;
        RECT 191.400 452.400 196.050 453.600 ;
        RECT 193.950 451.950 196.050 452.400 ;
        RECT 206.400 452.400 210.600 453.600 ;
        RECT 214.950 453.600 217.050 454.050 ;
        RECT 230.400 453.600 231.600 454.950 ;
        RECT 214.950 452.400 231.600 453.600 ;
        RECT 232.950 453.600 235.050 454.050 ;
        RECT 244.950 453.600 247.050 454.050 ;
        RECT 232.950 452.400 247.050 453.600 ;
        RECT 115.950 448.950 118.050 451.050 ;
        RECT 127.950 450.600 130.050 451.050 ;
        RECT 166.950 450.600 169.050 451.050 ;
        RECT 127.950 449.400 169.050 450.600 ;
        RECT 127.950 448.950 130.050 449.400 ;
        RECT 166.950 448.950 169.050 449.400 ;
        RECT 170.400 448.050 171.600 451.950 ;
        RECT 206.400 451.050 207.600 452.400 ;
        RECT 214.950 451.950 217.050 452.400 ;
        RECT 232.950 451.950 235.050 452.400 ;
        RECT 244.950 451.950 247.050 452.400 ;
        RECT 248.400 451.050 249.600 454.950 ;
        RECT 290.400 454.050 291.600 455.400 ;
        RECT 316.950 454.950 319.050 457.050 ;
        RECT 328.950 454.950 331.050 457.050 ;
        RECT 331.950 456.600 334.050 457.050 ;
        RECT 352.950 456.600 355.050 457.050 ;
        RECT 424.950 456.600 427.050 457.050 ;
        RECT 331.950 455.400 355.050 456.600 ;
        RECT 331.950 454.950 334.050 455.400 ;
        RECT 352.950 454.950 355.050 455.400 ;
        RECT 416.400 455.400 427.050 456.600 ;
        RECT 289.950 451.950 292.050 454.050 ;
        RECT 292.950 453.600 295.050 454.050 ;
        RECT 298.950 453.600 301.050 454.050 ;
        RECT 292.950 452.400 301.050 453.600 ;
        RECT 292.950 451.950 295.050 452.400 ;
        RECT 298.950 451.950 301.050 452.400 ;
        RECT 310.950 453.600 313.050 454.050 ;
        RECT 317.400 453.600 318.600 454.950 ;
        RECT 310.950 452.400 318.600 453.600 ;
        RECT 310.950 451.950 313.050 452.400 ;
        RECT 329.400 451.050 330.600 454.950 ;
        RECT 416.400 454.050 417.600 455.400 ;
        RECT 424.950 454.950 427.050 455.400 ;
        RECT 463.950 456.600 466.050 457.050 ;
        RECT 472.950 456.600 475.050 457.050 ;
        RECT 511.950 456.600 514.050 457.050 ;
        RECT 463.950 455.400 475.050 456.600 ;
        RECT 463.950 454.950 466.050 455.400 ;
        RECT 472.950 454.950 475.050 455.400 ;
        RECT 488.400 455.400 514.050 456.600 ;
        RECT 361.950 453.600 364.050 454.050 ;
        RECT 373.950 453.600 376.050 454.050 ;
        RECT 361.950 452.400 376.050 453.600 ;
        RECT 361.950 451.950 364.050 452.400 ;
        RECT 373.950 451.950 376.050 452.400 ;
        RECT 415.950 451.950 418.050 454.050 ;
        RECT 421.950 453.600 424.050 454.050 ;
        RECT 472.950 453.600 475.050 454.050 ;
        RECT 484.950 453.600 487.050 454.050 ;
        RECT 421.950 452.400 441.600 453.600 ;
        RECT 421.950 451.950 424.050 452.400 ;
        RECT 205.950 448.950 208.050 451.050 ;
        RECT 247.950 448.950 250.050 451.050 ;
        RECT 328.950 448.950 331.050 451.050 ;
        RECT 340.950 450.600 343.050 451.050 ;
        RECT 352.950 450.600 355.050 451.050 ;
        RECT 340.950 449.400 355.050 450.600 ;
        RECT 340.950 448.950 343.050 449.400 ;
        RECT 352.950 448.950 355.050 449.400 ;
        RECT 382.950 450.600 385.050 451.050 ;
        RECT 436.950 450.600 439.050 451.050 ;
        RECT 382.950 449.400 439.050 450.600 ;
        RECT 440.400 450.600 441.600 452.400 ;
        RECT 461.400 452.400 475.050 453.600 ;
        RECT 461.400 450.600 462.600 452.400 ;
        RECT 472.950 451.950 475.050 452.400 ;
        RECT 476.400 452.400 487.050 453.600 ;
        RECT 440.400 449.400 462.600 450.600 ;
        RECT 469.950 450.600 472.050 451.050 ;
        RECT 476.400 450.600 477.600 452.400 ;
        RECT 484.950 451.950 487.050 452.400 ;
        RECT 488.400 451.050 489.600 455.400 ;
        RECT 511.950 454.950 514.050 455.400 ;
        RECT 529.950 456.600 532.050 457.050 ;
        RECT 529.950 455.400 543.600 456.600 ;
        RECT 529.950 454.950 532.050 455.400 ;
        RECT 542.400 454.050 543.600 455.400 ;
        RECT 496.950 453.600 499.050 454.050 ;
        RECT 491.400 452.400 499.050 453.600 ;
        RECT 469.950 449.400 477.600 450.600 ;
        RECT 382.950 448.950 385.050 449.400 ;
        RECT 436.950 448.950 439.050 449.400 ;
        RECT 469.950 448.950 472.050 449.400 ;
        RECT 487.950 448.950 490.050 451.050 ;
        RECT 148.950 447.600 151.050 448.050 ;
        RECT 113.400 446.400 151.050 447.600 ;
        RECT 148.950 445.950 151.050 446.400 ;
        RECT 169.950 445.950 172.050 448.050 ;
        RECT 178.950 447.600 181.050 448.050 ;
        RECT 214.950 447.600 217.050 448.050 ;
        RECT 178.950 446.400 217.050 447.600 ;
        RECT 178.950 445.950 181.050 446.400 ;
        RECT 214.950 445.950 217.050 446.400 ;
        RECT 226.950 447.600 229.050 448.050 ;
        RECT 307.950 447.600 310.050 448.050 ;
        RECT 226.950 446.400 310.050 447.600 ;
        RECT 226.950 445.950 229.050 446.400 ;
        RECT 307.950 445.950 310.050 446.400 ;
        RECT 325.950 447.600 328.050 448.050 ;
        RECT 331.950 447.600 334.050 448.050 ;
        RECT 325.950 446.400 334.050 447.600 ;
        RECT 325.950 445.950 328.050 446.400 ;
        RECT 331.950 445.950 334.050 446.400 ;
        RECT 340.950 447.600 343.050 448.050 ;
        RECT 346.950 447.600 349.050 448.050 ;
        RECT 367.950 447.600 370.050 448.050 ;
        RECT 340.950 446.400 370.050 447.600 ;
        RECT 340.950 445.950 343.050 446.400 ;
        RECT 346.950 445.950 349.050 446.400 ;
        RECT 367.950 445.950 370.050 446.400 ;
        RECT 385.950 447.600 388.050 448.050 ;
        RECT 397.950 447.600 400.050 448.050 ;
        RECT 385.950 446.400 400.050 447.600 ;
        RECT 385.950 445.950 388.050 446.400 ;
        RECT 397.950 445.950 400.050 446.400 ;
        RECT 409.950 447.600 412.050 448.050 ;
        RECT 454.950 447.600 457.050 448.050 ;
        RECT 409.950 446.400 457.050 447.600 ;
        RECT 409.950 445.950 412.050 446.400 ;
        RECT 454.950 445.950 457.050 446.400 ;
        RECT 481.950 447.600 484.050 448.050 ;
        RECT 491.400 447.600 492.600 452.400 ;
        RECT 496.950 451.950 499.050 452.400 ;
        RECT 508.950 451.950 511.050 454.050 ;
        RECT 523.950 453.600 526.050 454.050 ;
        RECT 538.950 453.600 541.050 454.050 ;
        RECT 523.950 452.400 541.050 453.600 ;
        RECT 523.950 451.950 526.050 452.400 ;
        RECT 538.950 451.950 541.050 452.400 ;
        RECT 541.950 451.950 544.050 454.050 ;
        RECT 493.950 450.600 496.050 451.050 ;
        RECT 509.400 450.600 510.600 451.950 ;
        RECT 520.950 450.600 523.050 451.050 ;
        RECT 493.950 449.400 523.050 450.600 ;
        RECT 493.950 448.950 496.050 449.400 ;
        RECT 520.950 448.950 523.050 449.400 ;
        RECT 526.950 450.600 529.050 451.050 ;
        RECT 535.950 450.600 538.050 451.050 ;
        RECT 526.950 449.400 538.050 450.600 ;
        RECT 526.950 448.950 529.050 449.400 ;
        RECT 535.950 448.950 538.050 449.400 ;
        RECT 538.950 450.600 541.050 451.050 ;
        RECT 545.400 450.600 546.600 457.950 ;
        RECT 538.950 449.400 546.600 450.600 ;
        RECT 553.950 450.600 556.050 451.050 ;
        RECT 563.400 450.600 564.600 457.950 ;
        RECT 575.400 454.050 576.600 458.400 ;
        RECT 607.950 457.950 610.050 458.400 ;
        RECT 610.950 459.600 613.050 460.050 ;
        RECT 622.950 459.600 625.050 460.050 ;
        RECT 610.950 458.400 625.050 459.600 ;
        RECT 610.950 457.950 613.050 458.400 ;
        RECT 622.950 457.950 625.050 458.400 ;
        RECT 625.950 459.600 628.050 460.050 ;
        RECT 637.950 459.600 640.050 460.050 ;
        RECT 625.950 458.400 640.050 459.600 ;
        RECT 625.950 457.950 628.050 458.400 ;
        RECT 637.950 457.950 640.050 458.400 ;
        RECT 658.950 457.950 661.050 460.050 ;
        RECT 664.950 459.600 667.050 460.050 ;
        RECT 685.950 459.600 688.050 460.050 ;
        RECT 664.950 458.400 688.050 459.600 ;
        RECT 664.950 457.950 667.050 458.400 ;
        RECT 685.950 457.950 688.050 458.400 ;
        RECT 694.950 457.950 697.050 460.050 ;
        RECT 709.950 459.600 712.050 460.050 ;
        RECT 724.950 459.600 727.050 460.050 ;
        RECT 760.950 459.600 763.050 460.050 ;
        RECT 709.950 458.400 727.050 459.600 ;
        RECT 709.950 457.950 712.050 458.400 ;
        RECT 724.950 457.950 727.050 458.400 ;
        RECT 740.400 458.400 763.050 459.600 ;
        RECT 577.950 456.600 580.050 457.050 ;
        RECT 583.950 456.600 586.050 457.050 ;
        RECT 577.950 455.400 586.050 456.600 ;
        RECT 577.950 454.950 580.050 455.400 ;
        RECT 583.950 454.950 586.050 455.400 ;
        RECT 592.950 454.950 595.050 457.050 ;
        RECT 595.950 456.600 598.050 457.050 ;
        RECT 604.950 456.600 607.050 457.050 ;
        RECT 628.950 456.600 631.050 457.050 ;
        RECT 595.950 455.400 607.050 456.600 ;
        RECT 595.950 454.950 598.050 455.400 ;
        RECT 604.950 454.950 607.050 455.400 ;
        RECT 614.400 455.400 631.050 456.600 ;
        RECT 574.950 451.950 577.050 454.050 ;
        RECT 580.950 451.950 583.050 454.050 ;
        RECT 593.400 453.600 594.600 454.950 ;
        RECT 614.400 454.050 615.600 455.400 ;
        RECT 628.950 454.950 631.050 455.400 ;
        RECT 634.950 456.600 637.050 457.050 ;
        RECT 646.950 456.600 649.050 457.050 ;
        RECT 634.950 455.400 649.050 456.600 ;
        RECT 634.950 454.950 637.050 455.400 ;
        RECT 646.950 454.950 649.050 455.400 ;
        RECT 601.950 453.600 604.050 454.050 ;
        RECT 610.950 453.600 613.050 454.050 ;
        RECT 593.400 452.400 597.600 453.600 ;
        RECT 581.400 450.600 582.600 451.950 ;
        RECT 592.950 450.600 595.050 451.050 ;
        RECT 553.950 449.400 595.050 450.600 ;
        RECT 538.950 448.950 541.050 449.400 ;
        RECT 553.950 448.950 556.050 449.400 ;
        RECT 592.950 448.950 595.050 449.400 ;
        RECT 481.950 446.400 492.600 447.600 ;
        RECT 499.950 447.600 502.050 448.050 ;
        RECT 517.950 447.600 520.050 448.050 ;
        RECT 544.950 447.600 547.050 448.050 ;
        RECT 499.950 446.400 547.050 447.600 ;
        RECT 481.950 445.950 484.050 446.400 ;
        RECT 499.950 445.950 502.050 446.400 ;
        RECT 517.950 445.950 520.050 446.400 ;
        RECT 544.950 445.950 547.050 446.400 ;
        RECT 574.950 447.600 577.050 448.050 ;
        RECT 596.400 447.600 597.600 452.400 ;
        RECT 601.950 452.400 613.050 453.600 ;
        RECT 601.950 451.950 604.050 452.400 ;
        RECT 610.950 451.950 613.050 452.400 ;
        RECT 613.950 451.950 616.050 454.050 ;
        RECT 635.400 453.600 636.600 454.950 ;
        RECT 649.950 453.600 652.050 454.050 ;
        RECT 659.400 453.600 660.600 457.950 ;
        RECT 670.950 456.600 673.050 457.050 ;
        RECT 679.950 456.600 682.050 457.050 ;
        RECT 670.950 455.400 682.050 456.600 ;
        RECT 695.400 456.600 696.600 457.950 ;
        RECT 709.950 456.600 712.050 457.050 ;
        RECT 740.400 456.600 741.600 458.400 ;
        RECT 760.950 457.950 763.050 458.400 ;
        RECT 748.950 456.600 751.050 457.050 ;
        RECT 695.400 455.400 699.600 456.600 ;
        RECT 670.950 454.950 673.050 455.400 ;
        RECT 679.950 454.950 682.050 455.400 ;
        RECT 698.400 454.050 699.600 455.400 ;
        RECT 704.400 455.400 712.050 456.600 ;
        RECT 704.400 454.050 705.600 455.400 ;
        RECT 709.950 454.950 712.050 455.400 ;
        RECT 731.400 455.400 741.600 456.600 ;
        RECT 743.400 455.400 751.050 456.600 ;
        RECT 679.950 453.600 682.050 454.050 ;
        RECT 635.400 452.400 645.600 453.600 ;
        RECT 607.950 450.600 610.050 451.050 ;
        RECT 619.950 450.600 622.050 451.050 ;
        RECT 607.950 449.400 622.050 450.600 ;
        RECT 607.950 448.950 610.050 449.400 ;
        RECT 619.950 448.950 622.050 449.400 ;
        RECT 625.950 450.600 628.050 451.050 ;
        RECT 640.950 450.600 643.050 451.050 ;
        RECT 625.950 449.400 643.050 450.600 ;
        RECT 644.400 450.600 645.600 452.400 ;
        RECT 649.950 452.400 660.600 453.600 ;
        RECT 665.400 452.400 682.050 453.600 ;
        RECT 649.950 451.950 652.050 452.400 ;
        RECT 665.400 451.050 666.600 452.400 ;
        RECT 679.950 451.950 682.050 452.400 ;
        RECT 682.950 453.600 685.050 454.050 ;
        RECT 694.950 453.600 697.050 454.050 ;
        RECT 682.950 452.400 697.050 453.600 ;
        RECT 682.950 451.950 685.050 452.400 ;
        RECT 694.950 451.950 697.050 452.400 ;
        RECT 697.950 451.950 700.050 454.050 ;
        RECT 703.950 451.950 706.050 454.050 ;
        RECT 706.950 453.600 709.050 454.050 ;
        RECT 715.950 453.600 718.050 454.050 ;
        RECT 706.950 452.400 718.050 453.600 ;
        RECT 706.950 451.950 709.050 452.400 ;
        RECT 715.950 451.950 718.050 452.400 ;
        RECT 727.950 453.600 730.050 454.050 ;
        RECT 731.400 453.600 732.600 455.400 ;
        RECT 727.950 452.400 732.600 453.600 ;
        RECT 733.950 453.600 736.050 454.050 ;
        RECT 743.400 453.600 744.600 455.400 ;
        RECT 748.950 454.950 751.050 455.400 ;
        RECT 754.950 456.600 757.050 457.050 ;
        RECT 766.950 456.600 769.050 457.050 ;
        RECT 754.950 455.400 765.600 456.600 ;
        RECT 754.950 454.950 757.050 455.400 ;
        RECT 757.950 453.600 760.050 454.050 ;
        RECT 733.950 452.400 744.600 453.600 ;
        RECT 746.400 452.400 760.050 453.600 ;
        RECT 764.400 453.600 765.600 455.400 ;
        RECT 766.950 455.400 771.600 456.600 ;
        RECT 766.950 454.950 769.050 455.400 ;
        RECT 766.950 453.600 769.050 454.050 ;
        RECT 764.400 452.400 769.050 453.600 ;
        RECT 727.950 451.950 730.050 452.400 ;
        RECT 733.950 451.950 736.050 452.400 ;
        RECT 646.950 450.600 649.050 451.050 ;
        RECT 644.400 449.400 649.050 450.600 ;
        RECT 625.950 448.950 628.050 449.400 ;
        RECT 640.950 448.950 643.050 449.400 ;
        RECT 646.950 448.950 649.050 449.400 ;
        RECT 664.950 448.950 667.050 451.050 ;
        RECT 673.950 450.600 676.050 451.050 ;
        RECT 691.950 450.600 694.050 451.050 ;
        RECT 746.400 450.600 747.600 452.400 ;
        RECT 757.950 451.950 760.050 452.400 ;
        RECT 766.950 451.950 769.050 452.400 ;
        RECT 673.950 449.400 681.600 450.600 ;
        RECT 673.950 448.950 676.050 449.400 ;
        RECT 574.950 446.400 597.600 447.600 ;
        RECT 604.950 447.600 607.050 448.050 ;
        RECT 616.950 447.600 619.050 448.050 ;
        RECT 676.950 447.600 679.050 448.050 ;
        RECT 604.950 446.400 679.050 447.600 ;
        RECT 574.950 445.950 577.050 446.400 ;
        RECT 604.950 445.950 607.050 446.400 ;
        RECT 616.950 445.950 619.050 446.400 ;
        RECT 676.950 445.950 679.050 446.400 ;
        RECT 148.950 444.600 151.050 445.050 ;
        RECT 295.950 444.600 298.050 445.050 ;
        RECT 148.950 443.400 298.050 444.600 ;
        RECT 148.950 442.950 151.050 443.400 ;
        RECT 295.950 442.950 298.050 443.400 ;
        RECT 301.950 444.600 304.050 445.050 ;
        RECT 334.950 444.600 337.050 445.050 ;
        RECT 301.950 443.400 337.050 444.600 ;
        RECT 301.950 442.950 304.050 443.400 ;
        RECT 334.950 442.950 337.050 443.400 ;
        RECT 400.950 444.600 403.050 445.050 ;
        RECT 463.950 444.600 466.050 445.050 ;
        RECT 400.950 443.400 466.050 444.600 ;
        RECT 400.950 442.950 403.050 443.400 ;
        RECT 463.950 442.950 466.050 443.400 ;
        RECT 475.950 444.600 478.050 445.050 ;
        RECT 511.950 444.600 514.050 445.050 ;
        RECT 475.950 443.400 514.050 444.600 ;
        RECT 475.950 442.950 478.050 443.400 ;
        RECT 511.950 442.950 514.050 443.400 ;
        RECT 535.950 444.600 538.050 445.050 ;
        RECT 553.950 444.600 556.050 445.050 ;
        RECT 535.950 443.400 556.050 444.600 ;
        RECT 535.950 442.950 538.050 443.400 ;
        RECT 553.950 442.950 556.050 443.400 ;
        RECT 559.950 444.600 562.050 445.050 ;
        RECT 607.950 444.600 610.050 445.050 ;
        RECT 559.950 443.400 610.050 444.600 ;
        RECT 559.950 442.950 562.050 443.400 ;
        RECT 607.950 442.950 610.050 443.400 ;
        RECT 619.950 444.600 622.050 445.050 ;
        RECT 646.950 444.600 649.050 445.050 ;
        RECT 619.950 443.400 649.050 444.600 ;
        RECT 619.950 442.950 622.050 443.400 ;
        RECT 646.950 442.950 649.050 443.400 ;
        RECT 670.950 444.600 673.050 445.050 ;
        RECT 680.400 444.600 681.600 449.400 ;
        RECT 691.950 449.400 747.600 450.600 ;
        RECT 748.950 450.600 751.050 451.050 ;
        RECT 770.400 450.600 771.600 455.400 ;
        RECT 748.950 449.400 771.600 450.600 ;
        RECT 691.950 448.950 694.050 449.400 ;
        RECT 748.950 448.950 751.050 449.400 ;
        RECT 694.950 447.600 697.050 448.050 ;
        RECT 700.950 447.600 703.050 448.050 ;
        RECT 694.950 446.400 703.050 447.600 ;
        RECT 694.950 445.950 697.050 446.400 ;
        RECT 700.950 445.950 703.050 446.400 ;
        RECT 718.950 447.600 721.050 448.050 ;
        RECT 751.950 447.600 754.050 448.050 ;
        RECT 718.950 446.400 754.050 447.600 ;
        RECT 718.950 445.950 721.050 446.400 ;
        RECT 751.950 445.950 754.050 446.400 ;
        RECT 670.950 443.400 681.600 444.600 ;
        RECT 682.950 444.600 685.050 445.050 ;
        RECT 700.950 444.600 703.050 445.050 ;
        RECT 682.950 443.400 703.050 444.600 ;
        RECT 670.950 442.950 673.050 443.400 ;
        RECT 682.950 442.950 685.050 443.400 ;
        RECT 700.950 442.950 703.050 443.400 ;
        RECT 712.950 444.600 715.050 445.050 ;
        RECT 754.950 444.600 757.050 445.050 ;
        RECT 712.950 443.400 757.050 444.600 ;
        RECT 712.950 442.950 715.050 443.400 ;
        RECT 754.950 442.950 757.050 443.400 ;
        RECT 79.950 441.600 82.050 442.050 ;
        RECT 94.950 441.600 97.050 442.050 ;
        RECT 175.950 441.600 178.050 442.050 ;
        RECT 79.950 440.400 178.050 441.600 ;
        RECT 79.950 439.950 82.050 440.400 ;
        RECT 94.950 439.950 97.050 440.400 ;
        RECT 175.950 439.950 178.050 440.400 ;
        RECT 241.950 441.600 244.050 442.050 ;
        RECT 256.950 441.600 259.050 442.050 ;
        RECT 241.950 440.400 259.050 441.600 ;
        RECT 241.950 439.950 244.050 440.400 ;
        RECT 256.950 439.950 259.050 440.400 ;
        RECT 283.950 441.600 286.050 442.050 ;
        RECT 451.950 441.600 454.050 442.050 ;
        RECT 460.950 441.600 463.050 442.050 ;
        RECT 283.950 440.400 324.600 441.600 ;
        RECT 283.950 439.950 286.050 440.400 ;
        RECT 193.950 438.600 196.050 439.050 ;
        RECT 253.950 438.600 256.050 439.050 ;
        RECT 193.950 437.400 256.050 438.600 ;
        RECT 323.400 438.600 324.600 440.400 ;
        RECT 451.950 440.400 463.050 441.600 ;
        RECT 451.950 439.950 454.050 440.400 ;
        RECT 460.950 439.950 463.050 440.400 ;
        RECT 493.950 441.600 496.050 442.050 ;
        RECT 661.950 441.600 664.050 442.050 ;
        RECT 493.950 440.400 664.050 441.600 ;
        RECT 493.950 439.950 496.050 440.400 ;
        RECT 661.950 439.950 664.050 440.400 ;
        RECT 664.950 441.600 667.050 442.050 ;
        RECT 688.950 441.600 691.050 442.050 ;
        RECT 664.950 440.400 691.050 441.600 ;
        RECT 664.950 439.950 667.050 440.400 ;
        RECT 688.950 439.950 691.050 440.400 ;
        RECT 706.950 441.600 709.050 442.050 ;
        RECT 760.950 441.600 763.050 442.050 ;
        RECT 706.950 440.400 763.050 441.600 ;
        RECT 706.950 439.950 709.050 440.400 ;
        RECT 760.950 439.950 763.050 440.400 ;
        RECT 445.950 438.600 448.050 439.050 ;
        RECT 323.400 437.400 448.050 438.600 ;
        RECT 193.950 436.950 196.050 437.400 ;
        RECT 253.950 436.950 256.050 437.400 ;
        RECT 445.950 436.950 448.050 437.400 ;
        RECT 520.950 438.600 523.050 439.050 ;
        RECT 586.950 438.600 589.050 439.050 ;
        RECT 520.950 437.400 589.050 438.600 ;
        RECT 520.950 436.950 523.050 437.400 ;
        RECT 586.950 436.950 589.050 437.400 ;
        RECT 607.950 438.600 610.050 439.050 ;
        RECT 682.950 438.600 685.050 439.050 ;
        RECT 607.950 437.400 685.050 438.600 ;
        RECT 607.950 436.950 610.050 437.400 ;
        RECT 682.950 436.950 685.050 437.400 ;
        RECT 688.950 438.600 691.050 439.050 ;
        RECT 718.950 438.600 721.050 439.050 ;
        RECT 688.950 437.400 721.050 438.600 ;
        RECT 688.950 436.950 691.050 437.400 ;
        RECT 718.950 436.950 721.050 437.400 ;
        RECT 730.950 438.600 733.050 439.050 ;
        RECT 757.950 438.600 760.050 439.050 ;
        RECT 730.950 437.400 760.050 438.600 ;
        RECT 730.950 436.950 733.050 437.400 ;
        RECT 757.950 436.950 760.050 437.400 ;
        RECT 43.950 435.600 46.050 436.050 ;
        RECT 70.950 435.600 73.050 436.050 ;
        RECT 43.950 434.400 73.050 435.600 ;
        RECT 43.950 433.950 46.050 434.400 ;
        RECT 70.950 433.950 73.050 434.400 ;
        RECT 160.950 435.600 163.050 436.050 ;
        RECT 199.950 435.600 202.050 436.050 ;
        RECT 160.950 434.400 202.050 435.600 ;
        RECT 160.950 433.950 163.050 434.400 ;
        RECT 199.950 433.950 202.050 434.400 ;
        RECT 238.950 435.600 241.050 436.050 ;
        RECT 253.950 435.600 256.050 436.050 ;
        RECT 238.950 434.400 256.050 435.600 ;
        RECT 238.950 433.950 241.050 434.400 ;
        RECT 253.950 433.950 256.050 434.400 ;
        RECT 439.950 435.600 442.050 436.050 ;
        RECT 568.950 435.600 571.050 436.050 ;
        RECT 439.950 434.400 571.050 435.600 ;
        RECT 439.950 433.950 442.050 434.400 ;
        RECT 568.950 433.950 571.050 434.400 ;
        RECT 580.950 435.600 583.050 436.050 ;
        RECT 619.950 435.600 622.050 436.050 ;
        RECT 580.950 434.400 622.050 435.600 ;
        RECT 580.950 433.950 583.050 434.400 ;
        RECT 619.950 433.950 622.050 434.400 ;
        RECT 622.950 435.600 625.050 436.050 ;
        RECT 643.950 435.600 646.050 436.050 ;
        RECT 622.950 434.400 646.050 435.600 ;
        RECT 622.950 433.950 625.050 434.400 ;
        RECT 643.950 433.950 646.050 434.400 ;
        RECT 649.950 435.600 652.050 436.050 ;
        RECT 676.950 435.600 679.050 436.050 ;
        RECT 649.950 434.400 679.050 435.600 ;
        RECT 649.950 433.950 652.050 434.400 ;
        RECT 676.950 433.950 679.050 434.400 ;
        RECT 685.950 435.600 688.050 436.050 ;
        RECT 697.950 435.600 700.050 436.050 ;
        RECT 685.950 434.400 700.050 435.600 ;
        RECT 685.950 433.950 688.050 434.400 ;
        RECT 697.950 433.950 700.050 434.400 ;
        RECT 712.950 435.600 715.050 436.050 ;
        RECT 733.950 435.600 736.050 436.050 ;
        RECT 712.950 434.400 736.050 435.600 ;
        RECT 712.950 433.950 715.050 434.400 ;
        RECT 733.950 433.950 736.050 434.400 ;
        RECT 739.950 435.600 742.050 436.050 ;
        RECT 748.950 435.600 751.050 436.050 ;
        RECT 739.950 434.400 751.050 435.600 ;
        RECT 739.950 433.950 742.050 434.400 ;
        RECT 748.950 433.950 751.050 434.400 ;
        RECT 25.950 432.600 28.050 433.050 ;
        RECT 157.950 432.600 160.050 433.050 ;
        RECT 25.950 431.400 160.050 432.600 ;
        RECT 25.950 430.950 28.050 431.400 ;
        RECT 157.950 430.950 160.050 431.400 ;
        RECT 169.950 432.600 172.050 433.050 ;
        RECT 238.950 432.600 241.050 433.050 ;
        RECT 280.950 432.600 283.050 433.050 ;
        RECT 169.950 431.400 241.050 432.600 ;
        RECT 169.950 430.950 172.050 431.400 ;
        RECT 238.950 430.950 241.050 431.400 ;
        RECT 257.400 431.400 283.050 432.600 ;
        RECT 37.950 429.600 40.050 430.050 ;
        RECT 151.950 429.600 154.050 430.050 ;
        RECT 37.950 428.400 154.050 429.600 ;
        RECT 37.950 427.950 40.050 428.400 ;
        RECT 151.950 427.950 154.050 428.400 ;
        RECT 223.950 429.600 226.050 430.050 ;
        RECT 257.400 429.600 258.600 431.400 ;
        RECT 280.950 430.950 283.050 431.400 ;
        RECT 286.950 432.600 289.050 433.050 ;
        RECT 319.950 432.600 322.050 433.050 ;
        RECT 286.950 431.400 322.050 432.600 ;
        RECT 286.950 430.950 289.050 431.400 ;
        RECT 319.950 430.950 322.050 431.400 ;
        RECT 334.950 432.600 337.050 433.050 ;
        RECT 349.950 432.600 352.050 433.050 ;
        RECT 334.950 431.400 352.050 432.600 ;
        RECT 334.950 430.950 337.050 431.400 ;
        RECT 349.950 430.950 352.050 431.400 ;
        RECT 352.950 432.600 355.050 433.050 ;
        RECT 430.950 432.600 433.050 433.050 ;
        RECT 352.950 431.400 433.050 432.600 ;
        RECT 352.950 430.950 355.050 431.400 ;
        RECT 430.950 430.950 433.050 431.400 ;
        RECT 490.950 432.600 493.050 433.050 ;
        RECT 499.950 432.600 502.050 433.050 ;
        RECT 631.950 432.600 634.050 433.050 ;
        RECT 490.950 431.400 634.050 432.600 ;
        RECT 490.950 430.950 493.050 431.400 ;
        RECT 499.950 430.950 502.050 431.400 ;
        RECT 631.950 430.950 634.050 431.400 ;
        RECT 646.950 432.600 649.050 433.050 ;
        RECT 691.950 432.600 694.050 433.050 ;
        RECT 646.950 431.400 694.050 432.600 ;
        RECT 646.950 430.950 649.050 431.400 ;
        RECT 691.950 430.950 694.050 431.400 ;
        RECT 703.950 432.600 706.050 433.050 ;
        RECT 715.950 432.600 718.050 433.050 ;
        RECT 703.950 431.400 718.050 432.600 ;
        RECT 703.950 430.950 706.050 431.400 ;
        RECT 715.950 430.950 718.050 431.400 ;
        RECT 727.950 432.600 730.050 433.050 ;
        RECT 751.950 432.600 754.050 433.050 ;
        RECT 727.950 431.400 754.050 432.600 ;
        RECT 727.950 430.950 730.050 431.400 ;
        RECT 751.950 430.950 754.050 431.400 ;
        RECT 223.950 428.400 258.600 429.600 ;
        RECT 259.950 429.600 262.050 430.050 ;
        RECT 277.950 429.600 280.050 430.050 ;
        RECT 301.950 429.600 304.050 430.050 ;
        RECT 259.950 428.400 304.050 429.600 ;
        RECT 223.950 427.950 226.050 428.400 ;
        RECT 259.950 427.950 262.050 428.400 ;
        RECT 277.950 427.950 280.050 428.400 ;
        RECT 301.950 427.950 304.050 428.400 ;
        RECT 307.950 429.600 310.050 430.050 ;
        RECT 343.950 429.600 346.050 430.050 ;
        RECT 307.950 428.400 346.050 429.600 ;
        RECT 307.950 427.950 310.050 428.400 ;
        RECT 343.950 427.950 346.050 428.400 ;
        RECT 370.950 429.600 373.050 430.050 ;
        RECT 376.950 429.600 379.050 430.050 ;
        RECT 370.950 428.400 379.050 429.600 ;
        RECT 370.950 427.950 373.050 428.400 ;
        RECT 376.950 427.950 379.050 428.400 ;
        RECT 379.950 429.600 382.050 430.050 ;
        RECT 430.950 429.600 433.050 430.050 ;
        RECT 379.950 428.400 433.050 429.600 ;
        RECT 379.950 427.950 382.050 428.400 ;
        RECT 430.950 427.950 433.050 428.400 ;
        RECT 445.950 429.600 448.050 430.050 ;
        RECT 538.950 429.600 541.050 430.050 ;
        RECT 445.950 428.400 541.050 429.600 ;
        RECT 445.950 427.950 448.050 428.400 ;
        RECT 538.950 427.950 541.050 428.400 ;
        RECT 556.950 429.600 559.050 430.050 ;
        RECT 580.950 429.600 583.050 430.050 ;
        RECT 556.950 428.400 583.050 429.600 ;
        RECT 556.950 427.950 559.050 428.400 ;
        RECT 580.950 427.950 583.050 428.400 ;
        RECT 637.950 429.600 640.050 430.050 ;
        RECT 703.950 429.600 706.050 430.050 ;
        RECT 637.950 428.400 706.050 429.600 ;
        RECT 637.950 427.950 640.050 428.400 ;
        RECT 703.950 427.950 706.050 428.400 ;
        RECT 52.950 426.600 55.050 427.050 ;
        RECT 169.950 426.600 172.050 427.050 ;
        RECT 52.950 425.400 172.050 426.600 ;
        RECT 52.950 424.950 55.050 425.400 ;
        RECT 169.950 424.950 172.050 425.400 ;
        RECT 307.950 426.600 310.050 427.050 ;
        RECT 358.950 426.600 361.050 427.050 ;
        RECT 307.950 425.400 361.050 426.600 ;
        RECT 307.950 424.950 310.050 425.400 ;
        RECT 358.950 424.950 361.050 425.400 ;
        RECT 478.950 426.600 481.050 427.050 ;
        RECT 589.950 426.600 592.050 427.050 ;
        RECT 478.950 425.400 592.050 426.600 ;
        RECT 478.950 424.950 481.050 425.400 ;
        RECT 589.950 424.950 592.050 425.400 ;
        RECT 592.950 426.600 595.050 427.050 ;
        RECT 679.950 426.600 682.050 427.050 ;
        RECT 592.950 425.400 682.050 426.600 ;
        RECT 592.950 424.950 595.050 425.400 ;
        RECT 679.950 424.950 682.050 425.400 ;
        RECT 700.950 426.600 703.050 427.050 ;
        RECT 718.950 426.600 721.050 427.050 ;
        RECT 700.950 425.400 721.050 426.600 ;
        RECT 700.950 424.950 703.050 425.400 ;
        RECT 718.950 424.950 721.050 425.400 ;
        RECT 721.950 426.600 724.050 427.050 ;
        RECT 748.950 426.600 751.050 427.050 ;
        RECT 721.950 425.400 751.050 426.600 ;
        RECT 721.950 424.950 724.050 425.400 ;
        RECT 748.950 424.950 751.050 425.400 ;
        RECT 10.950 423.600 13.050 424.050 ;
        RECT 76.950 423.600 79.050 424.050 ;
        RECT 10.950 422.400 79.050 423.600 ;
        RECT 10.950 421.950 13.050 422.400 ;
        RECT 52.950 418.950 55.050 421.050 ;
        RECT 64.950 418.950 67.050 421.050 ;
        RECT 43.950 417.600 46.050 418.050 ;
        RECT 14.400 416.400 46.050 417.600 ;
        RECT 14.400 415.050 15.600 416.400 ;
        RECT 43.950 415.950 46.050 416.400 ;
        RECT 53.400 415.050 54.600 418.950 ;
        RECT 55.950 417.600 58.050 418.050 ;
        RECT 58.950 417.600 61.050 418.050 ;
        RECT 61.950 417.600 64.050 418.050 ;
        RECT 55.950 416.400 64.050 417.600 ;
        RECT 55.950 415.950 58.050 416.400 ;
        RECT 58.950 415.950 61.050 416.400 ;
        RECT 61.950 415.950 64.050 416.400 ;
        RECT 65.400 415.050 66.600 418.950 ;
        RECT 71.400 415.050 72.600 422.400 ;
        RECT 76.950 421.950 79.050 422.400 ;
        RECT 169.950 423.600 172.050 424.050 ;
        RECT 193.950 423.600 196.050 424.050 ;
        RECT 169.950 422.400 196.050 423.600 ;
        RECT 169.950 421.950 172.050 422.400 ;
        RECT 193.950 421.950 196.050 422.400 ;
        RECT 229.950 423.600 232.050 424.050 ;
        RECT 268.950 423.600 271.050 424.050 ;
        RECT 229.950 422.400 271.050 423.600 ;
        RECT 229.950 421.950 232.050 422.400 ;
        RECT 268.950 421.950 271.050 422.400 ;
        RECT 298.950 423.600 301.050 424.050 ;
        RECT 400.950 423.600 403.050 424.050 ;
        RECT 298.950 422.400 403.050 423.600 ;
        RECT 298.950 421.950 301.050 422.400 ;
        RECT 400.950 421.950 403.050 422.400 ;
        RECT 457.950 423.600 460.050 424.050 ;
        RECT 469.950 423.600 472.050 424.050 ;
        RECT 457.950 422.400 472.050 423.600 ;
        RECT 457.950 421.950 460.050 422.400 ;
        RECT 469.950 421.950 472.050 422.400 ;
        RECT 475.950 423.600 478.050 424.050 ;
        RECT 496.950 423.600 499.050 424.050 ;
        RECT 475.950 422.400 499.050 423.600 ;
        RECT 475.950 421.950 478.050 422.400 ;
        RECT 496.950 421.950 499.050 422.400 ;
        RECT 616.950 423.600 619.050 424.050 ;
        RECT 637.950 423.600 640.050 424.050 ;
        RECT 616.950 422.400 640.050 423.600 ;
        RECT 616.950 421.950 619.050 422.400 ;
        RECT 637.950 421.950 640.050 422.400 ;
        RECT 667.950 423.600 670.050 424.050 ;
        RECT 733.950 423.600 736.050 424.050 ;
        RECT 667.950 422.400 736.050 423.600 ;
        RECT 667.950 421.950 670.050 422.400 ;
        RECT 733.950 421.950 736.050 422.400 ;
        RECT 742.950 423.600 745.050 424.050 ;
        RECT 760.950 423.600 763.050 424.050 ;
        RECT 742.950 422.400 763.050 423.600 ;
        RECT 742.950 421.950 745.050 422.400 ;
        RECT 760.950 421.950 763.050 422.400 ;
        RECT 766.950 423.600 769.050 424.050 ;
        RECT 766.950 422.400 777.600 423.600 ;
        RECT 766.950 421.950 769.050 422.400 ;
        RECT 79.950 420.600 82.050 421.050 ;
        RECT 77.400 419.400 82.050 420.600 ;
        RECT 77.400 418.050 78.600 419.400 ;
        RECT 79.950 418.950 82.050 419.400 ;
        RECT 88.950 420.600 91.050 421.050 ;
        RECT 97.950 420.600 100.050 421.050 ;
        RECT 88.950 419.400 100.050 420.600 ;
        RECT 88.950 418.950 91.050 419.400 ;
        RECT 97.950 418.950 100.050 419.400 ;
        RECT 100.950 420.600 103.050 421.050 ;
        RECT 133.950 420.600 136.050 421.050 ;
        RECT 166.950 420.600 169.050 421.050 ;
        RECT 100.950 419.400 105.600 420.600 ;
        RECT 100.950 418.950 103.050 419.400 ;
        RECT 104.400 418.050 105.600 419.400 ;
        RECT 133.950 419.400 169.050 420.600 ;
        RECT 133.950 418.950 136.050 419.400 ;
        RECT 166.950 418.950 169.050 419.400 ;
        RECT 172.950 420.600 175.050 421.050 ;
        RECT 184.950 420.600 187.050 421.050 ;
        RECT 283.950 420.600 286.050 421.050 ;
        RECT 172.950 419.400 177.600 420.600 ;
        RECT 172.950 418.950 175.050 419.400 ;
        RECT 176.400 418.050 177.600 419.400 ;
        RECT 184.950 419.400 286.050 420.600 ;
        RECT 184.950 418.950 187.050 419.400 ;
        RECT 283.950 418.950 286.050 419.400 ;
        RECT 319.950 420.600 322.050 421.050 ;
        RECT 337.950 420.600 340.050 421.050 ;
        RECT 355.950 420.600 358.050 421.050 ;
        RECT 361.950 420.600 364.050 421.050 ;
        RECT 385.950 420.600 388.050 421.050 ;
        RECT 409.950 420.600 412.050 421.050 ;
        RECT 412.950 420.600 415.050 421.050 ;
        RECT 319.950 419.400 415.050 420.600 ;
        RECT 319.950 418.950 322.050 419.400 ;
        RECT 337.950 418.950 340.050 419.400 ;
        RECT 355.950 418.950 358.050 419.400 ;
        RECT 361.950 418.950 364.050 419.400 ;
        RECT 385.950 418.950 388.050 419.400 ;
        RECT 409.950 418.950 412.050 419.400 ;
        RECT 412.950 418.950 415.050 419.400 ;
        RECT 463.950 420.600 466.050 421.050 ;
        RECT 490.950 420.600 493.050 421.050 ;
        RECT 463.950 419.400 493.050 420.600 ;
        RECT 463.950 418.950 466.050 419.400 ;
        RECT 490.950 418.950 493.050 419.400 ;
        RECT 589.950 420.600 592.050 421.050 ;
        RECT 625.950 420.600 628.050 421.050 ;
        RECT 589.950 419.400 628.050 420.600 ;
        RECT 589.950 418.950 592.050 419.400 ;
        RECT 625.950 418.950 628.050 419.400 ;
        RECT 673.950 418.950 676.050 421.050 ;
        RECT 682.950 420.600 685.050 421.050 ;
        RECT 724.950 420.600 727.050 421.050 ;
        RECT 682.950 419.400 702.600 420.600 ;
        RECT 682.950 418.950 685.050 419.400 ;
        RECT 76.950 415.950 79.050 418.050 ;
        RECT 97.950 417.600 100.050 418.050 ;
        RECT 97.950 416.400 102.600 417.600 ;
        RECT 97.950 415.950 100.050 416.400 ;
        RECT 101.400 415.050 102.600 416.400 ;
        RECT 103.950 415.950 106.050 418.050 ;
        RECT 109.950 417.600 112.050 418.050 ;
        RECT 118.950 417.600 121.050 418.050 ;
        RECT 136.950 417.600 139.050 418.050 ;
        RECT 109.950 416.400 139.050 417.600 ;
        RECT 109.950 415.950 112.050 416.400 ;
        RECT 118.950 415.950 121.050 416.400 ;
        RECT 136.950 415.950 139.050 416.400 ;
        RECT 151.950 417.600 154.050 418.050 ;
        RECT 151.950 416.400 156.600 417.600 ;
        RECT 151.950 415.950 154.050 416.400 ;
        RECT 155.400 415.050 156.600 416.400 ;
        RECT 175.950 415.950 178.050 418.050 ;
        RECT 181.950 417.600 184.050 418.050 ;
        RECT 187.950 417.600 190.050 418.050 ;
        RECT 181.950 416.400 190.050 417.600 ;
        RECT 181.950 415.950 184.050 416.400 ;
        RECT 187.950 415.950 190.050 416.400 ;
        RECT 193.950 415.950 196.050 418.050 ;
        RECT 208.950 417.600 211.050 418.050 ;
        RECT 214.950 417.600 217.050 418.050 ;
        RECT 208.950 416.400 217.050 417.600 ;
        RECT 208.950 415.950 211.050 416.400 ;
        RECT 214.950 415.950 217.050 416.400 ;
        RECT 232.950 417.600 235.050 418.050 ;
        RECT 241.950 417.600 244.050 418.050 ;
        RECT 232.950 416.400 244.050 417.600 ;
        RECT 232.950 415.950 235.050 416.400 ;
        RECT 241.950 415.950 244.050 416.400 ;
        RECT 253.950 415.950 256.050 418.050 ;
        RECT 292.950 417.600 295.050 418.050 ;
        RECT 292.950 416.400 303.600 417.600 ;
        RECT 292.950 415.950 295.050 416.400 ;
        RECT 4.950 414.600 7.050 415.050 ;
        RECT 4.950 413.400 12.600 414.600 ;
        RECT 4.950 412.950 7.050 413.400 ;
        RECT 11.400 411.600 12.600 413.400 ;
        RECT 13.950 412.950 16.050 415.050 ;
        RECT 19.950 414.600 22.050 415.050 ;
        RECT 31.950 414.600 34.050 415.050 ;
        RECT 19.950 413.400 34.050 414.600 ;
        RECT 19.950 412.950 22.050 413.400 ;
        RECT 31.950 412.950 34.050 413.400 ;
        RECT 52.950 412.950 55.050 415.050 ;
        RECT 64.950 412.950 67.050 415.050 ;
        RECT 70.950 412.950 73.050 415.050 ;
        RECT 100.950 412.950 103.050 415.050 ;
        RECT 142.950 414.600 145.050 415.050 ;
        RECT 148.950 414.600 151.050 415.050 ;
        RECT 142.950 413.400 151.050 414.600 ;
        RECT 142.950 412.950 145.050 413.400 ;
        RECT 148.950 412.950 151.050 413.400 ;
        RECT 154.950 412.950 157.050 415.050 ;
        RECT 163.950 414.600 166.050 415.050 ;
        RECT 194.400 414.600 195.600 415.950 ;
        RECT 163.950 413.400 195.600 414.600 ;
        RECT 205.950 414.600 208.050 415.050 ;
        RECT 220.950 414.600 223.050 415.050 ;
        RECT 254.400 414.600 255.600 415.950 ;
        RECT 302.400 415.050 303.600 416.400 ;
        RECT 340.950 415.950 343.050 418.050 ;
        RECT 349.950 417.600 352.050 418.050 ;
        RECT 388.950 417.600 391.050 418.050 ;
        RECT 391.950 417.600 394.050 418.050 ;
        RECT 433.950 417.600 436.050 418.050 ;
        RECT 349.950 416.400 436.050 417.600 ;
        RECT 349.950 415.950 352.050 416.400 ;
        RECT 388.950 415.950 391.050 416.400 ;
        RECT 391.950 415.950 394.050 416.400 ;
        RECT 433.950 415.950 436.050 416.400 ;
        RECT 442.950 415.950 445.050 418.050 ;
        RECT 463.950 415.950 466.050 418.050 ;
        RECT 505.950 417.600 508.050 418.050 ;
        RECT 511.950 417.600 514.050 418.050 ;
        RECT 479.400 416.400 514.050 417.600 ;
        RECT 205.950 413.400 219.600 414.600 ;
        RECT 163.950 412.950 166.050 413.400 ;
        RECT 205.950 412.950 208.050 413.400 ;
        RECT 22.950 411.600 25.050 412.050 ;
        RECT 28.950 411.600 31.050 412.050 ;
        RECT 11.400 410.400 31.050 411.600 ;
        RECT 22.950 409.950 25.050 410.400 ;
        RECT 28.950 409.950 31.050 410.400 ;
        RECT 43.950 411.600 46.050 412.050 ;
        RECT 67.950 411.600 70.050 412.050 ;
        RECT 43.950 410.400 70.050 411.600 ;
        RECT 43.950 409.950 46.050 410.400 ;
        RECT 67.950 409.950 70.050 410.400 ;
        RECT 94.950 411.600 97.050 412.050 ;
        RECT 145.950 411.600 148.050 412.050 ;
        RECT 94.950 410.400 148.050 411.600 ;
        RECT 94.950 409.950 97.050 410.400 ;
        RECT 145.950 409.950 148.050 410.400 ;
        RECT 154.950 411.600 157.050 412.050 ;
        RECT 172.950 411.600 175.050 412.050 ;
        RECT 154.950 410.400 175.050 411.600 ;
        RECT 154.950 409.950 157.050 410.400 ;
        RECT 172.950 409.950 175.050 410.400 ;
        RECT 175.950 411.600 178.050 412.050 ;
        RECT 211.950 411.600 214.050 412.050 ;
        RECT 175.950 410.400 214.050 411.600 ;
        RECT 218.400 411.600 219.600 413.400 ;
        RECT 220.950 413.400 231.600 414.600 ;
        RECT 220.950 412.950 223.050 413.400 ;
        RECT 226.950 411.600 229.050 412.050 ;
        RECT 218.400 410.400 229.050 411.600 ;
        RECT 230.400 411.600 231.600 413.400 ;
        RECT 239.400 413.400 255.600 414.600 ;
        RECT 292.950 414.600 295.050 415.050 ;
        RECT 292.950 413.400 300.600 414.600 ;
        RECT 232.950 411.600 235.050 412.050 ;
        RECT 230.400 410.400 235.050 411.600 ;
        RECT 175.950 409.950 178.050 410.400 ;
        RECT 211.950 409.950 214.050 410.400 ;
        RECT 226.950 409.950 229.050 410.400 ;
        RECT 232.950 409.950 235.050 410.400 ;
        RECT 34.950 408.600 37.050 409.050 ;
        RECT 46.950 408.600 49.050 409.050 ;
        RECT 79.950 408.600 82.050 409.050 ;
        RECT 34.950 407.400 82.050 408.600 ;
        RECT 34.950 406.950 37.050 407.400 ;
        RECT 46.950 406.950 49.050 407.400 ;
        RECT 79.950 406.950 82.050 407.400 ;
        RECT 85.950 408.600 88.050 409.050 ;
        RECT 127.950 408.600 130.050 409.050 ;
        RECT 130.950 408.600 133.050 409.050 ;
        RECT 85.950 407.400 133.050 408.600 ;
        RECT 85.950 406.950 88.050 407.400 ;
        RECT 127.950 406.950 130.050 407.400 ;
        RECT 130.950 406.950 133.050 407.400 ;
        RECT 151.950 408.600 154.050 409.050 ;
        RECT 157.950 408.600 160.050 409.050 ;
        RECT 151.950 407.400 160.050 408.600 ;
        RECT 151.950 406.950 154.050 407.400 ;
        RECT 157.950 406.950 160.050 407.400 ;
        RECT 190.950 408.600 193.050 409.050 ;
        RECT 202.950 408.600 205.050 409.050 ;
        RECT 190.950 407.400 205.050 408.600 ;
        RECT 239.400 408.600 240.600 413.400 ;
        RECT 292.950 412.950 295.050 413.400 ;
        RECT 241.950 411.600 244.050 412.050 ;
        RECT 253.950 411.600 256.050 412.050 ;
        RECT 241.950 410.400 256.050 411.600 ;
        RECT 241.950 409.950 244.050 410.400 ;
        RECT 253.950 409.950 256.050 410.400 ;
        RECT 271.950 411.600 274.050 412.050 ;
        RECT 295.950 411.600 298.050 412.050 ;
        RECT 271.950 410.400 298.050 411.600 ;
        RECT 299.400 411.600 300.600 413.400 ;
        RECT 301.950 412.950 304.050 415.050 ;
        RECT 322.950 412.950 325.050 415.050 ;
        RECT 304.950 411.600 307.050 412.050 ;
        RECT 299.400 410.400 307.050 411.600 ;
        RECT 323.400 411.600 324.600 412.950 ;
        RECT 331.950 411.600 334.050 412.050 ;
        RECT 323.400 410.400 334.050 411.600 ;
        RECT 271.950 409.950 274.050 410.400 ;
        RECT 295.950 409.950 298.050 410.400 ;
        RECT 304.950 409.950 307.050 410.400 ;
        RECT 331.950 409.950 334.050 410.400 ;
        RECT 244.950 408.600 247.050 409.050 ;
        RECT 239.400 407.400 247.050 408.600 ;
        RECT 190.950 406.950 193.050 407.400 ;
        RECT 202.950 406.950 205.050 407.400 ;
        RECT 244.950 406.950 247.050 407.400 ;
        RECT 250.950 408.600 253.050 409.050 ;
        RECT 265.950 408.600 268.050 409.050 ;
        RECT 250.950 407.400 268.050 408.600 ;
        RECT 250.950 406.950 253.050 407.400 ;
        RECT 265.950 406.950 268.050 407.400 ;
        RECT 277.950 408.600 280.050 409.050 ;
        RECT 310.950 408.600 313.050 409.050 ;
        RECT 277.950 407.400 313.050 408.600 ;
        RECT 277.950 406.950 280.050 407.400 ;
        RECT 310.950 406.950 313.050 407.400 ;
        RECT 319.950 408.600 322.050 409.050 ;
        RECT 328.950 408.600 331.050 409.050 ;
        RECT 319.950 407.400 331.050 408.600 ;
        RECT 319.950 406.950 322.050 407.400 ;
        RECT 328.950 406.950 331.050 407.400 ;
        RECT 337.950 408.600 340.050 409.050 ;
        RECT 341.400 408.600 342.600 415.950 ;
        RECT 364.950 414.600 367.050 415.050 ;
        RECT 350.400 413.400 367.050 414.600 ;
        RECT 350.400 412.050 351.600 413.400 ;
        RECT 364.950 412.950 367.050 413.400 ;
        RECT 367.950 412.950 370.050 415.050 ;
        RECT 421.950 414.600 424.050 415.050 ;
        RECT 416.400 413.400 424.050 414.600 ;
        RECT 349.950 409.950 352.050 412.050 ;
        RECT 368.400 411.600 369.600 412.950 ;
        RECT 416.400 412.050 417.600 413.400 ;
        RECT 421.950 412.950 424.050 413.400 ;
        RECT 376.950 411.600 379.050 412.050 ;
        RECT 368.400 410.400 379.050 411.600 ;
        RECT 376.950 409.950 379.050 410.400 ;
        RECT 382.950 411.600 385.050 412.050 ;
        RECT 388.950 411.600 391.050 412.050 ;
        RECT 382.950 410.400 391.050 411.600 ;
        RECT 382.950 409.950 385.050 410.400 ;
        RECT 388.950 409.950 391.050 410.400 ;
        RECT 415.950 409.950 418.050 412.050 ;
        RECT 337.950 407.400 342.600 408.600 ;
        RECT 346.950 408.600 349.050 409.050 ;
        RECT 418.950 408.600 421.050 409.050 ;
        RECT 424.950 408.600 427.050 409.050 ;
        RECT 427.950 408.600 430.050 409.050 ;
        RECT 346.950 407.400 366.600 408.600 ;
        RECT 337.950 406.950 340.050 407.400 ;
        RECT 346.950 406.950 349.050 407.400 ;
        RECT 16.950 405.600 19.050 406.050 ;
        RECT 88.950 405.600 91.050 406.050 ;
        RECT 106.950 405.600 109.050 406.050 ;
        RECT 16.950 404.400 109.050 405.600 ;
        RECT 16.950 403.950 19.050 404.400 ;
        RECT 88.950 403.950 91.050 404.400 ;
        RECT 106.950 403.950 109.050 404.400 ;
        RECT 121.950 405.600 124.050 406.050 ;
        RECT 178.950 405.600 181.050 406.050 ;
        RECT 121.950 404.400 181.050 405.600 ;
        RECT 121.950 403.950 124.050 404.400 ;
        RECT 178.950 403.950 181.050 404.400 ;
        RECT 265.950 405.600 268.050 406.050 ;
        RECT 277.950 405.600 280.050 406.050 ;
        RECT 265.950 404.400 280.050 405.600 ;
        RECT 265.950 403.950 268.050 404.400 ;
        RECT 277.950 403.950 280.050 404.400 ;
        RECT 295.950 405.600 298.050 406.050 ;
        RECT 316.950 405.600 319.050 406.050 ;
        RECT 295.950 404.400 319.050 405.600 ;
        RECT 295.950 403.950 298.050 404.400 ;
        RECT 316.950 403.950 319.050 404.400 ;
        RECT 343.950 405.600 346.050 406.050 ;
        RECT 352.950 405.600 355.050 406.050 ;
        RECT 343.950 404.400 355.050 405.600 ;
        RECT 365.400 405.600 366.600 407.400 ;
        RECT 418.950 407.400 430.050 408.600 ;
        RECT 418.950 406.950 421.050 407.400 ;
        RECT 424.950 406.950 427.050 407.400 ;
        RECT 427.950 406.950 430.050 407.400 ;
        RECT 433.950 408.600 436.050 409.050 ;
        RECT 443.400 408.600 444.600 415.950 ;
        RECT 464.400 411.600 465.600 415.950 ;
        RECT 479.400 415.050 480.600 416.400 ;
        RECT 505.950 415.950 508.050 416.400 ;
        RECT 511.950 415.950 514.050 416.400 ;
        RECT 517.950 417.600 520.050 418.050 ;
        RECT 532.950 417.600 535.050 418.050 ;
        RECT 517.950 416.400 535.050 417.600 ;
        RECT 517.950 415.950 520.050 416.400 ;
        RECT 532.950 415.950 535.050 416.400 ;
        RECT 553.950 417.600 556.050 418.050 ;
        RECT 562.950 417.600 565.050 418.050 ;
        RECT 553.950 416.400 565.050 417.600 ;
        RECT 553.950 415.950 556.050 416.400 ;
        RECT 562.950 415.950 565.050 416.400 ;
        RECT 568.950 417.600 571.050 418.050 ;
        RECT 580.950 417.600 583.050 418.050 ;
        RECT 640.950 417.600 643.050 418.050 ;
        RECT 568.950 416.400 583.050 417.600 ;
        RECT 568.950 415.950 571.050 416.400 ;
        RECT 580.950 415.950 583.050 416.400 ;
        RECT 632.400 416.400 643.050 417.600 ;
        RECT 478.950 412.950 481.050 415.050 ;
        RECT 484.950 414.600 487.050 415.050 ;
        RECT 508.950 414.600 511.050 415.050 ;
        RECT 523.950 414.600 526.050 415.050 ;
        RECT 484.950 413.400 504.600 414.600 ;
        RECT 484.950 412.950 487.050 413.400 ;
        RECT 503.400 412.050 504.600 413.400 ;
        RECT 508.950 413.400 526.050 414.600 ;
        RECT 508.950 412.950 511.050 413.400 ;
        RECT 523.950 412.950 526.050 413.400 ;
        RECT 529.950 414.600 532.050 415.050 ;
        RECT 538.950 414.600 541.050 415.050 ;
        RECT 547.950 414.600 550.050 415.050 ;
        RECT 529.950 413.400 550.050 414.600 ;
        RECT 529.950 412.950 532.050 413.400 ;
        RECT 538.950 412.950 541.050 413.400 ;
        RECT 547.950 412.950 550.050 413.400 ;
        RECT 565.950 414.600 568.050 415.050 ;
        RECT 586.950 414.600 589.050 415.050 ;
        RECT 598.950 414.600 601.050 415.050 ;
        RECT 607.950 414.600 610.050 415.050 ;
        RECT 565.950 413.400 597.600 414.600 ;
        RECT 565.950 412.950 568.050 413.400 ;
        RECT 586.950 412.950 589.050 413.400 ;
        RECT 596.400 412.050 597.600 413.400 ;
        RECT 598.950 413.400 610.050 414.600 ;
        RECT 598.950 412.950 601.050 413.400 ;
        RECT 607.950 412.950 610.050 413.400 ;
        RECT 616.950 414.600 619.050 415.050 ;
        RECT 625.950 414.600 628.050 415.050 ;
        RECT 632.400 414.600 633.600 416.400 ;
        RECT 640.950 415.950 643.050 416.400 ;
        RECT 643.950 417.600 646.050 418.050 ;
        RECT 652.950 417.600 655.050 418.050 ;
        RECT 643.950 416.400 655.050 417.600 ;
        RECT 643.950 415.950 646.050 416.400 ;
        RECT 652.950 415.950 655.050 416.400 ;
        RECT 656.400 416.400 663.600 417.600 ;
        RECT 616.950 413.400 628.050 414.600 ;
        RECT 616.950 412.950 619.050 413.400 ;
        RECT 625.950 412.950 628.050 413.400 ;
        RECT 629.400 413.400 633.600 414.600 ;
        RECT 637.950 414.600 640.050 415.050 ;
        RECT 646.950 414.600 649.050 415.050 ;
        RECT 656.400 414.600 657.600 416.400 ;
        RECT 637.950 413.400 645.600 414.600 ;
        RECT 481.950 411.600 484.050 412.050 ;
        RECT 464.400 410.400 484.050 411.600 ;
        RECT 481.950 409.950 484.050 410.400 ;
        RECT 502.950 411.600 505.050 412.050 ;
        RECT 502.950 410.400 507.600 411.600 ;
        RECT 502.950 409.950 505.050 410.400 ;
        RECT 506.400 409.050 507.600 410.400 ;
        RECT 511.950 409.950 514.050 412.050 ;
        RECT 526.950 411.600 529.050 412.050 ;
        RECT 592.950 411.600 595.050 412.050 ;
        RECT 526.950 410.400 595.050 411.600 ;
        RECT 526.950 409.950 529.050 410.400 ;
        RECT 592.950 409.950 595.050 410.400 ;
        RECT 595.950 409.950 598.050 412.050 ;
        RECT 601.950 411.600 604.050 412.050 ;
        RECT 629.400 411.600 630.600 413.400 ;
        RECT 637.950 412.950 640.050 413.400 ;
        RECT 601.950 410.400 630.600 411.600 ;
        RECT 644.400 411.600 645.600 413.400 ;
        RECT 646.950 413.400 657.600 414.600 ;
        RECT 646.950 412.950 649.050 413.400 ;
        RECT 658.950 412.950 661.050 415.050 ;
        RECT 649.950 411.600 652.050 412.050 ;
        RECT 655.950 411.600 658.050 412.050 ;
        RECT 644.400 410.400 652.050 411.600 ;
        RECT 601.950 409.950 604.050 410.400 ;
        RECT 649.950 409.950 652.050 410.400 ;
        RECT 653.400 410.400 658.050 411.600 ;
        RECT 433.950 407.400 444.600 408.600 ;
        RECT 448.950 408.600 451.050 409.050 ;
        RECT 448.950 407.400 498.600 408.600 ;
        RECT 433.950 406.950 436.050 407.400 ;
        RECT 448.950 406.950 451.050 407.400 ;
        RECT 373.950 405.600 376.050 406.050 ;
        RECT 365.400 404.400 376.050 405.600 ;
        RECT 343.950 403.950 346.050 404.400 ;
        RECT 352.950 403.950 355.050 404.400 ;
        RECT 373.950 403.950 376.050 404.400 ;
        RECT 397.950 405.600 400.050 406.050 ;
        RECT 493.950 405.600 496.050 406.050 ;
        RECT 397.950 404.400 496.050 405.600 ;
        RECT 497.400 405.600 498.600 407.400 ;
        RECT 505.950 406.950 508.050 409.050 ;
        RECT 512.400 408.600 513.600 409.950 ;
        RECT 550.950 408.600 553.050 409.050 ;
        RECT 556.950 408.600 559.050 409.050 ;
        RECT 512.400 407.400 549.600 408.600 ;
        RECT 514.950 405.600 517.050 406.050 ;
        RECT 544.950 405.600 547.050 406.050 ;
        RECT 497.400 404.400 547.050 405.600 ;
        RECT 548.400 405.600 549.600 407.400 ;
        RECT 550.950 407.400 559.050 408.600 ;
        RECT 550.950 406.950 553.050 407.400 ;
        RECT 556.950 406.950 559.050 407.400 ;
        RECT 565.950 408.600 568.050 409.050 ;
        RECT 613.950 408.600 616.050 409.050 ;
        RECT 565.950 407.400 616.050 408.600 ;
        RECT 565.950 406.950 568.050 407.400 ;
        RECT 613.950 406.950 616.050 407.400 ;
        RECT 622.950 408.600 625.050 409.050 ;
        RECT 653.400 408.600 654.600 410.400 ;
        RECT 655.950 409.950 658.050 410.400 ;
        RECT 622.950 407.400 654.600 408.600 ;
        RECT 655.950 408.600 658.050 409.050 ;
        RECT 659.400 408.600 660.600 412.950 ;
        RECT 662.400 412.050 663.600 416.400 ;
        RECT 661.950 409.950 664.050 412.050 ;
        RECT 670.950 411.600 673.050 412.050 ;
        RECT 674.400 411.600 675.600 418.950 ;
        RECT 676.950 415.950 679.050 418.050 ;
        RECT 685.950 417.600 688.050 418.050 ;
        RECT 697.950 417.600 700.050 418.050 ;
        RECT 685.950 416.400 700.050 417.600 ;
        RECT 701.400 417.600 702.600 419.400 ;
        RECT 724.950 419.400 732.600 420.600 ;
        RECT 724.950 418.950 727.050 419.400 ;
        RECT 715.950 417.600 718.050 418.050 ;
        RECT 727.950 417.600 730.050 418.050 ;
        RECT 701.400 416.400 705.600 417.600 ;
        RECT 685.950 415.950 688.050 416.400 ;
        RECT 697.950 415.950 700.050 416.400 ;
        RECT 677.400 412.050 678.600 415.950 ;
        RECT 688.950 414.600 691.050 415.050 ;
        RECT 680.400 413.400 691.050 414.600 ;
        RECT 670.950 410.400 675.600 411.600 ;
        RECT 670.950 409.950 673.050 410.400 ;
        RECT 676.950 409.950 679.050 412.050 ;
        RECT 655.950 407.400 660.600 408.600 ;
        RECT 680.400 408.600 681.600 413.400 ;
        RECT 688.950 412.950 691.050 413.400 ;
        RECT 691.950 414.600 694.050 415.050 ;
        RECT 700.950 414.600 703.050 415.050 ;
        RECT 691.950 413.400 703.050 414.600 ;
        RECT 691.950 412.950 694.050 413.400 ;
        RECT 700.950 412.950 703.050 413.400 ;
        RECT 682.950 411.600 685.050 412.050 ;
        RECT 704.400 411.600 705.600 416.400 ;
        RECT 715.950 416.400 730.050 417.600 ;
        RECT 715.950 415.950 718.050 416.400 ;
        RECT 727.950 415.950 730.050 416.400 ;
        RECT 718.950 414.600 721.050 415.050 ;
        RECT 682.950 410.400 705.600 411.600 ;
        RECT 707.400 413.400 721.050 414.600 ;
        RECT 682.950 409.950 685.050 410.400 ;
        RECT 697.950 408.600 700.050 409.050 ;
        RECT 680.400 407.400 700.050 408.600 ;
        RECT 622.950 406.950 625.050 407.400 ;
        RECT 655.950 406.950 658.050 407.400 ;
        RECT 697.950 406.950 700.050 407.400 ;
        RECT 703.950 408.600 706.050 409.050 ;
        RECT 707.400 408.600 708.600 413.400 ;
        RECT 718.950 412.950 721.050 413.400 ;
        RECT 721.950 414.600 724.050 415.050 ;
        RECT 727.950 414.600 730.050 415.050 ;
        RECT 731.400 414.600 732.600 419.400 ;
        RECT 739.950 418.950 742.050 421.050 ;
        RECT 745.950 420.600 748.050 421.050 ;
        RECT 766.950 420.600 769.050 421.050 ;
        RECT 745.950 419.400 769.050 420.600 ;
        RECT 745.950 418.950 748.050 419.400 ;
        RECT 766.950 418.950 769.050 419.400 ;
        RECT 721.950 413.400 726.600 414.600 ;
        RECT 721.950 412.950 724.050 413.400 ;
        RECT 725.400 411.600 726.600 413.400 ;
        RECT 727.950 413.400 732.600 414.600 ;
        RECT 727.950 412.950 730.050 413.400 ;
        RECT 730.950 411.600 733.050 412.050 ;
        RECT 725.400 410.400 733.050 411.600 ;
        RECT 740.400 411.600 741.600 418.950 ;
        RECT 745.950 414.600 748.050 415.050 ;
        RECT 760.950 414.600 763.050 415.050 ;
        RECT 745.950 413.400 763.050 414.600 ;
        RECT 745.950 412.950 748.050 413.400 ;
        RECT 760.950 412.950 763.050 413.400 ;
        RECT 748.950 411.600 751.050 412.050 ;
        RECT 740.400 410.400 751.050 411.600 ;
        RECT 730.950 409.950 733.050 410.400 ;
        RECT 748.950 409.950 751.050 410.400 ;
        RECT 703.950 407.400 708.600 408.600 ;
        RECT 730.950 408.600 733.050 409.050 ;
        RECT 766.950 408.600 769.050 409.050 ;
        RECT 730.950 407.400 769.050 408.600 ;
        RECT 703.950 406.950 706.050 407.400 ;
        RECT 730.950 406.950 733.050 407.400 ;
        RECT 766.950 406.950 769.050 407.400 ;
        RECT 577.950 405.600 580.050 406.050 ;
        RECT 548.400 404.400 580.050 405.600 ;
        RECT 397.950 403.950 400.050 404.400 ;
        RECT 493.950 403.950 496.050 404.400 ;
        RECT 514.950 403.950 517.050 404.400 ;
        RECT 544.950 403.950 547.050 404.400 ;
        RECT 577.950 403.950 580.050 404.400 ;
        RECT 583.950 405.600 586.050 406.050 ;
        RECT 619.950 405.600 622.050 406.050 ;
        RECT 583.950 404.400 622.050 405.600 ;
        RECT 583.950 403.950 586.050 404.400 ;
        RECT 619.950 403.950 622.050 404.400 ;
        RECT 628.950 405.600 631.050 406.050 ;
        RECT 637.950 405.600 640.050 406.050 ;
        RECT 667.950 405.600 670.050 406.050 ;
        RECT 628.950 404.400 670.050 405.600 ;
        RECT 628.950 403.950 631.050 404.400 ;
        RECT 637.950 403.950 640.050 404.400 ;
        RECT 667.950 403.950 670.050 404.400 ;
        RECT 688.950 405.600 691.050 406.050 ;
        RECT 700.950 405.600 703.050 406.050 ;
        RECT 688.950 404.400 703.050 405.600 ;
        RECT 688.950 403.950 691.050 404.400 ;
        RECT 700.950 403.950 703.050 404.400 ;
        RECT 706.950 405.600 709.050 406.050 ;
        RECT 724.950 405.600 727.050 406.050 ;
        RECT 706.950 404.400 727.050 405.600 ;
        RECT 706.950 403.950 709.050 404.400 ;
        RECT 724.950 403.950 727.050 404.400 ;
        RECT 217.950 402.600 220.050 403.050 ;
        RECT 298.950 402.600 301.050 403.050 ;
        RECT 217.950 401.400 301.050 402.600 ;
        RECT 217.950 400.950 220.050 401.400 ;
        RECT 298.950 400.950 301.050 401.400 ;
        RECT 307.950 402.600 310.050 403.050 ;
        RECT 337.950 402.600 340.050 403.050 ;
        RECT 307.950 401.400 340.050 402.600 ;
        RECT 307.950 400.950 310.050 401.400 ;
        RECT 337.950 400.950 340.050 401.400 ;
        RECT 379.950 402.600 382.050 403.050 ;
        RECT 385.950 402.600 388.050 403.050 ;
        RECT 379.950 401.400 388.050 402.600 ;
        RECT 379.950 400.950 382.050 401.400 ;
        RECT 385.950 400.950 388.050 401.400 ;
        RECT 427.950 402.600 430.050 403.050 ;
        RECT 439.950 402.600 442.050 403.050 ;
        RECT 427.950 401.400 442.050 402.600 ;
        RECT 427.950 400.950 430.050 401.400 ;
        RECT 439.950 400.950 442.050 401.400 ;
        RECT 448.950 402.600 451.050 403.050 ;
        RECT 466.950 402.600 469.050 403.050 ;
        RECT 448.950 401.400 469.050 402.600 ;
        RECT 448.950 400.950 451.050 401.400 ;
        RECT 466.950 400.950 469.050 401.400 ;
        RECT 487.950 402.600 490.050 403.050 ;
        RECT 511.950 402.600 514.050 403.050 ;
        RECT 487.950 401.400 514.050 402.600 ;
        RECT 487.950 400.950 490.050 401.400 ;
        RECT 511.950 400.950 514.050 401.400 ;
        RECT 514.950 402.600 517.050 403.050 ;
        RECT 535.950 402.600 538.050 403.050 ;
        RECT 541.950 402.600 544.050 403.050 ;
        RECT 514.950 401.400 544.050 402.600 ;
        RECT 514.950 400.950 517.050 401.400 ;
        RECT 535.950 400.950 538.050 401.400 ;
        RECT 541.950 400.950 544.050 401.400 ;
        RECT 571.950 402.600 574.050 403.050 ;
        RECT 583.950 402.600 586.050 403.050 ;
        RECT 631.950 402.600 634.050 403.050 ;
        RECT 571.950 401.400 586.050 402.600 ;
        RECT 571.950 400.950 574.050 401.400 ;
        RECT 583.950 400.950 586.050 401.400 ;
        RECT 602.400 401.400 634.050 402.600 ;
        RECT 130.950 399.600 133.050 400.050 ;
        RECT 235.950 399.600 238.050 400.050 ;
        RECT 274.950 399.600 277.050 400.050 ;
        RECT 334.950 399.600 337.050 400.050 ;
        RECT 130.950 398.400 337.050 399.600 ;
        RECT 130.950 397.950 133.050 398.400 ;
        RECT 235.950 397.950 238.050 398.400 ;
        RECT 274.950 397.950 277.050 398.400 ;
        RECT 334.950 397.950 337.050 398.400 ;
        RECT 337.950 399.600 340.050 400.050 ;
        RECT 364.950 399.600 367.050 400.050 ;
        RECT 394.950 399.600 397.050 400.050 ;
        RECT 337.950 398.400 397.050 399.600 ;
        RECT 337.950 397.950 340.050 398.400 ;
        RECT 364.950 397.950 367.050 398.400 ;
        RECT 394.950 397.950 397.050 398.400 ;
        RECT 430.950 399.600 433.050 400.050 ;
        RECT 460.950 399.600 463.050 400.050 ;
        RECT 430.950 398.400 463.050 399.600 ;
        RECT 430.950 397.950 433.050 398.400 ;
        RECT 460.950 397.950 463.050 398.400 ;
        RECT 520.950 399.600 523.050 400.050 ;
        RECT 602.400 399.600 603.600 401.400 ;
        RECT 631.950 400.950 634.050 401.400 ;
        RECT 658.950 402.600 661.050 403.050 ;
        RECT 676.950 402.600 679.050 403.050 ;
        RECT 658.950 401.400 679.050 402.600 ;
        RECT 658.950 400.950 661.050 401.400 ;
        RECT 676.950 400.950 679.050 401.400 ;
        RECT 733.950 402.600 736.050 403.050 ;
        RECT 742.950 402.600 745.050 403.050 ;
        RECT 733.950 401.400 745.050 402.600 ;
        RECT 733.950 400.950 736.050 401.400 ;
        RECT 742.950 400.950 745.050 401.400 ;
        RECT 520.950 398.400 603.600 399.600 ;
        RECT 616.950 399.600 619.050 400.050 ;
        RECT 661.950 399.600 664.050 400.050 ;
        RECT 667.950 399.600 670.050 400.050 ;
        RECT 673.950 399.600 676.050 400.050 ;
        RECT 739.950 399.600 742.050 400.050 ;
        RECT 616.950 398.400 627.600 399.600 ;
        RECT 520.950 397.950 523.050 398.400 ;
        RECT 616.950 397.950 619.050 398.400 ;
        RECT 355.950 396.600 358.050 397.050 ;
        RECT 439.950 396.600 442.050 397.050 ;
        RECT 355.950 395.400 442.050 396.600 ;
        RECT 355.950 394.950 358.050 395.400 ;
        RECT 439.950 394.950 442.050 395.400 ;
        RECT 442.950 396.600 445.050 397.050 ;
        RECT 466.950 396.600 469.050 397.050 ;
        RECT 511.950 396.600 514.050 397.050 ;
        RECT 571.950 396.600 574.050 397.050 ;
        RECT 598.950 396.600 601.050 397.050 ;
        RECT 622.950 396.600 625.050 397.050 ;
        RECT 442.950 395.400 465.600 396.600 ;
        RECT 442.950 394.950 445.050 395.400 ;
        RECT 136.950 393.600 139.050 394.050 ;
        RECT 271.950 393.600 274.050 394.050 ;
        RECT 136.950 392.400 274.050 393.600 ;
        RECT 136.950 391.950 139.050 392.400 ;
        RECT 271.950 391.950 274.050 392.400 ;
        RECT 277.950 393.600 280.050 394.050 ;
        RECT 310.950 393.600 313.050 394.050 ;
        RECT 277.950 392.400 313.050 393.600 ;
        RECT 277.950 391.950 280.050 392.400 ;
        RECT 310.950 391.950 313.050 392.400 ;
        RECT 361.950 393.600 364.050 394.050 ;
        RECT 400.950 393.600 403.050 394.050 ;
        RECT 361.950 392.400 403.050 393.600 ;
        RECT 464.400 393.600 465.600 395.400 ;
        RECT 466.950 395.400 601.050 396.600 ;
        RECT 466.950 394.950 469.050 395.400 ;
        RECT 511.950 394.950 514.050 395.400 ;
        RECT 571.950 394.950 574.050 395.400 ;
        RECT 598.950 394.950 601.050 395.400 ;
        RECT 602.400 395.400 625.050 396.600 ;
        RECT 626.400 396.600 627.600 398.400 ;
        RECT 661.950 398.400 742.050 399.600 ;
        RECT 661.950 397.950 664.050 398.400 ;
        RECT 667.950 397.950 670.050 398.400 ;
        RECT 673.950 397.950 676.050 398.400 ;
        RECT 739.950 397.950 742.050 398.400 ;
        RECT 751.950 399.600 754.050 400.050 ;
        RECT 751.950 398.400 774.600 399.600 ;
        RECT 751.950 397.950 754.050 398.400 ;
        RECT 676.950 396.600 679.050 397.050 ;
        RECT 626.400 395.400 679.050 396.600 ;
        RECT 502.950 393.600 505.050 394.050 ;
        RECT 464.400 392.400 505.050 393.600 ;
        RECT 361.950 391.950 364.050 392.400 ;
        RECT 400.950 391.950 403.050 392.400 ;
        RECT 502.950 391.950 505.050 392.400 ;
        RECT 505.950 393.600 508.050 394.050 ;
        RECT 526.950 393.600 529.050 394.050 ;
        RECT 562.950 393.600 565.050 394.050 ;
        RECT 505.950 392.400 565.050 393.600 ;
        RECT 505.950 391.950 508.050 392.400 ;
        RECT 526.950 391.950 529.050 392.400 ;
        RECT 562.950 391.950 565.050 392.400 ;
        RECT 580.950 393.600 583.050 394.050 ;
        RECT 586.950 393.600 589.050 394.050 ;
        RECT 602.400 393.600 603.600 395.400 ;
        RECT 622.950 394.950 625.050 395.400 ;
        RECT 676.950 394.950 679.050 395.400 ;
        RECT 685.950 396.600 688.050 397.050 ;
        RECT 697.950 396.600 700.050 397.050 ;
        RECT 685.950 395.400 700.050 396.600 ;
        RECT 685.950 394.950 688.050 395.400 ;
        RECT 697.950 394.950 700.050 395.400 ;
        RECT 715.950 396.600 718.050 397.050 ;
        RECT 769.950 396.600 772.050 397.050 ;
        RECT 715.950 395.400 772.050 396.600 ;
        RECT 715.950 394.950 718.050 395.400 ;
        RECT 769.950 394.950 772.050 395.400 ;
        RECT 580.950 392.400 603.600 393.600 ;
        RECT 613.950 393.600 616.050 394.050 ;
        RECT 637.950 393.600 640.050 394.050 ;
        RECT 670.950 393.600 673.050 394.050 ;
        RECT 613.950 392.400 640.050 393.600 ;
        RECT 580.950 391.950 583.050 392.400 ;
        RECT 586.950 391.950 589.050 392.400 ;
        RECT 613.950 391.950 616.050 392.400 ;
        RECT 637.950 391.950 640.050 392.400 ;
        RECT 668.400 392.400 673.050 393.600 ;
        RECT 1.950 390.600 4.050 391.050 ;
        RECT 25.950 390.600 28.050 391.050 ;
        RECT 1.950 389.400 28.050 390.600 ;
        RECT 1.950 388.950 4.050 389.400 ;
        RECT 25.950 388.950 28.050 389.400 ;
        RECT 43.950 390.600 46.050 391.050 ;
        RECT 94.950 390.600 97.050 391.050 ;
        RECT 43.950 389.400 97.050 390.600 ;
        RECT 43.950 388.950 46.050 389.400 ;
        RECT 94.950 388.950 97.050 389.400 ;
        RECT 145.950 390.600 148.050 391.050 ;
        RECT 151.950 390.600 154.050 391.050 ;
        RECT 145.950 389.400 154.050 390.600 ;
        RECT 145.950 388.950 148.050 389.400 ;
        RECT 151.950 388.950 154.050 389.400 ;
        RECT 154.950 390.600 157.050 391.050 ;
        RECT 184.950 390.600 187.050 391.050 ;
        RECT 154.950 389.400 187.050 390.600 ;
        RECT 154.950 388.950 157.050 389.400 ;
        RECT 184.950 388.950 187.050 389.400 ;
        RECT 316.950 390.600 319.050 391.050 ;
        RECT 352.950 390.600 355.050 391.050 ;
        RECT 394.950 390.600 397.050 391.050 ;
        RECT 430.950 390.600 433.050 391.050 ;
        RECT 436.950 390.600 439.050 391.050 ;
        RECT 316.950 389.400 439.050 390.600 ;
        RECT 316.950 388.950 319.050 389.400 ;
        RECT 352.950 388.950 355.050 389.400 ;
        RECT 394.950 388.950 397.050 389.400 ;
        RECT 430.950 388.950 433.050 389.400 ;
        RECT 436.950 388.950 439.050 389.400 ;
        RECT 475.950 390.600 478.050 391.050 ;
        RECT 487.950 390.600 490.050 391.050 ;
        RECT 475.950 389.400 490.050 390.600 ;
        RECT 475.950 388.950 478.050 389.400 ;
        RECT 487.950 388.950 490.050 389.400 ;
        RECT 490.950 390.600 493.050 391.050 ;
        RECT 505.950 390.600 508.050 391.050 ;
        RECT 490.950 389.400 508.050 390.600 ;
        RECT 490.950 388.950 493.050 389.400 ;
        RECT 505.950 388.950 508.050 389.400 ;
        RECT 559.950 390.600 562.050 391.050 ;
        RECT 568.950 390.600 571.050 391.050 ;
        RECT 559.950 389.400 571.050 390.600 ;
        RECT 559.950 388.950 562.050 389.400 ;
        RECT 568.950 388.950 571.050 389.400 ;
        RECT 574.950 390.600 577.050 391.050 ;
        RECT 583.950 390.600 586.050 391.050 ;
        RECT 574.950 389.400 586.050 390.600 ;
        RECT 574.950 388.950 577.050 389.400 ;
        RECT 583.950 388.950 586.050 389.400 ;
        RECT 589.950 390.600 592.050 391.050 ;
        RECT 604.950 390.600 607.050 391.050 ;
        RECT 668.400 390.600 669.600 392.400 ;
        RECT 670.950 391.950 673.050 392.400 ;
        RECT 676.950 393.600 679.050 394.050 ;
        RECT 715.950 393.600 718.050 394.050 ;
        RECT 676.950 392.400 718.050 393.600 ;
        RECT 676.950 391.950 679.050 392.400 ;
        RECT 715.950 391.950 718.050 392.400 ;
        RECT 727.950 393.600 730.050 394.050 ;
        RECT 745.950 393.600 748.050 394.050 ;
        RECT 727.950 392.400 748.050 393.600 ;
        RECT 727.950 391.950 730.050 392.400 ;
        RECT 745.950 391.950 748.050 392.400 ;
        RECT 757.950 393.600 760.050 394.050 ;
        RECT 769.950 393.600 772.050 394.050 ;
        RECT 757.950 392.400 772.050 393.600 ;
        RECT 757.950 391.950 760.050 392.400 ;
        RECT 769.950 391.950 772.050 392.400 ;
        RECT 589.950 389.400 607.050 390.600 ;
        RECT 589.950 388.950 592.050 389.400 ;
        RECT 604.950 388.950 607.050 389.400 ;
        RECT 662.400 389.400 669.600 390.600 ;
        RECT 670.950 390.600 673.050 391.050 ;
        RECT 694.950 390.600 697.050 391.050 ;
        RECT 670.950 389.400 697.050 390.600 ;
        RECT 34.950 387.600 37.050 388.050 ;
        RECT 43.950 387.600 46.050 388.050 ;
        RECT 34.950 386.400 46.050 387.600 ;
        RECT 34.950 385.950 37.050 386.400 ;
        RECT 43.950 385.950 46.050 386.400 ;
        RECT 67.950 387.600 70.050 388.050 ;
        RECT 73.950 387.600 76.050 388.050 ;
        RECT 67.950 386.400 76.050 387.600 ;
        RECT 67.950 385.950 70.050 386.400 ;
        RECT 73.950 385.950 76.050 386.400 ;
        RECT 82.950 385.950 85.050 388.050 ;
        RECT 88.950 387.600 91.050 388.050 ;
        RECT 97.950 387.600 100.050 388.050 ;
        RECT 217.950 387.600 220.050 388.050 ;
        RECT 88.950 386.400 100.050 387.600 ;
        RECT 88.950 385.950 91.050 386.400 ;
        RECT 97.950 385.950 100.050 386.400 ;
        RECT 179.400 386.400 220.050 387.600 ;
        RECT 10.950 384.600 13.050 385.050 ;
        RECT 28.950 384.600 31.050 385.050 ;
        RECT 10.950 383.400 31.050 384.600 ;
        RECT 10.950 382.950 13.050 383.400 ;
        RECT 28.950 382.950 31.050 383.400 ;
        RECT 58.950 384.600 61.050 385.050 ;
        RECT 76.950 384.600 79.050 385.050 ;
        RECT 58.950 383.400 79.050 384.600 ;
        RECT 58.950 382.950 61.050 383.400 ;
        RECT 76.950 382.950 79.050 383.400 ;
        RECT 46.950 381.600 49.050 382.050 ;
        RECT 55.950 381.600 58.050 382.050 ;
        RECT 46.950 380.400 58.050 381.600 ;
        RECT 46.950 379.950 49.050 380.400 ;
        RECT 55.950 379.950 58.050 380.400 ;
        RECT 70.950 381.600 73.050 382.050 ;
        RECT 83.400 381.600 84.600 385.950 ;
        RECT 179.400 385.050 180.600 386.400 ;
        RECT 217.950 385.950 220.050 386.400 ;
        RECT 238.950 387.600 241.050 388.050 ;
        RECT 247.950 387.600 250.050 388.050 ;
        RECT 283.950 387.600 286.050 388.050 ;
        RECT 238.950 386.400 250.050 387.600 ;
        RECT 238.950 385.950 241.050 386.400 ;
        RECT 247.950 385.950 250.050 386.400 ;
        RECT 275.400 386.400 286.050 387.600 ;
        RECT 91.950 384.600 94.050 385.050 ;
        RECT 100.950 384.600 103.050 385.050 ;
        RECT 91.950 383.400 103.050 384.600 ;
        RECT 91.950 382.950 94.050 383.400 ;
        RECT 100.950 382.950 103.050 383.400 ;
        RECT 115.950 384.600 118.050 385.050 ;
        RECT 121.950 384.600 124.050 385.050 ;
        RECT 115.950 383.400 124.050 384.600 ;
        RECT 115.950 382.950 118.050 383.400 ;
        RECT 121.950 382.950 124.050 383.400 ;
        RECT 178.950 382.950 181.050 385.050 ;
        RECT 187.950 384.600 190.050 385.050 ;
        RECT 187.950 383.400 195.600 384.600 ;
        RECT 187.950 382.950 190.050 383.400 ;
        RECT 194.400 382.050 195.600 383.400 ;
        RECT 205.950 382.950 208.050 385.050 ;
        RECT 232.950 384.600 235.050 385.050 ;
        RECT 241.950 384.600 244.050 385.050 ;
        RECT 259.950 384.600 262.050 385.050 ;
        RECT 232.950 383.400 244.050 384.600 ;
        RECT 232.950 382.950 235.050 383.400 ;
        RECT 241.950 382.950 244.050 383.400 ;
        RECT 251.400 383.400 262.050 384.600 ;
        RECT 70.950 380.400 84.600 381.600 ;
        RECT 85.950 381.600 88.050 382.050 ;
        RECT 94.950 381.600 97.050 382.050 ;
        RECT 85.950 380.400 97.050 381.600 ;
        RECT 70.950 379.950 73.050 380.400 ;
        RECT 85.950 379.950 88.050 380.400 ;
        RECT 94.950 379.950 97.050 380.400 ;
        RECT 97.950 381.600 100.050 382.050 ;
        RECT 106.950 381.600 109.050 382.050 ;
        RECT 109.950 381.600 112.050 382.050 ;
        RECT 127.950 381.600 130.050 382.050 ;
        RECT 97.950 380.400 102.600 381.600 ;
        RECT 97.950 379.950 100.050 380.400 ;
        RECT 4.950 378.600 7.050 379.050 ;
        RECT 37.950 378.600 40.050 379.050 ;
        RECT 4.950 377.400 40.050 378.600 ;
        RECT 4.950 376.950 7.050 377.400 ;
        RECT 37.950 376.950 40.050 377.400 ;
        RECT 70.950 378.600 73.050 379.050 ;
        RECT 97.950 378.600 100.050 379.050 ;
        RECT 70.950 377.400 100.050 378.600 ;
        RECT 70.950 376.950 73.050 377.400 ;
        RECT 97.950 376.950 100.050 377.400 ;
        RECT 79.950 375.600 82.050 376.050 ;
        RECT 88.950 375.600 91.050 376.050 ;
        RECT 91.950 375.600 94.050 376.050 ;
        RECT 79.950 374.400 94.050 375.600 ;
        RECT 79.950 373.950 82.050 374.400 ;
        RECT 88.950 373.950 91.050 374.400 ;
        RECT 91.950 373.950 94.050 374.400 ;
        RECT 94.950 375.600 97.050 376.050 ;
        RECT 101.400 375.600 102.600 380.400 ;
        RECT 106.950 380.400 130.050 381.600 ;
        RECT 106.950 379.950 109.050 380.400 ;
        RECT 109.950 379.950 112.050 380.400 ;
        RECT 127.950 379.950 130.050 380.400 ;
        RECT 157.950 379.950 160.050 382.050 ;
        RECT 181.950 381.600 184.050 382.050 ;
        RECT 190.950 381.600 193.050 382.050 ;
        RECT 181.950 380.400 193.050 381.600 ;
        RECT 181.950 379.950 184.050 380.400 ;
        RECT 190.950 379.950 193.050 380.400 ;
        RECT 193.950 379.950 196.050 382.050 ;
        RECT 196.950 381.600 199.050 382.050 ;
        RECT 206.400 381.600 207.600 382.950 ;
        RECT 251.400 382.050 252.600 383.400 ;
        RECT 259.950 382.950 262.050 383.400 ;
        RECT 275.400 382.050 276.600 386.400 ;
        RECT 283.950 385.950 286.050 386.400 ;
        RECT 286.950 387.600 289.050 388.050 ;
        RECT 337.950 387.600 340.050 388.050 ;
        RECT 286.950 386.400 340.050 387.600 ;
        RECT 286.950 385.950 289.050 386.400 ;
        RECT 337.950 385.950 340.050 386.400 ;
        RECT 343.950 387.600 346.050 388.050 ;
        RECT 349.950 387.600 352.050 388.050 ;
        RECT 343.950 386.400 352.050 387.600 ;
        RECT 343.950 385.950 346.050 386.400 ;
        RECT 349.950 385.950 352.050 386.400 ;
        RECT 358.950 385.950 361.050 388.050 ;
        RECT 376.950 387.600 379.050 388.050 ;
        RECT 409.950 387.600 412.050 388.050 ;
        RECT 436.950 387.600 439.050 388.050 ;
        RECT 376.950 386.400 384.600 387.600 ;
        RECT 376.950 385.950 379.050 386.400 ;
        RECT 283.950 382.950 286.050 385.050 ;
        RECT 289.950 384.600 292.050 385.050 ;
        RECT 301.950 384.600 304.050 385.050 ;
        RECT 328.950 384.600 331.050 385.050 ;
        RECT 289.950 383.400 331.050 384.600 ;
        RECT 289.950 382.950 292.050 383.400 ;
        RECT 301.950 382.950 304.050 383.400 ;
        RECT 328.950 382.950 331.050 383.400 ;
        RECT 349.950 384.600 352.050 385.050 ;
        RECT 355.950 384.600 358.050 385.050 ;
        RECT 349.950 383.400 358.050 384.600 ;
        RECT 349.950 382.950 352.050 383.400 ;
        RECT 355.950 382.950 358.050 383.400 ;
        RECT 196.950 380.400 207.600 381.600 ;
        RECT 196.950 379.950 199.050 380.400 ;
        RECT 250.950 379.950 253.050 382.050 ;
        RECT 274.950 379.950 277.050 382.050 ;
        RECT 284.400 381.600 285.600 382.950 ;
        RECT 359.400 382.050 360.600 385.950 ;
        RECT 383.400 385.050 384.600 386.400 ;
        RECT 409.950 386.400 439.050 387.600 ;
        RECT 409.950 385.950 412.050 386.400 ;
        RECT 436.950 385.950 439.050 386.400 ;
        RECT 475.950 387.600 478.050 388.050 ;
        RECT 484.950 387.600 487.050 388.050 ;
        RECT 475.950 386.400 487.050 387.600 ;
        RECT 475.950 385.950 478.050 386.400 ;
        RECT 484.950 385.950 487.050 386.400 ;
        RECT 493.950 387.600 496.050 388.050 ;
        RECT 499.950 387.600 502.050 388.050 ;
        RECT 493.950 386.400 502.050 387.600 ;
        RECT 493.950 385.950 496.050 386.400 ;
        RECT 499.950 385.950 502.050 386.400 ;
        RECT 502.950 387.600 505.050 388.050 ;
        RECT 508.950 387.600 511.050 388.050 ;
        RECT 532.950 387.600 535.050 388.050 ;
        RECT 547.950 387.600 550.050 388.050 ;
        RECT 592.950 387.600 595.050 388.050 ;
        RECT 502.950 386.400 507.600 387.600 ;
        RECT 502.950 385.950 505.050 386.400 ;
        RECT 367.950 382.950 370.050 385.050 ;
        RECT 382.950 384.600 385.050 385.050 ;
        RECT 388.950 384.600 391.050 385.050 ;
        RECT 382.950 383.400 391.050 384.600 ;
        RECT 382.950 382.950 385.050 383.400 ;
        RECT 388.950 382.950 391.050 383.400 ;
        RECT 418.950 384.600 421.050 385.050 ;
        RECT 424.950 384.600 427.050 385.050 ;
        RECT 457.950 384.600 460.050 385.050 ;
        RECT 418.950 383.400 427.050 384.600 ;
        RECT 418.950 382.950 421.050 383.400 ;
        RECT 424.950 382.950 427.050 383.400 ;
        RECT 428.400 383.400 460.050 384.600 ;
        RECT 292.950 381.600 295.050 382.050 ;
        RECT 284.400 380.400 295.050 381.600 ;
        RECT 292.950 379.950 295.050 380.400 ;
        RECT 358.950 379.950 361.050 382.050 ;
        RECT 368.400 381.600 369.600 382.950 ;
        RECT 373.950 381.600 376.050 382.050 ;
        RECT 428.400 381.600 429.600 383.400 ;
        RECT 457.950 382.950 460.050 383.400 ;
        RECT 463.950 384.600 466.050 385.050 ;
        RECT 469.950 384.600 472.050 385.050 ;
        RECT 463.950 383.400 472.050 384.600 ;
        RECT 463.950 382.950 466.050 383.400 ;
        RECT 469.950 382.950 472.050 383.400 ;
        RECT 368.400 380.400 376.050 381.600 ;
        RECT 373.950 379.950 376.050 380.400 ;
        RECT 377.400 380.400 429.600 381.600 ;
        RECT 472.950 381.600 475.050 382.050 ;
        RECT 487.950 381.600 490.050 382.050 ;
        RECT 472.950 380.400 490.050 381.600 ;
        RECT 506.400 381.600 507.600 386.400 ;
        RECT 508.950 386.400 522.600 387.600 ;
        RECT 508.950 385.950 511.050 386.400 ;
        RECT 508.950 384.600 511.050 385.050 ;
        RECT 517.950 384.600 520.050 385.050 ;
        RECT 508.950 383.400 520.050 384.600 ;
        RECT 521.400 384.600 522.600 386.400 ;
        RECT 532.950 386.400 550.050 387.600 ;
        RECT 532.950 385.950 535.050 386.400 ;
        RECT 547.950 385.950 550.050 386.400 ;
        RECT 551.400 386.400 595.050 387.600 ;
        RECT 541.950 384.600 544.050 385.050 ;
        RECT 551.400 384.600 552.600 386.400 ;
        RECT 592.950 385.950 595.050 386.400 ;
        RECT 616.950 387.600 619.050 388.050 ;
        RECT 631.950 387.600 634.050 388.050 ;
        RECT 616.950 386.400 634.050 387.600 ;
        RECT 616.950 385.950 619.050 386.400 ;
        RECT 631.950 385.950 634.050 386.400 ;
        RECT 640.950 387.600 643.050 388.050 ;
        RECT 646.950 387.600 649.050 388.050 ;
        RECT 652.950 387.600 655.050 388.050 ;
        RECT 640.950 386.400 655.050 387.600 ;
        RECT 640.950 385.950 643.050 386.400 ;
        RECT 646.950 385.950 649.050 386.400 ;
        RECT 652.950 385.950 655.050 386.400 ;
        RECT 658.950 385.950 661.050 388.050 ;
        RECT 521.400 383.400 537.600 384.600 ;
        RECT 508.950 382.950 511.050 383.400 ;
        RECT 517.950 382.950 520.050 383.400 ;
        RECT 532.950 381.600 535.050 382.050 ;
        RECT 506.400 380.400 535.050 381.600 ;
        RECT 103.950 378.600 106.050 379.050 ;
        RECT 112.950 378.600 115.050 379.050 ;
        RECT 103.950 377.400 115.050 378.600 ;
        RECT 103.950 376.950 106.050 377.400 ;
        RECT 112.950 376.950 115.050 377.400 ;
        RECT 118.950 378.600 121.050 379.050 ;
        RECT 136.950 378.600 139.050 379.050 ;
        RECT 118.950 377.400 139.050 378.600 ;
        RECT 118.950 376.950 121.050 377.400 ;
        RECT 136.950 376.950 139.050 377.400 ;
        RECT 139.950 378.600 142.050 379.050 ;
        RECT 154.950 378.600 157.050 379.050 ;
        RECT 139.950 377.400 157.050 378.600 ;
        RECT 139.950 376.950 142.050 377.400 ;
        RECT 154.950 376.950 157.050 377.400 ;
        RECT 94.950 374.400 102.600 375.600 ;
        RECT 158.400 375.600 159.600 379.950 ;
        RECT 160.950 378.600 163.050 379.050 ;
        RECT 238.950 378.600 241.050 379.050 ;
        RECT 286.950 378.600 289.050 379.050 ;
        RECT 160.950 377.400 237.600 378.600 ;
        RECT 160.950 376.950 163.050 377.400 ;
        RECT 160.950 375.600 163.050 376.050 ;
        RECT 158.400 374.400 163.050 375.600 ;
        RECT 236.400 375.600 237.600 377.400 ;
        RECT 238.950 377.400 289.050 378.600 ;
        RECT 238.950 376.950 241.050 377.400 ;
        RECT 286.950 376.950 289.050 377.400 ;
        RECT 331.950 378.600 334.050 379.050 ;
        RECT 337.950 378.600 340.050 379.050 ;
        RECT 331.950 377.400 340.050 378.600 ;
        RECT 331.950 376.950 334.050 377.400 ;
        RECT 337.950 376.950 340.050 377.400 ;
        RECT 346.950 378.600 349.050 379.050 ;
        RECT 377.400 378.600 378.600 380.400 ;
        RECT 472.950 379.950 475.050 380.400 ;
        RECT 487.950 379.950 490.050 380.400 ;
        RECT 532.950 379.950 535.050 380.400 ;
        RECT 346.950 377.400 378.600 378.600 ;
        RECT 400.950 378.600 403.050 379.050 ;
        RECT 451.950 378.600 454.050 379.050 ;
        RECT 400.950 377.400 454.050 378.600 ;
        RECT 346.950 376.950 349.050 377.400 ;
        RECT 400.950 376.950 403.050 377.400 ;
        RECT 451.950 376.950 454.050 377.400 ;
        RECT 484.950 376.950 487.050 379.050 ;
        RECT 499.950 378.600 502.050 379.050 ;
        RECT 514.950 378.600 517.050 379.050 ;
        RECT 499.950 377.400 517.050 378.600 ;
        RECT 499.950 376.950 502.050 377.400 ;
        RECT 514.950 376.950 517.050 377.400 ;
        RECT 517.950 378.600 520.050 379.050 ;
        RECT 529.950 378.600 532.050 379.050 ;
        RECT 536.400 378.600 537.600 383.400 ;
        RECT 541.950 383.400 552.600 384.600 ;
        RECT 559.950 384.600 562.050 385.050 ;
        RECT 574.950 384.600 577.050 385.050 ;
        RECT 559.950 383.400 577.050 384.600 ;
        RECT 541.950 382.950 544.050 383.400 ;
        RECT 559.950 382.950 562.050 383.400 ;
        RECT 574.950 382.950 577.050 383.400 ;
        RECT 598.950 384.600 601.050 385.050 ;
        RECT 622.950 384.600 625.050 385.050 ;
        RECT 598.950 383.400 625.050 384.600 ;
        RECT 598.950 382.950 601.050 383.400 ;
        RECT 622.950 382.950 625.050 383.400 ;
        RECT 649.950 382.950 652.050 385.050 ;
        RECT 547.950 381.600 550.050 382.050 ;
        RECT 553.950 381.600 556.050 382.050 ;
        RECT 547.950 380.400 556.050 381.600 ;
        RECT 547.950 379.950 550.050 380.400 ;
        RECT 553.950 379.950 556.050 380.400 ;
        RECT 577.950 381.600 580.050 382.050 ;
        RECT 589.950 381.600 592.050 382.050 ;
        RECT 577.950 380.400 592.050 381.600 ;
        RECT 577.950 379.950 580.050 380.400 ;
        RECT 589.950 379.950 592.050 380.400 ;
        RECT 595.950 381.600 598.050 382.050 ;
        RECT 604.950 381.600 607.050 382.050 ;
        RECT 625.950 381.600 628.050 382.050 ;
        RECT 595.950 380.400 628.050 381.600 ;
        RECT 595.950 379.950 598.050 380.400 ;
        RECT 604.950 379.950 607.050 380.400 ;
        RECT 625.950 379.950 628.050 380.400 ;
        RECT 631.950 379.950 634.050 382.050 ;
        RECT 517.950 377.400 537.600 378.600 ;
        RECT 544.950 378.600 547.050 379.050 ;
        RECT 613.950 378.600 616.050 379.050 ;
        RECT 544.950 377.400 616.050 378.600 ;
        RECT 517.950 376.950 520.050 377.400 ;
        RECT 529.950 376.950 532.050 377.400 ;
        RECT 544.950 376.950 547.050 377.400 ;
        RECT 613.950 376.950 616.050 377.400 ;
        RECT 619.950 378.600 622.050 379.050 ;
        RECT 628.950 378.600 631.050 379.050 ;
        RECT 619.950 377.400 631.050 378.600 ;
        RECT 619.950 376.950 622.050 377.400 ;
        RECT 628.950 376.950 631.050 377.400 ;
        RECT 349.950 375.600 352.050 376.050 ;
        RECT 236.400 374.400 352.050 375.600 ;
        RECT 94.950 373.950 97.050 374.400 ;
        RECT 160.950 373.950 163.050 374.400 ;
        RECT 349.950 373.950 352.050 374.400 ;
        RECT 364.950 375.600 367.050 376.050 ;
        RECT 379.950 375.600 382.050 376.050 ;
        RECT 364.950 374.400 382.050 375.600 ;
        RECT 364.950 373.950 367.050 374.400 ;
        RECT 379.950 373.950 382.050 374.400 ;
        RECT 76.950 372.600 79.050 373.050 ;
        RECT 121.950 372.600 124.050 373.050 ;
        RECT 76.950 371.400 124.050 372.600 ;
        RECT 76.950 370.950 79.050 371.400 ;
        RECT 121.950 370.950 124.050 371.400 ;
        RECT 235.950 372.600 238.050 373.050 ;
        RECT 256.950 372.600 259.050 373.050 ;
        RECT 235.950 371.400 259.050 372.600 ;
        RECT 235.950 370.950 238.050 371.400 ;
        RECT 256.950 370.950 259.050 371.400 ;
        RECT 280.950 372.600 283.050 373.050 ;
        RECT 331.950 372.600 334.050 373.050 ;
        RECT 340.950 372.600 343.050 373.050 ;
        RECT 364.950 372.600 367.050 373.050 ;
        RECT 280.950 371.400 367.050 372.600 ;
        RECT 280.950 370.950 283.050 371.400 ;
        RECT 331.950 370.950 334.050 371.400 ;
        RECT 340.950 370.950 343.050 371.400 ;
        RECT 364.950 370.950 367.050 371.400 ;
        RECT 367.950 372.600 370.050 373.050 ;
        RECT 391.950 372.600 394.050 373.050 ;
        RECT 367.950 371.400 394.050 372.600 ;
        RECT 367.950 370.950 370.050 371.400 ;
        RECT 391.950 370.950 394.050 371.400 ;
        RECT 433.950 372.600 436.050 373.050 ;
        RECT 463.950 372.600 466.050 373.050 ;
        RECT 481.950 372.600 484.050 373.050 ;
        RECT 433.950 371.400 484.050 372.600 ;
        RECT 485.400 372.600 486.600 376.950 ;
        RECT 490.950 375.600 493.050 376.050 ;
        RECT 505.950 375.600 508.050 376.050 ;
        RECT 490.950 374.400 508.050 375.600 ;
        RECT 490.950 373.950 493.050 374.400 ;
        RECT 505.950 373.950 508.050 374.400 ;
        RECT 550.950 375.600 553.050 376.050 ;
        RECT 613.950 375.600 616.050 376.050 ;
        RECT 550.950 374.400 616.050 375.600 ;
        RECT 550.950 373.950 553.050 374.400 ;
        RECT 613.950 373.950 616.050 374.400 ;
        RECT 538.950 372.600 541.050 373.050 ;
        RECT 485.400 371.400 541.050 372.600 ;
        RECT 433.950 370.950 436.050 371.400 ;
        RECT 463.950 370.950 466.050 371.400 ;
        RECT 481.950 370.950 484.050 371.400 ;
        RECT 538.950 370.950 541.050 371.400 ;
        RECT 568.950 372.600 571.050 373.050 ;
        RECT 604.950 372.600 607.050 373.050 ;
        RECT 568.950 371.400 607.050 372.600 ;
        RECT 629.400 372.600 630.600 376.950 ;
        RECT 632.400 375.600 633.600 379.950 ;
        RECT 646.950 375.600 649.050 376.050 ;
        RECT 632.400 374.400 649.050 375.600 ;
        RECT 650.400 375.600 651.600 382.950 ;
        RECT 659.400 381.600 660.600 385.950 ;
        RECT 662.400 384.600 663.600 389.400 ;
        RECT 670.950 388.950 673.050 389.400 ;
        RECT 694.950 388.950 697.050 389.400 ;
        RECT 709.950 390.600 712.050 391.050 ;
        RECT 733.950 390.600 736.050 391.050 ;
        RECT 709.950 389.400 736.050 390.600 ;
        RECT 709.950 388.950 712.050 389.400 ;
        RECT 733.950 388.950 736.050 389.400 ;
        RECT 736.950 390.600 739.050 391.050 ;
        RECT 736.950 389.400 756.600 390.600 ;
        RECT 736.950 388.950 739.050 389.400 ;
        RECT 664.950 387.600 667.050 388.050 ;
        RECT 682.950 387.600 685.050 388.050 ;
        RECT 664.950 386.400 685.050 387.600 ;
        RECT 664.950 385.950 667.050 386.400 ;
        RECT 682.950 385.950 685.050 386.400 ;
        RECT 688.950 385.950 691.050 388.050 ;
        RECT 691.950 387.600 694.050 388.050 ;
        RECT 709.950 387.600 712.050 388.050 ;
        RECT 691.950 386.400 712.050 387.600 ;
        RECT 691.950 385.950 694.050 386.400 ;
        RECT 709.950 385.950 712.050 386.400 ;
        RECT 715.950 387.600 718.050 388.050 ;
        RECT 736.950 387.600 739.050 388.050 ;
        RECT 751.950 387.600 754.050 388.050 ;
        RECT 715.950 386.400 739.050 387.600 ;
        RECT 715.950 385.950 718.050 386.400 ;
        RECT 736.950 385.950 739.050 386.400 ;
        RECT 740.400 386.400 754.050 387.600 ;
        RECT 664.950 384.600 667.050 385.050 ;
        RECT 662.400 383.400 667.050 384.600 ;
        RECT 664.950 382.950 667.050 383.400 ;
        RECT 661.950 381.600 664.050 382.050 ;
        RECT 659.400 380.400 664.050 381.600 ;
        RECT 689.400 381.600 690.600 385.950 ;
        RECT 703.950 384.600 706.050 385.050 ;
        RECT 740.400 384.600 741.600 386.400 ;
        RECT 751.950 385.950 754.050 386.400 ;
        RECT 745.950 384.600 748.050 385.050 ;
        RECT 755.400 384.600 756.600 389.400 ;
        RECT 703.950 383.400 741.600 384.600 ;
        RECT 743.400 383.400 748.050 384.600 ;
        RECT 703.950 382.950 706.050 383.400 ;
        RECT 689.400 380.400 699.600 381.600 ;
        RECT 661.950 379.950 664.050 380.400 ;
        RECT 658.950 378.600 661.050 379.050 ;
        RECT 694.950 378.600 697.050 379.050 ;
        RECT 658.950 377.400 697.050 378.600 ;
        RECT 698.400 378.600 699.600 380.400 ;
        RECT 709.950 379.950 712.050 382.050 ;
        RECT 724.950 381.600 727.050 382.050 ;
        RECT 736.950 381.600 739.050 382.050 ;
        RECT 743.400 381.600 744.600 383.400 ;
        RECT 745.950 382.950 748.050 383.400 ;
        RECT 749.400 383.400 756.600 384.600 ;
        RECT 749.400 381.600 750.600 383.400 ;
        RECT 724.950 380.400 739.050 381.600 ;
        RECT 724.950 379.950 727.050 380.400 ;
        RECT 736.950 379.950 739.050 380.400 ;
        RECT 740.400 380.400 744.600 381.600 ;
        RECT 746.400 380.400 750.600 381.600 ;
        RECT 751.950 381.600 754.050 382.050 ;
        RECT 760.950 381.600 763.050 382.050 ;
        RECT 751.950 380.400 763.050 381.600 ;
        RECT 700.950 378.600 703.050 379.050 ;
        RECT 698.400 377.400 703.050 378.600 ;
        RECT 658.950 376.950 661.050 377.400 ;
        RECT 694.950 376.950 697.050 377.400 ;
        RECT 700.950 376.950 703.050 377.400 ;
        RECT 706.950 376.950 709.050 379.050 ;
        RECT 710.400 378.600 711.600 379.950 ;
        RECT 740.400 379.050 741.600 380.400 ;
        RECT 733.950 378.600 736.050 379.050 ;
        RECT 710.400 377.400 736.050 378.600 ;
        RECT 733.950 376.950 736.050 377.400 ;
        RECT 739.950 376.950 742.050 379.050 ;
        RECT 742.950 378.600 745.050 379.050 ;
        RECT 746.400 378.600 747.600 380.400 ;
        RECT 751.950 379.950 754.050 380.400 ;
        RECT 760.950 379.950 763.050 380.400 ;
        RECT 742.950 377.400 747.600 378.600 ;
        RECT 760.950 378.600 763.050 379.050 ;
        RECT 773.400 378.600 774.600 398.400 ;
        RECT 760.950 377.400 774.600 378.600 ;
        RECT 742.950 376.950 745.050 377.400 ;
        RECT 760.950 376.950 763.050 377.400 ;
        RECT 652.950 375.600 655.050 376.050 ;
        RECT 650.400 374.400 655.050 375.600 ;
        RECT 646.950 373.950 649.050 374.400 ;
        RECT 652.950 373.950 655.050 374.400 ;
        RECT 679.950 375.600 682.050 376.050 ;
        RECT 685.950 375.600 688.050 376.050 ;
        RECT 679.950 374.400 688.050 375.600 ;
        RECT 679.950 373.950 682.050 374.400 ;
        RECT 685.950 373.950 688.050 374.400 ;
        RECT 694.950 375.600 697.050 376.050 ;
        RECT 707.400 375.600 708.600 376.950 ;
        RECT 733.950 375.600 736.050 376.050 ;
        RECT 776.400 375.600 777.600 422.400 ;
        RECT 694.950 374.400 732.600 375.600 ;
        RECT 694.950 373.950 697.050 374.400 ;
        RECT 643.950 372.600 646.050 373.050 ;
        RECT 629.400 371.400 646.050 372.600 ;
        RECT 731.400 372.600 732.600 374.400 ;
        RECT 733.950 374.400 777.600 375.600 ;
        RECT 733.950 373.950 736.050 374.400 ;
        RECT 736.950 372.600 739.050 373.050 ;
        RECT 731.400 371.400 739.050 372.600 ;
        RECT 568.950 370.950 571.050 371.400 ;
        RECT 604.950 370.950 607.050 371.400 ;
        RECT 643.950 370.950 646.050 371.400 ;
        RECT 736.950 370.950 739.050 371.400 ;
        RECT 262.950 369.600 265.050 370.050 ;
        RECT 553.950 369.600 556.050 370.050 ;
        RECT 262.950 368.400 556.050 369.600 ;
        RECT 262.950 367.950 265.050 368.400 ;
        RECT 553.950 367.950 556.050 368.400 ;
        RECT 577.950 369.600 580.050 370.050 ;
        RECT 631.950 369.600 634.050 370.050 ;
        RECT 577.950 368.400 634.050 369.600 ;
        RECT 577.950 367.950 580.050 368.400 ;
        RECT 631.950 367.950 634.050 368.400 ;
        RECT 640.950 369.600 643.050 370.050 ;
        RECT 667.950 369.600 670.050 370.050 ;
        RECT 640.950 368.400 670.050 369.600 ;
        RECT 640.950 367.950 643.050 368.400 ;
        RECT 667.950 367.950 670.050 368.400 ;
        RECT 691.950 369.600 694.050 370.050 ;
        RECT 700.950 369.600 703.050 370.050 ;
        RECT 691.950 368.400 703.050 369.600 ;
        RECT 691.950 367.950 694.050 368.400 ;
        RECT 700.950 367.950 703.050 368.400 ;
        RECT 718.950 369.600 721.050 370.050 ;
        RECT 763.950 369.600 766.050 370.050 ;
        RECT 718.950 368.400 766.050 369.600 ;
        RECT 718.950 367.950 721.050 368.400 ;
        RECT 763.950 367.950 766.050 368.400 ;
        RECT 238.950 366.600 241.050 367.050 ;
        RECT 244.950 366.600 247.050 367.050 ;
        RECT 280.950 366.600 283.050 367.050 ;
        RECT 238.950 365.400 283.050 366.600 ;
        RECT 238.950 364.950 241.050 365.400 ;
        RECT 244.950 364.950 247.050 365.400 ;
        RECT 280.950 364.950 283.050 365.400 ;
        RECT 286.950 366.600 289.050 367.050 ;
        RECT 313.950 366.600 316.050 367.050 ;
        RECT 286.950 365.400 316.050 366.600 ;
        RECT 286.950 364.950 289.050 365.400 ;
        RECT 313.950 364.950 316.050 365.400 ;
        RECT 322.950 366.600 325.050 367.050 ;
        RECT 346.950 366.600 349.050 367.050 ;
        RECT 322.950 365.400 349.050 366.600 ;
        RECT 322.950 364.950 325.050 365.400 ;
        RECT 346.950 364.950 349.050 365.400 ;
        RECT 406.950 366.600 409.050 367.050 ;
        RECT 448.950 366.600 451.050 367.050 ;
        RECT 406.950 365.400 451.050 366.600 ;
        RECT 406.950 364.950 409.050 365.400 ;
        RECT 448.950 364.950 451.050 365.400 ;
        RECT 493.950 366.600 496.050 367.050 ;
        RECT 514.950 366.600 517.050 367.050 ;
        RECT 493.950 365.400 517.050 366.600 ;
        RECT 493.950 364.950 496.050 365.400 ;
        RECT 514.950 364.950 517.050 365.400 ;
        RECT 523.950 366.600 526.050 367.050 ;
        RECT 601.950 366.600 604.050 367.050 ;
        RECT 523.950 365.400 604.050 366.600 ;
        RECT 523.950 364.950 526.050 365.400 ;
        RECT 601.950 364.950 604.050 365.400 ;
        RECT 604.950 366.600 607.050 367.050 ;
        RECT 652.950 366.600 655.050 367.050 ;
        RECT 604.950 365.400 655.050 366.600 ;
        RECT 604.950 364.950 607.050 365.400 ;
        RECT 652.950 364.950 655.050 365.400 ;
        RECT 673.950 366.600 676.050 367.050 ;
        RECT 688.950 366.600 691.050 367.050 ;
        RECT 718.950 366.600 721.050 367.050 ;
        RECT 673.950 365.400 721.050 366.600 ;
        RECT 673.950 364.950 676.050 365.400 ;
        RECT 688.950 364.950 691.050 365.400 ;
        RECT 718.950 364.950 721.050 365.400 ;
        RECT 757.950 366.600 760.050 367.050 ;
        RECT 763.950 366.600 766.050 367.050 ;
        RECT 757.950 365.400 766.050 366.600 ;
        RECT 757.950 364.950 760.050 365.400 ;
        RECT 763.950 364.950 766.050 365.400 ;
        RECT 67.950 363.600 70.050 364.050 ;
        RECT 73.950 363.600 76.050 364.050 ;
        RECT 67.950 362.400 76.050 363.600 ;
        RECT 67.950 361.950 70.050 362.400 ;
        RECT 73.950 361.950 76.050 362.400 ;
        RECT 439.950 363.600 442.050 364.050 ;
        RECT 535.950 363.600 538.050 364.050 ;
        RECT 439.950 362.400 538.050 363.600 ;
        RECT 439.950 361.950 442.050 362.400 ;
        RECT 535.950 361.950 538.050 362.400 ;
        RECT 589.950 363.600 592.050 364.050 ;
        RECT 640.950 363.600 643.050 364.050 ;
        RECT 589.950 362.400 643.050 363.600 ;
        RECT 589.950 361.950 592.050 362.400 ;
        RECT 640.950 361.950 643.050 362.400 ;
        RECT 712.950 363.600 715.050 364.050 ;
        RECT 748.950 363.600 751.050 364.050 ;
        RECT 712.950 362.400 751.050 363.600 ;
        RECT 712.950 361.950 715.050 362.400 ;
        RECT 748.950 361.950 751.050 362.400 ;
        RECT 451.950 360.600 454.050 361.050 ;
        RECT 496.950 360.600 499.050 361.050 ;
        RECT 451.950 359.400 499.050 360.600 ;
        RECT 451.950 358.950 454.050 359.400 ;
        RECT 496.950 358.950 499.050 359.400 ;
        RECT 517.950 360.600 520.050 361.050 ;
        RECT 526.950 360.600 529.050 361.050 ;
        RECT 604.950 360.600 607.050 361.050 ;
        RECT 517.950 359.400 607.050 360.600 ;
        RECT 517.950 358.950 520.050 359.400 ;
        RECT 526.950 358.950 529.050 359.400 ;
        RECT 604.950 358.950 607.050 359.400 ;
        RECT 607.950 360.600 610.050 361.050 ;
        RECT 619.950 360.600 622.050 361.050 ;
        RECT 607.950 359.400 622.050 360.600 ;
        RECT 607.950 358.950 610.050 359.400 ;
        RECT 619.950 358.950 622.050 359.400 ;
        RECT 631.950 360.600 634.050 361.050 ;
        RECT 718.950 360.600 721.050 361.050 ;
        RECT 754.950 360.600 757.050 361.050 ;
        RECT 631.950 359.400 757.050 360.600 ;
        RECT 631.950 358.950 634.050 359.400 ;
        RECT 718.950 358.950 721.050 359.400 ;
        RECT 754.950 358.950 757.050 359.400 ;
        RECT 217.950 357.600 220.050 358.050 ;
        RECT 226.950 357.600 229.050 358.050 ;
        RECT 217.950 356.400 229.050 357.600 ;
        RECT 217.950 355.950 220.050 356.400 ;
        RECT 226.950 355.950 229.050 356.400 ;
        RECT 352.950 357.600 355.050 358.050 ;
        RECT 361.950 357.600 364.050 358.050 ;
        RECT 352.950 356.400 364.050 357.600 ;
        RECT 352.950 355.950 355.050 356.400 ;
        RECT 361.950 355.950 364.050 356.400 ;
        RECT 460.950 357.600 463.050 358.050 ;
        RECT 484.950 357.600 487.050 358.050 ;
        RECT 502.950 357.600 505.050 358.050 ;
        RECT 538.950 357.600 541.050 358.050 ;
        RECT 460.950 356.400 541.050 357.600 ;
        RECT 460.950 355.950 463.050 356.400 ;
        RECT 484.950 355.950 487.050 356.400 ;
        RECT 502.950 355.950 505.050 356.400 ;
        RECT 538.950 355.950 541.050 356.400 ;
        RECT 571.950 357.600 574.050 358.050 ;
        RECT 595.950 357.600 598.050 358.050 ;
        RECT 571.950 356.400 598.050 357.600 ;
        RECT 571.950 355.950 574.050 356.400 ;
        RECT 595.950 355.950 598.050 356.400 ;
        RECT 610.950 357.600 613.050 358.050 ;
        RECT 658.950 357.600 661.050 358.050 ;
        RECT 610.950 356.400 661.050 357.600 ;
        RECT 610.950 355.950 613.050 356.400 ;
        RECT 658.950 355.950 661.050 356.400 ;
        RECT 85.950 354.600 88.050 355.050 ;
        RECT 292.950 354.600 295.050 355.050 ;
        RECT 85.950 353.400 295.050 354.600 ;
        RECT 85.950 352.950 88.050 353.400 ;
        RECT 292.950 352.950 295.050 353.400 ;
        RECT 478.950 354.600 481.050 355.050 ;
        RECT 556.950 354.600 559.050 355.050 ;
        RECT 478.950 353.400 559.050 354.600 ;
        RECT 478.950 352.950 481.050 353.400 ;
        RECT 556.950 352.950 559.050 353.400 ;
        RECT 562.950 354.600 565.050 355.050 ;
        RECT 571.950 354.600 574.050 355.050 ;
        RECT 562.950 353.400 574.050 354.600 ;
        RECT 562.950 352.950 565.050 353.400 ;
        RECT 571.950 352.950 574.050 353.400 ;
        RECT 592.950 354.600 595.050 355.050 ;
        RECT 661.950 354.600 664.050 355.050 ;
        RECT 592.950 353.400 664.050 354.600 ;
        RECT 592.950 352.950 595.050 353.400 ;
        RECT 661.950 352.950 664.050 353.400 ;
        RECT 52.950 351.600 55.050 352.050 ;
        RECT 106.950 351.600 109.050 352.050 ;
        RECT 52.950 350.400 109.050 351.600 ;
        RECT 52.950 349.950 55.050 350.400 ;
        RECT 106.950 349.950 109.050 350.400 ;
        RECT 325.950 351.600 328.050 352.050 ;
        RECT 334.950 351.600 337.050 352.050 ;
        RECT 325.950 350.400 337.050 351.600 ;
        RECT 325.950 349.950 328.050 350.400 ;
        RECT 334.950 349.950 337.050 350.400 ;
        RECT 403.950 351.600 406.050 352.050 ;
        RECT 439.950 351.600 442.050 352.050 ;
        RECT 403.950 350.400 442.050 351.600 ;
        RECT 403.950 349.950 406.050 350.400 ;
        RECT 439.950 349.950 442.050 350.400 ;
        RECT 445.950 351.600 448.050 352.050 ;
        RECT 487.950 351.600 490.050 352.050 ;
        RECT 550.950 351.600 553.050 352.050 ;
        RECT 445.950 350.400 490.050 351.600 ;
        RECT 445.950 349.950 448.050 350.400 ;
        RECT 487.950 349.950 490.050 350.400 ;
        RECT 503.400 350.400 553.050 351.600 ;
        RECT 112.950 348.600 115.050 349.050 ;
        RECT 68.400 347.400 115.050 348.600 ;
        RECT 68.400 343.050 69.600 347.400 ;
        RECT 112.950 346.950 115.050 347.400 ;
        RECT 274.950 348.600 277.050 349.050 ;
        RECT 361.950 348.600 364.050 349.050 ;
        RECT 274.950 347.400 364.050 348.600 ;
        RECT 274.950 346.950 277.050 347.400 ;
        RECT 361.950 346.950 364.050 347.400 ;
        RECT 382.950 348.600 385.050 349.050 ;
        RECT 412.950 348.600 415.050 349.050 ;
        RECT 382.950 347.400 415.050 348.600 ;
        RECT 382.950 346.950 385.050 347.400 ;
        RECT 412.950 346.950 415.050 347.400 ;
        RECT 415.950 348.600 418.050 349.050 ;
        RECT 466.950 348.600 469.050 349.050 ;
        RECT 475.950 348.600 478.050 349.050 ;
        RECT 499.950 348.600 502.050 349.050 ;
        RECT 415.950 347.400 465.600 348.600 ;
        RECT 415.950 346.950 418.050 347.400 ;
        RECT 70.950 345.600 73.050 346.050 ;
        RECT 355.950 345.600 358.050 346.050 ;
        RECT 70.950 344.400 84.600 345.600 ;
        RECT 70.950 343.950 73.050 344.400 ;
        RECT 83.400 343.050 84.600 344.400 ;
        RECT 332.400 344.400 358.050 345.600 ;
        RECT 7.950 342.600 10.050 343.050 ;
        RECT 16.950 342.600 19.050 343.050 ;
        RECT 7.950 341.400 19.050 342.600 ;
        RECT 7.950 340.950 10.050 341.400 ;
        RECT 16.950 340.950 19.050 341.400 ;
        RECT 31.950 342.600 34.050 343.050 ;
        RECT 31.950 341.400 48.600 342.600 ;
        RECT 31.950 340.950 34.050 341.400 ;
        RECT 47.400 340.050 48.600 341.400 ;
        RECT 67.950 340.950 70.050 343.050 ;
        RECT 79.950 342.600 82.050 343.050 ;
        RECT 74.400 341.400 82.050 342.600 ;
        RECT 13.950 339.600 16.050 340.050 ;
        RECT 25.950 339.600 28.050 340.050 ;
        RECT 34.950 339.600 37.050 340.050 ;
        RECT 13.950 338.400 37.050 339.600 ;
        RECT 13.950 337.950 16.050 338.400 ;
        RECT 25.950 337.950 28.050 338.400 ;
        RECT 34.950 337.950 37.050 338.400 ;
        RECT 46.950 337.950 49.050 340.050 ;
        RECT 55.950 339.600 58.050 340.050 ;
        RECT 74.400 339.600 75.600 341.400 ;
        RECT 79.950 340.950 82.050 341.400 ;
        RECT 82.950 340.950 85.050 343.050 ;
        RECT 100.950 342.600 103.050 343.050 ;
        RECT 106.950 342.600 109.050 343.050 ;
        RECT 100.950 341.400 109.050 342.600 ;
        RECT 100.950 340.950 103.050 341.400 ;
        RECT 106.950 340.950 109.050 341.400 ;
        RECT 121.950 342.600 124.050 343.050 ;
        RECT 127.950 342.600 130.050 343.050 ;
        RECT 139.950 342.600 142.050 343.050 ;
        RECT 121.950 341.400 142.050 342.600 ;
        RECT 121.950 340.950 124.050 341.400 ;
        RECT 127.950 340.950 130.050 341.400 ;
        RECT 139.950 340.950 142.050 341.400 ;
        RECT 151.950 340.950 154.050 343.050 ;
        RECT 169.950 342.600 172.050 343.050 ;
        RECT 193.950 342.600 196.050 343.050 ;
        RECT 205.950 342.600 208.050 343.050 ;
        RECT 169.950 341.400 192.600 342.600 ;
        RECT 169.950 340.950 172.050 341.400 ;
        RECT 55.950 338.400 75.600 339.600 ;
        RECT 76.950 339.600 79.050 340.050 ;
        RECT 88.950 339.600 91.050 340.050 ;
        RECT 100.950 339.600 103.050 340.050 ;
        RECT 76.950 338.400 103.050 339.600 ;
        RECT 55.950 337.950 58.050 338.400 ;
        RECT 76.950 337.950 79.050 338.400 ;
        RECT 88.950 337.950 91.050 338.400 ;
        RECT 100.950 337.950 103.050 338.400 ;
        RECT 142.950 339.600 145.050 340.050 ;
        RECT 148.950 339.600 151.050 340.050 ;
        RECT 142.950 338.400 151.050 339.600 ;
        RECT 152.400 339.600 153.600 340.950 ;
        RECT 175.950 339.600 178.050 340.050 ;
        RECT 152.400 338.400 178.050 339.600 ;
        RECT 191.400 339.600 192.600 341.400 ;
        RECT 193.950 341.400 208.050 342.600 ;
        RECT 193.950 340.950 196.050 341.400 ;
        RECT 205.950 340.950 208.050 341.400 ;
        RECT 208.950 340.950 211.050 343.050 ;
        RECT 211.950 340.950 214.050 343.050 ;
        RECT 313.950 342.600 316.050 343.050 ;
        RECT 319.950 342.600 322.050 343.050 ;
        RECT 313.950 341.400 322.050 342.600 ;
        RECT 313.950 340.950 316.050 341.400 ;
        RECT 319.950 340.950 322.050 341.400 ;
        RECT 202.950 339.600 205.050 340.050 ;
        RECT 209.400 339.600 210.600 340.950 ;
        RECT 191.400 338.400 201.600 339.600 ;
        RECT 142.950 337.950 145.050 338.400 ;
        RECT 148.950 337.950 151.050 338.400 ;
        RECT 175.950 337.950 178.050 338.400 ;
        RECT 4.950 336.600 7.050 337.050 ;
        RECT 10.950 336.600 13.050 337.050 ;
        RECT 4.950 335.400 13.050 336.600 ;
        RECT 4.950 334.950 7.050 335.400 ;
        RECT 10.950 334.950 13.050 335.400 ;
        RECT 58.950 336.600 61.050 337.050 ;
        RECT 157.950 336.600 160.050 337.050 ;
        RECT 58.950 335.400 160.050 336.600 ;
        RECT 58.950 334.950 61.050 335.400 ;
        RECT 157.950 334.950 160.050 335.400 ;
        RECT 172.950 336.600 175.050 337.050 ;
        RECT 181.950 336.600 184.050 337.050 ;
        RECT 172.950 335.400 184.050 336.600 ;
        RECT 200.400 336.600 201.600 338.400 ;
        RECT 202.950 338.400 210.600 339.600 ;
        RECT 212.400 339.600 213.600 340.950 ;
        RECT 220.950 339.600 223.050 340.050 ;
        RECT 212.400 338.400 223.050 339.600 ;
        RECT 202.950 337.950 205.050 338.400 ;
        RECT 220.950 337.950 223.050 338.400 ;
        RECT 229.950 337.950 232.050 340.050 ;
        RECT 235.950 339.600 238.050 340.050 ;
        RECT 265.950 339.600 268.050 340.050 ;
        RECT 235.950 338.400 268.050 339.600 ;
        RECT 235.950 337.950 238.050 338.400 ;
        RECT 265.950 337.950 268.050 338.400 ;
        RECT 283.950 337.950 286.050 340.050 ;
        RECT 289.950 339.600 292.050 340.050 ;
        RECT 304.950 339.600 307.050 340.050 ;
        RECT 289.950 338.400 307.050 339.600 ;
        RECT 289.950 337.950 292.050 338.400 ;
        RECT 304.950 337.950 307.050 338.400 ;
        RECT 307.950 339.600 310.050 340.050 ;
        RECT 322.950 339.600 325.050 340.050 ;
        RECT 307.950 338.400 325.050 339.600 ;
        RECT 307.950 337.950 310.050 338.400 ;
        RECT 322.950 337.950 325.050 338.400 ;
        RECT 328.950 339.600 331.050 340.050 ;
        RECT 332.400 339.600 333.600 344.400 ;
        RECT 355.950 343.950 358.050 344.400 ;
        RECT 391.950 345.600 394.050 346.050 ;
        RECT 406.950 345.600 409.050 346.050 ;
        RECT 418.950 345.600 421.050 346.050 ;
        RECT 391.950 344.400 421.050 345.600 ;
        RECT 391.950 343.950 394.050 344.400 ;
        RECT 406.950 343.950 409.050 344.400 ;
        RECT 418.950 343.950 421.050 344.400 ;
        RECT 427.950 345.600 430.050 346.050 ;
        RECT 445.950 345.600 448.050 346.050 ;
        RECT 454.950 345.600 457.050 346.050 ;
        RECT 427.950 344.400 435.600 345.600 ;
        RECT 427.950 343.950 430.050 344.400 ;
        RECT 340.950 342.600 343.050 343.050 ;
        RECT 335.400 341.400 343.050 342.600 ;
        RECT 335.400 340.050 336.600 341.400 ;
        RECT 340.950 340.950 343.050 341.400 ;
        RECT 403.950 342.600 406.050 343.050 ;
        RECT 409.950 342.600 412.050 343.050 ;
        RECT 403.950 341.400 412.050 342.600 ;
        RECT 403.950 340.950 406.050 341.400 ;
        RECT 409.950 340.950 412.050 341.400 ;
        RECT 421.950 342.600 424.050 343.050 ;
        RECT 430.950 342.600 433.050 343.050 ;
        RECT 421.950 341.400 433.050 342.600 ;
        RECT 421.950 340.950 424.050 341.400 ;
        RECT 430.950 340.950 433.050 341.400 ;
        RECT 328.950 338.400 333.600 339.600 ;
        RECT 328.950 337.950 331.050 338.400 ;
        RECT 334.950 337.950 337.050 340.050 ;
        RECT 208.950 336.600 211.050 337.050 ;
        RECT 214.950 336.600 217.050 337.050 ;
        RECT 200.400 335.400 217.050 336.600 ;
        RECT 172.950 334.950 175.050 335.400 ;
        RECT 181.950 334.950 184.050 335.400 ;
        RECT 208.950 334.950 211.050 335.400 ;
        RECT 214.950 334.950 217.050 335.400 ;
        RECT 217.950 336.600 220.050 337.050 ;
        RECT 223.950 336.600 226.050 337.050 ;
        RECT 217.950 335.400 226.050 336.600 ;
        RECT 230.400 336.600 231.600 337.950 ;
        RECT 232.950 336.600 235.050 337.050 ;
        RECT 230.400 335.400 235.050 336.600 ;
        RECT 217.950 334.950 220.050 335.400 ;
        RECT 223.950 334.950 226.050 335.400 ;
        RECT 232.950 334.950 235.050 335.400 ;
        RECT 250.950 336.600 253.050 337.050 ;
        RECT 284.400 336.600 285.600 337.950 ;
        RECT 422.400 337.050 423.600 340.950 ;
        RECT 434.400 339.600 435.600 344.400 ;
        RECT 445.950 344.400 457.050 345.600 ;
        RECT 464.400 345.600 465.600 347.400 ;
        RECT 466.950 347.400 478.050 348.600 ;
        RECT 466.950 346.950 469.050 347.400 ;
        RECT 475.950 346.950 478.050 347.400 ;
        RECT 482.400 347.400 502.050 348.600 ;
        RECT 466.950 345.600 469.050 346.050 ;
        RECT 464.400 344.400 469.050 345.600 ;
        RECT 445.950 343.950 448.050 344.400 ;
        RECT 454.950 343.950 457.050 344.400 ;
        RECT 466.950 343.950 469.050 344.400 ;
        RECT 472.950 345.600 475.050 346.050 ;
        RECT 482.400 345.600 483.600 347.400 ;
        RECT 499.950 346.950 502.050 347.400 ;
        RECT 503.400 346.050 504.600 350.400 ;
        RECT 550.950 349.950 553.050 350.400 ;
        RECT 556.950 351.600 559.050 352.050 ;
        RECT 586.950 351.600 589.050 352.050 ;
        RECT 556.950 350.400 589.050 351.600 ;
        RECT 556.950 349.950 559.050 350.400 ;
        RECT 586.950 349.950 589.050 350.400 ;
        RECT 598.950 351.600 601.050 352.050 ;
        RECT 634.950 351.600 637.050 352.050 ;
        RECT 598.950 350.400 637.050 351.600 ;
        RECT 598.950 349.950 601.050 350.400 ;
        RECT 634.950 349.950 637.050 350.400 ;
        RECT 655.950 351.600 658.050 352.050 ;
        RECT 706.950 351.600 709.050 352.050 ;
        RECT 655.950 350.400 709.050 351.600 ;
        RECT 655.950 349.950 658.050 350.400 ;
        RECT 706.950 349.950 709.050 350.400 ;
        RECT 709.950 351.600 712.050 352.050 ;
        RECT 721.950 351.600 724.050 352.050 ;
        RECT 709.950 350.400 724.050 351.600 ;
        RECT 709.950 349.950 712.050 350.400 ;
        RECT 721.950 349.950 724.050 350.400 ;
        RECT 760.950 351.600 763.050 352.050 ;
        RECT 760.950 350.400 765.600 351.600 ;
        RECT 760.950 349.950 763.050 350.400 ;
        RECT 544.950 348.600 547.050 349.050 ;
        RECT 524.400 347.400 547.050 348.600 ;
        RECT 472.950 344.400 483.600 345.600 ;
        RECT 484.950 345.600 487.050 346.050 ;
        RECT 484.950 344.400 501.600 345.600 ;
        RECT 472.950 343.950 475.050 344.400 ;
        RECT 484.950 343.950 487.050 344.400 ;
        RECT 500.400 343.050 501.600 344.400 ;
        RECT 502.950 343.950 505.050 346.050 ;
        RECT 514.950 345.600 517.050 346.050 ;
        RECT 512.400 344.400 517.050 345.600 ;
        RECT 512.400 343.050 513.600 344.400 ;
        RECT 514.950 343.950 517.050 344.400 ;
        RECT 442.950 342.600 445.050 343.050 ;
        RECT 448.950 342.600 451.050 343.050 ;
        RECT 442.950 341.400 451.050 342.600 ;
        RECT 442.950 340.950 445.050 341.400 ;
        RECT 448.950 340.950 451.050 341.400 ;
        RECT 454.950 342.600 457.050 343.050 ;
        RECT 463.950 342.600 466.050 343.050 ;
        RECT 454.950 341.400 466.050 342.600 ;
        RECT 454.950 340.950 457.050 341.400 ;
        RECT 463.950 340.950 466.050 341.400 ;
        RECT 469.950 342.600 472.050 343.050 ;
        RECT 475.950 342.600 478.050 343.050 ;
        RECT 469.950 341.400 478.050 342.600 ;
        RECT 469.950 340.950 472.050 341.400 ;
        RECT 475.950 340.950 478.050 341.400 ;
        RECT 481.950 342.600 484.050 343.050 ;
        RECT 481.950 341.400 498.600 342.600 ;
        RECT 481.950 340.950 484.050 341.400 ;
        RECT 466.950 339.600 469.050 340.050 ;
        RECT 425.400 338.400 469.050 339.600 ;
        RECT 425.400 337.050 426.600 338.400 ;
        RECT 466.950 337.950 469.050 338.400 ;
        RECT 472.950 339.600 475.050 340.050 ;
        RECT 493.950 339.600 496.050 340.050 ;
        RECT 472.950 338.400 496.050 339.600 ;
        RECT 497.400 339.600 498.600 341.400 ;
        RECT 499.950 340.950 502.050 343.050 ;
        RECT 511.950 340.950 514.050 343.050 ;
        RECT 524.400 342.600 525.600 347.400 ;
        RECT 544.950 346.950 547.050 347.400 ;
        RECT 550.950 348.600 553.050 349.050 ;
        RECT 631.950 348.600 634.050 349.050 ;
        RECT 550.950 347.400 634.050 348.600 ;
        RECT 550.950 346.950 553.050 347.400 ;
        RECT 631.950 346.950 634.050 347.400 ;
        RECT 646.950 348.600 649.050 349.050 ;
        RECT 649.950 348.600 652.050 349.050 ;
        RECT 670.950 348.600 673.050 349.050 ;
        RECT 646.950 347.400 673.050 348.600 ;
        RECT 646.950 346.950 649.050 347.400 ;
        RECT 649.950 346.950 652.050 347.400 ;
        RECT 670.950 346.950 673.050 347.400 ;
        RECT 697.950 348.600 700.050 349.050 ;
        RECT 703.950 348.600 706.050 349.050 ;
        RECT 730.950 348.600 733.050 349.050 ;
        RECT 760.950 348.600 763.050 349.050 ;
        RECT 697.950 347.400 706.050 348.600 ;
        RECT 697.950 346.950 700.050 347.400 ;
        RECT 703.950 346.950 706.050 347.400 ;
        RECT 713.400 347.400 763.050 348.600 ;
        RECT 713.400 346.050 714.600 347.400 ;
        RECT 730.950 346.950 733.050 347.400 ;
        RECT 760.950 346.950 763.050 347.400 ;
        RECT 529.950 343.950 532.050 346.050 ;
        RECT 544.950 345.600 547.050 346.050 ;
        RECT 574.950 345.600 577.050 346.050 ;
        RECT 544.950 344.400 577.050 345.600 ;
        RECT 544.950 343.950 547.050 344.400 ;
        RECT 574.950 343.950 577.050 344.400 ;
        RECT 610.950 345.600 613.050 346.050 ;
        RECT 625.950 345.600 628.050 346.050 ;
        RECT 610.950 344.400 628.050 345.600 ;
        RECT 610.950 343.950 613.050 344.400 ;
        RECT 625.950 343.950 628.050 344.400 ;
        RECT 637.950 345.600 640.050 346.050 ;
        RECT 652.950 345.600 655.050 346.050 ;
        RECT 637.950 344.400 655.050 345.600 ;
        RECT 637.950 343.950 640.050 344.400 ;
        RECT 652.950 343.950 655.050 344.400 ;
        RECT 664.950 345.600 667.050 346.050 ;
        RECT 676.950 345.600 679.050 346.050 ;
        RECT 688.950 345.600 691.050 346.050 ;
        RECT 664.950 344.400 679.050 345.600 ;
        RECT 664.950 343.950 667.050 344.400 ;
        RECT 676.950 343.950 679.050 344.400 ;
        RECT 680.400 344.400 691.050 345.600 ;
        RECT 530.400 342.600 531.600 343.950 ;
        RECT 680.400 343.050 681.600 344.400 ;
        RECT 688.950 343.950 691.050 344.400 ;
        RECT 712.950 343.950 715.050 346.050 ;
        RECT 733.950 345.600 736.050 346.050 ;
        RECT 728.400 344.400 736.050 345.600 ;
        RECT 521.400 341.400 525.600 342.600 ;
        RECT 527.400 341.400 531.600 342.600 ;
        RECT 532.950 342.600 535.050 343.050 ;
        RECT 550.950 342.600 553.050 343.050 ;
        RECT 583.950 342.600 586.050 343.050 ;
        RECT 595.950 342.600 598.050 343.050 ;
        RECT 532.950 341.400 553.050 342.600 ;
        RECT 521.400 340.050 522.600 341.400 ;
        RECT 499.950 339.600 502.050 340.050 ;
        RECT 497.400 338.400 502.050 339.600 ;
        RECT 472.950 337.950 475.050 338.400 ;
        RECT 493.950 337.950 496.050 338.400 ;
        RECT 499.950 337.950 502.050 338.400 ;
        RECT 520.950 337.950 523.050 340.050 ;
        RECT 250.950 335.400 363.600 336.600 ;
        RECT 250.950 334.950 253.050 335.400 ;
        RECT 19.950 333.600 22.050 334.050 ;
        RECT 91.950 333.600 94.050 334.050 ;
        RECT 19.950 332.400 94.050 333.600 ;
        RECT 19.950 331.950 22.050 332.400 ;
        RECT 91.950 331.950 94.050 332.400 ;
        RECT 148.950 333.600 151.050 334.050 ;
        RECT 166.950 333.600 169.050 334.050 ;
        RECT 148.950 332.400 169.050 333.600 ;
        RECT 148.950 331.950 151.050 332.400 ;
        RECT 166.950 331.950 169.050 332.400 ;
        RECT 169.950 333.600 172.050 334.050 ;
        RECT 199.950 333.600 202.050 334.050 ;
        RECT 169.950 332.400 202.050 333.600 ;
        RECT 169.950 331.950 172.050 332.400 ;
        RECT 199.950 331.950 202.050 332.400 ;
        RECT 220.950 333.600 223.050 334.050 ;
        RECT 271.950 333.600 274.050 334.050 ;
        RECT 220.950 332.400 274.050 333.600 ;
        RECT 220.950 331.950 223.050 332.400 ;
        RECT 271.950 331.950 274.050 332.400 ;
        RECT 292.950 333.600 295.050 334.050 ;
        RECT 307.950 333.600 310.050 334.050 ;
        RECT 292.950 332.400 310.050 333.600 ;
        RECT 292.950 331.950 295.050 332.400 ;
        RECT 307.950 331.950 310.050 332.400 ;
        RECT 310.950 333.600 313.050 334.050 ;
        RECT 337.950 333.600 340.050 334.050 ;
        RECT 310.950 332.400 340.050 333.600 ;
        RECT 362.400 333.600 363.600 335.400 ;
        RECT 421.950 334.950 424.050 337.050 ;
        RECT 424.950 334.950 427.050 337.050 ;
        RECT 496.950 336.600 499.050 337.050 ;
        RECT 514.950 336.600 517.050 337.050 ;
        RECT 443.400 335.400 495.600 336.600 ;
        RECT 382.950 333.600 385.050 334.050 ;
        RECT 362.400 332.400 385.050 333.600 ;
        RECT 310.950 331.950 313.050 332.400 ;
        RECT 337.950 331.950 340.050 332.400 ;
        RECT 382.950 331.950 385.050 332.400 ;
        RECT 385.950 333.600 388.050 334.050 ;
        RECT 443.400 333.600 444.600 335.400 ;
        RECT 385.950 332.400 444.600 333.600 ;
        RECT 445.950 333.600 448.050 334.050 ;
        RECT 454.950 333.600 457.050 334.050 ;
        RECT 463.950 333.600 466.050 334.050 ;
        RECT 445.950 332.400 466.050 333.600 ;
        RECT 385.950 331.950 388.050 332.400 ;
        RECT 445.950 331.950 448.050 332.400 ;
        RECT 454.950 331.950 457.050 332.400 ;
        RECT 463.950 331.950 466.050 332.400 ;
        RECT 475.950 333.600 478.050 334.050 ;
        RECT 481.950 333.600 484.050 334.050 ;
        RECT 475.950 332.400 484.050 333.600 ;
        RECT 494.400 333.600 495.600 335.400 ;
        RECT 496.950 335.400 517.050 336.600 ;
        RECT 496.950 334.950 499.050 335.400 ;
        RECT 514.950 334.950 517.050 335.400 ;
        RECT 520.950 336.600 523.050 337.050 ;
        RECT 527.400 336.600 528.600 341.400 ;
        RECT 532.950 340.950 535.050 341.400 ;
        RECT 550.950 340.950 553.050 341.400 ;
        RECT 569.400 341.400 586.050 342.600 ;
        RECT 532.950 339.600 535.050 340.050 ;
        RECT 565.950 339.600 568.050 340.050 ;
        RECT 569.400 339.600 570.600 341.400 ;
        RECT 583.950 340.950 586.050 341.400 ;
        RECT 587.400 341.400 598.050 342.600 ;
        RECT 532.950 338.400 570.600 339.600 ;
        RECT 571.950 339.600 574.050 340.050 ;
        RECT 580.950 339.600 583.050 340.050 ;
        RECT 587.400 339.600 588.600 341.400 ;
        RECT 595.950 340.950 598.050 341.400 ;
        RECT 598.950 342.600 601.050 343.050 ;
        RECT 610.950 342.600 613.050 343.050 ;
        RECT 598.950 341.400 613.050 342.600 ;
        RECT 598.950 340.950 601.050 341.400 ;
        RECT 610.950 340.950 613.050 341.400 ;
        RECT 613.950 340.950 616.050 343.050 ;
        RECT 616.950 342.600 619.050 343.050 ;
        RECT 628.950 342.600 631.050 343.050 ;
        RECT 616.950 341.400 631.050 342.600 ;
        RECT 616.950 340.950 619.050 341.400 ;
        RECT 628.950 340.950 631.050 341.400 ;
        RECT 640.950 340.950 643.050 343.050 ;
        RECT 658.950 342.600 661.050 343.050 ;
        RECT 673.950 342.600 676.050 343.050 ;
        RECT 658.950 341.400 676.050 342.600 ;
        RECT 658.950 340.950 661.050 341.400 ;
        RECT 673.950 340.950 676.050 341.400 ;
        RECT 679.950 340.950 682.050 343.050 ;
        RECT 697.950 342.600 700.050 343.050 ;
        RECT 712.950 342.600 715.050 343.050 ;
        RECT 697.950 341.400 715.050 342.600 ;
        RECT 697.950 340.950 700.050 341.400 ;
        RECT 712.950 340.950 715.050 341.400 ;
        RECT 718.950 342.600 721.050 343.050 ;
        RECT 724.950 342.600 727.050 343.050 ;
        RECT 718.950 341.400 727.050 342.600 ;
        RECT 718.950 340.950 721.050 341.400 ;
        RECT 724.950 340.950 727.050 341.400 ;
        RECT 571.950 338.400 583.050 339.600 ;
        RECT 532.950 337.950 535.050 338.400 ;
        RECT 565.950 337.950 568.050 338.400 ;
        RECT 571.950 337.950 574.050 338.400 ;
        RECT 580.950 337.950 583.050 338.400 ;
        RECT 584.400 338.400 588.600 339.600 ;
        RECT 614.400 339.600 615.600 340.950 ;
        RECT 631.950 339.600 634.050 340.050 ;
        RECT 614.400 338.400 634.050 339.600 ;
        RECT 641.400 339.600 642.600 340.950 ;
        RECT 655.950 339.600 658.050 340.050 ;
        RECT 679.950 339.600 682.050 340.050 ;
        RECT 641.400 338.400 658.050 339.600 ;
        RECT 584.400 337.050 585.600 338.400 ;
        RECT 631.950 337.950 634.050 338.400 ;
        RECT 655.950 337.950 658.050 338.400 ;
        RECT 665.400 338.400 682.050 339.600 ;
        RECT 520.950 335.400 528.600 336.600 ;
        RECT 541.950 336.600 544.050 337.050 ;
        RECT 559.950 336.600 562.050 337.050 ;
        RECT 577.950 336.600 580.050 337.050 ;
        RECT 541.950 335.400 562.050 336.600 ;
        RECT 520.950 334.950 523.050 335.400 ;
        RECT 541.950 334.950 544.050 335.400 ;
        RECT 559.950 334.950 562.050 335.400 ;
        RECT 566.400 335.400 580.050 336.600 ;
        RECT 502.950 333.600 505.050 334.050 ;
        RECT 494.400 332.400 505.050 333.600 ;
        RECT 475.950 331.950 478.050 332.400 ;
        RECT 481.950 331.950 484.050 332.400 ;
        RECT 502.950 331.950 505.050 332.400 ;
        RECT 511.950 333.600 514.050 334.050 ;
        RECT 523.950 333.600 526.050 334.050 ;
        RECT 511.950 332.400 526.050 333.600 ;
        RECT 511.950 331.950 514.050 332.400 ;
        RECT 523.950 331.950 526.050 332.400 ;
        RECT 526.950 333.600 529.050 334.050 ;
        RECT 566.400 333.600 567.600 335.400 ;
        RECT 577.950 334.950 580.050 335.400 ;
        RECT 583.950 334.950 586.050 337.050 ;
        RECT 589.950 336.600 592.050 337.050 ;
        RECT 595.950 336.600 598.050 337.050 ;
        RECT 589.950 335.400 598.050 336.600 ;
        RECT 589.950 334.950 592.050 335.400 ;
        RECT 595.950 334.950 598.050 335.400 ;
        RECT 598.950 336.600 601.050 337.050 ;
        RECT 610.950 336.600 613.050 337.050 ;
        RECT 598.950 335.400 613.050 336.600 ;
        RECT 598.950 334.950 601.050 335.400 ;
        RECT 610.950 334.950 613.050 335.400 ;
        RECT 613.950 336.600 616.050 337.050 ;
        RECT 622.950 336.600 625.050 337.050 ;
        RECT 613.950 335.400 625.050 336.600 ;
        RECT 613.950 334.950 616.050 335.400 ;
        RECT 622.950 334.950 625.050 335.400 ;
        RECT 661.950 336.600 664.050 337.050 ;
        RECT 665.400 336.600 666.600 338.400 ;
        RECT 679.950 337.950 682.050 338.400 ;
        RECT 694.950 339.600 697.050 340.050 ;
        RECT 709.950 339.600 712.050 340.050 ;
        RECT 694.950 338.400 712.050 339.600 ;
        RECT 728.400 339.600 729.600 344.400 ;
        RECT 733.950 343.950 736.050 344.400 ;
        RECT 739.950 345.600 742.050 346.050 ;
        RECT 739.950 344.400 759.600 345.600 ;
        RECT 739.950 343.950 742.050 344.400 ;
        RECT 758.400 343.050 759.600 344.400 ;
        RECT 730.950 342.600 733.050 343.050 ;
        RECT 739.950 342.600 742.050 343.050 ;
        RECT 730.950 341.400 742.050 342.600 ;
        RECT 730.950 340.950 733.050 341.400 ;
        RECT 739.950 340.950 742.050 341.400 ;
        RECT 751.950 340.950 754.050 343.050 ;
        RECT 757.950 340.950 760.050 343.050 ;
        RECT 752.400 339.600 753.600 340.950 ;
        RECT 760.950 339.600 763.050 340.050 ;
        RECT 764.400 339.600 765.600 350.400 ;
        RECT 728.400 338.400 750.600 339.600 ;
        RECT 752.400 338.400 765.600 339.600 ;
        RECT 694.950 337.950 697.050 338.400 ;
        RECT 709.950 337.950 712.050 338.400 ;
        RECT 749.400 337.050 750.600 338.400 ;
        RECT 760.950 337.950 763.050 338.400 ;
        RECT 661.950 335.400 666.600 336.600 ;
        RECT 670.950 336.600 673.050 337.050 ;
        RECT 742.950 336.600 745.050 337.050 ;
        RECT 670.950 335.400 745.050 336.600 ;
        RECT 661.950 334.950 664.050 335.400 ;
        RECT 670.950 334.950 673.050 335.400 ;
        RECT 742.950 334.950 745.050 335.400 ;
        RECT 748.950 334.950 751.050 337.050 ;
        RECT 751.950 336.600 754.050 337.050 ;
        RECT 757.950 336.600 760.050 337.050 ;
        RECT 751.950 335.400 760.050 336.600 ;
        RECT 751.950 334.950 754.050 335.400 ;
        RECT 757.950 334.950 760.050 335.400 ;
        RECT 526.950 332.400 567.600 333.600 ;
        RECT 568.950 333.600 571.050 334.050 ;
        RECT 613.950 333.600 616.050 334.050 ;
        RECT 568.950 332.400 616.050 333.600 ;
        RECT 526.950 331.950 529.050 332.400 ;
        RECT 568.950 331.950 571.050 332.400 ;
        RECT 613.950 331.950 616.050 332.400 ;
        RECT 619.950 333.600 622.050 334.050 ;
        RECT 652.950 333.600 655.050 334.050 ;
        RECT 619.950 332.400 655.050 333.600 ;
        RECT 619.950 331.950 622.050 332.400 ;
        RECT 652.950 331.950 655.050 332.400 ;
        RECT 676.950 333.600 679.050 334.050 ;
        RECT 727.950 333.600 730.050 334.050 ;
        RECT 676.950 332.400 730.050 333.600 ;
        RECT 676.950 331.950 679.050 332.400 ;
        RECT 727.950 331.950 730.050 332.400 ;
        RECT 754.950 333.600 757.050 334.050 ;
        RECT 763.950 333.600 766.050 334.050 ;
        RECT 754.950 332.400 766.050 333.600 ;
        RECT 754.950 331.950 757.050 332.400 ;
        RECT 763.950 331.950 766.050 332.400 ;
        RECT 37.950 330.600 40.050 331.050 ;
        RECT 61.950 330.600 64.050 331.050 ;
        RECT 37.950 329.400 64.050 330.600 ;
        RECT 37.950 328.950 40.050 329.400 ;
        RECT 61.950 328.950 64.050 329.400 ;
        RECT 97.950 330.600 100.050 331.050 ;
        RECT 232.950 330.600 235.050 331.050 ;
        RECT 97.950 329.400 235.050 330.600 ;
        RECT 97.950 328.950 100.050 329.400 ;
        RECT 232.950 328.950 235.050 329.400 ;
        RECT 250.950 330.600 253.050 331.050 ;
        RECT 256.950 330.600 259.050 331.050 ;
        RECT 250.950 329.400 259.050 330.600 ;
        RECT 250.950 328.950 253.050 329.400 ;
        RECT 256.950 328.950 259.050 329.400 ;
        RECT 343.950 330.600 346.050 331.050 ;
        RECT 379.950 330.600 382.050 331.050 ;
        RECT 391.950 330.600 394.050 331.050 ;
        RECT 343.950 329.400 394.050 330.600 ;
        RECT 343.950 328.950 346.050 329.400 ;
        RECT 379.950 328.950 382.050 329.400 ;
        RECT 391.950 328.950 394.050 329.400 ;
        RECT 409.950 330.600 412.050 331.050 ;
        RECT 448.950 330.600 451.050 331.050 ;
        RECT 409.950 329.400 451.050 330.600 ;
        RECT 409.950 328.950 412.050 329.400 ;
        RECT 448.950 328.950 451.050 329.400 ;
        RECT 451.950 330.600 454.050 331.050 ;
        RECT 496.950 330.600 499.050 331.050 ;
        RECT 451.950 329.400 499.050 330.600 ;
        RECT 451.950 328.950 454.050 329.400 ;
        RECT 496.950 328.950 499.050 329.400 ;
        RECT 505.950 330.600 508.050 331.050 ;
        RECT 541.950 330.600 544.050 331.050 ;
        RECT 505.950 329.400 544.050 330.600 ;
        RECT 505.950 328.950 508.050 329.400 ;
        RECT 541.950 328.950 544.050 329.400 ;
        RECT 544.950 330.600 547.050 331.050 ;
        RECT 559.950 330.600 562.050 331.050 ;
        RECT 544.950 329.400 562.050 330.600 ;
        RECT 544.950 328.950 547.050 329.400 ;
        RECT 559.950 328.950 562.050 329.400 ;
        RECT 562.950 330.600 565.050 331.050 ;
        RECT 568.950 330.600 571.050 331.050 ;
        RECT 562.950 329.400 571.050 330.600 ;
        RECT 562.950 328.950 565.050 329.400 ;
        RECT 568.950 328.950 571.050 329.400 ;
        RECT 571.950 330.600 574.050 331.050 ;
        RECT 670.950 330.600 673.050 331.050 ;
        RECT 571.950 329.400 673.050 330.600 ;
        RECT 571.950 328.950 574.050 329.400 ;
        RECT 670.950 328.950 673.050 329.400 ;
        RECT 685.950 330.600 688.050 331.050 ;
        RECT 742.950 330.600 745.050 331.050 ;
        RECT 685.950 329.400 745.050 330.600 ;
        RECT 685.950 328.950 688.050 329.400 ;
        RECT 742.950 328.950 745.050 329.400 ;
        RECT 118.950 327.600 121.050 328.050 ;
        RECT 136.950 327.600 139.050 328.050 ;
        RECT 193.950 327.600 196.050 328.050 ;
        RECT 118.950 326.400 196.050 327.600 ;
        RECT 118.950 325.950 121.050 326.400 ;
        RECT 136.950 325.950 139.050 326.400 ;
        RECT 193.950 325.950 196.050 326.400 ;
        RECT 265.950 327.600 268.050 328.050 ;
        RECT 343.950 327.600 346.050 328.050 ;
        RECT 265.950 326.400 346.050 327.600 ;
        RECT 265.950 325.950 268.050 326.400 ;
        RECT 343.950 325.950 346.050 326.400 ;
        RECT 367.950 327.600 370.050 328.050 ;
        RECT 379.950 327.600 382.050 328.050 ;
        RECT 367.950 326.400 382.050 327.600 ;
        RECT 367.950 325.950 370.050 326.400 ;
        RECT 379.950 325.950 382.050 326.400 ;
        RECT 397.950 327.600 400.050 328.050 ;
        RECT 427.950 327.600 430.050 328.050 ;
        RECT 397.950 326.400 430.050 327.600 ;
        RECT 397.950 325.950 400.050 326.400 ;
        RECT 427.950 325.950 430.050 326.400 ;
        RECT 442.950 327.600 445.050 328.050 ;
        RECT 484.950 327.600 487.050 328.050 ;
        RECT 442.950 326.400 487.050 327.600 ;
        RECT 442.950 325.950 445.050 326.400 ;
        RECT 484.950 325.950 487.050 326.400 ;
        RECT 502.950 327.600 505.050 328.050 ;
        RECT 511.950 327.600 514.050 328.050 ;
        RECT 502.950 326.400 514.050 327.600 ;
        RECT 502.950 325.950 505.050 326.400 ;
        RECT 511.950 325.950 514.050 326.400 ;
        RECT 514.950 327.600 517.050 328.050 ;
        RECT 691.950 327.600 694.050 328.050 ;
        RECT 745.950 327.600 748.050 328.050 ;
        RECT 748.950 327.600 751.050 328.050 ;
        RECT 514.950 326.400 751.050 327.600 ;
        RECT 514.950 325.950 517.050 326.400 ;
        RECT 691.950 325.950 694.050 326.400 ;
        RECT 745.950 325.950 748.050 326.400 ;
        RECT 748.950 325.950 751.050 326.400 ;
        RECT 40.950 324.600 43.050 325.050 ;
        RECT 58.950 324.600 61.050 325.050 ;
        RECT 64.950 324.600 67.050 325.050 ;
        RECT 70.950 324.600 73.050 325.050 ;
        RECT 97.950 324.600 100.050 325.050 ;
        RECT 40.950 323.400 100.050 324.600 ;
        RECT 40.950 322.950 43.050 323.400 ;
        RECT 58.950 322.950 61.050 323.400 ;
        RECT 64.950 322.950 67.050 323.400 ;
        RECT 70.950 322.950 73.050 323.400 ;
        RECT 97.950 322.950 100.050 323.400 ;
        RECT 115.950 324.600 118.050 325.050 ;
        RECT 130.950 324.600 133.050 325.050 ;
        RECT 256.950 324.600 259.050 325.050 ;
        RECT 115.950 323.400 259.050 324.600 ;
        RECT 115.950 322.950 118.050 323.400 ;
        RECT 130.950 322.950 133.050 323.400 ;
        RECT 256.950 322.950 259.050 323.400 ;
        RECT 295.950 324.600 298.050 325.050 ;
        RECT 385.950 324.600 388.050 325.050 ;
        RECT 295.950 323.400 388.050 324.600 ;
        RECT 295.950 322.950 298.050 323.400 ;
        RECT 385.950 322.950 388.050 323.400 ;
        RECT 394.950 324.600 397.050 325.050 ;
        RECT 415.950 324.600 418.050 325.050 ;
        RECT 460.950 324.600 463.050 325.050 ;
        RECT 394.950 323.400 463.050 324.600 ;
        RECT 394.950 322.950 397.050 323.400 ;
        RECT 415.950 322.950 418.050 323.400 ;
        RECT 460.950 322.950 463.050 323.400 ;
        RECT 463.950 324.600 466.050 325.050 ;
        RECT 475.950 324.600 478.050 325.050 ;
        RECT 463.950 323.400 478.050 324.600 ;
        RECT 463.950 322.950 466.050 323.400 ;
        RECT 475.950 322.950 478.050 323.400 ;
        RECT 493.950 324.600 496.050 325.050 ;
        RECT 517.950 324.600 520.050 325.050 ;
        RECT 493.950 323.400 520.050 324.600 ;
        RECT 493.950 322.950 496.050 323.400 ;
        RECT 517.950 322.950 520.050 323.400 ;
        RECT 535.950 324.600 538.050 325.050 ;
        RECT 556.950 324.600 559.050 325.050 ;
        RECT 535.950 323.400 559.050 324.600 ;
        RECT 535.950 322.950 538.050 323.400 ;
        RECT 556.950 322.950 559.050 323.400 ;
        RECT 559.950 324.600 562.050 325.050 ;
        RECT 565.950 324.600 568.050 325.050 ;
        RECT 583.950 324.600 586.050 325.050 ;
        RECT 559.950 323.400 586.050 324.600 ;
        RECT 559.950 322.950 562.050 323.400 ;
        RECT 565.950 322.950 568.050 323.400 ;
        RECT 583.950 322.950 586.050 323.400 ;
        RECT 601.950 324.600 604.050 325.050 ;
        RECT 637.950 324.600 640.050 325.050 ;
        RECT 601.950 323.400 640.050 324.600 ;
        RECT 601.950 322.950 604.050 323.400 ;
        RECT 637.950 322.950 640.050 323.400 ;
        RECT 658.950 324.600 661.050 325.050 ;
        RECT 703.950 324.600 706.050 325.050 ;
        RECT 718.950 324.600 721.050 325.050 ;
        RECT 658.950 323.400 696.600 324.600 ;
        RECT 658.950 322.950 661.050 323.400 ;
        RECT 97.950 321.600 100.050 322.050 ;
        RECT 139.950 321.600 142.050 322.050 ;
        RECT 97.950 320.400 142.050 321.600 ;
        RECT 97.950 319.950 100.050 320.400 ;
        RECT 139.950 319.950 142.050 320.400 ;
        RECT 163.950 321.600 166.050 322.050 ;
        RECT 181.950 321.600 184.050 322.050 ;
        RECT 274.950 321.600 277.050 322.050 ;
        RECT 163.950 320.400 277.050 321.600 ;
        RECT 163.950 319.950 166.050 320.400 ;
        RECT 181.950 319.950 184.050 320.400 ;
        RECT 274.950 319.950 277.050 320.400 ;
        RECT 301.950 321.600 304.050 322.050 ;
        RECT 331.950 321.600 334.050 322.050 ;
        RECT 301.950 320.400 334.050 321.600 ;
        RECT 301.950 319.950 304.050 320.400 ;
        RECT 331.950 319.950 334.050 320.400 ;
        RECT 343.950 321.600 346.050 322.050 ;
        RECT 409.950 321.600 412.050 322.050 ;
        RECT 343.950 320.400 412.050 321.600 ;
        RECT 343.950 319.950 346.050 320.400 ;
        RECT 409.950 319.950 412.050 320.400 ;
        RECT 412.950 321.600 415.050 322.050 ;
        RECT 442.950 321.600 445.050 322.050 ;
        RECT 412.950 320.400 445.050 321.600 ;
        RECT 412.950 319.950 415.050 320.400 ;
        RECT 442.950 319.950 445.050 320.400 ;
        RECT 448.950 321.600 451.050 322.050 ;
        RECT 535.950 321.600 538.050 322.050 ;
        RECT 448.950 320.400 538.050 321.600 ;
        RECT 448.950 319.950 451.050 320.400 ;
        RECT 535.950 319.950 538.050 320.400 ;
        RECT 541.950 321.600 544.050 322.050 ;
        RECT 562.950 321.600 565.050 322.050 ;
        RECT 541.950 320.400 565.050 321.600 ;
        RECT 541.950 319.950 544.050 320.400 ;
        RECT 562.950 319.950 565.050 320.400 ;
        RECT 568.950 321.600 571.050 322.050 ;
        RECT 577.950 321.600 580.050 322.050 ;
        RECT 568.950 320.400 580.050 321.600 ;
        RECT 568.950 319.950 571.050 320.400 ;
        RECT 577.950 319.950 580.050 320.400 ;
        RECT 580.950 321.600 583.050 322.050 ;
        RECT 592.950 321.600 595.050 322.050 ;
        RECT 580.950 320.400 595.050 321.600 ;
        RECT 580.950 319.950 583.050 320.400 ;
        RECT 592.950 319.950 595.050 320.400 ;
        RECT 628.950 321.600 631.050 322.050 ;
        RECT 640.950 321.600 643.050 322.050 ;
        RECT 628.950 320.400 643.050 321.600 ;
        RECT 628.950 319.950 631.050 320.400 ;
        RECT 640.950 319.950 643.050 320.400 ;
        RECT 643.950 321.600 646.050 322.050 ;
        RECT 691.950 321.600 694.050 322.050 ;
        RECT 643.950 320.400 694.050 321.600 ;
        RECT 695.400 321.600 696.600 323.400 ;
        RECT 703.950 323.400 721.050 324.600 ;
        RECT 703.950 322.950 706.050 323.400 ;
        RECT 718.950 322.950 721.050 323.400 ;
        RECT 703.950 321.600 706.050 322.050 ;
        RECT 695.400 320.400 706.050 321.600 ;
        RECT 643.950 319.950 646.050 320.400 ;
        RECT 691.950 319.950 694.050 320.400 ;
        RECT 703.950 319.950 706.050 320.400 ;
        RECT 22.950 318.600 25.050 319.050 ;
        RECT 64.950 318.600 67.050 319.050 ;
        RECT 118.950 318.600 121.050 319.050 ;
        RECT 22.950 317.400 121.050 318.600 ;
        RECT 22.950 316.950 25.050 317.400 ;
        RECT 64.950 316.950 67.050 317.400 ;
        RECT 118.950 316.950 121.050 317.400 ;
        RECT 184.950 318.600 187.050 319.050 ;
        RECT 226.950 318.600 229.050 319.050 ;
        RECT 298.950 318.600 301.050 319.050 ;
        RECT 184.950 317.400 301.050 318.600 ;
        RECT 184.950 316.950 187.050 317.400 ;
        RECT 226.950 316.950 229.050 317.400 ;
        RECT 298.950 316.950 301.050 317.400 ;
        RECT 307.950 318.600 310.050 319.050 ;
        RECT 316.950 318.600 319.050 319.050 ;
        RECT 307.950 317.400 319.050 318.600 ;
        RECT 307.950 316.950 310.050 317.400 ;
        RECT 316.950 316.950 319.050 317.400 ;
        RECT 340.950 318.600 343.050 319.050 ;
        RECT 346.950 318.600 349.050 319.050 ;
        RECT 340.950 317.400 349.050 318.600 ;
        RECT 340.950 316.950 343.050 317.400 ;
        RECT 346.950 316.950 349.050 317.400 ;
        RECT 442.950 318.600 445.050 319.050 ;
        RECT 481.950 318.600 484.050 319.050 ;
        RECT 526.950 318.600 529.050 319.050 ;
        RECT 442.950 317.400 484.050 318.600 ;
        RECT 442.950 316.950 445.050 317.400 ;
        RECT 481.950 316.950 484.050 317.400 ;
        RECT 500.400 317.400 529.050 318.600 ;
        RECT 500.400 316.050 501.600 317.400 ;
        RECT 526.950 316.950 529.050 317.400 ;
        RECT 529.950 318.600 532.050 319.050 ;
        RECT 544.950 318.600 547.050 319.050 ;
        RECT 529.950 317.400 547.050 318.600 ;
        RECT 529.950 316.950 532.050 317.400 ;
        RECT 544.950 316.950 547.050 317.400 ;
        RECT 547.950 318.600 550.050 319.050 ;
        RECT 616.950 318.600 619.050 319.050 ;
        RECT 547.950 317.400 619.050 318.600 ;
        RECT 547.950 316.950 550.050 317.400 ;
        RECT 616.950 316.950 619.050 317.400 ;
        RECT 622.950 318.600 625.050 319.050 ;
        RECT 649.950 318.600 652.050 319.050 ;
        RECT 685.950 318.600 688.050 319.050 ;
        RECT 622.950 317.400 688.050 318.600 ;
        RECT 622.950 316.950 625.050 317.400 ;
        RECT 649.950 316.950 652.050 317.400 ;
        RECT 685.950 316.950 688.050 317.400 ;
        RECT 706.950 318.600 709.050 319.050 ;
        RECT 721.950 318.600 724.050 319.050 ;
        RECT 706.950 317.400 724.050 318.600 ;
        RECT 706.950 316.950 709.050 317.400 ;
        RECT 721.950 316.950 724.050 317.400 ;
        RECT 19.950 315.600 22.050 316.050 ;
        RECT 52.950 315.600 55.050 316.050 ;
        RECT 61.950 315.600 64.050 316.050 ;
        RECT 79.950 315.600 82.050 316.050 ;
        RECT 19.950 314.400 51.600 315.600 ;
        RECT 19.950 313.950 22.050 314.400 ;
        RECT 13.950 312.600 16.050 313.050 ;
        RECT 46.950 312.600 49.050 313.050 ;
        RECT 13.950 311.400 49.050 312.600 ;
        RECT 50.400 312.600 51.600 314.400 ;
        RECT 52.950 314.400 82.050 315.600 ;
        RECT 52.950 313.950 55.050 314.400 ;
        RECT 61.950 313.950 64.050 314.400 ;
        RECT 79.950 313.950 82.050 314.400 ;
        RECT 85.950 315.600 88.050 316.050 ;
        RECT 94.950 315.600 97.050 316.050 ;
        RECT 124.950 315.600 127.050 316.050 ;
        RECT 85.950 314.400 127.050 315.600 ;
        RECT 85.950 313.950 88.050 314.400 ;
        RECT 94.950 313.950 97.050 314.400 ;
        RECT 124.950 313.950 127.050 314.400 ;
        RECT 133.950 315.600 136.050 316.050 ;
        RECT 142.950 315.600 145.050 316.050 ;
        RECT 133.950 314.400 145.050 315.600 ;
        RECT 133.950 313.950 136.050 314.400 ;
        RECT 142.950 313.950 145.050 314.400 ;
        RECT 172.950 315.600 175.050 316.050 ;
        RECT 187.950 315.600 190.050 316.050 ;
        RECT 232.950 315.600 235.050 316.050 ;
        RECT 238.950 315.600 241.050 316.050 ;
        RECT 172.950 314.400 186.600 315.600 ;
        RECT 172.950 313.950 175.050 314.400 ;
        RECT 67.950 312.600 70.050 313.050 ;
        RECT 50.400 311.400 70.050 312.600 ;
        RECT 13.950 310.950 16.050 311.400 ;
        RECT 46.950 310.950 49.050 311.400 ;
        RECT 67.950 310.950 70.050 311.400 ;
        RECT 70.950 312.600 73.050 313.050 ;
        RECT 79.950 312.600 82.050 313.050 ;
        RECT 124.950 312.600 127.050 313.050 ;
        RECT 145.950 312.600 148.050 313.050 ;
        RECT 185.400 312.600 186.600 314.400 ;
        RECT 187.950 314.400 192.600 315.600 ;
        RECT 187.950 313.950 190.050 314.400 ;
        RECT 187.950 312.600 190.050 313.050 ;
        RECT 70.950 311.400 78.600 312.600 ;
        RECT 70.950 310.950 73.050 311.400 ;
        RECT 77.400 310.050 78.600 311.400 ;
        RECT 79.950 311.400 84.600 312.600 ;
        RECT 79.950 310.950 82.050 311.400 ;
        RECT 28.950 309.600 31.050 310.050 ;
        RECT 23.400 308.400 31.050 309.600 ;
        RECT 23.400 307.050 24.600 308.400 ;
        RECT 28.950 307.950 31.050 308.400 ;
        RECT 70.950 307.950 73.050 310.050 ;
        RECT 76.950 307.950 79.050 310.050 ;
        RECT 7.950 306.600 10.050 307.050 ;
        RECT 16.950 306.600 19.050 307.050 ;
        RECT 7.950 305.400 19.050 306.600 ;
        RECT 7.950 304.950 10.050 305.400 ;
        RECT 16.950 304.950 19.050 305.400 ;
        RECT 22.950 304.950 25.050 307.050 ;
        RECT 25.950 306.600 28.050 307.050 ;
        RECT 37.950 306.600 40.050 307.050 ;
        RECT 25.950 305.400 40.050 306.600 ;
        RECT 25.950 304.950 28.050 305.400 ;
        RECT 37.950 304.950 40.050 305.400 ;
        RECT 43.950 304.950 46.050 307.050 ;
        RECT 55.950 306.600 58.050 307.050 ;
        RECT 71.400 306.600 72.600 307.950 ;
        RECT 83.400 307.050 84.600 311.400 ;
        RECT 124.950 311.400 177.600 312.600 ;
        RECT 185.400 311.400 190.050 312.600 ;
        RECT 124.950 310.950 127.050 311.400 ;
        RECT 145.950 310.950 148.050 311.400 ;
        RECT 103.950 309.600 106.050 310.050 ;
        RECT 160.950 309.600 163.050 310.050 ;
        RECT 103.950 308.400 163.050 309.600 ;
        RECT 176.400 309.600 177.600 311.400 ;
        RECT 187.950 310.950 190.050 311.400 ;
        RECT 191.400 310.050 192.600 314.400 ;
        RECT 232.950 314.400 241.050 315.600 ;
        RECT 232.950 313.950 235.050 314.400 ;
        RECT 238.950 313.950 241.050 314.400 ;
        RECT 253.950 315.600 256.050 316.050 ;
        RECT 289.950 315.600 292.050 316.050 ;
        RECT 253.950 314.400 292.050 315.600 ;
        RECT 253.950 313.950 256.050 314.400 ;
        RECT 289.950 313.950 292.050 314.400 ;
        RECT 295.950 315.600 298.050 316.050 ;
        RECT 310.950 315.600 313.050 316.050 ;
        RECT 295.950 314.400 313.050 315.600 ;
        RECT 295.950 313.950 298.050 314.400 ;
        RECT 310.950 313.950 313.050 314.400 ;
        RECT 316.950 315.600 319.050 316.050 ;
        RECT 388.950 315.600 391.050 316.050 ;
        RECT 400.950 315.600 403.050 316.050 ;
        RECT 418.950 315.600 421.050 316.050 ;
        RECT 316.950 314.400 360.600 315.600 ;
        RECT 316.950 313.950 319.050 314.400 ;
        RECT 220.950 312.600 223.050 313.050 ;
        RECT 194.400 311.400 223.050 312.600 ;
        RECT 178.950 309.600 181.050 310.050 ;
        RECT 176.400 308.400 181.050 309.600 ;
        RECT 103.950 307.950 106.050 308.400 ;
        RECT 160.950 307.950 163.050 308.400 ;
        RECT 178.950 307.950 181.050 308.400 ;
        RECT 190.950 307.950 193.050 310.050 ;
        RECT 55.950 305.400 72.600 306.600 ;
        RECT 55.950 304.950 58.050 305.400 ;
        RECT 82.950 304.950 85.050 307.050 ;
        RECT 106.950 306.600 109.050 307.050 ;
        RECT 115.950 306.600 118.050 307.050 ;
        RECT 106.950 305.400 118.050 306.600 ;
        RECT 106.950 304.950 109.050 305.400 ;
        RECT 115.950 304.950 118.050 305.400 ;
        RECT 121.950 306.600 124.050 307.050 ;
        RECT 160.950 306.600 163.050 307.050 ;
        RECT 121.950 305.400 163.050 306.600 ;
        RECT 121.950 304.950 124.050 305.400 ;
        RECT 160.950 304.950 163.050 305.400 ;
        RECT 166.950 306.600 169.050 307.050 ;
        RECT 184.950 306.600 187.050 307.050 ;
        RECT 194.400 306.600 195.600 311.400 ;
        RECT 220.950 310.950 223.050 311.400 ;
        RECT 244.950 312.600 247.050 313.050 ;
        RECT 253.950 312.600 256.050 313.050 ;
        RECT 244.950 311.400 256.050 312.600 ;
        RECT 244.950 310.950 247.050 311.400 ;
        RECT 253.950 310.950 256.050 311.400 ;
        RECT 274.950 312.600 277.050 313.050 ;
        RECT 313.950 312.600 316.050 313.050 ;
        RECT 316.950 312.600 319.050 313.050 ;
        RECT 349.950 312.600 352.050 313.050 ;
        RECT 355.950 312.600 358.050 313.050 ;
        RECT 274.950 311.400 288.600 312.600 ;
        RECT 274.950 310.950 277.050 311.400 ;
        RECT 196.950 309.600 199.050 310.050 ;
        RECT 205.950 309.600 208.050 310.050 ;
        RECT 196.950 308.400 208.050 309.600 ;
        RECT 196.950 307.950 199.050 308.400 ;
        RECT 205.950 307.950 208.050 308.400 ;
        RECT 217.950 309.600 220.050 310.050 ;
        RECT 232.950 309.600 235.050 310.050 ;
        RECT 217.950 308.400 235.050 309.600 ;
        RECT 217.950 307.950 220.050 308.400 ;
        RECT 232.950 307.950 235.050 308.400 ;
        RECT 274.950 309.600 277.050 310.050 ;
        RECT 280.950 309.600 283.050 310.050 ;
        RECT 283.950 309.600 286.050 310.050 ;
        RECT 274.950 308.400 286.050 309.600 ;
        RECT 274.950 307.950 277.050 308.400 ;
        RECT 280.950 307.950 283.050 308.400 ;
        RECT 283.950 307.950 286.050 308.400 ;
        RECT 166.950 305.400 195.600 306.600 ;
        RECT 208.950 306.600 211.050 307.050 ;
        RECT 217.950 306.600 220.050 307.050 ;
        RECT 208.950 305.400 220.050 306.600 ;
        RECT 166.950 304.950 169.050 305.400 ;
        RECT 184.950 304.950 187.050 305.400 ;
        RECT 208.950 304.950 211.050 305.400 ;
        RECT 217.950 304.950 220.050 305.400 ;
        RECT 223.950 306.600 226.050 307.050 ;
        RECT 241.950 306.600 244.050 307.050 ;
        RECT 277.950 306.600 280.050 307.050 ;
        RECT 223.950 305.400 280.050 306.600 ;
        RECT 287.400 306.600 288.600 311.400 ;
        RECT 313.950 311.400 358.050 312.600 ;
        RECT 313.950 310.950 316.050 311.400 ;
        RECT 316.950 310.950 319.050 311.400 ;
        RECT 349.950 310.950 352.050 311.400 ;
        RECT 355.950 310.950 358.050 311.400 ;
        RECT 301.950 309.600 304.050 310.050 ;
        RECT 310.950 309.600 313.050 310.050 ;
        RECT 301.950 308.400 313.050 309.600 ;
        RECT 301.950 307.950 304.050 308.400 ;
        RECT 310.950 307.950 313.050 308.400 ;
        RECT 319.950 309.600 322.050 310.050 ;
        RECT 343.950 309.600 346.050 310.050 ;
        RECT 319.950 308.400 346.050 309.600 ;
        RECT 359.400 309.600 360.600 314.400 ;
        RECT 388.950 314.400 403.050 315.600 ;
        RECT 388.950 313.950 391.050 314.400 ;
        RECT 400.950 313.950 403.050 314.400 ;
        RECT 410.400 314.400 421.050 315.600 ;
        RECT 361.950 312.600 364.050 313.050 ;
        RECT 370.950 312.600 373.050 313.050 ;
        RECT 361.950 311.400 373.050 312.600 ;
        RECT 361.950 310.950 364.050 311.400 ;
        RECT 370.950 310.950 373.050 311.400 ;
        RECT 391.950 309.600 394.050 310.050 ;
        RECT 359.400 308.400 394.050 309.600 ;
        RECT 410.400 309.600 411.600 314.400 ;
        RECT 418.950 313.950 421.050 314.400 ;
        RECT 421.950 313.950 424.050 316.050 ;
        RECT 436.950 315.600 439.050 316.050 ;
        RECT 442.950 315.600 445.050 316.050 ;
        RECT 478.950 315.600 481.050 316.050 ;
        RECT 436.950 314.400 445.050 315.600 ;
        RECT 436.950 313.950 439.050 314.400 ;
        RECT 442.950 313.950 445.050 314.400 ;
        RECT 458.400 314.400 481.050 315.600 ;
        RECT 412.950 312.600 415.050 313.050 ;
        RECT 418.950 312.600 421.050 313.050 ;
        RECT 412.950 311.400 421.050 312.600 ;
        RECT 412.950 310.950 415.050 311.400 ;
        RECT 418.950 310.950 421.050 311.400 ;
        RECT 422.400 310.050 423.600 313.950 ;
        RECT 424.950 312.600 427.050 313.050 ;
        RECT 458.400 312.600 459.600 314.400 ;
        RECT 478.950 313.950 481.050 314.400 ;
        RECT 499.950 313.950 502.050 316.050 ;
        RECT 502.950 315.600 505.050 316.050 ;
        RECT 547.950 315.600 550.050 316.050 ;
        RECT 574.950 315.600 577.050 316.050 ;
        RECT 601.950 315.600 604.050 316.050 ;
        RECT 502.950 314.400 516.600 315.600 ;
        RECT 502.950 313.950 505.050 314.400 ;
        RECT 424.950 311.400 459.600 312.600 ;
        RECT 460.950 312.600 463.050 313.050 ;
        RECT 460.950 311.400 468.600 312.600 ;
        RECT 424.950 310.950 427.050 311.400 ;
        RECT 412.950 309.600 415.050 310.050 ;
        RECT 410.400 308.400 415.050 309.600 ;
        RECT 319.950 307.950 322.050 308.400 ;
        RECT 343.950 307.950 346.050 308.400 ;
        RECT 391.950 307.950 394.050 308.400 ;
        RECT 412.950 307.950 415.050 308.400 ;
        RECT 421.950 307.950 424.050 310.050 ;
        RECT 292.950 306.600 295.050 307.050 ;
        RECT 287.400 305.400 295.050 306.600 ;
        RECT 223.950 304.950 226.050 305.400 ;
        RECT 241.950 304.950 244.050 305.400 ;
        RECT 277.950 304.950 280.050 305.400 ;
        RECT 292.950 304.950 295.050 305.400 ;
        RECT 328.950 306.600 331.050 307.050 ;
        RECT 346.950 306.600 349.050 307.050 ;
        RECT 328.950 305.400 349.050 306.600 ;
        RECT 328.950 304.950 331.050 305.400 ;
        RECT 346.950 304.950 349.050 305.400 ;
        RECT 364.950 306.600 367.050 307.050 ;
        RECT 409.950 306.600 412.050 307.050 ;
        RECT 364.950 305.400 412.050 306.600 ;
        RECT 428.400 306.600 429.600 311.400 ;
        RECT 460.950 310.950 463.050 311.400 ;
        RECT 430.950 309.600 433.050 310.050 ;
        RECT 451.950 309.600 454.050 310.050 ;
        RECT 430.950 308.400 454.050 309.600 ;
        RECT 430.950 307.950 433.050 308.400 ;
        RECT 451.950 307.950 454.050 308.400 ;
        RECT 457.950 309.600 460.050 310.050 ;
        RECT 463.950 309.600 466.050 310.050 ;
        RECT 457.950 308.400 466.050 309.600 ;
        RECT 457.950 307.950 460.050 308.400 ;
        RECT 463.950 307.950 466.050 308.400 ;
        RECT 467.400 307.050 468.600 311.400 ;
        RECT 472.950 310.950 475.050 313.050 ;
        RECT 430.950 306.600 433.050 307.050 ;
        RECT 428.400 305.400 433.050 306.600 ;
        RECT 364.950 304.950 367.050 305.400 ;
        RECT 409.950 304.950 412.050 305.400 ;
        RECT 430.950 304.950 433.050 305.400 ;
        RECT 445.950 306.600 448.050 307.050 ;
        RECT 454.950 306.600 457.050 307.050 ;
        RECT 445.950 305.400 457.050 306.600 ;
        RECT 445.950 304.950 448.050 305.400 ;
        RECT 454.950 304.950 457.050 305.400 ;
        RECT 466.950 304.950 469.050 307.050 ;
        RECT 31.950 303.600 34.050 304.050 ;
        RECT 44.400 303.600 45.600 304.950 ;
        RECT 46.950 303.600 49.050 304.050 ;
        RECT 31.950 302.400 49.050 303.600 ;
        RECT 31.950 301.950 34.050 302.400 ;
        RECT 46.950 301.950 49.050 302.400 ;
        RECT 67.950 303.600 70.050 304.050 ;
        RECT 88.950 303.600 91.050 304.050 ;
        RECT 67.950 302.400 91.050 303.600 ;
        RECT 67.950 301.950 70.050 302.400 ;
        RECT 88.950 301.950 91.050 302.400 ;
        RECT 100.950 303.600 103.050 304.050 ;
        RECT 127.950 303.600 130.050 304.050 ;
        RECT 100.950 302.400 130.050 303.600 ;
        RECT 100.950 301.950 103.050 302.400 ;
        RECT 127.950 301.950 130.050 302.400 ;
        RECT 202.950 303.600 205.050 304.050 ;
        RECT 211.950 303.600 214.050 304.050 ;
        RECT 235.950 303.600 238.050 304.050 ;
        RECT 202.950 302.400 238.050 303.600 ;
        RECT 202.950 301.950 205.050 302.400 ;
        RECT 211.950 301.950 214.050 302.400 ;
        RECT 235.950 301.950 238.050 302.400 ;
        RECT 286.950 303.600 289.050 304.050 ;
        RECT 319.950 303.600 322.050 304.050 ;
        RECT 286.950 302.400 322.050 303.600 ;
        RECT 286.950 301.950 289.050 302.400 ;
        RECT 319.950 301.950 322.050 302.400 ;
        RECT 343.950 303.600 346.050 304.050 ;
        RECT 352.950 303.600 355.050 304.050 ;
        RECT 343.950 302.400 355.050 303.600 ;
        RECT 343.950 301.950 346.050 302.400 ;
        RECT 352.950 301.950 355.050 302.400 ;
        RECT 385.950 303.600 388.050 304.050 ;
        RECT 463.950 303.600 466.050 304.050 ;
        RECT 385.950 302.400 466.050 303.600 ;
        RECT 473.400 303.600 474.600 310.950 ;
        RECT 479.400 306.600 480.600 313.950 ;
        RECT 484.950 312.600 487.050 313.050 ;
        RECT 505.950 312.600 508.050 313.050 ;
        RECT 511.950 312.600 514.050 313.050 ;
        RECT 482.400 311.400 487.050 312.600 ;
        RECT 482.400 310.050 483.600 311.400 ;
        RECT 484.950 310.950 487.050 311.400 ;
        RECT 497.400 311.400 508.050 312.600 ;
        RECT 481.950 307.950 484.050 310.050 ;
        RECT 484.950 309.600 487.050 310.050 ;
        RECT 493.950 309.600 496.050 310.050 ;
        RECT 484.950 308.400 496.050 309.600 ;
        RECT 484.950 307.950 487.050 308.400 ;
        RECT 493.950 307.950 496.050 308.400 ;
        RECT 497.400 307.050 498.600 311.400 ;
        RECT 505.950 310.950 508.050 311.400 ;
        RECT 509.400 311.400 514.050 312.600 ;
        RECT 509.400 309.600 510.600 311.400 ;
        RECT 511.950 310.950 514.050 311.400 ;
        RECT 506.400 308.400 510.600 309.600 ;
        RECT 515.400 309.600 516.600 314.400 ;
        RECT 547.950 314.400 604.050 315.600 ;
        RECT 547.950 313.950 550.050 314.400 ;
        RECT 574.950 313.950 577.050 314.400 ;
        RECT 601.950 313.950 604.050 314.400 ;
        RECT 607.950 315.600 610.050 316.050 ;
        RECT 619.950 315.600 622.050 316.050 ;
        RECT 607.950 314.400 622.050 315.600 ;
        RECT 607.950 313.950 610.050 314.400 ;
        RECT 619.950 313.950 622.050 314.400 ;
        RECT 622.950 315.600 625.050 316.050 ;
        RECT 628.950 315.600 631.050 316.050 ;
        RECT 643.950 315.600 646.050 316.050 ;
        RECT 622.950 314.400 627.600 315.600 ;
        RECT 622.950 313.950 625.050 314.400 ;
        RECT 526.950 312.600 529.050 313.050 ;
        RECT 583.950 312.600 586.050 313.050 ;
        RECT 526.950 311.400 586.050 312.600 ;
        RECT 526.950 310.950 529.050 311.400 ;
        RECT 583.950 310.950 586.050 311.400 ;
        RECT 589.950 310.950 592.050 313.050 ;
        RECT 601.950 312.600 604.050 313.050 ;
        RECT 622.950 312.600 625.050 313.050 ;
        RECT 601.950 311.400 625.050 312.600 ;
        RECT 601.950 310.950 604.050 311.400 ;
        RECT 622.950 310.950 625.050 311.400 ;
        RECT 568.950 309.600 571.050 310.050 ;
        RECT 577.950 309.600 580.050 310.050 ;
        RECT 586.950 309.600 589.050 310.050 ;
        RECT 515.400 308.400 531.600 309.600 ;
        RECT 506.400 307.050 507.600 308.400 ;
        RECT 530.400 307.050 531.600 308.400 ;
        RECT 566.400 308.400 571.050 309.600 ;
        RECT 487.950 306.600 490.050 307.050 ;
        RECT 496.950 306.600 499.050 307.050 ;
        RECT 479.400 305.400 486.600 306.600 ;
        RECT 478.950 303.600 481.050 304.050 ;
        RECT 473.400 302.400 481.050 303.600 ;
        RECT 385.950 301.950 388.050 302.400 ;
        RECT 463.950 301.950 466.050 302.400 ;
        RECT 478.950 301.950 481.050 302.400 ;
        RECT 40.950 300.600 43.050 301.050 ;
        RECT 55.950 300.600 58.050 301.050 ;
        RECT 40.950 299.400 58.050 300.600 ;
        RECT 40.950 298.950 43.050 299.400 ;
        RECT 55.950 298.950 58.050 299.400 ;
        RECT 61.950 300.600 64.050 301.050 ;
        RECT 67.950 300.600 70.050 301.050 ;
        RECT 61.950 299.400 70.050 300.600 ;
        RECT 61.950 298.950 64.050 299.400 ;
        RECT 67.950 298.950 70.050 299.400 ;
        RECT 241.950 300.600 244.050 301.050 ;
        RECT 379.950 300.600 382.050 301.050 ;
        RECT 478.950 300.600 481.050 301.050 ;
        RECT 241.950 299.400 382.050 300.600 ;
        RECT 241.950 298.950 244.050 299.400 ;
        RECT 379.950 298.950 382.050 299.400 ;
        RECT 383.400 299.400 481.050 300.600 ;
        RECT 485.400 300.600 486.600 305.400 ;
        RECT 487.950 305.400 499.050 306.600 ;
        RECT 487.950 304.950 490.050 305.400 ;
        RECT 496.950 304.950 499.050 305.400 ;
        RECT 505.950 304.950 508.050 307.050 ;
        RECT 517.950 306.600 520.050 307.050 ;
        RECT 523.950 306.600 526.050 307.050 ;
        RECT 517.950 305.400 526.050 306.600 ;
        RECT 517.950 304.950 520.050 305.400 ;
        RECT 523.950 304.950 526.050 305.400 ;
        RECT 529.950 304.950 532.050 307.050 ;
        RECT 538.950 306.600 541.050 307.050 ;
        RECT 547.950 306.600 550.050 307.050 ;
        RECT 538.950 305.400 550.050 306.600 ;
        RECT 538.950 304.950 541.050 305.400 ;
        RECT 547.950 304.950 550.050 305.400 ;
        RECT 550.950 306.600 553.050 307.050 ;
        RECT 562.950 306.600 565.050 307.050 ;
        RECT 550.950 305.400 565.050 306.600 ;
        RECT 550.950 304.950 553.050 305.400 ;
        RECT 562.950 304.950 565.050 305.400 ;
        RECT 566.400 304.050 567.600 308.400 ;
        RECT 568.950 307.950 571.050 308.400 ;
        RECT 572.400 308.400 589.050 309.600 ;
        RECT 568.950 306.600 571.050 307.050 ;
        RECT 572.400 306.600 573.600 308.400 ;
        RECT 577.950 307.950 580.050 308.400 ;
        RECT 586.950 307.950 589.050 308.400 ;
        RECT 590.400 307.050 591.600 310.950 ;
        RECT 626.400 310.050 627.600 314.400 ;
        RECT 628.950 314.400 646.050 315.600 ;
        RECT 628.950 313.950 631.050 314.400 ;
        RECT 643.950 313.950 646.050 314.400 ;
        RECT 646.950 315.600 649.050 316.050 ;
        RECT 664.950 315.600 667.050 316.050 ;
        RECT 646.950 314.400 667.050 315.600 ;
        RECT 646.950 313.950 649.050 314.400 ;
        RECT 664.950 313.950 667.050 314.400 ;
        RECT 667.950 315.600 670.050 316.050 ;
        RECT 676.950 315.600 679.050 316.050 ;
        RECT 694.950 315.600 697.050 316.050 ;
        RECT 715.950 315.600 718.050 316.050 ;
        RECT 724.950 315.600 727.050 316.050 ;
        RECT 730.950 315.600 733.050 316.050 ;
        RECT 739.950 315.600 742.050 316.050 ;
        RECT 751.950 315.600 754.050 316.050 ;
        RECT 667.950 314.400 672.600 315.600 ;
        RECT 667.950 313.950 670.050 314.400 ;
        RECT 629.400 310.050 630.600 313.950 ;
        RECT 640.950 312.600 643.050 313.050 ;
        RECT 655.950 312.600 658.050 313.050 ;
        RECT 661.950 312.600 664.050 313.050 ;
        RECT 667.950 312.600 670.050 313.050 ;
        RECT 640.950 311.400 648.600 312.600 ;
        RECT 640.950 310.950 643.050 311.400 ;
        RECT 592.950 309.600 595.050 310.050 ;
        RECT 610.950 309.600 613.050 310.050 ;
        RECT 616.950 309.600 619.050 310.050 ;
        RECT 592.950 308.400 619.050 309.600 ;
        RECT 592.950 307.950 595.050 308.400 ;
        RECT 610.950 307.950 613.050 308.400 ;
        RECT 616.950 307.950 619.050 308.400 ;
        RECT 625.950 307.950 628.050 310.050 ;
        RECT 628.950 307.950 631.050 310.050 ;
        RECT 631.950 309.600 634.050 310.050 ;
        RECT 643.950 309.600 646.050 310.050 ;
        RECT 631.950 308.400 646.050 309.600 ;
        RECT 631.950 307.950 634.050 308.400 ;
        RECT 643.950 307.950 646.050 308.400 ;
        RECT 568.950 305.400 573.600 306.600 ;
        RECT 568.950 304.950 571.050 305.400 ;
        RECT 589.950 304.950 592.050 307.050 ;
        RECT 592.950 306.600 595.050 307.050 ;
        RECT 640.950 306.600 643.050 307.050 ;
        RECT 592.950 305.400 643.050 306.600 ;
        RECT 647.400 306.600 648.600 311.400 ;
        RECT 655.950 311.400 670.050 312.600 ;
        RECT 655.950 310.950 658.050 311.400 ;
        RECT 661.950 310.950 664.050 311.400 ;
        RECT 667.950 310.950 670.050 311.400 ;
        RECT 664.950 309.600 667.050 310.050 ;
        RECT 664.950 308.400 669.600 309.600 ;
        RECT 664.950 307.950 667.050 308.400 ;
        RECT 655.950 306.600 658.050 307.050 ;
        RECT 647.400 305.400 658.050 306.600 ;
        RECT 592.950 304.950 595.050 305.400 ;
        RECT 640.950 304.950 643.050 305.400 ;
        RECT 655.950 304.950 658.050 305.400 ;
        RECT 487.950 303.600 490.050 304.050 ;
        RECT 502.950 303.600 505.050 304.050 ;
        RECT 511.950 303.600 514.050 304.050 ;
        RECT 553.950 303.600 556.050 304.050 ;
        RECT 487.950 302.400 556.050 303.600 ;
        RECT 487.950 301.950 490.050 302.400 ;
        RECT 502.950 301.950 505.050 302.400 ;
        RECT 511.950 301.950 514.050 302.400 ;
        RECT 553.950 301.950 556.050 302.400 ;
        RECT 565.950 301.950 568.050 304.050 ;
        RECT 586.950 303.600 589.050 304.050 ;
        RECT 634.950 303.600 637.050 304.050 ;
        RECT 586.950 302.400 637.050 303.600 ;
        RECT 586.950 301.950 589.050 302.400 ;
        RECT 634.950 301.950 637.050 302.400 ;
        RECT 637.950 303.600 640.050 304.050 ;
        RECT 643.950 303.600 646.050 304.050 ;
        RECT 637.950 302.400 646.050 303.600 ;
        RECT 668.400 303.600 669.600 308.400 ;
        RECT 671.400 307.050 672.600 314.400 ;
        RECT 676.950 314.400 693.600 315.600 ;
        RECT 676.950 313.950 679.050 314.400 ;
        RECT 692.400 312.600 693.600 314.400 ;
        RECT 694.950 314.400 711.600 315.600 ;
        RECT 694.950 313.950 697.050 314.400 ;
        RECT 697.950 312.600 700.050 313.050 ;
        RECT 692.400 311.400 700.050 312.600 ;
        RECT 697.950 310.950 700.050 311.400 ;
        RECT 706.950 310.950 709.050 313.050 ;
        RECT 710.400 312.600 711.600 314.400 ;
        RECT 715.950 314.400 733.050 315.600 ;
        RECT 715.950 313.950 718.050 314.400 ;
        RECT 724.950 313.950 727.050 314.400 ;
        RECT 730.950 313.950 733.050 314.400 ;
        RECT 734.400 314.400 742.050 315.600 ;
        RECT 734.400 312.600 735.600 314.400 ;
        RECT 739.950 313.950 742.050 314.400 ;
        RECT 749.400 314.400 754.050 315.600 ;
        RECT 710.400 311.400 735.600 312.600 ;
        RECT 673.950 309.600 676.050 310.050 ;
        RECT 691.950 309.600 694.050 310.050 ;
        RECT 673.950 308.400 694.050 309.600 ;
        RECT 673.950 307.950 676.050 308.400 ;
        RECT 691.950 307.950 694.050 308.400 ;
        RECT 697.950 307.950 700.050 310.050 ;
        RECT 670.950 304.950 673.050 307.050 ;
        RECT 679.950 306.600 682.050 307.050 ;
        RECT 694.950 306.600 697.050 307.050 ;
        RECT 679.950 305.400 697.050 306.600 ;
        RECT 698.400 306.600 699.600 307.950 ;
        RECT 700.950 306.600 703.050 307.050 ;
        RECT 698.400 305.400 703.050 306.600 ;
        RECT 679.950 304.950 682.050 305.400 ;
        RECT 694.950 304.950 697.050 305.400 ;
        RECT 700.950 304.950 703.050 305.400 ;
        RECT 676.950 303.600 679.050 304.050 ;
        RECT 668.400 302.400 679.050 303.600 ;
        RECT 637.950 301.950 640.050 302.400 ;
        RECT 643.950 301.950 646.050 302.400 ;
        RECT 676.950 301.950 679.050 302.400 ;
        RECT 517.950 300.600 520.050 301.050 ;
        RECT 485.400 299.400 520.050 300.600 ;
        RECT 34.950 297.600 37.050 298.050 ;
        RECT 100.950 297.600 103.050 298.050 ;
        RECT 34.950 296.400 103.050 297.600 ;
        RECT 34.950 295.950 37.050 296.400 ;
        RECT 100.950 295.950 103.050 296.400 ;
        RECT 229.950 297.600 232.050 298.050 ;
        RECT 256.950 297.600 259.050 298.050 ;
        RECT 229.950 296.400 259.050 297.600 ;
        RECT 229.950 295.950 232.050 296.400 ;
        RECT 256.950 295.950 259.050 296.400 ;
        RECT 274.950 297.600 277.050 298.050 ;
        RECT 383.400 297.600 384.600 299.400 ;
        RECT 478.950 298.950 481.050 299.400 ;
        RECT 517.950 298.950 520.050 299.400 ;
        RECT 520.950 300.600 523.050 301.050 ;
        RECT 526.950 300.600 529.050 301.050 ;
        RECT 520.950 299.400 529.050 300.600 ;
        RECT 520.950 298.950 523.050 299.400 ;
        RECT 526.950 298.950 529.050 299.400 ;
        RECT 544.950 300.600 547.050 301.050 ;
        RECT 580.950 300.600 583.050 301.050 ;
        RECT 544.950 299.400 583.050 300.600 ;
        RECT 544.950 298.950 547.050 299.400 ;
        RECT 580.950 298.950 583.050 299.400 ;
        RECT 616.950 300.600 619.050 301.050 ;
        RECT 664.950 300.600 667.050 301.050 ;
        RECT 616.950 299.400 667.050 300.600 ;
        RECT 616.950 298.950 619.050 299.400 ;
        RECT 664.950 298.950 667.050 299.400 ;
        RECT 670.950 300.600 673.050 301.050 ;
        RECT 691.950 300.600 694.050 301.050 ;
        RECT 707.400 300.600 708.600 310.950 ;
        RECT 710.400 306.600 711.600 311.400 ;
        RECT 736.950 310.950 739.050 313.050 ;
        RECT 718.950 307.950 721.050 310.050 ;
        RECT 721.950 309.600 724.050 310.050 ;
        RECT 727.950 309.600 730.050 310.050 ;
        RECT 721.950 308.400 730.050 309.600 ;
        RECT 721.950 307.950 724.050 308.400 ;
        RECT 727.950 307.950 730.050 308.400 ;
        RECT 715.950 306.600 718.050 307.050 ;
        RECT 710.400 305.400 718.050 306.600 ;
        RECT 719.400 306.600 720.600 307.950 ;
        RECT 733.950 306.600 736.050 307.050 ;
        RECT 719.400 305.400 736.050 306.600 ;
        RECT 737.400 306.600 738.600 310.950 ;
        RECT 749.400 310.050 750.600 314.400 ;
        RECT 751.950 313.950 754.050 314.400 ;
        RECT 754.950 312.600 757.050 313.050 ;
        RECT 754.950 311.400 765.600 312.600 ;
        RECT 754.950 310.950 757.050 311.400 ;
        RECT 739.950 309.600 742.050 310.050 ;
        RECT 745.950 309.600 748.050 310.050 ;
        RECT 739.950 308.400 748.050 309.600 ;
        RECT 739.950 307.950 742.050 308.400 ;
        RECT 745.950 307.950 748.050 308.400 ;
        RECT 748.950 307.950 751.050 310.050 ;
        RECT 751.950 306.600 754.050 307.050 ;
        RECT 737.400 305.400 754.050 306.600 ;
        RECT 715.950 304.950 718.050 305.400 ;
        RECT 733.950 304.950 736.050 305.400 ;
        RECT 751.950 304.950 754.050 305.400 ;
        RECT 754.950 306.600 757.050 307.050 ;
        RECT 760.950 306.600 763.050 307.050 ;
        RECT 754.950 305.400 763.050 306.600 ;
        RECT 754.950 304.950 757.050 305.400 ;
        RECT 760.950 304.950 763.050 305.400 ;
        RECT 730.950 303.600 733.050 304.050 ;
        RECT 742.950 303.600 745.050 304.050 ;
        RECT 730.950 302.400 745.050 303.600 ;
        RECT 730.950 301.950 733.050 302.400 ;
        RECT 742.950 301.950 745.050 302.400 ;
        RECT 745.950 303.600 748.050 304.050 ;
        RECT 764.400 303.600 765.600 311.400 ;
        RECT 745.950 302.400 765.600 303.600 ;
        RECT 745.950 301.950 748.050 302.400 ;
        RECT 670.950 299.400 687.600 300.600 ;
        RECT 670.950 298.950 673.050 299.400 ;
        RECT 274.950 296.400 384.600 297.600 ;
        RECT 433.950 297.600 436.050 298.050 ;
        RECT 508.950 297.600 511.050 298.050 ;
        RECT 571.950 297.600 574.050 298.050 ;
        RECT 433.950 296.400 574.050 297.600 ;
        RECT 274.950 295.950 277.050 296.400 ;
        RECT 433.950 295.950 436.050 296.400 ;
        RECT 508.950 295.950 511.050 296.400 ;
        RECT 571.950 295.950 574.050 296.400 ;
        RECT 574.950 297.600 577.050 298.050 ;
        RECT 592.950 297.600 595.050 298.050 ;
        RECT 574.950 296.400 595.050 297.600 ;
        RECT 574.950 295.950 577.050 296.400 ;
        RECT 592.950 295.950 595.050 296.400 ;
        RECT 598.950 297.600 601.050 298.050 ;
        RECT 604.950 297.600 607.050 298.050 ;
        RECT 634.950 297.600 637.050 298.050 ;
        RECT 598.950 296.400 637.050 297.600 ;
        RECT 598.950 295.950 601.050 296.400 ;
        RECT 604.950 295.950 607.050 296.400 ;
        RECT 634.950 295.950 637.050 296.400 ;
        RECT 640.950 297.600 643.050 298.050 ;
        RECT 682.950 297.600 685.050 298.050 ;
        RECT 640.950 296.400 685.050 297.600 ;
        RECT 686.400 297.600 687.600 299.400 ;
        RECT 691.950 299.400 708.600 300.600 ;
        RECT 691.950 298.950 694.050 299.400 ;
        RECT 712.950 297.600 715.050 298.050 ;
        RECT 686.400 296.400 715.050 297.600 ;
        RECT 640.950 295.950 643.050 296.400 ;
        RECT 682.950 295.950 685.050 296.400 ;
        RECT 712.950 295.950 715.050 296.400 ;
        RECT 724.950 297.600 727.050 298.050 ;
        RECT 757.950 297.600 760.050 298.050 ;
        RECT 724.950 296.400 760.050 297.600 ;
        RECT 724.950 295.950 727.050 296.400 ;
        RECT 757.950 295.950 760.050 296.400 ;
        RECT 259.950 294.600 262.050 295.050 ;
        RECT 268.950 294.600 271.050 295.050 ;
        RECT 352.950 294.600 355.050 295.050 ;
        RECT 259.950 293.400 355.050 294.600 ;
        RECT 259.950 292.950 262.050 293.400 ;
        RECT 268.950 292.950 271.050 293.400 ;
        RECT 352.950 292.950 355.050 293.400 ;
        RECT 379.950 294.600 382.050 295.050 ;
        RECT 397.950 294.600 400.050 295.050 ;
        RECT 436.950 294.600 439.050 295.050 ;
        RECT 469.950 294.600 472.050 295.050 ;
        RECT 379.950 293.400 472.050 294.600 ;
        RECT 379.950 292.950 382.050 293.400 ;
        RECT 397.950 292.950 400.050 293.400 ;
        RECT 436.950 292.950 439.050 293.400 ;
        RECT 469.950 292.950 472.050 293.400 ;
        RECT 475.950 294.600 478.050 295.050 ;
        RECT 511.950 294.600 514.050 295.050 ;
        RECT 535.950 294.600 538.050 295.050 ;
        RECT 475.950 293.400 514.050 294.600 ;
        RECT 475.950 292.950 478.050 293.400 ;
        RECT 511.950 292.950 514.050 293.400 ;
        RECT 530.400 293.400 538.050 294.600 ;
        RECT 172.950 291.600 175.050 292.050 ;
        RECT 262.950 291.600 265.050 292.050 ;
        RECT 172.950 290.400 265.050 291.600 ;
        RECT 172.950 289.950 175.050 290.400 ;
        RECT 262.950 289.950 265.050 290.400 ;
        RECT 277.950 291.600 280.050 292.050 ;
        RECT 406.950 291.600 409.050 292.050 ;
        RECT 277.950 290.400 409.050 291.600 ;
        RECT 277.950 289.950 280.050 290.400 ;
        RECT 406.950 289.950 409.050 290.400 ;
        RECT 412.950 291.600 415.050 292.050 ;
        RECT 445.950 291.600 448.050 292.050 ;
        RECT 530.400 291.600 531.600 293.400 ;
        RECT 535.950 292.950 538.050 293.400 ;
        RECT 556.950 294.600 559.050 295.050 ;
        RECT 619.950 294.600 622.050 295.050 ;
        RECT 556.950 293.400 622.050 294.600 ;
        RECT 556.950 292.950 559.050 293.400 ;
        RECT 619.950 292.950 622.050 293.400 ;
        RECT 631.950 294.600 634.050 295.050 ;
        RECT 637.950 294.600 640.050 295.050 ;
        RECT 631.950 293.400 640.050 294.600 ;
        RECT 631.950 292.950 634.050 293.400 ;
        RECT 637.950 292.950 640.050 293.400 ;
        RECT 679.950 294.600 682.050 295.050 ;
        RECT 706.950 294.600 709.050 295.050 ;
        RECT 679.950 293.400 709.050 294.600 ;
        RECT 679.950 292.950 682.050 293.400 ;
        RECT 706.950 292.950 709.050 293.400 ;
        RECT 709.950 294.600 712.050 295.050 ;
        RECT 760.950 294.600 763.050 295.050 ;
        RECT 709.950 293.400 763.050 294.600 ;
        RECT 709.950 292.950 712.050 293.400 ;
        RECT 760.950 292.950 763.050 293.400 ;
        RECT 412.950 290.400 531.600 291.600 ;
        RECT 532.950 291.600 535.050 292.050 ;
        RECT 574.950 291.600 577.050 292.050 ;
        RECT 532.950 290.400 577.050 291.600 ;
        RECT 412.950 289.950 415.050 290.400 ;
        RECT 445.950 289.950 448.050 290.400 ;
        RECT 532.950 289.950 535.050 290.400 ;
        RECT 574.950 289.950 577.050 290.400 ;
        RECT 583.950 291.600 586.050 292.050 ;
        RECT 610.950 291.600 613.050 292.050 ;
        RECT 583.950 290.400 613.050 291.600 ;
        RECT 583.950 289.950 586.050 290.400 ;
        RECT 610.950 289.950 613.050 290.400 ;
        RECT 619.950 291.600 622.050 292.050 ;
        RECT 643.950 291.600 646.050 292.050 ;
        RECT 745.950 291.600 748.050 292.050 ;
        RECT 619.950 290.400 748.050 291.600 ;
        RECT 619.950 289.950 622.050 290.400 ;
        RECT 643.950 289.950 646.050 290.400 ;
        RECT 745.950 289.950 748.050 290.400 ;
        RECT 127.950 288.600 130.050 289.050 ;
        RECT 187.950 288.600 190.050 289.050 ;
        RECT 286.950 288.600 289.050 289.050 ;
        RECT 127.950 287.400 289.050 288.600 ;
        RECT 127.950 286.950 130.050 287.400 ;
        RECT 187.950 286.950 190.050 287.400 ;
        RECT 286.950 286.950 289.050 287.400 ;
        RECT 289.950 288.600 292.050 289.050 ;
        RECT 298.950 288.600 301.050 289.050 ;
        RECT 289.950 287.400 301.050 288.600 ;
        RECT 289.950 286.950 292.050 287.400 ;
        RECT 298.950 286.950 301.050 287.400 ;
        RECT 367.950 288.600 370.050 289.050 ;
        RECT 388.950 288.600 391.050 289.050 ;
        RECT 367.950 287.400 391.050 288.600 ;
        RECT 367.950 286.950 370.050 287.400 ;
        RECT 388.950 286.950 391.050 287.400 ;
        RECT 439.950 288.600 442.050 289.050 ;
        RECT 448.950 288.600 451.050 289.050 ;
        RECT 439.950 287.400 451.050 288.600 ;
        RECT 439.950 286.950 442.050 287.400 ;
        RECT 448.950 286.950 451.050 287.400 ;
        RECT 451.950 288.600 454.050 289.050 ;
        RECT 475.950 288.600 478.050 289.050 ;
        RECT 541.950 288.600 544.050 289.050 ;
        RECT 451.950 287.400 544.050 288.600 ;
        RECT 451.950 286.950 454.050 287.400 ;
        RECT 475.950 286.950 478.050 287.400 ;
        RECT 541.950 286.950 544.050 287.400 ;
        RECT 577.950 288.600 580.050 289.050 ;
        RECT 646.950 288.600 649.050 289.050 ;
        RECT 652.950 288.600 655.050 289.050 ;
        RECT 577.950 287.400 649.050 288.600 ;
        RECT 577.950 286.950 580.050 287.400 ;
        RECT 646.950 286.950 649.050 287.400 ;
        RECT 650.400 287.400 655.050 288.600 ;
        RECT 163.950 285.600 166.050 286.050 ;
        RECT 169.950 285.600 172.050 286.050 ;
        RECT 295.950 285.600 298.050 286.050 ;
        RECT 163.950 284.400 298.050 285.600 ;
        RECT 163.950 283.950 166.050 284.400 ;
        RECT 169.950 283.950 172.050 284.400 ;
        RECT 295.950 283.950 298.050 284.400 ;
        RECT 310.950 285.600 313.050 286.050 ;
        RECT 325.950 285.600 328.050 286.050 ;
        RECT 379.950 285.600 382.050 286.050 ;
        RECT 589.950 285.600 592.050 286.050 ;
        RECT 310.950 284.400 592.050 285.600 ;
        RECT 310.950 283.950 313.050 284.400 ;
        RECT 325.950 283.950 328.050 284.400 ;
        RECT 379.950 283.950 382.050 284.400 ;
        RECT 589.950 283.950 592.050 284.400 ;
        RECT 643.950 285.600 646.050 286.050 ;
        RECT 650.400 285.600 651.600 287.400 ;
        RECT 652.950 286.950 655.050 287.400 ;
        RECT 673.950 288.600 676.050 289.050 ;
        RECT 727.950 288.600 730.050 289.050 ;
        RECT 673.950 287.400 730.050 288.600 ;
        RECT 673.950 286.950 676.050 287.400 ;
        RECT 727.950 286.950 730.050 287.400 ;
        RECT 643.950 284.400 651.600 285.600 ;
        RECT 664.950 285.600 667.050 286.050 ;
        RECT 727.950 285.600 730.050 286.050 ;
        RECT 664.950 284.400 730.050 285.600 ;
        RECT 643.950 283.950 646.050 284.400 ;
        RECT 664.950 283.950 667.050 284.400 ;
        RECT 727.950 283.950 730.050 284.400 ;
        RECT 199.950 282.600 202.050 283.050 ;
        RECT 211.950 282.600 214.050 283.050 ;
        RECT 232.950 282.600 235.050 283.050 ;
        RECT 199.950 281.400 235.050 282.600 ;
        RECT 199.950 280.950 202.050 281.400 ;
        RECT 211.950 280.950 214.050 281.400 ;
        RECT 232.950 280.950 235.050 281.400 ;
        RECT 286.950 282.600 289.050 283.050 ;
        RECT 304.950 282.600 307.050 283.050 ;
        RECT 286.950 281.400 307.050 282.600 ;
        RECT 286.950 280.950 289.050 281.400 ;
        RECT 304.950 280.950 307.050 281.400 ;
        RECT 355.950 282.600 358.050 283.050 ;
        RECT 370.950 282.600 373.050 283.050 ;
        RECT 376.950 282.600 379.050 283.050 ;
        RECT 355.950 281.400 369.600 282.600 ;
        RECT 355.950 280.950 358.050 281.400 ;
        RECT 55.950 279.600 58.050 280.050 ;
        RECT 23.400 278.400 58.050 279.600 ;
        RECT 7.950 271.950 10.050 274.050 ;
        RECT 13.950 273.600 16.050 274.050 ;
        RECT 13.950 272.400 21.600 273.600 ;
        RECT 13.950 271.950 16.050 272.400 ;
        RECT 8.400 268.050 9.600 271.950 ;
        RECT 10.950 270.600 13.050 271.050 ;
        RECT 16.950 270.600 19.050 271.050 ;
        RECT 10.950 269.400 19.050 270.600 ;
        RECT 10.950 268.950 13.050 269.400 ;
        RECT 16.950 268.950 19.050 269.400 ;
        RECT 20.400 268.050 21.600 272.400 ;
        RECT 23.400 271.050 24.600 278.400 ;
        RECT 55.950 277.950 58.050 278.400 ;
        RECT 220.950 279.600 223.050 280.050 ;
        RECT 244.950 279.600 247.050 280.050 ;
        RECT 250.950 279.600 253.050 280.050 ;
        RECT 220.950 278.400 253.050 279.600 ;
        RECT 368.400 279.600 369.600 281.400 ;
        RECT 370.950 281.400 379.050 282.600 ;
        RECT 370.950 280.950 373.050 281.400 ;
        RECT 376.950 280.950 379.050 281.400 ;
        RECT 460.950 282.600 463.050 283.050 ;
        RECT 487.950 282.600 490.050 283.050 ;
        RECT 460.950 281.400 490.050 282.600 ;
        RECT 460.950 280.950 463.050 281.400 ;
        RECT 487.950 280.950 490.050 281.400 ;
        RECT 490.950 282.600 493.050 283.050 ;
        RECT 538.950 282.600 541.050 283.050 ;
        RECT 490.950 281.400 541.050 282.600 ;
        RECT 490.950 280.950 493.050 281.400 ;
        RECT 538.950 280.950 541.050 281.400 ;
        RECT 541.950 282.600 544.050 283.050 ;
        RECT 643.950 282.600 646.050 283.050 ;
        RECT 541.950 281.400 646.050 282.600 ;
        RECT 541.950 280.950 544.050 281.400 ;
        RECT 643.950 280.950 646.050 281.400 ;
        RECT 655.950 282.600 658.050 283.050 ;
        RECT 736.950 282.600 739.050 283.050 ;
        RECT 655.950 281.400 739.050 282.600 ;
        RECT 655.950 280.950 658.050 281.400 ;
        RECT 736.950 280.950 739.050 281.400 ;
        RECT 373.950 279.600 376.050 280.050 ;
        RECT 368.400 278.400 376.050 279.600 ;
        RECT 220.950 277.950 223.050 278.400 ;
        RECT 244.950 277.950 247.050 278.400 ;
        RECT 250.950 277.950 253.050 278.400 ;
        RECT 373.950 277.950 376.050 278.400 ;
        RECT 421.950 279.600 424.050 280.050 ;
        RECT 454.950 279.600 457.050 280.050 ;
        RECT 421.950 278.400 457.050 279.600 ;
        RECT 421.950 277.950 424.050 278.400 ;
        RECT 454.950 277.950 457.050 278.400 ;
        RECT 466.950 279.600 469.050 280.050 ;
        RECT 499.950 279.600 502.050 280.050 ;
        RECT 580.950 279.600 583.050 280.050 ;
        RECT 601.950 279.600 604.050 280.050 ;
        RECT 466.950 278.400 502.050 279.600 ;
        RECT 466.950 277.950 469.050 278.400 ;
        RECT 499.950 277.950 502.050 278.400 ;
        RECT 509.400 278.400 604.050 279.600 ;
        RECT 25.950 274.950 28.050 277.050 ;
        RECT 43.950 276.600 46.050 277.050 ;
        RECT 49.950 276.600 52.050 277.050 ;
        RECT 43.950 275.400 52.050 276.600 ;
        RECT 43.950 274.950 46.050 275.400 ;
        RECT 49.950 274.950 52.050 275.400 ;
        RECT 64.950 276.600 67.050 277.050 ;
        RECT 73.950 276.600 76.050 277.050 ;
        RECT 64.950 275.400 76.050 276.600 ;
        RECT 64.950 274.950 67.050 275.400 ;
        RECT 73.950 274.950 76.050 275.400 ;
        RECT 91.950 276.600 94.050 277.050 ;
        RECT 103.950 276.600 106.050 277.050 ;
        RECT 151.950 276.600 154.050 277.050 ;
        RECT 91.950 275.400 106.050 276.600 ;
        RECT 91.950 274.950 94.050 275.400 ;
        RECT 103.950 274.950 106.050 275.400 ;
        RECT 107.400 275.400 154.050 276.600 ;
        RECT 22.950 268.950 25.050 271.050 ;
        RECT 7.950 265.950 10.050 268.050 ;
        RECT 19.950 265.950 22.050 268.050 ;
        RECT 22.950 267.600 25.050 268.050 ;
        RECT 26.400 267.600 27.600 274.950 ;
        RECT 55.950 273.600 58.050 274.050 ;
        RECT 32.400 272.400 58.050 273.600 ;
        RECT 32.400 271.050 33.600 272.400 ;
        RECT 55.950 271.950 58.050 272.400 ;
        RECT 85.950 273.600 88.050 274.050 ;
        RECT 97.950 273.600 100.050 274.050 ;
        RECT 107.400 273.600 108.600 275.400 ;
        RECT 151.950 274.950 154.050 275.400 ;
        RECT 208.950 274.950 211.050 277.050 ;
        RECT 217.950 276.600 220.050 277.050 ;
        RECT 238.950 276.600 241.050 277.050 ;
        RECT 217.950 275.400 241.050 276.600 ;
        RECT 217.950 274.950 220.050 275.400 ;
        RECT 238.950 274.950 241.050 275.400 ;
        RECT 346.950 276.600 349.050 277.050 ;
        RECT 403.950 276.600 406.050 277.050 ;
        RECT 346.950 275.400 406.050 276.600 ;
        RECT 346.950 274.950 349.050 275.400 ;
        RECT 403.950 274.950 406.050 275.400 ;
        RECT 412.950 276.600 415.050 277.050 ;
        RECT 442.950 276.600 445.050 277.050 ;
        RECT 412.950 275.400 445.050 276.600 ;
        RECT 412.950 274.950 415.050 275.400 ;
        RECT 442.950 274.950 445.050 275.400 ;
        RECT 457.950 276.600 460.050 277.050 ;
        RECT 466.950 276.600 469.050 277.050 ;
        RECT 457.950 275.400 469.050 276.600 ;
        RECT 457.950 274.950 460.050 275.400 ;
        RECT 466.950 274.950 469.050 275.400 ;
        RECT 478.950 276.600 481.050 277.050 ;
        RECT 481.950 276.600 484.050 277.050 ;
        RECT 493.950 276.600 496.050 277.050 ;
        RECT 509.400 276.600 510.600 278.400 ;
        RECT 580.950 277.950 583.050 278.400 ;
        RECT 601.950 277.950 604.050 278.400 ;
        RECT 628.950 279.600 631.050 280.050 ;
        RECT 652.950 279.600 655.050 280.050 ;
        RECT 628.950 278.400 655.050 279.600 ;
        RECT 628.950 277.950 631.050 278.400 ;
        RECT 652.950 277.950 655.050 278.400 ;
        RECT 688.950 279.600 691.050 280.050 ;
        RECT 694.950 279.600 697.050 280.050 ;
        RECT 748.950 279.600 751.050 280.050 ;
        RECT 688.950 278.400 747.600 279.600 ;
        RECT 688.950 277.950 691.050 278.400 ;
        RECT 694.950 277.950 697.050 278.400 ;
        RECT 544.950 276.600 547.050 277.050 ;
        RECT 478.950 275.400 510.600 276.600 ;
        RECT 518.400 275.400 547.050 276.600 ;
        RECT 478.950 274.950 481.050 275.400 ;
        RECT 481.950 274.950 484.050 275.400 ;
        RECT 493.950 274.950 496.050 275.400 ;
        RECT 85.950 272.400 108.600 273.600 ;
        RECT 118.950 273.600 121.050 274.050 ;
        RECT 136.950 273.600 139.050 274.050 ;
        RECT 175.950 273.600 178.050 274.050 ;
        RECT 193.950 273.600 196.050 274.050 ;
        RECT 205.950 273.600 208.050 274.050 ;
        RECT 118.950 272.400 139.050 273.600 ;
        RECT 85.950 271.950 88.050 272.400 ;
        RECT 97.950 271.950 100.050 272.400 ;
        RECT 118.950 271.950 121.050 272.400 ;
        RECT 136.950 271.950 139.050 272.400 ;
        RECT 140.400 272.400 165.600 273.600 ;
        RECT 31.950 268.950 34.050 271.050 ;
        RECT 37.950 270.600 40.050 271.050 ;
        RECT 35.400 269.400 40.050 270.600 ;
        RECT 22.950 266.400 27.600 267.600 ;
        RECT 31.950 267.600 34.050 268.050 ;
        RECT 35.400 267.600 36.600 269.400 ;
        RECT 37.950 268.950 40.050 269.400 ;
        RECT 52.950 270.600 55.050 271.050 ;
        RECT 64.950 270.600 67.050 271.050 ;
        RECT 52.950 269.400 67.050 270.600 ;
        RECT 52.950 268.950 55.050 269.400 ;
        RECT 64.950 268.950 67.050 269.400 ;
        RECT 79.950 270.600 82.050 271.050 ;
        RECT 88.950 270.600 91.050 271.050 ;
        RECT 79.950 269.400 91.050 270.600 ;
        RECT 79.950 268.950 82.050 269.400 ;
        RECT 88.950 268.950 91.050 269.400 ;
        RECT 106.950 270.600 109.050 271.050 ;
        RECT 121.950 270.600 124.050 271.050 ;
        RECT 127.950 270.600 130.050 271.050 ;
        RECT 140.400 270.600 141.600 272.400 ;
        RECT 106.950 269.400 124.050 270.600 ;
        RECT 106.950 268.950 109.050 269.400 ;
        RECT 121.950 268.950 124.050 269.400 ;
        RECT 125.400 269.400 130.050 270.600 ;
        RECT 31.950 266.400 36.600 267.600 ;
        RECT 37.950 267.600 40.050 268.050 ;
        RECT 58.950 267.600 61.050 268.050 ;
        RECT 37.950 266.400 61.050 267.600 ;
        RECT 22.950 265.950 25.050 266.400 ;
        RECT 31.950 265.950 34.050 266.400 ;
        RECT 37.950 265.950 40.050 266.400 ;
        RECT 58.950 265.950 61.050 266.400 ;
        RECT 109.950 267.600 112.050 268.050 ;
        RECT 118.950 267.600 121.050 268.050 ;
        RECT 109.950 266.400 121.050 267.600 ;
        RECT 109.950 265.950 112.050 266.400 ;
        RECT 118.950 265.950 121.050 266.400 ;
        RECT 121.950 267.600 124.050 268.050 ;
        RECT 125.400 267.600 126.600 269.400 ;
        RECT 127.950 268.950 130.050 269.400 ;
        RECT 134.400 269.400 141.600 270.600 ;
        RECT 134.400 268.050 135.600 269.400 ;
        RECT 142.950 268.950 145.050 271.050 ;
        RECT 157.950 268.950 160.050 271.050 ;
        RECT 160.950 268.950 163.050 271.050 ;
        RECT 164.400 270.600 165.600 272.400 ;
        RECT 175.950 272.400 208.050 273.600 ;
        RECT 175.950 271.950 178.050 272.400 ;
        RECT 193.950 271.950 196.050 272.400 ;
        RECT 205.950 271.950 208.050 272.400 ;
        RECT 209.400 271.050 210.600 274.950 ;
        RECT 214.950 273.600 217.050 274.050 ;
        RECT 220.950 273.600 223.050 274.050 ;
        RECT 214.950 272.400 223.050 273.600 ;
        RECT 214.950 271.950 217.050 272.400 ;
        RECT 220.950 271.950 223.050 272.400 ;
        RECT 232.950 273.600 235.050 274.050 ;
        RECT 250.950 273.600 253.050 274.050 ;
        RECT 232.950 272.400 253.050 273.600 ;
        RECT 232.950 271.950 235.050 272.400 ;
        RECT 250.950 271.950 253.050 272.400 ;
        RECT 268.950 273.600 271.050 274.050 ;
        RECT 331.950 273.600 334.050 274.050 ;
        RECT 268.950 272.400 334.050 273.600 ;
        RECT 268.950 271.950 271.050 272.400 ;
        RECT 331.950 271.950 334.050 272.400 ;
        RECT 337.950 273.600 340.050 274.050 ;
        RECT 346.950 273.600 349.050 274.050 ;
        RECT 337.950 272.400 349.050 273.600 ;
        RECT 337.950 271.950 340.050 272.400 ;
        RECT 346.950 271.950 349.050 272.400 ;
        RECT 358.950 273.600 361.050 274.050 ;
        RECT 430.950 273.600 433.050 274.050 ;
        RECT 436.950 273.600 439.050 274.050 ;
        RECT 358.950 272.400 439.050 273.600 ;
        RECT 358.950 271.950 361.050 272.400 ;
        RECT 430.950 271.950 433.050 272.400 ;
        RECT 436.950 271.950 439.050 272.400 ;
        RECT 442.950 273.600 445.050 274.050 ;
        RECT 451.950 273.600 454.050 274.050 ;
        RECT 442.950 272.400 454.050 273.600 ;
        RECT 442.950 271.950 445.050 272.400 ;
        RECT 451.950 271.950 454.050 272.400 ;
        RECT 472.950 271.950 475.050 274.050 ;
        RECT 499.950 273.600 502.050 274.050 ;
        RECT 508.950 273.600 511.050 274.050 ;
        RECT 518.400 273.600 519.600 275.400 ;
        RECT 544.950 274.950 547.050 275.400 ;
        RECT 583.950 276.600 586.050 277.050 ;
        RECT 595.950 276.600 598.050 277.050 ;
        RECT 583.950 275.400 598.050 276.600 ;
        RECT 583.950 274.950 586.050 275.400 ;
        RECT 595.950 274.950 598.050 275.400 ;
        RECT 601.950 276.600 604.050 277.050 ;
        RECT 631.950 276.600 634.050 277.050 ;
        RECT 667.950 276.600 670.050 277.050 ;
        RECT 700.950 276.600 703.050 277.050 ;
        RECT 601.950 275.400 634.050 276.600 ;
        RECT 601.950 274.950 604.050 275.400 ;
        RECT 631.950 274.950 634.050 275.400 ;
        RECT 644.400 275.400 666.600 276.600 ;
        RECT 499.950 272.400 511.050 273.600 ;
        RECT 499.950 271.950 502.050 272.400 ;
        RECT 508.950 271.950 511.050 272.400 ;
        RECT 515.400 272.400 519.600 273.600 ;
        RECT 190.950 270.600 193.050 271.050 ;
        RECT 196.950 270.600 199.050 271.050 ;
        RECT 164.400 269.400 177.600 270.600 ;
        RECT 121.950 266.400 126.600 267.600 ;
        RECT 121.950 265.950 124.050 266.400 ;
        RECT 133.950 265.950 136.050 268.050 ;
        RECT 4.950 264.600 7.050 265.050 ;
        RECT 10.950 264.600 13.050 265.050 ;
        RECT 4.950 263.400 13.050 264.600 ;
        RECT 4.950 262.950 7.050 263.400 ;
        RECT 10.950 262.950 13.050 263.400 ;
        RECT 13.950 264.600 16.050 265.050 ;
        RECT 28.950 264.600 31.050 265.050 ;
        RECT 76.950 264.600 79.050 265.050 ;
        RECT 13.950 263.400 79.050 264.600 ;
        RECT 13.950 262.950 16.050 263.400 ;
        RECT 28.950 262.950 31.050 263.400 ;
        RECT 76.950 262.950 79.050 263.400 ;
        RECT 100.950 264.600 103.050 265.050 ;
        RECT 124.950 264.600 127.050 265.050 ;
        RECT 100.950 263.400 127.050 264.600 ;
        RECT 100.950 262.950 103.050 263.400 ;
        RECT 124.950 262.950 127.050 263.400 ;
        RECT 4.950 261.600 7.050 262.050 ;
        RECT 34.950 261.600 37.050 262.050 ;
        RECT 43.950 261.600 46.050 262.050 ;
        RECT 4.950 260.400 46.050 261.600 ;
        RECT 4.950 259.950 7.050 260.400 ;
        RECT 34.950 259.950 37.050 260.400 ;
        RECT 43.950 259.950 46.050 260.400 ;
        RECT 46.950 261.600 49.050 262.050 ;
        RECT 49.950 261.600 52.050 262.050 ;
        RECT 61.950 261.600 64.050 262.050 ;
        RECT 46.950 260.400 64.050 261.600 ;
        RECT 46.950 259.950 49.050 260.400 ;
        RECT 49.950 259.950 52.050 260.400 ;
        RECT 61.950 259.950 64.050 260.400 ;
        RECT 82.950 261.600 85.050 262.050 ;
        RECT 103.950 261.600 106.050 262.050 ;
        RECT 112.950 261.600 115.050 262.050 ;
        RECT 82.950 260.400 115.050 261.600 ;
        RECT 82.950 259.950 85.050 260.400 ;
        RECT 103.950 259.950 106.050 260.400 ;
        RECT 112.950 259.950 115.050 260.400 ;
        RECT 115.950 261.600 118.050 262.050 ;
        RECT 133.950 261.600 136.050 262.050 ;
        RECT 115.950 260.400 136.050 261.600 ;
        RECT 143.400 261.600 144.600 268.950 ;
        RECT 145.950 264.600 148.050 265.050 ;
        RECT 158.400 264.600 159.600 268.950 ;
        RECT 161.400 267.600 162.600 268.950 ;
        RECT 166.950 267.600 169.050 268.050 ;
        RECT 176.400 267.600 177.600 269.400 ;
        RECT 190.950 269.400 199.050 270.600 ;
        RECT 190.950 268.950 193.050 269.400 ;
        RECT 196.950 268.950 199.050 269.400 ;
        RECT 208.950 268.950 211.050 271.050 ;
        RECT 235.950 270.600 238.050 271.050 ;
        RECT 262.950 270.600 265.050 271.050 ;
        RECT 235.950 269.400 265.050 270.600 ;
        RECT 235.950 268.950 238.050 269.400 ;
        RECT 262.950 268.950 265.050 269.400 ;
        RECT 298.950 270.600 301.050 271.050 ;
        RECT 304.950 270.600 307.050 271.050 ;
        RECT 298.950 269.400 307.050 270.600 ;
        RECT 298.950 268.950 301.050 269.400 ;
        RECT 304.950 268.950 307.050 269.400 ;
        RECT 313.950 268.950 316.050 271.050 ;
        RECT 325.950 270.600 328.050 271.050 ;
        RECT 334.950 270.600 337.050 271.050 ;
        RECT 325.950 269.400 337.050 270.600 ;
        RECT 325.950 268.950 328.050 269.400 ;
        RECT 334.950 268.950 337.050 269.400 ;
        RECT 337.950 270.600 340.050 271.050 ;
        RECT 364.950 270.600 367.050 271.050 ;
        RECT 337.950 269.400 367.050 270.600 ;
        RECT 337.950 268.950 340.050 269.400 ;
        RECT 364.950 268.950 367.050 269.400 ;
        RECT 370.950 270.600 373.050 271.050 ;
        RECT 376.950 270.600 379.050 271.050 ;
        RECT 412.950 270.600 415.050 271.050 ;
        RECT 463.950 270.600 466.050 271.050 ;
        RECT 370.950 269.400 379.050 270.600 ;
        RECT 370.950 268.950 373.050 269.400 ;
        RECT 376.950 268.950 379.050 269.400 ;
        RECT 401.400 269.400 415.050 270.600 ;
        RECT 226.950 267.600 229.050 268.050 ;
        RECT 161.400 266.400 174.600 267.600 ;
        RECT 176.400 266.400 229.050 267.600 ;
        RECT 166.950 265.950 169.050 266.400 ;
        RECT 169.950 264.600 172.050 265.050 ;
        RECT 145.950 263.400 172.050 264.600 ;
        RECT 173.400 264.600 174.600 266.400 ;
        RECT 226.950 265.950 229.050 266.400 ;
        RECT 229.950 267.600 232.050 268.050 ;
        RECT 277.950 267.600 280.050 268.050 ;
        RECT 229.950 266.400 280.050 267.600 ;
        RECT 314.400 267.600 315.600 268.950 ;
        RECT 322.950 267.600 325.050 268.050 ;
        RECT 314.400 266.400 325.050 267.600 ;
        RECT 229.950 265.950 232.050 266.400 ;
        RECT 245.400 265.050 246.600 266.400 ;
        RECT 277.950 265.950 280.050 266.400 ;
        RECT 322.950 265.950 325.050 266.400 ;
        RECT 334.950 267.600 337.050 268.050 ;
        RECT 361.950 267.600 364.050 268.050 ;
        RECT 334.950 266.400 364.050 267.600 ;
        RECT 365.400 267.600 366.600 268.950 ;
        RECT 365.400 266.400 372.600 267.600 ;
        RECT 334.950 265.950 337.050 266.400 ;
        RECT 361.950 265.950 364.050 266.400 ;
        RECT 181.950 264.600 184.050 265.050 ;
        RECT 173.400 263.400 184.050 264.600 ;
        RECT 145.950 262.950 148.050 263.400 ;
        RECT 169.950 262.950 172.050 263.400 ;
        RECT 181.950 262.950 184.050 263.400 ;
        RECT 202.950 264.600 205.050 265.050 ;
        RECT 214.950 264.600 217.050 265.050 ;
        RECT 202.950 263.400 217.050 264.600 ;
        RECT 202.950 262.950 205.050 263.400 ;
        RECT 214.950 262.950 217.050 263.400 ;
        RECT 244.950 262.950 247.050 265.050 ;
        RECT 265.950 264.600 268.050 265.050 ;
        RECT 280.950 264.600 283.050 265.050 ;
        RECT 265.950 263.400 283.050 264.600 ;
        RECT 265.950 262.950 268.050 263.400 ;
        RECT 280.950 262.950 283.050 263.400 ;
        RECT 283.950 264.600 286.050 265.050 ;
        RECT 286.950 264.600 289.050 265.050 ;
        RECT 316.950 264.600 319.050 265.050 ;
        RECT 283.950 263.400 319.050 264.600 ;
        RECT 283.950 262.950 286.050 263.400 ;
        RECT 286.950 262.950 289.050 263.400 ;
        RECT 316.950 262.950 319.050 263.400 ;
        RECT 328.950 264.600 331.050 265.050 ;
        RECT 367.950 264.600 370.050 265.050 ;
        RECT 328.950 263.400 370.050 264.600 ;
        RECT 371.400 264.600 372.600 266.400 ;
        RECT 385.950 264.600 388.050 265.050 ;
        RECT 371.400 263.400 388.050 264.600 ;
        RECT 328.950 262.950 331.050 263.400 ;
        RECT 367.950 262.950 370.050 263.400 ;
        RECT 385.950 262.950 388.050 263.400 ;
        RECT 391.950 264.600 394.050 265.050 ;
        RECT 401.400 264.600 402.600 269.400 ;
        RECT 412.950 268.950 415.050 269.400 ;
        RECT 449.400 269.400 466.050 270.600 ;
        RECT 473.400 270.600 474.600 271.950 ;
        RECT 487.950 270.600 490.050 271.050 ;
        RECT 473.400 269.400 490.050 270.600 ;
        RECT 449.400 268.050 450.600 269.400 ;
        RECT 463.950 268.950 466.050 269.400 ;
        RECT 487.950 268.950 490.050 269.400 ;
        RECT 505.950 270.600 508.050 271.050 ;
        RECT 515.400 270.600 516.600 272.400 ;
        RECT 520.950 271.950 523.050 274.050 ;
        RECT 565.950 273.600 568.050 274.050 ;
        RECT 589.950 273.600 592.050 274.050 ;
        RECT 607.950 273.600 610.050 274.050 ;
        RECT 625.950 273.600 628.050 274.050 ;
        RECT 565.950 272.400 570.600 273.600 ;
        RECT 565.950 271.950 568.050 272.400 ;
        RECT 505.950 269.400 516.600 270.600 ;
        RECT 505.950 268.950 508.050 269.400 ;
        RECT 517.950 268.950 520.050 271.050 ;
        RECT 415.950 267.600 418.050 268.050 ;
        RECT 427.950 267.600 430.050 268.050 ;
        RECT 415.950 266.400 430.050 267.600 ;
        RECT 415.950 265.950 418.050 266.400 ;
        RECT 427.950 265.950 430.050 266.400 ;
        RECT 448.950 265.950 451.050 268.050 ;
        RECT 451.950 267.600 454.050 268.050 ;
        RECT 484.950 267.600 487.050 268.050 ;
        RECT 499.950 267.600 502.050 268.050 ;
        RECT 451.950 266.400 502.050 267.600 ;
        RECT 451.950 265.950 454.050 266.400 ;
        RECT 484.950 265.950 487.050 266.400 ;
        RECT 499.950 265.950 502.050 266.400 ;
        RECT 505.950 267.600 508.050 268.050 ;
        RECT 518.400 267.600 519.600 268.950 ;
        RECT 505.950 266.400 519.600 267.600 ;
        RECT 521.400 267.600 522.600 271.950 ;
        RECT 523.950 270.600 526.050 271.050 ;
        RECT 532.950 270.600 535.050 271.050 ;
        RECT 523.950 269.400 535.050 270.600 ;
        RECT 523.950 268.950 526.050 269.400 ;
        RECT 532.950 268.950 535.050 269.400 ;
        RECT 544.950 270.600 547.050 271.050 ;
        RECT 559.950 270.600 562.050 271.050 ;
        RECT 565.950 270.600 568.050 271.050 ;
        RECT 544.950 269.400 555.600 270.600 ;
        RECT 544.950 268.950 547.050 269.400 ;
        RECT 554.400 268.050 555.600 269.400 ;
        RECT 559.950 269.400 568.050 270.600 ;
        RECT 559.950 268.950 562.050 269.400 ;
        RECT 565.950 268.950 568.050 269.400 ;
        RECT 529.950 267.600 532.050 268.050 ;
        RECT 521.400 266.400 532.050 267.600 ;
        RECT 505.950 265.950 508.050 266.400 ;
        RECT 529.950 265.950 532.050 266.400 ;
        RECT 532.950 267.600 535.050 268.050 ;
        RECT 541.950 267.600 544.050 268.050 ;
        RECT 532.950 266.400 544.050 267.600 ;
        RECT 532.950 265.950 535.050 266.400 ;
        RECT 541.950 265.950 544.050 266.400 ;
        RECT 553.950 265.950 556.050 268.050 ;
        RECT 569.400 265.050 570.600 272.400 ;
        RECT 589.950 272.400 594.600 273.600 ;
        RECT 589.950 271.950 592.050 272.400 ;
        RECT 593.400 268.050 594.600 272.400 ;
        RECT 607.950 272.400 628.050 273.600 ;
        RECT 607.950 271.950 610.050 272.400 ;
        RECT 625.950 271.950 628.050 272.400 ;
        RECT 595.950 268.950 598.050 271.050 ;
        RECT 619.950 270.600 622.050 271.050 ;
        RECT 644.400 270.600 645.600 275.400 ;
        RECT 649.950 273.600 652.050 274.050 ;
        RECT 619.950 269.400 627.600 270.600 ;
        RECT 619.950 268.950 622.050 269.400 ;
        RECT 592.950 265.950 595.050 268.050 ;
        RECT 391.950 263.400 402.600 264.600 ;
        RECT 448.950 264.600 451.050 265.050 ;
        RECT 454.950 264.600 457.050 265.050 ;
        RECT 448.950 263.400 457.050 264.600 ;
        RECT 391.950 262.950 394.050 263.400 ;
        RECT 448.950 262.950 451.050 263.400 ;
        RECT 454.950 262.950 457.050 263.400 ;
        RECT 460.950 264.600 463.050 265.050 ;
        RECT 484.950 264.600 487.050 265.050 ;
        RECT 487.950 264.600 490.050 265.050 ;
        RECT 460.950 263.400 490.050 264.600 ;
        RECT 460.950 262.950 463.050 263.400 ;
        RECT 484.950 262.950 487.050 263.400 ;
        RECT 487.950 262.950 490.050 263.400 ;
        RECT 499.950 264.600 502.050 265.050 ;
        RECT 520.950 264.600 523.050 265.050 ;
        RECT 556.950 264.600 559.050 265.050 ;
        RECT 499.950 263.400 519.600 264.600 ;
        RECT 499.950 262.950 502.050 263.400 ;
        RECT 145.950 261.600 148.050 262.050 ;
        RECT 143.400 260.400 148.050 261.600 ;
        RECT 115.950 259.950 118.050 260.400 ;
        RECT 133.950 259.950 136.050 260.400 ;
        RECT 145.950 259.950 148.050 260.400 ;
        RECT 160.950 261.600 163.050 262.050 ;
        RECT 163.950 261.600 166.050 262.050 ;
        RECT 172.950 261.600 175.050 262.050 ;
        RECT 184.950 261.600 187.050 262.050 ;
        RECT 160.950 260.400 187.050 261.600 ;
        RECT 160.950 259.950 163.050 260.400 ;
        RECT 163.950 259.950 166.050 260.400 ;
        RECT 172.950 259.950 175.050 260.400 ;
        RECT 184.950 259.950 187.050 260.400 ;
        RECT 352.950 261.600 355.050 262.050 ;
        RECT 388.950 261.600 391.050 262.050 ;
        RECT 424.950 261.600 427.050 262.050 ;
        RECT 352.950 260.400 427.050 261.600 ;
        RECT 352.950 259.950 355.050 260.400 ;
        RECT 388.950 259.950 391.050 260.400 ;
        RECT 424.950 259.950 427.050 260.400 ;
        RECT 439.950 261.600 442.050 262.050 ;
        RECT 475.950 261.600 478.050 262.050 ;
        RECT 439.950 260.400 478.050 261.600 ;
        RECT 439.950 259.950 442.050 260.400 ;
        RECT 475.950 259.950 478.050 260.400 ;
        RECT 484.950 261.600 487.050 262.050 ;
        RECT 514.950 261.600 517.050 262.050 ;
        RECT 484.950 260.400 517.050 261.600 ;
        RECT 518.400 261.600 519.600 263.400 ;
        RECT 520.950 263.400 559.050 264.600 ;
        RECT 520.950 262.950 523.050 263.400 ;
        RECT 556.950 262.950 559.050 263.400 ;
        RECT 568.950 262.950 571.050 265.050 ;
        RECT 596.400 264.600 597.600 268.950 ;
        RECT 626.400 268.050 627.600 269.400 ;
        RECT 638.400 269.400 645.600 270.600 ;
        RECT 647.400 272.400 652.050 273.600 ;
        RECT 598.950 267.600 601.050 268.050 ;
        RECT 598.950 266.400 618.600 267.600 ;
        RECT 598.950 265.950 601.050 266.400 ;
        RECT 598.950 264.600 601.050 265.050 ;
        RECT 596.400 263.400 601.050 264.600 ;
        RECT 598.950 262.950 601.050 263.400 ;
        RECT 601.950 264.600 604.050 265.050 ;
        RECT 613.950 264.600 616.050 265.050 ;
        RECT 601.950 263.400 616.050 264.600 ;
        RECT 601.950 262.950 604.050 263.400 ;
        RECT 613.950 262.950 616.050 263.400 ;
        RECT 526.950 261.600 529.050 262.050 ;
        RECT 518.400 260.400 529.050 261.600 ;
        RECT 484.950 259.950 487.050 260.400 ;
        RECT 514.950 259.950 517.050 260.400 ;
        RECT 526.950 259.950 529.050 260.400 ;
        RECT 532.950 261.600 535.050 262.050 ;
        RECT 538.950 261.600 541.050 262.050 ;
        RECT 532.950 260.400 541.050 261.600 ;
        RECT 532.950 259.950 535.050 260.400 ;
        RECT 538.950 259.950 541.050 260.400 ;
        RECT 571.950 261.600 574.050 262.050 ;
        RECT 574.950 261.600 577.050 262.050 ;
        RECT 604.950 261.600 607.050 262.050 ;
        RECT 571.950 260.400 607.050 261.600 ;
        RECT 617.400 261.600 618.600 266.400 ;
        RECT 625.950 265.950 628.050 268.050 ;
        RECT 619.950 264.600 622.050 265.050 ;
        RECT 638.400 264.600 639.600 269.400 ;
        RECT 643.950 267.600 646.050 268.050 ;
        RECT 647.400 267.600 648.600 272.400 ;
        RECT 649.950 271.950 652.050 272.400 ;
        RECT 652.950 271.950 655.050 274.050 ;
        RECT 665.400 273.600 666.600 275.400 ;
        RECT 667.950 275.400 703.050 276.600 ;
        RECT 667.950 274.950 670.050 275.400 ;
        RECT 700.950 274.950 703.050 275.400 ;
        RECT 715.950 276.600 718.050 277.050 ;
        RECT 733.950 276.600 736.050 277.050 ;
        RECT 715.950 275.400 736.050 276.600 ;
        RECT 715.950 274.950 718.050 275.400 ;
        RECT 733.950 274.950 736.050 275.400 ;
        RECT 736.950 276.600 739.050 277.050 ;
        RECT 746.400 276.600 747.600 278.400 ;
        RECT 748.950 278.400 774.600 279.600 ;
        RECT 748.950 277.950 751.050 278.400 ;
        RECT 763.950 276.600 766.050 277.050 ;
        RECT 736.950 275.400 741.600 276.600 ;
        RECT 746.400 275.400 766.050 276.600 ;
        RECT 736.950 274.950 739.050 275.400 ;
        RECT 740.400 274.050 741.600 275.400 ;
        RECT 763.950 274.950 766.050 275.400 ;
        RECT 682.950 273.600 685.050 274.050 ;
        RECT 665.400 272.400 685.050 273.600 ;
        RECT 682.950 271.950 685.050 272.400 ;
        RECT 691.950 273.600 694.050 274.050 ;
        RECT 706.950 273.600 709.050 274.050 ;
        RECT 691.950 272.400 709.050 273.600 ;
        RECT 691.950 271.950 694.050 272.400 ;
        RECT 706.950 271.950 709.050 272.400 ;
        RECT 739.950 271.950 742.050 274.050 ;
        RECT 653.400 270.600 654.600 271.950 ;
        RECT 650.400 269.400 654.600 270.600 ;
        RECT 650.400 268.050 651.600 269.400 ;
        RECT 655.950 268.950 658.050 271.050 ;
        RECT 661.950 268.950 664.050 271.050 ;
        RECT 670.950 270.600 673.050 271.050 ;
        RECT 682.950 270.600 685.050 271.050 ;
        RECT 703.950 270.600 706.050 271.050 ;
        RECT 718.950 270.600 721.050 271.050 ;
        RECT 670.950 269.400 675.600 270.600 ;
        RECT 670.950 268.950 673.050 269.400 ;
        RECT 643.950 266.400 648.600 267.600 ;
        RECT 643.950 265.950 646.050 266.400 ;
        RECT 649.950 265.950 652.050 268.050 ;
        RECT 619.950 263.400 639.600 264.600 ;
        RECT 646.950 264.600 649.050 265.050 ;
        RECT 656.400 264.600 657.600 268.950 ;
        RECT 662.400 267.600 663.600 268.950 ;
        RECT 662.400 266.400 672.600 267.600 ;
        RECT 671.400 265.050 672.600 266.400 ;
        RECT 667.950 264.600 670.050 265.050 ;
        RECT 646.950 263.400 670.050 264.600 ;
        RECT 619.950 262.950 622.050 263.400 ;
        RECT 646.950 262.950 649.050 263.400 ;
        RECT 667.950 262.950 670.050 263.400 ;
        RECT 670.950 262.950 673.050 265.050 ;
        RECT 674.400 264.600 675.600 269.400 ;
        RECT 682.950 269.400 721.050 270.600 ;
        RECT 682.950 268.950 685.050 269.400 ;
        RECT 703.950 268.950 706.050 269.400 ;
        RECT 718.950 268.950 721.050 269.400 ;
        RECT 736.950 270.600 739.050 271.050 ;
        RECT 751.950 270.600 754.050 271.050 ;
        RECT 736.950 269.400 754.050 270.600 ;
        RECT 736.950 268.950 739.050 269.400 ;
        RECT 751.950 268.950 754.050 269.400 ;
        RECT 700.950 267.600 703.050 268.050 ;
        RECT 715.950 267.600 718.050 268.050 ;
        RECT 700.950 266.400 718.050 267.600 ;
        RECT 700.950 265.950 703.050 266.400 ;
        RECT 715.950 265.950 718.050 266.400 ;
        RECT 724.950 267.600 727.050 268.050 ;
        RECT 739.950 267.600 742.050 268.050 ;
        RECT 748.950 267.600 751.050 268.050 ;
        RECT 724.950 266.400 742.050 267.600 ;
        RECT 724.950 265.950 727.050 266.400 ;
        RECT 739.950 265.950 742.050 266.400 ;
        RECT 743.400 266.400 751.050 267.600 ;
        RECT 685.950 264.600 688.050 265.050 ;
        RECT 709.950 264.600 712.050 265.050 ;
        RECT 743.400 264.600 744.600 266.400 ;
        RECT 748.950 265.950 751.050 266.400 ;
        RECT 754.950 267.600 757.050 268.050 ;
        RECT 769.950 267.600 772.050 268.050 ;
        RECT 754.950 266.400 772.050 267.600 ;
        RECT 754.950 265.950 757.050 266.400 ;
        RECT 769.950 265.950 772.050 266.400 ;
        RECT 674.400 263.400 744.600 264.600 ;
        RECT 745.950 264.600 748.050 265.050 ;
        RECT 763.950 264.600 766.050 265.050 ;
        RECT 773.400 264.600 774.600 278.400 ;
        RECT 745.950 263.400 766.050 264.600 ;
        RECT 685.950 262.950 688.050 263.400 ;
        RECT 709.950 262.950 712.050 263.400 ;
        RECT 745.950 262.950 748.050 263.400 ;
        RECT 763.950 262.950 766.050 263.400 ;
        RECT 767.400 263.400 774.600 264.600 ;
        RECT 619.950 261.600 622.050 262.050 ;
        RECT 617.400 260.400 622.050 261.600 ;
        RECT 571.950 259.950 574.050 260.400 ;
        RECT 574.950 259.950 577.050 260.400 ;
        RECT 604.950 259.950 607.050 260.400 ;
        RECT 619.950 259.950 622.050 260.400 ;
        RECT 622.950 261.600 625.050 262.050 ;
        RECT 628.950 261.600 631.050 262.050 ;
        RECT 640.950 261.600 643.050 262.050 ;
        RECT 622.950 260.400 643.050 261.600 ;
        RECT 622.950 259.950 625.050 260.400 ;
        RECT 628.950 259.950 631.050 260.400 ;
        RECT 640.950 259.950 643.050 260.400 ;
        RECT 661.950 261.600 664.050 262.050 ;
        RECT 685.950 261.600 688.050 262.050 ;
        RECT 661.950 260.400 688.050 261.600 ;
        RECT 661.950 259.950 664.050 260.400 ;
        RECT 685.950 259.950 688.050 260.400 ;
        RECT 688.950 261.600 691.050 262.050 ;
        RECT 700.950 261.600 703.050 262.050 ;
        RECT 688.950 260.400 703.050 261.600 ;
        RECT 688.950 259.950 691.050 260.400 ;
        RECT 700.950 259.950 703.050 260.400 ;
        RECT 730.950 261.600 733.050 262.050 ;
        RECT 751.950 261.600 754.050 262.050 ;
        RECT 730.950 260.400 754.050 261.600 ;
        RECT 730.950 259.950 733.050 260.400 ;
        RECT 751.950 259.950 754.050 260.400 ;
        RECT 763.950 261.600 766.050 262.050 ;
        RECT 767.400 261.600 768.600 263.400 ;
        RECT 763.950 260.400 768.600 261.600 ;
        RECT 763.950 259.950 766.050 260.400 ;
        RECT 88.950 258.600 91.050 259.050 ;
        RECT 145.950 258.600 148.050 259.050 ;
        RECT 88.950 257.400 148.050 258.600 ;
        RECT 88.950 256.950 91.050 257.400 ;
        RECT 145.950 256.950 148.050 257.400 ;
        RECT 166.950 258.600 169.050 259.050 ;
        RECT 175.950 258.600 178.050 259.050 ;
        RECT 223.950 258.600 226.050 259.050 ;
        RECT 166.950 257.400 178.050 258.600 ;
        RECT 166.950 256.950 169.050 257.400 ;
        RECT 175.950 256.950 178.050 257.400 ;
        RECT 179.400 257.400 226.050 258.600 ;
        RECT 76.950 255.600 79.050 256.050 ;
        RECT 100.950 255.600 103.050 256.050 ;
        RECT 139.950 255.600 142.050 256.050 ;
        RECT 76.950 254.400 142.050 255.600 ;
        RECT 76.950 253.950 79.050 254.400 ;
        RECT 100.950 253.950 103.050 254.400 ;
        RECT 139.950 253.950 142.050 254.400 ;
        RECT 175.950 255.600 178.050 256.050 ;
        RECT 179.400 255.600 180.600 257.400 ;
        RECT 223.950 256.950 226.050 257.400 ;
        RECT 226.950 258.600 229.050 259.050 ;
        RECT 277.950 258.600 280.050 259.050 ;
        RECT 226.950 257.400 280.050 258.600 ;
        RECT 226.950 256.950 229.050 257.400 ;
        RECT 277.950 256.950 280.050 257.400 ;
        RECT 340.950 258.600 343.050 259.050 ;
        RECT 355.950 258.600 358.050 259.050 ;
        RECT 400.950 258.600 403.050 259.050 ;
        RECT 340.950 257.400 403.050 258.600 ;
        RECT 340.950 256.950 343.050 257.400 ;
        RECT 355.950 256.950 358.050 257.400 ;
        RECT 400.950 256.950 403.050 257.400 ;
        RECT 421.950 258.600 424.050 259.050 ;
        RECT 436.950 258.600 439.050 259.050 ;
        RECT 421.950 257.400 439.050 258.600 ;
        RECT 421.950 256.950 424.050 257.400 ;
        RECT 436.950 256.950 439.050 257.400 ;
        RECT 454.950 258.600 457.050 259.050 ;
        RECT 466.950 258.600 469.050 259.050 ;
        RECT 454.950 257.400 469.050 258.600 ;
        RECT 454.950 256.950 457.050 257.400 ;
        RECT 466.950 256.950 469.050 257.400 ;
        RECT 487.950 258.600 490.050 259.050 ;
        RECT 496.950 258.600 499.050 259.050 ;
        RECT 487.950 257.400 499.050 258.600 ;
        RECT 487.950 256.950 490.050 257.400 ;
        RECT 496.950 256.950 499.050 257.400 ;
        RECT 586.950 258.600 589.050 259.050 ;
        RECT 616.950 258.600 619.050 259.050 ;
        RECT 586.950 257.400 619.050 258.600 ;
        RECT 586.950 256.950 589.050 257.400 ;
        RECT 616.950 256.950 619.050 257.400 ;
        RECT 628.950 258.600 631.050 259.050 ;
        RECT 643.950 258.600 646.050 259.050 ;
        RECT 628.950 257.400 646.050 258.600 ;
        RECT 628.950 256.950 631.050 257.400 ;
        RECT 643.950 256.950 646.050 257.400 ;
        RECT 670.950 258.600 673.050 259.050 ;
        RECT 709.950 258.600 712.050 259.050 ;
        RECT 670.950 257.400 712.050 258.600 ;
        RECT 670.950 256.950 673.050 257.400 ;
        RECT 709.950 256.950 712.050 257.400 ;
        RECT 760.950 258.600 763.050 259.050 ;
        RECT 769.950 258.600 772.050 259.050 ;
        RECT 760.950 257.400 772.050 258.600 ;
        RECT 760.950 256.950 763.050 257.400 ;
        RECT 769.950 256.950 772.050 257.400 ;
        RECT 175.950 254.400 180.600 255.600 ;
        RECT 187.950 255.600 190.050 256.050 ;
        RECT 241.950 255.600 244.050 256.050 ;
        RECT 187.950 254.400 244.050 255.600 ;
        RECT 175.950 253.950 178.050 254.400 ;
        RECT 187.950 253.950 190.050 254.400 ;
        RECT 241.950 253.950 244.050 254.400 ;
        RECT 268.950 255.600 271.050 256.050 ;
        RECT 289.950 255.600 292.050 256.050 ;
        RECT 268.950 254.400 292.050 255.600 ;
        RECT 268.950 253.950 271.050 254.400 ;
        RECT 289.950 253.950 292.050 254.400 ;
        RECT 301.950 255.600 304.050 256.050 ;
        RECT 340.950 255.600 343.050 256.050 ;
        RECT 301.950 254.400 343.050 255.600 ;
        RECT 301.950 253.950 304.050 254.400 ;
        RECT 340.950 253.950 343.050 254.400 ;
        RECT 343.950 255.600 346.050 256.050 ;
        RECT 409.950 255.600 412.050 256.050 ;
        RECT 343.950 254.400 412.050 255.600 ;
        RECT 343.950 253.950 346.050 254.400 ;
        RECT 409.950 253.950 412.050 254.400 ;
        RECT 436.950 255.600 439.050 256.050 ;
        RECT 583.950 255.600 586.050 256.050 ;
        RECT 436.950 254.400 586.050 255.600 ;
        RECT 436.950 253.950 439.050 254.400 ;
        RECT 583.950 253.950 586.050 254.400 ;
        RECT 589.950 255.600 592.050 256.050 ;
        RECT 616.950 255.600 619.050 256.050 ;
        RECT 589.950 254.400 619.050 255.600 ;
        RECT 589.950 253.950 592.050 254.400 ;
        RECT 616.950 253.950 619.050 254.400 ;
        RECT 619.950 255.600 622.050 256.050 ;
        RECT 652.950 255.600 655.050 256.050 ;
        RECT 697.950 255.600 700.050 256.050 ;
        RECT 619.950 254.400 700.050 255.600 ;
        RECT 619.950 253.950 622.050 254.400 ;
        RECT 652.950 253.950 655.050 254.400 ;
        RECT 697.950 253.950 700.050 254.400 ;
        RECT 718.950 255.600 721.050 256.050 ;
        RECT 724.950 255.600 727.050 256.050 ;
        RECT 730.950 255.600 733.050 256.050 ;
        RECT 718.950 254.400 733.050 255.600 ;
        RECT 718.950 253.950 721.050 254.400 ;
        RECT 724.950 253.950 727.050 254.400 ;
        RECT 730.950 253.950 733.050 254.400 ;
        RECT 64.950 252.600 67.050 253.050 ;
        RECT 115.950 252.600 118.050 253.050 ;
        RECT 181.950 252.600 184.050 253.050 ;
        RECT 190.950 252.600 193.050 253.050 ;
        RECT 64.950 251.400 118.050 252.600 ;
        RECT 64.950 250.950 67.050 251.400 ;
        RECT 115.950 250.950 118.050 251.400 ;
        RECT 128.400 251.400 193.050 252.600 ;
        RECT 61.950 249.600 64.050 250.050 ;
        RECT 70.950 249.600 73.050 250.050 ;
        RECT 128.400 249.600 129.600 251.400 ;
        RECT 181.950 250.950 184.050 251.400 ;
        RECT 190.950 250.950 193.050 251.400 ;
        RECT 394.950 252.600 397.050 253.050 ;
        RECT 400.950 252.600 403.050 253.050 ;
        RECT 394.950 251.400 403.050 252.600 ;
        RECT 394.950 250.950 397.050 251.400 ;
        RECT 400.950 250.950 403.050 251.400 ;
        RECT 430.950 252.600 433.050 253.050 ;
        RECT 451.950 252.600 454.050 253.050 ;
        RECT 430.950 251.400 454.050 252.600 ;
        RECT 430.950 250.950 433.050 251.400 ;
        RECT 451.950 250.950 454.050 251.400 ;
        RECT 466.950 252.600 469.050 253.050 ;
        RECT 472.950 252.600 475.050 253.050 ;
        RECT 508.950 252.600 511.050 253.050 ;
        RECT 466.950 251.400 511.050 252.600 ;
        RECT 466.950 250.950 469.050 251.400 ;
        RECT 472.950 250.950 475.050 251.400 ;
        RECT 508.950 250.950 511.050 251.400 ;
        RECT 529.950 252.600 532.050 253.050 ;
        RECT 538.950 252.600 541.050 253.050 ;
        RECT 529.950 251.400 541.050 252.600 ;
        RECT 529.950 250.950 532.050 251.400 ;
        RECT 538.950 250.950 541.050 251.400 ;
        RECT 547.950 252.600 550.050 253.050 ;
        RECT 595.950 252.600 598.050 253.050 ;
        RECT 607.950 252.600 610.050 253.050 ;
        RECT 547.950 251.400 610.050 252.600 ;
        RECT 547.950 250.950 550.050 251.400 ;
        RECT 595.950 250.950 598.050 251.400 ;
        RECT 607.950 250.950 610.050 251.400 ;
        RECT 658.950 252.600 661.050 253.050 ;
        RECT 670.950 252.600 673.050 253.050 ;
        RECT 658.950 251.400 673.050 252.600 ;
        RECT 658.950 250.950 661.050 251.400 ;
        RECT 670.950 250.950 673.050 251.400 ;
        RECT 673.950 252.600 676.050 253.050 ;
        RECT 706.950 252.600 709.050 253.050 ;
        RECT 673.950 251.400 709.050 252.600 ;
        RECT 673.950 250.950 676.050 251.400 ;
        RECT 706.950 250.950 709.050 251.400 ;
        RECT 709.950 252.600 712.050 253.050 ;
        RECT 736.950 252.600 739.050 253.050 ;
        RECT 709.950 251.400 739.050 252.600 ;
        RECT 709.950 250.950 712.050 251.400 ;
        RECT 736.950 250.950 739.050 251.400 ;
        RECT 61.950 248.400 129.600 249.600 ;
        RECT 130.950 249.600 133.050 250.050 ;
        RECT 136.950 249.600 139.050 250.050 ;
        RECT 151.950 249.600 154.050 250.050 ;
        RECT 178.950 249.600 181.050 250.050 ;
        RECT 247.950 249.600 250.050 250.050 ;
        RECT 259.950 249.600 262.050 250.050 ;
        RECT 130.950 248.400 262.050 249.600 ;
        RECT 61.950 247.950 64.050 248.400 ;
        RECT 70.950 247.950 73.050 248.400 ;
        RECT 130.950 247.950 133.050 248.400 ;
        RECT 136.950 247.950 139.050 248.400 ;
        RECT 151.950 247.950 154.050 248.400 ;
        RECT 178.950 247.950 181.050 248.400 ;
        RECT 247.950 247.950 250.050 248.400 ;
        RECT 259.950 247.950 262.050 248.400 ;
        RECT 274.950 249.600 277.050 250.050 ;
        RECT 280.950 249.600 283.050 250.050 ;
        RECT 274.950 248.400 283.050 249.600 ;
        RECT 274.950 247.950 277.050 248.400 ;
        RECT 280.950 247.950 283.050 248.400 ;
        RECT 286.950 249.600 289.050 250.050 ;
        RECT 310.950 249.600 313.050 250.050 ;
        RECT 286.950 248.400 313.050 249.600 ;
        RECT 286.950 247.950 289.050 248.400 ;
        RECT 310.950 247.950 313.050 248.400 ;
        RECT 322.950 249.600 325.050 250.050 ;
        RECT 328.950 249.600 331.050 250.050 ;
        RECT 364.950 249.600 367.050 250.050 ;
        RECT 322.950 248.400 367.050 249.600 ;
        RECT 322.950 247.950 325.050 248.400 ;
        RECT 328.950 247.950 331.050 248.400 ;
        RECT 364.950 247.950 367.050 248.400 ;
        RECT 409.950 249.600 412.050 250.050 ;
        RECT 415.950 249.600 418.050 250.050 ;
        RECT 409.950 248.400 418.050 249.600 ;
        RECT 409.950 247.950 412.050 248.400 ;
        RECT 415.950 247.950 418.050 248.400 ;
        RECT 427.950 249.600 430.050 250.050 ;
        RECT 445.950 249.600 448.050 250.050 ;
        RECT 481.950 249.600 484.050 250.050 ;
        RECT 427.950 248.400 444.600 249.600 ;
        RECT 427.950 247.950 430.050 248.400 ;
        RECT 40.950 246.600 43.050 247.050 ;
        RECT 52.950 246.600 55.050 247.050 ;
        RECT 106.950 246.600 109.050 247.050 ;
        RECT 40.950 245.400 109.050 246.600 ;
        RECT 40.950 244.950 43.050 245.400 ;
        RECT 52.950 244.950 55.050 245.400 ;
        RECT 106.950 244.950 109.050 245.400 ;
        RECT 109.950 246.600 112.050 247.050 ;
        RECT 115.950 246.600 118.050 247.050 ;
        RECT 109.950 245.400 118.050 246.600 ;
        RECT 109.950 244.950 112.050 245.400 ;
        RECT 115.950 244.950 118.050 245.400 ;
        RECT 124.950 246.600 127.050 247.050 ;
        RECT 157.950 246.600 160.050 247.050 ;
        RECT 124.950 245.400 160.050 246.600 ;
        RECT 124.950 244.950 127.050 245.400 ;
        RECT 157.950 244.950 160.050 245.400 ;
        RECT 172.950 246.600 175.050 247.050 ;
        RECT 214.950 246.600 217.050 247.050 ;
        RECT 172.950 245.400 217.050 246.600 ;
        RECT 172.950 244.950 175.050 245.400 ;
        RECT 214.950 244.950 217.050 245.400 ;
        RECT 220.950 246.600 223.050 247.050 ;
        RECT 298.950 246.600 301.050 247.050 ;
        RECT 304.950 246.600 307.050 247.050 ;
        RECT 220.950 245.400 307.050 246.600 ;
        RECT 220.950 244.950 223.050 245.400 ;
        RECT 298.950 244.950 301.050 245.400 ;
        RECT 304.950 244.950 307.050 245.400 ;
        RECT 319.950 246.600 322.050 247.050 ;
        RECT 331.950 246.600 334.050 247.050 ;
        RECT 319.950 245.400 334.050 246.600 ;
        RECT 319.950 244.950 322.050 245.400 ;
        RECT 331.950 244.950 334.050 245.400 ;
        RECT 340.950 246.600 343.050 247.050 ;
        RECT 355.950 246.600 358.050 247.050 ;
        RECT 340.950 245.400 358.050 246.600 ;
        RECT 340.950 244.950 343.050 245.400 ;
        RECT 355.950 244.950 358.050 245.400 ;
        RECT 358.950 246.600 361.050 247.050 ;
        RECT 376.950 246.600 379.050 247.050 ;
        RECT 358.950 245.400 379.050 246.600 ;
        RECT 358.950 244.950 361.050 245.400 ;
        RECT 376.950 244.950 379.050 245.400 ;
        RECT 391.950 246.600 394.050 247.050 ;
        RECT 439.950 246.600 442.050 247.050 ;
        RECT 391.950 245.400 442.050 246.600 ;
        RECT 443.400 246.600 444.600 248.400 ;
        RECT 445.950 248.400 484.050 249.600 ;
        RECT 445.950 247.950 448.050 248.400 ;
        RECT 481.950 247.950 484.050 248.400 ;
        RECT 490.950 249.600 493.050 250.050 ;
        RECT 496.950 249.600 499.050 250.050 ;
        RECT 490.950 248.400 499.050 249.600 ;
        RECT 490.950 247.950 493.050 248.400 ;
        RECT 496.950 247.950 499.050 248.400 ;
        RECT 559.950 249.600 562.050 250.050 ;
        RECT 613.950 249.600 616.050 250.050 ;
        RECT 559.950 248.400 616.050 249.600 ;
        RECT 559.950 247.950 562.050 248.400 ;
        RECT 613.950 247.950 616.050 248.400 ;
        RECT 619.950 249.600 622.050 250.050 ;
        RECT 625.950 249.600 628.050 250.050 ;
        RECT 619.950 248.400 628.050 249.600 ;
        RECT 619.950 247.950 622.050 248.400 ;
        RECT 625.950 247.950 628.050 248.400 ;
        RECT 637.950 249.600 640.050 250.050 ;
        RECT 688.950 249.600 691.050 250.050 ;
        RECT 637.950 248.400 691.050 249.600 ;
        RECT 637.950 247.950 640.050 248.400 ;
        RECT 688.950 247.950 691.050 248.400 ;
        RECT 691.950 249.600 694.050 250.050 ;
        RECT 718.950 249.600 721.050 250.050 ;
        RECT 691.950 248.400 721.050 249.600 ;
        RECT 691.950 247.950 694.050 248.400 ;
        RECT 718.950 247.950 721.050 248.400 ;
        RECT 721.950 249.600 724.050 250.050 ;
        RECT 766.950 249.600 769.050 250.050 ;
        RECT 721.950 248.400 769.050 249.600 ;
        RECT 721.950 247.950 724.050 248.400 ;
        RECT 766.950 247.950 769.050 248.400 ;
        RECT 559.950 246.600 562.050 247.050 ;
        RECT 443.400 245.400 562.050 246.600 ;
        RECT 391.950 244.950 394.050 245.400 ;
        RECT 439.950 244.950 442.050 245.400 ;
        RECT 559.950 244.950 562.050 245.400 ;
        RECT 610.950 246.600 613.050 247.050 ;
        RECT 622.950 246.600 625.050 247.050 ;
        RECT 610.950 245.400 625.050 246.600 ;
        RECT 610.950 244.950 613.050 245.400 ;
        RECT 622.950 244.950 625.050 245.400 ;
        RECT 637.950 246.600 640.050 247.050 ;
        RECT 643.950 246.600 646.050 247.050 ;
        RECT 676.950 246.600 679.050 247.050 ;
        RECT 637.950 245.400 646.050 246.600 ;
        RECT 637.950 244.950 640.050 245.400 ;
        RECT 643.950 244.950 646.050 245.400 ;
        RECT 671.400 245.400 679.050 246.600 ;
        RECT 671.400 244.050 672.600 245.400 ;
        RECT 676.950 244.950 679.050 245.400 ;
        RECT 700.950 246.600 703.050 247.050 ;
        RECT 718.950 246.600 721.050 247.050 ;
        RECT 733.950 246.600 736.050 247.050 ;
        RECT 700.950 245.400 717.600 246.600 ;
        RECT 700.950 244.950 703.050 245.400 ;
        RECT 16.950 243.600 19.050 244.050 ;
        RECT 25.950 243.600 28.050 244.050 ;
        RECT 16.950 242.400 28.050 243.600 ;
        RECT 16.950 241.950 19.050 242.400 ;
        RECT 25.950 241.950 28.050 242.400 ;
        RECT 43.950 243.600 46.050 244.050 ;
        RECT 79.950 243.600 82.050 244.050 ;
        RECT 88.950 243.600 91.050 244.050 ;
        RECT 94.950 243.600 97.050 244.050 ;
        RECT 43.950 242.400 60.600 243.600 ;
        RECT 43.950 241.950 46.050 242.400 ;
        RECT 22.950 238.950 25.050 241.050 ;
        RECT 55.950 240.600 58.050 241.050 ;
        RECT 32.400 239.400 58.050 240.600 ;
        RECT 23.400 237.600 24.600 238.950 ;
        RECT 32.400 238.050 33.600 239.400 ;
        RECT 55.950 238.950 58.050 239.400 ;
        RECT 8.400 236.400 24.600 237.600 ;
        RECT 8.400 235.050 9.600 236.400 ;
        RECT 31.950 235.950 34.050 238.050 ;
        RECT 59.400 237.600 60.600 242.400 ;
        RECT 79.950 242.400 97.050 243.600 ;
        RECT 79.950 241.950 82.050 242.400 ;
        RECT 88.950 241.950 91.050 242.400 ;
        RECT 94.950 241.950 97.050 242.400 ;
        RECT 121.950 243.600 124.050 244.050 ;
        RECT 139.950 243.600 142.050 244.050 ;
        RECT 142.950 243.600 145.050 244.050 ;
        RECT 121.950 242.400 145.050 243.600 ;
        RECT 121.950 241.950 124.050 242.400 ;
        RECT 139.950 241.950 142.050 242.400 ;
        RECT 142.950 241.950 145.050 242.400 ;
        RECT 148.950 243.600 151.050 244.050 ;
        RECT 154.950 243.600 157.050 244.050 ;
        RECT 172.950 243.600 175.050 244.050 ;
        RECT 148.950 242.400 175.050 243.600 ;
        RECT 148.950 241.950 151.050 242.400 ;
        RECT 154.950 241.950 157.050 242.400 ;
        RECT 172.950 241.950 175.050 242.400 ;
        RECT 175.950 243.600 178.050 244.050 ;
        RECT 202.950 243.600 205.050 244.050 ;
        RECT 223.950 243.600 226.050 244.050 ;
        RECT 268.950 243.600 271.050 244.050 ;
        RECT 175.950 242.400 192.600 243.600 ;
        RECT 175.950 241.950 178.050 242.400 ;
        RECT 73.950 240.600 76.050 241.050 ;
        RECT 85.950 240.600 88.050 241.050 ;
        RECT 73.950 239.400 88.050 240.600 ;
        RECT 73.950 238.950 76.050 239.400 ;
        RECT 85.950 238.950 88.050 239.400 ;
        RECT 112.950 240.600 115.050 241.050 ;
        RECT 124.950 240.600 127.050 241.050 ;
        RECT 130.950 240.600 133.050 241.050 ;
        RECT 112.950 239.400 127.050 240.600 ;
        RECT 112.950 238.950 115.050 239.400 ;
        RECT 116.400 238.050 117.600 239.400 ;
        RECT 124.950 238.950 127.050 239.400 ;
        RECT 128.400 239.400 133.050 240.600 ;
        RECT 70.950 237.600 73.050 238.050 ;
        RECT 59.400 236.400 73.050 237.600 ;
        RECT 70.950 235.950 73.050 236.400 ;
        RECT 73.950 235.950 76.050 238.050 ;
        RECT 94.950 237.600 97.050 238.050 ;
        RECT 94.950 236.400 99.600 237.600 ;
        RECT 94.950 235.950 97.050 236.400 ;
        RECT 7.950 232.950 10.050 235.050 ;
        RECT 10.950 234.600 13.050 235.050 ;
        RECT 22.950 234.600 25.050 235.050 ;
        RECT 34.950 234.600 37.050 235.050 ;
        RECT 10.950 233.400 37.050 234.600 ;
        RECT 10.950 232.950 13.050 233.400 ;
        RECT 22.950 232.950 25.050 233.400 ;
        RECT 34.950 232.950 37.050 233.400 ;
        RECT 67.950 234.600 70.050 235.050 ;
        RECT 74.400 234.600 75.600 235.950 ;
        RECT 67.950 233.400 75.600 234.600 ;
        RECT 67.950 232.950 70.050 233.400 ;
        RECT 98.400 232.050 99.600 236.400 ;
        RECT 115.950 235.950 118.050 238.050 ;
        RECT 128.400 237.600 129.600 239.400 ;
        RECT 130.950 238.950 133.050 239.400 ;
        RECT 148.950 238.950 151.050 241.050 ;
        RECT 184.950 240.600 187.050 241.050 ;
        RECT 182.400 239.400 187.050 240.600 ;
        RECT 119.400 236.400 129.600 237.600 ;
        RECT 149.400 237.600 150.600 238.950 ;
        RECT 160.950 237.600 163.050 238.050 ;
        RECT 149.400 236.400 163.050 237.600 ;
        RECT 109.950 234.600 112.050 235.050 ;
        RECT 119.400 234.600 120.600 236.400 ;
        RECT 160.950 235.950 163.050 236.400 ;
        RECT 172.950 237.600 175.050 238.050 ;
        RECT 182.400 237.600 183.600 239.400 ;
        RECT 184.950 238.950 187.050 239.400 ;
        RECT 187.950 238.950 190.050 241.050 ;
        RECT 191.400 240.600 192.600 242.400 ;
        RECT 202.950 242.400 271.050 243.600 ;
        RECT 202.950 241.950 205.050 242.400 ;
        RECT 223.950 241.950 226.050 242.400 ;
        RECT 268.950 241.950 271.050 242.400 ;
        RECT 277.950 243.600 280.050 244.050 ;
        RECT 301.950 243.600 304.050 244.050 ;
        RECT 277.950 242.400 304.050 243.600 ;
        RECT 277.950 241.950 280.050 242.400 ;
        RECT 301.950 241.950 304.050 242.400 ;
        RECT 325.950 243.600 328.050 244.050 ;
        RECT 352.950 243.600 355.050 244.050 ;
        RECT 325.950 242.400 355.050 243.600 ;
        RECT 325.950 241.950 328.050 242.400 ;
        RECT 352.950 241.950 355.050 242.400 ;
        RECT 373.950 243.600 376.050 244.050 ;
        RECT 412.950 243.600 415.050 244.050 ;
        RECT 373.950 242.400 415.050 243.600 ;
        RECT 373.950 241.950 376.050 242.400 ;
        RECT 412.950 241.950 415.050 242.400 ;
        RECT 442.950 243.600 445.050 244.050 ;
        RECT 460.950 243.600 463.050 244.050 ;
        RECT 478.950 243.600 481.050 244.050 ;
        RECT 490.950 243.600 493.050 244.050 ;
        RECT 442.950 242.400 463.050 243.600 ;
        RECT 442.950 241.950 445.050 242.400 ;
        RECT 460.950 241.950 463.050 242.400 ;
        RECT 464.400 242.400 474.600 243.600 ;
        RECT 208.950 240.600 211.050 241.050 ;
        RECT 191.400 239.400 211.050 240.600 ;
        RECT 208.950 238.950 211.050 239.400 ;
        RECT 220.950 238.950 223.050 241.050 ;
        RECT 229.950 240.600 232.050 241.050 ;
        RECT 250.950 240.600 253.050 241.050 ;
        RECT 229.950 239.400 253.050 240.600 ;
        RECT 229.950 238.950 232.050 239.400 ;
        RECT 172.950 236.400 183.600 237.600 ;
        RECT 188.400 237.600 189.600 238.950 ;
        RECT 188.400 236.400 195.600 237.600 ;
        RECT 172.950 235.950 175.050 236.400 ;
        RECT 194.400 235.050 195.600 236.400 ;
        RECT 221.400 235.050 222.600 238.950 ;
        RECT 236.400 235.050 237.600 239.400 ;
        RECT 250.950 238.950 253.050 239.400 ;
        RECT 253.950 240.600 256.050 241.050 ;
        RECT 262.950 240.600 265.050 241.050 ;
        RECT 253.950 239.400 265.050 240.600 ;
        RECT 253.950 238.950 256.050 239.400 ;
        RECT 262.950 238.950 265.050 239.400 ;
        RECT 265.950 240.600 268.050 241.050 ;
        RECT 271.950 240.600 274.050 241.050 ;
        RECT 283.950 240.600 286.050 241.050 ;
        RECT 265.950 239.400 274.050 240.600 ;
        RECT 265.950 238.950 268.050 239.400 ;
        RECT 271.950 238.950 274.050 239.400 ;
        RECT 275.400 239.400 286.050 240.600 ;
        RECT 268.950 237.600 271.050 238.050 ;
        RECT 275.400 237.600 276.600 239.400 ;
        RECT 283.950 238.950 286.050 239.400 ;
        RECT 286.950 238.950 289.050 241.050 ;
        RECT 304.950 240.600 307.050 241.050 ;
        RECT 290.400 239.400 307.050 240.600 ;
        RECT 287.400 237.600 288.600 238.950 ;
        RECT 290.400 238.050 291.600 239.400 ;
        RECT 304.950 238.950 307.050 239.400 ;
        RECT 310.950 240.600 313.050 241.050 ;
        RECT 322.950 240.600 325.050 241.050 ;
        RECT 310.950 239.400 325.050 240.600 ;
        RECT 310.950 238.950 313.050 239.400 ;
        RECT 322.950 238.950 325.050 239.400 ;
        RECT 346.950 240.600 349.050 241.050 ;
        RECT 382.950 240.600 385.050 241.050 ;
        RECT 346.950 239.400 385.050 240.600 ;
        RECT 346.950 238.950 349.050 239.400 ;
        RECT 362.400 238.050 363.600 239.400 ;
        RECT 382.950 238.950 385.050 239.400 ;
        RECT 415.950 240.600 418.050 241.050 ;
        RECT 448.950 240.600 451.050 241.050 ;
        RECT 464.400 240.600 465.600 242.400 ;
        RECT 415.950 239.400 444.600 240.600 ;
        RECT 415.950 238.950 418.050 239.400 ;
        RECT 242.400 236.400 276.600 237.600 ;
        RECT 278.400 236.400 288.600 237.600 ;
        RECT 242.400 235.050 243.600 236.400 ;
        RECT 268.950 235.950 271.050 236.400 ;
        RECT 109.950 233.400 120.600 234.600 ;
        RECT 127.950 234.600 130.050 235.050 ;
        RECT 139.950 234.600 142.050 235.050 ;
        RECT 127.950 233.400 142.050 234.600 ;
        RECT 109.950 232.950 112.050 233.400 ;
        RECT 127.950 232.950 130.050 233.400 ;
        RECT 139.950 232.950 142.050 233.400 ;
        RECT 157.950 234.600 160.050 235.050 ;
        RECT 169.950 234.600 172.050 235.050 ;
        RECT 157.950 233.400 172.050 234.600 ;
        RECT 157.950 232.950 160.050 233.400 ;
        RECT 169.950 232.950 172.050 233.400 ;
        RECT 193.950 232.950 196.050 235.050 ;
        RECT 220.950 232.950 223.050 235.050 ;
        RECT 235.950 232.950 238.050 235.050 ;
        RECT 241.950 232.950 244.050 235.050 ;
        RECT 274.950 234.600 277.050 235.050 ;
        RECT 278.400 234.600 279.600 236.400 ;
        RECT 289.950 235.950 292.050 238.050 ;
        RECT 301.950 237.600 304.050 238.050 ;
        RECT 361.950 237.600 364.050 238.050 ;
        RECT 394.950 237.600 397.050 238.050 ;
        RECT 301.950 236.400 364.050 237.600 ;
        RECT 301.950 235.950 304.050 236.400 ;
        RECT 361.950 235.950 364.050 236.400 ;
        RECT 389.400 236.400 397.050 237.600 ;
        RECT 389.400 235.050 390.600 236.400 ;
        RECT 394.950 235.950 397.050 236.400 ;
        RECT 412.950 237.600 415.050 238.050 ;
        RECT 439.950 237.600 442.050 238.050 ;
        RECT 412.950 236.400 426.600 237.600 ;
        RECT 412.950 235.950 415.050 236.400 ;
        RECT 425.400 235.050 426.600 236.400 ;
        RECT 431.400 236.400 442.050 237.600 ;
        RECT 431.400 235.050 432.600 236.400 ;
        RECT 439.950 235.950 442.050 236.400 ;
        RECT 310.950 234.600 313.050 235.050 ;
        RECT 274.950 233.400 313.050 234.600 ;
        RECT 274.950 232.950 277.050 233.400 ;
        RECT 310.950 232.950 313.050 233.400 ;
        RECT 316.950 234.600 319.050 235.050 ;
        RECT 364.950 234.600 367.050 235.050 ;
        RECT 316.950 233.400 367.050 234.600 ;
        RECT 316.950 232.950 319.050 233.400 ;
        RECT 364.950 232.950 367.050 233.400 ;
        RECT 379.950 234.600 382.050 235.050 ;
        RECT 388.950 234.600 391.050 235.050 ;
        RECT 379.950 233.400 391.050 234.600 ;
        RECT 379.950 232.950 382.050 233.400 ;
        RECT 388.950 232.950 391.050 233.400 ;
        RECT 409.950 234.600 412.050 235.050 ;
        RECT 415.950 234.600 418.050 235.050 ;
        RECT 418.950 234.600 421.050 235.050 ;
        RECT 409.950 233.400 421.050 234.600 ;
        RECT 409.950 232.950 412.050 233.400 ;
        RECT 415.950 232.950 418.050 233.400 ;
        RECT 418.950 232.950 421.050 233.400 ;
        RECT 424.950 232.950 427.050 235.050 ;
        RECT 430.950 232.950 433.050 235.050 ;
        RECT 443.400 234.600 444.600 239.400 ;
        RECT 448.950 239.400 465.600 240.600 ;
        RECT 448.950 238.950 451.050 239.400 ;
        RECT 469.950 238.950 472.050 241.050 ;
        RECT 473.400 240.600 474.600 242.400 ;
        RECT 478.950 242.400 493.050 243.600 ;
        RECT 478.950 241.950 481.050 242.400 ;
        RECT 490.950 241.950 493.050 242.400 ;
        RECT 529.950 243.600 532.050 244.050 ;
        RECT 544.950 243.600 547.050 244.050 ;
        RECT 529.950 242.400 547.050 243.600 ;
        RECT 529.950 241.950 532.050 242.400 ;
        RECT 544.950 241.950 547.050 242.400 ;
        RECT 547.950 243.600 550.050 244.050 ;
        RECT 553.950 243.600 556.050 244.050 ;
        RECT 583.950 243.600 586.050 244.050 ;
        RECT 547.950 242.400 556.050 243.600 ;
        RECT 547.950 241.950 550.050 242.400 ;
        RECT 553.950 241.950 556.050 242.400 ;
        RECT 575.400 242.400 586.050 243.600 ;
        RECT 493.950 240.600 496.050 241.050 ;
        RECT 505.950 240.600 508.050 241.050 ;
        RECT 514.950 240.600 517.050 241.050 ;
        RECT 473.400 239.400 517.050 240.600 ;
        RECT 493.950 238.950 496.050 239.400 ;
        RECT 505.950 238.950 508.050 239.400 ;
        RECT 514.950 238.950 517.050 239.400 ;
        RECT 523.950 240.600 526.050 241.050 ;
        RECT 535.950 240.600 538.050 241.050 ;
        RECT 523.950 239.400 538.050 240.600 ;
        RECT 523.950 238.950 526.050 239.400 ;
        RECT 535.950 238.950 538.050 239.400 ;
        RECT 544.950 240.600 547.050 241.050 ;
        RECT 553.950 240.600 556.050 241.050 ;
        RECT 544.950 239.400 556.050 240.600 ;
        RECT 544.950 238.950 547.050 239.400 ;
        RECT 553.950 238.950 556.050 239.400 ;
        RECT 562.950 238.950 565.050 241.050 ;
        RECT 445.950 237.600 448.050 238.050 ;
        RECT 451.950 237.600 454.050 238.050 ;
        RECT 445.950 236.400 454.050 237.600 ;
        RECT 445.950 235.950 448.050 236.400 ;
        RECT 451.950 235.950 454.050 236.400 ;
        RECT 470.400 235.050 471.600 238.950 ;
        RECT 502.950 237.600 505.050 238.050 ;
        RECT 494.400 236.400 505.050 237.600 ;
        RECT 494.400 235.050 495.600 236.400 ;
        RECT 502.950 235.950 505.050 236.400 ;
        RECT 511.950 237.600 514.050 238.050 ;
        RECT 526.950 237.600 529.050 238.050 ;
        RECT 563.400 237.600 564.600 238.950 ;
        RECT 565.950 237.600 568.050 238.050 ;
        RECT 511.950 236.400 529.050 237.600 ;
        RECT 511.950 235.950 514.050 236.400 ;
        RECT 526.950 235.950 529.050 236.400 ;
        RECT 548.400 236.400 568.050 237.600 ;
        RECT 463.950 234.600 466.050 235.050 ;
        RECT 443.400 233.400 466.050 234.600 ;
        RECT 463.950 232.950 466.050 233.400 ;
        RECT 469.950 232.950 472.050 235.050 ;
        RECT 493.950 232.950 496.050 235.050 ;
        RECT 523.950 234.600 526.050 235.050 ;
        RECT 548.400 234.600 549.600 236.400 ;
        RECT 565.950 235.950 568.050 236.400 ;
        RECT 571.950 235.950 574.050 238.050 ;
        RECT 575.400 237.600 576.600 242.400 ;
        RECT 583.950 241.950 586.050 242.400 ;
        RECT 586.950 243.600 589.050 244.050 ;
        RECT 592.950 243.600 595.050 244.050 ;
        RECT 619.950 243.600 622.050 244.050 ;
        RECT 586.950 242.400 595.050 243.600 ;
        RECT 586.950 241.950 589.050 242.400 ;
        RECT 592.950 241.950 595.050 242.400 ;
        RECT 617.400 242.400 622.050 243.600 ;
        RECT 577.950 240.600 580.050 241.050 ;
        RECT 577.950 239.400 582.600 240.600 ;
        RECT 577.950 238.950 580.050 239.400 ;
        RECT 577.950 237.600 580.050 238.050 ;
        RECT 575.400 236.400 580.050 237.600 ;
        RECT 581.400 237.600 582.600 239.400 ;
        RECT 601.950 238.950 604.050 241.050 ;
        RECT 613.950 238.950 616.050 241.050 ;
        RECT 589.950 237.600 592.050 238.050 ;
        RECT 602.400 237.600 603.600 238.950 ;
        RECT 581.400 236.400 592.050 237.600 ;
        RECT 577.950 235.950 580.050 236.400 ;
        RECT 589.950 235.950 592.050 236.400 ;
        RECT 593.400 236.400 603.600 237.600 ;
        RECT 604.950 237.600 607.050 238.050 ;
        RECT 610.950 237.600 613.050 238.050 ;
        RECT 604.950 236.400 613.050 237.600 ;
        RECT 523.950 233.400 549.600 234.600 ;
        RECT 562.950 234.600 565.050 235.050 ;
        RECT 568.950 234.600 571.050 235.050 ;
        RECT 562.950 233.400 571.050 234.600 ;
        RECT 572.400 234.600 573.600 235.950 ;
        RECT 593.400 235.050 594.600 236.400 ;
        RECT 604.950 235.950 607.050 236.400 ;
        RECT 610.950 235.950 613.050 236.400 ;
        RECT 580.950 234.600 583.050 235.050 ;
        RECT 572.400 233.400 583.050 234.600 ;
        RECT 523.950 232.950 526.050 233.400 ;
        RECT 562.950 232.950 565.050 233.400 ;
        RECT 568.950 232.950 571.050 233.400 ;
        RECT 580.950 232.950 583.050 233.400 ;
        RECT 592.950 232.950 595.050 235.050 ;
        RECT 595.950 234.600 598.050 235.050 ;
        RECT 601.950 234.600 604.050 235.050 ;
        RECT 595.950 233.400 604.050 234.600 ;
        RECT 595.950 232.950 598.050 233.400 ;
        RECT 601.950 232.950 604.050 233.400 ;
        RECT 607.950 234.600 610.050 235.050 ;
        RECT 614.400 234.600 615.600 238.950 ;
        RECT 607.950 233.400 615.600 234.600 ;
        RECT 617.400 234.600 618.600 242.400 ;
        RECT 619.950 241.950 622.050 242.400 ;
        RECT 625.950 243.600 628.050 244.050 ;
        RECT 649.950 243.600 652.050 244.050 ;
        RECT 625.950 242.400 652.050 243.600 ;
        RECT 625.950 241.950 628.050 242.400 ;
        RECT 649.950 241.950 652.050 242.400 ;
        RECT 655.950 243.600 658.050 244.050 ;
        RECT 667.950 243.600 670.050 244.050 ;
        RECT 655.950 242.400 670.050 243.600 ;
        RECT 655.950 241.950 658.050 242.400 ;
        RECT 667.950 241.950 670.050 242.400 ;
        RECT 670.950 241.950 673.050 244.050 ;
        RECT 673.950 243.600 676.050 244.050 ;
        RECT 691.950 243.600 694.050 244.050 ;
        RECT 673.950 242.400 694.050 243.600 ;
        RECT 673.950 241.950 676.050 242.400 ;
        RECT 691.950 241.950 694.050 242.400 ;
        RECT 694.950 243.600 697.050 244.050 ;
        RECT 709.950 243.600 712.050 244.050 ;
        RECT 694.950 242.400 712.050 243.600 ;
        RECT 716.400 243.600 717.600 245.400 ;
        RECT 718.950 245.400 736.050 246.600 ;
        RECT 718.950 244.950 721.050 245.400 ;
        RECT 733.950 244.950 736.050 245.400 ;
        RECT 721.950 243.600 724.050 244.050 ;
        RECT 727.950 243.600 730.050 244.050 ;
        RECT 716.400 242.400 720.600 243.600 ;
        RECT 694.950 241.950 697.050 242.400 ;
        RECT 709.950 241.950 712.050 242.400 ;
        RECT 655.950 240.600 658.050 241.050 ;
        RECT 647.400 239.400 658.050 240.600 ;
        RECT 619.950 237.600 622.050 238.050 ;
        RECT 647.400 237.600 648.600 239.400 ;
        RECT 655.950 238.950 658.050 239.400 ;
        RECT 661.950 240.600 664.050 241.050 ;
        RECT 661.950 239.400 675.600 240.600 ;
        RECT 661.950 238.950 664.050 239.400 ;
        RECT 674.400 238.050 675.600 239.400 ;
        RECT 676.950 238.950 679.050 241.050 ;
        RECT 682.950 240.600 685.050 241.050 ;
        RECT 694.950 240.600 697.050 241.050 ;
        RECT 712.950 240.600 715.050 241.050 ;
        RECT 682.950 239.400 697.050 240.600 ;
        RECT 682.950 238.950 685.050 239.400 ;
        RECT 694.950 238.950 697.050 239.400 ;
        RECT 704.400 239.400 715.050 240.600 ;
        RECT 719.400 240.600 720.600 242.400 ;
        RECT 721.950 242.400 730.050 243.600 ;
        RECT 721.950 241.950 724.050 242.400 ;
        RECT 727.950 241.950 730.050 242.400 ;
        RECT 736.950 243.600 739.050 244.050 ;
        RECT 760.950 243.600 763.050 244.050 ;
        RECT 736.950 242.400 763.050 243.600 ;
        RECT 736.950 241.950 739.050 242.400 ;
        RECT 760.950 241.950 763.050 242.400 ;
        RECT 745.950 240.600 748.050 241.050 ;
        RECT 719.400 239.400 748.050 240.600 ;
        RECT 619.950 236.400 648.600 237.600 ;
        RECT 649.950 237.600 652.050 238.050 ;
        RECT 649.950 236.400 660.600 237.600 ;
        RECT 619.950 235.950 622.050 236.400 ;
        RECT 619.950 234.600 622.050 235.050 ;
        RECT 617.400 233.400 622.050 234.600 ;
        RECT 638.400 234.600 639.600 236.400 ;
        RECT 649.950 235.950 652.050 236.400 ;
        RECT 646.950 234.600 649.050 235.050 ;
        RECT 638.400 233.400 649.050 234.600 ;
        RECT 607.950 232.950 610.050 233.400 ;
        RECT 619.950 232.950 622.050 233.400 ;
        RECT 646.950 232.950 649.050 233.400 ;
        RECT 70.950 231.600 73.050 232.050 ;
        RECT 82.950 231.600 85.050 232.050 ;
        RECT 70.950 230.400 85.050 231.600 ;
        RECT 70.950 229.950 73.050 230.400 ;
        RECT 82.950 229.950 85.050 230.400 ;
        RECT 97.950 229.950 100.050 232.050 ;
        RECT 112.950 231.600 115.050 232.050 ;
        RECT 121.950 231.600 124.050 232.050 ;
        RECT 133.950 231.600 136.050 232.050 ;
        RECT 112.950 230.400 136.050 231.600 ;
        RECT 112.950 229.950 115.050 230.400 ;
        RECT 121.950 229.950 124.050 230.400 ;
        RECT 133.950 229.950 136.050 230.400 ;
        RECT 202.950 231.600 205.050 232.050 ;
        RECT 205.950 231.600 208.050 232.050 ;
        RECT 226.950 231.600 229.050 232.050 ;
        RECT 241.950 231.600 244.050 232.050 ;
        RECT 244.950 231.600 247.050 232.050 ;
        RECT 202.950 230.400 247.050 231.600 ;
        RECT 202.950 229.950 205.050 230.400 ;
        RECT 205.950 229.950 208.050 230.400 ;
        RECT 226.950 229.950 229.050 230.400 ;
        RECT 241.950 229.950 244.050 230.400 ;
        RECT 244.950 229.950 247.050 230.400 ;
        RECT 286.950 231.600 289.050 232.050 ;
        RECT 301.950 231.600 304.050 232.050 ;
        RECT 286.950 230.400 304.050 231.600 ;
        RECT 286.950 229.950 289.050 230.400 ;
        RECT 301.950 229.950 304.050 230.400 ;
        RECT 319.950 231.600 322.050 232.050 ;
        RECT 376.950 231.600 379.050 232.050 ;
        RECT 319.950 230.400 379.050 231.600 ;
        RECT 319.950 229.950 322.050 230.400 ;
        RECT 376.950 229.950 379.050 230.400 ;
        RECT 403.950 231.600 406.050 232.050 ;
        RECT 451.950 231.600 454.050 232.050 ;
        RECT 403.950 230.400 454.050 231.600 ;
        RECT 403.950 229.950 406.050 230.400 ;
        RECT 451.950 229.950 454.050 230.400 ;
        RECT 475.950 231.600 478.050 232.050 ;
        RECT 481.950 231.600 484.050 232.050 ;
        RECT 475.950 230.400 484.050 231.600 ;
        RECT 475.950 229.950 478.050 230.400 ;
        RECT 481.950 229.950 484.050 230.400 ;
        RECT 628.950 231.600 631.050 232.050 ;
        RECT 637.950 231.600 640.050 232.050 ;
        RECT 628.950 230.400 640.050 231.600 ;
        RECT 659.400 231.600 660.600 236.400 ;
        RECT 673.950 235.950 676.050 238.050 ;
        RECT 664.950 234.600 667.050 235.050 ;
        RECT 677.400 234.600 678.600 238.950 ;
        RECT 704.400 237.600 705.600 239.400 ;
        RECT 712.950 238.950 715.050 239.400 ;
        RECT 745.950 238.950 748.050 239.400 ;
        RECT 760.950 240.600 763.050 241.050 ;
        RECT 760.950 239.400 771.600 240.600 ;
        RECT 760.950 238.950 763.050 239.400 ;
        RECT 712.950 237.600 715.050 238.050 ;
        RECT 736.950 237.600 739.050 238.050 ;
        RECT 683.400 236.400 705.600 237.600 ;
        RECT 707.400 236.400 739.050 237.600 ;
        RECT 683.400 235.050 684.600 236.400 ;
        RECT 664.950 233.400 678.600 234.600 ;
        RECT 664.950 232.950 667.050 233.400 ;
        RECT 682.950 232.950 685.050 235.050 ;
        RECT 703.950 234.600 706.050 235.050 ;
        RECT 707.400 234.600 708.600 236.400 ;
        RECT 712.950 235.950 715.050 236.400 ;
        RECT 736.950 235.950 739.050 236.400 ;
        RECT 742.950 235.950 745.050 238.050 ;
        RECT 748.950 237.600 751.050 238.050 ;
        RECT 763.950 237.600 766.050 238.050 ;
        RECT 748.950 236.400 766.050 237.600 ;
        RECT 748.950 235.950 751.050 236.400 ;
        RECT 763.950 235.950 766.050 236.400 ;
        RECT 766.950 235.950 769.050 238.050 ;
        RECT 686.400 233.400 708.600 234.600 ;
        RECT 721.950 234.600 724.050 235.050 ;
        RECT 743.400 234.600 744.600 235.950 ;
        RECT 757.950 234.600 760.050 235.050 ;
        RECT 767.400 234.600 768.600 235.950 ;
        RECT 721.950 233.400 760.050 234.600 ;
        RECT 686.400 231.600 687.600 233.400 ;
        RECT 703.950 232.950 706.050 233.400 ;
        RECT 721.950 232.950 724.050 233.400 ;
        RECT 725.400 232.050 726.600 233.400 ;
        RECT 757.950 232.950 760.050 233.400 ;
        RECT 764.400 233.400 768.600 234.600 ;
        RECT 659.400 230.400 687.600 231.600 ;
        RECT 697.950 231.600 700.050 232.050 ;
        RECT 706.950 231.600 709.050 232.050 ;
        RECT 697.950 230.400 709.050 231.600 ;
        RECT 628.950 229.950 631.050 230.400 ;
        RECT 637.950 229.950 640.050 230.400 ;
        RECT 697.950 229.950 700.050 230.400 ;
        RECT 706.950 229.950 709.050 230.400 ;
        RECT 724.950 229.950 727.050 232.050 ;
        RECT 742.950 231.600 745.050 232.050 ;
        RECT 748.950 231.600 751.050 232.050 ;
        RECT 742.950 230.400 751.050 231.600 ;
        RECT 742.950 229.950 745.050 230.400 ;
        RECT 748.950 229.950 751.050 230.400 ;
        RECT 760.950 231.600 763.050 232.050 ;
        RECT 764.400 231.600 765.600 233.400 ;
        RECT 760.950 230.400 765.600 231.600 ;
        RECT 766.950 231.600 769.050 232.050 ;
        RECT 770.400 231.600 771.600 239.400 ;
        RECT 766.950 230.400 771.600 231.600 ;
        RECT 760.950 229.950 763.050 230.400 ;
        RECT 766.950 229.950 769.050 230.400 ;
        RECT 85.950 228.600 88.050 229.050 ;
        RECT 103.950 228.600 106.050 229.050 ;
        RECT 85.950 227.400 106.050 228.600 ;
        RECT 85.950 226.950 88.050 227.400 ;
        RECT 103.950 226.950 106.050 227.400 ;
        RECT 199.950 228.600 202.050 229.050 ;
        RECT 205.950 228.600 208.050 229.050 ;
        RECT 199.950 227.400 208.050 228.600 ;
        RECT 199.950 226.950 202.050 227.400 ;
        RECT 205.950 226.950 208.050 227.400 ;
        RECT 208.950 228.600 211.050 229.050 ;
        RECT 223.950 228.600 226.050 229.050 ;
        RECT 208.950 227.400 226.050 228.600 ;
        RECT 208.950 226.950 211.050 227.400 ;
        RECT 223.950 226.950 226.050 227.400 ;
        RECT 256.950 228.600 259.050 229.050 ;
        RECT 316.950 228.600 319.050 229.050 ;
        RECT 334.950 228.600 337.050 229.050 ;
        RECT 256.950 227.400 319.050 228.600 ;
        RECT 256.950 226.950 259.050 227.400 ;
        RECT 316.950 226.950 319.050 227.400 ;
        RECT 320.400 227.400 337.050 228.600 ;
        RECT 58.950 225.600 61.050 226.050 ;
        RECT 97.950 225.600 100.050 226.050 ;
        RECT 58.950 224.400 100.050 225.600 ;
        RECT 58.950 223.950 61.050 224.400 ;
        RECT 97.950 223.950 100.050 224.400 ;
        RECT 154.950 225.600 157.050 226.050 ;
        RECT 187.950 225.600 190.050 226.050 ;
        RECT 190.950 225.600 193.050 226.050 ;
        RECT 259.950 225.600 262.050 226.050 ;
        RECT 154.950 224.400 262.050 225.600 ;
        RECT 154.950 223.950 157.050 224.400 ;
        RECT 187.950 223.950 190.050 224.400 ;
        RECT 190.950 223.950 193.050 224.400 ;
        RECT 259.950 223.950 262.050 224.400 ;
        RECT 280.950 225.600 283.050 226.050 ;
        RECT 307.950 225.600 310.050 226.050 ;
        RECT 320.400 225.600 321.600 227.400 ;
        RECT 334.950 226.950 337.050 227.400 ;
        RECT 412.950 228.600 415.050 229.050 ;
        RECT 523.950 228.600 526.050 229.050 ;
        RECT 412.950 227.400 526.050 228.600 ;
        RECT 412.950 226.950 415.050 227.400 ;
        RECT 523.950 226.950 526.050 227.400 ;
        RECT 526.950 228.600 529.050 229.050 ;
        RECT 550.950 228.600 553.050 229.050 ;
        RECT 595.950 228.600 598.050 229.050 ;
        RECT 526.950 227.400 553.050 228.600 ;
        RECT 526.950 226.950 529.050 227.400 ;
        RECT 550.950 226.950 553.050 227.400 ;
        RECT 584.400 227.400 598.050 228.600 ;
        RECT 280.950 224.400 321.600 225.600 ;
        RECT 322.950 225.600 325.050 226.050 ;
        RECT 343.950 225.600 346.050 226.050 ;
        RECT 322.950 224.400 346.050 225.600 ;
        RECT 280.950 223.950 283.050 224.400 ;
        RECT 307.950 223.950 310.050 224.400 ;
        RECT 322.950 223.950 325.050 224.400 ;
        RECT 343.950 223.950 346.050 224.400 ;
        RECT 367.950 225.600 370.050 226.050 ;
        RECT 406.950 225.600 409.050 226.050 ;
        RECT 367.950 224.400 409.050 225.600 ;
        RECT 367.950 223.950 370.050 224.400 ;
        RECT 406.950 223.950 409.050 224.400 ;
        RECT 418.950 225.600 421.050 226.050 ;
        RECT 538.950 225.600 541.050 226.050 ;
        RECT 584.400 225.600 585.600 227.400 ;
        RECT 595.950 226.950 598.050 227.400 ;
        RECT 610.950 228.600 613.050 229.050 ;
        RECT 631.950 228.600 634.050 229.050 ;
        RECT 652.950 228.600 655.050 229.050 ;
        RECT 661.950 228.600 664.050 229.050 ;
        RECT 610.950 227.400 664.050 228.600 ;
        RECT 610.950 226.950 613.050 227.400 ;
        RECT 631.950 226.950 634.050 227.400 ;
        RECT 652.950 226.950 655.050 227.400 ;
        RECT 661.950 226.950 664.050 227.400 ;
        RECT 676.950 228.600 679.050 229.050 ;
        RECT 682.950 228.600 685.050 229.050 ;
        RECT 676.950 227.400 685.050 228.600 ;
        RECT 676.950 226.950 679.050 227.400 ;
        RECT 682.950 226.950 685.050 227.400 ;
        RECT 700.950 228.600 703.050 229.050 ;
        RECT 757.950 228.600 760.050 229.050 ;
        RECT 700.950 227.400 760.050 228.600 ;
        RECT 700.950 226.950 703.050 227.400 ;
        RECT 757.950 226.950 760.050 227.400 ;
        RECT 418.950 224.400 585.600 225.600 ;
        RECT 589.950 225.600 592.050 226.050 ;
        RECT 634.950 225.600 637.050 226.050 ;
        RECT 664.950 225.600 667.050 226.050 ;
        RECT 589.950 224.400 667.050 225.600 ;
        RECT 418.950 223.950 421.050 224.400 ;
        RECT 538.950 223.950 541.050 224.400 ;
        RECT 589.950 223.950 592.050 224.400 ;
        RECT 634.950 223.950 637.050 224.400 ;
        RECT 664.950 223.950 667.050 224.400 ;
        RECT 685.950 225.600 688.050 226.050 ;
        RECT 727.950 225.600 730.050 226.050 ;
        RECT 685.950 224.400 730.050 225.600 ;
        RECT 685.950 223.950 688.050 224.400 ;
        RECT 727.950 223.950 730.050 224.400 ;
        RECT 757.950 225.600 760.050 226.050 ;
        RECT 769.950 225.600 772.050 226.050 ;
        RECT 757.950 224.400 772.050 225.600 ;
        RECT 757.950 223.950 760.050 224.400 ;
        RECT 769.950 223.950 772.050 224.400 ;
        RECT 133.950 222.600 136.050 223.050 ;
        RECT 193.950 222.600 196.050 223.050 ;
        RECT 226.950 222.600 229.050 223.050 ;
        RECT 253.950 222.600 256.050 223.050 ;
        RECT 133.950 221.400 256.050 222.600 ;
        RECT 133.950 220.950 136.050 221.400 ;
        RECT 193.950 220.950 196.050 221.400 ;
        RECT 226.950 220.950 229.050 221.400 ;
        RECT 253.950 220.950 256.050 221.400 ;
        RECT 307.950 222.600 310.050 223.050 ;
        RECT 379.950 222.600 382.050 223.050 ;
        RECT 307.950 221.400 382.050 222.600 ;
        RECT 307.950 220.950 310.050 221.400 ;
        RECT 379.950 220.950 382.050 221.400 ;
        RECT 385.950 222.600 388.050 223.050 ;
        RECT 421.950 222.600 424.050 223.050 ;
        RECT 385.950 221.400 424.050 222.600 ;
        RECT 385.950 220.950 388.050 221.400 ;
        RECT 421.950 220.950 424.050 221.400 ;
        RECT 484.950 222.600 487.050 223.050 ;
        RECT 541.950 222.600 544.050 223.050 ;
        RECT 484.950 221.400 544.050 222.600 ;
        RECT 484.950 220.950 487.050 221.400 ;
        RECT 541.950 220.950 544.050 221.400 ;
        RECT 595.950 222.600 598.050 223.050 ;
        RECT 637.950 222.600 640.050 223.050 ;
        RECT 595.950 221.400 640.050 222.600 ;
        RECT 595.950 220.950 598.050 221.400 ;
        RECT 637.950 220.950 640.050 221.400 ;
        RECT 640.950 222.600 643.050 223.050 ;
        RECT 661.950 222.600 664.050 223.050 ;
        RECT 640.950 221.400 664.050 222.600 ;
        RECT 640.950 220.950 643.050 221.400 ;
        RECT 661.950 220.950 664.050 221.400 ;
        RECT 679.950 222.600 682.050 223.050 ;
        RECT 745.950 222.600 748.050 223.050 ;
        RECT 679.950 221.400 748.050 222.600 ;
        RECT 679.950 220.950 682.050 221.400 ;
        RECT 745.950 220.950 748.050 221.400 ;
        RECT 193.950 219.600 196.050 220.050 ;
        RECT 217.950 219.600 220.050 220.050 ;
        RECT 193.950 218.400 220.050 219.600 ;
        RECT 193.950 217.950 196.050 218.400 ;
        RECT 217.950 217.950 220.050 218.400 ;
        RECT 229.950 219.600 232.050 220.050 ;
        RECT 274.950 219.600 277.050 220.050 ;
        RECT 229.950 218.400 277.050 219.600 ;
        RECT 229.950 217.950 232.050 218.400 ;
        RECT 274.950 217.950 277.050 218.400 ;
        RECT 295.950 219.600 298.050 220.050 ;
        RECT 373.950 219.600 376.050 220.050 ;
        RECT 295.950 218.400 376.050 219.600 ;
        RECT 295.950 217.950 298.050 218.400 ;
        RECT 373.950 217.950 376.050 218.400 ;
        RECT 385.950 219.600 388.050 220.050 ;
        RECT 454.950 219.600 457.050 220.050 ;
        RECT 385.950 218.400 457.050 219.600 ;
        RECT 385.950 217.950 388.050 218.400 ;
        RECT 454.950 217.950 457.050 218.400 ;
        RECT 478.950 219.600 481.050 220.050 ;
        RECT 505.950 219.600 508.050 220.050 ;
        RECT 520.950 219.600 523.050 220.050 ;
        RECT 478.950 218.400 523.050 219.600 ;
        RECT 478.950 217.950 481.050 218.400 ;
        RECT 505.950 217.950 508.050 218.400 ;
        RECT 520.950 217.950 523.050 218.400 ;
        RECT 583.950 219.600 586.050 220.050 ;
        RECT 646.950 219.600 649.050 220.050 ;
        RECT 583.950 218.400 649.050 219.600 ;
        RECT 583.950 217.950 586.050 218.400 ;
        RECT 646.950 217.950 649.050 218.400 ;
        RECT 658.950 219.600 661.050 220.050 ;
        RECT 688.950 219.600 691.050 220.050 ;
        RECT 658.950 218.400 691.050 219.600 ;
        RECT 658.950 217.950 661.050 218.400 ;
        RECT 688.950 217.950 691.050 218.400 ;
        RECT 745.950 219.600 748.050 220.050 ;
        RECT 751.950 219.600 754.050 220.050 ;
        RECT 745.950 218.400 754.050 219.600 ;
        RECT 745.950 217.950 748.050 218.400 ;
        RECT 751.950 217.950 754.050 218.400 ;
        RECT 220.950 216.600 223.050 217.050 ;
        RECT 238.950 216.600 241.050 217.050 ;
        RECT 220.950 215.400 241.050 216.600 ;
        RECT 220.950 214.950 223.050 215.400 ;
        RECT 238.950 214.950 241.050 215.400 ;
        RECT 367.950 216.600 370.050 217.050 ;
        RECT 397.950 216.600 400.050 217.050 ;
        RECT 367.950 215.400 400.050 216.600 ;
        RECT 367.950 214.950 370.050 215.400 ;
        RECT 397.950 214.950 400.050 215.400 ;
        RECT 400.950 216.600 403.050 217.050 ;
        RECT 442.950 216.600 445.050 217.050 ;
        RECT 400.950 215.400 445.050 216.600 ;
        RECT 400.950 214.950 403.050 215.400 ;
        RECT 442.950 214.950 445.050 215.400 ;
        RECT 481.950 216.600 484.050 217.050 ;
        RECT 508.950 216.600 511.050 217.050 ;
        RECT 481.950 215.400 511.050 216.600 ;
        RECT 481.950 214.950 484.050 215.400 ;
        RECT 508.950 214.950 511.050 215.400 ;
        RECT 532.950 216.600 535.050 217.050 ;
        RECT 610.950 216.600 613.050 217.050 ;
        RECT 532.950 215.400 613.050 216.600 ;
        RECT 532.950 214.950 535.050 215.400 ;
        RECT 610.950 214.950 613.050 215.400 ;
        RECT 673.950 216.600 676.050 217.050 ;
        RECT 700.950 216.600 703.050 217.050 ;
        RECT 673.950 215.400 703.050 216.600 ;
        RECT 673.950 214.950 676.050 215.400 ;
        RECT 700.950 214.950 703.050 215.400 ;
        RECT 748.950 216.600 751.050 217.050 ;
        RECT 763.950 216.600 766.050 217.050 ;
        RECT 748.950 215.400 766.050 216.600 ;
        RECT 748.950 214.950 751.050 215.400 ;
        RECT 763.950 214.950 766.050 215.400 ;
        RECT 259.950 213.600 262.050 214.050 ;
        RECT 304.950 213.600 307.050 214.050 ;
        RECT 259.950 212.400 307.050 213.600 ;
        RECT 259.950 211.950 262.050 212.400 ;
        RECT 304.950 211.950 307.050 212.400 ;
        RECT 310.950 213.600 313.050 214.050 ;
        RECT 319.950 213.600 322.050 214.050 ;
        RECT 310.950 212.400 322.050 213.600 ;
        RECT 310.950 211.950 313.050 212.400 ;
        RECT 319.950 211.950 322.050 212.400 ;
        RECT 349.950 213.600 352.050 214.050 ;
        RECT 370.950 213.600 373.050 214.050 ;
        RECT 385.950 213.600 388.050 214.050 ;
        RECT 349.950 212.400 388.050 213.600 ;
        RECT 349.950 211.950 352.050 212.400 ;
        RECT 370.950 211.950 373.050 212.400 ;
        RECT 385.950 211.950 388.050 212.400 ;
        RECT 457.950 213.600 460.050 214.050 ;
        RECT 553.950 213.600 556.050 214.050 ;
        RECT 457.950 212.400 556.050 213.600 ;
        RECT 457.950 211.950 460.050 212.400 ;
        RECT 553.950 211.950 556.050 212.400 ;
        RECT 592.950 213.600 595.050 214.050 ;
        RECT 604.950 213.600 607.050 214.050 ;
        RECT 697.950 213.600 700.050 214.050 ;
        RECT 592.950 212.400 700.050 213.600 ;
        RECT 592.950 211.950 595.050 212.400 ;
        RECT 604.950 211.950 607.050 212.400 ;
        RECT 697.950 211.950 700.050 212.400 ;
        RECT 706.950 213.600 709.050 214.050 ;
        RECT 712.950 213.600 715.050 214.050 ;
        RECT 736.950 213.600 739.050 214.050 ;
        RECT 706.950 212.400 739.050 213.600 ;
        RECT 706.950 211.950 709.050 212.400 ;
        RECT 712.950 211.950 715.050 212.400 ;
        RECT 736.950 211.950 739.050 212.400 ;
        RECT 748.950 213.600 751.050 214.050 ;
        RECT 760.950 213.600 763.050 214.050 ;
        RECT 769.950 213.600 772.050 214.050 ;
        RECT 748.950 212.400 772.050 213.600 ;
        RECT 748.950 211.950 751.050 212.400 ;
        RECT 760.950 211.950 763.050 212.400 ;
        RECT 769.950 211.950 772.050 212.400 ;
        RECT 1.950 210.600 4.050 211.050 ;
        RECT 52.950 210.600 55.050 211.050 ;
        RECT 1.950 209.400 55.050 210.600 ;
        RECT 1.950 208.950 4.050 209.400 ;
        RECT 52.950 208.950 55.050 209.400 ;
        RECT 211.950 210.600 214.050 211.050 ;
        RECT 214.950 210.600 217.050 211.050 ;
        RECT 235.950 210.600 238.050 211.050 ;
        RECT 274.950 210.600 277.050 211.050 ;
        RECT 307.950 210.600 310.050 211.050 ;
        RECT 211.950 209.400 273.600 210.600 ;
        RECT 211.950 208.950 214.050 209.400 ;
        RECT 214.950 208.950 217.050 209.400 ;
        RECT 235.950 208.950 238.050 209.400 ;
        RECT 250.950 207.600 253.050 208.050 ;
        RECT 268.950 207.600 271.050 208.050 ;
        RECT 250.950 206.400 271.050 207.600 ;
        RECT 272.400 207.600 273.600 209.400 ;
        RECT 274.950 209.400 310.050 210.600 ;
        RECT 274.950 208.950 277.050 209.400 ;
        RECT 307.950 208.950 310.050 209.400 ;
        RECT 310.950 210.600 313.050 211.050 ;
        RECT 346.950 210.600 349.050 211.050 ;
        RECT 400.950 210.600 403.050 211.050 ;
        RECT 310.950 209.400 403.050 210.600 ;
        RECT 310.950 208.950 313.050 209.400 ;
        RECT 346.950 208.950 349.050 209.400 ;
        RECT 400.950 208.950 403.050 209.400 ;
        RECT 403.950 210.600 406.050 211.050 ;
        RECT 418.950 210.600 421.050 211.050 ;
        RECT 403.950 209.400 421.050 210.600 ;
        RECT 403.950 208.950 406.050 209.400 ;
        RECT 418.950 208.950 421.050 209.400 ;
        RECT 475.950 210.600 478.050 211.050 ;
        RECT 520.950 210.600 523.050 211.050 ;
        RECT 475.950 209.400 523.050 210.600 ;
        RECT 475.950 208.950 478.050 209.400 ;
        RECT 520.950 208.950 523.050 209.400 ;
        RECT 535.950 210.600 538.050 211.050 ;
        RECT 547.950 210.600 550.050 211.050 ;
        RECT 535.950 209.400 550.050 210.600 ;
        RECT 535.950 208.950 538.050 209.400 ;
        RECT 547.950 208.950 550.050 209.400 ;
        RECT 550.950 208.950 553.050 211.050 ;
        RECT 574.950 210.600 577.050 211.050 ;
        RECT 592.950 210.600 595.050 211.050 ;
        RECT 574.950 209.400 595.050 210.600 ;
        RECT 574.950 208.950 577.050 209.400 ;
        RECT 592.950 208.950 595.050 209.400 ;
        RECT 598.950 210.600 601.050 211.050 ;
        RECT 640.950 210.600 643.050 211.050 ;
        RECT 598.950 209.400 643.050 210.600 ;
        RECT 598.950 208.950 601.050 209.400 ;
        RECT 640.950 208.950 643.050 209.400 ;
        RECT 670.950 210.600 673.050 211.050 ;
        RECT 691.950 210.600 694.050 211.050 ;
        RECT 670.950 209.400 694.050 210.600 ;
        RECT 670.950 208.950 673.050 209.400 ;
        RECT 691.950 208.950 694.050 209.400 ;
        RECT 733.950 210.600 736.050 211.050 ;
        RECT 745.950 210.600 748.050 211.050 ;
        RECT 733.950 209.400 748.050 210.600 ;
        RECT 733.950 208.950 736.050 209.400 ;
        RECT 745.950 208.950 748.050 209.400 ;
        RECT 313.950 207.600 316.050 208.050 ;
        RECT 331.950 207.600 334.050 208.050 ;
        RECT 272.400 206.400 334.050 207.600 ;
        RECT 250.950 205.950 253.050 206.400 ;
        RECT 268.950 205.950 271.050 206.400 ;
        RECT 313.950 205.950 316.050 206.400 ;
        RECT 331.950 205.950 334.050 206.400 ;
        RECT 355.950 207.600 358.050 208.050 ;
        RECT 373.950 207.600 376.050 208.050 ;
        RECT 406.950 207.600 409.050 208.050 ;
        RECT 421.950 207.600 424.050 208.050 ;
        RECT 355.950 206.400 372.600 207.600 ;
        RECT 355.950 205.950 358.050 206.400 ;
        RECT 1.950 204.600 4.050 205.050 ;
        RECT 10.950 204.600 13.050 205.050 ;
        RECT 1.950 203.400 13.050 204.600 ;
        RECT 1.950 202.950 4.050 203.400 ;
        RECT 10.950 202.950 13.050 203.400 ;
        RECT 64.950 204.600 67.050 205.050 ;
        RECT 94.950 204.600 97.050 205.050 ;
        RECT 160.950 204.600 163.050 205.050 ;
        RECT 64.950 203.400 97.050 204.600 ;
        RECT 64.950 202.950 67.050 203.400 ;
        RECT 94.950 202.950 97.050 203.400 ;
        RECT 149.400 203.400 163.050 204.600 ;
        RECT 1.950 201.600 4.050 202.050 ;
        RECT 7.950 201.600 10.050 202.050 ;
        RECT 1.950 200.400 10.050 201.600 ;
        RECT 1.950 199.950 4.050 200.400 ;
        RECT 7.950 199.950 10.050 200.400 ;
        RECT 31.950 199.950 34.050 202.050 ;
        RECT 67.950 201.600 70.050 202.050 ;
        RECT 82.950 201.600 85.050 202.050 ;
        RECT 67.950 200.400 85.050 201.600 ;
        RECT 67.950 199.950 70.050 200.400 ;
        RECT 82.950 199.950 85.050 200.400 ;
        RECT 136.950 201.600 139.050 202.050 ;
        RECT 142.950 201.600 145.050 202.050 ;
        RECT 136.950 200.400 145.050 201.600 ;
        RECT 136.950 199.950 139.050 200.400 ;
        RECT 142.950 199.950 145.050 200.400 ;
        RECT 4.950 198.600 7.050 199.050 ;
        RECT 19.950 198.600 22.050 199.050 ;
        RECT 4.950 197.400 27.600 198.600 ;
        RECT 4.950 196.950 7.050 197.400 ;
        RECT 19.950 196.950 22.050 197.400 ;
        RECT 26.400 196.050 27.600 197.400 ;
        RECT 28.950 196.950 31.050 199.050 ;
        RECT 1.950 195.600 4.050 196.050 ;
        RECT 7.950 195.600 10.050 196.050 ;
        RECT 1.950 194.400 10.050 195.600 ;
        RECT 1.950 193.950 4.050 194.400 ;
        RECT 7.950 193.950 10.050 194.400 ;
        RECT 25.950 193.950 28.050 196.050 ;
        RECT 4.950 192.600 7.050 193.050 ;
        RECT 10.950 192.600 13.050 193.050 ;
        RECT 4.950 191.400 13.050 192.600 ;
        RECT 4.950 190.950 7.050 191.400 ;
        RECT 10.950 190.950 13.050 191.400 ;
        RECT 13.950 189.600 16.050 190.050 ;
        RECT 29.400 189.600 30.600 196.950 ;
        RECT 32.400 196.050 33.600 199.950 ;
        RECT 34.950 198.600 37.050 199.050 ;
        RECT 37.950 198.600 40.050 199.050 ;
        RECT 43.950 198.600 46.050 199.050 ;
        RECT 34.950 197.400 46.050 198.600 ;
        RECT 34.950 196.950 37.050 197.400 ;
        RECT 37.950 196.950 40.050 197.400 ;
        RECT 43.950 196.950 46.050 197.400 ;
        RECT 46.950 198.600 49.050 199.050 ;
        RECT 61.950 198.600 64.050 199.050 ;
        RECT 46.950 197.400 64.050 198.600 ;
        RECT 46.950 196.950 49.050 197.400 ;
        RECT 61.950 196.950 64.050 197.400 ;
        RECT 73.950 196.950 76.050 199.050 ;
        RECT 79.950 198.600 82.050 199.050 ;
        RECT 91.950 198.600 94.050 199.050 ;
        RECT 79.950 197.400 94.050 198.600 ;
        RECT 79.950 196.950 82.050 197.400 ;
        RECT 91.950 196.950 94.050 197.400 ;
        RECT 106.950 198.600 109.050 199.050 ;
        RECT 130.950 198.600 133.050 199.050 ;
        RECT 145.950 198.600 148.050 199.050 ;
        RECT 106.950 197.400 148.050 198.600 ;
        RECT 106.950 196.950 109.050 197.400 ;
        RECT 130.950 196.950 133.050 197.400 ;
        RECT 145.950 196.950 148.050 197.400 ;
        RECT 31.950 193.950 34.050 196.050 ;
        RECT 58.950 195.600 61.050 196.050 ;
        RECT 74.400 195.600 75.600 196.950 ;
        RECT 149.400 196.050 150.600 203.400 ;
        RECT 160.950 202.950 163.050 203.400 ;
        RECT 253.950 204.600 256.050 205.050 ;
        RECT 286.950 204.600 289.050 205.050 ;
        RECT 253.950 203.400 289.050 204.600 ;
        RECT 253.950 202.950 256.050 203.400 ;
        RECT 286.950 202.950 289.050 203.400 ;
        RECT 292.950 204.600 295.050 205.050 ;
        RECT 331.950 204.600 334.050 205.050 ;
        RECT 340.950 204.600 343.050 205.050 ;
        RECT 367.950 204.600 370.050 205.050 ;
        RECT 292.950 203.400 330.600 204.600 ;
        RECT 292.950 202.950 295.050 203.400 ;
        RECT 151.950 199.950 154.050 202.050 ;
        RECT 166.950 201.600 169.050 202.050 ;
        RECT 175.950 201.600 178.050 202.050 ;
        RECT 187.950 201.600 190.050 202.050 ;
        RECT 166.950 200.400 190.050 201.600 ;
        RECT 166.950 199.950 169.050 200.400 ;
        RECT 175.950 199.950 178.050 200.400 ;
        RECT 187.950 199.950 190.050 200.400 ;
        RECT 190.950 201.600 193.050 202.050 ;
        RECT 196.950 201.600 199.050 202.050 ;
        RECT 190.950 200.400 199.050 201.600 ;
        RECT 190.950 199.950 193.050 200.400 ;
        RECT 196.950 199.950 199.050 200.400 ;
        RECT 208.950 199.950 211.050 202.050 ;
        RECT 217.950 201.600 220.050 202.050 ;
        RECT 232.950 201.600 235.050 202.050 ;
        RECT 217.950 200.400 235.050 201.600 ;
        RECT 217.950 199.950 220.050 200.400 ;
        RECT 232.950 199.950 235.050 200.400 ;
        RECT 238.950 199.950 241.050 202.050 ;
        RECT 247.950 201.600 250.050 202.050 ;
        RECT 265.950 201.600 268.050 202.050 ;
        RECT 247.950 200.400 268.050 201.600 ;
        RECT 247.950 199.950 250.050 200.400 ;
        RECT 265.950 199.950 268.050 200.400 ;
        RECT 280.950 201.600 283.050 202.050 ;
        RECT 286.950 201.600 289.050 202.050 ;
        RECT 295.950 201.600 298.050 202.050 ;
        RECT 280.950 200.400 285.600 201.600 ;
        RECT 280.950 199.950 283.050 200.400 ;
        RECT 152.400 196.050 153.600 199.950 ;
        RECT 154.950 196.950 157.050 199.050 ;
        RECT 160.950 198.600 163.050 199.050 ;
        RECT 181.950 198.600 184.050 199.050 ;
        RECT 199.950 198.600 202.050 199.050 ;
        RECT 160.950 197.400 202.050 198.600 ;
        RECT 160.950 196.950 163.050 197.400 ;
        RECT 58.950 194.400 75.600 195.600 ;
        RECT 91.950 195.600 94.050 196.050 ;
        RECT 103.950 195.600 106.050 196.050 ;
        RECT 91.950 194.400 106.050 195.600 ;
        RECT 58.950 193.950 61.050 194.400 ;
        RECT 91.950 193.950 94.050 194.400 ;
        RECT 103.950 193.950 106.050 194.400 ;
        RECT 109.950 195.600 112.050 196.050 ;
        RECT 115.950 195.600 118.050 196.050 ;
        RECT 109.950 194.400 118.050 195.600 ;
        RECT 109.950 193.950 112.050 194.400 ;
        RECT 115.950 193.950 118.050 194.400 ;
        RECT 118.950 195.600 121.050 196.050 ;
        RECT 127.950 195.600 130.050 196.050 ;
        RECT 118.950 194.400 130.050 195.600 ;
        RECT 118.950 193.950 121.050 194.400 ;
        RECT 127.950 193.950 130.050 194.400 ;
        RECT 136.950 195.600 139.050 196.050 ;
        RECT 142.950 195.600 145.050 196.050 ;
        RECT 136.950 194.400 145.050 195.600 ;
        RECT 136.950 193.950 139.050 194.400 ;
        RECT 142.950 193.950 145.050 194.400 ;
        RECT 148.950 193.950 151.050 196.050 ;
        RECT 151.950 193.950 154.050 196.050 ;
        RECT 67.950 192.600 70.050 193.050 ;
        RECT 76.950 192.600 79.050 193.050 ;
        RECT 67.950 191.400 79.050 192.600 ;
        RECT 67.950 190.950 70.050 191.400 ;
        RECT 76.950 190.950 79.050 191.400 ;
        RECT 94.950 192.600 97.050 193.050 ;
        RECT 124.950 192.600 127.050 193.050 ;
        RECT 94.950 191.400 127.050 192.600 ;
        RECT 94.950 190.950 97.050 191.400 ;
        RECT 124.950 190.950 127.050 191.400 ;
        RECT 145.950 192.600 148.050 193.050 ;
        RECT 155.400 192.600 156.600 196.950 ;
        RECT 170.400 196.050 171.600 197.400 ;
        RECT 181.950 196.950 184.050 197.400 ;
        RECT 199.950 196.950 202.050 197.400 ;
        RECT 169.950 193.950 172.050 196.050 ;
        RECT 209.400 195.600 210.600 199.950 ;
        RECT 232.950 195.600 235.050 196.050 ;
        RECT 209.400 194.400 235.050 195.600 ;
        RECT 239.400 195.600 240.600 199.950 ;
        RECT 247.950 198.600 250.050 199.050 ;
        RECT 256.950 198.600 259.050 199.050 ;
        RECT 247.950 197.400 259.050 198.600 ;
        RECT 247.950 196.950 250.050 197.400 ;
        RECT 256.950 196.950 259.050 197.400 ;
        RECT 259.950 196.950 262.050 199.050 ;
        RECT 262.950 198.600 265.050 199.050 ;
        RECT 274.950 198.600 277.050 199.050 ;
        RECT 262.950 197.400 277.050 198.600 ;
        RECT 284.400 198.600 285.600 200.400 ;
        RECT 286.950 200.400 298.050 201.600 ;
        RECT 286.950 199.950 289.050 200.400 ;
        RECT 295.950 199.950 298.050 200.400 ;
        RECT 301.950 201.600 304.050 202.050 ;
        RECT 307.950 201.600 310.050 202.050 ;
        RECT 301.950 200.400 310.050 201.600 ;
        RECT 301.950 199.950 304.050 200.400 ;
        RECT 307.950 199.950 310.050 200.400 ;
        RECT 319.950 201.600 322.050 202.050 ;
        RECT 329.400 201.600 330.600 203.400 ;
        RECT 331.950 203.400 370.050 204.600 ;
        RECT 371.400 204.600 372.600 206.400 ;
        RECT 373.950 206.400 405.600 207.600 ;
        RECT 373.950 205.950 376.050 206.400 ;
        RECT 382.950 204.600 385.050 205.050 ;
        RECT 371.400 203.400 385.050 204.600 ;
        RECT 331.950 202.950 334.050 203.400 ;
        RECT 340.950 202.950 343.050 203.400 ;
        RECT 367.950 202.950 370.050 203.400 ;
        RECT 382.950 202.950 385.050 203.400 ;
        RECT 388.950 204.600 391.050 205.050 ;
        RECT 400.950 204.600 403.050 205.050 ;
        RECT 388.950 203.400 403.050 204.600 ;
        RECT 404.400 204.600 405.600 206.400 ;
        RECT 406.950 206.400 424.050 207.600 ;
        RECT 406.950 205.950 409.050 206.400 ;
        RECT 421.950 205.950 424.050 206.400 ;
        RECT 430.950 207.600 433.050 208.050 ;
        RECT 436.950 207.600 439.050 208.050 ;
        RECT 430.950 206.400 439.050 207.600 ;
        RECT 430.950 205.950 433.050 206.400 ;
        RECT 436.950 205.950 439.050 206.400 ;
        RECT 463.950 207.600 466.050 208.050 ;
        RECT 469.950 207.600 472.050 208.050 ;
        RECT 463.950 206.400 472.050 207.600 ;
        RECT 463.950 205.950 466.050 206.400 ;
        RECT 469.950 205.950 472.050 206.400 ;
        RECT 493.950 207.600 496.050 208.050 ;
        RECT 544.950 207.600 547.050 208.050 ;
        RECT 493.950 206.400 547.050 207.600 ;
        RECT 551.400 207.600 552.600 208.950 ;
        RECT 568.950 207.600 571.050 208.050 ;
        RECT 551.400 206.400 571.050 207.600 ;
        RECT 493.950 205.950 496.050 206.400 ;
        RECT 544.950 205.950 547.050 206.400 ;
        RECT 568.950 205.950 571.050 206.400 ;
        RECT 580.950 207.600 583.050 208.050 ;
        RECT 598.950 207.600 601.050 208.050 ;
        RECT 580.950 206.400 601.050 207.600 ;
        RECT 580.950 205.950 583.050 206.400 ;
        RECT 598.950 205.950 601.050 206.400 ;
        RECT 625.950 207.600 628.050 208.050 ;
        RECT 631.950 207.600 634.050 208.050 ;
        RECT 625.950 206.400 634.050 207.600 ;
        RECT 625.950 205.950 628.050 206.400 ;
        RECT 631.950 205.950 634.050 206.400 ;
        RECT 643.950 207.600 646.050 208.050 ;
        RECT 691.950 207.600 694.050 208.050 ;
        RECT 643.950 206.400 694.050 207.600 ;
        RECT 643.950 205.950 646.050 206.400 ;
        RECT 691.950 205.950 694.050 206.400 ;
        RECT 694.950 207.600 697.050 208.050 ;
        RECT 721.950 207.600 724.050 208.050 ;
        RECT 694.950 206.400 724.050 207.600 ;
        RECT 694.950 205.950 697.050 206.400 ;
        RECT 721.950 205.950 724.050 206.400 ;
        RECT 742.950 207.600 745.050 208.050 ;
        RECT 754.950 207.600 757.050 208.050 ;
        RECT 742.950 206.400 757.050 207.600 ;
        RECT 742.950 205.950 745.050 206.400 ;
        RECT 754.950 205.950 757.050 206.400 ;
        RECT 412.950 204.600 415.050 205.050 ;
        RECT 404.400 203.400 415.050 204.600 ;
        RECT 388.950 202.950 391.050 203.400 ;
        RECT 400.950 202.950 403.050 203.400 ;
        RECT 412.950 202.950 415.050 203.400 ;
        RECT 415.950 204.600 418.050 205.050 ;
        RECT 484.950 204.600 487.050 205.050 ;
        RECT 538.950 204.600 541.050 205.050 ;
        RECT 415.950 203.400 487.050 204.600 ;
        RECT 415.950 202.950 418.050 203.400 ;
        RECT 484.950 202.950 487.050 203.400 ;
        RECT 536.400 203.400 541.050 204.600 ;
        RECT 349.950 201.600 352.050 202.050 ;
        RECT 319.950 200.400 327.600 201.600 ;
        RECT 329.400 200.400 352.050 201.600 ;
        RECT 319.950 199.950 322.050 200.400 ;
        RECT 326.400 198.600 327.600 200.400 ;
        RECT 349.950 199.950 352.050 200.400 ;
        RECT 355.950 201.600 358.050 202.050 ;
        RECT 355.950 200.400 369.600 201.600 ;
        RECT 355.950 199.950 358.050 200.400 ;
        RECT 364.950 198.600 367.050 199.050 ;
        RECT 284.400 197.400 288.600 198.600 ;
        RECT 326.400 197.400 351.600 198.600 ;
        RECT 262.950 196.950 265.050 197.400 ;
        RECT 274.950 196.950 277.050 197.400 ;
        RECT 244.950 195.600 247.050 196.050 ;
        RECT 239.400 194.400 247.050 195.600 ;
        RECT 232.950 193.950 235.050 194.400 ;
        RECT 244.950 193.950 247.050 194.400 ;
        RECT 260.400 195.600 261.600 196.950 ;
        RECT 271.950 195.600 274.050 196.050 ;
        RECT 260.400 194.400 274.050 195.600 ;
        RECT 260.400 193.050 261.600 194.400 ;
        RECT 271.950 193.950 274.050 194.400 ;
        RECT 277.950 195.600 280.050 196.050 ;
        RECT 283.950 195.600 286.050 196.050 ;
        RECT 277.950 194.400 286.050 195.600 ;
        RECT 277.950 193.950 280.050 194.400 ;
        RECT 283.950 193.950 286.050 194.400 ;
        RECT 145.950 191.400 156.600 192.600 ;
        RECT 160.950 192.600 163.050 193.050 ;
        RECT 175.950 192.600 178.050 193.050 ;
        RECT 160.950 191.400 178.050 192.600 ;
        RECT 145.950 190.950 148.050 191.400 ;
        RECT 160.950 190.950 163.050 191.400 ;
        RECT 175.950 190.950 178.050 191.400 ;
        RECT 187.950 192.600 190.050 193.050 ;
        RECT 190.950 192.600 193.050 193.050 ;
        RECT 223.950 192.600 226.050 193.050 ;
        RECT 187.950 191.400 226.050 192.600 ;
        RECT 187.950 190.950 190.050 191.400 ;
        RECT 190.950 190.950 193.050 191.400 ;
        RECT 223.950 190.950 226.050 191.400 ;
        RECT 259.950 190.950 262.050 193.050 ;
        RECT 262.950 192.600 265.050 193.050 ;
        RECT 277.950 192.600 280.050 193.050 ;
        RECT 262.950 191.400 280.050 192.600 ;
        RECT 262.950 190.950 265.050 191.400 ;
        RECT 277.950 190.950 280.050 191.400 ;
        RECT 280.950 192.600 283.050 193.050 ;
        RECT 287.400 192.600 288.600 197.400 ;
        RECT 350.400 196.050 351.600 197.400 ;
        RECT 359.400 197.400 367.050 198.600 ;
        RECT 359.400 196.050 360.600 197.400 ;
        RECT 364.950 196.950 367.050 197.400 ;
        RECT 316.950 195.600 319.050 196.050 ;
        RECT 319.950 195.600 322.050 196.050 ;
        RECT 340.950 195.600 343.050 196.050 ;
        RECT 316.950 194.400 343.050 195.600 ;
        RECT 316.950 193.950 319.050 194.400 ;
        RECT 319.950 193.950 322.050 194.400 ;
        RECT 340.950 193.950 343.050 194.400 ;
        RECT 349.950 193.950 352.050 196.050 ;
        RECT 358.950 193.950 361.050 196.050 ;
        RECT 368.400 195.600 369.600 200.400 ;
        RECT 373.950 199.950 376.050 202.050 ;
        RECT 376.950 201.600 379.050 202.050 ;
        RECT 424.950 201.600 427.050 202.050 ;
        RECT 433.950 201.600 436.050 202.050 ;
        RECT 376.950 200.400 423.600 201.600 ;
        RECT 376.950 199.950 379.050 200.400 ;
        RECT 374.400 198.600 375.600 199.950 ;
        RECT 382.950 198.600 385.050 199.050 ;
        RECT 388.950 198.600 391.050 199.050 ;
        RECT 415.950 198.600 418.050 199.050 ;
        RECT 374.400 197.400 381.600 198.600 ;
        RECT 373.950 195.600 376.050 196.050 ;
        RECT 368.400 194.400 376.050 195.600 ;
        RECT 380.400 195.600 381.600 197.400 ;
        RECT 382.950 197.400 391.050 198.600 ;
        RECT 382.950 196.950 385.050 197.400 ;
        RECT 388.950 196.950 391.050 197.400 ;
        RECT 392.400 197.400 418.050 198.600 ;
        RECT 422.400 198.600 423.600 200.400 ;
        RECT 424.950 200.400 436.050 201.600 ;
        RECT 424.950 199.950 427.050 200.400 ;
        RECT 433.950 199.950 436.050 200.400 ;
        RECT 436.950 201.600 439.050 202.050 ;
        RECT 445.950 201.600 448.050 202.050 ;
        RECT 478.950 201.600 481.050 202.050 ;
        RECT 496.950 201.600 499.050 202.050 ;
        RECT 436.950 200.400 448.050 201.600 ;
        RECT 436.950 199.950 439.050 200.400 ;
        RECT 445.950 199.950 448.050 200.400 ;
        RECT 449.400 200.400 481.050 201.600 ;
        RECT 449.400 199.050 450.600 200.400 ;
        RECT 478.950 199.950 481.050 200.400 ;
        RECT 491.400 200.400 499.050 201.600 ;
        RECT 491.400 199.050 492.600 200.400 ;
        RECT 496.950 199.950 499.050 200.400 ;
        RECT 499.950 201.600 502.050 202.050 ;
        RECT 517.950 201.600 520.050 202.050 ;
        RECT 499.950 200.400 516.600 201.600 ;
        RECT 499.950 199.950 502.050 200.400 ;
        RECT 422.400 197.400 441.600 198.600 ;
        RECT 392.400 196.050 393.600 197.400 ;
        RECT 415.950 196.950 418.050 197.400 ;
        RECT 440.400 196.050 441.600 197.400 ;
        RECT 448.950 196.950 451.050 199.050 ;
        RECT 460.950 198.600 463.050 199.050 ;
        RECT 466.950 198.600 469.050 199.050 ;
        RECT 460.950 197.400 469.050 198.600 ;
        RECT 460.950 196.950 463.050 197.400 ;
        RECT 466.950 196.950 469.050 197.400 ;
        RECT 472.950 198.600 475.050 199.050 ;
        RECT 478.950 198.600 481.050 199.050 ;
        RECT 472.950 197.400 481.050 198.600 ;
        RECT 472.950 196.950 475.050 197.400 ;
        RECT 478.950 196.950 481.050 197.400 ;
        RECT 490.950 196.950 493.050 199.050 ;
        RECT 493.950 198.600 496.050 199.050 ;
        RECT 505.950 198.600 508.050 199.050 ;
        RECT 493.950 197.400 508.050 198.600 ;
        RECT 515.400 198.600 516.600 200.400 ;
        RECT 517.950 200.400 534.600 201.600 ;
        RECT 517.950 199.950 520.050 200.400 ;
        RECT 533.400 199.050 534.600 200.400 ;
        RECT 529.950 198.600 532.050 199.050 ;
        RECT 515.400 197.400 532.050 198.600 ;
        RECT 493.950 196.950 496.050 197.400 ;
        RECT 505.950 196.950 508.050 197.400 ;
        RECT 529.950 196.950 532.050 197.400 ;
        RECT 532.950 196.950 535.050 199.050 ;
        RECT 385.950 195.600 388.050 196.050 ;
        RECT 380.400 194.400 388.050 195.600 ;
        RECT 373.950 193.950 376.050 194.400 ;
        RECT 385.950 193.950 388.050 194.400 ;
        RECT 391.950 193.950 394.050 196.050 ;
        RECT 397.950 195.600 400.050 196.050 ;
        RECT 409.950 195.600 412.050 196.050 ;
        RECT 397.950 194.400 412.050 195.600 ;
        RECT 397.950 193.950 400.050 194.400 ;
        RECT 409.950 193.950 412.050 194.400 ;
        RECT 418.950 193.950 421.050 196.050 ;
        RECT 424.950 195.600 427.050 196.050 ;
        RECT 433.950 195.600 436.050 196.050 ;
        RECT 424.950 194.400 436.050 195.600 ;
        RECT 424.950 193.950 427.050 194.400 ;
        RECT 433.950 193.950 436.050 194.400 ;
        RECT 439.950 193.950 442.050 196.050 ;
        RECT 445.950 195.600 448.050 196.050 ;
        RECT 469.950 195.600 472.050 196.050 ;
        RECT 445.950 194.400 472.050 195.600 ;
        RECT 445.950 193.950 448.050 194.400 ;
        RECT 469.950 193.950 472.050 194.400 ;
        RECT 475.950 195.600 478.050 196.050 ;
        RECT 481.950 195.600 484.050 196.050 ;
        RECT 511.950 195.600 514.050 196.050 ;
        RECT 475.950 194.400 514.050 195.600 ;
        RECT 475.950 193.950 478.050 194.400 ;
        RECT 481.950 193.950 484.050 194.400 ;
        RECT 511.950 193.950 514.050 194.400 ;
        RECT 532.950 195.600 535.050 196.050 ;
        RECT 536.400 195.600 537.600 203.400 ;
        RECT 538.950 202.950 541.050 203.400 ;
        RECT 541.950 204.600 544.050 205.050 ;
        RECT 589.950 204.600 592.050 205.050 ;
        RECT 541.950 203.400 592.050 204.600 ;
        RECT 541.950 202.950 544.050 203.400 ;
        RECT 589.950 202.950 592.050 203.400 ;
        RECT 607.950 204.600 610.050 205.050 ;
        RECT 613.950 204.600 616.050 205.050 ;
        RECT 607.950 203.400 616.050 204.600 ;
        RECT 607.950 202.950 610.050 203.400 ;
        RECT 613.950 202.950 616.050 203.400 ;
        RECT 619.950 204.600 622.050 205.050 ;
        RECT 619.950 203.400 633.600 204.600 ;
        RECT 619.950 202.950 622.050 203.400 ;
        RECT 550.950 199.950 553.050 202.050 ;
        RECT 556.950 201.600 559.050 202.050 ;
        RECT 565.950 201.600 568.050 202.050 ;
        RECT 556.950 200.400 568.050 201.600 ;
        RECT 556.950 199.950 559.050 200.400 ;
        RECT 565.950 199.950 568.050 200.400 ;
        RECT 571.950 201.600 574.050 202.050 ;
        RECT 577.950 201.600 580.050 202.050 ;
        RECT 571.950 200.400 580.050 201.600 ;
        RECT 571.950 199.950 574.050 200.400 ;
        RECT 577.950 199.950 580.050 200.400 ;
        RECT 583.950 201.600 586.050 202.050 ;
        RECT 595.950 201.600 598.050 202.050 ;
        RECT 601.950 201.600 604.050 202.050 ;
        RECT 583.950 200.400 604.050 201.600 ;
        RECT 583.950 199.950 586.050 200.400 ;
        RECT 595.950 199.950 598.050 200.400 ;
        RECT 601.950 199.950 604.050 200.400 ;
        RECT 604.950 199.950 607.050 202.050 ;
        RECT 610.950 199.950 613.050 202.050 ;
        RECT 538.950 198.600 541.050 199.050 ;
        RECT 544.950 198.600 547.050 199.050 ;
        RECT 538.950 197.400 547.050 198.600 ;
        RECT 538.950 196.950 541.050 197.400 ;
        RECT 544.950 196.950 547.050 197.400 ;
        RECT 532.950 194.400 537.600 195.600 ;
        RECT 551.400 195.600 552.600 199.950 ;
        RECT 553.950 198.600 556.050 199.050 ;
        RECT 605.400 198.600 606.600 199.950 ;
        RECT 553.950 197.400 606.600 198.600 ;
        RECT 553.950 196.950 556.050 197.400 ;
        RECT 559.950 195.600 562.050 196.050 ;
        RECT 551.400 194.400 562.050 195.600 ;
        RECT 532.950 193.950 535.050 194.400 ;
        RECT 559.950 193.950 562.050 194.400 ;
        RECT 586.950 195.600 589.050 196.050 ;
        RECT 598.950 195.600 601.050 196.050 ;
        RECT 586.950 194.400 601.050 195.600 ;
        RECT 611.400 195.600 612.600 199.950 ;
        RECT 619.950 198.600 622.050 199.050 ;
        RECT 628.950 198.600 631.050 199.050 ;
        RECT 619.950 197.400 631.050 198.600 ;
        RECT 632.400 198.600 633.600 203.400 ;
        RECT 637.950 202.950 640.050 205.050 ;
        RECT 646.950 204.600 649.050 205.050 ;
        RECT 664.950 204.600 667.050 205.050 ;
        RECT 730.950 204.600 733.050 205.050 ;
        RECT 646.950 203.400 651.600 204.600 ;
        RECT 646.950 202.950 649.050 203.400 ;
        RECT 634.950 201.600 637.050 202.050 ;
        RECT 638.400 201.600 639.600 202.950 ;
        RECT 650.400 202.050 651.600 203.400 ;
        RECT 664.950 203.400 684.600 204.600 ;
        RECT 664.950 202.950 667.050 203.400 ;
        RECT 683.400 202.050 684.600 203.400 ;
        RECT 728.400 203.400 733.050 204.600 ;
        RECT 634.950 200.400 639.600 201.600 ;
        RECT 640.950 201.600 643.050 202.050 ;
        RECT 649.950 201.600 652.050 202.050 ;
        RECT 640.950 200.400 652.050 201.600 ;
        RECT 634.950 199.950 637.050 200.400 ;
        RECT 640.950 199.950 643.050 200.400 ;
        RECT 649.950 199.950 652.050 200.400 ;
        RECT 673.950 199.950 676.050 202.050 ;
        RECT 682.950 199.950 685.050 202.050 ;
        RECT 688.950 201.600 691.050 202.050 ;
        RECT 694.950 201.600 697.050 202.050 ;
        RECT 688.950 200.400 697.050 201.600 ;
        RECT 688.950 199.950 691.050 200.400 ;
        RECT 694.950 199.950 697.050 200.400 ;
        RECT 715.950 199.950 718.050 202.050 ;
        RECT 649.950 198.600 652.050 199.050 ;
        RECT 632.400 197.400 652.050 198.600 ;
        RECT 619.950 196.950 622.050 197.400 ;
        RECT 628.950 196.950 631.050 197.400 ;
        RECT 649.950 196.950 652.050 197.400 ;
        RECT 664.950 196.950 667.050 199.050 ;
        RECT 667.950 196.950 670.050 199.050 ;
        RECT 670.950 196.950 673.050 199.050 ;
        RECT 646.950 195.600 649.050 196.050 ;
        RECT 611.400 194.400 649.050 195.600 ;
        RECT 586.950 193.950 589.050 194.400 ;
        RECT 598.950 193.950 601.050 194.400 ;
        RECT 646.950 193.950 649.050 194.400 ;
        RECT 655.950 195.600 658.050 196.050 ;
        RECT 665.400 195.600 666.600 196.950 ;
        RECT 655.950 194.400 666.600 195.600 ;
        RECT 655.950 193.950 658.050 194.400 ;
        RECT 307.950 192.600 310.050 193.050 ;
        RECT 319.950 192.600 322.050 193.050 ;
        RECT 280.950 191.400 288.600 192.600 ;
        RECT 290.400 191.400 322.050 192.600 ;
        RECT 280.950 190.950 283.050 191.400 ;
        RECT 64.950 189.600 67.050 190.050 ;
        RECT 70.950 189.600 73.050 190.050 ;
        RECT 13.950 188.400 73.050 189.600 ;
        RECT 13.950 187.950 16.050 188.400 ;
        RECT 64.950 187.950 67.050 188.400 ;
        RECT 70.950 187.950 73.050 188.400 ;
        RECT 73.950 189.600 76.050 190.050 ;
        RECT 112.950 189.600 115.050 190.050 ;
        RECT 73.950 188.400 115.050 189.600 ;
        RECT 73.950 187.950 76.050 188.400 ;
        RECT 112.950 187.950 115.050 188.400 ;
        RECT 142.950 189.600 145.050 190.050 ;
        RECT 157.950 189.600 160.050 190.050 ;
        RECT 181.950 189.600 184.050 190.050 ;
        RECT 142.950 188.400 160.050 189.600 ;
        RECT 142.950 187.950 145.050 188.400 ;
        RECT 157.950 187.950 160.050 188.400 ;
        RECT 173.400 188.400 184.050 189.600 ;
        RECT 1.950 186.600 4.050 187.050 ;
        RECT 16.950 186.600 19.050 187.050 ;
        RECT 1.950 185.400 19.050 186.600 ;
        RECT 1.950 184.950 4.050 185.400 ;
        RECT 16.950 184.950 19.050 185.400 ;
        RECT 22.950 186.600 25.050 187.050 ;
        RECT 40.950 186.600 43.050 187.050 ;
        RECT 85.950 186.600 88.050 187.050 ;
        RECT 22.950 185.400 43.050 186.600 ;
        RECT 22.950 184.950 25.050 185.400 ;
        RECT 40.950 184.950 43.050 185.400 ;
        RECT 44.400 185.400 88.050 186.600 ;
        RECT 7.950 183.600 10.050 184.050 ;
        RECT 16.950 183.600 19.050 184.050 ;
        RECT 44.400 183.600 45.600 185.400 ;
        RECT 85.950 184.950 88.050 185.400 ;
        RECT 154.950 186.600 157.050 187.050 ;
        RECT 173.400 186.600 174.600 188.400 ;
        RECT 181.950 187.950 184.050 188.400 ;
        RECT 244.950 189.600 247.050 190.050 ;
        RECT 290.400 189.600 291.600 191.400 ;
        RECT 307.950 190.950 310.050 191.400 ;
        RECT 319.950 190.950 322.050 191.400 ;
        RECT 343.950 192.600 346.050 193.050 ;
        RECT 355.950 192.600 358.050 193.050 ;
        RECT 343.950 191.400 358.050 192.600 ;
        RECT 343.950 190.950 346.050 191.400 ;
        RECT 355.950 190.950 358.050 191.400 ;
        RECT 376.950 192.600 379.050 193.050 ;
        RECT 382.950 192.600 385.050 193.050 ;
        RECT 376.950 191.400 385.050 192.600 ;
        RECT 419.400 192.600 420.600 193.950 ;
        RECT 460.950 192.600 463.050 193.050 ;
        RECT 419.400 191.400 463.050 192.600 ;
        RECT 376.950 190.950 379.050 191.400 ;
        RECT 382.950 190.950 385.050 191.400 ;
        RECT 460.950 190.950 463.050 191.400 ;
        RECT 466.950 192.600 469.050 193.050 ;
        RECT 496.950 192.600 499.050 193.050 ;
        RECT 514.950 192.600 517.050 193.050 ;
        RECT 466.950 191.400 517.050 192.600 ;
        RECT 466.950 190.950 469.050 191.400 ;
        RECT 496.950 190.950 499.050 191.400 ;
        RECT 514.950 190.950 517.050 191.400 ;
        RECT 523.950 192.600 526.050 193.050 ;
        RECT 529.950 192.600 532.050 193.050 ;
        RECT 523.950 191.400 532.050 192.600 ;
        RECT 523.950 190.950 526.050 191.400 ;
        RECT 529.950 190.950 532.050 191.400 ;
        RECT 580.950 192.600 583.050 193.050 ;
        RECT 610.950 192.600 613.050 193.050 ;
        RECT 580.950 191.400 613.050 192.600 ;
        RECT 580.950 190.950 583.050 191.400 ;
        RECT 610.950 190.950 613.050 191.400 ;
        RECT 625.950 192.600 628.050 193.050 ;
        RECT 628.950 192.600 631.050 193.050 ;
        RECT 637.950 192.600 640.050 193.050 ;
        RECT 625.950 191.400 640.050 192.600 ;
        RECT 625.950 190.950 628.050 191.400 ;
        RECT 628.950 190.950 631.050 191.400 ;
        RECT 637.950 190.950 640.050 191.400 ;
        RECT 643.950 192.600 646.050 193.050 ;
        RECT 664.950 192.600 667.050 193.050 ;
        RECT 643.950 191.400 667.050 192.600 ;
        RECT 643.950 190.950 646.050 191.400 ;
        RECT 664.950 190.950 667.050 191.400 ;
        RECT 244.950 188.400 291.600 189.600 ;
        RECT 304.950 189.600 307.050 190.050 ;
        RECT 334.950 189.600 337.050 190.050 ;
        RECT 304.950 188.400 337.050 189.600 ;
        RECT 244.950 187.950 247.050 188.400 ;
        RECT 304.950 187.950 307.050 188.400 ;
        RECT 334.950 187.950 337.050 188.400 ;
        RECT 349.950 189.600 352.050 190.050 ;
        RECT 424.950 189.600 427.050 190.050 ;
        RECT 430.950 189.600 433.050 190.050 ;
        RECT 475.950 189.600 478.050 190.050 ;
        RECT 349.950 188.400 423.600 189.600 ;
        RECT 349.950 187.950 352.050 188.400 ;
        RECT 154.950 185.400 174.600 186.600 ;
        RECT 178.950 186.600 181.050 187.050 ;
        RECT 211.950 186.600 214.050 187.050 ;
        RECT 247.950 186.600 250.050 187.050 ;
        RECT 262.950 186.600 265.050 187.050 ;
        RECT 178.950 185.400 214.050 186.600 ;
        RECT 154.950 184.950 157.050 185.400 ;
        RECT 178.950 184.950 181.050 185.400 ;
        RECT 211.950 184.950 214.050 185.400 ;
        RECT 215.400 185.400 265.050 186.600 ;
        RECT 7.950 182.400 45.600 183.600 ;
        RECT 52.950 183.600 55.050 184.050 ;
        RECT 79.950 183.600 82.050 184.050 ;
        RECT 52.950 182.400 82.050 183.600 ;
        RECT 7.950 181.950 10.050 182.400 ;
        RECT 16.950 181.950 19.050 182.400 ;
        RECT 52.950 181.950 55.050 182.400 ;
        RECT 79.950 181.950 82.050 182.400 ;
        RECT 85.950 183.600 88.050 184.050 ;
        RECT 97.950 183.600 100.050 184.050 ;
        RECT 184.950 183.600 187.050 184.050 ;
        RECT 85.950 182.400 187.050 183.600 ;
        RECT 85.950 181.950 88.050 182.400 ;
        RECT 97.950 181.950 100.050 182.400 ;
        RECT 184.950 181.950 187.050 182.400 ;
        RECT 190.950 183.600 193.050 184.050 ;
        RECT 205.950 183.600 208.050 184.050 ;
        RECT 215.400 183.600 216.600 185.400 ;
        RECT 247.950 184.950 250.050 185.400 ;
        RECT 262.950 184.950 265.050 185.400 ;
        RECT 268.950 186.600 271.050 187.050 ;
        RECT 283.950 186.600 286.050 187.050 ;
        RECT 340.950 186.600 343.050 187.050 ;
        RECT 268.950 185.400 343.050 186.600 ;
        RECT 268.950 184.950 271.050 185.400 ;
        RECT 283.950 184.950 286.050 185.400 ;
        RECT 340.950 184.950 343.050 185.400 ;
        RECT 364.950 186.600 367.050 187.050 ;
        RECT 394.950 186.600 397.050 187.050 ;
        RECT 364.950 185.400 397.050 186.600 ;
        RECT 422.400 186.600 423.600 188.400 ;
        RECT 424.950 188.400 433.050 189.600 ;
        RECT 424.950 187.950 427.050 188.400 ;
        RECT 430.950 187.950 433.050 188.400 ;
        RECT 455.400 188.400 478.050 189.600 ;
        RECT 455.400 186.600 456.600 188.400 ;
        RECT 475.950 187.950 478.050 188.400 ;
        RECT 490.950 189.600 493.050 190.050 ;
        RECT 574.950 189.600 577.050 190.050 ;
        RECT 592.950 189.600 595.050 190.050 ;
        RECT 490.950 188.400 595.050 189.600 ;
        RECT 490.950 187.950 493.050 188.400 ;
        RECT 574.950 187.950 577.050 188.400 ;
        RECT 592.950 187.950 595.050 188.400 ;
        RECT 604.950 189.600 607.050 190.050 ;
        RECT 625.950 189.600 628.050 190.050 ;
        RECT 652.950 189.600 655.050 190.050 ;
        RECT 604.950 188.400 655.050 189.600 ;
        RECT 668.400 189.600 669.600 196.950 ;
        RECT 671.400 192.600 672.600 196.950 ;
        RECT 674.400 196.050 675.600 199.950 ;
        RECT 682.950 198.600 685.050 199.050 ;
        RECT 697.950 198.600 700.050 199.050 ;
        RECT 682.950 197.400 700.050 198.600 ;
        RECT 682.950 196.950 685.050 197.400 ;
        RECT 697.950 196.950 700.050 197.400 ;
        RECT 673.950 193.950 676.050 196.050 ;
        RECT 676.950 195.600 679.050 196.050 ;
        RECT 688.950 195.600 691.050 196.050 ;
        RECT 676.950 194.400 691.050 195.600 ;
        RECT 676.950 193.950 679.050 194.400 ;
        RECT 688.950 193.950 691.050 194.400 ;
        RECT 685.950 192.600 688.050 193.050 ;
        RECT 671.400 191.400 688.050 192.600 ;
        RECT 685.950 190.950 688.050 191.400 ;
        RECT 712.950 192.600 715.050 193.050 ;
        RECT 716.400 192.600 717.600 199.950 ;
        RECT 728.400 195.600 729.600 203.400 ;
        RECT 730.950 202.950 733.050 203.400 ;
        RECT 739.950 202.950 742.050 205.050 ;
        RECT 745.950 204.600 748.050 205.050 ;
        RECT 763.950 204.600 766.050 205.050 ;
        RECT 745.950 203.400 750.600 204.600 ;
        RECT 745.950 202.950 748.050 203.400 ;
        RECT 740.400 201.600 741.600 202.950 ;
        RECT 740.400 200.400 747.600 201.600 ;
        RECT 730.950 198.600 733.050 199.050 ;
        RECT 742.950 198.600 745.050 199.050 ;
        RECT 730.950 197.400 745.050 198.600 ;
        RECT 730.950 196.950 733.050 197.400 ;
        RECT 742.950 196.950 745.050 197.400 ;
        RECT 733.950 195.600 736.050 196.050 ;
        RECT 746.400 195.600 747.600 200.400 ;
        RECT 749.400 196.050 750.600 203.400 ;
        RECT 763.950 203.400 771.600 204.600 ;
        RECT 763.950 202.950 766.050 203.400 ;
        RECT 766.950 201.600 769.050 202.050 ;
        RECT 761.400 200.400 769.050 201.600 ;
        RECT 728.400 194.400 736.050 195.600 ;
        RECT 733.950 193.950 736.050 194.400 ;
        RECT 740.400 194.400 747.600 195.600 ;
        RECT 712.950 191.400 717.600 192.600 ;
        RECT 721.950 192.600 724.050 193.050 ;
        RECT 730.950 192.600 733.050 193.050 ;
        RECT 721.950 191.400 733.050 192.600 ;
        RECT 712.950 190.950 715.050 191.400 ;
        RECT 721.950 190.950 724.050 191.400 ;
        RECT 730.950 190.950 733.050 191.400 ;
        RECT 670.950 189.600 673.050 190.050 ;
        RECT 668.400 188.400 673.050 189.600 ;
        RECT 604.950 187.950 607.050 188.400 ;
        RECT 625.950 187.950 628.050 188.400 ;
        RECT 652.950 187.950 655.050 188.400 ;
        RECT 670.950 187.950 673.050 188.400 ;
        RECT 676.950 189.600 679.050 190.050 ;
        RECT 721.950 189.600 724.050 190.050 ;
        RECT 676.950 188.400 724.050 189.600 ;
        RECT 676.950 187.950 679.050 188.400 ;
        RECT 721.950 187.950 724.050 188.400 ;
        RECT 730.950 189.600 733.050 190.050 ;
        RECT 740.400 189.600 741.600 194.400 ;
        RECT 748.950 193.950 751.050 196.050 ;
        RECT 742.950 192.600 745.050 193.050 ;
        RECT 754.950 192.600 757.050 193.050 ;
        RECT 742.950 191.400 757.050 192.600 ;
        RECT 742.950 190.950 745.050 191.400 ;
        RECT 754.950 190.950 757.050 191.400 ;
        RECT 761.400 190.050 762.600 200.400 ;
        RECT 766.950 199.950 769.050 200.400 ;
        RECT 730.950 188.400 741.600 189.600 ;
        RECT 745.950 189.600 748.050 190.050 ;
        RECT 757.950 189.600 760.050 190.050 ;
        RECT 745.950 188.400 760.050 189.600 ;
        RECT 730.950 187.950 733.050 188.400 ;
        RECT 745.950 187.950 748.050 188.400 ;
        RECT 757.950 187.950 760.050 188.400 ;
        RECT 760.950 187.950 763.050 190.050 ;
        RECT 422.400 185.400 456.600 186.600 ;
        RECT 568.950 186.600 571.050 187.050 ;
        RECT 643.950 186.600 646.050 187.050 ;
        RECT 568.950 185.400 646.050 186.600 ;
        RECT 364.950 184.950 367.050 185.400 ;
        RECT 394.950 184.950 397.050 185.400 ;
        RECT 568.950 184.950 571.050 185.400 ;
        RECT 643.950 184.950 646.050 185.400 ;
        RECT 646.950 186.600 649.050 187.050 ;
        RECT 652.950 186.600 655.050 187.050 ;
        RECT 646.950 185.400 655.050 186.600 ;
        RECT 646.950 184.950 649.050 185.400 ;
        RECT 652.950 184.950 655.050 185.400 ;
        RECT 664.950 186.600 667.050 187.050 ;
        RECT 697.950 186.600 700.050 187.050 ;
        RECT 664.950 185.400 700.050 186.600 ;
        RECT 664.950 184.950 667.050 185.400 ;
        RECT 697.950 184.950 700.050 185.400 ;
        RECT 706.950 186.600 709.050 187.050 ;
        RECT 712.950 186.600 715.050 187.050 ;
        RECT 766.950 186.600 769.050 187.050 ;
        RECT 706.950 185.400 769.050 186.600 ;
        RECT 706.950 184.950 709.050 185.400 ;
        RECT 712.950 184.950 715.050 185.400 ;
        RECT 766.950 184.950 769.050 185.400 ;
        RECT 190.950 182.400 216.600 183.600 ;
        RECT 232.950 183.600 235.050 184.050 ;
        RECT 271.950 183.600 274.050 184.050 ;
        RECT 232.950 182.400 274.050 183.600 ;
        RECT 190.950 181.950 193.050 182.400 ;
        RECT 205.950 181.950 208.050 182.400 ;
        RECT 232.950 181.950 235.050 182.400 ;
        RECT 271.950 181.950 274.050 182.400 ;
        RECT 274.950 183.600 277.050 184.050 ;
        RECT 310.950 183.600 313.050 184.050 ;
        RECT 274.950 182.400 313.050 183.600 ;
        RECT 274.950 181.950 277.050 182.400 ;
        RECT 310.950 181.950 313.050 182.400 ;
        RECT 322.950 183.600 325.050 184.050 ;
        RECT 352.950 183.600 355.050 184.050 ;
        RECT 322.950 182.400 355.050 183.600 ;
        RECT 322.950 181.950 325.050 182.400 ;
        RECT 352.950 181.950 355.050 182.400 ;
        RECT 379.950 183.600 382.050 184.050 ;
        RECT 430.950 183.600 433.050 184.050 ;
        RECT 379.950 182.400 433.050 183.600 ;
        RECT 379.950 181.950 382.050 182.400 ;
        RECT 430.950 181.950 433.050 182.400 ;
        RECT 556.950 183.600 559.050 184.050 ;
        RECT 601.950 183.600 604.050 184.050 ;
        RECT 556.950 182.400 604.050 183.600 ;
        RECT 556.950 181.950 559.050 182.400 ;
        RECT 601.950 181.950 604.050 182.400 ;
        RECT 616.950 183.600 619.050 184.050 ;
        RECT 655.950 183.600 658.050 184.050 ;
        RECT 616.950 182.400 658.050 183.600 ;
        RECT 616.950 181.950 619.050 182.400 ;
        RECT 655.950 181.950 658.050 182.400 ;
        RECT 667.950 183.600 670.050 184.050 ;
        RECT 679.950 183.600 682.050 184.050 ;
        RECT 685.950 183.600 688.050 184.050 ;
        RECT 667.950 182.400 688.050 183.600 ;
        RECT 667.950 181.950 670.050 182.400 ;
        RECT 679.950 181.950 682.050 182.400 ;
        RECT 685.950 181.950 688.050 182.400 ;
        RECT 688.950 183.600 691.050 184.050 ;
        RECT 763.950 183.600 766.050 184.050 ;
        RECT 688.950 182.400 766.050 183.600 ;
        RECT 688.950 181.950 691.050 182.400 ;
        RECT 763.950 181.950 766.050 182.400 ;
        RECT 766.950 183.600 769.050 184.050 ;
        RECT 770.400 183.600 771.600 203.400 ;
        RECT 766.950 182.400 771.600 183.600 ;
        RECT 766.950 181.950 769.050 182.400 ;
        RECT 160.950 180.600 163.050 181.050 ;
        RECT 172.950 180.600 175.050 181.050 ;
        RECT 187.950 180.600 190.050 181.050 ;
        RECT 160.950 179.400 190.050 180.600 ;
        RECT 160.950 178.950 163.050 179.400 ;
        RECT 172.950 178.950 175.050 179.400 ;
        RECT 187.950 178.950 190.050 179.400 ;
        RECT 196.950 180.600 199.050 181.050 ;
        RECT 238.950 180.600 241.050 181.050 ;
        RECT 196.950 179.400 241.050 180.600 ;
        RECT 196.950 178.950 199.050 179.400 ;
        RECT 238.950 178.950 241.050 179.400 ;
        RECT 241.950 180.600 244.050 181.050 ;
        RECT 265.950 180.600 268.050 181.050 ;
        RECT 241.950 179.400 268.050 180.600 ;
        RECT 241.950 178.950 244.050 179.400 ;
        RECT 265.950 178.950 268.050 179.400 ;
        RECT 289.950 180.600 292.050 181.050 ;
        RECT 301.950 180.600 304.050 181.050 ;
        RECT 307.950 180.600 310.050 181.050 ;
        RECT 289.950 179.400 310.050 180.600 ;
        RECT 289.950 178.950 292.050 179.400 ;
        RECT 301.950 178.950 304.050 179.400 ;
        RECT 307.950 178.950 310.050 179.400 ;
        RECT 340.950 180.600 343.050 181.050 ;
        RECT 400.950 180.600 403.050 181.050 ;
        RECT 499.950 180.600 502.050 181.050 ;
        RECT 340.950 179.400 502.050 180.600 ;
        RECT 340.950 178.950 343.050 179.400 ;
        RECT 400.950 178.950 403.050 179.400 ;
        RECT 499.950 178.950 502.050 179.400 ;
        RECT 517.950 180.600 520.050 181.050 ;
        RECT 571.950 180.600 574.050 181.050 ;
        RECT 517.950 179.400 574.050 180.600 ;
        RECT 517.950 178.950 520.050 179.400 ;
        RECT 571.950 178.950 574.050 179.400 ;
        RECT 589.950 180.600 592.050 181.050 ;
        RECT 637.950 180.600 640.050 181.050 ;
        RECT 589.950 179.400 640.050 180.600 ;
        RECT 589.950 178.950 592.050 179.400 ;
        RECT 637.950 178.950 640.050 179.400 ;
        RECT 649.950 180.600 652.050 181.050 ;
        RECT 676.950 180.600 679.050 181.050 ;
        RECT 649.950 179.400 679.050 180.600 ;
        RECT 649.950 178.950 652.050 179.400 ;
        RECT 676.950 178.950 679.050 179.400 ;
        RECT 697.950 180.600 700.050 181.050 ;
        RECT 745.950 180.600 748.050 181.050 ;
        RECT 697.950 179.400 748.050 180.600 ;
        RECT 697.950 178.950 700.050 179.400 ;
        RECT 745.950 178.950 748.050 179.400 ;
        RECT 751.950 180.600 754.050 181.050 ;
        RECT 760.950 180.600 763.050 181.050 ;
        RECT 751.950 179.400 763.050 180.600 ;
        RECT 751.950 178.950 754.050 179.400 ;
        RECT 760.950 178.950 763.050 179.400 ;
        RECT 4.950 177.600 7.050 178.050 ;
        RECT 58.950 177.600 61.050 178.050 ;
        RECT 4.950 176.400 61.050 177.600 ;
        RECT 4.950 175.950 7.050 176.400 ;
        RECT 58.950 175.950 61.050 176.400 ;
        RECT 82.950 177.600 85.050 178.050 ;
        RECT 121.950 177.600 124.050 178.050 ;
        RECT 82.950 176.400 124.050 177.600 ;
        RECT 82.950 175.950 85.050 176.400 ;
        RECT 121.950 175.950 124.050 176.400 ;
        RECT 127.950 177.600 130.050 178.050 ;
        RECT 151.950 177.600 154.050 178.050 ;
        RECT 169.950 177.600 172.050 178.050 ;
        RECT 127.950 176.400 172.050 177.600 ;
        RECT 127.950 175.950 130.050 176.400 ;
        RECT 151.950 175.950 154.050 176.400 ;
        RECT 169.950 175.950 172.050 176.400 ;
        RECT 178.950 177.600 181.050 178.050 ;
        RECT 193.950 177.600 196.050 178.050 ;
        RECT 178.950 176.400 196.050 177.600 ;
        RECT 178.950 175.950 181.050 176.400 ;
        RECT 193.950 175.950 196.050 176.400 ;
        RECT 211.950 177.600 214.050 178.050 ;
        RECT 217.950 177.600 220.050 178.050 ;
        RECT 238.950 177.600 241.050 178.050 ;
        RECT 211.950 176.400 241.050 177.600 ;
        RECT 211.950 175.950 214.050 176.400 ;
        RECT 217.950 175.950 220.050 176.400 ;
        RECT 238.950 175.950 241.050 176.400 ;
        RECT 244.950 177.600 247.050 178.050 ;
        RECT 292.950 177.600 295.050 178.050 ;
        RECT 244.950 176.400 295.050 177.600 ;
        RECT 244.950 175.950 247.050 176.400 ;
        RECT 292.950 175.950 295.050 176.400 ;
        RECT 316.950 177.600 319.050 178.050 ;
        RECT 349.950 177.600 352.050 178.050 ;
        RECT 316.950 176.400 352.050 177.600 ;
        RECT 316.950 175.950 319.050 176.400 ;
        RECT 349.950 175.950 352.050 176.400 ;
        RECT 367.950 177.600 370.050 178.050 ;
        RECT 403.950 177.600 406.050 178.050 ;
        RECT 367.950 176.400 406.050 177.600 ;
        RECT 367.950 175.950 370.050 176.400 ;
        RECT 403.950 175.950 406.050 176.400 ;
        RECT 427.950 177.600 430.050 178.050 ;
        RECT 472.950 177.600 475.050 178.050 ;
        RECT 478.950 177.600 481.050 178.050 ;
        RECT 427.950 176.400 481.050 177.600 ;
        RECT 427.950 175.950 430.050 176.400 ;
        RECT 472.950 175.950 475.050 176.400 ;
        RECT 478.950 175.950 481.050 176.400 ;
        RECT 502.950 177.600 505.050 178.050 ;
        RECT 535.950 177.600 538.050 178.050 ;
        RECT 502.950 176.400 538.050 177.600 ;
        RECT 502.950 175.950 505.050 176.400 ;
        RECT 535.950 175.950 538.050 176.400 ;
        RECT 565.950 177.600 568.050 178.050 ;
        RECT 586.950 177.600 589.050 178.050 ;
        RECT 565.950 176.400 589.050 177.600 ;
        RECT 565.950 175.950 568.050 176.400 ;
        RECT 586.950 175.950 589.050 176.400 ;
        RECT 589.950 177.600 592.050 178.050 ;
        RECT 598.950 177.600 601.050 178.050 ;
        RECT 619.950 177.600 622.050 178.050 ;
        RECT 589.950 176.400 622.050 177.600 ;
        RECT 589.950 175.950 592.050 176.400 ;
        RECT 598.950 175.950 601.050 176.400 ;
        RECT 619.950 175.950 622.050 176.400 ;
        RECT 643.950 177.600 646.050 178.050 ;
        RECT 658.950 177.600 661.050 178.050 ;
        RECT 643.950 176.400 661.050 177.600 ;
        RECT 643.950 175.950 646.050 176.400 ;
        RECT 658.950 175.950 661.050 176.400 ;
        RECT 682.950 177.600 685.050 178.050 ;
        RECT 703.950 177.600 706.050 178.050 ;
        RECT 724.950 177.600 727.050 178.050 ;
        RECT 682.950 176.400 727.050 177.600 ;
        RECT 682.950 175.950 685.050 176.400 ;
        RECT 703.950 175.950 706.050 176.400 ;
        RECT 724.950 175.950 727.050 176.400 ;
        RECT 730.950 177.600 733.050 178.050 ;
        RECT 754.950 177.600 757.050 178.050 ;
        RECT 730.950 176.400 757.050 177.600 ;
        RECT 730.950 175.950 733.050 176.400 ;
        RECT 754.950 175.950 757.050 176.400 ;
        RECT 49.950 174.600 52.050 175.050 ;
        RECT 58.950 174.600 61.050 175.050 ;
        RECT 145.950 174.600 148.050 175.050 ;
        RECT 49.950 173.400 148.050 174.600 ;
        RECT 49.950 172.950 52.050 173.400 ;
        RECT 58.950 172.950 61.050 173.400 ;
        RECT 145.950 172.950 148.050 173.400 ;
        RECT 181.950 174.600 184.050 175.050 ;
        RECT 280.950 174.600 283.050 175.050 ;
        RECT 181.950 173.400 283.050 174.600 ;
        RECT 181.950 172.950 184.050 173.400 ;
        RECT 280.950 172.950 283.050 173.400 ;
        RECT 289.950 174.600 292.050 175.050 ;
        RECT 328.950 174.600 331.050 175.050 ;
        RECT 289.950 173.400 331.050 174.600 ;
        RECT 289.950 172.950 292.050 173.400 ;
        RECT 328.950 172.950 331.050 173.400 ;
        RECT 346.950 174.600 349.050 175.050 ;
        RECT 355.950 174.600 358.050 175.050 ;
        RECT 346.950 173.400 358.050 174.600 ;
        RECT 346.950 172.950 349.050 173.400 ;
        RECT 355.950 172.950 358.050 173.400 ;
        RECT 361.950 174.600 364.050 175.050 ;
        RECT 385.950 174.600 388.050 175.050 ;
        RECT 361.950 173.400 388.050 174.600 ;
        RECT 361.950 172.950 364.050 173.400 ;
        RECT 385.950 172.950 388.050 173.400 ;
        RECT 388.950 174.600 391.050 175.050 ;
        RECT 391.950 174.600 394.050 175.050 ;
        RECT 415.950 174.600 418.050 175.050 ;
        RECT 427.950 174.600 430.050 175.050 ;
        RECT 559.950 174.600 562.050 175.050 ;
        RECT 592.950 174.600 595.050 175.050 ;
        RECT 388.950 173.400 430.050 174.600 ;
        RECT 388.950 172.950 391.050 173.400 ;
        RECT 391.950 172.950 394.050 173.400 ;
        RECT 415.950 172.950 418.050 173.400 ;
        RECT 427.950 172.950 430.050 173.400 ;
        RECT 434.400 173.400 595.050 174.600 ;
        RECT 136.950 171.600 139.050 172.050 ;
        RECT 163.950 171.600 166.050 172.050 ;
        RECT 136.950 170.400 166.050 171.600 ;
        RECT 136.950 169.950 139.050 170.400 ;
        RECT 163.950 169.950 166.050 170.400 ;
        RECT 181.950 171.600 184.050 172.050 ;
        RECT 211.950 171.600 214.050 172.050 ;
        RECT 181.950 170.400 214.050 171.600 ;
        RECT 181.950 169.950 184.050 170.400 ;
        RECT 211.950 169.950 214.050 170.400 ;
        RECT 217.950 171.600 220.050 172.050 ;
        RECT 235.950 171.600 238.050 172.050 ;
        RECT 217.950 170.400 238.050 171.600 ;
        RECT 217.950 169.950 220.050 170.400 ;
        RECT 235.950 169.950 238.050 170.400 ;
        RECT 250.950 171.600 253.050 172.050 ;
        RECT 256.950 171.600 259.050 172.050 ;
        RECT 250.950 170.400 259.050 171.600 ;
        RECT 250.950 169.950 253.050 170.400 ;
        RECT 256.950 169.950 259.050 170.400 ;
        RECT 259.950 171.600 262.050 172.050 ;
        RECT 265.950 171.600 268.050 172.050 ;
        RECT 259.950 170.400 268.050 171.600 ;
        RECT 259.950 169.950 262.050 170.400 ;
        RECT 265.950 169.950 268.050 170.400 ;
        RECT 298.950 171.600 301.050 172.050 ;
        RECT 316.950 171.600 319.050 172.050 ;
        RECT 298.950 170.400 319.050 171.600 ;
        RECT 298.950 169.950 301.050 170.400 ;
        RECT 316.950 169.950 319.050 170.400 ;
        RECT 370.950 171.600 373.050 172.050 ;
        RECT 424.950 171.600 427.050 172.050 ;
        RECT 370.950 170.400 427.050 171.600 ;
        RECT 370.950 169.950 373.050 170.400 ;
        RECT 424.950 169.950 427.050 170.400 ;
        RECT 427.950 171.600 430.050 172.050 ;
        RECT 434.400 171.600 435.600 173.400 ;
        RECT 559.950 172.950 562.050 173.400 ;
        RECT 592.950 172.950 595.050 173.400 ;
        RECT 616.950 174.600 619.050 175.050 ;
        RECT 676.950 174.600 679.050 175.050 ;
        RECT 616.950 173.400 679.050 174.600 ;
        RECT 616.950 172.950 619.050 173.400 ;
        RECT 676.950 172.950 679.050 173.400 ;
        RECT 682.950 174.600 685.050 175.050 ;
        RECT 712.950 174.600 715.050 175.050 ;
        RECT 727.950 174.600 730.050 175.050 ;
        RECT 739.950 174.600 742.050 175.050 ;
        RECT 682.950 173.400 742.050 174.600 ;
        RECT 682.950 172.950 685.050 173.400 ;
        RECT 712.950 172.950 715.050 173.400 ;
        RECT 727.950 172.950 730.050 173.400 ;
        RECT 739.950 172.950 742.050 173.400 ;
        RECT 427.950 170.400 435.600 171.600 ;
        RECT 442.950 171.600 445.050 172.050 ;
        RECT 451.950 171.600 454.050 172.050 ;
        RECT 442.950 170.400 454.050 171.600 ;
        RECT 427.950 169.950 430.050 170.400 ;
        RECT 442.950 169.950 445.050 170.400 ;
        RECT 451.950 169.950 454.050 170.400 ;
        RECT 454.950 171.600 457.050 172.050 ;
        RECT 475.950 171.600 478.050 172.050 ;
        RECT 454.950 170.400 478.050 171.600 ;
        RECT 454.950 169.950 457.050 170.400 ;
        RECT 475.950 169.950 478.050 170.400 ;
        RECT 484.950 171.600 487.050 172.050 ;
        RECT 505.950 171.600 508.050 172.050 ;
        RECT 484.950 170.400 508.050 171.600 ;
        RECT 484.950 169.950 487.050 170.400 ;
        RECT 505.950 169.950 508.050 170.400 ;
        RECT 547.950 171.600 550.050 172.050 ;
        RECT 601.950 171.600 604.050 172.050 ;
        RECT 619.950 171.600 622.050 172.050 ;
        RECT 628.950 171.600 631.050 172.050 ;
        RECT 547.950 170.400 600.600 171.600 ;
        RECT 547.950 169.950 550.050 170.400 ;
        RECT 13.950 168.600 16.050 169.050 ;
        RECT 19.950 168.600 22.050 169.050 ;
        RECT 13.950 167.400 22.050 168.600 ;
        RECT 13.950 166.950 16.050 167.400 ;
        RECT 19.950 166.950 22.050 167.400 ;
        RECT 40.950 168.600 43.050 169.050 ;
        RECT 64.950 168.600 67.050 169.050 ;
        RECT 40.950 167.400 67.050 168.600 ;
        RECT 40.950 166.950 43.050 167.400 ;
        RECT 64.950 166.950 67.050 167.400 ;
        RECT 82.950 168.600 85.050 169.050 ;
        RECT 109.950 168.600 112.050 169.050 ;
        RECT 121.950 168.600 124.050 169.050 ;
        RECT 169.950 168.600 172.050 169.050 ;
        RECT 82.950 167.400 87.600 168.600 ;
        RECT 82.950 166.950 85.050 167.400 ;
        RECT 86.400 166.050 87.600 167.400 ;
        RECT 109.950 167.400 120.600 168.600 ;
        RECT 109.950 166.950 112.050 167.400 ;
        RECT 1.950 165.600 4.050 166.050 ;
        RECT 10.950 165.600 13.050 166.050 ;
        RECT 1.950 164.400 13.050 165.600 ;
        RECT 1.950 163.950 4.050 164.400 ;
        RECT 10.950 163.950 13.050 164.400 ;
        RECT 25.950 165.600 28.050 166.050 ;
        RECT 34.950 165.600 37.050 166.050 ;
        RECT 25.950 164.400 37.050 165.600 ;
        RECT 25.950 163.950 28.050 164.400 ;
        RECT 34.950 163.950 37.050 164.400 ;
        RECT 40.950 165.600 43.050 166.050 ;
        RECT 55.950 165.600 58.050 166.050 ;
        RECT 40.950 164.400 58.050 165.600 ;
        RECT 40.950 163.950 43.050 164.400 ;
        RECT 55.950 163.950 58.050 164.400 ;
        RECT 67.950 163.950 70.050 166.050 ;
        RECT 85.950 163.950 88.050 166.050 ;
        RECT 91.950 165.600 94.050 166.050 ;
        RECT 89.400 164.400 94.050 165.600 ;
        RECT 43.950 162.600 46.050 163.050 ;
        RECT 68.400 162.600 69.600 163.950 ;
        RECT 89.400 162.600 90.600 164.400 ;
        RECT 91.950 163.950 94.050 164.400 ;
        RECT 115.950 163.950 118.050 166.050 ;
        RECT 119.400 165.600 120.600 167.400 ;
        RECT 121.950 167.400 172.050 168.600 ;
        RECT 121.950 166.950 124.050 167.400 ;
        RECT 169.950 166.950 172.050 167.400 ;
        RECT 184.950 166.950 187.050 169.050 ;
        RECT 241.950 166.950 244.050 169.050 ;
        RECT 247.950 168.600 250.050 169.050 ;
        RECT 253.950 168.600 256.050 169.050 ;
        RECT 247.950 167.400 256.050 168.600 ;
        RECT 247.950 166.950 250.050 167.400 ;
        RECT 253.950 166.950 256.050 167.400 ;
        RECT 262.950 166.950 265.050 169.050 ;
        RECT 292.950 168.600 295.050 169.050 ;
        RECT 281.400 167.400 295.050 168.600 ;
        RECT 124.950 165.600 127.050 166.050 ;
        RECT 119.400 164.400 127.050 165.600 ;
        RECT 124.950 163.950 127.050 164.400 ;
        RECT 151.950 165.600 154.050 166.050 ;
        RECT 166.950 165.600 169.050 166.050 ;
        RECT 151.950 164.400 169.050 165.600 ;
        RECT 151.950 163.950 154.050 164.400 ;
        RECT 166.950 163.950 169.050 164.400 ;
        RECT 43.950 161.400 90.600 162.600 ;
        RECT 43.950 160.950 46.050 161.400 ;
        RECT 62.400 160.050 63.600 161.400 ;
        RECT 112.950 160.950 115.050 163.050 ;
        RECT 116.400 162.600 117.600 163.950 ;
        RECT 185.400 163.050 186.600 166.950 ;
        RECT 187.950 165.600 190.050 166.050 ;
        RECT 193.950 165.600 196.050 166.050 ;
        RECT 187.950 164.400 196.050 165.600 ;
        RECT 187.950 163.950 190.050 164.400 ;
        RECT 193.950 163.950 196.050 164.400 ;
        RECT 199.950 165.600 202.050 166.050 ;
        RECT 208.950 165.600 211.050 166.050 ;
        RECT 220.950 165.600 223.050 166.050 ;
        RECT 232.950 165.600 235.050 166.050 ;
        RECT 242.400 165.600 243.600 166.950 ;
        RECT 199.950 164.400 207.600 165.600 ;
        RECT 199.950 163.950 202.050 164.400 ;
        RECT 157.950 162.600 160.050 163.050 ;
        RECT 116.400 161.400 160.050 162.600 ;
        RECT 157.950 160.950 160.050 161.400 ;
        RECT 169.950 162.600 172.050 163.050 ;
        RECT 175.950 162.600 178.050 163.050 ;
        RECT 169.950 161.400 178.050 162.600 ;
        RECT 169.950 160.950 172.050 161.400 ;
        RECT 175.950 160.950 178.050 161.400 ;
        RECT 184.950 160.950 187.050 163.050 ;
        RECT 206.400 162.600 207.600 164.400 ;
        RECT 208.950 164.400 235.050 165.600 ;
        RECT 208.950 163.950 211.050 164.400 ;
        RECT 220.950 163.950 223.050 164.400 ;
        RECT 232.950 163.950 235.050 164.400 ;
        RECT 239.400 164.400 243.600 165.600 ;
        RECT 263.400 165.600 264.600 166.950 ;
        RECT 281.400 166.050 282.600 167.400 ;
        RECT 292.950 166.950 295.050 167.400 ;
        RECT 319.950 168.600 322.050 169.050 ;
        RECT 331.950 168.600 334.050 169.050 ;
        RECT 319.950 167.400 334.050 168.600 ;
        RECT 319.950 166.950 322.050 167.400 ;
        RECT 331.950 166.950 334.050 167.400 ;
        RECT 334.950 168.600 337.050 169.050 ;
        RECT 364.950 168.600 367.050 169.050 ;
        RECT 382.950 168.600 385.050 169.050 ;
        RECT 334.950 167.400 345.600 168.600 ;
        RECT 334.950 166.950 337.050 167.400 ;
        RECT 265.950 165.600 268.050 166.050 ;
        RECT 263.400 164.400 268.050 165.600 ;
        RECT 235.950 162.600 238.050 163.050 ;
        RECT 206.400 161.400 238.050 162.600 ;
        RECT 235.950 160.950 238.050 161.400 ;
        RECT 61.950 157.950 64.050 160.050 ;
        RECT 113.400 159.600 114.600 160.950 ;
        RECT 239.400 160.050 240.600 164.400 ;
        RECT 265.950 163.950 268.050 164.400 ;
        RECT 280.950 163.950 283.050 166.050 ;
        RECT 295.950 165.600 298.050 166.050 ;
        RECT 307.950 165.600 310.050 166.050 ;
        RECT 295.950 164.400 310.050 165.600 ;
        RECT 295.950 163.950 298.050 164.400 ;
        RECT 307.950 163.950 310.050 164.400 ;
        RECT 313.950 165.600 316.050 166.050 ;
        RECT 319.950 165.600 322.050 166.050 ;
        RECT 313.950 164.400 322.050 165.600 ;
        RECT 313.950 163.950 316.050 164.400 ;
        RECT 319.950 163.950 322.050 164.400 ;
        RECT 334.950 165.600 337.050 166.050 ;
        RECT 340.950 165.600 343.050 166.050 ;
        RECT 334.950 164.400 343.050 165.600 ;
        RECT 334.950 163.950 337.050 164.400 ;
        RECT 340.950 163.950 343.050 164.400 ;
        RECT 344.400 163.050 345.600 167.400 ;
        RECT 347.400 167.400 367.050 168.600 ;
        RECT 347.400 166.050 348.600 167.400 ;
        RECT 364.950 166.950 367.050 167.400 ;
        RECT 371.400 167.400 385.050 168.600 ;
        RECT 346.950 163.950 349.050 166.050 ;
        RECT 349.950 165.600 352.050 166.050 ;
        RECT 361.950 165.600 364.050 166.050 ;
        RECT 349.950 164.400 364.050 165.600 ;
        RECT 349.950 163.950 352.050 164.400 ;
        RECT 361.950 163.950 364.050 164.400 ;
        RECT 371.400 163.050 372.600 167.400 ;
        RECT 382.950 166.950 385.050 167.400 ;
        RECT 421.950 166.950 424.050 169.050 ;
        RECT 430.950 168.600 433.050 169.050 ;
        RECT 425.400 167.400 433.050 168.600 ;
        RECT 412.950 165.600 415.050 166.050 ;
        RECT 422.400 165.600 423.600 166.950 ;
        RECT 425.400 166.050 426.600 167.400 ;
        RECT 430.950 166.950 433.050 167.400 ;
        RECT 457.950 168.600 460.050 169.050 ;
        RECT 466.950 168.600 469.050 169.050 ;
        RECT 457.950 167.400 469.050 168.600 ;
        RECT 457.950 166.950 460.050 167.400 ;
        RECT 466.950 166.950 469.050 167.400 ;
        RECT 496.950 168.600 499.050 169.050 ;
        RECT 526.950 168.600 529.050 169.050 ;
        RECT 547.950 168.600 550.050 169.050 ;
        RECT 496.950 167.400 516.600 168.600 ;
        RECT 496.950 166.950 499.050 167.400 ;
        RECT 515.400 166.050 516.600 167.400 ;
        RECT 526.950 167.400 550.050 168.600 ;
        RECT 526.950 166.950 529.050 167.400 ;
        RECT 547.950 166.950 550.050 167.400 ;
        RECT 571.950 168.600 574.050 169.050 ;
        RECT 571.950 167.400 591.600 168.600 ;
        RECT 571.950 166.950 574.050 167.400 ;
        RECT 412.950 164.400 423.600 165.600 ;
        RECT 412.950 163.950 415.050 164.400 ;
        RECT 424.950 163.950 427.050 166.050 ;
        RECT 430.950 165.600 433.050 166.050 ;
        RECT 442.950 165.600 445.050 166.050 ;
        RECT 493.950 165.600 496.050 166.050 ;
        RECT 430.950 164.400 445.050 165.600 ;
        RECT 430.950 163.950 433.050 164.400 ;
        RECT 442.950 163.950 445.050 164.400 ;
        RECT 458.400 164.400 496.050 165.600 ;
        RECT 241.950 162.600 244.050 163.050 ;
        RECT 256.950 162.600 259.050 163.050 ;
        RECT 241.950 161.400 259.050 162.600 ;
        RECT 241.950 160.950 244.050 161.400 ;
        RECT 256.950 160.950 259.050 161.400 ;
        RECT 304.950 162.600 307.050 163.050 ;
        RECT 322.950 162.600 325.050 163.050 ;
        RECT 304.950 161.400 325.050 162.600 ;
        RECT 304.950 160.950 307.050 161.400 ;
        RECT 322.950 160.950 325.050 161.400 ;
        RECT 343.950 160.950 346.050 163.050 ;
        RECT 370.950 160.950 373.050 163.050 ;
        RECT 376.950 162.600 379.050 163.050 ;
        RECT 379.950 162.600 382.050 163.050 ;
        RECT 397.950 162.600 400.050 163.050 ;
        RECT 439.950 162.600 442.050 163.050 ;
        RECT 376.950 161.400 442.050 162.600 ;
        RECT 376.950 160.950 379.050 161.400 ;
        RECT 379.950 160.950 382.050 161.400 ;
        RECT 397.950 160.950 400.050 161.400 ;
        RECT 439.950 160.950 442.050 161.400 ;
        RECT 445.950 162.600 448.050 163.050 ;
        RECT 458.400 162.600 459.600 164.400 ;
        RECT 493.950 163.950 496.050 164.400 ;
        RECT 499.950 165.600 502.050 166.050 ;
        RECT 499.950 164.400 513.600 165.600 ;
        RECT 499.950 163.950 502.050 164.400 ;
        RECT 445.950 161.400 459.600 162.600 ;
        RECT 463.950 162.600 466.050 163.050 ;
        RECT 472.950 162.600 475.050 163.050 ;
        RECT 463.950 161.400 475.050 162.600 ;
        RECT 445.950 160.950 448.050 161.400 ;
        RECT 463.950 160.950 466.050 161.400 ;
        RECT 472.950 160.950 475.050 161.400 ;
        RECT 487.950 162.600 490.050 163.050 ;
        RECT 496.950 162.600 499.050 163.050 ;
        RECT 487.950 161.400 499.050 162.600 ;
        RECT 512.400 162.600 513.600 164.400 ;
        RECT 514.950 163.950 517.050 166.050 ;
        RECT 541.950 165.600 544.050 166.050 ;
        RECT 553.950 165.600 556.050 166.050 ;
        RECT 568.950 165.600 571.050 166.050 ;
        RECT 580.950 165.600 583.050 166.050 ;
        RECT 586.950 165.600 589.050 166.050 ;
        RECT 541.950 164.400 589.050 165.600 ;
        RECT 541.950 163.950 544.050 164.400 ;
        RECT 553.950 163.950 556.050 164.400 ;
        RECT 568.950 163.950 571.050 164.400 ;
        RECT 580.950 163.950 583.050 164.400 ;
        RECT 586.950 163.950 589.050 164.400 ;
        RECT 523.950 162.600 526.050 163.050 ;
        RECT 532.950 162.600 535.050 163.050 ;
        RECT 512.400 161.400 522.600 162.600 ;
        RECT 487.950 160.950 490.050 161.400 ;
        RECT 496.950 160.950 499.050 161.400 ;
        RECT 133.950 159.600 136.050 160.050 ;
        RECT 113.400 158.400 136.050 159.600 ;
        RECT 133.950 157.950 136.050 158.400 ;
        RECT 148.950 159.600 151.050 160.050 ;
        RECT 154.950 159.600 157.050 160.050 ;
        RECT 148.950 158.400 157.050 159.600 ;
        RECT 148.950 157.950 151.050 158.400 ;
        RECT 154.950 157.950 157.050 158.400 ;
        RECT 178.950 159.600 181.050 160.050 ;
        RECT 196.950 159.600 199.050 160.050 ;
        RECT 178.950 158.400 199.050 159.600 ;
        RECT 178.950 157.950 181.050 158.400 ;
        RECT 196.950 157.950 199.050 158.400 ;
        RECT 214.950 159.600 217.050 160.050 ;
        RECT 226.950 159.600 229.050 160.050 ;
        RECT 214.950 158.400 229.050 159.600 ;
        RECT 214.950 157.950 217.050 158.400 ;
        RECT 226.950 157.950 229.050 158.400 ;
        RECT 238.950 157.950 241.050 160.050 ;
        RECT 337.950 159.600 340.050 160.050 ;
        RECT 373.950 159.600 376.050 160.050 ;
        RECT 337.950 158.400 376.050 159.600 ;
        RECT 337.950 157.950 340.050 158.400 ;
        RECT 373.950 157.950 376.050 158.400 ;
        RECT 385.950 159.600 388.050 160.050 ;
        RECT 436.950 159.600 439.050 160.050 ;
        RECT 385.950 158.400 439.050 159.600 ;
        RECT 385.950 157.950 388.050 158.400 ;
        RECT 436.950 157.950 439.050 158.400 ;
        RECT 439.950 159.600 442.050 160.050 ;
        RECT 481.950 159.600 484.050 160.050 ;
        RECT 517.950 159.600 520.050 160.050 ;
        RECT 439.950 158.400 520.050 159.600 ;
        RECT 521.400 159.600 522.600 161.400 ;
        RECT 523.950 161.400 535.050 162.600 ;
        RECT 523.950 160.950 526.050 161.400 ;
        RECT 532.950 160.950 535.050 161.400 ;
        RECT 544.950 160.950 547.050 163.050 ;
        RECT 556.950 162.600 559.050 163.050 ;
        RECT 574.950 162.600 577.050 163.050 ;
        RECT 556.950 161.400 577.050 162.600 ;
        RECT 590.400 162.600 591.600 167.400 ;
        RECT 599.400 166.050 600.600 170.400 ;
        RECT 601.950 170.400 631.050 171.600 ;
        RECT 601.950 169.950 604.050 170.400 ;
        RECT 619.950 169.950 622.050 170.400 ;
        RECT 628.950 169.950 631.050 170.400 ;
        RECT 631.950 171.600 634.050 172.050 ;
        RECT 655.950 171.600 658.050 172.050 ;
        RECT 631.950 170.400 658.050 171.600 ;
        RECT 631.950 169.950 634.050 170.400 ;
        RECT 604.950 168.600 607.050 169.050 ;
        RECT 604.950 167.400 618.600 168.600 ;
        RECT 604.950 166.950 607.050 167.400 ;
        RECT 598.950 163.950 601.050 166.050 ;
        RECT 601.950 165.600 604.050 166.050 ;
        RECT 607.950 165.600 610.050 166.050 ;
        RECT 613.950 165.600 616.050 166.050 ;
        RECT 601.950 164.400 616.050 165.600 ;
        RECT 601.950 163.950 604.050 164.400 ;
        RECT 607.950 163.950 610.050 164.400 ;
        RECT 613.950 163.950 616.050 164.400 ;
        RECT 617.400 163.050 618.600 167.400 ;
        RECT 628.950 165.600 631.050 166.050 ;
        RECT 640.950 165.600 643.050 166.050 ;
        RECT 628.950 164.400 643.050 165.600 ;
        RECT 628.950 163.950 631.050 164.400 ;
        RECT 640.950 163.950 643.050 164.400 ;
        RECT 613.950 162.600 616.050 163.050 ;
        RECT 590.400 161.400 616.050 162.600 ;
        RECT 556.950 160.950 559.050 161.400 ;
        RECT 574.950 160.950 577.050 161.400 ;
        RECT 613.950 160.950 616.050 161.400 ;
        RECT 616.950 160.950 619.050 163.050 ;
        RECT 644.400 162.600 645.600 170.400 ;
        RECT 655.950 169.950 658.050 170.400 ;
        RECT 673.950 171.600 676.050 172.050 ;
        RECT 691.950 171.600 694.050 172.050 ;
        RECT 673.950 170.400 694.050 171.600 ;
        RECT 673.950 169.950 676.050 170.400 ;
        RECT 691.950 169.950 694.050 170.400 ;
        RECT 694.950 169.950 697.050 172.050 ;
        RECT 697.950 171.600 700.050 172.050 ;
        RECT 706.950 171.600 709.050 172.050 ;
        RECT 697.950 170.400 709.050 171.600 ;
        RECT 697.950 169.950 700.050 170.400 ;
        RECT 706.950 169.950 709.050 170.400 ;
        RECT 721.950 171.600 724.050 172.050 ;
        RECT 748.950 171.600 751.050 172.050 ;
        RECT 721.950 170.400 751.050 171.600 ;
        RECT 721.950 169.950 724.050 170.400 ;
        RECT 748.950 169.950 751.050 170.400 ;
        RECT 649.950 168.600 652.050 169.050 ;
        RECT 664.950 168.600 667.050 169.050 ;
        RECT 649.950 167.400 667.050 168.600 ;
        RECT 649.950 166.950 652.050 167.400 ;
        RECT 664.950 166.950 667.050 167.400 ;
        RECT 665.400 165.600 666.600 166.950 ;
        RECT 662.400 164.400 666.600 165.600 ;
        RECT 676.950 165.600 679.050 166.050 ;
        RECT 688.950 165.600 691.050 166.050 ;
        RECT 676.950 164.400 691.050 165.600 ;
        RECT 649.950 162.600 652.050 163.050 ;
        RECT 644.400 161.400 652.050 162.600 ;
        RECT 649.950 160.950 652.050 161.400 ;
        RECT 658.950 162.600 661.050 163.050 ;
        RECT 662.400 162.600 663.600 164.400 ;
        RECT 676.950 163.950 679.050 164.400 ;
        RECT 688.950 163.950 691.050 164.400 ;
        RECT 691.950 165.600 694.050 166.050 ;
        RECT 695.400 165.600 696.600 169.950 ;
        RECT 697.950 168.600 700.050 169.050 ;
        RECT 709.950 168.600 712.050 169.050 ;
        RECT 721.950 168.600 724.050 169.050 ;
        RECT 697.950 167.400 708.600 168.600 ;
        RECT 697.950 166.950 700.050 167.400 ;
        RECT 707.400 166.050 708.600 167.400 ;
        RECT 709.950 167.400 724.050 168.600 ;
        RECT 709.950 166.950 712.050 167.400 ;
        RECT 721.950 166.950 724.050 167.400 ;
        RECT 724.950 168.600 727.050 169.050 ;
        RECT 736.950 168.600 739.050 169.050 ;
        RECT 742.950 168.600 745.050 169.050 ;
        RECT 724.950 167.400 732.600 168.600 ;
        RECT 724.950 166.950 727.050 167.400 ;
        RECT 731.400 166.050 732.600 167.400 ;
        RECT 736.950 167.400 745.050 168.600 ;
        RECT 736.950 166.950 739.050 167.400 ;
        RECT 742.950 166.950 745.050 167.400 ;
        RECT 691.950 164.400 696.600 165.600 ;
        RECT 691.950 163.950 694.050 164.400 ;
        RECT 706.950 163.950 709.050 166.050 ;
        RECT 730.950 163.950 733.050 166.050 ;
        RECT 745.950 165.600 748.050 166.050 ;
        RECT 763.950 165.600 766.050 166.050 ;
        RECT 745.950 164.400 766.050 165.600 ;
        RECT 745.950 163.950 748.050 164.400 ;
        RECT 763.950 163.950 766.050 164.400 ;
        RECT 658.950 161.400 663.600 162.600 ;
        RECT 664.950 162.600 667.050 163.050 ;
        RECT 673.950 162.600 676.050 163.050 ;
        RECT 664.950 161.400 676.050 162.600 ;
        RECT 658.950 160.950 661.050 161.400 ;
        RECT 664.950 160.950 667.050 161.400 ;
        RECT 673.950 160.950 676.050 161.400 ;
        RECT 733.950 162.600 736.050 163.050 ;
        RECT 742.950 162.600 745.050 163.050 ;
        RECT 754.950 162.600 757.050 163.050 ;
        RECT 733.950 161.400 757.050 162.600 ;
        RECT 733.950 160.950 736.050 161.400 ;
        RECT 742.950 160.950 745.050 161.400 ;
        RECT 754.950 160.950 757.050 161.400 ;
        RECT 538.950 159.600 541.050 160.050 ;
        RECT 521.400 158.400 541.050 159.600 ;
        RECT 545.400 159.600 546.600 160.950 ;
        RECT 625.950 159.600 628.050 160.050 ;
        RECT 545.400 158.400 628.050 159.600 ;
        RECT 439.950 157.950 442.050 158.400 ;
        RECT 481.950 157.950 484.050 158.400 ;
        RECT 517.950 157.950 520.050 158.400 ;
        RECT 538.950 157.950 541.050 158.400 ;
        RECT 625.950 157.950 628.050 158.400 ;
        RECT 646.950 159.600 649.050 160.050 ;
        RECT 661.950 159.600 664.050 160.050 ;
        RECT 697.950 159.600 700.050 160.050 ;
        RECT 646.950 158.400 700.050 159.600 ;
        RECT 646.950 157.950 649.050 158.400 ;
        RECT 661.950 157.950 664.050 158.400 ;
        RECT 697.950 157.950 700.050 158.400 ;
        RECT 727.950 159.600 730.050 160.050 ;
        RECT 766.950 159.600 769.050 160.050 ;
        RECT 727.950 158.400 769.050 159.600 ;
        RECT 727.950 157.950 730.050 158.400 ;
        RECT 766.950 157.950 769.050 158.400 ;
        RECT 79.950 156.600 82.050 157.050 ;
        RECT 142.950 156.600 145.050 157.050 ;
        RECT 79.950 155.400 145.050 156.600 ;
        RECT 79.950 154.950 82.050 155.400 ;
        RECT 142.950 154.950 145.050 155.400 ;
        RECT 223.950 156.600 226.050 157.050 ;
        RECT 283.950 156.600 286.050 157.050 ;
        RECT 223.950 155.400 286.050 156.600 ;
        RECT 223.950 154.950 226.050 155.400 ;
        RECT 283.950 154.950 286.050 155.400 ;
        RECT 331.950 156.600 334.050 157.050 ;
        RECT 397.950 156.600 400.050 157.050 ;
        RECT 331.950 155.400 400.050 156.600 ;
        RECT 331.950 154.950 334.050 155.400 ;
        RECT 397.950 154.950 400.050 155.400 ;
        RECT 544.950 156.600 547.050 157.050 ;
        RECT 550.950 156.600 553.050 157.050 ;
        RECT 592.950 156.600 595.050 157.050 ;
        RECT 544.950 155.400 549.600 156.600 ;
        RECT 544.950 154.950 547.050 155.400 ;
        RECT 172.950 153.600 175.050 154.050 ;
        RECT 394.950 153.600 397.050 154.050 ;
        RECT 490.950 153.600 493.050 154.050 ;
        RECT 172.950 152.400 393.600 153.600 ;
        RECT 172.950 151.950 175.050 152.400 ;
        RECT 226.950 150.600 229.050 151.050 ;
        RECT 238.950 150.600 241.050 151.050 ;
        RECT 226.950 149.400 241.050 150.600 ;
        RECT 226.950 148.950 229.050 149.400 ;
        RECT 238.950 148.950 241.050 149.400 ;
        RECT 277.950 150.600 280.050 151.050 ;
        RECT 355.950 150.600 358.050 151.050 ;
        RECT 370.950 150.600 373.050 151.050 ;
        RECT 277.950 149.400 373.050 150.600 ;
        RECT 392.400 150.600 393.600 152.400 ;
        RECT 394.950 152.400 493.050 153.600 ;
        RECT 394.950 151.950 397.050 152.400 ;
        RECT 490.950 151.950 493.050 152.400 ;
        RECT 535.950 153.600 538.050 154.050 ;
        RECT 544.950 153.600 547.050 154.050 ;
        RECT 535.950 152.400 547.050 153.600 ;
        RECT 548.400 153.600 549.600 155.400 ;
        RECT 550.950 155.400 595.050 156.600 ;
        RECT 550.950 154.950 553.050 155.400 ;
        RECT 592.950 154.950 595.050 155.400 ;
        RECT 595.950 156.600 598.050 157.050 ;
        RECT 664.950 156.600 667.050 157.050 ;
        RECT 595.950 155.400 667.050 156.600 ;
        RECT 595.950 154.950 598.050 155.400 ;
        RECT 664.950 154.950 667.050 155.400 ;
        RECT 667.950 156.600 670.050 157.050 ;
        RECT 694.950 156.600 697.050 157.050 ;
        RECT 667.950 155.400 697.050 156.600 ;
        RECT 667.950 154.950 670.050 155.400 ;
        RECT 694.950 154.950 697.050 155.400 ;
        RECT 670.950 153.600 673.050 154.050 ;
        RECT 548.400 152.400 673.050 153.600 ;
        RECT 535.950 151.950 538.050 152.400 ;
        RECT 544.950 151.950 547.050 152.400 ;
        RECT 670.950 151.950 673.050 152.400 ;
        RECT 673.950 153.600 676.050 154.050 ;
        RECT 691.950 153.600 694.050 154.050 ;
        RECT 673.950 152.400 694.050 153.600 ;
        RECT 673.950 151.950 676.050 152.400 ;
        RECT 691.950 151.950 694.050 152.400 ;
        RECT 748.950 153.600 751.050 154.050 ;
        RECT 757.950 153.600 760.050 154.050 ;
        RECT 748.950 152.400 760.050 153.600 ;
        RECT 748.950 151.950 751.050 152.400 ;
        RECT 757.950 151.950 760.050 152.400 ;
        RECT 493.950 150.600 496.050 151.050 ;
        RECT 392.400 149.400 496.050 150.600 ;
        RECT 277.950 148.950 280.050 149.400 ;
        RECT 355.950 148.950 358.050 149.400 ;
        RECT 370.950 148.950 373.050 149.400 ;
        RECT 493.950 148.950 496.050 149.400 ;
        RECT 499.950 150.600 502.050 151.050 ;
        RECT 529.950 150.600 532.050 151.050 ;
        RECT 565.950 150.600 568.050 151.050 ;
        RECT 499.950 149.400 568.050 150.600 ;
        RECT 499.950 148.950 502.050 149.400 ;
        RECT 529.950 148.950 532.050 149.400 ;
        RECT 565.950 148.950 568.050 149.400 ;
        RECT 598.950 150.600 601.050 151.050 ;
        RECT 607.950 150.600 610.050 151.050 ;
        RECT 598.950 149.400 610.050 150.600 ;
        RECT 598.950 148.950 601.050 149.400 ;
        RECT 607.950 148.950 610.050 149.400 ;
        RECT 634.950 150.600 637.050 151.050 ;
        RECT 682.950 150.600 685.050 151.050 ;
        RECT 634.950 149.400 685.050 150.600 ;
        RECT 634.950 148.950 637.050 149.400 ;
        RECT 682.950 148.950 685.050 149.400 ;
        RECT 205.950 147.600 208.050 148.050 ;
        RECT 361.950 147.600 364.050 148.050 ;
        RECT 205.950 146.400 364.050 147.600 ;
        RECT 205.950 145.950 208.050 146.400 ;
        RECT 361.950 145.950 364.050 146.400 ;
        RECT 382.950 147.600 385.050 148.050 ;
        RECT 403.950 147.600 406.050 148.050 ;
        RECT 382.950 146.400 406.050 147.600 ;
        RECT 382.950 145.950 385.050 146.400 ;
        RECT 403.950 145.950 406.050 146.400 ;
        RECT 436.950 147.600 439.050 148.050 ;
        RECT 469.950 147.600 472.050 148.050 ;
        RECT 487.950 147.600 490.050 148.050 ;
        RECT 436.950 146.400 490.050 147.600 ;
        RECT 436.950 145.950 439.050 146.400 ;
        RECT 469.950 145.950 472.050 146.400 ;
        RECT 487.950 145.950 490.050 146.400 ;
        RECT 490.950 147.600 493.050 148.050 ;
        RECT 613.950 147.600 616.050 148.050 ;
        RECT 634.950 147.600 637.050 148.050 ;
        RECT 490.950 146.400 600.600 147.600 ;
        RECT 490.950 145.950 493.050 146.400 ;
        RECT 43.950 144.600 46.050 145.050 ;
        RECT 49.950 144.600 52.050 145.050 ;
        RECT 139.950 144.600 142.050 145.050 ;
        RECT 43.950 143.400 142.050 144.600 ;
        RECT 43.950 142.950 46.050 143.400 ;
        RECT 49.950 142.950 52.050 143.400 ;
        RECT 139.950 142.950 142.050 143.400 ;
        RECT 241.950 144.600 244.050 145.050 ;
        RECT 247.950 144.600 250.050 145.050 ;
        RECT 241.950 143.400 250.050 144.600 ;
        RECT 241.950 142.950 244.050 143.400 ;
        RECT 247.950 142.950 250.050 143.400 ;
        RECT 271.950 144.600 274.050 145.050 ;
        RECT 313.950 144.600 316.050 145.050 ;
        RECT 379.950 144.600 382.050 145.050 ;
        RECT 271.950 143.400 282.600 144.600 ;
        RECT 271.950 142.950 274.050 143.400 ;
        RECT 139.950 141.600 142.050 142.050 ;
        RECT 274.950 141.600 277.050 142.050 ;
        RECT 139.950 140.400 277.050 141.600 ;
        RECT 281.400 141.600 282.600 143.400 ;
        RECT 313.950 143.400 382.050 144.600 ;
        RECT 313.950 142.950 316.050 143.400 ;
        RECT 379.950 142.950 382.050 143.400 ;
        RECT 409.950 144.600 412.050 145.050 ;
        RECT 415.950 144.600 418.050 145.050 ;
        RECT 529.950 144.600 532.050 145.050 ;
        RECT 538.950 144.600 541.050 145.050 ;
        RECT 409.950 143.400 418.050 144.600 ;
        RECT 409.950 142.950 412.050 143.400 ;
        RECT 415.950 142.950 418.050 143.400 ;
        RECT 503.400 143.400 541.050 144.600 ;
        RECT 328.950 141.600 331.050 142.050 ;
        RECT 281.400 140.400 331.050 141.600 ;
        RECT 139.950 139.950 142.050 140.400 ;
        RECT 274.950 139.950 277.050 140.400 ;
        RECT 328.950 139.950 331.050 140.400 ;
        RECT 331.950 141.600 334.050 142.050 ;
        RECT 391.950 141.600 394.050 142.050 ;
        RECT 331.950 140.400 394.050 141.600 ;
        RECT 331.950 139.950 334.050 140.400 ;
        RECT 391.950 139.950 394.050 140.400 ;
        RECT 397.950 141.600 400.050 142.050 ;
        RECT 454.950 141.600 457.050 142.050 ;
        RECT 397.950 140.400 457.050 141.600 ;
        RECT 397.950 139.950 400.050 140.400 ;
        RECT 454.950 139.950 457.050 140.400 ;
        RECT 475.950 141.600 478.050 142.050 ;
        RECT 503.400 141.600 504.600 143.400 ;
        RECT 529.950 142.950 532.050 143.400 ;
        RECT 538.950 142.950 541.050 143.400 ;
        RECT 583.950 144.600 586.050 145.050 ;
        RECT 595.950 144.600 598.050 145.050 ;
        RECT 583.950 143.400 598.050 144.600 ;
        RECT 599.400 144.600 600.600 146.400 ;
        RECT 613.950 146.400 637.050 147.600 ;
        RECT 613.950 145.950 616.050 146.400 ;
        RECT 634.950 145.950 637.050 146.400 ;
        RECT 652.950 147.600 655.050 148.050 ;
        RECT 676.950 147.600 679.050 148.050 ;
        RECT 652.950 146.400 679.050 147.600 ;
        RECT 652.950 145.950 655.050 146.400 ;
        RECT 676.950 145.950 679.050 146.400 ;
        RECT 757.950 147.600 760.050 148.050 ;
        RECT 769.950 147.600 772.050 148.050 ;
        RECT 757.950 146.400 772.050 147.600 ;
        RECT 757.950 145.950 760.050 146.400 ;
        RECT 769.950 145.950 772.050 146.400 ;
        RECT 628.950 144.600 631.050 145.050 ;
        RECT 661.950 144.600 664.050 145.050 ;
        RECT 599.400 143.400 618.600 144.600 ;
        RECT 583.950 142.950 586.050 143.400 ;
        RECT 595.950 142.950 598.050 143.400 ;
        RECT 475.950 140.400 504.600 141.600 ;
        RECT 505.950 141.600 508.050 142.050 ;
        RECT 517.950 141.600 520.050 142.050 ;
        RECT 505.950 140.400 520.050 141.600 ;
        RECT 475.950 139.950 478.050 140.400 ;
        RECT 505.950 139.950 508.050 140.400 ;
        RECT 517.950 139.950 520.050 140.400 ;
        RECT 520.950 141.600 523.050 142.050 ;
        RECT 583.950 141.600 586.050 142.050 ;
        RECT 520.950 140.400 586.050 141.600 ;
        RECT 520.950 139.950 523.050 140.400 ;
        RECT 583.950 139.950 586.050 140.400 ;
        RECT 589.950 141.600 592.050 142.050 ;
        RECT 613.950 141.600 616.050 142.050 ;
        RECT 589.950 140.400 616.050 141.600 ;
        RECT 617.400 141.600 618.600 143.400 ;
        RECT 628.950 143.400 664.050 144.600 ;
        RECT 628.950 142.950 631.050 143.400 ;
        RECT 661.950 142.950 664.050 143.400 ;
        RECT 679.950 141.600 682.050 142.050 ;
        RECT 617.400 140.400 682.050 141.600 ;
        RECT 589.950 139.950 592.050 140.400 ;
        RECT 613.950 139.950 616.050 140.400 ;
        RECT 679.950 139.950 682.050 140.400 ;
        RECT 148.950 138.600 151.050 139.050 ;
        RECT 229.950 138.600 232.050 139.050 ;
        RECT 148.950 137.400 232.050 138.600 ;
        RECT 148.950 136.950 151.050 137.400 ;
        RECT 229.950 136.950 232.050 137.400 ;
        RECT 235.950 138.600 238.050 139.050 ;
        RECT 247.950 138.600 250.050 139.050 ;
        RECT 265.950 138.600 268.050 139.050 ;
        RECT 334.950 138.600 337.050 139.050 ;
        RECT 367.950 138.600 370.050 139.050 ;
        RECT 646.950 138.600 649.050 139.050 ;
        RECT 685.950 138.600 688.050 139.050 ;
        RECT 235.950 137.400 370.050 138.600 ;
        RECT 235.950 136.950 238.050 137.400 ;
        RECT 247.950 136.950 250.050 137.400 ;
        RECT 265.950 136.950 268.050 137.400 ;
        RECT 334.950 136.950 337.050 137.400 ;
        RECT 367.950 136.950 370.050 137.400 ;
        RECT 434.400 137.400 649.050 138.600 ;
        RECT 434.400 136.050 435.600 137.400 ;
        RECT 646.950 136.950 649.050 137.400 ;
        RECT 677.400 137.400 688.050 138.600 ;
        RECT 88.950 135.600 91.050 136.050 ;
        RECT 118.950 135.600 121.050 136.050 ;
        RECT 88.950 134.400 121.050 135.600 ;
        RECT 88.950 133.950 91.050 134.400 ;
        RECT 118.950 133.950 121.050 134.400 ;
        RECT 229.950 135.600 232.050 136.050 ;
        RECT 268.950 135.600 271.050 136.050 ;
        RECT 229.950 134.400 271.050 135.600 ;
        RECT 229.950 133.950 232.050 134.400 ;
        RECT 268.950 133.950 271.050 134.400 ;
        RECT 340.950 135.600 343.050 136.050 ;
        RECT 376.950 135.600 379.050 136.050 ;
        RECT 340.950 134.400 379.050 135.600 ;
        RECT 340.950 133.950 343.050 134.400 ;
        RECT 376.950 133.950 379.050 134.400 ;
        RECT 397.950 135.600 400.050 136.050 ;
        RECT 412.950 135.600 415.050 136.050 ;
        RECT 397.950 134.400 415.050 135.600 ;
        RECT 397.950 133.950 400.050 134.400 ;
        RECT 412.950 133.950 415.050 134.400 ;
        RECT 433.950 133.950 436.050 136.050 ;
        RECT 502.950 135.600 505.050 136.050 ;
        RECT 562.950 135.600 565.050 136.050 ;
        RECT 502.950 134.400 565.050 135.600 ;
        RECT 502.950 133.950 505.050 134.400 ;
        RECT 562.950 133.950 565.050 134.400 ;
        RECT 568.950 135.600 571.050 136.050 ;
        RECT 589.950 135.600 592.050 136.050 ;
        RECT 568.950 134.400 592.050 135.600 ;
        RECT 568.950 133.950 571.050 134.400 ;
        RECT 589.950 133.950 592.050 134.400 ;
        RECT 592.950 135.600 595.050 136.050 ;
        RECT 677.400 135.600 678.600 137.400 ;
        RECT 685.950 136.950 688.050 137.400 ;
        RECT 736.950 138.600 739.050 139.050 ;
        RECT 754.950 138.600 757.050 139.050 ;
        RECT 736.950 137.400 757.050 138.600 ;
        RECT 736.950 136.950 739.050 137.400 ;
        RECT 754.950 136.950 757.050 137.400 ;
        RECT 592.950 134.400 678.600 135.600 ;
        RECT 679.950 135.600 682.050 136.050 ;
        RECT 730.950 135.600 733.050 136.050 ;
        RECT 763.950 135.600 766.050 136.050 ;
        RECT 679.950 134.400 766.050 135.600 ;
        RECT 592.950 133.950 595.050 134.400 ;
        RECT 679.950 133.950 682.050 134.400 ;
        RECT 730.950 133.950 733.050 134.400 ;
        RECT 763.950 133.950 766.050 134.400 ;
        RECT 55.950 132.600 58.050 133.050 ;
        RECT 76.950 132.600 79.050 133.050 ;
        RECT 55.950 131.400 79.050 132.600 ;
        RECT 55.950 130.950 58.050 131.400 ;
        RECT 76.950 130.950 79.050 131.400 ;
        RECT 115.950 132.600 118.050 133.050 ;
        RECT 121.950 132.600 124.050 133.050 ;
        RECT 115.950 131.400 124.050 132.600 ;
        RECT 115.950 130.950 118.050 131.400 ;
        RECT 121.950 130.950 124.050 131.400 ;
        RECT 178.950 132.600 181.050 133.050 ;
        RECT 244.950 132.600 247.050 133.050 ;
        RECT 178.950 131.400 247.050 132.600 ;
        RECT 178.950 130.950 181.050 131.400 ;
        RECT 244.950 130.950 247.050 131.400 ;
        RECT 250.950 132.600 253.050 133.050 ;
        RECT 253.950 132.600 256.050 133.050 ;
        RECT 262.950 132.600 265.050 133.050 ;
        RECT 250.950 131.400 265.050 132.600 ;
        RECT 250.950 130.950 253.050 131.400 ;
        RECT 253.950 130.950 256.050 131.400 ;
        RECT 262.950 130.950 265.050 131.400 ;
        RECT 307.950 132.600 310.050 133.050 ;
        RECT 313.950 132.600 316.050 133.050 ;
        RECT 307.950 131.400 316.050 132.600 ;
        RECT 307.950 130.950 310.050 131.400 ;
        RECT 313.950 130.950 316.050 131.400 ;
        RECT 325.950 132.600 328.050 133.050 ;
        RECT 337.950 132.600 340.050 133.050 ;
        RECT 349.950 132.600 352.050 133.050 ;
        RECT 325.950 131.400 352.050 132.600 ;
        RECT 325.950 130.950 328.050 131.400 ;
        RECT 337.950 130.950 340.050 131.400 ;
        RECT 349.950 130.950 352.050 131.400 ;
        RECT 352.950 132.600 355.050 133.050 ;
        RECT 460.950 132.600 463.050 133.050 ;
        RECT 352.950 131.400 423.600 132.600 ;
        RECT 352.950 130.950 355.050 131.400 ;
        RECT 28.950 129.600 31.050 130.050 ;
        RECT 34.950 129.600 37.050 130.050 ;
        RECT 37.950 129.600 40.050 130.050 ;
        RECT 28.950 128.400 40.050 129.600 ;
        RECT 28.950 127.950 31.050 128.400 ;
        RECT 34.950 127.950 37.050 128.400 ;
        RECT 37.950 127.950 40.050 128.400 ;
        RECT 100.950 129.600 103.050 130.050 ;
        RECT 115.950 129.600 118.050 130.050 ;
        RECT 127.950 129.600 130.050 130.050 ;
        RECT 100.950 128.400 118.050 129.600 ;
        RECT 100.950 127.950 103.050 128.400 ;
        RECT 115.950 127.950 118.050 128.400 ;
        RECT 125.400 128.400 130.050 129.600 ;
        RECT 13.950 126.600 16.050 127.050 ;
        RECT 28.950 126.600 31.050 127.050 ;
        RECT 13.950 125.400 31.050 126.600 ;
        RECT 13.950 124.950 16.050 125.400 ;
        RECT 28.950 124.950 31.050 125.400 ;
        RECT 37.950 124.950 40.050 127.050 ;
        RECT 58.950 126.600 61.050 127.050 ;
        RECT 64.950 126.600 67.050 127.050 ;
        RECT 67.950 126.600 70.050 127.050 ;
        RECT 58.950 125.400 70.050 126.600 ;
        RECT 58.950 124.950 61.050 125.400 ;
        RECT 64.950 124.950 67.050 125.400 ;
        RECT 67.950 124.950 70.050 125.400 ;
        RECT 73.950 124.950 76.050 127.050 ;
        RECT 112.950 126.600 115.050 127.050 ;
        RECT 125.400 126.600 126.600 128.400 ;
        RECT 127.950 127.950 130.050 128.400 ;
        RECT 136.950 129.600 139.050 130.050 ;
        RECT 142.950 129.600 145.050 130.050 ;
        RECT 172.950 129.600 175.050 130.050 ;
        RECT 136.950 128.400 175.050 129.600 ;
        RECT 136.950 127.950 139.050 128.400 ;
        RECT 142.950 127.950 145.050 128.400 ;
        RECT 172.950 127.950 175.050 128.400 ;
        RECT 217.950 129.600 220.050 130.050 ;
        RECT 229.950 129.600 232.050 130.050 ;
        RECT 256.950 129.600 259.050 130.050 ;
        RECT 217.950 128.400 232.050 129.600 ;
        RECT 217.950 127.950 220.050 128.400 ;
        RECT 229.950 127.950 232.050 128.400 ;
        RECT 251.400 128.400 259.050 129.600 ;
        RECT 112.950 125.400 126.600 126.600 ;
        RECT 175.950 126.600 178.050 127.050 ;
        RECT 184.950 126.600 187.050 127.050 ;
        RECT 175.950 125.400 187.050 126.600 ;
        RECT 112.950 124.950 115.050 125.400 ;
        RECT 175.950 124.950 178.050 125.400 ;
        RECT 184.950 124.950 187.050 125.400 ;
        RECT 190.950 124.950 193.050 127.050 ;
        RECT 25.950 123.600 28.050 124.050 ;
        RECT 38.400 123.600 39.600 124.950 ;
        RECT 70.950 123.600 73.050 124.050 ;
        RECT 25.950 122.400 73.050 123.600 ;
        RECT 74.400 123.600 75.600 124.950 ;
        RECT 133.950 123.600 136.050 124.050 ;
        RECT 74.400 122.400 136.050 123.600 ;
        RECT 191.400 123.600 192.600 124.950 ;
        RECT 202.950 123.600 205.050 124.050 ;
        RECT 191.400 122.400 205.050 123.600 ;
        RECT 25.950 121.950 28.050 122.400 ;
        RECT 70.950 121.950 73.050 122.400 ;
        RECT 133.950 121.950 136.050 122.400 ;
        RECT 202.950 121.950 205.050 122.400 ;
        RECT 214.950 123.600 217.050 124.050 ;
        RECT 238.950 123.600 241.050 124.050 ;
        RECT 214.950 122.400 241.050 123.600 ;
        RECT 214.950 121.950 217.050 122.400 ;
        RECT 238.950 121.950 241.050 122.400 ;
        RECT 244.950 123.600 247.050 124.050 ;
        RECT 251.400 123.600 252.600 128.400 ;
        RECT 256.950 127.950 259.050 128.400 ;
        RECT 265.950 129.600 268.050 130.050 ;
        RECT 283.950 129.600 286.050 130.050 ;
        RECT 265.950 128.400 286.050 129.600 ;
        RECT 265.950 127.950 268.050 128.400 ;
        RECT 283.950 127.950 286.050 128.400 ;
        RECT 310.950 129.600 313.050 130.050 ;
        RECT 319.950 129.600 322.050 130.050 ;
        RECT 322.950 129.600 325.050 130.050 ;
        RECT 310.950 128.400 325.050 129.600 ;
        RECT 310.950 127.950 313.050 128.400 ;
        RECT 319.950 127.950 322.050 128.400 ;
        RECT 322.950 127.950 325.050 128.400 ;
        RECT 346.950 129.600 349.050 130.050 ;
        RECT 370.950 129.600 373.050 130.050 ;
        RECT 373.950 129.600 376.050 130.050 ;
        RECT 346.950 128.400 376.050 129.600 ;
        RECT 346.950 127.950 349.050 128.400 ;
        RECT 370.950 127.950 373.050 128.400 ;
        RECT 373.950 127.950 376.050 128.400 ;
        RECT 391.950 129.600 394.050 130.050 ;
        RECT 403.950 129.600 406.050 130.050 ;
        RECT 391.950 128.400 406.050 129.600 ;
        RECT 391.950 127.950 394.050 128.400 ;
        RECT 403.950 127.950 406.050 128.400 ;
        RECT 409.950 129.600 412.050 130.050 ;
        RECT 418.950 129.600 421.050 130.050 ;
        RECT 409.950 128.400 421.050 129.600 ;
        RECT 422.400 129.600 423.600 131.400 ;
        RECT 452.400 131.400 463.050 132.600 ;
        RECT 422.400 128.400 450.600 129.600 ;
        RECT 409.950 127.950 412.050 128.400 ;
        RECT 418.950 127.950 421.050 128.400 ;
        RECT 283.950 126.600 286.050 127.050 ;
        RECT 292.950 126.600 295.050 127.050 ;
        RECT 283.950 125.400 295.050 126.600 ;
        RECT 283.950 124.950 286.050 125.400 ;
        RECT 292.950 124.950 295.050 125.400 ;
        RECT 343.950 124.950 346.050 127.050 ;
        RECT 244.950 122.400 252.600 123.600 ;
        RECT 277.950 123.600 280.050 124.050 ;
        RECT 298.950 123.600 301.050 124.050 ;
        RECT 310.950 123.600 313.050 124.050 ;
        RECT 277.950 122.400 313.050 123.600 ;
        RECT 244.950 121.950 247.050 122.400 ;
        RECT 277.950 121.950 280.050 122.400 ;
        RECT 298.950 121.950 301.050 122.400 ;
        RECT 310.950 121.950 313.050 122.400 ;
        RECT 331.950 123.600 334.050 124.050 ;
        RECT 340.950 123.600 343.050 124.050 ;
        RECT 331.950 122.400 343.050 123.600 ;
        RECT 331.950 121.950 334.050 122.400 ;
        RECT 340.950 121.950 343.050 122.400 ;
        RECT 7.950 120.600 10.050 121.050 ;
        RECT 19.950 120.600 22.050 121.050 ;
        RECT 7.950 119.400 22.050 120.600 ;
        RECT 7.950 118.950 10.050 119.400 ;
        RECT 19.950 118.950 22.050 119.400 ;
        RECT 34.950 120.600 37.050 121.050 ;
        RECT 40.950 120.600 43.050 121.050 ;
        RECT 34.950 119.400 43.050 120.600 ;
        RECT 34.950 118.950 37.050 119.400 ;
        RECT 40.950 118.950 43.050 119.400 ;
        RECT 76.950 120.600 79.050 121.050 ;
        RECT 79.950 120.600 82.050 121.050 ;
        RECT 139.950 120.600 142.050 121.050 ;
        RECT 76.950 119.400 142.050 120.600 ;
        RECT 76.950 118.950 79.050 119.400 ;
        RECT 79.950 118.950 82.050 119.400 ;
        RECT 139.950 118.950 142.050 119.400 ;
        RECT 166.950 120.600 169.050 121.050 ;
        RECT 220.950 120.600 223.050 121.050 ;
        RECT 166.950 119.400 223.050 120.600 ;
        RECT 166.950 118.950 169.050 119.400 ;
        RECT 220.950 118.950 223.050 119.400 ;
        RECT 226.950 120.600 229.050 121.050 ;
        RECT 238.950 120.600 241.050 121.050 ;
        RECT 226.950 119.400 241.050 120.600 ;
        RECT 226.950 118.950 229.050 119.400 ;
        RECT 238.950 118.950 241.050 119.400 ;
        RECT 250.950 120.600 253.050 121.050 ;
        RECT 265.950 120.600 268.050 121.050 ;
        RECT 271.950 120.600 274.050 121.050 ;
        RECT 250.950 119.400 274.050 120.600 ;
        RECT 250.950 118.950 253.050 119.400 ;
        RECT 265.950 118.950 268.050 119.400 ;
        RECT 271.950 118.950 274.050 119.400 ;
        RECT 295.950 120.600 298.050 121.050 ;
        RECT 331.950 120.600 334.050 121.050 ;
        RECT 295.950 119.400 334.050 120.600 ;
        RECT 344.400 120.600 345.600 124.950 ;
        RECT 347.400 124.050 348.600 127.950 ;
        RECT 352.950 126.600 355.050 127.050 ;
        RECT 391.950 126.600 394.050 127.050 ;
        RECT 352.950 125.400 394.050 126.600 ;
        RECT 352.950 124.950 355.050 125.400 ;
        RECT 391.950 124.950 394.050 125.400 ;
        RECT 406.950 126.600 409.050 127.050 ;
        RECT 412.950 126.600 415.050 127.050 ;
        RECT 430.950 126.600 433.050 127.050 ;
        RECT 406.950 125.400 415.050 126.600 ;
        RECT 406.950 124.950 409.050 125.400 ;
        RECT 412.950 124.950 415.050 125.400 ;
        RECT 422.400 125.400 433.050 126.600 ;
        RECT 422.400 124.050 423.600 125.400 ;
        RECT 430.950 124.950 433.050 125.400 ;
        RECT 433.950 126.600 436.050 127.050 ;
        RECT 445.950 126.600 448.050 127.050 ;
        RECT 433.950 125.400 448.050 126.600 ;
        RECT 433.950 124.950 436.050 125.400 ;
        RECT 445.950 124.950 448.050 125.400 ;
        RECT 346.950 121.950 349.050 124.050 ;
        RECT 385.950 123.600 388.050 124.050 ;
        RECT 350.400 122.400 388.050 123.600 ;
        RECT 350.400 120.600 351.600 122.400 ;
        RECT 385.950 121.950 388.050 122.400 ;
        RECT 421.950 121.950 424.050 124.050 ;
        RECT 424.950 123.600 427.050 124.050 ;
        RECT 442.950 123.600 445.050 124.050 ;
        RECT 449.400 123.600 450.600 128.400 ;
        RECT 424.950 122.400 432.600 123.600 ;
        RECT 424.950 121.950 427.050 122.400 ;
        RECT 431.400 121.050 432.600 122.400 ;
        RECT 442.950 122.400 450.600 123.600 ;
        RECT 452.400 123.600 453.600 131.400 ;
        RECT 460.950 130.950 463.050 131.400 ;
        RECT 487.950 132.600 490.050 133.050 ;
        RECT 508.950 132.600 511.050 133.050 ;
        RECT 487.950 131.400 511.050 132.600 ;
        RECT 487.950 130.950 490.050 131.400 ;
        RECT 508.950 130.950 511.050 131.400 ;
        RECT 547.950 132.600 550.050 133.050 ;
        RECT 607.950 132.600 610.050 133.050 ;
        RECT 616.950 132.600 619.050 133.050 ;
        RECT 547.950 131.400 573.600 132.600 ;
        RECT 547.950 130.950 550.050 131.400 ;
        RECT 572.400 130.050 573.600 131.400 ;
        RECT 605.400 131.400 610.050 132.600 ;
        RECT 454.950 129.600 457.050 130.050 ;
        RECT 499.950 129.600 502.050 130.050 ;
        RECT 454.950 128.400 502.050 129.600 ;
        RECT 454.950 127.950 457.050 128.400 ;
        RECT 499.950 127.950 502.050 128.400 ;
        RECT 514.950 129.600 517.050 130.050 ;
        RECT 559.950 129.600 562.050 130.050 ;
        RECT 565.950 129.600 568.050 130.050 ;
        RECT 514.950 128.400 549.600 129.600 ;
        RECT 514.950 127.950 517.050 128.400 ;
        RECT 457.950 126.600 460.050 127.050 ;
        RECT 469.950 126.600 472.050 127.050 ;
        RECT 457.950 125.400 472.050 126.600 ;
        RECT 457.950 124.950 460.050 125.400 ;
        RECT 469.950 124.950 472.050 125.400 ;
        RECT 481.950 126.600 484.050 127.050 ;
        RECT 499.950 126.600 502.050 127.050 ;
        RECT 502.950 126.600 505.050 127.050 ;
        RECT 481.950 125.400 505.050 126.600 ;
        RECT 481.950 124.950 484.050 125.400 ;
        RECT 499.950 124.950 502.050 125.400 ;
        RECT 502.950 124.950 505.050 125.400 ;
        RECT 514.950 126.600 517.050 127.050 ;
        RECT 544.950 126.600 547.050 127.050 ;
        RECT 514.950 125.400 547.050 126.600 ;
        RECT 514.950 124.950 517.050 125.400 ;
        RECT 544.950 124.950 547.050 125.400 ;
        RECT 548.400 124.050 549.600 128.400 ;
        RECT 559.950 128.400 568.050 129.600 ;
        RECT 559.950 127.950 562.050 128.400 ;
        RECT 565.950 127.950 568.050 128.400 ;
        RECT 571.950 127.950 574.050 130.050 ;
        RECT 577.950 129.600 580.050 130.050 ;
        RECT 589.950 129.600 592.050 130.050 ;
        RECT 577.950 128.400 603.600 129.600 ;
        RECT 577.950 127.950 580.050 128.400 ;
        RECT 589.950 127.950 592.050 128.400 ;
        RECT 602.400 127.050 603.600 128.400 ;
        RECT 556.950 126.600 559.050 127.050 ;
        RECT 562.950 126.600 565.050 127.050 ;
        RECT 574.950 126.600 577.050 127.050 ;
        RECT 556.950 125.400 577.050 126.600 ;
        RECT 556.950 124.950 559.050 125.400 ;
        RECT 562.950 124.950 565.050 125.400 ;
        RECT 574.950 124.950 577.050 125.400 ;
        RECT 580.950 126.600 583.050 127.050 ;
        RECT 580.950 125.400 600.600 126.600 ;
        RECT 580.950 124.950 583.050 125.400 ;
        RECT 599.400 124.050 600.600 125.400 ;
        RECT 601.950 124.950 604.050 127.050 ;
        RECT 520.950 123.600 523.050 124.050 ;
        RECT 532.950 123.600 535.050 124.050 ;
        RECT 535.950 123.600 538.050 124.050 ;
        RECT 452.400 122.400 459.600 123.600 ;
        RECT 442.950 121.950 445.050 122.400 ;
        RECT 458.400 121.050 459.600 122.400 ;
        RECT 497.400 122.400 538.050 123.600 ;
        RECT 497.400 121.050 498.600 122.400 ;
        RECT 520.950 121.950 523.050 122.400 ;
        RECT 532.950 121.950 535.050 122.400 ;
        RECT 535.950 121.950 538.050 122.400 ;
        RECT 547.950 121.950 550.050 124.050 ;
        RECT 550.950 123.600 553.050 124.050 ;
        RECT 568.950 123.600 571.050 124.050 ;
        RECT 550.950 122.400 571.050 123.600 ;
        RECT 550.950 121.950 553.050 122.400 ;
        RECT 568.950 121.950 571.050 122.400 ;
        RECT 598.950 121.950 601.050 124.050 ;
        RECT 601.950 123.600 604.050 124.050 ;
        RECT 605.400 123.600 606.600 131.400 ;
        RECT 607.950 130.950 610.050 131.400 ;
        RECT 614.400 131.400 619.050 132.600 ;
        RECT 610.950 127.950 613.050 130.050 ;
        RECT 611.400 124.050 612.600 127.950 ;
        RECT 601.950 122.400 606.600 123.600 ;
        RECT 601.950 121.950 604.050 122.400 ;
        RECT 610.950 121.950 613.050 124.050 ;
        RECT 344.400 119.400 351.600 120.600 ;
        RECT 376.950 120.600 379.050 121.050 ;
        RECT 394.950 120.600 397.050 121.050 ;
        RECT 400.950 120.600 403.050 121.050 ;
        RECT 376.950 119.400 403.050 120.600 ;
        RECT 295.950 118.950 298.050 119.400 ;
        RECT 331.950 118.950 334.050 119.400 ;
        RECT 376.950 118.950 379.050 119.400 ;
        RECT 394.950 118.950 397.050 119.400 ;
        RECT 400.950 118.950 403.050 119.400 ;
        RECT 430.950 118.950 433.050 121.050 ;
        RECT 448.950 120.600 451.050 121.050 ;
        RECT 454.950 120.600 457.050 121.050 ;
        RECT 448.950 119.400 457.050 120.600 ;
        RECT 448.950 118.950 451.050 119.400 ;
        RECT 454.950 118.950 457.050 119.400 ;
        RECT 457.950 118.950 460.050 121.050 ;
        RECT 469.950 120.600 472.050 121.050 ;
        RECT 475.950 120.600 478.050 121.050 ;
        RECT 469.950 119.400 478.050 120.600 ;
        RECT 469.950 118.950 472.050 119.400 ;
        RECT 475.950 118.950 478.050 119.400 ;
        RECT 496.950 118.950 499.050 121.050 ;
        RECT 502.950 120.600 505.050 121.050 ;
        RECT 550.950 120.600 553.050 121.050 ;
        RECT 502.950 119.400 553.050 120.600 ;
        RECT 502.950 118.950 505.050 119.400 ;
        RECT 550.950 118.950 553.050 119.400 ;
        RECT 553.950 120.600 556.050 121.050 ;
        RECT 583.950 120.600 586.050 121.050 ;
        RECT 553.950 119.400 586.050 120.600 ;
        RECT 553.950 118.950 556.050 119.400 ;
        RECT 583.950 118.950 586.050 119.400 ;
        RECT 607.950 120.600 610.050 121.050 ;
        RECT 614.400 120.600 615.600 131.400 ;
        RECT 616.950 130.950 619.050 131.400 ;
        RECT 622.950 132.600 625.050 133.050 ;
        RECT 643.950 132.600 646.050 133.050 ;
        RECT 622.950 131.400 646.050 132.600 ;
        RECT 622.950 130.950 625.050 131.400 ;
        RECT 643.950 130.950 646.050 131.400 ;
        RECT 670.950 132.600 673.050 133.050 ;
        RECT 700.950 132.600 703.050 133.050 ;
        RECT 706.950 132.600 709.050 133.050 ;
        RECT 670.950 131.400 690.600 132.600 ;
        RECT 670.950 130.950 673.050 131.400 ;
        RECT 689.400 130.050 690.600 131.400 ;
        RECT 700.950 131.400 709.050 132.600 ;
        RECT 700.950 130.950 703.050 131.400 ;
        RECT 706.950 130.950 709.050 131.400 ;
        RECT 721.950 132.600 724.050 133.050 ;
        RECT 742.950 132.600 745.050 133.050 ;
        RECT 721.950 131.400 745.050 132.600 ;
        RECT 721.950 130.950 724.050 131.400 ;
        RECT 742.950 130.950 745.050 131.400 ;
        RECT 631.950 129.600 634.050 130.050 ;
        RECT 637.950 129.600 640.050 130.050 ;
        RECT 617.400 128.400 634.050 129.600 ;
        RECT 617.400 127.050 618.600 128.400 ;
        RECT 631.950 127.950 634.050 128.400 ;
        RECT 635.400 128.400 640.050 129.600 ;
        RECT 616.950 124.950 619.050 127.050 ;
        RECT 622.950 126.600 625.050 127.050 ;
        RECT 631.950 126.600 634.050 127.050 ;
        RECT 622.950 125.400 634.050 126.600 ;
        RECT 622.950 124.950 625.050 125.400 ;
        RECT 631.950 124.950 634.050 125.400 ;
        RECT 625.950 123.600 628.050 124.050 ;
        RECT 635.400 123.600 636.600 128.400 ;
        RECT 637.950 127.950 640.050 128.400 ;
        RECT 649.950 129.600 652.050 130.050 ;
        RECT 676.950 129.600 679.050 130.050 ;
        RECT 649.950 128.400 679.050 129.600 ;
        RECT 649.950 127.950 652.050 128.400 ;
        RECT 676.950 127.950 679.050 128.400 ;
        RECT 688.950 127.950 691.050 130.050 ;
        RECT 697.950 129.600 700.050 130.050 ;
        RECT 709.950 129.600 712.050 130.050 ;
        RECT 697.950 128.400 712.050 129.600 ;
        RECT 697.950 127.950 700.050 128.400 ;
        RECT 709.950 127.950 712.050 128.400 ;
        RECT 715.950 129.600 718.050 130.050 ;
        RECT 715.950 128.400 732.600 129.600 ;
        RECT 715.950 127.950 718.050 128.400 ;
        RECT 731.400 127.050 732.600 128.400 ;
        RECT 649.950 126.600 652.050 127.050 ;
        RECT 655.950 126.600 658.050 127.050 ;
        RECT 658.950 126.600 661.050 127.050 ;
        RECT 649.950 125.400 661.050 126.600 ;
        RECT 649.950 124.950 652.050 125.400 ;
        RECT 655.950 124.950 658.050 125.400 ;
        RECT 658.950 124.950 661.050 125.400 ;
        RECT 670.950 126.600 673.050 127.050 ;
        RECT 685.950 126.600 688.050 127.050 ;
        RECT 703.950 126.600 706.050 127.050 ;
        RECT 670.950 125.400 706.050 126.600 ;
        RECT 670.950 124.950 673.050 125.400 ;
        RECT 685.950 124.950 688.050 125.400 ;
        RECT 703.950 124.950 706.050 125.400 ;
        RECT 721.950 126.600 724.050 127.050 ;
        RECT 727.950 126.600 730.050 127.050 ;
        RECT 721.950 125.400 730.050 126.600 ;
        RECT 721.950 124.950 724.050 125.400 ;
        RECT 727.950 124.950 730.050 125.400 ;
        RECT 730.950 124.950 733.050 127.050 ;
        RECT 625.950 122.400 636.600 123.600 ;
        RECT 676.950 123.600 679.050 124.050 ;
        RECT 691.950 123.600 694.050 124.050 ;
        RECT 694.950 123.600 697.050 124.050 ;
        RECT 676.950 122.400 697.050 123.600 ;
        RECT 625.950 121.950 628.050 122.400 ;
        RECT 676.950 121.950 679.050 122.400 ;
        RECT 691.950 121.950 694.050 122.400 ;
        RECT 694.950 121.950 697.050 122.400 ;
        RECT 703.950 123.600 706.050 124.050 ;
        RECT 736.950 123.600 739.050 124.050 ;
        RECT 703.950 122.400 739.050 123.600 ;
        RECT 703.950 121.950 706.050 122.400 ;
        RECT 736.950 121.950 739.050 122.400 ;
        RECT 739.950 123.600 742.050 124.050 ;
        RECT 745.950 123.600 748.050 124.050 ;
        RECT 739.950 122.400 748.050 123.600 ;
        RECT 739.950 121.950 742.050 122.400 ;
        RECT 745.950 121.950 748.050 122.400 ;
        RECT 607.950 119.400 615.600 120.600 ;
        RECT 658.950 120.600 661.050 121.050 ;
        RECT 667.950 120.600 670.050 121.050 ;
        RECT 688.950 120.600 691.050 121.050 ;
        RECT 658.950 119.400 691.050 120.600 ;
        RECT 607.950 118.950 610.050 119.400 ;
        RECT 658.950 118.950 661.050 119.400 ;
        RECT 667.950 118.950 670.050 119.400 ;
        RECT 688.950 118.950 691.050 119.400 ;
        RECT 718.950 120.600 721.050 121.050 ;
        RECT 724.950 120.600 727.050 121.050 ;
        RECT 718.950 119.400 727.050 120.600 ;
        RECT 718.950 118.950 721.050 119.400 ;
        RECT 724.950 118.950 727.050 119.400 ;
        RECT 751.950 120.600 754.050 121.050 ;
        RECT 757.950 120.600 760.050 121.050 ;
        RECT 751.950 119.400 760.050 120.600 ;
        RECT 751.950 118.950 754.050 119.400 ;
        RECT 757.950 118.950 760.050 119.400 ;
        RECT 31.950 117.600 34.050 118.050 ;
        RECT 49.950 117.600 52.050 118.050 ;
        RECT 31.950 116.400 52.050 117.600 ;
        RECT 31.950 115.950 34.050 116.400 ;
        RECT 49.950 115.950 52.050 116.400 ;
        RECT 187.950 117.600 190.050 118.050 ;
        RECT 250.950 117.600 253.050 118.050 ;
        RECT 187.950 116.400 253.050 117.600 ;
        RECT 187.950 115.950 190.050 116.400 ;
        RECT 250.950 115.950 253.050 116.400 ;
        RECT 286.950 117.600 289.050 118.050 ;
        RECT 316.950 117.600 319.050 118.050 ;
        RECT 286.950 116.400 319.050 117.600 ;
        RECT 286.950 115.950 289.050 116.400 ;
        RECT 316.950 115.950 319.050 116.400 ;
        RECT 340.950 117.600 343.050 118.050 ;
        RECT 361.950 117.600 364.050 118.050 ;
        RECT 472.950 117.600 475.050 118.050 ;
        RECT 340.950 116.400 475.050 117.600 ;
        RECT 340.950 115.950 343.050 116.400 ;
        RECT 361.950 115.950 364.050 116.400 ;
        RECT 472.950 115.950 475.050 116.400 ;
        RECT 478.950 117.600 481.050 118.050 ;
        RECT 523.950 117.600 526.050 118.050 ;
        RECT 553.950 117.600 556.050 118.050 ;
        RECT 478.950 116.400 556.050 117.600 ;
        RECT 478.950 115.950 481.050 116.400 ;
        RECT 523.950 115.950 526.050 116.400 ;
        RECT 553.950 115.950 556.050 116.400 ;
        RECT 565.950 117.600 568.050 118.050 ;
        RECT 619.950 117.600 622.050 118.050 ;
        RECT 634.950 117.600 637.050 118.050 ;
        RECT 565.950 116.400 637.050 117.600 ;
        RECT 565.950 115.950 568.050 116.400 ;
        RECT 619.950 115.950 622.050 116.400 ;
        RECT 634.950 115.950 637.050 116.400 ;
        RECT 646.950 117.600 649.050 118.050 ;
        RECT 700.950 117.600 703.050 118.050 ;
        RECT 646.950 116.400 703.050 117.600 ;
        RECT 646.950 115.950 649.050 116.400 ;
        RECT 700.950 115.950 703.050 116.400 ;
        RECT 16.950 114.600 19.050 115.050 ;
        RECT 46.950 114.600 49.050 115.050 ;
        RECT 16.950 113.400 49.050 114.600 ;
        RECT 16.950 112.950 19.050 113.400 ;
        RECT 46.950 112.950 49.050 113.400 ;
        RECT 97.950 114.600 100.050 115.050 ;
        RECT 118.950 114.600 121.050 115.050 ;
        RECT 148.950 114.600 151.050 115.050 ;
        RECT 160.950 114.600 163.050 115.050 ;
        RECT 97.950 113.400 163.050 114.600 ;
        RECT 97.950 112.950 100.050 113.400 ;
        RECT 118.950 112.950 121.050 113.400 ;
        RECT 148.950 112.950 151.050 113.400 ;
        RECT 160.950 112.950 163.050 113.400 ;
        RECT 196.950 114.600 199.050 115.050 ;
        RECT 235.950 114.600 238.050 115.050 ;
        RECT 196.950 113.400 238.050 114.600 ;
        RECT 196.950 112.950 199.050 113.400 ;
        RECT 235.950 112.950 238.050 113.400 ;
        RECT 259.950 114.600 262.050 115.050 ;
        RECT 277.950 114.600 280.050 115.050 ;
        RECT 259.950 113.400 280.050 114.600 ;
        RECT 259.950 112.950 262.050 113.400 ;
        RECT 277.950 112.950 280.050 113.400 ;
        RECT 283.950 114.600 286.050 115.050 ;
        RECT 301.950 114.600 304.050 115.050 ;
        RECT 283.950 113.400 304.050 114.600 ;
        RECT 283.950 112.950 286.050 113.400 ;
        RECT 301.950 112.950 304.050 113.400 ;
        RECT 304.950 114.600 307.050 115.050 ;
        RECT 307.950 114.600 310.050 115.050 ;
        RECT 511.950 114.600 514.050 115.050 ;
        RECT 304.950 113.400 514.050 114.600 ;
        RECT 304.950 112.950 307.050 113.400 ;
        RECT 307.950 112.950 310.050 113.400 ;
        RECT 511.950 112.950 514.050 113.400 ;
        RECT 541.950 114.600 544.050 115.050 ;
        RECT 622.950 114.600 625.050 115.050 ;
        RECT 541.950 113.400 625.050 114.600 ;
        RECT 541.950 112.950 544.050 113.400 ;
        RECT 622.950 112.950 625.050 113.400 ;
        RECT 649.950 114.600 652.050 115.050 ;
        RECT 751.950 114.600 754.050 115.050 ;
        RECT 649.950 113.400 754.050 114.600 ;
        RECT 649.950 112.950 652.050 113.400 ;
        RECT 751.950 112.950 754.050 113.400 ;
        RECT 211.950 111.600 214.050 112.050 ;
        RECT 220.950 111.600 223.050 112.050 ;
        RECT 241.950 111.600 244.050 112.050 ;
        RECT 211.950 110.400 244.050 111.600 ;
        RECT 211.950 109.950 214.050 110.400 ;
        RECT 220.950 109.950 223.050 110.400 ;
        RECT 241.950 109.950 244.050 110.400 ;
        RECT 244.950 111.600 247.050 112.050 ;
        RECT 265.950 111.600 268.050 112.050 ;
        RECT 244.950 110.400 268.050 111.600 ;
        RECT 244.950 109.950 247.050 110.400 ;
        RECT 265.950 109.950 268.050 110.400 ;
        RECT 271.950 111.600 274.050 112.050 ;
        RECT 283.950 111.600 286.050 112.050 ;
        RECT 289.950 111.600 292.050 112.050 ;
        RECT 271.950 110.400 292.050 111.600 ;
        RECT 271.950 109.950 274.050 110.400 ;
        RECT 283.950 109.950 286.050 110.400 ;
        RECT 289.950 109.950 292.050 110.400 ;
        RECT 316.950 111.600 319.050 112.050 ;
        RECT 379.950 111.600 382.050 112.050 ;
        RECT 316.950 110.400 382.050 111.600 ;
        RECT 316.950 109.950 319.050 110.400 ;
        RECT 379.950 109.950 382.050 110.400 ;
        RECT 382.950 111.600 385.050 112.050 ;
        RECT 394.950 111.600 397.050 112.050 ;
        RECT 382.950 110.400 397.050 111.600 ;
        RECT 382.950 109.950 385.050 110.400 ;
        RECT 394.950 109.950 397.050 110.400 ;
        RECT 397.950 111.600 400.050 112.050 ;
        RECT 418.950 111.600 421.050 112.050 ;
        RECT 397.950 110.400 421.050 111.600 ;
        RECT 397.950 109.950 400.050 110.400 ;
        RECT 418.950 109.950 421.050 110.400 ;
        RECT 433.950 111.600 436.050 112.050 ;
        RECT 487.950 111.600 490.050 112.050 ;
        RECT 433.950 110.400 490.050 111.600 ;
        RECT 433.950 109.950 436.050 110.400 ;
        RECT 487.950 109.950 490.050 110.400 ;
        RECT 526.950 111.600 529.050 112.050 ;
        RECT 586.950 111.600 589.050 112.050 ;
        RECT 604.950 111.600 607.050 112.050 ;
        RECT 526.950 110.400 607.050 111.600 ;
        RECT 526.950 109.950 529.050 110.400 ;
        RECT 586.950 109.950 589.050 110.400 ;
        RECT 604.950 109.950 607.050 110.400 ;
        RECT 628.950 111.600 631.050 112.050 ;
        RECT 646.950 111.600 649.050 112.050 ;
        RECT 694.950 111.600 697.050 112.050 ;
        RECT 628.950 110.400 697.050 111.600 ;
        RECT 628.950 109.950 631.050 110.400 ;
        RECT 646.950 109.950 649.050 110.400 ;
        RECT 694.950 109.950 697.050 110.400 ;
        RECT 241.950 108.600 244.050 109.050 ;
        RECT 262.950 108.600 265.050 109.050 ;
        RECT 241.950 107.400 265.050 108.600 ;
        RECT 241.950 106.950 244.050 107.400 ;
        RECT 262.950 106.950 265.050 107.400 ;
        RECT 277.950 108.600 280.050 109.050 ;
        RECT 316.950 108.600 319.050 109.050 ;
        RECT 277.950 107.400 319.050 108.600 ;
        RECT 277.950 106.950 280.050 107.400 ;
        RECT 316.950 106.950 319.050 107.400 ;
        RECT 325.950 108.600 328.050 109.050 ;
        RECT 406.950 108.600 409.050 109.050 ;
        RECT 325.950 107.400 409.050 108.600 ;
        RECT 325.950 106.950 328.050 107.400 ;
        RECT 406.950 106.950 409.050 107.400 ;
        RECT 439.950 108.600 442.050 109.050 ;
        RECT 652.950 108.600 655.050 109.050 ;
        RECT 439.950 107.400 655.050 108.600 ;
        RECT 439.950 106.950 442.050 107.400 ;
        RECT 652.950 106.950 655.050 107.400 ;
        RECT 679.950 108.600 682.050 109.050 ;
        RECT 703.950 108.600 706.050 109.050 ;
        RECT 679.950 107.400 706.050 108.600 ;
        RECT 679.950 106.950 682.050 107.400 ;
        RECT 703.950 106.950 706.050 107.400 ;
        RECT 19.950 105.600 22.050 106.050 ;
        RECT 46.950 105.600 49.050 106.050 ;
        RECT 19.950 104.400 49.050 105.600 ;
        RECT 19.950 103.950 22.050 104.400 ;
        RECT 46.950 103.950 49.050 104.400 ;
        RECT 172.950 105.600 175.050 106.050 ;
        RECT 190.950 105.600 193.050 106.050 ;
        RECT 172.950 104.400 193.050 105.600 ;
        RECT 172.950 103.950 175.050 104.400 ;
        RECT 190.950 103.950 193.050 104.400 ;
        RECT 193.950 105.600 196.050 106.050 ;
        RECT 196.950 105.600 199.050 106.050 ;
        RECT 244.950 105.600 247.050 106.050 ;
        RECT 193.950 104.400 247.050 105.600 ;
        RECT 193.950 103.950 196.050 104.400 ;
        RECT 196.950 103.950 199.050 104.400 ;
        RECT 244.950 103.950 247.050 104.400 ;
        RECT 262.950 105.600 265.050 106.050 ;
        RECT 280.950 105.600 283.050 106.050 ;
        RECT 262.950 104.400 283.050 105.600 ;
        RECT 262.950 103.950 265.050 104.400 ;
        RECT 280.950 103.950 283.050 104.400 ;
        RECT 325.950 105.600 328.050 106.050 ;
        RECT 343.950 105.600 346.050 106.050 ;
        RECT 325.950 104.400 346.050 105.600 ;
        RECT 325.950 103.950 328.050 104.400 ;
        RECT 343.950 103.950 346.050 104.400 ;
        RECT 346.950 105.600 349.050 106.050 ;
        RECT 388.950 105.600 391.050 106.050 ;
        RECT 346.950 104.400 391.050 105.600 ;
        RECT 346.950 103.950 349.050 104.400 ;
        RECT 388.950 103.950 391.050 104.400 ;
        RECT 427.950 105.600 430.050 106.050 ;
        RECT 442.950 105.600 445.050 106.050 ;
        RECT 484.950 105.600 487.050 106.050 ;
        RECT 427.950 104.400 487.050 105.600 ;
        RECT 427.950 103.950 430.050 104.400 ;
        RECT 442.950 103.950 445.050 104.400 ;
        RECT 484.950 103.950 487.050 104.400 ;
        RECT 487.950 105.600 490.050 106.050 ;
        RECT 550.950 105.600 553.050 106.050 ;
        RECT 487.950 104.400 553.050 105.600 ;
        RECT 487.950 103.950 490.050 104.400 ;
        RECT 550.950 103.950 553.050 104.400 ;
        RECT 610.950 105.600 613.050 106.050 ;
        RECT 637.950 105.600 640.050 106.050 ;
        RECT 697.950 105.600 700.050 106.050 ;
        RECT 712.950 105.600 715.050 106.050 ;
        RECT 610.950 104.400 715.050 105.600 ;
        RECT 610.950 103.950 613.050 104.400 ;
        RECT 637.950 103.950 640.050 104.400 ;
        RECT 697.950 103.950 700.050 104.400 ;
        RECT 712.950 103.950 715.050 104.400 ;
        RECT 46.950 102.600 49.050 103.050 ;
        RECT 82.950 102.600 85.050 103.050 ;
        RECT 46.950 101.400 85.050 102.600 ;
        RECT 46.950 100.950 49.050 101.400 ;
        RECT 82.950 100.950 85.050 101.400 ;
        RECT 112.950 102.600 115.050 103.050 ;
        RECT 145.950 102.600 148.050 103.050 ;
        RECT 112.950 101.400 148.050 102.600 ;
        RECT 112.950 100.950 115.050 101.400 ;
        RECT 145.950 100.950 148.050 101.400 ;
        RECT 154.950 102.600 157.050 103.050 ;
        RECT 160.950 102.600 163.050 103.050 ;
        RECT 178.950 102.600 181.050 103.050 ;
        RECT 253.950 102.600 256.050 103.050 ;
        RECT 154.950 101.400 256.050 102.600 ;
        RECT 154.950 100.950 157.050 101.400 ;
        RECT 160.950 100.950 163.050 101.400 ;
        RECT 178.950 100.950 181.050 101.400 ;
        RECT 253.950 100.950 256.050 101.400 ;
        RECT 274.950 102.600 277.050 103.050 ;
        RECT 292.950 102.600 295.050 103.050 ;
        RECT 301.950 102.600 304.050 103.050 ;
        RECT 274.950 101.400 304.050 102.600 ;
        RECT 274.950 100.950 277.050 101.400 ;
        RECT 292.950 100.950 295.050 101.400 ;
        RECT 301.950 100.950 304.050 101.400 ;
        RECT 337.950 102.600 340.050 103.050 ;
        RECT 355.950 102.600 358.050 103.050 ;
        RECT 337.950 101.400 358.050 102.600 ;
        RECT 337.950 100.950 340.050 101.400 ;
        RECT 355.950 100.950 358.050 101.400 ;
        RECT 391.950 102.600 394.050 103.050 ;
        RECT 412.950 102.600 415.050 103.050 ;
        RECT 391.950 101.400 415.050 102.600 ;
        RECT 391.950 100.950 394.050 101.400 ;
        RECT 412.950 100.950 415.050 101.400 ;
        RECT 439.950 102.600 442.050 103.050 ;
        RECT 466.950 102.600 469.050 103.050 ;
        RECT 481.950 102.600 484.050 103.050 ;
        RECT 439.950 101.400 484.050 102.600 ;
        RECT 439.950 100.950 442.050 101.400 ;
        RECT 466.950 100.950 469.050 101.400 ;
        RECT 481.950 100.950 484.050 101.400 ;
        RECT 490.950 102.600 493.050 103.050 ;
        RECT 502.950 102.600 505.050 103.050 ;
        RECT 490.950 101.400 505.050 102.600 ;
        RECT 490.950 100.950 493.050 101.400 ;
        RECT 502.950 100.950 505.050 101.400 ;
        RECT 514.950 102.600 517.050 103.050 ;
        RECT 547.950 102.600 550.050 103.050 ;
        RECT 574.950 102.600 577.050 103.050 ;
        RECT 514.950 101.400 546.600 102.600 ;
        RECT 514.950 100.950 517.050 101.400 ;
        RECT 10.950 99.600 13.050 100.050 ;
        RECT 28.950 99.600 31.050 100.050 ;
        RECT 10.950 98.400 31.050 99.600 ;
        RECT 10.950 97.950 13.050 98.400 ;
        RECT 28.950 97.950 31.050 98.400 ;
        RECT 67.950 97.950 70.050 100.050 ;
        RECT 109.950 99.600 112.050 100.050 ;
        RECT 115.950 99.600 118.050 100.050 ;
        RECT 109.950 98.400 118.050 99.600 ;
        RECT 109.950 97.950 112.050 98.400 ;
        RECT 115.950 97.950 118.050 98.400 ;
        RECT 124.950 99.600 127.050 100.050 ;
        RECT 130.950 99.600 133.050 100.050 ;
        RECT 124.950 98.400 133.050 99.600 ;
        RECT 124.950 97.950 127.050 98.400 ;
        RECT 130.950 97.950 133.050 98.400 ;
        RECT 145.950 99.600 148.050 100.050 ;
        RECT 175.950 99.600 178.050 100.050 ;
        RECT 145.950 98.400 178.050 99.600 ;
        RECT 145.950 97.950 148.050 98.400 ;
        RECT 175.950 97.950 178.050 98.400 ;
        RECT 187.950 99.600 190.050 100.050 ;
        RECT 202.950 99.600 205.050 100.050 ;
        RECT 187.950 98.400 205.050 99.600 ;
        RECT 187.950 97.950 190.050 98.400 ;
        RECT 202.950 97.950 205.050 98.400 ;
        RECT 205.950 99.600 208.050 100.050 ;
        RECT 247.950 99.600 250.050 100.050 ;
        RECT 205.950 98.400 250.050 99.600 ;
        RECT 205.950 97.950 208.050 98.400 ;
        RECT 247.950 97.950 250.050 98.400 ;
        RECT 253.950 99.600 256.050 100.050 ;
        RECT 274.950 99.600 277.050 100.050 ;
        RECT 253.950 98.400 277.050 99.600 ;
        RECT 253.950 97.950 256.050 98.400 ;
        RECT 274.950 97.950 277.050 98.400 ;
        RECT 277.950 99.600 280.050 100.050 ;
        RECT 298.950 99.600 301.050 100.050 ;
        RECT 277.950 98.400 301.050 99.600 ;
        RECT 277.950 97.950 280.050 98.400 ;
        RECT 298.950 97.950 301.050 98.400 ;
        RECT 337.950 99.600 340.050 100.050 ;
        RECT 367.950 99.600 370.050 100.050 ;
        RECT 373.950 99.600 376.050 100.050 ;
        RECT 382.950 99.600 385.050 100.050 ;
        RECT 337.950 98.400 385.050 99.600 ;
        RECT 337.950 97.950 340.050 98.400 ;
        RECT 367.950 97.950 370.050 98.400 ;
        RECT 373.950 97.950 376.050 98.400 ;
        RECT 382.950 97.950 385.050 98.400 ;
        RECT 403.950 99.600 406.050 100.050 ;
        RECT 412.950 99.600 415.050 100.050 ;
        RECT 436.950 99.600 439.050 100.050 ;
        RECT 454.950 99.600 457.050 100.050 ;
        RECT 403.950 98.400 415.050 99.600 ;
        RECT 403.950 97.950 406.050 98.400 ;
        RECT 412.950 97.950 415.050 98.400 ;
        RECT 431.400 98.400 439.050 99.600 ;
        RECT 4.950 96.600 7.050 97.050 ;
        RECT 25.950 96.600 28.050 97.050 ;
        RECT 4.950 95.400 28.050 96.600 ;
        RECT 4.950 94.950 7.050 95.400 ;
        RECT 25.950 94.950 28.050 95.400 ;
        RECT 31.950 96.600 34.050 97.050 ;
        RECT 40.950 96.600 43.050 97.050 ;
        RECT 31.950 95.400 43.050 96.600 ;
        RECT 31.950 94.950 34.050 95.400 ;
        RECT 40.950 94.950 43.050 95.400 ;
        RECT 55.950 96.600 58.050 97.050 ;
        RECT 64.950 96.600 67.050 97.050 ;
        RECT 55.950 95.400 67.050 96.600 ;
        RECT 55.950 94.950 58.050 95.400 ;
        RECT 64.950 94.950 67.050 95.400 ;
        RECT 68.400 94.050 69.600 97.950 ;
        RECT 73.950 96.600 76.050 97.050 ;
        RECT 79.950 96.600 82.050 97.050 ;
        RECT 73.950 95.400 82.050 96.600 ;
        RECT 73.950 94.950 76.050 95.400 ;
        RECT 79.950 94.950 82.050 95.400 ;
        RECT 88.950 96.600 91.050 97.050 ;
        RECT 100.950 96.600 103.050 97.050 ;
        RECT 88.950 95.400 103.050 96.600 ;
        RECT 88.950 94.950 91.050 95.400 ;
        RECT 100.950 94.950 103.050 95.400 ;
        RECT 106.950 94.950 109.050 97.050 ;
        RECT 145.950 96.600 148.050 97.050 ;
        RECT 172.950 96.600 175.050 97.050 ;
        RECT 196.950 96.600 199.050 97.050 ;
        RECT 223.950 96.600 226.050 97.050 ;
        RECT 145.950 95.400 159.600 96.600 ;
        RECT 145.950 94.950 148.050 95.400 ;
        RECT 13.950 93.600 16.050 94.050 ;
        RECT 11.400 92.400 16.050 93.600 ;
        RECT 7.950 84.600 10.050 85.050 ;
        RECT 11.400 84.600 12.600 92.400 ;
        RECT 13.950 91.950 16.050 92.400 ;
        RECT 16.950 93.600 19.050 94.050 ;
        RECT 37.950 93.600 40.050 94.050 ;
        RECT 16.950 92.400 40.050 93.600 ;
        RECT 16.950 91.950 19.050 92.400 ;
        RECT 37.950 91.950 40.050 92.400 ;
        RECT 67.950 91.950 70.050 94.050 ;
        RECT 70.950 93.600 73.050 94.050 ;
        RECT 76.950 93.600 79.050 94.050 ;
        RECT 70.950 92.400 79.050 93.600 ;
        RECT 70.950 91.950 73.050 92.400 ;
        RECT 76.950 91.950 79.050 92.400 ;
        RECT 82.950 91.950 85.050 94.050 ;
        RECT 91.950 93.600 94.050 94.050 ;
        RECT 97.950 93.600 100.050 94.050 ;
        RECT 91.950 92.400 100.050 93.600 ;
        RECT 107.400 93.600 108.600 94.950 ;
        RECT 158.400 94.050 159.600 95.400 ;
        RECT 172.950 95.400 189.600 96.600 ;
        RECT 172.950 94.950 175.050 95.400 ;
        RECT 127.950 93.600 130.050 94.050 ;
        RECT 107.400 92.400 130.050 93.600 ;
        RECT 91.950 91.950 94.050 92.400 ;
        RECT 97.950 91.950 100.050 92.400 ;
        RECT 127.950 91.950 130.050 92.400 ;
        RECT 133.950 93.600 136.050 94.050 ;
        RECT 139.950 93.600 142.050 94.050 ;
        RECT 133.950 92.400 142.050 93.600 ;
        RECT 133.950 91.950 136.050 92.400 ;
        RECT 139.950 91.950 142.050 92.400 ;
        RECT 157.950 91.950 160.050 94.050 ;
        RECT 166.950 93.600 169.050 94.050 ;
        RECT 181.950 93.600 184.050 94.050 ;
        RECT 166.950 92.400 184.050 93.600 ;
        RECT 166.950 91.950 169.050 92.400 ;
        RECT 181.950 91.950 184.050 92.400 ;
        RECT 13.950 88.950 16.050 91.050 ;
        RECT 43.950 90.600 46.050 91.050 ;
        RECT 83.400 90.600 84.600 91.950 ;
        RECT 43.950 89.400 84.600 90.600 ;
        RECT 103.950 90.600 106.050 91.050 ;
        RECT 109.950 90.600 112.050 91.050 ;
        RECT 103.950 89.400 112.050 90.600 ;
        RECT 43.950 88.950 46.050 89.400 ;
        RECT 103.950 88.950 106.050 89.400 ;
        RECT 109.950 88.950 112.050 89.400 ;
        RECT 112.950 90.600 115.050 91.050 ;
        RECT 115.950 90.600 118.050 91.050 ;
        RECT 172.950 90.600 175.050 91.050 ;
        RECT 112.950 89.400 175.050 90.600 ;
        RECT 188.400 90.600 189.600 95.400 ;
        RECT 191.400 95.400 199.050 96.600 ;
        RECT 191.400 94.050 192.600 95.400 ;
        RECT 196.950 94.950 199.050 95.400 ;
        RECT 212.400 95.400 226.050 96.600 ;
        RECT 190.950 91.950 193.050 94.050 ;
        RECT 196.950 91.950 199.050 94.050 ;
        RECT 205.950 93.600 208.050 94.050 ;
        RECT 212.400 93.600 213.600 95.400 ;
        RECT 223.950 94.950 226.050 95.400 ;
        RECT 247.950 96.600 250.050 97.050 ;
        RECT 256.950 96.600 259.050 97.050 ;
        RECT 259.950 96.600 262.050 97.050 ;
        RECT 286.950 96.600 289.050 97.050 ;
        RECT 247.950 95.400 262.050 96.600 ;
        RECT 247.950 94.950 250.050 95.400 ;
        RECT 256.950 94.950 259.050 95.400 ;
        RECT 259.950 94.950 262.050 95.400 ;
        RECT 263.400 95.400 289.050 96.600 ;
        RECT 263.400 94.050 264.600 95.400 ;
        RECT 286.950 94.950 289.050 95.400 ;
        RECT 319.950 94.950 322.050 97.050 ;
        RECT 325.950 96.600 328.050 97.050 ;
        RECT 343.950 96.600 346.050 97.050 ;
        RECT 349.950 96.600 352.050 97.050 ;
        RECT 325.950 95.400 336.600 96.600 ;
        RECT 325.950 94.950 328.050 95.400 ;
        RECT 205.950 92.400 213.600 93.600 ;
        RECT 214.950 93.600 217.050 94.050 ;
        RECT 226.950 93.600 229.050 94.050 ;
        RECT 214.950 92.400 229.050 93.600 ;
        RECT 205.950 91.950 208.050 92.400 ;
        RECT 214.950 91.950 217.050 92.400 ;
        RECT 226.950 91.950 229.050 92.400 ;
        RECT 229.950 93.600 232.050 94.050 ;
        RECT 253.950 93.600 256.050 94.050 ;
        RECT 229.950 92.400 256.050 93.600 ;
        RECT 229.950 91.950 232.050 92.400 ;
        RECT 253.950 91.950 256.050 92.400 ;
        RECT 262.950 91.950 265.050 94.050 ;
        RECT 265.950 93.600 268.050 94.050 ;
        RECT 277.950 93.600 280.050 94.050 ;
        RECT 265.950 92.400 280.050 93.600 ;
        RECT 265.950 91.950 268.050 92.400 ;
        RECT 277.950 91.950 280.050 92.400 ;
        RECT 283.950 93.600 286.050 94.050 ;
        RECT 289.950 93.600 292.050 94.050 ;
        RECT 283.950 92.400 292.050 93.600 ;
        RECT 283.950 91.950 286.050 92.400 ;
        RECT 289.950 91.950 292.050 92.400 ;
        RECT 304.950 91.950 307.050 94.050 ;
        RECT 190.950 90.600 193.050 91.050 ;
        RECT 188.400 89.400 193.050 90.600 ;
        RECT 197.400 90.600 198.600 91.950 ;
        RECT 215.400 90.600 216.600 91.950 ;
        RECT 197.400 89.400 216.600 90.600 ;
        RECT 235.950 90.600 238.050 91.050 ;
        RECT 286.950 90.600 289.050 91.050 ;
        RECT 235.950 89.400 289.050 90.600 ;
        RECT 112.950 88.950 115.050 89.400 ;
        RECT 115.950 88.950 118.050 89.400 ;
        RECT 172.950 88.950 175.050 89.400 ;
        RECT 190.950 88.950 193.050 89.400 ;
        RECT 235.950 88.950 238.050 89.400 ;
        RECT 286.950 88.950 289.050 89.400 ;
        RECT 14.400 87.600 15.600 88.950 ;
        RECT 61.950 87.600 64.050 88.050 ;
        RECT 88.950 87.600 91.050 88.050 ;
        RECT 14.400 86.400 91.050 87.600 ;
        RECT 61.950 85.950 64.050 86.400 ;
        RECT 88.950 85.950 91.050 86.400 ;
        RECT 163.950 87.600 166.050 88.050 ;
        RECT 199.950 87.600 202.050 88.050 ;
        RECT 163.950 86.400 202.050 87.600 ;
        RECT 163.950 85.950 166.050 86.400 ;
        RECT 199.950 85.950 202.050 86.400 ;
        RECT 220.950 87.600 223.050 88.050 ;
        RECT 238.950 87.600 241.050 88.050 ;
        RECT 220.950 86.400 241.050 87.600 ;
        RECT 220.950 85.950 223.050 86.400 ;
        RECT 238.950 85.950 241.050 86.400 ;
        RECT 259.950 87.600 262.050 88.050 ;
        RECT 298.950 87.600 301.050 88.050 ;
        RECT 305.400 87.600 306.600 91.950 ;
        RECT 320.400 91.050 321.600 94.950 ;
        RECT 335.400 94.050 336.600 95.400 ;
        RECT 343.950 95.400 352.050 96.600 ;
        RECT 343.950 94.950 346.050 95.400 ;
        RECT 349.950 94.950 352.050 95.400 ;
        RECT 367.950 96.600 370.050 97.050 ;
        RECT 376.950 96.600 379.050 97.050 ;
        RECT 367.950 95.400 379.050 96.600 ;
        RECT 367.950 94.950 370.050 95.400 ;
        RECT 376.950 94.950 379.050 95.400 ;
        RECT 397.950 94.950 400.050 97.050 ;
        RECT 334.950 91.950 337.050 94.050 ;
        RECT 343.950 93.600 346.050 94.050 ;
        RECT 355.950 93.600 358.050 94.050 ;
        RECT 364.950 93.600 367.050 94.050 ;
        RECT 343.950 92.400 354.600 93.600 ;
        RECT 343.950 91.950 346.050 92.400 ;
        RECT 319.950 88.950 322.050 91.050 ;
        RECT 322.950 90.600 325.050 91.050 ;
        RECT 346.950 90.600 349.050 91.050 ;
        RECT 322.950 89.400 349.050 90.600 ;
        RECT 353.400 90.600 354.600 92.400 ;
        RECT 355.950 92.400 367.050 93.600 ;
        RECT 355.950 91.950 358.050 92.400 ;
        RECT 364.950 91.950 367.050 92.400 ;
        RECT 370.950 93.600 373.050 94.050 ;
        RECT 379.950 93.600 382.050 94.050 ;
        RECT 370.950 92.400 382.050 93.600 ;
        RECT 370.950 91.950 373.050 92.400 ;
        RECT 379.950 91.950 382.050 92.400 ;
        RECT 385.950 91.950 388.050 94.050 ;
        RECT 386.400 90.600 387.600 91.950 ;
        RECT 353.400 89.400 387.600 90.600 ;
        RECT 398.400 90.600 399.600 94.950 ;
        RECT 400.950 93.600 403.050 94.050 ;
        RECT 415.950 93.600 418.050 94.050 ;
        RECT 400.950 92.400 418.050 93.600 ;
        RECT 431.400 93.600 432.600 98.400 ;
        RECT 436.950 97.950 439.050 98.400 ;
        RECT 449.400 98.400 457.050 99.600 ;
        RECT 433.950 96.600 436.050 97.050 ;
        RECT 449.400 96.600 450.600 98.400 ;
        RECT 454.950 97.950 457.050 98.400 ;
        RECT 457.950 99.600 460.050 100.050 ;
        RECT 460.950 99.600 463.050 100.050 ;
        RECT 469.950 99.600 472.050 100.050 ;
        RECT 457.950 98.400 472.050 99.600 ;
        RECT 457.950 97.950 460.050 98.400 ;
        RECT 460.950 97.950 463.050 98.400 ;
        RECT 469.950 97.950 472.050 98.400 ;
        RECT 481.950 99.600 484.050 100.050 ;
        RECT 490.950 99.600 493.050 100.050 ;
        RECT 505.950 99.600 508.050 100.050 ;
        RECT 517.950 99.600 520.050 100.050 ;
        RECT 481.950 98.400 520.050 99.600 ;
        RECT 481.950 97.950 484.050 98.400 ;
        RECT 490.950 97.950 493.050 98.400 ;
        RECT 505.950 97.950 508.050 98.400 ;
        RECT 517.950 97.950 520.050 98.400 ;
        RECT 526.950 99.600 529.050 100.050 ;
        RECT 541.950 99.600 544.050 100.050 ;
        RECT 526.950 98.400 544.050 99.600 ;
        RECT 526.950 97.950 529.050 98.400 ;
        RECT 541.950 97.950 544.050 98.400 ;
        RECT 433.950 95.400 450.600 96.600 ;
        RECT 451.950 96.600 454.050 97.050 ;
        RECT 460.950 96.600 463.050 97.050 ;
        RECT 451.950 95.400 463.050 96.600 ;
        RECT 433.950 94.950 436.050 95.400 ;
        RECT 451.950 94.950 454.050 95.400 ;
        RECT 460.950 94.950 463.050 95.400 ;
        RECT 463.950 94.950 466.050 97.050 ;
        RECT 508.950 96.600 511.050 97.050 ;
        RECT 535.950 96.600 538.050 97.050 ;
        RECT 482.400 95.400 511.050 96.600 ;
        RECT 436.950 93.600 439.050 94.050 ;
        RECT 442.950 93.600 445.050 94.050 ;
        RECT 431.400 92.400 435.600 93.600 ;
        RECT 400.950 91.950 403.050 92.400 ;
        RECT 415.950 91.950 418.050 92.400 ;
        RECT 412.950 90.600 415.050 91.050 ;
        RECT 398.400 89.400 415.050 90.600 ;
        RECT 434.400 90.600 435.600 92.400 ;
        RECT 436.950 92.400 445.050 93.600 ;
        RECT 436.950 91.950 439.050 92.400 ;
        RECT 442.950 91.950 445.050 92.400 ;
        RECT 451.950 93.600 454.050 94.050 ;
        RECT 464.400 93.600 465.600 94.950 ;
        RECT 482.400 94.050 483.600 95.400 ;
        RECT 508.950 94.950 511.050 95.400 ;
        RECT 512.400 95.400 538.050 96.600 ;
        RECT 545.400 96.600 546.600 101.400 ;
        RECT 547.950 101.400 577.050 102.600 ;
        RECT 547.950 100.950 550.050 101.400 ;
        RECT 574.950 100.950 577.050 101.400 ;
        RECT 592.950 102.600 595.050 103.050 ;
        RECT 628.950 102.600 631.050 103.050 ;
        RECT 661.950 102.600 664.050 103.050 ;
        RECT 676.950 102.600 679.050 103.050 ;
        RECT 592.950 101.400 679.050 102.600 ;
        RECT 592.950 100.950 595.050 101.400 ;
        RECT 628.950 100.950 631.050 101.400 ;
        RECT 661.950 100.950 664.050 101.400 ;
        RECT 676.950 100.950 679.050 101.400 ;
        RECT 682.950 102.600 685.050 103.050 ;
        RECT 745.950 102.600 748.050 103.050 ;
        RECT 682.950 101.400 748.050 102.600 ;
        RECT 682.950 100.950 685.050 101.400 ;
        RECT 745.950 100.950 748.050 101.400 ;
        RECT 556.950 99.600 559.050 100.050 ;
        RECT 565.950 99.600 568.050 100.050 ;
        RECT 556.950 98.400 568.050 99.600 ;
        RECT 556.950 97.950 559.050 98.400 ;
        RECT 565.950 97.950 568.050 98.400 ;
        RECT 571.950 99.600 574.050 100.050 ;
        RECT 577.950 99.600 580.050 100.050 ;
        RECT 571.950 98.400 580.050 99.600 ;
        RECT 571.950 97.950 574.050 98.400 ;
        RECT 577.950 97.950 580.050 98.400 ;
        RECT 580.950 99.600 583.050 100.050 ;
        RECT 598.950 99.600 601.050 100.050 ;
        RECT 625.950 99.600 628.050 100.050 ;
        RECT 580.950 98.400 597.600 99.600 ;
        RECT 580.950 97.950 583.050 98.400 ;
        RECT 596.400 97.050 597.600 98.400 ;
        RECT 598.950 98.400 628.050 99.600 ;
        RECT 598.950 97.950 601.050 98.400 ;
        RECT 625.950 97.950 628.050 98.400 ;
        RECT 631.950 99.600 634.050 100.050 ;
        RECT 640.950 99.600 643.050 100.050 ;
        RECT 667.950 99.600 670.050 100.050 ;
        RECT 673.950 99.600 676.050 100.050 ;
        RECT 727.950 99.600 730.050 100.050 ;
        RECT 631.950 98.400 639.600 99.600 ;
        RECT 631.950 97.950 634.050 98.400 ;
        RECT 562.950 96.600 565.050 97.050 ;
        RECT 595.950 96.600 598.050 97.050 ;
        RECT 613.950 96.600 616.050 97.050 ;
        RECT 545.400 95.400 573.600 96.600 ;
        RECT 512.400 94.050 513.600 95.400 ;
        RECT 535.950 94.950 538.050 95.400 ;
        RECT 554.400 94.050 555.600 95.400 ;
        RECT 562.950 94.950 565.050 95.400 ;
        RECT 451.950 92.400 465.600 93.600 ;
        RECT 466.950 93.600 469.050 94.050 ;
        RECT 478.950 93.600 481.050 94.050 ;
        RECT 466.950 92.400 481.050 93.600 ;
        RECT 451.950 91.950 454.050 92.400 ;
        RECT 466.950 91.950 469.050 92.400 ;
        RECT 478.950 91.950 481.050 92.400 ;
        RECT 481.950 91.950 484.050 94.050 ;
        RECT 511.950 91.950 514.050 94.050 ;
        RECT 523.950 93.600 526.050 94.050 ;
        RECT 538.950 93.600 541.050 94.050 ;
        RECT 523.950 92.400 541.050 93.600 ;
        RECT 523.950 91.950 526.050 92.400 ;
        RECT 538.950 91.950 541.050 92.400 ;
        RECT 553.950 91.950 556.050 94.050 ;
        RECT 559.950 93.600 562.050 94.050 ;
        RECT 568.950 93.600 571.050 94.050 ;
        RECT 559.950 92.400 571.050 93.600 ;
        RECT 572.400 93.600 573.600 95.400 ;
        RECT 595.950 95.400 616.050 96.600 ;
        RECT 595.950 94.950 598.050 95.400 ;
        RECT 613.950 94.950 616.050 95.400 ;
        RECT 628.950 96.600 631.050 97.050 ;
        RECT 628.950 95.400 636.600 96.600 ;
        RECT 628.950 94.950 631.050 95.400 ;
        RECT 635.400 94.050 636.600 95.400 ;
        RECT 638.400 94.050 639.600 98.400 ;
        RECT 640.950 98.400 654.600 99.600 ;
        RECT 640.950 97.950 643.050 98.400 ;
        RECT 653.400 96.600 654.600 98.400 ;
        RECT 667.950 98.400 676.050 99.600 ;
        RECT 667.950 97.950 670.050 98.400 ;
        RECT 673.950 97.950 676.050 98.400 ;
        RECT 719.400 98.400 730.050 99.600 ;
        RECT 715.950 96.600 718.050 97.050 ;
        RECT 653.400 95.400 681.600 96.600 ;
        RECT 653.400 94.050 654.600 95.400 ;
        RECT 680.400 94.050 681.600 95.400 ;
        RECT 713.400 95.400 718.050 96.600 ;
        RECT 592.950 93.600 595.050 94.050 ;
        RECT 572.400 92.400 595.050 93.600 ;
        RECT 559.950 91.950 562.050 92.400 ;
        RECT 568.950 91.950 571.050 92.400 ;
        RECT 592.950 91.950 595.050 92.400 ;
        RECT 607.950 93.600 610.050 94.050 ;
        RECT 628.950 93.600 631.050 94.050 ;
        RECT 607.950 92.400 631.050 93.600 ;
        RECT 607.950 91.950 610.050 92.400 ;
        RECT 628.950 91.950 631.050 92.400 ;
        RECT 634.950 91.950 637.050 94.050 ;
        RECT 637.950 91.950 640.050 94.050 ;
        RECT 652.950 93.600 655.050 94.050 ;
        RECT 664.950 93.600 667.050 94.050 ;
        RECT 652.950 92.400 667.050 93.600 ;
        RECT 652.950 91.950 655.050 92.400 ;
        RECT 664.950 91.950 667.050 92.400 ;
        RECT 670.950 91.950 673.050 94.050 ;
        RECT 679.950 91.950 682.050 94.050 ;
        RECT 694.950 93.600 697.050 94.050 ;
        RECT 709.950 93.600 712.050 94.050 ;
        RECT 694.950 92.400 712.050 93.600 ;
        RECT 694.950 91.950 697.050 92.400 ;
        RECT 709.950 91.950 712.050 92.400 ;
        RECT 439.950 90.600 442.050 91.050 ;
        RECT 434.400 89.400 442.050 90.600 ;
        RECT 322.950 88.950 325.050 89.400 ;
        RECT 346.950 88.950 349.050 89.400 ;
        RECT 412.950 88.950 415.050 89.400 ;
        RECT 439.950 88.950 442.050 89.400 ;
        RECT 442.950 90.600 445.050 91.050 ;
        RECT 448.950 90.600 451.050 91.050 ;
        RECT 442.950 89.400 451.050 90.600 ;
        RECT 442.950 88.950 445.050 89.400 ;
        RECT 448.950 88.950 451.050 89.400 ;
        RECT 454.950 90.600 457.050 91.050 ;
        RECT 460.950 90.600 463.050 91.050 ;
        RECT 454.950 89.400 463.050 90.600 ;
        RECT 454.950 88.950 457.050 89.400 ;
        RECT 460.950 88.950 463.050 89.400 ;
        RECT 493.950 88.950 496.050 91.050 ;
        RECT 514.950 90.600 517.050 91.050 ;
        RECT 526.950 90.600 529.050 91.050 ;
        RECT 514.950 89.400 529.050 90.600 ;
        RECT 514.950 88.950 517.050 89.400 ;
        RECT 526.950 88.950 529.050 89.400 ;
        RECT 532.950 90.600 535.050 91.050 ;
        RECT 544.950 90.600 547.050 91.050 ;
        RECT 532.950 89.400 547.050 90.600 ;
        RECT 532.950 88.950 535.050 89.400 ;
        RECT 544.950 88.950 547.050 89.400 ;
        RECT 565.950 88.950 568.050 91.050 ;
        RECT 595.950 90.600 598.050 91.050 ;
        RECT 604.950 90.600 607.050 91.050 ;
        RECT 595.950 89.400 607.050 90.600 ;
        RECT 595.950 88.950 598.050 89.400 ;
        RECT 604.950 88.950 607.050 89.400 ;
        RECT 625.950 90.600 628.050 91.050 ;
        RECT 640.950 90.600 643.050 91.050 ;
        RECT 671.400 90.600 672.600 91.950 ;
        RECT 713.400 90.600 714.600 95.400 ;
        RECT 715.950 94.950 718.050 95.400 ;
        RECT 719.400 93.600 720.600 98.400 ;
        RECT 727.950 97.950 730.050 98.400 ;
        RECT 733.950 99.600 736.050 100.050 ;
        RECT 739.950 99.600 742.050 100.050 ;
        RECT 733.950 98.400 742.050 99.600 ;
        RECT 733.950 97.950 736.050 98.400 ;
        RECT 739.950 97.950 742.050 98.400 ;
        RECT 721.950 96.600 724.050 97.050 ;
        RECT 727.950 96.600 730.050 97.050 ;
        RECT 739.950 96.600 742.050 97.050 ;
        RECT 721.950 95.400 730.050 96.600 ;
        RECT 721.950 94.950 724.050 95.400 ;
        RECT 727.950 94.950 730.050 95.400 ;
        RECT 734.400 95.400 742.050 96.600 ;
        RECT 734.400 93.600 735.600 95.400 ;
        RECT 739.950 94.950 742.050 95.400 ;
        RECT 625.950 89.400 714.600 90.600 ;
        RECT 716.400 92.400 720.600 93.600 ;
        RECT 728.400 92.400 735.600 93.600 ;
        RECT 736.950 93.600 739.050 94.050 ;
        RECT 745.950 93.600 748.050 94.050 ;
        RECT 736.950 92.400 748.050 93.600 ;
        RECT 625.950 88.950 628.050 89.400 ;
        RECT 640.950 88.950 643.050 89.400 ;
        RECT 328.950 87.600 331.050 88.050 ;
        RECT 259.950 86.400 331.050 87.600 ;
        RECT 259.950 85.950 262.050 86.400 ;
        RECT 298.950 85.950 301.050 86.400 ;
        RECT 328.950 85.950 331.050 86.400 ;
        RECT 358.950 87.600 361.050 88.050 ;
        RECT 430.950 87.600 433.050 88.050 ;
        RECT 445.950 87.600 448.050 88.050 ;
        RECT 358.950 86.400 448.050 87.600 ;
        RECT 358.950 85.950 361.050 86.400 ;
        RECT 430.950 85.950 433.050 86.400 ;
        RECT 445.950 85.950 448.050 86.400 ;
        RECT 457.950 87.600 460.050 88.050 ;
        RECT 494.400 87.600 495.600 88.950 ;
        RECT 544.950 87.600 547.050 88.050 ;
        RECT 457.950 86.400 547.050 87.600 ;
        RECT 457.950 85.950 460.050 86.400 ;
        RECT 544.950 85.950 547.050 86.400 ;
        RECT 562.950 87.600 565.050 88.050 ;
        RECT 566.400 87.600 567.600 88.950 ;
        RECT 716.400 88.050 717.600 92.400 ;
        RECT 718.950 90.600 721.050 91.050 ;
        RECT 728.400 90.600 729.600 92.400 ;
        RECT 736.950 91.950 739.050 92.400 ;
        RECT 745.950 91.950 748.050 92.400 ;
        RECT 718.950 89.400 729.600 90.600 ;
        RECT 730.950 90.600 733.050 91.050 ;
        RECT 742.950 90.600 745.050 91.050 ;
        RECT 730.950 89.400 745.050 90.600 ;
        RECT 718.950 88.950 721.050 89.400 ;
        RECT 730.950 88.950 733.050 89.400 ;
        RECT 742.950 88.950 745.050 89.400 ;
        RECT 562.950 86.400 567.600 87.600 ;
        RECT 598.950 87.600 601.050 88.050 ;
        RECT 610.950 87.600 613.050 88.050 ;
        RECT 619.950 87.600 622.050 88.050 ;
        RECT 598.950 86.400 622.050 87.600 ;
        RECT 562.950 85.950 565.050 86.400 ;
        RECT 598.950 85.950 601.050 86.400 ;
        RECT 610.950 85.950 613.050 86.400 ;
        RECT 619.950 85.950 622.050 86.400 ;
        RECT 628.950 87.600 631.050 88.050 ;
        RECT 658.950 87.600 661.050 88.050 ;
        RECT 688.950 87.600 691.050 88.050 ;
        RECT 628.950 86.400 691.050 87.600 ;
        RECT 628.950 85.950 631.050 86.400 ;
        RECT 658.950 85.950 661.050 86.400 ;
        RECT 688.950 85.950 691.050 86.400 ;
        RECT 715.950 85.950 718.050 88.050 ;
        RECT 7.950 83.400 12.600 84.600 ;
        RECT 64.950 84.600 67.050 85.050 ;
        RECT 73.950 84.600 76.050 85.050 ;
        RECT 64.950 83.400 76.050 84.600 ;
        RECT 7.950 82.950 10.050 83.400 ;
        RECT 64.950 82.950 67.050 83.400 ;
        RECT 73.950 82.950 76.050 83.400 ;
        RECT 211.950 84.600 214.050 85.050 ;
        RECT 256.950 84.600 259.050 85.050 ;
        RECT 211.950 83.400 259.050 84.600 ;
        RECT 211.950 82.950 214.050 83.400 ;
        RECT 256.950 82.950 259.050 83.400 ;
        RECT 397.950 84.600 400.050 85.050 ;
        RECT 424.950 84.600 427.050 85.050 ;
        RECT 442.950 84.600 445.050 85.050 ;
        RECT 397.950 83.400 445.050 84.600 ;
        RECT 397.950 82.950 400.050 83.400 ;
        RECT 424.950 82.950 427.050 83.400 ;
        RECT 442.950 82.950 445.050 83.400 ;
        RECT 472.950 84.600 475.050 85.050 ;
        RECT 475.950 84.600 478.050 85.050 ;
        RECT 499.950 84.600 502.050 85.050 ;
        RECT 586.950 84.600 589.050 85.050 ;
        RECT 472.950 83.400 589.050 84.600 ;
        RECT 472.950 82.950 475.050 83.400 ;
        RECT 475.950 82.950 478.050 83.400 ;
        RECT 499.950 82.950 502.050 83.400 ;
        RECT 586.950 82.950 589.050 83.400 ;
        RECT 703.950 84.600 706.050 85.050 ;
        RECT 748.950 84.600 751.050 85.050 ;
        RECT 703.950 83.400 751.050 84.600 ;
        RECT 703.950 82.950 706.050 83.400 ;
        RECT 748.950 82.950 751.050 83.400 ;
        RECT 1.950 81.600 4.050 82.050 ;
        RECT 22.950 81.600 25.050 82.050 ;
        RECT 52.950 81.600 55.050 82.050 ;
        RECT 1.950 80.400 55.050 81.600 ;
        RECT 1.950 79.950 4.050 80.400 ;
        RECT 22.950 79.950 25.050 80.400 ;
        RECT 52.950 79.950 55.050 80.400 ;
        RECT 334.950 81.600 337.050 82.050 ;
        RECT 409.950 81.600 412.050 82.050 ;
        RECT 334.950 80.400 412.050 81.600 ;
        RECT 334.950 79.950 337.050 80.400 ;
        RECT 409.950 79.950 412.050 80.400 ;
        RECT 415.950 81.600 418.050 82.050 ;
        RECT 481.950 81.600 484.050 82.050 ;
        RECT 415.950 80.400 484.050 81.600 ;
        RECT 415.950 79.950 418.050 80.400 ;
        RECT 481.950 79.950 484.050 80.400 ;
        RECT 1.950 78.600 4.050 79.050 ;
        RECT 7.950 78.600 10.050 79.050 ;
        RECT 1.950 77.400 10.050 78.600 ;
        RECT 1.950 76.950 4.050 77.400 ;
        RECT 7.950 76.950 10.050 77.400 ;
        RECT 31.950 78.600 34.050 79.050 ;
        RECT 103.950 78.600 106.050 79.050 ;
        RECT 31.950 77.400 106.050 78.600 ;
        RECT 31.950 76.950 34.050 77.400 ;
        RECT 103.950 76.950 106.050 77.400 ;
        RECT 121.950 78.600 124.050 79.050 ;
        RECT 160.950 78.600 163.050 79.050 ;
        RECT 121.950 77.400 163.050 78.600 ;
        RECT 121.950 76.950 124.050 77.400 ;
        RECT 160.950 76.950 163.050 77.400 ;
        RECT 460.950 78.600 463.050 79.050 ;
        RECT 514.950 78.600 517.050 79.050 ;
        RECT 541.950 78.600 544.050 79.050 ;
        RECT 460.950 77.400 544.050 78.600 ;
        RECT 460.950 76.950 463.050 77.400 ;
        RECT 514.950 76.950 517.050 77.400 ;
        RECT 541.950 76.950 544.050 77.400 ;
        RECT 40.950 75.600 43.050 76.050 ;
        RECT 67.950 75.600 70.050 76.050 ;
        RECT 40.950 74.400 70.050 75.600 ;
        RECT 40.950 73.950 43.050 74.400 ;
        RECT 67.950 73.950 70.050 74.400 ;
        RECT 421.950 75.600 424.050 76.050 ;
        RECT 571.950 75.600 574.050 76.050 ;
        RECT 421.950 74.400 574.050 75.600 ;
        RECT 421.950 73.950 424.050 74.400 ;
        RECT 571.950 73.950 574.050 74.400 ;
        RECT 85.950 72.600 88.050 73.050 ;
        RECT 133.950 72.600 136.050 73.050 ;
        RECT 85.950 71.400 136.050 72.600 ;
        RECT 85.950 70.950 88.050 71.400 ;
        RECT 133.950 70.950 136.050 71.400 ;
        RECT 307.950 72.600 310.050 73.050 ;
        RECT 316.950 72.600 319.050 73.050 ;
        RECT 307.950 71.400 319.050 72.600 ;
        RECT 307.950 70.950 310.050 71.400 ;
        RECT 316.950 70.950 319.050 71.400 ;
        RECT 382.950 72.600 385.050 73.050 ;
        RECT 391.950 72.600 394.050 73.050 ;
        RECT 382.950 71.400 394.050 72.600 ;
        RECT 382.950 70.950 385.050 71.400 ;
        RECT 391.950 70.950 394.050 71.400 ;
        RECT 463.950 72.600 466.050 73.050 ;
        RECT 637.950 72.600 640.050 73.050 ;
        RECT 463.950 71.400 640.050 72.600 ;
        RECT 463.950 70.950 466.050 71.400 ;
        RECT 637.950 70.950 640.050 71.400 ;
        RECT 694.950 72.600 697.050 73.050 ;
        RECT 700.950 72.600 703.050 73.050 ;
        RECT 694.950 71.400 703.050 72.600 ;
        RECT 694.950 70.950 697.050 71.400 ;
        RECT 700.950 70.950 703.050 71.400 ;
        RECT 106.950 69.600 109.050 70.050 ;
        RECT 151.950 69.600 154.050 70.050 ;
        RECT 106.950 68.400 154.050 69.600 ;
        RECT 106.950 67.950 109.050 68.400 ;
        RECT 151.950 67.950 154.050 68.400 ;
        RECT 226.950 69.600 229.050 70.050 ;
        RECT 244.950 69.600 247.050 70.050 ;
        RECT 250.950 69.600 253.050 70.050 ;
        RECT 226.950 68.400 253.050 69.600 ;
        RECT 226.950 67.950 229.050 68.400 ;
        RECT 244.950 67.950 247.050 68.400 ;
        RECT 250.950 67.950 253.050 68.400 ;
        RECT 253.950 69.600 256.050 70.050 ;
        RECT 262.950 69.600 265.050 70.050 ;
        RECT 253.950 68.400 265.050 69.600 ;
        RECT 253.950 67.950 256.050 68.400 ;
        RECT 262.950 67.950 265.050 68.400 ;
        RECT 304.950 69.600 307.050 70.050 ;
        RECT 334.950 69.600 337.050 70.050 ;
        RECT 304.950 68.400 337.050 69.600 ;
        RECT 304.950 67.950 307.050 68.400 ;
        RECT 334.950 67.950 337.050 68.400 ;
        RECT 346.950 69.600 349.050 70.050 ;
        RECT 409.950 69.600 412.050 70.050 ;
        RECT 346.950 68.400 412.050 69.600 ;
        RECT 346.950 67.950 349.050 68.400 ;
        RECT 409.950 67.950 412.050 68.400 ;
        RECT 418.950 69.600 421.050 70.050 ;
        RECT 427.950 69.600 430.050 70.050 ;
        RECT 466.950 69.600 469.050 70.050 ;
        RECT 658.950 69.600 661.050 70.050 ;
        RECT 418.950 68.400 661.050 69.600 ;
        RECT 418.950 67.950 421.050 68.400 ;
        RECT 427.950 67.950 430.050 68.400 ;
        RECT 466.950 67.950 469.050 68.400 ;
        RECT 658.950 67.950 661.050 68.400 ;
        RECT 82.950 66.600 85.050 67.050 ;
        RECT 142.950 66.600 145.050 67.050 ;
        RECT 82.950 65.400 145.050 66.600 ;
        RECT 82.950 64.950 85.050 65.400 ;
        RECT 142.950 64.950 145.050 65.400 ;
        RECT 151.950 66.600 154.050 67.050 ;
        RECT 169.950 66.600 172.050 67.050 ;
        RECT 151.950 65.400 172.050 66.600 ;
        RECT 151.950 64.950 154.050 65.400 ;
        RECT 169.950 64.950 172.050 65.400 ;
        RECT 538.950 66.600 541.050 67.050 ;
        RECT 571.950 66.600 574.050 67.050 ;
        RECT 538.950 65.400 574.050 66.600 ;
        RECT 538.950 64.950 541.050 65.400 ;
        RECT 571.950 64.950 574.050 65.400 ;
        RECT 586.950 66.600 589.050 67.050 ;
        RECT 604.950 66.600 607.050 67.050 ;
        RECT 586.950 65.400 607.050 66.600 ;
        RECT 586.950 64.950 589.050 65.400 ;
        RECT 604.950 64.950 607.050 65.400 ;
        RECT 13.950 63.600 16.050 64.050 ;
        RECT 43.950 63.600 46.050 64.050 ;
        RECT 130.950 63.600 133.050 64.050 ;
        RECT 184.950 63.600 187.050 64.050 ;
        RECT 13.950 62.400 187.050 63.600 ;
        RECT 13.950 61.950 16.050 62.400 ;
        RECT 43.950 61.950 46.050 62.400 ;
        RECT 130.950 61.950 133.050 62.400 ;
        RECT 184.950 61.950 187.050 62.400 ;
        RECT 250.950 63.600 253.050 64.050 ;
        RECT 268.950 63.600 271.050 64.050 ;
        RECT 250.950 62.400 271.050 63.600 ;
        RECT 250.950 61.950 253.050 62.400 ;
        RECT 268.950 61.950 271.050 62.400 ;
        RECT 376.950 63.600 379.050 64.050 ;
        RECT 385.950 63.600 388.050 64.050 ;
        RECT 376.950 62.400 388.050 63.600 ;
        RECT 376.950 61.950 379.050 62.400 ;
        RECT 385.950 61.950 388.050 62.400 ;
        RECT 424.950 63.600 427.050 64.050 ;
        RECT 481.950 63.600 484.050 64.050 ;
        RECT 424.950 62.400 484.050 63.600 ;
        RECT 424.950 61.950 427.050 62.400 ;
        RECT 481.950 61.950 484.050 62.400 ;
        RECT 547.950 63.600 550.050 64.050 ;
        RECT 583.950 63.600 586.050 64.050 ;
        RECT 547.950 62.400 586.050 63.600 ;
        RECT 547.950 61.950 550.050 62.400 ;
        RECT 583.950 61.950 586.050 62.400 ;
        RECT 4.950 60.600 7.050 61.050 ;
        RECT 16.950 60.600 19.050 61.050 ;
        RECT 46.950 60.600 49.050 61.050 ;
        RECT 52.950 60.600 55.050 61.050 ;
        RECT 58.950 60.600 61.050 61.050 ;
        RECT 139.950 60.600 142.050 61.050 ;
        RECT 4.950 59.400 45.600 60.600 ;
        RECT 4.950 58.950 7.050 59.400 ;
        RECT 16.950 58.950 19.050 59.400 ;
        RECT 10.950 57.600 13.050 58.050 ;
        RECT 22.950 57.600 25.050 58.050 ;
        RECT 40.950 57.600 43.050 58.050 ;
        RECT 10.950 56.400 25.050 57.600 ;
        RECT 10.950 55.950 13.050 56.400 ;
        RECT 22.950 55.950 25.050 56.400 ;
        RECT 26.400 56.400 43.050 57.600 ;
        RECT 44.400 57.600 45.600 59.400 ;
        RECT 46.950 59.400 61.050 60.600 ;
        RECT 46.950 58.950 49.050 59.400 ;
        RECT 52.950 58.950 55.050 59.400 ;
        RECT 58.950 58.950 61.050 59.400 ;
        RECT 95.400 59.400 142.050 60.600 ;
        RECT 95.400 57.600 96.600 59.400 ;
        RECT 139.950 58.950 142.050 59.400 ;
        RECT 388.950 60.600 391.050 61.050 ;
        RECT 424.950 60.600 427.050 61.050 ;
        RECT 388.950 59.400 427.050 60.600 ;
        RECT 388.950 58.950 391.050 59.400 ;
        RECT 424.950 58.950 427.050 59.400 ;
        RECT 439.950 60.600 442.050 61.050 ;
        RECT 586.950 60.600 589.050 61.050 ;
        RECT 439.950 59.400 589.050 60.600 ;
        RECT 439.950 58.950 442.050 59.400 ;
        RECT 586.950 58.950 589.050 59.400 ;
        RECT 640.950 60.600 643.050 61.050 ;
        RECT 649.950 60.600 652.050 61.050 ;
        RECT 640.950 59.400 652.050 60.600 ;
        RECT 640.950 58.950 643.050 59.400 ;
        RECT 649.950 58.950 652.050 59.400 ;
        RECT 691.950 60.600 694.050 61.050 ;
        RECT 706.950 60.600 709.050 61.050 ;
        RECT 691.950 59.400 709.050 60.600 ;
        RECT 691.950 58.950 694.050 59.400 ;
        RECT 706.950 58.950 709.050 59.400 ;
        RECT 724.950 58.950 727.050 61.050 ;
        RECT 745.950 60.600 748.050 61.050 ;
        RECT 740.400 59.400 748.050 60.600 ;
        RECT 44.400 56.400 96.600 57.600 ;
        RECT 109.950 57.600 112.050 58.050 ;
        RECT 118.950 57.600 121.050 58.050 ;
        RECT 109.950 56.400 121.050 57.600 ;
        RECT 26.400 55.050 27.600 56.400 ;
        RECT 40.950 55.950 43.050 56.400 ;
        RECT 109.950 55.950 112.050 56.400 ;
        RECT 118.950 55.950 121.050 56.400 ;
        RECT 133.950 57.600 136.050 58.050 ;
        RECT 139.950 57.600 142.050 58.050 ;
        RECT 145.950 57.600 148.050 58.050 ;
        RECT 133.950 56.400 138.600 57.600 ;
        RECT 133.950 55.950 136.050 56.400 ;
        RECT 1.950 54.600 4.050 55.050 ;
        RECT 7.950 54.600 10.050 55.050 ;
        RECT 1.950 53.400 10.050 54.600 ;
        RECT 1.950 52.950 4.050 53.400 ;
        RECT 7.950 52.950 10.050 53.400 ;
        RECT 25.950 52.950 28.050 55.050 ;
        RECT 31.950 52.950 34.050 55.050 ;
        RECT 37.950 54.600 40.050 55.050 ;
        RECT 49.950 54.600 52.050 55.050 ;
        RECT 37.950 53.400 52.050 54.600 ;
        RECT 37.950 52.950 40.050 53.400 ;
        RECT 49.950 52.950 52.050 53.400 ;
        RECT 61.950 54.600 64.050 55.050 ;
        RECT 67.950 54.600 70.050 55.050 ;
        RECT 61.950 53.400 70.050 54.600 ;
        RECT 61.950 52.950 64.050 53.400 ;
        RECT 67.950 52.950 70.050 53.400 ;
        RECT 73.950 54.600 76.050 55.050 ;
        RECT 88.950 54.600 91.050 55.050 ;
        RECT 73.950 53.400 91.050 54.600 ;
        RECT 73.950 52.950 76.050 53.400 ;
        RECT 88.950 52.950 91.050 53.400 ;
        RECT 100.950 52.950 103.050 55.050 ;
        RECT 103.950 52.950 106.050 55.050 ;
        RECT 106.950 54.600 109.050 55.050 ;
        RECT 137.400 54.600 138.600 56.400 ;
        RECT 139.950 56.400 148.050 57.600 ;
        RECT 139.950 55.950 142.050 56.400 ;
        RECT 145.950 55.950 148.050 56.400 ;
        RECT 169.950 57.600 172.050 58.050 ;
        RECT 178.950 57.600 181.050 58.050 ;
        RECT 199.950 57.600 202.050 58.050 ;
        RECT 214.950 57.600 217.050 58.050 ;
        RECT 169.950 56.400 217.050 57.600 ;
        RECT 169.950 55.950 172.050 56.400 ;
        RECT 178.950 55.950 181.050 56.400 ;
        RECT 199.950 55.950 202.050 56.400 ;
        RECT 214.950 55.950 217.050 56.400 ;
        RECT 265.950 57.600 268.050 58.050 ;
        RECT 268.950 57.600 271.050 58.050 ;
        RECT 280.950 57.600 283.050 58.050 ;
        RECT 265.950 56.400 283.050 57.600 ;
        RECT 265.950 55.950 268.050 56.400 ;
        RECT 268.950 55.950 271.050 56.400 ;
        RECT 280.950 55.950 283.050 56.400 ;
        RECT 292.950 57.600 295.050 58.050 ;
        RECT 304.950 57.600 307.050 58.050 ;
        RECT 292.950 56.400 307.050 57.600 ;
        RECT 292.950 55.950 295.050 56.400 ;
        RECT 304.950 55.950 307.050 56.400 ;
        RECT 313.950 57.600 316.050 58.050 ;
        RECT 328.950 57.600 331.050 58.050 ;
        RECT 313.950 56.400 331.050 57.600 ;
        RECT 313.950 55.950 316.050 56.400 ;
        RECT 328.950 55.950 331.050 56.400 ;
        RECT 364.950 57.600 367.050 58.050 ;
        RECT 376.950 57.600 379.050 58.050 ;
        RECT 385.950 57.600 388.050 58.050 ;
        RECT 409.950 57.600 412.050 58.050 ;
        RECT 364.950 56.400 384.600 57.600 ;
        RECT 364.950 55.950 367.050 56.400 ;
        RECT 376.950 55.950 379.050 56.400 ;
        RECT 142.950 54.600 145.050 55.050 ;
        RECT 106.950 53.400 117.600 54.600 ;
        RECT 137.400 53.400 145.050 54.600 ;
        RECT 106.950 52.950 109.050 53.400 ;
        RECT 1.950 51.600 4.050 52.050 ;
        RECT 19.950 51.600 22.050 52.050 ;
        RECT 1.950 50.400 22.050 51.600 ;
        RECT 1.950 49.950 4.050 50.400 ;
        RECT 19.950 49.950 22.050 50.400 ;
        RECT 25.950 51.600 28.050 52.050 ;
        RECT 32.400 51.600 33.600 52.950 ;
        RECT 25.950 50.400 33.600 51.600 ;
        RECT 34.950 51.600 37.050 52.050 ;
        RECT 40.950 51.600 43.050 52.050 ;
        RECT 34.950 50.400 43.050 51.600 ;
        RECT 25.950 49.950 28.050 50.400 ;
        RECT 34.950 49.950 37.050 50.400 ;
        RECT 40.950 49.950 43.050 50.400 ;
        RECT 58.950 51.600 61.050 52.050 ;
        RECT 94.950 51.600 97.050 52.050 ;
        RECT 58.950 50.400 97.050 51.600 ;
        RECT 58.950 49.950 61.050 50.400 ;
        RECT 94.950 49.950 97.050 50.400 ;
        RECT 101.400 49.050 102.600 52.950 ;
        RECT 104.400 51.600 105.600 52.950 ;
        RECT 116.400 52.050 117.600 53.400 ;
        RECT 142.950 52.950 145.050 53.400 ;
        RECT 175.950 54.600 178.050 55.050 ;
        RECT 181.950 54.600 184.050 55.050 ;
        RECT 175.950 53.400 184.050 54.600 ;
        RECT 175.950 52.950 178.050 53.400 ;
        RECT 181.950 52.950 184.050 53.400 ;
        RECT 202.950 54.600 205.050 55.050 ;
        RECT 289.950 54.600 292.050 55.050 ;
        RECT 202.950 53.400 292.050 54.600 ;
        RECT 202.950 52.950 205.050 53.400 ;
        RECT 289.950 52.950 292.050 53.400 ;
        RECT 295.950 54.600 298.050 55.050 ;
        RECT 301.950 54.600 304.050 55.050 ;
        RECT 295.950 53.400 304.050 54.600 ;
        RECT 295.950 52.950 298.050 53.400 ;
        RECT 301.950 52.950 304.050 53.400 ;
        RECT 307.950 52.950 310.050 55.050 ;
        RECT 319.950 52.950 322.050 55.050 ;
        RECT 322.950 52.950 325.050 55.050 ;
        RECT 337.950 54.600 340.050 55.050 ;
        RECT 355.950 54.600 358.050 55.050 ;
        RECT 337.950 53.400 358.050 54.600 ;
        RECT 337.950 52.950 340.050 53.400 ;
        RECT 355.950 52.950 358.050 53.400 ;
        RECT 367.950 54.600 370.050 55.050 ;
        RECT 373.950 54.600 376.050 55.050 ;
        RECT 367.950 53.400 376.050 54.600 ;
        RECT 383.400 54.600 384.600 56.400 ;
        RECT 385.950 56.400 412.050 57.600 ;
        RECT 385.950 55.950 388.050 56.400 ;
        RECT 409.950 55.950 412.050 56.400 ;
        RECT 412.950 57.600 415.050 58.050 ;
        RECT 421.950 57.600 424.050 58.050 ;
        RECT 433.950 57.600 436.050 58.050 ;
        RECT 412.950 56.400 436.050 57.600 ;
        RECT 412.950 55.950 415.050 56.400 ;
        RECT 421.950 55.950 424.050 56.400 ;
        RECT 433.950 55.950 436.050 56.400 ;
        RECT 454.950 57.600 457.050 58.050 ;
        RECT 469.950 57.600 472.050 58.050 ;
        RECT 454.950 56.400 472.050 57.600 ;
        RECT 454.950 55.950 457.050 56.400 ;
        RECT 469.950 55.950 472.050 56.400 ;
        RECT 475.950 57.600 478.050 58.050 ;
        RECT 481.950 57.600 484.050 58.050 ;
        RECT 487.950 57.600 490.050 58.050 ;
        RECT 475.950 56.400 490.050 57.600 ;
        RECT 475.950 55.950 478.050 56.400 ;
        RECT 481.950 55.950 484.050 56.400 ;
        RECT 487.950 55.950 490.050 56.400 ;
        RECT 493.950 57.600 496.050 58.050 ;
        RECT 496.950 57.600 499.050 58.050 ;
        RECT 499.950 57.600 502.050 58.050 ;
        RECT 493.950 56.400 502.050 57.600 ;
        RECT 493.950 55.950 496.050 56.400 ;
        RECT 496.950 55.950 499.050 56.400 ;
        RECT 499.950 55.950 502.050 56.400 ;
        RECT 502.950 57.600 505.050 58.050 ;
        RECT 511.950 57.600 514.050 58.050 ;
        RECT 502.950 56.400 514.050 57.600 ;
        RECT 502.950 55.950 505.050 56.400 ;
        RECT 511.950 55.950 514.050 56.400 ;
        RECT 523.950 57.600 526.050 58.050 ;
        RECT 532.950 57.600 535.050 58.050 ;
        RECT 553.950 57.600 556.050 58.050 ;
        RECT 559.950 57.600 562.050 58.050 ;
        RECT 523.950 56.400 546.600 57.600 ;
        RECT 523.950 55.950 526.050 56.400 ;
        RECT 532.950 55.950 535.050 56.400 ;
        RECT 545.400 55.050 546.600 56.400 ;
        RECT 553.950 56.400 562.050 57.600 ;
        RECT 553.950 55.950 556.050 56.400 ;
        RECT 559.950 55.950 562.050 56.400 ;
        RECT 562.950 57.600 565.050 58.050 ;
        RECT 562.950 56.400 567.600 57.600 ;
        RECT 562.950 55.950 565.050 56.400 ;
        RECT 391.950 54.600 394.050 55.050 ;
        RECT 383.400 53.400 394.050 54.600 ;
        RECT 367.950 52.950 370.050 53.400 ;
        RECT 373.950 52.950 376.050 53.400 ;
        RECT 391.950 52.950 394.050 53.400 ;
        RECT 424.950 52.950 427.050 55.050 ;
        RECT 439.950 52.950 442.050 55.050 ;
        RECT 445.950 54.600 448.050 55.050 ;
        RECT 454.950 54.600 457.050 55.050 ;
        RECT 445.950 53.400 457.050 54.600 ;
        RECT 445.950 52.950 448.050 53.400 ;
        RECT 454.950 52.950 457.050 53.400 ;
        RECT 466.950 54.600 469.050 55.050 ;
        RECT 472.950 54.600 475.050 55.050 ;
        RECT 466.950 53.400 475.050 54.600 ;
        RECT 466.950 52.950 469.050 53.400 ;
        RECT 472.950 52.950 475.050 53.400 ;
        RECT 505.950 54.600 508.050 55.050 ;
        RECT 514.950 54.600 517.050 55.050 ;
        RECT 505.950 53.400 517.050 54.600 ;
        RECT 505.950 52.950 508.050 53.400 ;
        RECT 514.950 52.950 517.050 53.400 ;
        RECT 526.950 54.600 529.050 55.050 ;
        RECT 532.950 54.600 535.050 55.050 ;
        RECT 526.950 53.400 535.050 54.600 ;
        RECT 526.950 52.950 529.050 53.400 ;
        RECT 532.950 52.950 535.050 53.400 ;
        RECT 538.950 52.950 541.050 55.050 ;
        RECT 544.950 52.950 547.050 55.050 ;
        RECT 556.950 54.600 559.050 55.050 ;
        RECT 562.950 54.600 565.050 55.050 ;
        RECT 556.950 53.400 565.050 54.600 ;
        RECT 556.950 52.950 559.050 53.400 ;
        RECT 562.950 52.950 565.050 53.400 ;
        RECT 109.950 51.600 112.050 52.050 ;
        RECT 104.400 50.400 112.050 51.600 ;
        RECT 109.950 49.950 112.050 50.400 ;
        RECT 115.950 49.950 118.050 52.050 ;
        RECT 136.950 51.600 139.050 52.050 ;
        RECT 166.950 51.600 169.050 52.050 ;
        RECT 136.950 50.400 169.050 51.600 ;
        RECT 136.950 49.950 139.050 50.400 ;
        RECT 166.950 49.950 169.050 50.400 ;
        RECT 277.950 51.600 280.050 52.050 ;
        RECT 298.950 51.600 301.050 52.050 ;
        RECT 277.950 50.400 301.050 51.600 ;
        RECT 277.950 49.950 280.050 50.400 ;
        RECT 298.950 49.950 301.050 50.400 ;
        RECT 28.950 48.600 31.050 49.050 ;
        RECT 40.950 48.600 43.050 49.050 ;
        RECT 64.950 48.600 67.050 49.050 ;
        RECT 82.950 48.600 85.050 49.050 ;
        RECT 28.950 47.400 85.050 48.600 ;
        RECT 28.950 46.950 31.050 47.400 ;
        RECT 40.950 46.950 43.050 47.400 ;
        RECT 64.950 46.950 67.050 47.400 ;
        RECT 82.950 46.950 85.050 47.400 ;
        RECT 100.950 46.950 103.050 49.050 ;
        RECT 103.950 48.600 106.050 49.050 ;
        RECT 112.950 48.600 115.050 49.050 ;
        RECT 103.950 47.400 115.050 48.600 ;
        RECT 103.950 46.950 106.050 47.400 ;
        RECT 112.950 46.950 115.050 47.400 ;
        RECT 142.950 48.600 145.050 49.050 ;
        RECT 148.950 48.600 151.050 49.050 ;
        RECT 142.950 47.400 151.050 48.600 ;
        RECT 142.950 46.950 145.050 47.400 ;
        RECT 148.950 46.950 151.050 47.400 ;
        RECT 217.950 48.600 220.050 49.050 ;
        RECT 304.950 48.600 307.050 49.050 ;
        RECT 217.950 47.400 307.050 48.600 ;
        RECT 308.400 48.600 309.600 52.950 ;
        RECT 320.400 49.050 321.600 52.950 ;
        RECT 323.400 49.050 324.600 52.950 ;
        RECT 328.950 51.600 331.050 52.050 ;
        RECT 349.950 51.600 352.050 52.050 ;
        RECT 373.950 51.600 376.050 52.050 ;
        RECT 406.950 51.600 409.050 52.050 ;
        RECT 328.950 50.400 376.050 51.600 ;
        RECT 328.950 49.950 331.050 50.400 ;
        RECT 349.950 49.950 352.050 50.400 ;
        RECT 373.950 49.950 376.050 50.400 ;
        RECT 392.400 50.400 409.050 51.600 ;
        RECT 392.400 49.050 393.600 50.400 ;
        RECT 406.950 49.950 409.050 50.400 ;
        RECT 425.400 49.050 426.600 52.950 ;
        RECT 430.950 51.600 433.050 52.050 ;
        RECT 440.400 51.600 441.600 52.950 ;
        RECT 430.950 50.400 441.600 51.600 ;
        RECT 448.950 51.600 451.050 52.050 ;
        RECT 463.950 51.600 466.050 52.050 ;
        RECT 490.950 51.600 493.050 52.050 ;
        RECT 448.950 50.400 493.050 51.600 ;
        RECT 430.950 49.950 433.050 50.400 ;
        RECT 448.950 49.950 451.050 50.400 ;
        RECT 463.950 49.950 466.050 50.400 ;
        RECT 490.950 49.950 493.050 50.400 ;
        RECT 496.950 51.600 499.050 52.050 ;
        RECT 520.950 51.600 523.050 52.050 ;
        RECT 496.950 50.400 523.050 51.600 ;
        RECT 496.950 49.950 499.050 50.400 ;
        RECT 520.950 49.950 523.050 50.400 ;
        RECT 313.950 48.600 316.050 49.050 ;
        RECT 308.400 47.400 316.050 48.600 ;
        RECT 217.950 46.950 220.050 47.400 ;
        RECT 304.950 46.950 307.050 47.400 ;
        RECT 313.950 46.950 316.050 47.400 ;
        RECT 319.950 46.950 322.050 49.050 ;
        RECT 322.950 46.950 325.050 49.050 ;
        RECT 379.950 48.600 382.050 49.050 ;
        RECT 385.950 48.600 388.050 49.050 ;
        RECT 379.950 47.400 388.050 48.600 ;
        RECT 379.950 46.950 382.050 47.400 ;
        RECT 385.950 46.950 388.050 47.400 ;
        RECT 391.950 46.950 394.050 49.050 ;
        RECT 424.950 46.950 427.050 49.050 ;
        RECT 436.950 48.600 439.050 49.050 ;
        RECT 475.950 48.600 478.050 49.050 ;
        RECT 436.950 47.400 478.050 48.600 ;
        RECT 436.950 46.950 439.050 47.400 ;
        RECT 475.950 46.950 478.050 47.400 ;
        RECT 487.950 48.600 490.050 49.050 ;
        RECT 502.950 48.600 505.050 49.050 ;
        RECT 517.950 48.600 520.050 49.050 ;
        RECT 487.950 47.400 520.050 48.600 ;
        RECT 539.400 48.600 540.600 52.950 ;
        RECT 566.400 52.050 567.600 56.400 ;
        RECT 577.950 55.950 580.050 58.050 ;
        RECT 625.950 57.600 628.050 58.050 ;
        RECT 658.950 57.600 661.050 58.050 ;
        RECT 625.950 56.400 661.050 57.600 ;
        RECT 625.950 55.950 628.050 56.400 ;
        RECT 658.950 55.950 661.050 56.400 ;
        RECT 673.950 57.600 676.050 58.050 ;
        RECT 697.950 57.600 700.050 58.050 ;
        RECT 703.950 57.600 706.050 58.050 ;
        RECT 673.950 56.400 706.050 57.600 ;
        RECT 673.950 55.950 676.050 56.400 ;
        RECT 697.950 55.950 700.050 56.400 ;
        RECT 703.950 55.950 706.050 56.400 ;
        RECT 578.400 54.600 579.600 55.950 ;
        RECT 707.400 55.050 708.600 58.950 ;
        RECT 721.950 57.600 724.050 58.050 ;
        RECT 725.400 57.600 726.600 58.950 ;
        RECT 721.950 56.400 726.600 57.600 ;
        RECT 721.950 55.950 724.050 56.400 ;
        RECT 740.400 55.050 741.600 59.400 ;
        RECT 745.950 58.950 748.050 59.400 ;
        RECT 742.950 57.600 745.050 58.050 ;
        RECT 760.950 57.600 763.050 58.050 ;
        RECT 742.950 56.400 763.050 57.600 ;
        RECT 742.950 55.950 745.050 56.400 ;
        RECT 760.950 55.950 763.050 56.400 ;
        RECT 625.950 54.600 628.050 55.050 ;
        RECT 572.400 53.400 579.600 54.600 ;
        RECT 614.400 53.400 628.050 54.600 ;
        RECT 572.400 52.050 573.600 53.400 ;
        RECT 541.950 51.600 544.050 52.050 ;
        RECT 547.950 51.600 550.050 52.050 ;
        RECT 541.950 50.400 550.050 51.600 ;
        RECT 541.950 49.950 544.050 50.400 ;
        RECT 547.950 49.950 550.050 50.400 ;
        RECT 565.950 49.950 568.050 52.050 ;
        RECT 571.950 49.950 574.050 52.050 ;
        RECT 574.950 51.600 577.050 52.050 ;
        RECT 607.950 51.600 610.050 52.050 ;
        RECT 614.400 51.600 615.600 53.400 ;
        RECT 625.950 52.950 628.050 53.400 ;
        RECT 649.950 54.600 652.050 55.050 ;
        RECT 664.950 54.600 667.050 55.050 ;
        RECT 649.950 53.400 667.050 54.600 ;
        RECT 649.950 52.950 652.050 53.400 ;
        RECT 664.950 52.950 667.050 53.400 ;
        RECT 676.950 52.950 679.050 55.050 ;
        RECT 682.950 54.600 685.050 55.050 ;
        RECT 694.950 54.600 697.050 55.050 ;
        RECT 700.950 54.600 703.050 55.050 ;
        RECT 682.950 53.400 693.600 54.600 ;
        RECT 682.950 52.950 685.050 53.400 ;
        RECT 574.950 50.400 615.600 51.600 ;
        RECT 616.950 51.600 619.050 52.050 ;
        RECT 628.950 51.600 631.050 52.050 ;
        RECT 655.950 51.600 658.050 52.050 ;
        RECT 616.950 50.400 658.050 51.600 ;
        RECT 677.400 51.600 678.600 52.950 ;
        RECT 688.950 51.600 691.050 52.050 ;
        RECT 677.400 50.400 691.050 51.600 ;
        RECT 692.400 51.600 693.600 53.400 ;
        RECT 694.950 53.400 703.050 54.600 ;
        RECT 694.950 52.950 697.050 53.400 ;
        RECT 700.950 52.950 703.050 53.400 ;
        RECT 706.950 52.950 709.050 55.050 ;
        RECT 724.950 54.600 727.050 55.050 ;
        RECT 739.950 54.600 742.050 55.050 ;
        RECT 724.950 53.400 742.050 54.600 ;
        RECT 724.950 52.950 727.050 53.400 ;
        RECT 739.950 52.950 742.050 53.400 ;
        RECT 751.950 52.950 754.050 55.050 ;
        RECT 754.950 54.600 757.050 55.050 ;
        RECT 763.950 54.600 766.050 55.050 ;
        RECT 754.950 53.400 766.050 54.600 ;
        RECT 754.950 52.950 757.050 53.400 ;
        RECT 763.950 52.950 766.050 53.400 ;
        RECT 712.950 51.600 715.050 52.050 ;
        RECT 727.950 51.600 730.050 52.050 ;
        RECT 736.950 51.600 739.050 52.050 ;
        RECT 692.400 50.400 739.050 51.600 ;
        RECT 752.400 51.600 753.600 52.950 ;
        RECT 757.950 51.600 760.050 52.050 ;
        RECT 752.400 50.400 760.050 51.600 ;
        RECT 574.950 49.950 577.050 50.400 ;
        RECT 607.950 49.950 610.050 50.400 ;
        RECT 616.950 49.950 619.050 50.400 ;
        RECT 628.950 49.950 631.050 50.400 ;
        RECT 655.950 49.950 658.050 50.400 ;
        RECT 688.950 49.950 691.050 50.400 ;
        RECT 712.950 49.950 715.050 50.400 ;
        RECT 727.950 49.950 730.050 50.400 ;
        RECT 736.950 49.950 739.050 50.400 ;
        RECT 757.950 49.950 760.050 50.400 ;
        RECT 550.950 48.600 553.050 49.050 ;
        RECT 539.400 47.400 553.050 48.600 ;
        RECT 487.950 46.950 490.050 47.400 ;
        RECT 502.950 46.950 505.050 47.400 ;
        RECT 517.950 46.950 520.050 47.400 ;
        RECT 550.950 46.950 553.050 47.400 ;
        RECT 562.950 48.600 565.050 49.050 ;
        RECT 580.950 48.600 583.050 49.050 ;
        RECT 562.950 47.400 583.050 48.600 ;
        RECT 562.950 46.950 565.050 47.400 ;
        RECT 580.950 46.950 583.050 47.400 ;
        RECT 595.950 48.600 598.050 49.050 ;
        RECT 613.950 48.600 616.050 49.050 ;
        RECT 595.950 47.400 616.050 48.600 ;
        RECT 595.950 46.950 598.050 47.400 ;
        RECT 613.950 46.950 616.050 47.400 ;
        RECT 649.950 48.600 652.050 49.050 ;
        RECT 679.950 48.600 682.050 49.050 ;
        RECT 649.950 47.400 682.050 48.600 ;
        RECT 649.950 46.950 652.050 47.400 ;
        RECT 679.950 46.950 682.050 47.400 ;
        RECT 694.950 48.600 697.050 49.050 ;
        RECT 700.950 48.600 703.050 49.050 ;
        RECT 694.950 47.400 703.050 48.600 ;
        RECT 694.950 46.950 697.050 47.400 ;
        RECT 700.950 46.950 703.050 47.400 ;
        RECT 751.950 48.600 754.050 49.050 ;
        RECT 760.950 48.600 763.050 49.050 ;
        RECT 751.950 47.400 763.050 48.600 ;
        RECT 751.950 46.950 754.050 47.400 ;
        RECT 760.950 46.950 763.050 47.400 ;
        RECT 49.950 45.600 52.050 46.050 ;
        RECT 70.950 45.600 73.050 46.050 ;
        RECT 49.950 44.400 73.050 45.600 ;
        RECT 49.950 43.950 52.050 44.400 ;
        RECT 70.950 43.950 73.050 44.400 ;
        RECT 97.950 45.600 100.050 46.050 ;
        RECT 130.950 45.600 133.050 46.050 ;
        RECT 97.950 44.400 133.050 45.600 ;
        RECT 97.950 43.950 100.050 44.400 ;
        RECT 130.950 43.950 133.050 44.400 ;
        RECT 304.950 45.600 307.050 46.050 ;
        RECT 340.950 45.600 343.050 46.050 ;
        RECT 352.950 45.600 355.050 46.050 ;
        RECT 304.950 44.400 355.050 45.600 ;
        RECT 304.950 43.950 307.050 44.400 ;
        RECT 340.950 43.950 343.050 44.400 ;
        RECT 352.950 43.950 355.050 44.400 ;
        RECT 376.950 45.600 379.050 46.050 ;
        RECT 394.950 45.600 397.050 46.050 ;
        RECT 376.950 44.400 397.050 45.600 ;
        RECT 376.950 43.950 379.050 44.400 ;
        RECT 394.950 43.950 397.050 44.400 ;
        RECT 412.950 45.600 415.050 46.050 ;
        RECT 472.950 45.600 475.050 46.050 ;
        RECT 412.950 44.400 475.050 45.600 ;
        RECT 412.950 43.950 415.050 44.400 ;
        RECT 472.950 43.950 475.050 44.400 ;
        RECT 475.950 45.600 478.050 46.050 ;
        RECT 514.950 45.600 517.050 46.050 ;
        RECT 475.950 44.400 517.050 45.600 ;
        RECT 475.950 43.950 478.050 44.400 ;
        RECT 514.950 43.950 517.050 44.400 ;
        RECT 529.950 45.600 532.050 46.050 ;
        RECT 559.950 45.600 562.050 46.050 ;
        RECT 529.950 44.400 562.050 45.600 ;
        RECT 529.950 43.950 532.050 44.400 ;
        RECT 559.950 43.950 562.050 44.400 ;
        RECT 571.950 45.600 574.050 46.050 ;
        RECT 580.950 45.600 583.050 46.050 ;
        RECT 592.950 45.600 595.050 46.050 ;
        RECT 571.950 44.400 595.050 45.600 ;
        RECT 571.950 43.950 574.050 44.400 ;
        RECT 580.950 43.950 583.050 44.400 ;
        RECT 592.950 43.950 595.050 44.400 ;
        RECT 598.950 45.600 601.050 46.050 ;
        RECT 601.950 45.600 604.050 46.050 ;
        RECT 619.950 45.600 622.050 46.050 ;
        RECT 646.950 45.600 649.050 46.050 ;
        RECT 598.950 44.400 649.050 45.600 ;
        RECT 598.950 43.950 601.050 44.400 ;
        RECT 601.950 43.950 604.050 44.400 ;
        RECT 619.950 43.950 622.050 44.400 ;
        RECT 646.950 43.950 649.050 44.400 ;
        RECT 679.950 45.600 682.050 46.050 ;
        RECT 730.950 45.600 733.050 46.050 ;
        RECT 748.950 45.600 751.050 46.050 ;
        RECT 679.950 44.400 751.050 45.600 ;
        RECT 679.950 43.950 682.050 44.400 ;
        RECT 730.950 43.950 733.050 44.400 ;
        RECT 748.950 43.950 751.050 44.400 ;
        RECT 67.950 42.600 70.050 43.050 ;
        RECT 124.950 42.600 127.050 43.050 ;
        RECT 67.950 41.400 127.050 42.600 ;
        RECT 67.950 40.950 70.050 41.400 ;
        RECT 124.950 40.950 127.050 41.400 ;
        RECT 139.950 42.600 142.050 43.050 ;
        RECT 172.950 42.600 175.050 43.050 ;
        RECT 184.950 42.600 187.050 43.050 ;
        RECT 139.950 41.400 187.050 42.600 ;
        RECT 139.950 40.950 142.050 41.400 ;
        RECT 172.950 40.950 175.050 41.400 ;
        RECT 184.950 40.950 187.050 41.400 ;
        RECT 232.950 42.600 235.050 43.050 ;
        RECT 253.950 42.600 256.050 43.050 ;
        RECT 277.950 42.600 280.050 43.050 ;
        RECT 232.950 41.400 280.050 42.600 ;
        RECT 232.950 40.950 235.050 41.400 ;
        RECT 253.950 40.950 256.050 41.400 ;
        RECT 277.950 40.950 280.050 41.400 ;
        RECT 286.950 42.600 289.050 43.050 ;
        RECT 322.950 42.600 325.050 43.050 ;
        RECT 286.950 41.400 325.050 42.600 ;
        RECT 286.950 40.950 289.050 41.400 ;
        RECT 322.950 40.950 325.050 41.400 ;
        RECT 343.950 42.600 346.050 43.050 ;
        RECT 370.950 42.600 373.050 43.050 ;
        RECT 343.950 41.400 373.050 42.600 ;
        RECT 343.950 40.950 346.050 41.400 ;
        RECT 370.950 40.950 373.050 41.400 ;
        RECT 439.950 42.600 442.050 43.050 ;
        RECT 457.950 42.600 460.050 43.050 ;
        RECT 439.950 41.400 460.050 42.600 ;
        RECT 439.950 40.950 442.050 41.400 ;
        RECT 457.950 40.950 460.050 41.400 ;
        RECT 463.950 42.600 466.050 43.050 ;
        RECT 529.950 42.600 532.050 43.050 ;
        RECT 463.950 41.400 532.050 42.600 ;
        RECT 463.950 40.950 466.050 41.400 ;
        RECT 529.950 40.950 532.050 41.400 ;
        RECT 550.950 42.600 553.050 43.050 ;
        RECT 673.950 42.600 676.050 43.050 ;
        RECT 550.950 41.400 676.050 42.600 ;
        RECT 550.950 40.950 553.050 41.400 ;
        RECT 673.950 40.950 676.050 41.400 ;
        RECT 715.950 42.600 718.050 43.050 ;
        RECT 730.950 42.600 733.050 43.050 ;
        RECT 715.950 41.400 733.050 42.600 ;
        RECT 715.950 40.950 718.050 41.400 ;
        RECT 730.950 40.950 733.050 41.400 ;
        RECT 10.950 39.600 13.050 40.050 ;
        RECT 16.950 39.600 19.050 40.050 ;
        RECT 58.950 39.600 61.050 40.050 ;
        RECT 10.950 38.400 61.050 39.600 ;
        RECT 10.950 37.950 13.050 38.400 ;
        RECT 16.950 37.950 19.050 38.400 ;
        RECT 58.950 37.950 61.050 38.400 ;
        RECT 220.950 39.600 223.050 40.050 ;
        RECT 250.950 39.600 253.050 40.050 ;
        RECT 220.950 38.400 253.050 39.600 ;
        RECT 220.950 37.950 223.050 38.400 ;
        RECT 250.950 37.950 253.050 38.400 ;
        RECT 340.950 39.600 343.050 40.050 ;
        RECT 376.950 39.600 379.050 40.050 ;
        RECT 340.950 38.400 379.050 39.600 ;
        RECT 340.950 37.950 343.050 38.400 ;
        RECT 376.950 37.950 379.050 38.400 ;
        RECT 391.950 39.600 394.050 40.050 ;
        RECT 412.950 39.600 415.050 40.050 ;
        RECT 391.950 38.400 415.050 39.600 ;
        RECT 391.950 37.950 394.050 38.400 ;
        RECT 412.950 37.950 415.050 38.400 ;
        RECT 433.950 39.600 436.050 40.050 ;
        RECT 478.950 39.600 481.050 40.050 ;
        RECT 484.950 39.600 487.050 40.050 ;
        RECT 433.950 38.400 487.050 39.600 ;
        RECT 433.950 37.950 436.050 38.400 ;
        RECT 478.950 37.950 481.050 38.400 ;
        RECT 484.950 37.950 487.050 38.400 ;
        RECT 508.950 39.600 511.050 40.050 ;
        RECT 526.950 39.600 529.050 40.050 ;
        RECT 556.950 39.600 559.050 40.050 ;
        RECT 508.950 38.400 559.050 39.600 ;
        RECT 508.950 37.950 511.050 38.400 ;
        RECT 526.950 37.950 529.050 38.400 ;
        RECT 556.950 37.950 559.050 38.400 ;
        RECT 592.950 39.600 595.050 40.050 ;
        RECT 604.950 39.600 607.050 40.050 ;
        RECT 592.950 38.400 607.050 39.600 ;
        RECT 592.950 37.950 595.050 38.400 ;
        RECT 604.950 37.950 607.050 38.400 ;
        RECT 610.950 39.600 613.050 40.050 ;
        RECT 631.950 39.600 634.050 40.050 ;
        RECT 610.950 38.400 634.050 39.600 ;
        RECT 610.950 37.950 613.050 38.400 ;
        RECT 631.950 37.950 634.050 38.400 ;
        RECT 58.950 36.600 61.050 37.050 ;
        RECT 73.950 36.600 76.050 37.050 ;
        RECT 79.950 36.600 82.050 37.050 ;
        RECT 58.950 35.400 82.050 36.600 ;
        RECT 58.950 34.950 61.050 35.400 ;
        RECT 73.950 34.950 76.050 35.400 ;
        RECT 79.950 34.950 82.050 35.400 ;
        RECT 157.950 36.600 160.050 37.050 ;
        RECT 202.950 36.600 205.050 37.050 ;
        RECT 157.950 35.400 205.050 36.600 ;
        RECT 157.950 34.950 160.050 35.400 ;
        RECT 202.950 34.950 205.050 35.400 ;
        RECT 238.950 36.600 241.050 37.050 ;
        RECT 274.950 36.600 277.050 37.050 ;
        RECT 238.950 35.400 277.050 36.600 ;
        RECT 238.950 34.950 241.050 35.400 ;
        RECT 274.950 34.950 277.050 35.400 ;
        RECT 325.950 36.600 328.050 37.050 ;
        RECT 358.950 36.600 361.050 37.050 ;
        RECT 325.950 35.400 361.050 36.600 ;
        RECT 325.950 34.950 328.050 35.400 ;
        RECT 358.950 34.950 361.050 35.400 ;
        RECT 370.950 36.600 373.050 37.050 ;
        RECT 388.950 36.600 391.050 37.050 ;
        RECT 535.950 36.600 538.050 37.050 ;
        RECT 370.950 35.400 538.050 36.600 ;
        RECT 370.950 34.950 373.050 35.400 ;
        RECT 388.950 34.950 391.050 35.400 ;
        RECT 535.950 34.950 538.050 35.400 ;
        RECT 568.950 36.600 571.050 37.050 ;
        RECT 715.950 36.600 718.050 37.050 ;
        RECT 568.950 35.400 718.050 36.600 ;
        RECT 568.950 34.950 571.050 35.400 ;
        RECT 715.950 34.950 718.050 35.400 ;
        RECT 79.950 33.600 82.050 34.050 ;
        RECT 151.950 33.600 154.050 34.050 ;
        RECT 169.950 33.600 172.050 34.050 ;
        RECT 79.950 32.400 172.050 33.600 ;
        RECT 79.950 31.950 82.050 32.400 ;
        RECT 151.950 31.950 154.050 32.400 ;
        RECT 169.950 31.950 172.050 32.400 ;
        RECT 241.950 33.600 244.050 34.050 ;
        RECT 256.950 33.600 259.050 34.050 ;
        RECT 262.950 33.600 265.050 34.050 ;
        RECT 241.950 32.400 265.050 33.600 ;
        RECT 241.950 31.950 244.050 32.400 ;
        RECT 256.950 31.950 259.050 32.400 ;
        RECT 262.950 31.950 265.050 32.400 ;
        RECT 271.950 33.600 274.050 34.050 ;
        RECT 355.950 33.600 358.050 34.050 ;
        RECT 271.950 32.400 358.050 33.600 ;
        RECT 271.950 31.950 274.050 32.400 ;
        RECT 355.950 31.950 358.050 32.400 ;
        RECT 412.950 33.600 415.050 34.050 ;
        RECT 448.950 33.600 451.050 34.050 ;
        RECT 412.950 32.400 451.050 33.600 ;
        RECT 412.950 31.950 415.050 32.400 ;
        RECT 448.950 31.950 451.050 32.400 ;
        RECT 487.950 33.600 490.050 34.050 ;
        RECT 511.950 33.600 514.050 34.050 ;
        RECT 529.950 33.600 532.050 34.050 ;
        RECT 547.950 33.600 550.050 34.050 ;
        RECT 487.950 32.400 550.050 33.600 ;
        RECT 487.950 31.950 490.050 32.400 ;
        RECT 511.950 31.950 514.050 32.400 ;
        RECT 529.950 31.950 532.050 32.400 ;
        RECT 547.950 31.950 550.050 32.400 ;
        RECT 148.950 30.600 151.050 31.050 ;
        RECT 196.950 30.600 199.050 31.050 ;
        RECT 148.950 29.400 199.050 30.600 ;
        RECT 148.950 28.950 151.050 29.400 ;
        RECT 196.950 28.950 199.050 29.400 ;
        RECT 229.950 30.600 232.050 31.050 ;
        RECT 286.950 30.600 289.050 31.050 ;
        RECT 229.950 29.400 289.050 30.600 ;
        RECT 229.950 28.950 232.050 29.400 ;
        RECT 286.950 28.950 289.050 29.400 ;
        RECT 298.950 30.600 301.050 31.050 ;
        RECT 367.950 30.600 370.050 31.050 ;
        RECT 442.950 30.600 445.050 31.050 ;
        RECT 298.950 29.400 445.050 30.600 ;
        RECT 298.950 28.950 301.050 29.400 ;
        RECT 367.950 28.950 370.050 29.400 ;
        RECT 442.950 28.950 445.050 29.400 ;
        RECT 508.950 30.600 511.050 31.050 ;
        RECT 526.950 30.600 529.050 31.050 ;
        RECT 580.950 30.600 583.050 31.050 ;
        RECT 508.950 29.400 583.050 30.600 ;
        RECT 508.950 28.950 511.050 29.400 ;
        RECT 526.950 28.950 529.050 29.400 ;
        RECT 580.950 28.950 583.050 29.400 ;
        RECT 661.950 30.600 664.050 31.050 ;
        RECT 685.950 30.600 688.050 31.050 ;
        RECT 661.950 29.400 688.050 30.600 ;
        RECT 661.950 28.950 664.050 29.400 ;
        RECT 685.950 28.950 688.050 29.400 ;
        RECT 709.950 30.600 712.050 31.050 ;
        RECT 727.950 30.600 730.050 31.050 ;
        RECT 733.950 30.600 736.050 31.050 ;
        RECT 709.950 29.400 736.050 30.600 ;
        RECT 709.950 28.950 712.050 29.400 ;
        RECT 727.950 28.950 730.050 29.400 ;
        RECT 733.950 28.950 736.050 29.400 ;
        RECT 7.950 27.600 10.050 28.050 ;
        RECT 25.950 27.600 28.050 28.050 ;
        RECT 31.950 27.600 34.050 28.050 ;
        RECT 7.950 26.400 34.050 27.600 ;
        RECT 7.950 25.950 10.050 26.400 ;
        RECT 25.950 25.950 28.050 26.400 ;
        RECT 31.950 25.950 34.050 26.400 ;
        RECT 49.950 27.600 52.050 28.050 ;
        RECT 97.950 27.600 100.050 28.050 ;
        RECT 100.950 27.600 103.050 28.050 ;
        RECT 49.950 26.400 103.050 27.600 ;
        RECT 49.950 25.950 52.050 26.400 ;
        RECT 97.950 25.950 100.050 26.400 ;
        RECT 100.950 25.950 103.050 26.400 ;
        RECT 115.950 27.600 118.050 28.050 ;
        RECT 121.950 27.600 124.050 28.050 ;
        RECT 184.950 27.600 187.050 28.050 ;
        RECT 115.950 26.400 187.050 27.600 ;
        RECT 115.950 25.950 118.050 26.400 ;
        RECT 121.950 25.950 124.050 26.400 ;
        RECT 184.950 25.950 187.050 26.400 ;
        RECT 190.950 27.600 193.050 28.050 ;
        RECT 235.950 27.600 238.050 28.050 ;
        RECT 190.950 26.400 238.050 27.600 ;
        RECT 190.950 25.950 193.050 26.400 ;
        RECT 235.950 25.950 238.050 26.400 ;
        RECT 238.950 25.950 241.050 28.050 ;
        RECT 250.950 27.600 253.050 28.050 ;
        RECT 265.950 27.600 268.050 28.050 ;
        RECT 250.950 26.400 268.050 27.600 ;
        RECT 250.950 25.950 253.050 26.400 ;
        RECT 265.950 25.950 268.050 26.400 ;
        RECT 292.950 27.600 295.050 28.050 ;
        RECT 319.950 27.600 322.050 28.050 ;
        RECT 331.950 27.600 334.050 28.050 ;
        RECT 292.950 26.400 334.050 27.600 ;
        RECT 292.950 25.950 295.050 26.400 ;
        RECT 319.950 25.950 322.050 26.400 ;
        RECT 331.950 25.950 334.050 26.400 ;
        RECT 334.950 27.600 337.050 28.050 ;
        RECT 346.950 27.600 349.050 28.050 ;
        RECT 373.950 27.600 376.050 28.050 ;
        RECT 403.950 27.600 406.050 28.050 ;
        RECT 334.950 26.400 360.600 27.600 ;
        RECT 334.950 25.950 337.050 26.400 ;
        RECT 346.950 25.950 349.050 26.400 ;
        RECT 4.950 24.600 7.050 25.050 ;
        RECT 13.950 24.600 16.050 25.050 ;
        RECT 4.950 23.400 16.050 24.600 ;
        RECT 4.950 22.950 7.050 23.400 ;
        RECT 13.950 22.950 16.050 23.400 ;
        RECT 22.950 24.600 25.050 25.050 ;
        RECT 37.950 24.600 40.050 25.050 ;
        RECT 55.950 24.600 58.050 25.050 ;
        RECT 22.950 23.400 36.600 24.600 ;
        RECT 22.950 22.950 25.050 23.400 ;
        RECT 35.400 22.050 36.600 23.400 ;
        RECT 37.950 23.400 58.050 24.600 ;
        RECT 37.950 22.950 40.050 23.400 ;
        RECT 55.950 22.950 58.050 23.400 ;
        RECT 85.950 24.600 88.050 25.050 ;
        RECT 91.950 24.600 94.050 25.050 ;
        RECT 85.950 23.400 94.050 24.600 ;
        RECT 85.950 22.950 88.050 23.400 ;
        RECT 91.950 22.950 94.050 23.400 ;
        RECT 127.950 24.600 130.050 25.050 ;
        RECT 160.950 24.600 163.050 25.050 ;
        RECT 223.950 24.600 226.050 25.050 ;
        RECT 127.950 23.400 226.050 24.600 ;
        RECT 127.950 22.950 130.050 23.400 ;
        RECT 160.950 22.950 163.050 23.400 ;
        RECT 223.950 22.950 226.050 23.400 ;
        RECT 239.400 22.050 240.600 25.950 ;
        RECT 247.950 24.600 250.050 25.050 ;
        RECT 253.950 24.600 256.050 25.050 ;
        RECT 283.950 24.600 286.050 25.050 ;
        RECT 295.950 24.600 298.050 25.050 ;
        RECT 328.950 24.600 331.050 25.050 ;
        RECT 247.950 23.400 270.600 24.600 ;
        RECT 247.950 22.950 250.050 23.400 ;
        RECT 253.950 22.950 256.050 23.400 ;
        RECT 34.950 19.950 37.050 22.050 ;
        RECT 82.950 21.600 85.050 22.050 ;
        RECT 94.950 21.600 97.050 22.050 ;
        RECT 103.950 21.600 106.050 22.050 ;
        RECT 82.950 20.400 106.050 21.600 ;
        RECT 82.950 19.950 85.050 20.400 ;
        RECT 94.950 19.950 97.050 20.400 ;
        RECT 103.950 19.950 106.050 20.400 ;
        RECT 112.950 21.600 115.050 22.050 ;
        RECT 127.950 21.600 130.050 22.050 ;
        RECT 112.950 20.400 130.050 21.600 ;
        RECT 112.950 19.950 115.050 20.400 ;
        RECT 127.950 19.950 130.050 20.400 ;
        RECT 139.950 19.950 142.050 22.050 ;
        RECT 154.950 21.600 157.050 22.050 ;
        RECT 163.950 21.600 166.050 22.050 ;
        RECT 172.950 21.600 175.050 22.050 ;
        RECT 154.950 20.400 175.050 21.600 ;
        RECT 154.950 19.950 157.050 20.400 ;
        RECT 163.950 19.950 166.050 20.400 ;
        RECT 172.950 19.950 175.050 20.400 ;
        RECT 178.950 21.600 181.050 22.050 ;
        RECT 190.950 21.600 193.050 22.050 ;
        RECT 178.950 20.400 193.050 21.600 ;
        RECT 178.950 19.950 181.050 20.400 ;
        RECT 190.950 19.950 193.050 20.400 ;
        RECT 205.950 19.950 208.050 22.050 ;
        RECT 226.950 21.600 229.050 22.050 ;
        RECT 232.950 21.600 235.050 22.050 ;
        RECT 226.950 20.400 235.050 21.600 ;
        RECT 226.950 19.950 229.050 20.400 ;
        RECT 232.950 19.950 235.050 20.400 ;
        RECT 238.950 19.950 241.050 22.050 ;
        RECT 244.950 21.600 247.050 22.050 ;
        RECT 248.400 21.600 249.600 22.950 ;
        RECT 269.400 22.050 270.600 23.400 ;
        RECT 283.950 23.400 331.050 24.600 ;
        RECT 283.950 22.950 286.050 23.400 ;
        RECT 295.950 22.950 298.050 23.400 ;
        RECT 328.950 22.950 331.050 23.400 ;
        RECT 355.950 22.950 358.050 25.050 ;
        RECT 359.400 24.600 360.600 26.400 ;
        RECT 373.950 26.400 406.050 27.600 ;
        RECT 373.950 25.950 376.050 26.400 ;
        RECT 403.950 25.950 406.050 26.400 ;
        RECT 409.950 27.600 412.050 28.050 ;
        RECT 430.950 27.600 433.050 28.050 ;
        RECT 451.950 27.600 454.050 28.050 ;
        RECT 469.950 27.600 472.050 28.050 ;
        RECT 481.950 27.600 484.050 28.050 ;
        RECT 409.950 26.400 454.050 27.600 ;
        RECT 409.950 25.950 412.050 26.400 ;
        RECT 430.950 25.950 433.050 26.400 ;
        RECT 451.950 25.950 454.050 26.400 ;
        RECT 455.400 26.400 484.050 27.600 ;
        RECT 424.950 24.600 427.050 25.050 ;
        RECT 359.400 23.400 427.050 24.600 ;
        RECT 424.950 22.950 427.050 23.400 ;
        RECT 448.950 24.600 451.050 25.050 ;
        RECT 455.400 24.600 456.600 26.400 ;
        RECT 469.950 25.950 472.050 26.400 ;
        RECT 481.950 25.950 484.050 26.400 ;
        RECT 496.950 27.600 499.050 28.050 ;
        RECT 517.950 27.600 520.050 28.050 ;
        RECT 523.950 27.600 526.050 28.050 ;
        RECT 496.950 26.400 526.050 27.600 ;
        RECT 496.950 25.950 499.050 26.400 ;
        RECT 517.950 25.950 520.050 26.400 ;
        RECT 523.950 25.950 526.050 26.400 ;
        RECT 538.950 27.600 541.050 28.050 ;
        RECT 559.950 27.600 562.050 28.050 ;
        RECT 538.950 26.400 562.050 27.600 ;
        RECT 538.950 25.950 541.050 26.400 ;
        RECT 559.950 25.950 562.050 26.400 ;
        RECT 616.950 27.600 619.050 28.050 ;
        RECT 631.950 27.600 634.050 28.050 ;
        RECT 637.950 27.600 640.050 28.050 ;
        RECT 616.950 26.400 640.050 27.600 ;
        RECT 616.950 25.950 619.050 26.400 ;
        RECT 631.950 25.950 634.050 26.400 ;
        RECT 637.950 25.950 640.050 26.400 ;
        RECT 670.950 25.950 673.050 28.050 ;
        RECT 688.950 27.600 691.050 28.050 ;
        RECT 688.950 26.400 744.600 27.600 ;
        RECT 688.950 25.950 691.050 26.400 ;
        RECT 490.950 24.600 493.050 25.050 ;
        RECT 502.950 24.600 505.050 25.050 ;
        RECT 448.950 23.400 456.600 24.600 ;
        RECT 467.400 23.400 493.050 24.600 ;
        RECT 448.950 22.950 451.050 23.400 ;
        RECT 244.950 20.400 249.600 21.600 ;
        RECT 244.950 19.950 247.050 20.400 ;
        RECT 268.950 19.950 271.050 22.050 ;
        RECT 274.950 21.600 277.050 22.050 ;
        RECT 280.950 21.600 283.050 22.050 ;
        RECT 274.950 20.400 283.050 21.600 ;
        RECT 274.950 19.950 277.050 20.400 ;
        RECT 280.950 19.950 283.050 20.400 ;
        RECT 292.950 19.950 295.050 22.050 ;
        RECT 298.950 21.600 301.050 22.050 ;
        RECT 316.950 21.600 319.050 22.050 ;
        RECT 298.950 20.400 319.050 21.600 ;
        RECT 298.950 19.950 301.050 20.400 ;
        RECT 316.950 19.950 319.050 20.400 ;
        RECT 322.950 21.600 325.050 22.050 ;
        RECT 328.950 21.600 331.050 22.050 ;
        RECT 322.950 20.400 331.050 21.600 ;
        RECT 356.400 21.600 357.600 22.950 ;
        RECT 467.400 22.050 468.600 23.400 ;
        RECT 490.950 22.950 493.050 23.400 ;
        RECT 494.400 23.400 505.050 24.600 ;
        RECT 494.400 22.050 495.600 23.400 ;
        RECT 502.950 22.950 505.050 23.400 ;
        RECT 511.950 24.600 514.050 25.050 ;
        RECT 520.950 24.600 523.050 25.050 ;
        RECT 586.950 24.600 589.050 25.050 ;
        RECT 616.950 24.600 619.050 25.050 ;
        RECT 511.950 23.400 589.050 24.600 ;
        RECT 511.950 22.950 514.050 23.400 ;
        RECT 520.950 22.950 523.050 23.400 ;
        RECT 586.950 22.950 589.050 23.400 ;
        RECT 599.400 23.400 619.050 24.600 ;
        RECT 361.950 21.600 364.050 22.050 ;
        RECT 356.400 20.400 364.050 21.600 ;
        RECT 322.950 19.950 325.050 20.400 ;
        RECT 328.950 19.950 331.050 20.400 ;
        RECT 361.950 19.950 364.050 20.400 ;
        RECT 391.950 21.600 394.050 22.050 ;
        RECT 427.950 21.600 430.050 22.050 ;
        RECT 391.950 20.400 430.050 21.600 ;
        RECT 391.950 19.950 394.050 20.400 ;
        RECT 427.950 19.950 430.050 20.400 ;
        RECT 451.950 21.600 454.050 22.050 ;
        RECT 460.950 21.600 463.050 22.050 ;
        RECT 451.950 20.400 463.050 21.600 ;
        RECT 451.950 19.950 454.050 20.400 ;
        RECT 460.950 19.950 463.050 20.400 ;
        RECT 466.950 19.950 469.050 22.050 ;
        RECT 493.950 19.950 496.050 22.050 ;
        RECT 517.950 21.600 520.050 22.050 ;
        RECT 532.950 21.600 535.050 22.050 ;
        RECT 517.950 20.400 535.050 21.600 ;
        RECT 517.950 19.950 520.050 20.400 ;
        RECT 532.950 19.950 535.050 20.400 ;
        RECT 550.950 21.600 553.050 22.050 ;
        RECT 556.950 21.600 559.050 22.050 ;
        RECT 550.950 20.400 559.050 21.600 ;
        RECT 550.950 19.950 553.050 20.400 ;
        RECT 556.950 19.950 559.050 20.400 ;
        RECT 562.950 21.600 565.050 22.050 ;
        RECT 574.950 21.600 577.050 22.050 ;
        RECT 599.400 21.600 600.600 23.400 ;
        RECT 616.950 22.950 619.050 23.400 ;
        RECT 625.950 24.600 628.050 25.050 ;
        RECT 643.950 24.600 646.050 25.050 ;
        RECT 671.400 24.600 672.600 25.950 ;
        RECT 682.950 24.600 685.050 25.050 ;
        RECT 625.950 23.400 685.050 24.600 ;
        RECT 625.950 22.950 628.050 23.400 ;
        RECT 643.950 22.950 646.050 23.400 ;
        RECT 682.950 22.950 685.050 23.400 ;
        RECT 700.950 24.600 703.050 25.050 ;
        RECT 709.950 24.600 712.050 25.050 ;
        RECT 718.950 24.600 721.050 25.050 ;
        RECT 736.950 24.600 739.050 25.050 ;
        RECT 739.950 24.600 742.050 25.050 ;
        RECT 700.950 23.400 712.050 24.600 ;
        RECT 700.950 22.950 703.050 23.400 ;
        RECT 709.950 22.950 712.050 23.400 ;
        RECT 713.400 23.400 742.050 24.600 ;
        RECT 713.400 22.050 714.600 23.400 ;
        RECT 718.950 22.950 721.050 23.400 ;
        RECT 736.950 22.950 739.050 23.400 ;
        RECT 739.950 22.950 742.050 23.400 ;
        RECT 743.400 22.050 744.600 26.400 ;
        RECT 562.950 20.400 577.050 21.600 ;
        RECT 562.950 19.950 565.050 20.400 ;
        RECT 574.950 19.950 577.050 20.400 ;
        RECT 596.400 20.400 600.600 21.600 ;
        RECT 604.950 21.600 607.050 22.050 ;
        RECT 622.950 21.600 625.050 22.050 ;
        RECT 643.950 21.600 646.050 22.050 ;
        RECT 649.950 21.600 652.050 22.050 ;
        RECT 664.950 21.600 667.050 22.050 ;
        RECT 673.950 21.600 676.050 22.050 ;
        RECT 604.950 20.400 618.600 21.600 ;
        RECT 55.950 18.600 58.050 19.050 ;
        RECT 70.950 18.600 73.050 19.050 ;
        RECT 76.950 18.600 79.050 19.050 ;
        RECT 55.950 17.400 79.050 18.600 ;
        RECT 55.950 16.950 58.050 17.400 ;
        RECT 70.950 16.950 73.050 17.400 ;
        RECT 76.950 16.950 79.050 17.400 ;
        RECT 100.950 18.600 103.050 19.050 ;
        RECT 118.950 18.600 121.050 19.050 ;
        RECT 124.950 18.600 127.050 19.050 ;
        RECT 100.950 17.400 127.050 18.600 ;
        RECT 100.950 16.950 103.050 17.400 ;
        RECT 118.950 16.950 121.050 17.400 ;
        RECT 124.950 16.950 127.050 17.400 ;
        RECT 130.950 18.600 133.050 19.050 ;
        RECT 140.400 18.600 141.600 19.950 ;
        RECT 130.950 17.400 141.600 18.600 ;
        RECT 130.950 16.950 133.050 17.400 ;
        RECT 187.950 16.950 190.050 19.050 ;
        RECT 193.950 18.600 196.050 19.050 ;
        RECT 206.400 18.600 207.600 19.950 ;
        RECT 193.950 17.400 207.600 18.600 ;
        RECT 250.950 18.600 253.050 19.050 ;
        RECT 262.950 18.600 265.050 19.050 ;
        RECT 250.950 17.400 265.050 18.600 ;
        RECT 193.950 16.950 196.050 17.400 ;
        RECT 250.950 16.950 253.050 17.400 ;
        RECT 262.950 16.950 265.050 17.400 ;
        RECT 268.950 18.600 271.050 19.050 ;
        RECT 293.400 18.600 294.600 19.950 ;
        RECT 596.400 19.050 597.600 20.400 ;
        RECT 604.950 19.950 607.050 20.400 ;
        RECT 268.950 17.400 294.600 18.600 ;
        RECT 325.950 18.600 328.050 19.050 ;
        RECT 352.950 18.600 355.050 19.050 ;
        RECT 325.950 17.400 355.050 18.600 ;
        RECT 268.950 16.950 271.050 17.400 ;
        RECT 325.950 16.950 328.050 17.400 ;
        RECT 352.950 16.950 355.050 17.400 ;
        RECT 382.950 18.600 385.050 19.050 ;
        RECT 406.950 18.600 409.050 19.050 ;
        RECT 382.950 17.400 409.050 18.600 ;
        RECT 382.950 16.950 385.050 17.400 ;
        RECT 406.950 16.950 409.050 17.400 ;
        RECT 442.950 18.600 445.050 19.050 ;
        RECT 466.950 18.600 469.050 19.050 ;
        RECT 472.950 18.600 475.050 19.050 ;
        RECT 442.950 17.400 475.050 18.600 ;
        RECT 442.950 16.950 445.050 17.400 ;
        RECT 466.950 16.950 469.050 17.400 ;
        RECT 472.950 16.950 475.050 17.400 ;
        RECT 478.950 18.600 481.050 19.050 ;
        RECT 481.950 18.600 484.050 19.050 ;
        RECT 565.950 18.600 568.050 19.050 ;
        RECT 478.950 17.400 568.050 18.600 ;
        RECT 478.950 16.950 481.050 17.400 ;
        RECT 481.950 16.950 484.050 17.400 ;
        RECT 565.950 16.950 568.050 17.400 ;
        RECT 595.950 16.950 598.050 19.050 ;
        RECT 118.950 15.600 121.050 16.050 ;
        RECT 188.400 15.600 189.600 16.950 ;
        RECT 118.950 14.400 189.600 15.600 ;
        RECT 589.950 15.600 592.050 16.050 ;
        RECT 613.950 15.600 616.050 16.050 ;
        RECT 589.950 14.400 616.050 15.600 ;
        RECT 617.400 15.600 618.600 20.400 ;
        RECT 622.950 20.400 633.600 21.600 ;
        RECT 622.950 19.950 625.050 20.400 ;
        RECT 619.950 18.600 622.050 19.050 ;
        RECT 628.950 18.600 631.050 19.050 ;
        RECT 619.950 17.400 631.050 18.600 ;
        RECT 632.400 18.600 633.600 20.400 ;
        RECT 643.950 20.400 652.050 21.600 ;
        RECT 643.950 19.950 646.050 20.400 ;
        RECT 649.950 19.950 652.050 20.400 ;
        RECT 653.400 20.400 676.050 21.600 ;
        RECT 653.400 18.600 654.600 20.400 ;
        RECT 664.950 19.950 667.050 20.400 ;
        RECT 673.950 19.950 676.050 20.400 ;
        RECT 712.950 19.950 715.050 22.050 ;
        RECT 718.950 21.600 721.050 22.050 ;
        RECT 724.950 21.600 727.050 22.050 ;
        RECT 718.950 20.400 727.050 21.600 ;
        RECT 718.950 19.950 721.050 20.400 ;
        RECT 724.950 19.950 727.050 20.400 ;
        RECT 733.950 21.600 736.050 22.050 ;
        RECT 742.950 21.600 745.050 22.050 ;
        RECT 733.950 20.400 745.050 21.600 ;
        RECT 733.950 19.950 736.050 20.400 ;
        RECT 742.950 19.950 745.050 20.400 ;
        RECT 632.400 17.400 654.600 18.600 ;
        RECT 661.950 18.600 664.050 19.050 ;
        RECT 685.950 18.600 688.050 19.050 ;
        RECT 661.950 17.400 688.050 18.600 ;
        RECT 619.950 16.950 622.050 17.400 ;
        RECT 628.950 16.950 631.050 17.400 ;
        RECT 661.950 16.950 664.050 17.400 ;
        RECT 685.950 16.950 688.050 17.400 ;
        RECT 691.950 18.600 694.050 19.050 ;
        RECT 703.950 18.600 706.050 19.050 ;
        RECT 691.950 17.400 706.050 18.600 ;
        RECT 691.950 16.950 694.050 17.400 ;
        RECT 703.950 16.950 706.050 17.400 ;
        RECT 662.400 15.600 663.600 16.950 ;
        RECT 617.400 14.400 663.600 15.600 ;
        RECT 118.950 13.950 121.050 14.400 ;
        RECT 589.950 13.950 592.050 14.400 ;
        RECT 613.950 13.950 616.050 14.400 ;
        RECT 106.950 12.600 109.050 13.050 ;
        RECT 145.950 12.600 148.050 13.050 ;
        RECT 106.950 11.400 148.050 12.600 ;
        RECT 106.950 10.950 109.050 11.400 ;
        RECT 145.950 10.950 148.050 11.400 ;
        RECT 613.950 12.600 616.050 13.050 ;
        RECT 697.950 12.600 700.050 13.050 ;
        RECT 613.950 11.400 700.050 12.600 ;
        RECT 613.950 10.950 616.050 11.400 ;
        RECT 697.950 10.950 700.050 11.400 ;
  END
END ALU_wrapper
END LIBRARY

