magic
tech scmos
magscale 1 3
timestamp 1723012252
<< checkpaint >>
rect -15 -15 425 425
<< nwell >>
rect 110 110 300 300
<< pdiffusion >>
rect 195 195 215 215
<< psubstratepdiff >>
rect 45 345 365 365
rect 45 65 65 345
rect 345 65 365 345
rect 45 45 365 65
<< nsubstratendiff >>
rect 130 260 280 280
rect 130 150 150 260
rect 260 150 280 260
rect 130 130 280 150
<< metal1 >>
rect 45 345 365 365
rect 45 65 65 345
rect 130 260 280 280
rect 130 150 150 260
rect 195 195 215 215
rect 260 150 280 260
rect 130 130 280 150
rect 345 65 365 345
rect 45 45 365 65
use ntap_CDNS_7230122529113  ntap_CDNS_7230122529113_0
timestamp 1723012252
transform 1 0 256 0 1 146
box 4 4 24 114
use ntap_CDNS_7230122529113  ntap_CDNS_7230122529113_1
timestamp 1723012252
transform 0 1 146 1 0 256
box 4 4 24 114
use ntap_CDNS_7230122529113  ntap_CDNS_7230122529113_2
timestamp 1723012252
transform 0 1 146 1 0 126
box 4 4 24 114
use ntap_CDNS_7230122529113  ntap_CDNS_7230122529113_3
timestamp 1723012252
transform 1 0 126 0 1 146
box 4 4 24 114
use ptap_CDNS_7230122529114  ptap_CDNS_7230122529114_0
timestamp 1723012252
transform 0 1 71 1 0 41
box 4 4 24 264
use ptap_CDNS_7230122529114  ptap_CDNS_7230122529114_1
timestamp 1723012252
transform 1 0 41 0 1 71
box 4 4 24 264
use ptap_CDNS_7230122529114  ptap_CDNS_7230122529114_2
timestamp 1723012252
transform 0 1 71 1 0 341
box 4 4 24 264
use ptap_CDNS_7230122529114  ptap_CDNS_7230122529114_3
timestamp 1723012252
transform 1 0 341 0 1 71
box 4 4 24 264
use ptap_CDNS_7230122529115  ptap_CDNS_7230122529115_0
timestamp 1723012252
transform 1 0 191 0 1 191
box 4 4 24 24
<< end >>
