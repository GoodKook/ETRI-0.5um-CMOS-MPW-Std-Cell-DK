magic
tech scmos
magscale 1 3
timestamp 1555596690
<< checkpaint >>
rect -50 -50 300 300
use ndiode_CDNS_7230122529120  ndiode_CDNS_7230122529120_0
timestamp 1555596690
transform 1 0 0 0 1 0
box 10 10 240 240
<< end >>
