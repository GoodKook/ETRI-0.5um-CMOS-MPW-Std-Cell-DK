magic
tech scmos
magscale 1 3
timestamp 1726995271
<< checkpaint >>
rect 682 462 1826 472
rect -8 442 1826 462
rect -8 322 2056 442
rect 102 302 2056 322
rect 102 242 1552 302
rect -88 92 1552 242
rect -88 2 2596 92
rect -58 -48 2596 2
rect -58 -58 293 -48
use ndiode  ndiode_0
timestamp 1555596690
transform 1 0 962 0 1 2
box 10 10 240 240
use NMOS4  NMOS4_0
timestamp 1555596690
transform 1 0 157 0 1 0
box 5 2 76 134
use p2res  p2res_0
timestamp 1555596690
transform 1 0 44 0 1 374
box 8 8 1032 28
use pdiode  pdiode_0
timestamp 1555596690
transform 1 0 1222 0 1 12
box 0 0 270 270
use pipcap_CDNS_723012252914  pipcap_CDNS_723012252914_0
timestamp 1555596690
transform 1 0 0 0 1 0
box 2 2 142 122
use PMOS4  PMOS4_0
timestamp 1555596690
transform 1 0 162 0 1 152
box 0 0 88 142
use pnp2  pnp2_0
timestamp 1555596690
transform 1 0 217 0 1 -33
box 45 45 365 365
use pnp5  pnp5_0
timestamp 1555596690
transform 1 0 557 0 1 -33
box 45 45 395 395
<< end >>
