magic
tech scmos
magscale 1 2
timestamp 1727494898
<< nwell >>
rect -6 154 106 272
<< ntransistor >>
rect 20 14 24 74
rect 30 14 34 74
rect 44 14 48 74
<< ptransistor >>
rect 20 206 24 246
rect 40 206 44 246
rect 60 206 64 246
<< ndiffusion >>
rect 18 14 20 74
rect 24 14 30 74
rect 34 14 44 74
rect 48 72 62 74
rect 48 14 50 72
<< pdiffusion >>
rect 18 206 20 246
rect 24 206 26 246
rect 38 206 40 246
rect 44 210 46 246
rect 58 210 60 246
rect 44 206 60 210
rect 64 206 66 246
<< ndcontact >>
rect 6 14 18 74
rect 50 14 62 72
<< pdcontact >>
rect 6 206 18 246
rect 26 206 38 246
rect 46 210 58 246
rect 66 206 78 246
<< psubstratepcontact >>
rect 0 -6 100 6
<< nsubstratencontact >>
rect 0 254 100 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 20 194 24 206
rect 40 194 44 206
rect 10 190 24 194
rect 30 190 44 194
rect 10 123 16 190
rect 30 129 34 190
rect 60 123 64 206
rect 10 82 16 111
rect 10 78 24 82
rect 20 74 24 78
rect 30 74 34 117
rect 56 111 64 123
rect 53 82 57 111
rect 44 78 57 82
rect 44 74 48 78
rect 20 10 24 14
rect 30 10 34 14
rect 44 10 48 14
<< polycontact >>
rect 4 111 16 123
rect 24 117 36 129
rect 44 111 56 123
<< metal1 >>
rect 0 266 100 268
rect 0 252 100 254
rect 6 246 18 252
rect 46 246 58 252
rect 28 204 38 206
rect 66 204 72 206
rect 28 198 72 204
rect 66 117 72 198
rect 66 78 72 103
rect 50 72 72 78
rect 62 70 72 72
rect 6 8 18 14
rect 0 6 100 8
rect 0 -8 100 -6
<< m2contact >>
rect 3 123 17 137
rect 43 123 57 137
rect 23 103 37 117
rect 63 103 77 117
<< metal2 >>
rect 3 143 17 157
rect 3 137 16 143
rect 43 137 57 157
rect 23 83 37 103
rect 63 83 77 103
<< m2p >>
rect 3 143 17 157
rect 43 143 57 157
rect 23 83 37 97
rect 63 83 77 97
<< labels >>
rlabel metal2 3 143 17 157 0 A
port 0 nsew signal input
rlabel metal2 23 83 37 97 0 B
port 1 nsew signal input
rlabel metal2 43 143 57 157 0 C
port 2 nsew signal input
rlabel metal2 63 83 77 97 0 Y
port 3 nsew signal output
rlabel metal1 0 266 100 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 0 254 100 266 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 0 252 100 254 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 0 6 100 8 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 0 -6 100 6 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 0 -8 100 -6 0 gnd
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
