magic
tech scmos
magscale 1 2
timestamp 1728171741
<< nwell >>
rect -12 174 492 252
<< ntransistor >>
rect 24 14 28 54
rect 36 14 40 54
rect 60 14 64 54
rect 72 14 76 54
rect 122 14 126 34
rect 142 14 146 34
rect 162 14 166 34
rect 212 14 216 34
rect 232 14 236 34
rect 276 14 280 34
rect 296 14 300 34
rect 350 14 354 54
rect 362 14 366 54
rect 384 14 388 54
rect 396 14 400 54
rect 444 14 448 34
<< ptransistor >>
rect 22 186 26 226
rect 42 186 46 226
rect 62 186 66 226
rect 82 186 86 226
rect 126 206 130 226
rect 146 206 150 226
rect 166 186 170 226
rect 212 186 216 226
rect 232 186 236 226
rect 276 206 280 226
rect 296 206 300 226
rect 340 186 344 226
rect 360 186 364 226
rect 380 186 384 226
rect 400 186 404 226
rect 444 186 448 226
<< ndiffusion >>
rect 20 14 24 54
rect 28 14 36 54
rect 40 14 44 54
rect 56 14 60 54
rect 64 14 72 54
rect 76 14 80 54
rect 120 14 122 34
rect 126 14 128 34
rect 140 14 142 34
rect 146 14 148 34
rect 160 14 162 34
rect 166 14 168 34
rect 210 14 212 34
rect 216 14 218 34
rect 230 14 232 34
rect 236 14 238 34
rect 274 14 276 34
rect 280 14 282 34
rect 294 14 296 34
rect 300 14 302 34
rect 346 14 350 54
rect 354 14 362 54
rect 366 14 368 54
rect 380 14 384 54
rect 388 14 396 54
rect 400 14 404 54
rect 442 14 444 34
rect 448 14 450 34
<< pdiffusion >>
rect 20 186 22 226
rect 26 186 28 226
rect 40 186 42 226
rect 46 186 48 226
rect 60 186 62 226
rect 66 186 68 226
rect 80 186 82 226
rect 86 203 88 226
rect 124 206 126 226
rect 130 206 132 226
rect 144 206 146 226
rect 150 206 152 226
rect 164 206 166 226
rect 86 186 100 203
rect 154 186 166 206
rect 170 186 172 226
rect 210 186 212 226
rect 216 186 218 226
rect 230 186 232 226
rect 236 186 238 226
rect 274 206 276 226
rect 280 206 282 226
rect 294 206 296 226
rect 300 206 302 226
rect 338 186 340 226
rect 344 186 346 226
rect 358 186 360 226
rect 364 186 366 226
rect 378 186 380 226
rect 384 186 386 226
rect 398 186 400 226
rect 404 186 406 226
rect 442 186 444 226
rect 448 186 450 226
<< ndcontact >>
rect 8 14 20 54
rect 44 14 56 54
rect 80 14 92 54
rect 108 14 120 34
rect 128 14 140 34
rect 148 14 160 34
rect 168 14 180 34
rect 198 14 210 34
rect 218 14 230 34
rect 238 14 250 34
rect 262 14 274 34
rect 282 14 294 34
rect 302 14 314 34
rect 334 14 346 54
rect 368 14 380 54
rect 404 14 416 54
rect 430 14 442 34
rect 450 14 462 34
<< pdcontact >>
rect 8 186 20 226
rect 28 186 40 226
rect 48 186 60 226
rect 68 186 80 226
rect 88 203 100 226
rect 112 206 124 226
rect 132 206 144 226
rect 152 206 164 226
rect 172 186 184 226
rect 198 186 210 226
rect 218 186 230 226
rect 238 186 250 226
rect 262 206 274 226
rect 282 206 294 226
rect 302 206 314 226
rect 326 186 338 226
rect 346 186 358 226
rect 366 186 378 226
rect 386 186 398 226
rect 406 186 418 226
rect 430 186 442 226
rect 450 186 462 226
<< psubstratepcontact >>
rect -6 -6 486 6
<< nsubstratencontact >>
rect -6 234 486 246
<< polysilicon >>
rect 22 226 26 230
rect 42 226 46 230
rect 62 226 66 230
rect 82 226 86 230
rect 126 226 130 230
rect 146 226 150 230
rect 166 226 170 230
rect 212 226 216 230
rect 232 226 236 230
rect 276 226 280 230
rect 296 226 300 230
rect 340 226 344 230
rect 360 226 364 230
rect 380 226 384 230
rect 400 226 404 230
rect 444 226 448 230
rect 22 123 26 186
rect 42 168 46 186
rect 22 111 24 123
rect 24 54 28 111
rect 44 72 48 156
rect 62 151 66 186
rect 36 54 40 60
rect 60 54 64 139
rect 82 116 86 186
rect 126 107 130 206
rect 82 84 86 104
rect 127 95 130 107
rect 146 117 150 206
rect 146 87 150 105
rect 166 87 170 186
rect 212 105 216 186
rect 232 128 236 186
rect 276 171 280 206
rect 256 159 280 171
rect 232 122 244 128
rect 212 93 219 105
rect 72 80 86 84
rect 122 83 150 87
rect 72 54 76 80
rect 122 34 126 83
rect 142 34 146 63
rect 162 34 166 75
rect 212 54 216 93
rect 240 72 244 122
rect 276 88 280 159
rect 296 117 300 206
rect 340 168 344 186
rect 300 105 314 117
rect 276 82 300 88
rect 236 66 244 72
rect 192 42 216 54
rect 212 34 216 42
rect 232 34 236 60
rect 276 34 280 60
rect 296 34 300 82
rect 308 72 314 105
rect 328 62 334 168
rect 360 166 364 186
rect 380 180 384 186
rect 350 160 364 166
rect 350 122 356 160
rect 380 150 384 168
rect 370 144 384 150
rect 344 70 350 110
rect 370 90 374 144
rect 400 143 404 186
rect 400 102 404 131
rect 372 78 374 90
rect 344 66 366 70
rect 328 58 354 62
rect 350 54 354 58
rect 362 54 366 66
rect 370 62 374 78
rect 380 98 404 102
rect 380 70 384 98
rect 444 90 448 186
rect 404 78 448 90
rect 380 66 400 70
rect 370 58 388 62
rect 384 54 388 58
rect 396 54 400 66
rect 444 34 448 78
rect 24 10 28 14
rect 36 10 40 14
rect 60 10 64 14
rect 72 10 76 14
rect 122 10 126 14
rect 142 10 146 14
rect 162 10 166 14
rect 212 10 216 14
rect 232 10 236 14
rect 276 10 280 14
rect 296 10 300 14
rect 350 10 354 14
rect 362 10 366 14
rect 384 10 388 14
rect 396 10 400 14
rect 444 10 448 14
<< polycontact >>
rect 38 156 50 168
rect 24 111 36 123
rect 36 60 48 72
rect 60 139 72 151
rect 77 104 89 116
rect 115 95 127 107
rect 146 105 158 117
rect 244 159 256 171
rect 219 93 231 105
rect 162 75 174 87
rect 137 63 149 75
rect 328 168 340 180
rect 288 105 300 117
rect 224 60 236 72
rect 180 42 192 54
rect 276 60 288 72
rect 308 60 320 72
rect 372 168 384 180
rect 344 110 356 122
rect 392 131 404 143
rect 360 78 372 90
rect 392 78 404 90
<< metal1 >>
rect -6 246 486 248
rect -6 232 486 234
rect 8 226 20 232
rect 48 226 60 232
rect 88 226 100 232
rect 172 226 184 232
rect 218 226 230 232
rect 326 226 338 232
rect 366 226 378 232
rect 406 226 418 232
rect 450 226 462 232
rect 109 206 112 226
rect 130 206 132 226
rect 151 206 152 226
rect 109 197 115 206
rect 130 197 137 206
rect 151 197 159 206
rect 28 180 35 186
rect 8 174 35 180
rect 8 84 16 174
rect 68 166 80 186
rect 157 183 159 197
rect 263 186 271 206
rect 283 186 294 206
rect 303 198 311 206
rect 203 180 210 186
rect 346 180 358 186
rect 297 172 328 177
rect 237 171 251 172
rect 50 158 187 166
rect 237 159 244 171
rect 283 169 328 172
rect 346 172 372 180
rect 174 152 187 158
rect 72 143 123 151
rect 174 145 263 152
rect 390 155 398 186
rect 317 149 416 155
rect 23 123 37 137
rect 174 131 392 139
rect 77 125 187 131
rect 77 117 89 125
rect 63 116 89 117
rect 27 97 35 111
rect 63 103 77 116
rect 95 113 140 119
rect 95 97 103 113
rect 27 90 103 97
rect 8 78 110 84
rect 8 54 16 78
rect 48 60 92 68
rect 82 54 92 60
rect 103 57 110 78
rect 120 72 127 95
rect 133 99 140 113
rect 158 111 203 113
rect 217 117 300 121
rect 217 113 288 117
rect 158 105 213 111
rect 133 93 213 99
rect 309 110 344 122
rect 309 99 315 110
rect 363 104 377 117
rect 206 87 213 93
rect 251 92 315 99
rect 322 97 377 104
rect 251 87 257 92
rect 174 75 197 85
rect 206 78 257 87
rect 322 85 329 97
rect 263 78 329 85
rect 352 78 360 88
rect 372 78 392 88
rect 120 64 137 72
rect 149 63 171 69
rect 183 63 197 75
rect 263 72 270 78
rect 165 54 171 63
rect 236 60 270 72
rect 288 60 308 72
rect 352 54 362 78
rect 410 54 416 149
rect 165 45 180 54
rect 108 34 117 43
rect 128 34 137 43
rect 148 34 157 43
rect 203 34 210 40
rect 239 34 250 40
rect 263 34 274 40
rect 283 34 294 40
rect 305 34 314 40
rect 346 46 362 54
rect 430 117 440 186
rect 430 103 457 117
rect 430 34 440 103
rect 44 8 56 14
rect 168 8 180 14
rect 218 8 230 14
rect 368 8 380 14
rect 450 8 462 14
rect -6 6 486 8
rect -6 -8 486 -6
<< m2contact >>
rect 103 183 117 197
rect 123 183 137 197
rect 143 183 157 197
rect 203 166 217 180
rect 237 172 251 186
rect 263 172 277 186
rect 283 172 297 186
rect 303 184 317 198
rect 123 137 137 151
rect 263 145 277 159
rect 303 145 317 159
rect 203 111 217 125
rect 231 93 245 107
rect 103 43 117 57
rect 123 43 137 57
rect 143 43 157 57
rect 203 40 217 54
rect 237 40 251 54
rect 263 40 277 54
rect 283 40 297 54
rect 303 40 317 54
<< metal2 >>
rect 107 57 115 183
rect 127 151 135 183
rect 127 57 135 137
rect 147 57 155 183
rect 205 125 213 166
rect 205 54 213 111
rect 241 107 249 172
rect 267 159 275 172
rect 245 93 249 107
rect 243 54 249 93
rect 265 54 275 145
rect 289 54 297 172
rect 305 159 313 184
rect 305 54 313 145
<< m1p >>
rect 23 123 37 137
rect 63 103 77 117
rect 363 103 377 117
rect 443 103 457 117
rect 183 63 197 77
<< labels >>
rlabel metal1 -6 -8 486 8 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal1 443 103 457 117 0 Q
port 4 nsew signal output
rlabel metal1 183 63 197 77 0 D
port 2 nsew signal input
rlabel metal1 63 103 77 117 0 S
port 1 nsew signal input
rlabel metal1 -6 232 486 248 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 363 103 377 117 0 CLK
port 3 nsew clock input
rlabel metal1 23 123 37 137 0 R
port 0 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 480 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
