magic
tech scmos
magscale 1 2
timestamp 1727851015
<< metal1 >>
rect -63 5762 30 5778
rect -63 5298 -3 5762
rect 37 5657 73 5663
rect 37 5567 43 5657
rect 833 5663 847 5673
rect 267 5657 303 5663
rect 833 5660 873 5663
rect 837 5657 873 5660
rect 297 5607 303 5657
rect 767 5633 773 5647
rect 407 5613 413 5627
rect 1237 5623 1243 5733
rect 4197 5717 4223 5723
rect 1447 5653 1453 5667
rect 1527 5653 1533 5667
rect 1307 5633 1313 5647
rect 1777 5643 1783 5673
rect 3157 5657 3193 5663
rect 1777 5637 1813 5643
rect 2047 5633 2053 5647
rect 1207 5617 1243 5623
rect 1637 5567 1643 5633
rect 2517 5627 2523 5653
rect 2567 5633 2573 5647
rect 2757 5623 2763 5653
rect 2757 5617 2793 5623
rect 2997 5587 3003 5653
rect 3107 5633 3113 5647
rect 3157 5607 3163 5657
rect 3327 5633 3333 5647
rect 3517 5567 3523 5653
rect 3737 5643 3743 5673
rect 4217 5667 4223 5717
rect 3707 5637 3743 5643
rect 4847 5643 4860 5647
rect 4847 5637 4873 5643
rect 4847 5633 4860 5637
rect 5160 5643 5173 5647
rect 5147 5637 5173 5643
rect 5160 5633 5173 5637
rect 5067 5613 5073 5627
rect 5723 5538 5783 5778
rect 5690 5522 5783 5538
rect 47 5443 60 5447
rect 47 5437 73 5443
rect 47 5433 60 5437
rect 317 5407 323 5433
rect 457 5427 463 5473
rect 597 5423 603 5493
rect 837 5443 843 5473
rect 4133 5467 4147 5473
rect 837 5437 873 5443
rect 597 5417 633 5423
rect 1007 5413 1013 5427
rect 2380 5423 2392 5427
rect 2367 5417 2392 5423
rect 2380 5413 2392 5417
rect 2607 5413 2613 5427
rect 3057 5423 3063 5453
rect 3837 5437 3873 5443
rect 3057 5417 3093 5423
rect 177 5397 213 5403
rect 177 5367 183 5397
rect 787 5397 823 5403
rect 817 5347 823 5397
rect 1607 5397 1643 5403
rect 1237 5347 1243 5373
rect 1637 5327 1643 5397
rect 1747 5397 1783 5403
rect 1777 5367 1783 5397
rect 1947 5393 1953 5407
rect 2160 5403 2172 5407
rect 2147 5397 2172 5403
rect 2160 5393 2172 5397
rect 2507 5397 2543 5403
rect 1873 5387 1887 5393
rect 2537 5367 2543 5397
rect 2687 5393 2693 5407
rect 2807 5403 2820 5407
rect 2807 5397 2833 5403
rect 2807 5393 2820 5397
rect 3177 5387 3183 5413
rect 3577 5407 3583 5433
rect 3057 5327 3063 5373
rect 3837 5327 3843 5437
rect 4867 5433 4873 5447
rect 3977 5387 3983 5433
rect 4127 5413 4133 5427
rect 4317 5417 4353 5423
rect 4267 5397 4303 5403
rect 4297 5347 4303 5397
rect 4317 5387 4323 5417
rect 4677 5367 4683 5413
rect 5077 5327 5083 5493
rect 5517 5387 5523 5453
rect -63 5282 30 5298
rect -63 4818 -3 5282
rect 157 5127 163 5253
rect 277 5207 283 5233
rect 277 5167 283 5193
rect 507 5173 513 5187
rect 697 5147 703 5173
rect 587 5133 593 5147
rect 977 5143 983 5193
rect 1407 5173 1413 5187
rect 1777 5183 1783 5253
rect 1777 5177 1813 5183
rect 2607 5173 2613 5187
rect 3147 5173 3153 5187
rect 3197 5183 3203 5253
rect 3197 5177 3233 5183
rect 2747 5153 2753 5167
rect 2917 5147 2923 5173
rect 977 5137 1013 5143
rect 1267 5133 1273 5147
rect 1667 5133 1673 5147
rect 3457 5087 3463 5213
rect 3617 5127 3623 5153
rect 3757 5143 3763 5193
rect 3927 5153 3933 5167
rect 3757 5137 3793 5143
rect 4257 5107 4263 5193
rect 4277 5143 4283 5233
rect 4417 5163 4423 5253
rect 4417 5157 4453 5163
rect 4277 5137 4313 5143
rect 4353 5127 4367 5133
rect 4497 5127 4503 5233
rect 5537 5127 5543 5213
rect 5640 5163 5653 5167
rect 5627 5157 5653 5163
rect 5640 5153 5653 5157
rect 5723 5058 5783 5522
rect 5690 5042 5783 5058
rect 1180 5023 1193 5027
rect 1177 5013 1193 5023
rect 157 4867 163 5013
rect 437 4867 443 4993
rect 467 4953 473 4967
rect 577 4867 583 5013
rect 1177 4987 1183 5013
rect 887 4933 893 4947
rect 1177 4927 1183 4973
rect 1357 4967 1363 4993
rect 1747 4933 1753 4947
rect 1937 4937 1973 4943
rect 607 4913 613 4927
rect 1827 4913 1833 4927
rect 1937 4907 1943 4937
rect 2537 4943 2543 5013
rect 2613 4987 2627 4993
rect 4017 4967 4023 5013
rect 5347 4953 5353 4967
rect 5437 4957 5473 4963
rect 2620 4943 2633 4947
rect 2507 4937 2543 4943
rect 2607 4937 2633 4943
rect 2620 4933 2633 4937
rect 3360 4943 3373 4947
rect 3347 4937 3373 4943
rect 3360 4933 3373 4937
rect 3767 4933 3773 4947
rect 697 4867 703 4893
rect 2877 4867 2883 4933
rect 4017 4867 4023 4953
rect 4227 4937 4263 4943
rect 4257 4887 4263 4937
rect 4617 4907 4623 4953
rect 4477 4867 4483 4893
rect 4957 4847 4963 4913
rect 5437 4847 5443 4957
rect -63 4802 30 4818
rect -63 4338 -3 4802
rect 37 4697 73 4703
rect 37 4647 43 4697
rect 397 4687 403 4733
rect 2613 4720 2627 4733
rect 687 4697 723 4703
rect 267 4653 273 4667
rect 717 4607 723 4697
rect 827 4697 863 4703
rect 857 4607 863 4697
rect 1367 4697 1403 4703
rect 997 4663 1003 4693
rect 967 4657 1003 4663
rect 1397 4607 1403 4697
rect 1567 4693 1573 4707
rect 1867 4693 1873 4707
rect 2147 4673 2153 4687
rect 2217 4683 2223 4713
rect 2617 4707 2623 4720
rect 2217 4677 2253 4683
rect 2657 4667 2663 4773
rect 2873 4707 2887 4713
rect 3287 4693 3292 4707
rect 3047 4673 3053 4687
rect 3147 4673 3153 4687
rect 3607 4673 3613 4687
rect 3777 4667 3783 4713
rect 2006 4653 2013 4667
rect 3487 4653 3493 4667
rect 5187 4653 5193 4667
rect 5247 4653 5253 4667
rect 3997 4607 4003 4653
rect 5723 4578 5783 5042
rect 5690 4562 5783 4578
rect 177 4483 183 4533
rect 2157 4487 2163 4533
rect 177 4477 213 4483
rect 1827 4473 1833 4487
rect 887 4453 893 4467
rect 557 4437 593 4443
rect 557 4367 563 4437
rect 787 4437 823 4443
rect 817 4407 823 4437
rect 1027 4437 1063 4443
rect 1057 4367 1063 4437
rect 1167 4433 1173 4447
rect 1337 4443 1343 4473
rect 1307 4437 1343 4443
rect 1457 4427 1463 4473
rect 1508 4453 1513 4467
rect 1947 4443 1960 4447
rect 1947 4437 1973 4443
rect 1947 4433 1960 4437
rect 2337 4387 2343 4533
rect 2457 4477 2493 4483
rect 2457 4447 2463 4477
rect 3087 4473 3093 4487
rect 3307 4473 3313 4487
rect 4087 4477 4113 4483
rect 5207 4473 5213 4487
rect 3237 4447 3243 4473
rect 4117 4447 4123 4473
rect 4397 4457 4433 4463
rect 2417 4420 2423 4433
rect 3157 4420 3163 4433
rect 2413 4407 2427 4420
rect 3153 4407 3167 4420
rect 4397 4407 4403 4457
rect -63 4322 30 4338
rect -63 3858 -3 4322
rect 207 4213 213 4227
rect 447 4223 460 4227
rect 447 4217 473 4223
rect 447 4213 460 4217
rect 577 4187 583 4293
rect 113 4167 127 4173
rect 126 4157 127 4167
rect 717 4127 723 4193
rect 1117 4183 1123 4293
rect 1167 4213 1173 4227
rect 1307 4193 1313 4207
rect 1377 4203 1383 4233
rect 1377 4197 1413 4203
rect 1087 4177 1123 4183
rect 1617 4147 1623 4253
rect 1647 4213 1653 4227
rect 2397 4207 2403 4273
rect 2137 4147 2143 4173
rect 2417 4167 2423 4233
rect 2697 4187 2703 4293
rect 2927 4197 2963 4203
rect 2447 4173 2453 4187
rect 2697 4147 2703 4173
rect 1617 4137 1633 4147
rect 1620 4133 1633 4137
rect 2957 4127 2963 4197
rect 3097 4183 3103 4273
rect 3097 4177 3133 4183
rect 3237 4167 3243 4273
rect 3547 4193 3553 4207
rect 4057 4147 4063 4273
rect 4177 4227 4183 4253
rect 4177 4183 4183 4213
rect 4573 4187 4587 4193
rect 4147 4177 4183 4183
rect 4726 4173 4733 4187
rect 5140 4183 5152 4187
rect 5127 4177 5152 4183
rect 5140 4173 5152 4177
rect 5723 4098 5783 4562
rect 5690 4082 5783 4098
rect 697 4007 703 4033
rect 267 3993 273 4007
rect 1307 3993 1313 4007
rect 1357 3997 1393 4003
rect 407 3953 413 3967
rect 697 3927 703 3993
rect 1077 3957 1113 3963
rect 1077 3907 1083 3957
rect 1357 3927 1363 3997
rect 1617 3967 1623 4033
rect 2077 4003 2083 4033
rect 2047 3997 2083 4003
rect 2257 4003 2263 4053
rect 2257 3997 2293 4003
rect 2447 3997 2483 4003
rect 1667 3973 1673 3987
rect 2477 3947 2483 3997
rect 2497 3967 2503 4033
rect 2527 3993 2533 4007
rect 3627 3993 3633 4007
rect 3687 3993 3693 4007
rect 3947 3993 3953 4007
rect 3347 3973 3353 3987
rect 4297 3983 4303 4053
rect 5077 4003 5083 4033
rect 5077 3997 5113 4003
rect 4267 3977 4303 3983
rect 3427 3953 3433 3967
rect 4017 3927 4023 3973
rect 4357 3940 4363 3953
rect 4353 3927 4367 3940
rect 5037 3940 5043 3953
rect 4717 3907 4723 3933
rect 5033 3927 5047 3940
rect 5217 3887 5223 4053
rect 5677 3987 5683 4053
rect 5467 3973 5473 3987
rect 5527 3977 5563 3983
rect 5557 3887 5563 3977
rect -63 3842 30 3858
rect -63 3378 -3 3842
rect 297 3707 303 3753
rect 797 3737 833 3743
rect 587 3713 593 3727
rect 67 3693 73 3707
rect 687 3693 693 3707
rect 533 3687 547 3692
rect 797 3647 803 3737
rect 1267 3733 1273 3747
rect 1407 3713 1413 3727
rect 1757 3717 1793 3723
rect 1097 3697 1133 3703
rect 1097 3667 1103 3697
rect 1757 3667 1763 3717
rect 1997 3667 2003 3813
rect 2086 3773 2087 3780
rect 2073 3760 2087 3773
rect 2077 3747 2083 3760
rect 2117 3687 2123 3773
rect 2257 3703 2263 3813
rect 2953 3760 2967 3773
rect 2957 3747 2963 3760
rect 2997 3747 3003 3793
rect 3627 3733 3633 3747
rect 3767 3737 3803 3743
rect 2547 3713 2553 3727
rect 2227 3697 2263 3703
rect 3137 3647 3143 3713
rect 3797 3707 3803 3737
rect 3907 3733 3913 3747
rect 5607 3713 5613 3727
rect 4593 3707 4607 3713
rect 5723 3618 5783 4082
rect 5690 3602 5783 3618
rect 267 3473 273 3487
rect 437 3483 443 3553
rect 547 3513 553 3527
rect 967 3517 1003 3523
rect 407 3477 443 3483
rect 827 3473 833 3487
rect 997 3447 1003 3517
rect 1566 3513 1573 3527
rect 1787 3513 1793 3527
rect 1047 3493 1053 3507
rect 2217 3497 2253 3503
rect 1593 3487 1607 3493
rect 1367 3473 1373 3487
rect 1537 3447 1543 3473
rect 2217 3427 2223 3497
rect 2297 3427 2303 3553
rect 2527 3513 2533 3527
rect 2627 3493 2633 3507
rect 2777 3447 2783 3513
rect 2987 3493 2993 3507
rect 3157 3483 3163 3533
rect 3267 3513 3273 3527
rect 3297 3507 3303 3573
rect 3507 3513 3513 3527
rect 3367 3500 3403 3503
rect 3367 3497 3407 3500
rect 3127 3477 3163 3483
rect 3393 3487 3407 3497
rect 3677 3483 3683 3573
rect 4587 3513 4593 3527
rect 5167 3517 5203 3523
rect 3867 3493 3873 3507
rect 4127 3493 4133 3507
rect 3647 3477 3683 3483
rect 4437 3447 4443 3513
rect 5197 3407 5203 3517
rect 5407 3493 5413 3507
rect 5297 3447 5303 3493
rect 5537 3480 5543 3493
rect 5533 3467 5547 3480
rect 5697 3407 5703 3493
rect -63 3362 30 3378
rect -63 2898 -3 3362
rect 2107 3343 2120 3347
rect 2107 3333 2123 3343
rect 407 3253 413 3267
rect 457 3263 463 3313
rect 457 3257 493 3263
rect 717 3223 723 3273
rect 1237 3263 1243 3313
rect 1207 3257 1243 3263
rect 1647 3253 1653 3267
rect 1913 3247 1927 3253
rect 767 3233 773 3247
rect 847 3233 853 3247
rect 1427 3233 1433 3247
rect 1787 3233 1793 3247
rect 687 3217 723 3223
rect 927 3213 933 3227
rect 1527 3213 1533 3227
rect 1587 3213 1594 3227
rect 1977 3223 1983 3253
rect 2117 3247 2123 3333
rect 2273 3267 2287 3273
rect 2286 3260 2287 3267
rect 2447 3253 2453 3267
rect 2637 3227 2643 3273
rect 1947 3217 1983 3223
rect 2587 3217 2623 3223
rect 1257 3167 1263 3193
rect 2617 3167 2623 3217
rect 2777 3187 2783 3333
rect 4657 3267 4663 3293
rect 2927 3233 2933 3247
rect 3213 3240 3227 3253
rect 3217 3237 3223 3240
rect 3287 3233 3293 3247
rect 3420 3243 3433 3247
rect 3407 3237 3433 3243
rect 3420 3233 3433 3237
rect 3713 3233 3714 3243
rect 3713 3227 3727 3233
rect 3953 3227 3967 3233
rect 4917 3227 4923 3273
rect 5077 3243 5083 3273
rect 5077 3237 5113 3243
rect 3087 3213 3093 3227
rect 3467 3213 3473 3227
rect 5560 3223 5573 3227
rect 5547 3217 5573 3223
rect 5560 3213 5573 3217
rect 5697 3223 5703 3333
rect 5667 3217 5703 3223
rect 3233 3207 3247 3212
rect 5723 3138 5783 3602
rect 5690 3122 5783 3138
rect 37 3037 73 3043
rect 37 2927 43 3037
rect 277 3007 283 3093
rect 297 2947 303 3053
rect 467 3033 473 3047
rect 1617 3037 1653 3043
rect 747 3013 753 3027
rect 327 2993 333 3007
rect 577 2997 613 3003
rect 577 2967 583 2997
rect 1197 2997 1233 3003
rect 1197 2967 1203 2997
rect 1437 2967 1443 3033
rect 1617 2967 1623 3037
rect 1737 3003 1743 3093
rect 1737 2997 1773 3003
rect 1957 2967 1963 3013
rect 1997 3007 2003 3033
rect 2017 2967 2023 3073
rect 2277 3043 2283 3093
rect 2417 3067 2423 3093
rect 2247 3037 2283 3043
rect 2437 2967 2443 3093
rect 2557 3007 2563 3053
rect 2817 3027 2823 3073
rect 2913 3007 2927 3013
rect 2977 2927 2983 3073
rect 3837 3043 3843 3093
rect 3807 3037 3843 3043
rect 3027 3013 3033 3027
rect 3907 3013 3913 3027
rect 4127 3013 4133 3027
rect 3197 2947 3203 3013
rect 4377 3000 4383 3013
rect 3597 2927 3603 2973
rect 4057 2947 4063 2993
rect 4373 2987 4387 3000
rect 4277 2927 4283 2973
rect 4837 2947 4843 2993
rect 4957 2967 4963 3013
rect 5080 3003 5093 3007
rect 5067 2997 5093 3003
rect 5080 2993 5093 2997
rect 5237 3003 5243 3033
rect 5207 2997 5243 3003
rect 5397 2927 5403 3033
rect -63 2882 30 2898
rect -63 2418 -3 2882
rect 1233 2800 1247 2813
rect 17 2747 23 2793
rect 1237 2787 1243 2800
rect 177 2747 183 2773
rect 373 2767 387 2773
rect 647 2753 653 2767
rect 347 2733 353 2747
rect 977 2727 983 2773
rect 1393 2767 1407 2773
rect 1337 2740 1373 2743
rect 1333 2737 1373 2740
rect 1333 2727 1347 2737
rect 1617 2727 1623 2853
rect 1877 2767 1883 2853
rect 2117 2787 2123 2813
rect 1997 2707 2003 2753
rect 2257 2743 2263 2773
rect 2533 2767 2547 2773
rect 2257 2737 2293 2743
rect 2607 2737 2643 2743
rect 2637 2707 2643 2737
rect 2657 2737 2693 2743
rect 2657 2687 2663 2737
rect 3377 2743 3383 2793
rect 3553 2787 3567 2793
rect 3547 2773 3553 2787
rect 3377 2737 3413 2743
rect 3153 2727 3167 2733
rect 3777 2707 3783 2853
rect 4533 2800 4547 2813
rect 3933 2787 3947 2793
rect 4537 2787 4543 2800
rect 3807 2733 3813 2747
rect 4697 2727 4703 2753
rect 4717 2707 4723 2833
rect 4997 2707 5003 2813
rect 5167 2733 5173 2747
rect 5237 2707 5243 2853
rect 5433 2823 5447 2833
rect 5417 2820 5447 2823
rect 5417 2817 5443 2820
rect 5293 2767 5307 2773
rect 5337 2687 5343 2813
rect 5417 2787 5423 2817
rect 5557 2747 5563 2813
rect 5697 2807 5703 2833
rect 5667 2737 5703 2743
rect 5697 2687 5703 2737
rect 5723 2658 5783 3122
rect 5690 2642 5783 2658
rect 267 2553 273 2567
rect 67 2513 73 2527
rect 317 2507 323 2573
rect 337 2567 343 2613
rect 860 2603 873 2607
rect 857 2593 873 2603
rect 627 2563 640 2567
rect 627 2557 653 2563
rect 627 2553 640 2557
rect 757 2543 763 2573
rect 857 2547 863 2593
rect 757 2537 793 2543
rect 347 2513 353 2527
rect 757 2447 763 2537
rect 887 2513 893 2527
rect 977 2517 1013 2523
rect 977 2447 983 2517
rect 1217 2447 1223 2613
rect 2267 2553 2273 2567
rect 2377 2563 2383 2613
rect 2767 2573 2773 2587
rect 2377 2557 2413 2563
rect 2637 2557 2673 2563
rect 1407 2533 1413 2547
rect 1857 2537 1893 2543
rect 1567 2523 1580 2527
rect 1567 2517 1593 2523
rect 1567 2513 1580 2517
rect 1857 2467 1863 2537
rect 1957 2517 1993 2523
rect 1957 2447 1963 2517
rect 2637 2507 2643 2557
rect 2807 2533 2813 2547
rect 2837 2467 2843 2613
rect 3237 2557 3273 2563
rect 3237 2507 3243 2557
rect 3377 2547 3383 2613
rect 3517 2563 3523 2593
rect 3487 2557 3523 2563
rect 3537 2547 3543 2573
rect 3787 2557 3823 2563
rect 3377 2467 3383 2533
rect 3677 2527 3683 2553
rect 3817 2467 3823 2557
rect 4077 2527 4083 2613
rect 4547 2553 4553 2567
rect 4607 2557 4643 2563
rect 4217 2447 4223 2553
rect 4397 2523 4403 2553
rect 4397 2517 4433 2523
rect 4637 2447 4643 2557
rect 5067 2553 5073 2567
rect 4807 2533 4813 2547
rect 4687 2513 4693 2527
rect 4877 2467 4883 2533
rect 5517 2467 5523 2593
rect 5637 2527 5643 2593
rect 5697 2467 5703 2613
rect -63 2402 30 2418
rect -63 1938 -3 2402
rect 457 2297 493 2303
rect 457 2207 463 2297
rect 1047 2293 1053 2307
rect 1157 2297 1193 2303
rect 1157 2247 1163 2297
rect 1657 2267 1663 2333
rect 1817 2247 1823 2373
rect 2393 2307 2407 2313
rect 2217 2257 2253 2263
rect 2217 2207 2223 2257
rect 2557 2227 2563 2353
rect 2677 2307 2683 2373
rect 3317 2347 3323 2373
rect 2660 2303 2673 2307
rect 2647 2297 2673 2303
rect 2660 2293 2673 2297
rect 2847 2273 2853 2287
rect 2917 2267 2923 2333
rect 2767 2253 2773 2267
rect 3197 2257 3233 2263
rect 2873 2227 2887 2233
rect 3197 2207 3203 2257
rect 3317 2263 3323 2333
rect 3317 2257 3353 2263
rect 3437 2263 3443 2333
rect 3657 2283 3663 2313
rect 3627 2277 3663 2283
rect 3817 2267 3823 2373
rect 3437 2257 3473 2263
rect 3437 2227 3443 2257
rect 4057 2207 4063 2373
rect 4077 2207 4083 2253
rect 4337 2227 4343 2353
rect 4617 2327 4623 2373
rect 4757 2267 4763 2313
rect 4777 2207 4783 2273
rect 5177 2267 5183 2313
rect 4927 2253 4933 2267
rect 5357 2207 5363 2333
rect 5637 2327 5643 2373
rect 5587 2277 5623 2283
rect 5617 2207 5623 2277
rect 5723 2178 5783 2642
rect 5690 2162 5783 2178
rect 347 2073 353 2087
rect 267 2033 273 2047
rect 457 1967 463 2133
rect 597 2077 633 2083
rect 597 1967 603 2077
rect 1407 2053 1413 2067
rect 2737 2060 2773 2063
rect 2733 2057 2773 2060
rect 837 2007 843 2053
rect 2733 2047 2747 2057
rect 1127 2033 1133 2047
rect 1237 2037 1273 2043
rect 1237 2007 1243 2037
rect 2317 2037 2353 2043
rect 1897 2007 1903 2033
rect 2273 2027 2287 2033
rect 2317 1967 2323 2037
rect 2937 2043 2943 2113
rect 2907 2037 2943 2043
rect 2857 2020 2863 2033
rect 2853 2007 2867 2020
rect 2937 1967 2943 2037
rect 3013 2027 3027 2033
rect 3233 2027 3247 2033
rect 3317 1967 3323 2133
rect 3427 2077 3463 2083
rect 3457 1967 3463 2077
rect 3597 2047 3603 2133
rect 3687 2077 3723 2083
rect 3717 1987 3723 2077
rect 3977 2047 3983 2093
rect 3767 2033 3773 2047
rect 4277 1987 4283 2133
rect 4417 2080 4453 2083
rect 4413 2077 4453 2080
rect 4413 2067 4427 2077
rect 4677 2007 4683 2133
rect 5337 2087 5343 2113
rect 5357 2077 5393 2083
rect 4677 1997 4693 2007
rect 4680 1993 4693 1997
rect 4797 1967 4803 2033
rect 4817 2027 4823 2073
rect 4866 2033 4867 2040
rect 4853 2027 4867 2033
rect 5157 2007 5163 2053
rect 5357 2047 5363 2077
rect 5617 2083 5623 2133
rect 5587 2077 5623 2083
rect 5617 1987 5623 2077
rect 5677 1987 5683 2033
rect 5697 1967 5703 2013
rect 5680 1966 5703 1967
rect 5687 1956 5703 1966
rect 5687 1953 5700 1956
rect -63 1922 30 1938
rect -63 1458 -3 1922
rect 297 1823 303 1893
rect 267 1817 303 1823
rect 437 1787 443 1833
rect 687 1817 723 1823
rect 577 1747 583 1773
rect 717 1747 723 1817
rect 827 1817 863 1823
rect 857 1727 863 1817
rect 980 1823 993 1827
rect 967 1817 993 1823
rect 980 1813 993 1817
rect 1107 1773 1113 1787
rect 1137 1747 1143 1873
rect 1297 1783 1303 1893
rect 1467 1793 1473 1807
rect 1297 1777 1333 1783
rect 1567 1773 1573 1787
rect 1537 1727 1543 1753
rect 1777 1747 1783 1853
rect 1827 1793 1833 1807
rect 2057 1727 2063 1893
rect 2833 1840 2847 1853
rect 2837 1827 2843 1840
rect 3197 1827 3203 1893
rect 2557 1787 2563 1813
rect 2327 1773 2333 1787
rect 2797 1747 2803 1793
rect 2917 1787 2923 1813
rect 3057 1787 3063 1813
rect 2993 1767 3007 1773
rect 3437 1747 3443 1813
rect 3577 1807 3583 1893
rect 3467 1773 3473 1787
rect 3527 1777 3563 1783
rect 3557 1727 3563 1777
rect 3717 1747 3723 1893
rect 4407 1803 4420 1807
rect 4407 1797 4433 1803
rect 4407 1793 4420 1797
rect 5017 1787 5023 1833
rect 3967 1773 3973 1787
rect 4740 1783 4752 1787
rect 4727 1777 4752 1783
rect 4740 1773 4752 1777
rect 5157 1727 5163 1813
rect 5277 1727 5283 1813
rect 5297 1727 5303 1873
rect 5447 1773 5453 1787
rect 5537 1727 5543 1873
rect 5677 1787 5683 1813
rect 5697 1727 5703 1893
rect 5157 1717 5173 1727
rect 5160 1713 5173 1717
rect 5687 1717 5703 1727
rect 5687 1713 5700 1717
rect 5723 1698 5783 2162
rect 5690 1682 5783 1698
rect 177 1603 183 1653
rect 177 1597 213 1603
rect 317 1597 353 1603
rect 317 1567 323 1597
rect 766 1593 773 1607
rect 997 1587 1003 1653
rect 1107 1593 1113 1607
rect 1137 1587 1143 1633
rect 597 1557 633 1563
rect 597 1507 603 1557
rect 997 1547 1003 1573
rect 1277 1563 1283 1653
rect 1247 1557 1283 1563
rect 1557 1507 1563 1633
rect 1807 1597 1843 1603
rect 1697 1563 1703 1593
rect 1667 1557 1703 1563
rect 1837 1527 1843 1597
rect 2117 1603 2123 1633
rect 2087 1597 2123 1603
rect 2307 1593 2313 1607
rect 3267 1597 3303 1603
rect 2607 1573 2613 1587
rect 1947 1553 1953 1567
rect 2227 1553 2233 1567
rect 2507 1557 2543 1563
rect 2697 1560 2703 1573
rect 2537 1487 2543 1557
rect 2693 1547 2707 1560
rect 3097 1540 3103 1553
rect 3297 1547 3303 1597
rect 3093 1527 3107 1540
rect 3437 1507 3443 1633
rect 3577 1563 3583 1593
rect 3827 1583 3840 1587
rect 3827 1577 3853 1583
rect 3827 1573 3840 1577
rect 3577 1557 3613 1563
rect 4137 1487 4143 1613
rect 4237 1487 4243 1633
rect 4357 1547 4363 1573
rect 4657 1527 4663 1653
rect 4917 1487 4923 1633
rect 5197 1587 5203 1653
rect 5337 1603 5343 1653
rect 5307 1597 5343 1603
rect 5057 1547 5063 1573
rect 5337 1507 5343 1597
rect 5357 1597 5393 1603
rect 5357 1527 5363 1597
rect 5617 1507 5623 1653
rect 5677 1487 5683 1653
rect -63 1442 30 1458
rect -63 978 -3 1442
rect 4837 1420 4874 1423
rect 4833 1417 4874 1420
rect 280 1343 293 1347
rect 267 1337 293 1343
rect 280 1333 293 1337
rect 407 1333 413 1347
rect 457 1303 463 1413
rect 967 1333 973 1347
rect 457 1297 493 1303
rect 1047 1293 1053 1307
rect 1257 1267 1263 1413
rect 1453 1347 1467 1353
rect 1407 1333 1413 1347
rect 2037 1327 2043 1373
rect 2333 1343 2347 1353
rect 2333 1340 2373 1343
rect 2337 1337 2373 1340
rect 2253 1327 2267 1333
rect 2457 1327 2463 1413
rect 4833 1407 4847 1417
rect 4557 1347 4563 1393
rect 4227 1343 4240 1347
rect 4227 1337 4253 1343
rect 4227 1333 4240 1337
rect 1787 1317 1823 1323
rect 1733 1287 1747 1292
rect 1746 1277 1747 1287
rect 1817 1247 1823 1317
rect 1907 1313 1913 1327
rect 2147 1313 2153 1327
rect 3267 1313 3273 1327
rect 3627 1313 3633 1327
rect 4927 1313 4933 1327
rect 2287 1293 2293 1307
rect 3817 1287 3823 1313
rect 4077 1297 4113 1303
rect 3633 1267 3647 1273
rect 4077 1247 4083 1297
rect 4957 1247 4963 1353
rect 4977 1347 4983 1373
rect 5097 1347 5103 1373
rect 5667 1313 5673 1327
rect 5406 1293 5413 1307
rect 5723 1218 5783 1682
rect 5690 1202 5783 1218
rect 177 1127 183 1173
rect 407 1113 413 1127
rect 577 1123 583 1153
rect 547 1117 583 1123
rect 717 1107 723 1153
rect 1437 1123 1443 1153
rect 1407 1117 1443 1123
rect 1697 1087 1703 1153
rect 687 1073 693 1087
rect 967 1073 973 1087
rect 1267 1073 1273 1087
rect 1837 1027 1843 1153
rect 2187 1113 2193 1127
rect 3227 1113 3233 1127
rect 1907 1093 1913 1107
rect 2927 1093 2933 1107
rect 2047 1080 2083 1083
rect 2047 1077 2087 1080
rect 2073 1067 2087 1077
rect 2607 1073 2613 1087
rect 3257 1007 3263 1133
rect 3397 1067 3403 1113
rect 3417 1007 3423 1133
rect 3577 1067 3583 1153
rect 3607 1093 3613 1107
rect 4157 1047 4163 1153
rect 4487 1093 4493 1107
rect 4707 1093 4713 1107
rect 4827 1093 4833 1107
rect 5047 1093 5053 1107
rect 4187 1083 4200 1087
rect 4187 1077 4213 1083
rect 4187 1073 4200 1077
rect 4373 1067 4387 1073
rect 5097 1067 5103 1133
rect 5237 1007 5243 1173
rect 5377 1027 5383 1153
rect 5497 1047 5503 1173
rect 5637 1067 5643 1113
rect 5657 1007 5663 1153
rect -63 962 30 978
rect -63 498 -3 962
rect 87 833 93 847
rect 257 823 263 933
rect 697 887 703 933
rect 380 863 393 867
rect 367 857 393 863
rect 380 853 393 857
rect 507 853 513 867
rect 787 853 793 867
rect 227 817 263 823
rect 817 807 823 893
rect 927 817 963 823
rect 873 807 887 813
rect 957 767 963 817
rect 977 807 983 933
rect 2227 857 2263 863
rect 1237 807 1243 853
rect 1427 833 1433 847
rect 1488 843 1500 847
rect 1488 837 1513 843
rect 1488 833 1500 837
rect 1827 813 1833 827
rect 1587 793 1593 807
rect 2257 787 2263 857
rect 2417 843 2423 873
rect 2973 847 2987 853
rect 2417 837 2453 843
rect 3037 823 3043 933
rect 3147 857 3183 863
rect 3007 817 3043 823
rect 2953 807 2967 813
rect 2473 787 2487 793
rect 3177 767 3183 857
rect 3407 813 3413 827
rect 3457 767 3463 833
rect 3597 767 3603 853
rect 3628 833 3633 847
rect 4317 807 4323 893
rect 4400 843 4413 847
rect 4387 837 4413 843
rect 4400 833 4413 837
rect 4437 807 4443 893
rect 4577 817 4613 823
rect 3667 793 3673 807
rect 4577 767 4583 817
rect 4717 767 4723 893
rect 4747 853 4753 867
rect 4857 843 4863 893
rect 4857 837 4893 843
rect 5007 833 5014 847
rect 5057 827 5063 933
rect 5197 807 5203 853
rect 5317 767 5323 893
rect 5457 767 5463 933
rect 5673 860 5687 873
rect 5677 847 5683 860
rect 3457 757 3473 767
rect 3460 753 3473 757
rect 5723 738 5783 1202
rect 5690 722 5783 738
rect 507 633 513 647
rect 557 643 563 673
rect 557 637 593 643
rect 87 613 93 627
rect 727 593 733 607
rect 837 597 873 603
rect 837 567 843 597
rect 977 587 983 613
rect 1197 600 1203 613
rect 1193 587 1207 600
rect 1237 527 1243 653
rect 1397 627 1403 673
rect 2487 653 2493 667
rect 1547 643 1560 647
rect 1547 637 1573 643
rect 1547 633 1560 637
rect 1677 607 1683 653
rect 1867 613 1873 627
rect 2507 613 2513 627
rect 1397 597 1433 603
rect 1397 567 1403 597
rect 2007 593 2013 607
rect 2057 597 2093 603
rect 2057 547 2063 597
rect 2377 567 2383 613
rect 2577 527 2583 633
rect 2857 627 2863 673
rect 2857 597 2893 603
rect 2857 547 2863 597
rect 3117 527 3123 673
rect 3257 617 3293 623
rect 3257 567 3263 617
rect 3357 607 3363 673
rect 3487 643 3500 647
rect 3487 637 3513 643
rect 3487 633 3500 637
rect 3737 607 3743 673
rect 4117 607 4123 633
rect 3847 593 3853 607
rect 3437 580 3443 593
rect 3433 567 3447 580
rect 4477 527 4483 673
rect 4953 667 4967 673
rect 4587 637 4623 643
rect 4617 587 4623 637
rect 5117 627 5123 693
rect 4927 613 4933 627
rect 5467 613 5473 627
rect 5667 613 5673 627
rect 5167 593 5173 607
rect 5573 587 5587 593
rect -63 482 30 498
rect -63 18 -3 482
rect 757 387 763 433
rect 37 377 73 383
rect 37 287 43 377
rect 927 373 933 387
rect 297 343 303 373
rect 597 347 603 373
rect 267 337 303 343
rect 297 307 303 337
rect 327 333 333 347
rect 1157 343 1163 393
rect 1177 347 1183 453
rect 1317 347 1323 453
rect 1347 373 1353 387
rect 1127 337 1163 343
rect 1457 343 1463 433
rect 1873 367 1887 373
rect 1457 337 1493 343
rect 1627 333 1633 347
rect 1977 343 1983 433
rect 2117 383 2123 413
rect 2087 377 2123 383
rect 2337 363 2343 413
rect 2447 377 2483 383
rect 2477 367 2483 377
rect 2527 373 2533 387
rect 2737 367 2743 453
rect 3827 373 3833 387
rect 2307 357 2343 363
rect 2477 357 2493 367
rect 2480 353 2493 357
rect 1947 337 1983 343
rect 2877 343 2883 373
rect 3347 353 3353 367
rect 4127 353 4133 367
rect 4437 347 4443 433
rect 4677 383 4683 413
rect 4677 377 4713 383
rect 4937 367 4943 433
rect 5077 377 5113 383
rect 2847 337 2883 343
rect 3640 343 3653 347
rect 3627 337 3653 343
rect 3640 333 3653 337
rect 4907 337 4943 343
rect 1073 327 1087 333
rect 2097 287 2103 333
rect 3307 313 3313 327
rect 4937 307 4943 337
rect 5077 287 5083 377
rect 5227 383 5240 387
rect 5227 377 5253 383
rect 5227 373 5240 377
rect 5357 327 5363 413
rect 5497 347 5503 413
rect 5667 353 5673 367
rect 5723 258 5783 722
rect 5690 242 5783 258
rect 87 133 93 147
rect 1007 133 1013 147
rect 227 117 263 123
rect 257 47 263 117
rect 647 113 653 127
rect 800 123 813 127
rect 787 117 813 123
rect 800 113 813 117
rect 1077 123 1083 173
rect 1453 168 1467 173
rect 1307 154 1313 167
rect 1307 153 1323 154
rect 1537 143 1543 193
rect 2647 173 2653 187
rect 3447 177 3483 183
rect 3257 157 3293 163
rect 1507 137 1543 143
rect 1780 143 1793 147
rect 1767 137 1793 143
rect 1780 133 1793 137
rect 2007 133 2013 147
rect 2627 133 2633 147
rect 927 117 963 123
rect 1077 117 1113 123
rect 957 87 963 117
rect 2547 113 2553 127
rect 3257 67 3263 157
rect 3477 147 3483 177
rect 4087 153 4093 167
rect 4117 157 4153 163
rect 3407 133 3413 147
rect 3597 87 3603 133
rect 3747 113 3753 127
rect 4117 87 4123 157
rect 4357 147 4363 173
rect 5357 163 5363 213
rect 5327 157 5363 163
rect 5497 163 5503 193
rect 5497 157 5533 163
rect 4667 133 4673 147
rect 5667 133 5673 147
rect 4497 120 4533 123
rect 4493 117 4533 120
rect 4493 107 4507 117
rect 4737 117 4773 123
rect 4737 87 4743 117
rect -63 2 30 18
rect 5723 2 5783 242
<< m2contact >>
rect 1233 5733 1247 5747
rect 833 5673 847 5687
rect 113 5653 127 5667
rect 213 5653 227 5667
rect 93 5633 107 5647
rect 133 5633 147 5647
rect 193 5633 207 5647
rect 233 5633 247 5647
rect 913 5653 927 5667
rect 333 5633 347 5647
rect 373 5633 387 5647
rect 492 5633 506 5647
rect 533 5633 547 5647
rect 633 5633 647 5647
rect 673 5633 687 5647
rect 753 5633 767 5647
rect 894 5633 908 5647
rect 933 5633 947 5647
rect 1013 5633 1027 5647
rect 1053 5633 1067 5647
rect 1133 5633 1147 5647
rect 1173 5633 1187 5647
rect 353 5613 367 5627
rect 413 5613 427 5627
rect 473 5613 487 5627
rect 514 5613 528 5627
rect 654 5613 668 5627
rect 693 5613 707 5627
rect 993 5613 1007 5627
rect 1033 5613 1047 5627
rect 1153 5613 1167 5627
rect 1773 5673 1787 5687
rect 3733 5673 3747 5687
rect 1393 5653 1407 5667
rect 1453 5653 1467 5667
rect 1513 5653 1527 5667
rect 1573 5653 1587 5667
rect 1313 5633 1327 5647
rect 1373 5633 1387 5647
rect 1413 5633 1427 5647
rect 1553 5633 1567 5647
rect 1593 5633 1607 5647
rect 1634 5633 1648 5647
rect 1673 5633 1687 5647
rect 1713 5633 1727 5647
rect 2513 5653 2527 5667
rect 2753 5653 2767 5667
rect 2913 5653 2927 5667
rect 2953 5653 2967 5667
rect 2993 5653 3007 5667
rect 1913 5633 1927 5647
rect 1953 5633 1967 5647
rect 2033 5633 2047 5647
rect 2154 5633 2168 5647
rect 2413 5633 2427 5647
rect 2454 5633 2468 5647
rect 293 5593 307 5607
rect 793 5593 807 5607
rect 1313 5593 1327 5607
rect 2573 5633 2587 5647
rect 2653 5633 2667 5647
rect 2693 5633 2707 5647
rect 1693 5613 1707 5627
rect 1733 5613 1747 5627
rect 1933 5613 1947 5627
rect 1973 5613 1987 5627
rect 2193 5613 2207 5627
rect 2293 5613 2307 5627
rect 2333 5613 2347 5627
rect 2433 5613 2447 5627
rect 2473 5613 2487 5627
rect 2513 5613 2527 5627
rect 2633 5613 2647 5627
rect 2673 5613 2687 5627
rect 2813 5633 2827 5647
rect 2853 5633 2867 5647
rect 2933 5633 2947 5647
rect 2833 5613 2847 5627
rect 1833 5593 1847 5607
rect 2033 5593 2047 5607
rect 2214 5593 2228 5607
rect 2314 5593 2328 5607
rect 2573 5593 2587 5607
rect 3113 5633 3127 5647
rect 3053 5613 3067 5627
rect 3233 5653 3247 5667
rect 3433 5653 3447 5667
rect 3473 5653 3487 5667
rect 3513 5653 3527 5667
rect 3213 5633 3227 5647
rect 3253 5633 3267 5647
rect 3313 5633 3327 5647
rect 3453 5633 3467 5647
rect 3033 5593 3047 5607
rect 3153 5593 3167 5607
rect 3353 5593 3367 5607
rect 2993 5573 3007 5587
rect 3553 5633 3567 5647
rect 4749 5713 4763 5727
rect 4213 5653 4227 5667
rect 4272 5653 4286 5667
rect 4313 5653 4327 5667
rect 4293 5633 4307 5647
rect 4833 5633 4847 5647
rect 4912 5633 4926 5647
rect 5173 5633 5187 5647
rect 5233 5633 5247 5647
rect 5553 5633 5567 5647
rect 4893 5613 4907 5627
rect 4933 5613 4947 5627
rect 5013 5613 5027 5627
rect 5073 5613 5087 5627
rect 5293 5613 5307 5627
rect 5372 5613 5386 5627
rect 5413 5613 5427 5627
rect 5573 5613 5587 5627
rect 5033 5593 5047 5607
rect 5113 5593 5127 5607
rect 5252 5593 5266 5607
rect 33 5553 47 5567
rect 1633 5553 1647 5567
rect 3513 5553 3527 5567
rect 593 5493 607 5507
rect 5073 5493 5087 5507
rect 453 5473 467 5487
rect 33 5433 47 5447
rect 113 5433 127 5447
rect 313 5433 327 5447
rect 373 5433 387 5447
rect 413 5433 427 5447
rect 93 5413 107 5427
rect 133 5413 147 5427
rect 233 5413 247 5427
rect 273 5413 287 5427
rect 513 5433 527 5447
rect 554 5433 568 5447
rect 353 5413 367 5427
rect 393 5413 407 5427
rect 453 5413 467 5427
rect 493 5413 507 5427
rect 533 5413 547 5427
rect 833 5473 847 5487
rect 4133 5473 4147 5487
rect 653 5453 667 5467
rect 1073 5453 1087 5467
rect 2373 5453 2387 5467
rect 2573 5453 2587 5467
rect 3053 5453 3067 5467
rect 3153 5453 3167 5467
rect 4033 5453 4047 5467
rect 4373 5453 4387 5467
rect 5013 5453 5027 5467
rect 913 5433 927 5447
rect 1053 5433 1067 5447
rect 1273 5433 1287 5447
rect 1313 5433 1327 5447
rect 1353 5433 1367 5447
rect 713 5413 727 5427
rect 753 5413 767 5427
rect 893 5413 907 5427
rect 933 5413 947 5427
rect 993 5413 1007 5427
rect 1153 5413 1167 5427
rect 1293 5413 1307 5427
rect 1333 5413 1347 5427
rect 1433 5413 1447 5427
rect 1533 5413 1547 5427
rect 1573 5413 1587 5427
rect 1673 5413 1687 5427
rect 1713 5413 1727 5427
rect 1853 5413 1867 5427
rect 1973 5413 1987 5427
rect 2013 5413 2027 5427
rect 2074 5413 2088 5427
rect 2113 5413 2127 5427
rect 2233 5413 2247 5427
rect 2392 5413 2406 5427
rect 2433 5413 2447 5427
rect 2473 5413 2487 5427
rect 2613 5413 2627 5427
rect 2713 5413 2727 5427
rect 2753 5413 2767 5427
rect 2853 5413 2867 5427
rect 2893 5413 2907 5427
rect 2993 5413 3007 5427
rect 3133 5433 3147 5447
rect 3374 5433 3388 5447
rect 3413 5433 3427 5447
rect 3573 5433 3587 5447
rect 3633 5433 3647 5447
rect 3673 5433 3687 5447
rect 3173 5413 3187 5427
rect 3233 5413 3247 5427
rect 3353 5413 3367 5427
rect 3393 5413 3407 5427
rect 3513 5413 3527 5427
rect 253 5393 267 5407
rect 313 5393 327 5407
rect 733 5393 747 5407
rect 173 5353 187 5367
rect 1133 5393 1147 5407
rect 1173 5393 1187 5407
rect 1413 5393 1427 5407
rect 1453 5393 1467 5407
rect 1553 5393 1567 5407
rect 1233 5373 1247 5387
rect 813 5333 827 5347
rect 1233 5333 1247 5347
rect 1693 5393 1707 5407
rect 1833 5393 1847 5407
rect 1873 5393 1887 5407
rect 1933 5393 1947 5407
rect 1993 5393 2007 5407
rect 2093 5393 2107 5407
rect 2172 5393 2186 5407
rect 2213 5393 2227 5407
rect 2253 5393 2267 5407
rect 2453 5393 2467 5407
rect 1873 5373 1887 5387
rect 2673 5393 2687 5407
rect 2733 5393 2747 5407
rect 2793 5393 2807 5407
rect 2872 5393 2886 5407
rect 2973 5393 2987 5407
rect 3013 5393 3027 5407
rect 3612 5413 3626 5427
rect 3653 5413 3667 5427
rect 3772 5413 3786 5427
rect 3212 5393 3226 5407
rect 3253 5393 3267 5407
rect 3493 5393 3507 5407
rect 3533 5393 3547 5407
rect 3573 5393 3587 5407
rect 3752 5393 3766 5407
rect 3794 5393 3808 5407
rect 3053 5373 3067 5387
rect 3173 5373 3187 5387
rect 1773 5353 1787 5367
rect 2533 5353 2547 5367
rect 3913 5433 3927 5447
rect 3973 5433 3987 5447
rect 4432 5433 4446 5447
rect 4474 5433 4488 5447
rect 4573 5433 4587 5447
rect 4613 5433 4627 5447
rect 4713 5433 4727 5447
rect 4754 5433 4768 5447
rect 4853 5433 4867 5447
rect 4933 5433 4947 5447
rect 4993 5433 5007 5447
rect 5033 5433 5047 5447
rect 3893 5413 3907 5427
rect 3933 5413 3947 5427
rect 4013 5413 4027 5427
rect 4133 5413 4147 5427
rect 4193 5413 4207 5427
rect 4234 5413 4248 5427
rect 4213 5393 4227 5407
rect 3973 5373 3987 5387
rect 4453 5413 4467 5427
rect 4493 5413 4507 5427
rect 4593 5413 4607 5427
rect 4634 5413 4648 5427
rect 4673 5413 4687 5427
rect 4733 5413 4747 5427
rect 4773 5413 4787 5427
rect 4893 5413 4907 5427
rect 4313 5373 4327 5387
rect 4673 5353 4687 5367
rect 4293 5333 4307 5347
rect 5133 5453 5147 5467
rect 5232 5453 5246 5467
rect 5513 5453 5527 5467
rect 5113 5433 5127 5447
rect 5153 5433 5167 5447
rect 5253 5433 5267 5447
rect 5373 5433 5387 5447
rect 5413 5433 5427 5447
rect 5453 5433 5467 5447
rect 5293 5413 5307 5427
rect 5393 5413 5407 5427
rect 5433 5413 5447 5427
rect 5553 5433 5567 5447
rect 5593 5433 5607 5447
rect 5633 5433 5647 5447
rect 5574 5413 5588 5427
rect 5612 5413 5626 5427
rect 5513 5373 5527 5387
rect 1633 5313 1647 5327
rect 3053 5313 3067 5327
rect 3832 5313 3846 5327
rect 5073 5313 5087 5327
rect 153 5253 167 5267
rect 1773 5253 1787 5267
rect 3193 5253 3207 5267
rect 4413 5253 4427 5267
rect 73 5133 87 5147
rect 113 5133 127 5147
rect 273 5233 287 5247
rect 273 5193 287 5207
rect 973 5193 987 5207
rect 193 5173 207 5187
rect 233 5173 247 5187
rect 453 5173 467 5187
rect 513 5173 527 5187
rect 693 5173 707 5187
rect 213 5153 227 5167
rect 273 5153 287 5167
rect 333 5153 347 5167
rect 373 5153 387 5167
rect 433 5153 447 5167
rect 473 5153 487 5167
rect 613 5153 627 5167
rect 733 5153 747 5167
rect 774 5153 788 5167
rect 872 5153 886 5167
rect 914 5153 928 5167
rect 313 5133 327 5147
rect 353 5133 367 5147
rect 573 5133 587 5147
rect 653 5133 667 5147
rect 694 5133 708 5147
rect 753 5133 767 5147
rect 793 5133 807 5147
rect 853 5133 867 5147
rect 892 5133 906 5147
rect 1393 5173 1407 5187
rect 1453 5173 1467 5187
rect 1533 5173 1547 5187
rect 1573 5173 1587 5187
rect 1852 5173 1866 5187
rect 1933 5173 1947 5187
rect 1973 5173 1987 5187
rect 2593 5173 2607 5187
rect 2653 5173 2667 5187
rect 2833 5173 2847 5187
rect 2873 5173 2887 5187
rect 2913 5173 2927 5187
rect 2952 5173 2966 5187
rect 2993 5173 3007 5187
rect 3093 5173 3107 5187
rect 3153 5173 3167 5187
rect 4272 5233 4286 5247
rect 3453 5213 3467 5227
rect 3273 5173 3287 5187
rect 1033 5153 1047 5167
rect 1293 5153 1307 5167
rect 1333 5153 1347 5167
rect 1433 5153 1447 5167
rect 1473 5153 1487 5167
rect 1552 5153 1566 5167
rect 1693 5153 1707 5167
rect 1833 5153 1847 5167
rect 1873 5153 1887 5167
rect 1953 5153 1967 5167
rect 2073 5153 2087 5167
rect 2113 5153 2127 5167
rect 2213 5153 2227 5167
rect 2253 5153 2267 5167
rect 2493 5153 2507 5167
rect 2633 5153 2647 5167
rect 2673 5153 2687 5167
rect 2733 5153 2747 5167
rect 2853 5153 2867 5167
rect 2973 5153 2987 5167
rect 3073 5153 3087 5167
rect 3113 5153 3127 5167
rect 3253 5153 3267 5167
rect 3293 5153 3307 5167
rect 3353 5153 3367 5167
rect 3393 5153 3407 5167
rect 1073 5133 1087 5147
rect 1133 5133 1147 5147
rect 1172 5133 1186 5147
rect 1253 5133 1267 5147
rect 1313 5133 1327 5147
rect 1653 5133 1667 5147
rect 1733 5133 1747 5147
rect 2093 5133 2107 5147
rect 2133 5133 2147 5147
rect 2233 5133 2247 5147
rect 2273 5133 2287 5147
rect 2332 5133 2346 5147
rect 2374 5133 2388 5147
rect 2453 5133 2467 5147
rect 2513 5133 2527 5147
rect 2913 5133 2927 5147
rect 3372 5133 3386 5147
rect 3413 5133 3427 5147
rect 93 5113 107 5127
rect 153 5113 167 5127
rect 1152 5113 1166 5127
rect 2352 5113 2366 5127
rect 2733 5113 2747 5127
rect 3753 5193 3767 5207
rect 4254 5193 4268 5207
rect 3513 5153 3527 5167
rect 3553 5153 3567 5167
rect 3613 5153 3627 5167
rect 3653 5153 3667 5167
rect 3692 5153 3706 5167
rect 3533 5133 3547 5147
rect 3573 5133 3587 5147
rect 3673 5133 3687 5147
rect 3714 5133 3728 5147
rect 3813 5153 3827 5167
rect 3913 5153 3927 5167
rect 4153 5153 4167 5167
rect 4194 5153 4208 5167
rect 3853 5133 3867 5147
rect 4013 5133 4027 5147
rect 4053 5133 4067 5147
rect 4132 5133 4146 5147
rect 4173 5133 4187 5147
rect 4213 5133 4227 5147
rect 3613 5113 3627 5127
rect 3953 5113 3967 5127
rect 4033 5113 4047 5127
rect 4332 5153 4346 5167
rect 4373 5153 4387 5167
rect 4493 5233 4507 5247
rect 5117 5233 5131 5247
rect 4353 5133 4367 5147
rect 5533 5213 5547 5227
rect 4552 5153 4566 5167
rect 4593 5153 4607 5167
rect 4713 5153 4727 5167
rect 4753 5153 4767 5167
rect 4833 5153 4847 5167
rect 4873 5153 4887 5167
rect 4993 5153 5007 5167
rect 5033 5153 5047 5167
rect 4533 5133 4547 5147
rect 4573 5133 4587 5147
rect 4613 5133 4627 5147
rect 4693 5133 4707 5147
rect 4733 5133 4747 5147
rect 4853 5133 4867 5147
rect 4893 5133 4907 5147
rect 4973 5133 4987 5147
rect 5013 5133 5027 5147
rect 5653 5153 5667 5167
rect 4353 5113 4367 5127
rect 4433 5113 4447 5127
rect 4493 5113 4507 5127
rect 5533 5113 5547 5127
rect 5593 5113 5607 5127
rect 4253 5093 4267 5107
rect 3453 5073 3467 5087
rect 153 5013 167 5027
rect 573 5013 587 5027
rect 1193 5013 1207 5027
rect 2533 5013 2547 5027
rect 4013 5013 4027 5027
rect 93 4933 107 4947
rect 73 4913 87 4927
rect 113 4913 127 4927
rect 433 4993 447 5007
rect 213 4953 227 4967
rect 253 4953 267 4967
rect 313 4953 327 4967
rect 354 4953 368 4967
rect 193 4933 207 4947
rect 234 4933 248 4947
rect 333 4933 347 4947
rect 373 4933 387 4947
rect 453 4953 467 4967
rect 513 4953 527 4967
rect 493 4933 507 4947
rect 533 4933 547 4947
rect 1353 4993 1367 5007
rect 853 4973 867 4987
rect 1173 4973 1187 4987
rect 1213 4973 1227 4987
rect 633 4933 647 4947
rect 673 4933 687 4947
rect 753 4933 767 4947
rect 893 4933 907 4947
rect 952 4933 966 4947
rect 994 4933 1008 4947
rect 1113 4933 1127 4947
rect 1513 4973 1527 4987
rect 1713 4973 1727 4987
rect 2033 4973 2047 4987
rect 2233 4973 2247 4987
rect 2473 4973 2487 4987
rect 1233 4953 1247 4967
rect 1353 4953 1367 4967
rect 1493 4953 1507 4967
rect 1533 4953 1547 4967
rect 2013 4953 2027 4967
rect 2212 4953 2226 4967
rect 2252 4953 2266 4967
rect 2372 4953 2386 4967
rect 2414 4953 2428 4967
rect 1273 4933 1287 4947
rect 1393 4933 1407 4947
rect 1633 4933 1647 4947
rect 1753 4933 1767 4947
rect 1853 4933 1867 4947
rect 1893 4933 1907 4947
rect 593 4913 607 4927
rect 652 4913 666 4927
rect 733 4913 747 4927
rect 773 4913 787 4927
rect 973 4913 987 4927
rect 1013 4913 1027 4927
rect 1093 4913 1107 4927
rect 1133 4913 1147 4927
rect 1173 4913 1187 4927
rect 1373 4913 1387 4927
rect 1413 4913 1427 4927
rect 1613 4913 1627 4927
rect 1653 4913 1667 4927
rect 1813 4913 1827 4927
rect 1874 4913 1888 4927
rect 2113 4933 2127 4947
rect 2353 4933 2367 4947
rect 2393 4933 2407 4947
rect 2613 4993 2627 5007
rect 2613 4973 2627 4987
rect 2693 4973 2707 4987
rect 3353 4973 3367 4987
rect 3833 4973 3847 4987
rect 3953 4973 3967 4987
rect 4194 4973 4208 4987
rect 4333 4973 4347 4987
rect 4414 4973 4428 4987
rect 4534 4973 4548 4987
rect 5293 4973 5307 4987
rect 2674 4953 2688 4967
rect 2714 4953 2728 4967
rect 2952 4953 2966 4967
rect 2993 4953 3007 4967
rect 3213 4953 3227 4967
rect 3254 4953 3268 4967
rect 3433 4953 3447 4967
rect 3473 4953 3487 4967
rect 3513 4953 3527 4967
rect 3813 4953 3827 4967
rect 3853 4953 3867 4967
rect 3933 4953 3947 4967
rect 3973 4953 3987 4967
rect 4013 4953 4027 4967
rect 4093 4953 4107 4967
rect 4134 4953 4148 4967
rect 4393 4953 4407 4967
rect 4433 4953 4447 4967
rect 4514 4953 4528 4967
rect 4553 4953 4567 4967
rect 4613 4953 4627 4967
rect 4733 4953 4747 4967
rect 4813 4953 4827 4967
rect 4853 4953 4867 4967
rect 5153 4953 5167 4967
rect 5193 4953 5207 4967
rect 5333 4953 5347 4967
rect 5393 4953 5407 4967
rect 2633 4933 2647 4947
rect 2813 4933 2827 4947
rect 2873 4933 2887 4947
rect 2933 4933 2947 4947
rect 2973 4933 2987 4947
rect 3073 4933 3087 4947
rect 3193 4933 3207 4947
rect 3233 4933 3247 4947
rect 3373 4933 3387 4947
rect 3453 4933 3467 4947
rect 3493 4933 3507 4947
rect 3593 4933 3607 4947
rect 3713 4933 3727 4947
rect 3773 4933 3787 4947
rect 2093 4913 2107 4927
rect 2133 4913 2147 4927
rect 2793 4913 2807 4927
rect 2833 4913 2847 4927
rect 693 4893 707 4907
rect 1933 4893 1947 4907
rect 3053 4913 3067 4927
rect 3093 4913 3107 4927
rect 3573 4913 3587 4927
rect 3613 4913 3627 4927
rect 4073 4933 4087 4947
rect 4113 4933 4127 4947
rect 4313 4933 4327 4947
rect 4673 4933 4687 4947
rect 5013 4933 5027 4947
rect 5133 4933 5147 4947
rect 5172 4933 5186 4947
rect 5273 4933 5287 4947
rect 4653 4913 4667 4927
rect 4693 4913 4707 4927
rect 4953 4913 4967 4927
rect 4993 4913 5007 4927
rect 5033 4913 5047 4927
rect 4473 4893 4487 4907
rect 4613 4893 4627 4907
rect 4253 4873 4267 4887
rect 153 4853 167 4867
rect 433 4853 447 4867
rect 573 4853 587 4867
rect 693 4853 707 4867
rect 2873 4853 2887 4867
rect 4013 4853 4027 4867
rect 4473 4853 4487 4867
rect 5513 4953 5527 4967
rect 5494 4933 5508 4947
rect 5533 4933 5547 4947
rect 5633 4933 5647 4947
rect 5613 4913 5627 4927
rect 5653 4913 5667 4927
rect 4953 4833 4967 4847
rect 5433 4833 5447 4847
rect 2653 4773 2667 4787
rect 393 4733 407 4747
rect 2613 4733 2627 4747
rect 113 4693 127 4707
rect 2213 4713 2227 4727
rect 634 4693 648 4707
rect 93 4673 107 4687
rect 133 4673 147 4687
rect 192 4673 206 4687
rect 233 4673 247 4687
rect 353 4673 367 4687
rect 394 4673 408 4687
rect 493 4673 507 4687
rect 533 4673 547 4687
rect 613 4673 627 4687
rect 653 4673 667 4687
rect 213 4653 227 4667
rect 273 4653 287 4667
rect 333 4653 347 4667
rect 373 4653 387 4667
rect 473 4653 487 4667
rect 513 4653 527 4667
rect 33 4633 47 4647
rect 773 4693 787 4707
rect 753 4673 767 4687
rect 793 4673 807 4687
rect 993 4693 1007 4707
rect 1193 4693 1207 4707
rect 1233 4693 1247 4707
rect 1313 4693 1327 4707
rect 893 4673 907 4687
rect 933 4673 947 4687
rect 912 4653 926 4667
rect 1053 4673 1067 4687
rect 1093 4673 1107 4687
rect 1213 4673 1227 4687
rect 1293 4673 1307 4687
rect 1333 4673 1347 4687
rect 1033 4653 1047 4667
rect 1073 4653 1087 4667
rect 1553 4693 1567 4707
rect 1614 4693 1628 4707
rect 1853 4693 1867 4707
rect 1913 4693 1927 4707
rect 1593 4673 1607 4687
rect 1633 4673 1647 4687
rect 1713 4673 1727 4687
rect 1753 4673 1767 4687
rect 1893 4673 1907 4687
rect 1934 4673 1948 4687
rect 2033 4673 2047 4687
rect 2073 4673 2087 4687
rect 2133 4673 2147 4687
rect 2573 4693 2587 4707
rect 2613 4693 2627 4707
rect 2353 4673 2367 4687
rect 2393 4673 2407 4687
rect 2513 4673 2527 4687
rect 2592 4673 2606 4687
rect 2873 4713 2887 4727
rect 3773 4713 3787 4727
rect 2873 4693 2887 4707
rect 2913 4693 2927 4707
rect 3233 4693 3247 4707
rect 3292 4693 3306 4707
rect 3353 4693 3367 4707
rect 3393 4693 3407 4707
rect 2733 4673 2747 4687
rect 2773 4673 2787 4687
rect 2893 4673 2907 4687
rect 3053 4673 3067 4687
rect 3153 4673 3167 4687
rect 3213 4673 3227 4687
rect 3253 4673 3267 4687
rect 3373 4673 3387 4687
rect 3513 4673 3527 4687
rect 3613 4673 3627 4687
rect 3813 4693 3827 4707
rect 3853 4693 3867 4707
rect 4153 4693 4167 4707
rect 4193 4693 4207 4707
rect 4513 4693 4527 4707
rect 4553 4693 4567 4707
rect 4973 4693 4987 4707
rect 5013 4693 5027 4707
rect 3833 4673 3847 4687
rect 4173 4673 4187 4687
rect 4533 4673 4547 4687
rect 4653 4673 4667 4687
rect 4993 4673 5007 4687
rect 5113 4673 5127 4687
rect 5153 4673 5167 4687
rect 5373 4673 5387 4687
rect 1453 4653 1467 4667
rect 1493 4653 1507 4667
rect 1692 4653 1706 4667
rect 1734 4653 1748 4667
rect 1774 4653 1788 4667
rect 1992 4653 2006 4667
rect 2052 4653 2066 4667
rect 2332 4653 2346 4667
rect 2374 4653 2388 4667
rect 2493 4653 2507 4667
rect 2653 4653 2667 4667
rect 2713 4653 2727 4667
rect 2752 4653 2766 4667
rect 2793 4653 2807 4667
rect 2993 4653 3007 4667
rect 3473 4653 3487 4667
rect 3673 4653 3687 4667
rect 3713 4653 3727 4667
rect 3773 4653 3787 4667
rect 3912 4653 3926 4667
rect 3954 4653 3968 4667
rect 3993 4653 4007 4667
rect 4033 4653 4047 4667
rect 4073 4653 4087 4667
rect 4313 4653 4327 4667
rect 4353 4653 4367 4667
rect 4433 4653 4447 4667
rect 4713 4653 4727 4667
rect 4793 4653 4807 4667
rect 4833 4653 4847 4667
rect 5133 4653 5147 4667
rect 5193 4653 5207 4667
rect 5233 4653 5247 4667
rect 5293 4653 5307 4667
rect 5492 4653 5506 4667
rect 5533 4653 5547 4667
rect 5613 4653 5627 4667
rect 1472 4633 1486 4647
rect 2133 4633 2147 4647
rect 2233 4633 2247 4647
rect 2973 4633 2987 4647
rect 3153 4633 3167 4647
rect 3573 4633 3587 4647
rect 3693 4633 3707 4647
rect 3932 4633 3946 4647
rect 4053 4633 4067 4647
rect 4633 4633 4647 4647
rect 5393 4633 5407 4647
rect 713 4593 727 4607
rect 853 4593 867 4607
rect 1393 4593 1407 4607
rect 3993 4593 4007 4607
rect 173 4533 187 4547
rect 2153 4533 2167 4547
rect 2333 4533 2347 4547
rect 93 4473 107 4487
rect 133 4473 147 4487
rect 373 4493 387 4507
rect 853 4493 867 4507
rect 1493 4493 1507 4507
rect 253 4473 267 4487
rect 353 4473 367 4487
rect 393 4473 407 4487
rect 1333 4473 1347 4487
rect 1453 4473 1467 4487
rect 1733 4473 1747 4487
rect 1813 4473 1827 4487
rect 1874 4473 1888 4487
rect 2153 4473 2167 4487
rect 2253 4473 2267 4487
rect 2293 4473 2307 4487
rect 73 4453 87 4467
rect 113 4453 127 4467
rect 234 4453 248 4467
rect 273 4453 287 4467
rect 493 4453 507 4467
rect 613 4453 627 4467
rect 653 4453 667 4467
rect 713 4453 727 4467
rect 753 4453 767 4467
rect 893 4453 907 4467
rect 953 4453 967 4467
rect 993 4453 1007 4467
rect 1093 4453 1107 4467
rect 1133 4453 1147 4467
rect 1233 4453 1247 4467
rect 1273 4453 1287 4467
rect 473 4433 487 4447
rect 513 4433 527 4447
rect 633 4433 647 4447
rect 733 4433 747 4447
rect 973 4433 987 4447
rect 813 4393 827 4407
rect 1113 4433 1127 4447
rect 1173 4433 1187 4447
rect 1253 4433 1267 4447
rect 1393 4453 1407 4467
rect 1373 4433 1387 4447
rect 1414 4433 1428 4447
rect 1494 4453 1508 4467
rect 1632 4453 1646 4467
rect 1713 4453 1727 4467
rect 1853 4453 1867 4467
rect 1893 4453 1907 4467
rect 1993 4453 2007 4467
rect 2033 4453 2047 4467
rect 2113 4453 2127 4467
rect 2232 4453 2246 4467
rect 2273 4453 2287 4467
rect 1613 4433 1627 4447
rect 1653 4433 1667 4447
rect 1933 4433 1947 4447
rect 2014 4433 2028 4447
rect 2093 4433 2107 4447
rect 2133 4433 2147 4447
rect 1453 4413 1467 4427
rect 2934 4493 2948 4507
rect 3513 4493 3527 4507
rect 2393 4453 2407 4467
rect 2553 4473 2567 4487
rect 2633 4473 2647 4487
rect 2673 4473 2687 4487
rect 2714 4473 2728 4487
rect 2913 4473 2927 4487
rect 2953 4473 2967 4487
rect 3033 4473 3047 4487
rect 3093 4473 3107 4487
rect 3234 4473 3248 4487
rect 3313 4473 3327 4487
rect 3373 4473 3387 4487
rect 3413 4473 3427 4487
rect 3533 4473 3547 4487
rect 3653 4473 3667 4487
rect 3694 4473 3708 4487
rect 3933 4473 3947 4487
rect 3974 4473 3988 4487
rect 4033 4473 4047 4487
rect 4113 4473 4127 4487
rect 4314 4473 4328 4487
rect 4353 4473 4367 4487
rect 4634 4473 4648 4487
rect 4712 4473 4726 4487
rect 4753 4473 4767 4487
rect 4933 4473 4947 4487
rect 4973 4473 4987 4487
rect 5153 4473 5167 4487
rect 5213 4473 5227 4487
rect 5253 4473 5267 4487
rect 5333 4473 5347 4487
rect 5373 4473 5387 4487
rect 5513 4473 5527 4487
rect 5553 4473 5567 4487
rect 2513 4453 2527 4467
rect 2654 4453 2668 4467
rect 2693 4453 2707 4467
rect 2793 4453 2807 4467
rect 3174 4453 3188 4467
rect 3273 4453 3287 4467
rect 3393 4453 3407 4467
rect 3433 4453 3447 4467
rect 3573 4453 3587 4467
rect 3673 4453 3687 4467
rect 3713 4453 3727 4467
rect 3833 4453 3847 4467
rect 4193 4453 4207 4467
rect 4292 4453 4306 4467
rect 4333 4453 4347 4467
rect 2373 4433 2387 4447
rect 2413 4433 2427 4447
rect 2453 4433 2467 4447
rect 2773 4433 2787 4447
rect 2813 4433 2827 4447
rect 3153 4433 3167 4447
rect 3193 4433 3207 4447
rect 3233 4433 3247 4447
rect 3813 4433 3827 4447
rect 3854 4433 3868 4447
rect 4113 4433 4127 4447
rect 4173 4433 4187 4447
rect 4213 4433 4227 4447
rect 2413 4393 2427 4407
rect 4573 4453 4587 4467
rect 4913 4453 4927 4467
rect 4953 4453 4967 4467
rect 5052 4453 5066 4467
rect 5533 4453 5547 4467
rect 5573 4453 5587 4467
rect 5033 4433 5047 4447
rect 5073 4433 5087 4447
rect 3153 4393 3167 4407
rect 4393 4393 4407 4407
rect 2333 4373 2347 4387
rect 553 4353 567 4367
rect 1053 4353 1067 4367
rect 573 4293 587 4307
rect 1113 4293 1127 4307
rect 2693 4293 2707 4307
rect 193 4213 207 4227
rect 253 4213 267 4227
rect 353 4213 367 4227
rect 393 4213 407 4227
rect 433 4213 447 4227
rect 513 4213 527 4227
rect 93 4193 107 4207
rect 133 4193 147 4207
rect 233 4193 247 4207
rect 273 4193 287 4207
rect 372 4193 386 4207
rect 493 4193 507 4207
rect 533 4193 547 4207
rect 893 4213 907 4227
rect 933 4213 947 4227
rect 613 4193 627 4207
rect 654 4193 668 4207
rect 713 4193 727 4207
rect 773 4193 787 4207
rect 813 4193 827 4207
rect 912 4193 926 4207
rect 1053 4193 1067 4207
rect 73 4173 87 4187
rect 573 4173 587 4187
rect 633 4173 647 4187
rect 674 4173 688 4187
rect 112 4153 126 4167
rect 752 4173 766 4187
rect 794 4173 808 4187
rect 834 4173 848 4187
rect 1013 4173 1027 4187
rect 2393 4273 2407 4287
rect 1613 4253 1627 4267
rect 1373 4233 1387 4247
rect 1153 4213 1167 4227
rect 1212 4213 1226 4227
rect 1193 4193 1207 4207
rect 1233 4193 1247 4207
rect 1293 4193 1307 4207
rect 1513 4193 1527 4207
rect 1553 4193 1567 4207
rect 1533 4173 1547 4187
rect 1573 4173 1587 4187
rect 1333 4153 1347 4167
rect 1433 4153 1447 4167
rect 1633 4213 1647 4227
rect 1693 4213 1707 4227
rect 1773 4213 1787 4227
rect 1814 4213 1828 4227
rect 2033 4213 2047 4227
rect 2073 4213 2087 4227
rect 2413 4233 2427 4247
rect 1673 4193 1687 4207
rect 1714 4193 1728 4207
rect 1792 4193 1806 4207
rect 1912 4193 1926 4207
rect 1953 4193 1967 4207
rect 2052 4193 2066 4207
rect 2173 4193 2187 4207
rect 2213 4193 2227 4207
rect 2314 4193 2328 4207
rect 2353 4193 2367 4207
rect 2393 4193 2407 4207
rect 1933 4173 1947 4187
rect 1973 4173 1987 4187
rect 2134 4173 2148 4187
rect 2193 4173 2207 4187
rect 2233 4173 2247 4187
rect 2293 4173 2307 4187
rect 2333 4173 2347 4187
rect 2473 4193 2487 4207
rect 2593 4193 2607 4207
rect 2634 4193 2648 4207
rect 3093 4273 3107 4287
rect 3233 4273 3247 4287
rect 4053 4273 4067 4287
rect 3013 4213 3027 4227
rect 3053 4213 3067 4227
rect 2753 4193 2767 4207
rect 2793 4193 2807 4207
rect 2433 4173 2447 4187
rect 2513 4173 2527 4187
rect 2573 4173 2587 4187
rect 2613 4173 2627 4187
rect 2653 4173 2667 4187
rect 2694 4173 2708 4187
rect 2732 4173 2746 4187
rect 2772 4173 2786 4187
rect 2814 4173 2828 4187
rect 2413 4153 2427 4167
rect 2893 4153 2907 4167
rect 1633 4133 1647 4147
rect 2133 4133 2147 4147
rect 2693 4133 2707 4147
rect 3033 4193 3047 4207
rect 3153 4193 3167 4207
rect 3193 4173 3207 4187
rect 3653 4213 3667 4227
rect 3693 4213 3707 4227
rect 3753 4213 3767 4227
rect 3793 4213 3807 4227
rect 3893 4213 3907 4227
rect 3933 4213 3947 4227
rect 3272 4193 3286 4207
rect 3314 4193 3328 4207
rect 3413 4193 3427 4207
rect 3453 4193 3467 4207
rect 3533 4193 3547 4207
rect 3673 4193 3687 4207
rect 3773 4193 3787 4207
rect 3913 4193 3927 4207
rect 4013 4193 4027 4207
rect 3294 4173 3308 4187
rect 3333 4173 3347 4187
rect 3392 4173 3406 4187
rect 3433 4173 3447 4187
rect 3233 4153 3247 4167
rect 3573 4153 3587 4167
rect 3993 4153 4007 4167
rect 4173 4253 4187 4267
rect 4173 4213 4187 4227
rect 4213 4213 4227 4227
rect 4253 4213 4267 4227
rect 5333 4213 5347 4227
rect 5373 4213 5387 4227
rect 5473 4213 5487 4227
rect 5513 4213 5527 4227
rect 4093 4173 4107 4187
rect 4233 4193 4247 4207
rect 4352 4193 4366 4207
rect 4392 4193 4406 4207
rect 4573 4193 4587 4207
rect 5213 4193 5227 4207
rect 5253 4193 5267 4207
rect 5353 4193 5367 4207
rect 5492 4193 5506 4207
rect 5593 4193 5607 4207
rect 5633 4193 5647 4207
rect 4373 4173 4387 4187
rect 4413 4173 4427 4187
rect 4453 4173 4467 4187
rect 4533 4173 4547 4187
rect 4712 4173 4726 4187
rect 4773 4173 4787 4187
rect 4873 4173 4887 4187
rect 4913 4173 4927 4187
rect 4993 4173 5007 4187
rect 5073 4173 5087 4187
rect 5152 4173 5166 4187
rect 5193 4173 5207 4187
rect 5233 4173 5247 4187
rect 5573 4173 5587 4187
rect 5613 4173 5627 4187
rect 4053 4133 4067 4147
rect 713 4113 727 4127
rect 2953 4113 2967 4127
rect 2253 4053 2267 4067
rect 4293 4053 4307 4067
rect 5213 4053 5227 4067
rect 5673 4053 5687 4067
rect 693 4033 707 4047
rect 1613 4033 1627 4047
rect 2073 4033 2087 4047
rect 753 4013 767 4027
rect 214 3993 228 4007
rect 273 3993 287 4007
rect 473 3993 487 4007
rect 514 3993 528 4007
rect 693 3993 707 4007
rect 733 3993 747 4007
rect 773 3993 787 4007
rect 1253 3993 1267 4007
rect 1313 3993 1327 4007
rect 93 3973 107 3987
rect 133 3973 147 3987
rect 193 3973 207 3987
rect 233 3973 247 3987
rect 333 3973 347 3987
rect 373 3973 387 3987
rect 493 3973 507 3987
rect 533 3973 547 3987
rect 634 3973 648 3987
rect 73 3953 87 3967
rect 113 3953 127 3967
rect 353 3953 367 3967
rect 413 3953 427 3967
rect 613 3953 627 3967
rect 653 3953 667 3967
rect 873 3973 887 3987
rect 1013 3973 1027 3987
rect 1132 3973 1146 3987
rect 1173 3973 1187 3987
rect 1233 3973 1247 3987
rect 1273 3973 1287 3987
rect 853 3953 867 3967
rect 894 3953 908 3967
rect 993 3953 1007 3967
rect 1033 3953 1047 3967
rect 693 3913 707 3927
rect 1153 3953 1167 3967
rect 1433 3993 1447 4007
rect 1512 3993 1526 4007
rect 1552 3993 1566 4007
rect 1413 3973 1427 3987
rect 1453 3973 1467 3987
rect 1533 3973 1547 3987
rect 1574 3973 1588 3987
rect 1653 4013 1667 4027
rect 1893 3993 1907 4007
rect 1953 3993 1967 4007
rect 2133 3993 2147 4007
rect 2173 3993 2187 4007
rect 2213 3993 2227 4007
rect 2493 4033 2507 4047
rect 2333 3993 2347 4007
rect 2393 3993 2407 4007
rect 1653 3973 1667 3987
rect 1773 3973 1787 3987
rect 1913 3973 1927 3987
rect 2013 3973 2027 3987
rect 2153 3973 2167 3987
rect 2193 3973 2207 3987
rect 1613 3953 1627 3967
rect 1752 3953 1766 3967
rect 1793 3953 1807 3967
rect 2833 4013 2847 4027
rect 2973 4013 2987 4027
rect 3353 4013 3367 4027
rect 3853 4013 3867 4027
rect 2513 3993 2527 4007
rect 2573 3993 2587 4007
rect 2813 3993 2827 4007
rect 2953 3993 2967 4007
rect 3053 3993 3067 4007
rect 3093 3993 3107 4007
rect 3573 3993 3587 4007
rect 3633 3993 3647 4007
rect 3673 3993 3687 4007
rect 3733 3993 3747 4007
rect 3833 3993 3847 4007
rect 3873 3993 3887 4007
rect 3933 3993 3947 4007
rect 3994 3993 4008 4007
rect 2673 3973 2687 3987
rect 2773 3973 2787 3987
rect 2913 3973 2927 3987
rect 3072 3973 3086 3987
rect 3114 3973 3128 3987
rect 3213 3973 3227 3987
rect 3253 3973 3267 3987
rect 3353 3973 3367 3987
rect 3453 3973 3467 3987
rect 3494 3973 3508 3987
rect 3553 3973 3567 3987
rect 3593 3973 3607 3987
rect 3713 3973 3727 3987
rect 3753 3973 3767 3987
rect 3973 3973 3987 3987
rect 4113 3973 4127 3987
rect 5073 4033 5087 4047
rect 4493 3993 4507 4007
rect 4533 3993 4547 4007
rect 4753 3993 4767 4007
rect 4793 3993 4807 4007
rect 4852 3993 4866 4007
rect 4893 3993 4907 4007
rect 5154 3993 5168 4007
rect 4373 3973 4387 3987
rect 4473 3973 4487 3987
rect 4513 3973 4527 3987
rect 4613 3973 4627 3987
rect 4733 3973 4747 3987
rect 4773 3973 4787 3987
rect 4873 3973 4887 3987
rect 4913 3973 4927 3987
rect 5013 3973 5027 3987
rect 5133 3973 5147 3987
rect 5173 3973 5187 3987
rect 2493 3953 2507 3967
rect 2652 3953 2666 3967
rect 2693 3953 2707 3967
rect 3193 3953 3207 3967
rect 3232 3953 3246 3967
rect 3413 3953 3427 3967
rect 3473 3953 3487 3967
rect 2473 3933 2487 3947
rect 4353 3953 4367 3967
rect 4393 3953 4407 3967
rect 4592 3953 4606 3967
rect 4633 3953 4647 3967
rect 4993 3953 5007 3967
rect 5034 3953 5048 3967
rect 4713 3933 4727 3947
rect 1353 3913 1367 3927
rect 4013 3913 4027 3927
rect 4353 3913 4367 3927
rect 5033 3913 5047 3927
rect 1073 3893 1087 3907
rect 4712 3893 4726 3907
rect 5413 4013 5427 4027
rect 5593 3993 5607 4007
rect 5633 3993 5647 4007
rect 5273 3973 5287 3987
rect 5392 3973 5406 3987
rect 5453 3973 5467 3987
rect 5253 3953 5267 3967
rect 5293 3953 5307 3967
rect 5673 3973 5687 3987
rect 5213 3873 5227 3887
rect 5553 3873 5567 3887
rect 1992 3813 2006 3827
rect 2253 3813 2267 3827
rect 293 3753 307 3767
rect 193 3713 207 3727
rect 233 3713 247 3727
rect 332 3713 346 3727
rect 373 3713 387 3727
rect 513 3713 527 3727
rect 593 3713 607 3727
rect 713 3713 727 3727
rect 753 3713 767 3727
rect 53 3693 67 3707
rect 113 3693 127 3707
rect 213 3693 227 3707
rect 253 3693 267 3707
rect 292 3693 306 3707
rect 353 3693 367 3707
rect 394 3693 408 3707
rect 473 3692 487 3706
rect 673 3693 687 3707
rect 733 3693 747 3707
rect 533 3673 547 3687
rect 873 3733 887 3747
rect 1253 3733 1267 3747
rect 1313 3733 1327 3747
rect 853 3713 867 3727
rect 894 3713 908 3727
rect 994 3713 1008 3727
rect 1034 3713 1048 3727
rect 1153 3713 1167 3727
rect 1293 3713 1307 3727
rect 1333 3713 1347 3727
rect 1393 3713 1407 3727
rect 1513 3713 1527 3727
rect 1553 3713 1567 3727
rect 1653 3713 1667 3727
rect 1693 3713 1707 3727
rect 973 3693 987 3707
rect 1014 3693 1028 3707
rect 1053 3693 1067 3707
rect 1193 3693 1207 3707
rect 1533 3693 1547 3707
rect 1573 3693 1587 3707
rect 1674 3693 1688 3707
rect 1713 3693 1727 3707
rect 1433 3673 1447 3687
rect 1833 3693 1847 3707
rect 1913 3693 1927 3707
rect 1953 3693 1967 3707
rect 1853 3673 1867 3687
rect 1933 3673 1947 3687
rect 2072 3773 2086 3787
rect 2113 3773 2127 3787
rect 2033 3733 2047 3747
rect 2074 3733 2088 3747
rect 2053 3713 2067 3727
rect 2193 3713 2207 3727
rect 2153 3693 2167 3707
rect 2993 3793 3007 3807
rect 2953 3773 2967 3787
rect 2413 3733 2427 3747
rect 2453 3733 2467 3747
rect 2653 3733 2667 3747
rect 2693 3733 2707 3747
rect 2913 3733 2927 3747
rect 2993 3733 3007 3747
rect 3573 3733 3587 3747
rect 3633 3733 3647 3747
rect 3713 3733 3727 3747
rect 2433 3713 2447 3727
rect 2533 3713 2547 3727
rect 2673 3713 2687 3727
rect 2793 3713 2807 3727
rect 2834 3713 2848 3727
rect 2933 3713 2947 3727
rect 3032 3713 3046 3727
rect 3074 3713 3088 3727
rect 3133 3713 3147 3727
rect 3313 3713 3327 3727
rect 3353 3713 3367 3727
rect 3553 3713 3567 3727
rect 3593 3713 3607 3727
rect 3693 3713 3707 3727
rect 3733 3713 3747 3727
rect 2313 3693 2327 3707
rect 2353 3693 2367 3707
rect 2773 3693 2787 3707
rect 2813 3693 2827 3707
rect 3013 3693 3027 3707
rect 3052 3693 3066 3707
rect 3094 3693 3108 3707
rect 2113 3673 2127 3687
rect 2333 3673 2347 3687
rect 2533 3673 2547 3687
rect 1093 3653 1107 3667
rect 1753 3653 1767 3667
rect 1993 3653 2007 3667
rect 3853 3733 3867 3747
rect 3913 3733 3927 3747
rect 5113 3733 5127 3747
rect 5153 3733 5167 3747
rect 3832 3713 3846 3727
rect 3874 3713 3888 3727
rect 4013 3713 4027 3727
rect 4133 3713 4147 3727
rect 4173 3713 4187 3727
rect 4593 3713 4607 3727
rect 4993 3713 5007 3727
rect 5033 3713 5047 3727
rect 5133 3713 5147 3727
rect 5253 3713 5267 3727
rect 5613 3713 5627 3727
rect 3172 3693 3186 3707
rect 3213 3693 3227 3707
rect 3293 3693 3307 3707
rect 3333 3693 3347 3707
rect 3453 3693 3467 3707
rect 3493 3693 3507 3707
rect 3793 3693 3807 3707
rect 3973 3693 3987 3707
rect 4033 3693 4047 3707
rect 4113 3693 4127 3707
rect 4153 3693 4167 3707
rect 4233 3693 4247 3707
rect 4313 3693 4327 3707
rect 4353 3693 4367 3707
rect 4473 3693 4487 3707
rect 4553 3693 4567 3707
rect 4713 3693 4727 3707
rect 4792 3693 4806 3707
rect 4833 3693 4847 3707
rect 4972 3693 4986 3707
rect 5013 3693 5027 3707
rect 5313 3693 5327 3707
rect 5392 3693 5406 3707
rect 5433 3693 5447 3707
rect 3193 3673 3207 3687
rect 3473 3673 3487 3687
rect 5233 3673 5247 3687
rect 5573 3673 5587 3687
rect 793 3633 807 3647
rect 3133 3633 3147 3647
rect 3293 3573 3307 3587
rect 3673 3573 3687 3587
rect 433 3553 447 3567
rect 2293 3553 2307 3567
rect 72 3513 86 3527
rect 112 3513 126 3527
rect 93 3493 107 3507
rect 134 3493 148 3507
rect 193 3493 207 3507
rect 233 3493 247 3507
rect 333 3493 347 3507
rect 373 3493 387 3507
rect 214 3473 228 3487
rect 273 3473 287 3487
rect 352 3473 366 3487
rect 1073 3533 1087 3547
rect 1992 3533 2006 3547
rect 2233 3533 2247 3547
rect 493 3513 507 3527
rect 553 3513 567 3527
rect 613 3513 627 3527
rect 654 3513 668 3527
rect 913 3513 927 3527
rect 473 3493 487 3507
rect 513 3493 527 3507
rect 633 3493 647 3507
rect 673 3493 687 3507
rect 753 3493 767 3507
rect 793 3493 807 3507
rect 893 3493 907 3507
rect 933 3493 947 3507
rect 773 3473 787 3487
rect 833 3473 847 3487
rect 1133 3513 1147 3527
rect 1173 3513 1187 3527
rect 1213 3513 1227 3527
rect 1552 3513 1566 3527
rect 1633 3513 1647 3527
rect 1693 3513 1707 3527
rect 1733 3513 1747 3527
rect 1793 3513 1807 3527
rect 1973 3513 1987 3527
rect 2013 3513 2027 3527
rect 2133 3513 2147 3527
rect 2173 3513 2187 3527
rect 1033 3493 1047 3507
rect 1153 3493 1167 3507
rect 1193 3493 1207 3507
rect 1293 3493 1307 3507
rect 1333 3493 1347 3507
rect 1473 3493 1487 3507
rect 1713 3493 1727 3507
rect 1753 3493 1767 3507
rect 1893 3493 1907 3507
rect 2113 3493 2127 3507
rect 2153 3493 2167 3507
rect 1313 3473 1327 3487
rect 1373 3473 1387 3487
rect 1454 3473 1468 3487
rect 1493 3473 1507 3487
rect 1533 3473 1547 3487
rect 1593 3473 1607 3487
rect 1873 3473 1887 3487
rect 1913 3473 1927 3487
rect 993 3433 1007 3447
rect 1534 3433 1548 3447
rect 2593 3533 2607 3547
rect 2713 3533 2727 3547
rect 2953 3533 2967 3547
rect 3153 3533 3167 3547
rect 2473 3513 2487 3527
rect 2533 3513 2547 3527
rect 2692 3513 2706 3527
rect 2733 3513 2747 3527
rect 2773 3513 2787 3527
rect 2813 3513 2827 3527
rect 2853 3513 2867 3527
rect 2353 3493 2367 3507
rect 2453 3493 2467 3507
rect 2493 3493 2507 3507
rect 2633 3493 2647 3507
rect 2333 3473 2347 3487
rect 2373 3473 2387 3487
rect 2833 3493 2847 3507
rect 2873 3493 2887 3507
rect 2993 3493 3007 3507
rect 3054 3493 3068 3507
rect 3093 3493 3107 3507
rect 3073 3473 3087 3487
rect 3212 3513 3226 3527
rect 3273 3513 3287 3527
rect 3333 3533 3347 3547
rect 3453 3513 3467 3527
rect 3513 3513 3527 3527
rect 3193 3493 3207 3507
rect 3233 3493 3247 3507
rect 3293 3493 3307 3507
rect 3433 3493 3447 3507
rect 3473 3493 3487 3507
rect 3572 3493 3586 3507
rect 3613 3493 3627 3507
rect 3393 3473 3407 3487
rect 3593 3473 3607 3487
rect 5373 3533 5387 3547
rect 3713 3513 3727 3527
rect 3753 3513 3767 3527
rect 4333 3513 4347 3527
rect 4373 3513 4387 3527
rect 4433 3513 4447 3527
rect 4573 3513 4587 3527
rect 4633 3513 4647 3527
rect 4833 3513 4847 3527
rect 4913 3513 4927 3527
rect 4953 3513 4967 3527
rect 5113 3513 5127 3527
rect 3732 3493 3746 3507
rect 3773 3493 3787 3507
rect 3853 3493 3867 3507
rect 4012 3493 4026 3507
rect 4133 3493 4147 3507
rect 4253 3493 4267 3507
rect 4353 3493 4367 3507
rect 4393 3493 4407 3507
rect 4493 3493 4507 3507
rect 4613 3493 4627 3507
rect 4653 3493 4667 3507
rect 4753 3493 4767 3507
rect 5093 3493 5107 3507
rect 5133 3493 5147 3507
rect 4473 3473 4487 3487
rect 4513 3473 4527 3487
rect 4733 3473 4747 3487
rect 4773 3473 4787 3487
rect 2773 3433 2787 3447
rect 4433 3433 4447 3447
rect 2212 3413 2226 3427
rect 2293 3413 2307 3427
rect 5232 3513 5246 3527
rect 5273 3513 5287 3527
rect 5473 3513 5487 3527
rect 5513 3513 5527 3527
rect 5253 3493 5267 3507
rect 5293 3493 5307 3507
rect 5413 3493 5427 3507
rect 5493 3493 5507 3507
rect 5633 3493 5647 3507
rect 5693 3493 5707 3507
rect 5613 3473 5627 3487
rect 5653 3473 5667 3487
rect 5533 3453 5547 3467
rect 5293 3433 5307 3447
rect 5193 3393 5207 3407
rect 5693 3393 5707 3407
rect 2093 3333 2107 3347
rect 2773 3333 2787 3347
rect 5693 3333 5707 3347
rect 453 3313 467 3327
rect 1233 3313 1247 3327
rect 354 3253 368 3267
rect 413 3253 427 3267
rect 713 3273 727 3287
rect 533 3253 547 3267
rect 73 3233 87 3247
rect 113 3233 127 3247
rect 214 3233 228 3247
rect 254 3233 268 3247
rect 333 3233 347 3247
rect 373 3233 387 3247
rect 513 3233 527 3247
rect 552 3233 566 3247
rect 612 3233 626 3247
rect 653 3233 667 3247
rect 93 3213 107 3227
rect 134 3213 148 3227
rect 193 3213 207 3227
rect 233 3213 247 3227
rect 634 3213 648 3227
rect 1154 3253 1168 3267
rect 1633 3253 1647 3267
rect 1693 3253 1707 3267
rect 1913 3253 1927 3267
rect 1973 3253 1987 3267
rect 2013 3253 2027 3267
rect 2053 3253 2067 3267
rect 753 3233 767 3247
rect 833 3233 847 3247
rect 893 3233 907 3247
rect 1013 3233 1027 3247
rect 1053 3233 1067 3247
rect 1133 3233 1147 3247
rect 1173 3233 1187 3247
rect 1293 3233 1307 3247
rect 1333 3233 1347 3247
rect 1413 3233 1427 3247
rect 1673 3233 1687 3247
rect 1713 3233 1727 3247
rect 1773 3233 1787 3247
rect 1913 3233 1927 3247
rect 873 3213 887 3227
rect 933 3213 947 3227
rect 993 3213 1007 3227
rect 1032 3213 1046 3227
rect 1313 3213 1327 3227
rect 1353 3213 1367 3227
rect 1513 3213 1527 3227
rect 1594 3213 1608 3227
rect 1873 3213 1887 3227
rect 2273 3273 2287 3287
rect 2633 3273 2647 3287
rect 2153 3253 2167 3267
rect 2193 3253 2207 3267
rect 2272 3253 2286 3267
rect 2314 3253 2328 3267
rect 2393 3253 2407 3267
rect 2453 3253 2467 3267
rect 2033 3233 2047 3247
rect 2113 3233 2127 3247
rect 2173 3233 2187 3247
rect 2292 3233 2306 3247
rect 2373 3233 2387 3247
rect 2413 3233 2427 3247
rect 2513 3233 2527 3247
rect 2553 3233 2567 3247
rect 2673 3233 2687 3247
rect 2713 3233 2727 3247
rect 2533 3213 2547 3227
rect 793 3193 807 3207
rect 1253 3193 1267 3207
rect 1453 3193 1467 3207
rect 1813 3193 1827 3207
rect 2633 3213 2647 3227
rect 2693 3213 2707 3227
rect 2733 3213 2747 3227
rect 4654 3293 4668 3307
rect 4913 3273 4927 3287
rect 5073 3273 5087 3287
rect 3213 3253 3227 3267
rect 4113 3253 4127 3267
rect 4153 3253 4167 3267
rect 4573 3253 4587 3267
rect 4613 3253 4627 3267
rect 4653 3253 4667 3267
rect 4693 3253 4707 3267
rect 4733 3253 4747 3267
rect 2913 3233 2927 3247
rect 3013 3233 3027 3247
rect 3053 3233 3067 3247
rect 3293 3233 3307 3247
rect 3433 3233 3447 3247
rect 3493 3233 3507 3247
rect 3533 3233 3547 3247
rect 3714 3233 3728 3247
rect 3953 3233 3967 3247
rect 4133 3233 4147 3247
rect 4232 3233 4246 3247
rect 4273 3233 4287 3247
rect 4373 3233 4387 3247
rect 4473 3233 4487 3247
rect 4593 3233 4607 3247
rect 4713 3233 4727 3247
rect 4813 3233 4827 3247
rect 4853 3233 4867 3247
rect 4973 3233 4987 3247
rect 5013 3233 5027 3247
rect 5333 3233 5347 3247
rect 5373 3233 5387 3247
rect 5473 3233 5487 3247
rect 5513 3233 5527 3247
rect 2813 3213 2827 3227
rect 2853 3213 2867 3227
rect 3033 3213 3047 3227
rect 3093 3213 3107 3227
rect 3173 3212 3187 3226
rect 3453 3213 3467 3227
rect 3513 3213 3527 3227
rect 3593 3213 3607 3227
rect 3673 3213 3687 3227
rect 3833 3213 3847 3227
rect 3913 3213 3927 3227
rect 4253 3213 4267 3227
rect 4293 3213 4307 3227
rect 4793 3213 4807 3227
rect 4833 3213 4847 3227
rect 4873 3213 4887 3227
rect 4913 3213 4927 3227
rect 4993 3213 5007 3227
rect 5033 3213 5047 3227
rect 5213 3213 5227 3227
rect 5253 3213 5267 3227
rect 5313 3213 5327 3227
rect 5353 3213 5367 3227
rect 5493 3213 5507 3227
rect 5573 3213 5587 3227
rect 5614 3213 5628 3227
rect 2833 3193 2847 3207
rect 2953 3193 2967 3207
rect 3233 3193 3247 3207
rect 3413 3193 3427 3207
rect 4353 3193 4367 3207
rect 4493 3193 4507 3207
rect 5133 3193 5147 3207
rect 5233 3193 5247 3207
rect 5633 3193 5647 3207
rect 2773 3173 2787 3187
rect 1253 3153 1267 3167
rect 2613 3153 2627 3167
rect 273 3093 287 3107
rect 1733 3093 1747 3107
rect 2273 3093 2287 3107
rect 2412 3093 2426 3107
rect 2434 3093 2448 3107
rect 3833 3093 3847 3107
rect 133 3033 147 3047
rect 93 3013 107 3027
rect 213 3013 227 3027
rect 293 3053 307 3067
rect 733 3053 747 3067
rect 1012 3053 1026 3067
rect 193 2993 207 3007
rect 233 2993 247 3007
rect 272 2993 286 3007
rect 453 3033 467 3047
rect 512 3033 526 3047
rect 872 3033 886 3047
rect 913 3033 927 3047
rect 993 3033 1007 3047
rect 1033 3033 1047 3047
rect 1433 3033 1447 3047
rect 1473 3033 1487 3047
rect 1513 3033 1527 3047
rect 1553 3033 1567 3047
rect 353 3013 367 3027
rect 393 3013 407 3027
rect 493 3013 507 3027
rect 533 3013 547 3027
rect 633 3013 647 3027
rect 673 3013 687 3027
rect 733 3013 747 3027
rect 852 3013 866 3027
rect 893 3013 907 3027
rect 1113 3013 1127 3027
rect 1253 3013 1267 3027
rect 1293 3013 1307 3027
rect 1373 3013 1387 3027
rect 313 2993 327 3007
rect 373 2993 387 3007
rect 653 2993 667 3007
rect 1093 2993 1107 3007
rect 1133 2993 1147 3007
rect 1273 2993 1287 3007
rect 1353 2993 1367 3007
rect 1393 2993 1407 3007
rect 1492 3013 1506 3027
rect 1533 3013 1547 3027
rect 1693 3033 1707 3047
rect 2014 3073 2028 3087
rect 1893 3033 1907 3047
rect 1933 3033 1947 3047
rect 1993 3033 2007 3047
rect 1793 3013 1807 3027
rect 1833 3013 1847 3027
rect 1913 3013 1927 3027
rect 1953 3013 1967 3027
rect 1813 2993 1827 3007
rect 1993 2993 2007 3007
rect 2074 3033 2088 3047
rect 2114 3033 2128 3047
rect 2173 3033 2187 3047
rect 2413 3053 2427 3067
rect 2313 3033 2327 3047
rect 2374 3033 2388 3047
rect 2052 3013 2066 3027
rect 2093 3013 2107 3027
rect 2213 3013 2227 3027
rect 2353 3013 2367 3027
rect 2813 3073 2827 3087
rect 2973 3073 2987 3087
rect 2553 3053 2567 3067
rect 2493 3013 2507 3027
rect 2612 3033 2626 3047
rect 2653 3033 2667 3047
rect 2713 3033 2727 3047
rect 2753 3033 2767 3047
rect 2853 3033 2867 3047
rect 2893 3033 2907 3047
rect 2593 3013 2607 3027
rect 2633 3013 2647 3027
rect 2733 3013 2747 3027
rect 2773 3013 2787 3027
rect 2813 3013 2827 3027
rect 2873 3013 2887 3027
rect 2913 3013 2927 3027
rect 2473 2993 2487 3007
rect 2513 2993 2527 3007
rect 2553 2993 2567 3007
rect 2913 2993 2927 3007
rect 573 2953 587 2967
rect 1193 2953 1207 2967
rect 1433 2953 1447 2967
rect 1613 2953 1627 2967
rect 1953 2953 1967 2967
rect 2013 2953 2027 2967
rect 2433 2953 2447 2967
rect 293 2933 307 2947
rect 3033 3053 3047 3067
rect 3093 3033 3107 3047
rect 3133 3033 3147 3047
rect 3233 3033 3247 3047
rect 3272 3033 3286 3047
rect 3373 3033 3387 3047
rect 3413 3033 3427 3047
rect 3533 3033 3547 3047
rect 3574 3033 3588 3047
rect 3753 3033 3767 3047
rect 3873 3053 3887 3067
rect 4013 3053 4027 3067
rect 4093 3053 4107 3067
rect 4232 3053 4246 3067
rect 5553 3053 5567 3067
rect 3993 3033 4007 3047
rect 4033 3033 4047 3047
rect 4213 3033 4227 3047
rect 4253 3033 4267 3047
rect 4313 3033 4327 3047
rect 4353 3033 4367 3047
rect 4573 3033 4587 3047
rect 4613 3033 4627 3047
rect 4653 3033 4667 3047
rect 4733 3033 4747 3047
rect 4773 3033 4787 3047
rect 5233 3033 5247 3047
rect 5312 3033 5326 3047
rect 5354 3033 5368 3047
rect 5393 3033 5407 3047
rect 5453 3033 5467 3047
rect 5493 3033 5507 3047
rect 5573 3033 5587 3047
rect 3033 3013 3047 3027
rect 3113 3013 3127 3027
rect 3154 3013 3168 3027
rect 3193 3013 3207 3027
rect 3253 3013 3267 3027
rect 3293 3013 3307 3027
rect 3393 3013 3407 3027
rect 3433 3013 3447 3027
rect 3653 3013 3667 3027
rect 3693 3013 3707 3027
rect 3913 3013 3927 3027
rect 4133 3013 4147 3027
rect 4334 3013 4348 3027
rect 4373 3013 4387 3027
rect 4493 3013 4507 3027
rect 4593 3013 4607 3027
rect 4633 3013 4647 3027
rect 4752 3013 4766 3027
rect 4793 3013 4807 3027
rect 4894 3013 4908 3027
rect 4952 3013 4966 3027
rect 4993 3013 5007 3027
rect 5033 3013 5047 3027
rect 5133 3013 5147 3027
rect 5173 3013 5187 3027
rect 4053 2993 4067 3007
rect 3592 2973 3606 2987
rect 3193 2933 3207 2947
rect 4473 2993 4487 3007
rect 4514 2993 4528 3007
rect 4833 2993 4847 3007
rect 4874 2993 4888 3007
rect 4913 2993 4927 3007
rect 4274 2973 4288 2987
rect 4373 2973 4387 2987
rect 4052 2933 4066 2947
rect 5013 2993 5027 3007
rect 5093 2993 5107 3007
rect 5153 2993 5167 3007
rect 5293 3013 5307 3027
rect 5332 3013 5346 3027
rect 4953 2953 4967 2967
rect 4833 2933 4847 2947
rect 5433 3013 5447 3027
rect 5473 3013 5487 3027
rect 5613 3013 5627 3027
rect 33 2913 47 2927
rect 2973 2913 2987 2927
rect 3593 2913 3607 2927
rect 4272 2913 4286 2927
rect 5393 2913 5407 2927
rect 1613 2853 1627 2867
rect 1873 2853 1887 2867
rect 3773 2853 3787 2867
rect 5233 2853 5247 2867
rect 1233 2813 1247 2827
rect 13 2793 27 2807
rect 173 2773 187 2787
rect 213 2773 227 2787
rect 253 2773 267 2787
rect 373 2773 387 2787
rect 974 2773 988 2787
rect 1013 2773 1027 2787
rect 1053 2773 1067 2787
rect 1113 2773 1127 2787
rect 1153 2773 1167 2787
rect 1233 2773 1247 2787
rect 1273 2773 1287 2787
rect 1393 2773 1407 2787
rect 72 2753 86 2767
rect 114 2753 128 2767
rect 233 2753 247 2767
rect 273 2753 287 2767
rect 373 2753 387 2767
rect 414 2753 428 2767
rect 493 2753 507 2767
rect 533 2753 547 2767
rect 653 2753 667 2767
rect 733 2753 747 2767
rect 773 2753 787 2767
rect 873 2753 887 2767
rect 913 2753 927 2767
rect 13 2733 27 2747
rect 92 2733 106 2747
rect 133 2733 147 2747
rect 174 2733 188 2747
rect 333 2733 347 2747
rect 393 2733 407 2747
rect 513 2733 527 2747
rect 553 2733 567 2747
rect 753 2733 767 2747
rect 793 2733 807 2747
rect 853 2733 867 2747
rect 894 2733 908 2747
rect 1032 2753 1046 2767
rect 1133 2753 1147 2767
rect 1254 2753 1268 2767
rect 1513 2753 1527 2767
rect 1553 2753 1567 2767
rect 1433 2733 1447 2747
rect 1492 2733 1506 2747
rect 1533 2733 1547 2747
rect 1573 2733 1587 2747
rect 2114 2813 2128 2827
rect 3373 2793 3387 2807
rect 3553 2793 3567 2807
rect 1913 2773 1927 2787
rect 1953 2773 1967 2787
rect 2113 2773 2127 2787
rect 2153 2773 2167 2787
rect 2194 2773 2208 2787
rect 2253 2773 2267 2787
rect 2412 2773 2426 2787
rect 2453 2773 2467 2787
rect 2533 2773 2547 2787
rect 1873 2753 1887 2767
rect 1933 2753 1947 2767
rect 1993 2753 2007 2767
rect 2033 2753 2047 2767
rect 2073 2753 2087 2767
rect 2173 2753 2187 2767
rect 1653 2733 1667 2747
rect 1693 2733 1707 2747
rect 1773 2733 1787 2747
rect 1813 2733 1827 2747
rect 653 2713 667 2727
rect 973 2713 987 2727
rect 1333 2713 1347 2727
rect 1613 2713 1627 2727
rect 2053 2733 2067 2747
rect 2093 2733 2107 2747
rect 2313 2753 2327 2767
rect 2433 2753 2447 2767
rect 2533 2753 2547 2767
rect 2573 2753 2587 2767
rect 2813 2753 2827 2767
rect 2853 2753 2867 2767
rect 2953 2753 2967 2767
rect 2993 2753 3007 2767
rect 3093 2753 3107 2767
rect 2353 2733 2367 2747
rect 2552 2733 2566 2747
rect 1993 2693 2007 2707
rect 2633 2693 2647 2707
rect 2733 2733 2747 2747
rect 2793 2733 2807 2747
rect 2833 2733 2847 2747
rect 2933 2733 2947 2747
rect 2973 2733 2987 2747
rect 3233 2733 3247 2747
rect 3273 2733 3287 2747
rect 3533 2773 3547 2787
rect 3593 2773 3607 2787
rect 3433 2753 3447 2767
rect 3473 2753 3487 2767
rect 3572 2753 3586 2767
rect 3453 2733 3467 2747
rect 3693 2733 3707 2747
rect 3733 2733 3747 2747
rect 3113 2713 3127 2727
rect 3153 2713 3167 2727
rect 3713 2713 3727 2727
rect 4713 2833 4727 2847
rect 4533 2813 4547 2827
rect 3933 2793 3947 2807
rect 3933 2773 3947 2787
rect 3973 2773 3987 2787
rect 4493 2773 4507 2787
rect 4533 2773 4547 2787
rect 3953 2753 3967 2767
rect 4053 2753 4067 2767
rect 4093 2753 4107 2767
rect 4213 2753 4227 2767
rect 4253 2753 4267 2767
rect 4353 2753 4367 2767
rect 4393 2753 4407 2767
rect 4513 2753 4527 2767
rect 4612 2753 4626 2767
rect 4653 2753 4667 2767
rect 4693 2753 4707 2767
rect 3793 2733 3807 2747
rect 3853 2733 3867 2747
rect 4032 2733 4046 2747
rect 4073 2733 4087 2747
rect 4193 2733 4207 2747
rect 4233 2733 4247 2747
rect 4273 2733 4287 2747
rect 4333 2733 4347 2747
rect 4373 2733 4387 2747
rect 4592 2733 4606 2747
rect 4634 2733 4648 2747
rect 4693 2713 4707 2727
rect 4993 2813 5007 2827
rect 4753 2753 4767 2767
rect 4793 2753 4807 2767
rect 4873 2753 4887 2767
rect 4933 2753 4947 2767
rect 4773 2733 4787 2747
rect 4813 2733 4827 2747
rect 4894 2733 4908 2747
rect 4953 2733 4967 2747
rect 5032 2773 5046 2787
rect 5073 2773 5087 2787
rect 5054 2753 5068 2767
rect 5194 2753 5208 2767
rect 5153 2733 5167 2747
rect 5433 2833 5447 2847
rect 5693 2833 5707 2847
rect 5333 2813 5347 2827
rect 5293 2773 5307 2787
rect 5273 2733 5287 2747
rect 3773 2693 3787 2707
rect 4713 2693 4727 2707
rect 4993 2693 5007 2707
rect 5233 2693 5247 2707
rect 5553 2813 5567 2827
rect 5373 2773 5387 2787
rect 5473 2773 5487 2787
rect 5513 2773 5527 2787
rect 5393 2753 5407 2767
rect 5492 2753 5506 2767
rect 5693 2793 5707 2807
rect 5633 2753 5647 2767
rect 5553 2733 5567 2747
rect 5593 2733 5607 2747
rect 2653 2673 2667 2687
rect 5332 2673 5346 2687
rect 5693 2673 5707 2687
rect 333 2613 347 2627
rect 1213 2613 1227 2627
rect 2373 2613 2387 2627
rect 2833 2613 2847 2627
rect 3373 2613 3387 2627
rect 4074 2613 4088 2627
rect 5693 2613 5707 2627
rect 312 2573 326 2587
rect 214 2553 228 2567
rect 273 2553 287 2567
rect 93 2533 107 2547
rect 133 2533 147 2547
rect 192 2533 206 2547
rect 234 2533 248 2547
rect 53 2513 67 2527
rect 113 2513 127 2527
rect 873 2593 887 2607
rect 753 2573 767 2587
rect 813 2573 827 2587
rect 334 2553 348 2567
rect 493 2553 507 2567
rect 533 2553 547 2567
rect 573 2553 587 2567
rect 613 2553 627 2567
rect 693 2553 707 2567
rect 373 2533 387 2547
rect 413 2533 427 2547
rect 513 2533 527 2547
rect 553 2533 567 2547
rect 673 2533 687 2547
rect 713 2533 727 2547
rect 1153 2573 1167 2587
rect 1133 2553 1147 2567
rect 1174 2553 1188 2567
rect 333 2513 347 2527
rect 393 2513 407 2527
rect 313 2493 327 2507
rect 853 2533 867 2547
rect 913 2533 927 2547
rect 1033 2533 1047 2547
rect 1073 2533 1087 2547
rect 873 2513 887 2527
rect 933 2513 947 2527
rect 1053 2513 1067 2527
rect 1413 2573 1427 2587
rect 1513 2573 1527 2587
rect 1913 2573 1927 2587
rect 1733 2553 1747 2567
rect 1774 2553 1788 2567
rect 1813 2553 1827 2567
rect 2113 2553 2127 2567
rect 2152 2553 2166 2567
rect 2253 2553 2267 2567
rect 2333 2553 2347 2567
rect 2753 2573 2767 2587
rect 2453 2553 2467 2567
rect 2513 2553 2527 2567
rect 2573 2553 2587 2567
rect 1293 2533 1307 2547
rect 1413 2533 1427 2547
rect 1493 2533 1507 2547
rect 1613 2533 1627 2547
rect 1653 2533 1667 2547
rect 1753 2533 1767 2547
rect 1793 2533 1807 2547
rect 1273 2513 1287 2527
rect 1313 2513 1327 2527
rect 1553 2513 1567 2527
rect 1633 2513 1647 2527
rect 2013 2533 2027 2547
rect 2053 2533 2067 2547
rect 2133 2533 2147 2547
rect 2174 2533 2188 2547
rect 2293 2533 2307 2547
rect 2553 2533 2567 2547
rect 1853 2453 1867 2467
rect 2033 2513 2047 2527
rect 2713 2553 2727 2567
rect 2813 2533 2827 2547
rect 2633 2493 2647 2507
rect 2873 2553 2887 2567
rect 2912 2553 2926 2567
rect 2953 2553 2967 2567
rect 3013 2553 3027 2567
rect 3093 2553 3107 2567
rect 3133 2553 3147 2567
rect 2892 2533 2906 2547
rect 2934 2533 2948 2547
rect 3314 2553 3328 2567
rect 3513 2593 3527 2607
rect 3433 2553 3447 2567
rect 3533 2573 3547 2587
rect 3593 2553 3607 2567
rect 3633 2553 3647 2567
rect 3673 2553 3687 2567
rect 3733 2553 3747 2567
rect 3293 2533 3307 2547
rect 3333 2533 3347 2547
rect 3373 2533 3387 2547
rect 3412 2533 3426 2547
rect 3453 2533 3467 2547
rect 3533 2533 3547 2547
rect 3573 2533 3587 2547
rect 3613 2533 3627 2547
rect 3233 2493 3247 2507
rect 3713 2533 3727 2547
rect 3753 2533 3767 2547
rect 3673 2513 3687 2527
rect 3853 2553 3867 2567
rect 3913 2553 3927 2567
rect 3873 2533 3887 2547
rect 3933 2533 3947 2547
rect 4013 2533 4027 2547
rect 5513 2593 5527 2607
rect 5633 2593 5647 2607
rect 4793 2573 4807 2587
rect 4933 2573 4947 2587
rect 4112 2553 4126 2567
rect 4154 2553 4168 2567
rect 4212 2553 4226 2567
rect 4253 2553 4267 2567
rect 4293 2553 4307 2567
rect 4333 2553 4347 2567
rect 4393 2553 4407 2567
rect 4533 2553 4547 2567
rect 4133 2533 4147 2547
rect 4173 2533 4187 2547
rect 3993 2513 4007 2527
rect 4033 2513 4047 2527
rect 4073 2513 4087 2527
rect 2833 2453 2847 2467
rect 3373 2453 3387 2467
rect 3813 2453 3827 2467
rect 4273 2533 4287 2547
rect 4314 2533 4328 2547
rect 4453 2533 4467 2547
rect 4493 2533 4507 2547
rect 4473 2513 4487 2527
rect 5013 2553 5027 2567
rect 5073 2553 5087 2567
rect 5293 2553 5307 2567
rect 5333 2553 5347 2567
rect 5393 2553 5407 2567
rect 5433 2553 5447 2567
rect 5473 2553 5487 2567
rect 4713 2533 4727 2547
rect 4793 2533 4807 2547
rect 4873 2533 4887 2547
rect 4913 2533 4927 2547
rect 5153 2533 5167 2547
rect 5273 2533 5287 2547
rect 5313 2533 5327 2547
rect 5413 2533 5427 2547
rect 5453 2533 5467 2547
rect 4673 2513 4687 2527
rect 4733 2513 4747 2527
rect 5132 2513 5146 2527
rect 5173 2513 5187 2527
rect 5573 2533 5587 2547
rect 5553 2513 5567 2527
rect 5593 2513 5607 2527
rect 5633 2513 5647 2527
rect 4873 2453 4887 2467
rect 5513 2453 5527 2467
rect 5693 2453 5707 2467
rect 753 2433 767 2447
rect 973 2433 987 2447
rect 1213 2433 1227 2447
rect 1953 2433 1967 2447
rect 4213 2433 4227 2447
rect 4633 2433 4647 2447
rect 1813 2373 1827 2387
rect 2673 2373 2687 2387
rect 3313 2373 3327 2387
rect 3813 2373 3827 2387
rect 4053 2373 4067 2387
rect 4613 2373 4627 2387
rect 5633 2373 5647 2387
rect 1653 2333 1667 2347
rect 72 2293 86 2307
rect 113 2293 127 2307
rect 93 2273 107 2287
rect 133 2273 147 2287
rect 213 2273 227 2287
rect 253 2273 267 2287
rect 352 2273 366 2287
rect 394 2273 408 2287
rect 233 2253 247 2267
rect 273 2253 287 2267
rect 333 2253 347 2267
rect 372 2253 386 2267
rect 533 2293 547 2307
rect 773 2293 787 2307
rect 813 2293 827 2307
rect 1033 2293 1047 2307
rect 1093 2293 1107 2307
rect 513 2273 527 2287
rect 553 2273 567 2287
rect 632 2273 646 2287
rect 672 2273 686 2287
rect 753 2273 767 2287
rect 793 2273 807 2287
rect 914 2273 928 2287
rect 953 2273 967 2287
rect 1073 2273 1087 2287
rect 1113 2273 1127 2287
rect 653 2253 667 2267
rect 694 2253 708 2267
rect 893 2253 907 2267
rect 933 2253 947 2267
rect 1233 2293 1247 2307
rect 1313 2293 1327 2307
rect 1353 2293 1367 2307
rect 1213 2273 1227 2287
rect 1253 2273 1267 2287
rect 1333 2273 1347 2287
rect 1453 2273 1467 2287
rect 1493 2273 1507 2287
rect 1713 2273 1727 2287
rect 1753 2273 1767 2287
rect 1473 2253 1487 2267
rect 1513 2253 1527 2267
rect 1573 2253 1587 2267
rect 1613 2253 1627 2267
rect 1653 2253 1667 2267
rect 1733 2253 1747 2267
rect 1773 2253 1787 2267
rect 2553 2353 2567 2367
rect 2393 2313 2407 2327
rect 2133 2293 2147 2307
rect 2173 2293 2187 2307
rect 2433 2293 2447 2307
rect 1853 2273 1867 2287
rect 1893 2273 1907 2287
rect 1993 2273 2007 2287
rect 2033 2273 2047 2287
rect 2153 2273 2167 2287
rect 2273 2273 2287 2287
rect 2413 2273 2427 2287
rect 2493 2273 2507 2287
rect 1874 2253 1888 2267
rect 1914 2253 1928 2267
rect 1973 2253 1987 2267
rect 2013 2253 2027 2267
rect 1153 2233 1167 2247
rect 1593 2233 1607 2247
rect 1813 2233 1827 2247
rect 2314 2253 2328 2267
rect 2513 2253 2527 2267
rect 2913 2333 2927 2347
rect 3313 2333 3327 2347
rect 3433 2333 3447 2347
rect 2593 2293 2607 2307
rect 2673 2293 2687 2307
rect 2613 2273 2627 2287
rect 2833 2273 2847 2287
rect 3093 2273 3107 2287
rect 3133 2273 3147 2287
rect 2713 2253 2727 2267
rect 2773 2253 2787 2267
rect 2913 2253 2927 2267
rect 2953 2253 2967 2267
rect 2993 2253 3007 2267
rect 3072 2253 3086 2267
rect 3113 2253 3127 2267
rect 3153 2253 3167 2267
rect 2973 2233 2987 2247
rect 2553 2213 2567 2227
rect 2873 2213 2887 2227
rect 3273 2253 3287 2267
rect 3394 2253 3408 2267
rect 3653 2313 3667 2327
rect 3493 2273 3507 2287
rect 3533 2273 3547 2287
rect 3712 2273 3726 2287
rect 3753 2273 3767 2287
rect 3853 2293 3867 2307
rect 3893 2293 3907 2307
rect 3874 2273 3888 2287
rect 3973 2273 3987 2287
rect 4013 2273 4027 2287
rect 3253 2233 3267 2247
rect 3373 2233 3387 2247
rect 3514 2253 3528 2267
rect 3693 2253 3707 2267
rect 3733 2253 3747 2267
rect 3813 2253 3827 2267
rect 3953 2253 3967 2267
rect 3993 2253 4007 2267
rect 3633 2233 3647 2247
rect 3433 2213 3447 2227
rect 4333 2353 4347 2367
rect 4113 2273 4127 2287
rect 4153 2273 4167 2287
rect 4073 2253 4087 2267
rect 4133 2253 4147 2267
rect 4173 2253 4187 2267
rect 4232 2253 4246 2267
rect 4274 2253 4288 2267
rect 4252 2233 4266 2247
rect 5353 2333 5367 2347
rect 4613 2313 4627 2327
rect 4753 2313 4767 2327
rect 5173 2313 5187 2327
rect 4373 2293 4387 2307
rect 4413 2293 4427 2307
rect 4393 2273 4407 2287
rect 4513 2273 4527 2287
rect 4553 2273 4567 2287
rect 4653 2273 4667 2287
rect 4694 2273 4708 2287
rect 4813 2293 4827 2307
rect 4853 2293 4867 2307
rect 4773 2273 4787 2287
rect 4834 2273 4848 2287
rect 4953 2273 4967 2287
rect 5073 2273 5087 2287
rect 5113 2273 5127 2287
rect 4492 2253 4506 2267
rect 4533 2253 4547 2267
rect 4573 2253 4587 2267
rect 4633 2253 4647 2267
rect 4673 2253 4687 2267
rect 4713 2253 4727 2267
rect 4753 2253 4767 2267
rect 4333 2213 4347 2227
rect 5233 2273 5247 2287
rect 5272 2273 5286 2287
rect 4913 2253 4927 2267
rect 4993 2253 5007 2267
rect 5052 2253 5066 2267
rect 5093 2253 5107 2267
rect 5133 2253 5147 2267
rect 5173 2253 5187 2267
rect 5213 2253 5227 2267
rect 5253 2253 5267 2267
rect 5293 2253 5307 2267
rect 5633 2313 5647 2327
rect 5393 2273 5407 2287
rect 5433 2273 5447 2287
rect 5533 2273 5547 2287
rect 5573 2273 5587 2287
rect 5413 2253 5427 2267
rect 5453 2253 5467 2267
rect 5512 2253 5526 2267
rect 5554 2253 5568 2267
rect 453 2193 467 2207
rect 2213 2193 2227 2207
rect 3193 2193 3207 2207
rect 4052 2193 4066 2207
rect 4074 2193 4088 2207
rect 4773 2193 4787 2207
rect 5353 2193 5367 2207
rect 5613 2193 5627 2207
rect 453 2133 467 2147
rect 3313 2133 3327 2147
rect 3593 2133 3607 2147
rect 4273 2133 4287 2147
rect 4673 2133 4687 2147
rect 5613 2133 5627 2147
rect 73 2073 87 2087
rect 114 2073 128 2087
rect 333 2073 347 2087
rect 393 2073 407 2087
rect 93 2053 107 2067
rect 133 2053 147 2067
rect 194 2053 208 2067
rect 233 2053 247 2067
rect 372 2053 386 2067
rect 413 2053 427 2067
rect 213 2033 227 2047
rect 273 2033 287 2047
rect 2933 2113 2947 2127
rect 1433 2093 1447 2107
rect 2753 2093 2767 2107
rect 513 2073 527 2087
rect 553 2073 567 2087
rect 493 2053 507 2067
rect 533 2053 547 2067
rect 693 2073 707 2087
rect 1513 2073 1527 2087
rect 1553 2073 1567 2087
rect 1593 2073 1607 2087
rect 1793 2073 1807 2087
rect 1833 2073 1847 2087
rect 1873 2073 1887 2087
rect 2073 2073 2087 2087
rect 2113 2073 2127 2087
rect 2473 2073 2487 2087
rect 2513 2073 2527 2087
rect 2613 2073 2627 2087
rect 2673 2073 2687 2087
rect 652 2053 666 2067
rect 773 2053 787 2067
rect 833 2053 847 2067
rect 893 2053 907 2067
rect 1033 2053 1047 2067
rect 1153 2053 1167 2067
rect 1193 2053 1207 2067
rect 1293 2053 1307 2067
rect 1333 2053 1347 2067
rect 1393 2053 1407 2067
rect 1533 2053 1547 2067
rect 1573 2053 1587 2067
rect 1693 2053 1707 2067
rect 1813 2053 1827 2067
rect 1854 2053 1868 2067
rect 1973 2053 1987 2067
rect 2013 2053 2027 2067
rect 2093 2053 2107 2067
rect 2133 2053 2147 2067
rect 2253 2053 2267 2067
rect 2373 2053 2387 2067
rect 2413 2053 2427 2067
rect 2493 2053 2507 2067
rect 2533 2053 2547 2067
rect 2653 2053 2667 2067
rect 753 2033 767 2047
rect 793 2033 807 2047
rect 2873 2053 2887 2067
rect 873 2033 887 2047
rect 913 2033 927 2047
rect 1013 2033 1027 2047
rect 1053 2033 1067 2047
rect 1113 2033 1127 2047
rect 1173 2033 1187 2047
rect 1313 2033 1327 2047
rect 1672 2033 1686 2047
rect 1713 2033 1727 2047
rect 1893 2033 1907 2047
rect 1953 2033 1967 2047
rect 1994 2033 2008 2047
rect 2233 2033 2247 2047
rect 2273 2013 2287 2027
rect 833 1993 847 2007
rect 1233 1993 1247 2007
rect 1893 1993 1907 2007
rect 2393 2033 2407 2047
rect 2733 2033 2747 2047
rect 3093 2073 3107 2087
rect 3134 2073 3148 2087
rect 2993 2053 3007 2067
rect 3113 2053 3127 2067
rect 3153 2053 3167 2067
rect 3252 2053 3266 2067
rect 2853 1993 2867 2007
rect 2973 2033 2987 2047
rect 3233 2033 3247 2047
rect 3273 2033 3287 2047
rect 3013 2013 3027 2027
rect 3233 2013 3247 2027
rect 3373 2073 3387 2087
rect 3353 2053 3367 2067
rect 3393 2053 3407 2067
rect 3493 2073 3507 2087
rect 3534 2073 3548 2087
rect 3513 2053 3527 2067
rect 3553 2053 3567 2067
rect 3653 2093 3667 2107
rect 3973 2093 3987 2107
rect 3633 2073 3647 2087
rect 3593 2033 3607 2047
rect 3793 2053 3807 2067
rect 3833 2053 3847 2067
rect 3914 2053 3928 2067
rect 4193 2073 4207 2087
rect 4233 2073 4247 2087
rect 4052 2053 4066 2067
rect 4093 2053 4107 2067
rect 4173 2053 4187 2067
rect 4213 2053 4227 2067
rect 3753 2033 3767 2047
rect 3813 2033 3827 2047
rect 3893 2033 3907 2047
rect 3933 2033 3947 2047
rect 3973 2033 3987 2047
rect 4033 2033 4047 2047
rect 4073 2033 4087 2047
rect 4333 2073 4347 2087
rect 4373 2073 4387 2087
rect 4513 2073 4527 2087
rect 4573 2073 4587 2087
rect 4613 2073 4627 2087
rect 4313 2053 4327 2067
rect 4353 2053 4367 2067
rect 4413 2053 4427 2067
rect 4473 2053 4487 2067
rect 4593 2053 4607 2067
rect 4633 2053 4647 2067
rect 5332 2113 5346 2127
rect 4813 2073 4827 2087
rect 4993 2073 5007 2087
rect 5033 2073 5047 2087
rect 5093 2073 5107 2087
rect 5133 2073 5147 2087
rect 5232 2073 5246 2087
rect 5272 2073 5286 2087
rect 5333 2073 5347 2087
rect 4733 2053 4747 2067
rect 4713 2033 4727 2047
rect 4753 2033 4767 2047
rect 4792 2033 4806 2047
rect 4693 1993 4707 2007
rect 3713 1973 3727 1987
rect 4273 1973 4287 1987
rect 4873 2053 4887 2067
rect 4973 2053 4987 2067
rect 5013 2053 5027 2067
rect 5113 2053 5127 2067
rect 5154 2053 5168 2067
rect 5253 2053 5267 2067
rect 5293 2053 5307 2067
rect 4852 2033 4866 2047
rect 4892 2033 4906 2047
rect 4813 2013 4827 2027
rect 4853 2013 4867 2027
rect 5453 2073 5467 2087
rect 5513 2073 5527 2087
rect 5413 2053 5427 2067
rect 5553 2053 5567 2067
rect 5353 2033 5367 2047
rect 5152 1993 5166 2007
rect 5673 2033 5687 2047
rect 5693 2013 5707 2027
rect 5613 1973 5627 1987
rect 5673 1973 5687 1987
rect 453 1953 467 1967
rect 593 1953 607 1967
rect 2313 1953 2327 1967
rect 2933 1953 2947 1967
rect 3313 1953 3327 1967
rect 3453 1953 3467 1967
rect 4793 1953 4807 1967
rect 5673 1952 5687 1966
rect 293 1893 307 1907
rect 1293 1893 1307 1907
rect 2053 1893 2067 1907
rect 3193 1893 3207 1907
rect 3573 1893 3587 1907
rect 3713 1893 3727 1907
rect 5693 1893 5707 1907
rect 213 1813 227 1827
rect 1133 1873 1147 1887
rect 433 1833 447 1847
rect 93 1793 107 1807
rect 132 1793 146 1807
rect 193 1793 207 1807
rect 233 1793 247 1807
rect 354 1793 368 1807
rect 393 1793 407 1807
rect 633 1813 647 1827
rect 493 1793 507 1807
rect 533 1793 547 1807
rect 613 1793 627 1807
rect 653 1793 667 1807
rect 73 1773 87 1787
rect 112 1773 126 1787
rect 333 1773 347 1787
rect 373 1773 387 1787
rect 433 1773 447 1787
rect 473 1773 487 1787
rect 513 1773 527 1787
rect 573 1773 587 1787
rect 773 1813 787 1827
rect 753 1793 767 1807
rect 793 1793 807 1807
rect 573 1733 587 1747
rect 713 1733 727 1747
rect 913 1813 927 1827
rect 993 1813 1007 1827
rect 893 1793 907 1807
rect 933 1793 947 1807
rect 1033 1793 1047 1807
rect 1073 1793 1087 1807
rect 1052 1773 1066 1787
rect 1113 1773 1127 1787
rect 1193 1793 1207 1807
rect 1233 1793 1247 1807
rect 1173 1773 1187 1787
rect 1213 1773 1227 1787
rect 1774 1853 1788 1867
rect 1693 1813 1707 1827
rect 1733 1813 1747 1827
rect 1353 1793 1367 1807
rect 1393 1793 1407 1807
rect 1453 1793 1467 1807
rect 1593 1793 1607 1807
rect 1713 1793 1727 1807
rect 1373 1773 1387 1787
rect 1553 1773 1567 1787
rect 1633 1773 1647 1787
rect 1493 1753 1507 1767
rect 1533 1753 1547 1767
rect 1133 1733 1147 1747
rect 1953 1813 1967 1827
rect 1993 1813 2007 1827
rect 1813 1793 1827 1807
rect 1972 1793 1986 1807
rect 1873 1773 1887 1787
rect 1894 1753 1908 1767
rect 1773 1733 1787 1747
rect 2833 1853 2847 1867
rect 2553 1813 2567 1827
rect 2593 1813 2607 1827
rect 2633 1813 2647 1827
rect 2833 1813 2847 1827
rect 2873 1813 2887 1827
rect 2913 1813 2927 1827
rect 3053 1813 3067 1827
rect 3192 1813 3206 1827
rect 3233 1813 3247 1827
rect 3273 1813 3287 1827
rect 3433 1813 3447 1827
rect 2093 1793 2107 1807
rect 2133 1793 2147 1807
rect 2353 1793 2367 1807
rect 2393 1793 2407 1807
rect 2613 1793 2627 1807
rect 2733 1793 2747 1807
rect 2793 1793 2807 1807
rect 2852 1793 2866 1807
rect 2113 1773 2127 1787
rect 2153 1773 2167 1787
rect 2233 1773 2247 1787
rect 2273 1773 2287 1787
rect 2313 1773 2327 1787
rect 2372 1773 2386 1787
rect 2473 1773 2487 1787
rect 2513 1773 2527 1787
rect 2553 1773 2567 1787
rect 2253 1753 2267 1767
rect 2493 1753 2507 1767
rect 2753 1753 2767 1767
rect 2973 1793 2987 1807
rect 3013 1793 3027 1807
rect 3113 1793 3127 1807
rect 3153 1793 3167 1807
rect 3253 1793 3267 1807
rect 2913 1773 2927 1787
rect 2953 1773 2967 1787
rect 3053 1773 3067 1787
rect 3093 1773 3107 1787
rect 3133 1773 3147 1787
rect 3173 1773 3187 1787
rect 3353 1773 3367 1787
rect 3393 1773 3407 1787
rect 2993 1753 3007 1767
rect 3373 1753 3387 1767
rect 3573 1793 3587 1807
rect 3613 1793 3627 1807
rect 3652 1793 3666 1807
rect 3453 1773 3467 1787
rect 3493 1753 3507 1767
rect 2793 1733 2807 1747
rect 3433 1733 3447 1747
rect 3633 1773 3647 1787
rect 3673 1773 3687 1787
rect 5293 1873 5307 1887
rect 5534 1873 5548 1887
rect 5013 1833 5027 1847
rect 3772 1793 3786 1807
rect 3813 1793 3827 1807
rect 3892 1793 3906 1807
rect 3933 1793 3947 1807
rect 4053 1793 4067 1807
rect 4093 1793 4107 1807
rect 4193 1793 4207 1807
rect 4233 1793 4247 1807
rect 4333 1793 4347 1807
rect 4393 1793 4407 1807
rect 4533 1793 4547 1807
rect 4573 1793 4587 1807
rect 4652 1793 4666 1807
rect 4693 1793 4707 1807
rect 4933 1793 4947 1807
rect 4973 1793 4987 1807
rect 5153 1813 5167 1827
rect 5272 1813 5286 1827
rect 5053 1793 5067 1807
rect 5093 1793 5107 1807
rect 3752 1773 3766 1787
rect 3793 1773 3807 1787
rect 3833 1773 3847 1787
rect 3913 1773 3927 1787
rect 3973 1773 3987 1787
rect 4072 1773 4086 1787
rect 4112 1773 4126 1787
rect 4212 1773 4226 1787
rect 4254 1773 4268 1787
rect 4553 1773 4567 1787
rect 4593 1773 4607 1787
rect 4673 1773 4687 1787
rect 4752 1773 4766 1787
rect 4792 1773 4806 1787
rect 4833 1773 4847 1787
rect 4913 1773 4927 1787
rect 4953 1773 4967 1787
rect 5013 1773 5027 1787
rect 5072 1773 5086 1787
rect 5113 1773 5127 1787
rect 4313 1753 4327 1767
rect 4413 1753 4427 1767
rect 3713 1733 3727 1747
rect 5193 1773 5207 1787
rect 5234 1773 5248 1787
rect 5333 1773 5347 1787
rect 5373 1773 5387 1787
rect 5433 1773 5447 1787
rect 5493 1773 5507 1787
rect 5353 1753 5367 1767
rect 5673 1813 5687 1827
rect 5573 1793 5587 1807
rect 5613 1793 5627 1807
rect 5593 1773 5607 1787
rect 5633 1773 5647 1787
rect 5673 1773 5687 1787
rect 853 1713 867 1727
rect 1533 1713 1547 1727
rect 2053 1713 2067 1727
rect 3553 1713 3567 1727
rect 5173 1713 5187 1727
rect 5272 1713 5286 1727
rect 5294 1713 5308 1727
rect 5533 1713 5547 1727
rect 5673 1713 5687 1727
rect 173 1653 187 1667
rect 993 1653 1007 1667
rect 1273 1653 1287 1667
rect 4654 1653 4668 1667
rect 5193 1653 5207 1667
rect 5333 1653 5347 1667
rect 5613 1653 5627 1667
rect 5673 1653 5687 1667
rect 93 1593 107 1607
rect 133 1593 147 1607
rect 254 1593 268 1607
rect 73 1573 87 1587
rect 113 1573 127 1587
rect 233 1573 247 1587
rect 273 1573 287 1587
rect 393 1593 407 1607
rect 752 1593 766 1607
rect 812 1593 826 1607
rect 893 1593 907 1607
rect 933 1593 947 1607
rect 1133 1633 1147 1647
rect 1053 1593 1067 1607
rect 1113 1593 1127 1607
rect 373 1573 387 1587
rect 413 1573 427 1587
rect 473 1573 487 1587
rect 513 1573 527 1587
rect 653 1573 667 1587
rect 693 1573 707 1587
rect 793 1573 807 1587
rect 833 1573 847 1587
rect 913 1573 927 1587
rect 953 1573 967 1587
rect 993 1573 1007 1587
rect 1033 1573 1047 1587
rect 1073 1573 1087 1587
rect 1133 1573 1147 1587
rect 1173 1573 1187 1587
rect 1213 1573 1227 1587
rect 313 1553 327 1567
rect 492 1553 506 1567
rect 533 1553 547 1567
rect 673 1553 687 1567
rect 1193 1553 1207 1567
rect 1553 1633 1567 1647
rect 2113 1633 2127 1647
rect 3433 1633 3447 1647
rect 4233 1633 4247 1647
rect 1313 1593 1327 1607
rect 1353 1593 1367 1607
rect 1452 1593 1466 1607
rect 1493 1593 1507 1607
rect 1333 1573 1347 1587
rect 1373 1573 1387 1587
rect 1473 1573 1487 1587
rect 1513 1573 1527 1587
rect 993 1533 1007 1547
rect 1693 1593 1707 1607
rect 1753 1593 1767 1607
rect 1592 1573 1606 1587
rect 1634 1573 1648 1587
rect 1613 1553 1627 1567
rect 1733 1573 1747 1587
rect 1773 1573 1787 1587
rect 2033 1593 2047 1607
rect 2613 1613 2627 1627
rect 2293 1593 2307 1607
rect 2353 1593 2367 1607
rect 2713 1593 2727 1607
rect 2753 1593 2767 1607
rect 2813 1593 2827 1607
rect 2852 1593 2866 1607
rect 3193 1593 3207 1607
rect 1873 1573 1887 1587
rect 1913 1573 1927 1587
rect 2013 1573 2027 1587
rect 2053 1573 2067 1587
rect 2153 1573 2167 1587
rect 2193 1573 2207 1587
rect 2333 1573 2347 1587
rect 2373 1573 2387 1587
rect 2433 1573 2447 1587
rect 2473 1573 2487 1587
rect 2613 1573 2627 1587
rect 2693 1573 2707 1587
rect 2733 1573 2747 1587
rect 2833 1573 2847 1587
rect 2873 1573 2887 1587
rect 2973 1573 2987 1587
rect 3112 1573 3126 1587
rect 3233 1573 3247 1587
rect 1893 1553 1907 1567
rect 1953 1553 1967 1567
rect 2173 1553 2187 1567
rect 2233 1553 2247 1567
rect 2453 1553 2467 1567
rect 1833 1513 1847 1527
rect 593 1493 607 1507
rect 1553 1493 1567 1507
rect 2952 1553 2966 1567
rect 2993 1553 3007 1567
rect 3093 1553 3107 1567
rect 3133 1553 3147 1567
rect 2693 1533 2707 1547
rect 3333 1593 3347 1607
rect 3373 1593 3387 1607
rect 3353 1573 3367 1587
rect 3393 1573 3407 1587
rect 3293 1533 3307 1547
rect 3093 1513 3107 1527
rect 3773 1613 3787 1627
rect 3873 1613 3887 1627
rect 4133 1613 4147 1627
rect 4173 1613 4187 1627
rect 3473 1593 3487 1607
rect 3513 1593 3527 1607
rect 3573 1593 3587 1607
rect 3913 1593 3927 1607
rect 3993 1593 4007 1607
rect 4033 1593 4047 1607
rect 3493 1573 3507 1587
rect 3533 1573 3547 1587
rect 3633 1573 3647 1587
rect 3753 1573 3767 1587
rect 3813 1573 3827 1587
rect 3653 1553 3667 1567
rect 3433 1493 3447 1507
rect 4192 1573 4206 1587
rect 4533 1593 4547 1607
rect 4593 1593 4607 1607
rect 4292 1573 4306 1587
rect 4353 1573 4367 1587
rect 4433 1573 4447 1587
rect 4513 1573 4527 1587
rect 4573 1573 4587 1587
rect 4273 1553 4287 1567
rect 4312 1553 4326 1567
rect 4413 1553 4427 1567
rect 4453 1553 4467 1567
rect 4353 1533 4367 1547
rect 4913 1633 4927 1647
rect 4713 1593 4727 1607
rect 4753 1593 4767 1607
rect 4814 1593 4828 1607
rect 4853 1593 4867 1607
rect 4693 1573 4707 1587
rect 4733 1573 4747 1587
rect 4834 1573 4848 1587
rect 4873 1573 4887 1587
rect 4653 1513 4667 1527
rect 4952 1593 4966 1607
rect 4993 1593 5007 1607
rect 5093 1593 5107 1607
rect 5133 1593 5147 1607
rect 5253 1593 5267 1607
rect 4974 1573 4988 1587
rect 5013 1573 5027 1587
rect 5053 1573 5067 1587
rect 5113 1573 5127 1587
rect 5153 1573 5167 1587
rect 5193 1573 5207 1587
rect 5233 1573 5247 1587
rect 5273 1573 5287 1587
rect 5053 1533 5067 1547
rect 5433 1593 5447 1607
rect 5513 1593 5527 1607
rect 5553 1593 5567 1607
rect 5413 1573 5427 1587
rect 5453 1573 5467 1587
rect 5532 1573 5546 1587
rect 5573 1573 5587 1587
rect 5353 1513 5367 1527
rect 5334 1493 5348 1507
rect 5613 1493 5627 1507
rect 2533 1473 2547 1487
rect 4133 1473 4147 1487
rect 4233 1473 4247 1487
rect 4913 1473 4927 1487
rect 5673 1473 5687 1487
rect 453 1413 467 1427
rect 1254 1413 1268 1427
rect 2453 1413 2467 1427
rect 214 1333 228 1347
rect 293 1333 307 1347
rect 353 1333 367 1347
rect 413 1333 427 1347
rect 73 1313 87 1327
rect 113 1313 127 1327
rect 193 1313 207 1327
rect 233 1313 247 1327
rect 332 1313 346 1327
rect 373 1313 387 1327
rect 92 1293 106 1307
rect 134 1293 148 1307
rect 913 1333 927 1347
rect 973 1333 987 1347
rect 1173 1333 1187 1347
rect 1213 1333 1227 1347
rect 512 1313 526 1327
rect 553 1313 567 1327
rect 633 1313 647 1327
rect 673 1313 687 1327
rect 773 1313 787 1327
rect 814 1313 828 1327
rect 893 1313 907 1327
rect 933 1313 947 1327
rect 1073 1313 1087 1327
rect 1194 1313 1208 1327
rect 533 1293 547 1307
rect 652 1293 666 1307
rect 694 1293 708 1307
rect 793 1293 807 1307
rect 833 1293 847 1307
rect 1033 1293 1047 1307
rect 1113 1293 1127 1307
rect 2033 1373 2047 1387
rect 1453 1353 1467 1367
rect 1313 1333 1327 1347
rect 1353 1333 1367 1347
rect 1393 1333 1407 1347
rect 1553 1333 1567 1347
rect 1593 1333 1607 1347
rect 2333 1353 2347 1367
rect 2253 1333 2267 1347
rect 2412 1333 2426 1347
rect 4874 1413 4888 1427
rect 4553 1393 4567 1407
rect 4833 1393 4847 1407
rect 4973 1373 4987 1387
rect 5093 1373 5107 1387
rect 4953 1353 4967 1367
rect 2493 1333 2507 1347
rect 2533 1333 2547 1347
rect 4213 1333 4227 1347
rect 4293 1333 4307 1347
rect 4373 1333 4387 1347
rect 4413 1333 4427 1347
rect 4553 1333 4567 1347
rect 1333 1313 1347 1327
rect 1433 1313 1447 1327
rect 1573 1313 1587 1327
rect 1713 1313 1727 1327
rect 1673 1292 1687 1306
rect 1732 1273 1746 1287
rect 1253 1253 1267 1267
rect 1913 1313 1927 1327
rect 1992 1313 2006 1327
rect 2033 1313 2047 1327
rect 2153 1313 2167 1327
rect 2213 1313 2227 1327
rect 2393 1313 2407 1327
rect 2453 1313 2467 1327
rect 2513 1313 2527 1327
rect 2732 1313 2746 1327
rect 2774 1313 2788 1327
rect 2913 1313 2927 1327
rect 3132 1313 3146 1327
rect 3174 1313 3188 1327
rect 3253 1313 3267 1327
rect 3633 1313 3647 1327
rect 3733 1313 3747 1327
rect 3773 1313 3787 1327
rect 3814 1313 3828 1327
rect 3853 1313 3867 1327
rect 3893 1313 3907 1327
rect 4133 1313 4147 1327
rect 4273 1313 4287 1327
rect 4313 1313 4327 1327
rect 4393 1313 4407 1327
rect 4633 1313 4647 1327
rect 4673 1313 4687 1327
rect 4773 1313 4787 1327
rect 4814 1313 4828 1327
rect 4933 1313 4947 1327
rect 1973 1293 1987 1307
rect 2013 1293 2027 1307
rect 2233 1293 2247 1307
rect 2293 1293 2307 1307
rect 2613 1293 2627 1307
rect 2653 1293 2667 1307
rect 2713 1293 2727 1307
rect 2752 1293 2766 1307
rect 2793 1293 2807 1307
rect 2893 1293 2907 1307
rect 2973 1293 2987 1307
rect 3013 1293 3027 1307
rect 3113 1293 3127 1307
rect 3152 1293 3166 1307
rect 3193 1293 3207 1307
rect 3333 1293 3347 1307
rect 3413 1293 3427 1307
rect 3454 1293 3468 1307
rect 3713 1293 3727 1307
rect 3753 1293 3767 1307
rect 3873 1293 3887 1307
rect 3913 1293 3927 1307
rect 3993 1293 4007 1307
rect 4033 1293 4047 1307
rect 1873 1273 1887 1287
rect 2153 1273 2167 1287
rect 2633 1273 2647 1287
rect 2993 1273 3007 1287
rect 3293 1273 3307 1287
rect 3813 1273 3827 1287
rect 4013 1273 4027 1287
rect 3633 1253 3647 1267
rect 4173 1293 4187 1307
rect 4493 1293 4507 1307
rect 4533 1293 4547 1307
rect 4612 1293 4626 1307
rect 4653 1293 4667 1307
rect 4753 1293 4767 1307
rect 4793 1293 4807 1307
rect 4513 1273 4527 1287
rect 4893 1273 4907 1287
rect 4973 1333 4987 1347
rect 5093 1333 5107 1347
rect 5293 1333 5307 1347
rect 5333 1333 5347 1347
rect 5533 1333 5547 1347
rect 5573 1333 5587 1347
rect 5013 1313 5027 1327
rect 5053 1313 5067 1327
rect 5313 1313 5327 1327
rect 5432 1313 5446 1327
rect 5473 1313 5487 1327
rect 5553 1313 5567 1327
rect 5653 1313 5667 1327
rect 4993 1293 5007 1307
rect 5033 1293 5047 1307
rect 5073 1293 5087 1307
rect 5172 1293 5186 1307
rect 5213 1293 5227 1307
rect 5392 1293 5406 1307
rect 5453 1293 5467 1307
rect 5193 1273 5207 1287
rect 5693 1273 5707 1287
rect 1814 1233 1828 1247
rect 4073 1233 4087 1247
rect 4953 1233 4967 1247
rect 173 1173 187 1187
rect 5233 1173 5247 1187
rect 5493 1173 5507 1187
rect 573 1153 587 1167
rect 713 1153 727 1167
rect 1433 1153 1447 1167
rect 1693 1153 1707 1167
rect 1833 1153 1847 1167
rect 3573 1153 3587 1167
rect 4153 1153 4167 1167
rect 93 1113 107 1127
rect 133 1113 147 1127
rect 173 1113 187 1127
rect 353 1113 367 1127
rect 413 1113 427 1127
rect 493 1113 507 1127
rect 753 1113 767 1127
rect 793 1113 807 1127
rect 1052 1113 1066 1127
rect 1092 1113 1106 1127
rect 1133 1113 1147 1127
rect 1353 1113 1367 1127
rect 73 1093 87 1107
rect 113 1093 127 1107
rect 233 1093 247 1107
rect 272 1093 286 1107
rect 333 1093 347 1107
rect 373 1093 387 1107
rect 473 1093 487 1107
rect 513 1093 527 1107
rect 613 1093 627 1107
rect 653 1093 667 1107
rect 713 1093 727 1107
rect 773 1093 787 1107
rect 813 1093 827 1107
rect 893 1093 907 1107
rect 933 1093 947 1107
rect 1073 1093 1087 1107
rect 1113 1093 1127 1107
rect 1192 1093 1206 1107
rect 1233 1093 1247 1107
rect 1333 1093 1347 1107
rect 1373 1093 1387 1107
rect 1493 1093 1507 1107
rect 1593 1093 1607 1107
rect 1633 1093 1647 1107
rect 1733 1113 1747 1127
rect 1773 1113 1787 1127
rect 1753 1093 1767 1107
rect 1793 1093 1807 1107
rect 213 1073 227 1087
rect 254 1073 268 1087
rect 633 1073 647 1087
rect 693 1073 707 1087
rect 913 1073 927 1087
rect 973 1073 987 1087
rect 1213 1073 1227 1087
rect 1273 1073 1287 1087
rect 1473 1073 1487 1087
rect 1513 1073 1527 1087
rect 1614 1073 1628 1087
rect 1653 1073 1667 1087
rect 1693 1073 1707 1087
rect 1873 1133 1887 1147
rect 2813 1133 2827 1147
rect 2913 1133 2927 1147
rect 3253 1133 3267 1147
rect 3413 1133 3427 1147
rect 2133 1113 2147 1127
rect 2193 1113 2207 1127
rect 2253 1113 2267 1127
rect 2293 1113 2307 1127
rect 2393 1113 2407 1127
rect 2433 1113 2447 1127
rect 2793 1113 2807 1127
rect 2833 1113 2847 1127
rect 3053 1113 3067 1127
rect 3093 1113 3107 1127
rect 3173 1113 3187 1127
rect 3233 1113 3247 1127
rect 1913 1093 1927 1107
rect 1973 1093 1987 1107
rect 2013 1093 2027 1107
rect 2113 1093 2127 1107
rect 2153 1093 2167 1107
rect 2273 1093 2287 1107
rect 2314 1093 2328 1107
rect 2413 1093 2427 1107
rect 2453 1093 2467 1107
rect 2532 1093 2546 1107
rect 2573 1093 2587 1107
rect 2693 1093 2707 1107
rect 2913 1093 2927 1107
rect 3033 1093 3047 1107
rect 3073 1093 3087 1107
rect 3153 1093 3167 1107
rect 3193 1093 3207 1107
rect 1993 1073 2007 1087
rect 2553 1073 2567 1087
rect 2613 1073 2627 1087
rect 2673 1073 2687 1087
rect 2713 1073 2727 1087
rect 2073 1053 2087 1067
rect 1833 1013 1847 1027
rect 3292 1113 3306 1127
rect 3334 1113 3348 1127
rect 3393 1113 3407 1127
rect 3313 1093 3327 1107
rect 3353 1093 3367 1107
rect 3393 1053 3407 1067
rect 3453 1113 3467 1127
rect 3493 1113 3507 1127
rect 3533 1113 3547 1127
rect 3472 1093 3486 1107
rect 3513 1093 3527 1107
rect 3633 1133 3647 1147
rect 3973 1133 3987 1147
rect 4053 1133 4067 1147
rect 3673 1113 3687 1127
rect 3753 1113 3767 1127
rect 3793 1113 3807 1127
rect 3952 1113 3966 1127
rect 3993 1113 4007 1127
rect 4073 1113 4087 1127
rect 3593 1093 3607 1107
rect 4113 1093 4127 1107
rect 3573 1053 3587 1067
rect 4453 1133 4467 1147
rect 4733 1133 4747 1147
rect 4793 1133 4807 1147
rect 5033 1133 5047 1147
rect 5093 1133 5107 1147
rect 4553 1113 4567 1127
rect 4593 1113 4607 1127
rect 4913 1113 4927 1127
rect 4953 1113 4967 1127
rect 4233 1093 4247 1107
rect 4273 1093 4287 1107
rect 4353 1093 4367 1107
rect 4493 1093 4507 1107
rect 4573 1093 4587 1107
rect 4612 1093 4626 1107
rect 4693 1093 4707 1107
rect 4833 1093 4847 1107
rect 4893 1093 4907 1107
rect 4933 1093 4947 1107
rect 5033 1093 5047 1107
rect 4173 1073 4187 1087
rect 4252 1073 4266 1087
rect 4333 1073 4347 1087
rect 4373 1073 4387 1087
rect 5133 1113 5147 1127
rect 5173 1113 5187 1127
rect 5153 1093 5167 1107
rect 5193 1093 5207 1107
rect 4373 1053 4387 1067
rect 5093 1053 5107 1067
rect 4153 1033 4167 1047
rect 5373 1153 5387 1167
rect 5273 1113 5287 1127
rect 5313 1113 5327 1127
rect 5293 1093 5307 1107
rect 5333 1093 5347 1107
rect 5433 1133 5447 1147
rect 5413 1113 5427 1127
rect 5453 1113 5467 1127
rect 5653 1153 5667 1167
rect 5533 1113 5547 1127
rect 5573 1113 5587 1127
rect 5633 1113 5647 1127
rect 5553 1093 5567 1107
rect 5593 1093 5607 1107
rect 5633 1053 5647 1067
rect 5493 1033 5507 1047
rect 5373 1013 5387 1027
rect 3253 993 3267 1007
rect 3413 993 3427 1007
rect 5233 993 5247 1007
rect 5653 993 5667 1007
rect 253 933 267 947
rect 693 933 707 947
rect 973 933 987 947
rect 3033 933 3047 947
rect 5053 933 5067 947
rect 5453 933 5467 947
rect 93 833 107 847
rect 153 833 167 847
rect 193 833 207 847
rect 173 813 187 827
rect 813 893 827 907
rect 693 873 707 887
rect 313 853 327 867
rect 393 853 407 867
rect 453 853 467 867
rect 513 853 527 867
rect 733 853 747 867
rect 793 853 807 867
rect 293 833 307 847
rect 333 833 347 847
rect 432 833 446 847
rect 474 833 488 847
rect 593 833 607 847
rect 634 833 648 847
rect 714 833 728 847
rect 753 833 767 847
rect 613 813 627 827
rect 654 813 668 827
rect 853 833 867 847
rect 893 833 907 847
rect 93 793 107 807
rect 813 793 827 807
rect 873 793 887 807
rect 2413 873 2427 887
rect 1233 853 1247 867
rect 2173 853 2187 867
rect 1013 833 1027 847
rect 1053 833 1067 847
rect 1032 813 1046 827
rect 1074 813 1088 827
rect 1154 813 1168 827
rect 1193 813 1207 827
rect 1274 833 1288 847
rect 1313 833 1327 847
rect 1433 833 1447 847
rect 1474 833 1488 847
rect 1933 833 1947 847
rect 2053 833 2067 847
rect 2093 833 2107 847
rect 2153 833 2167 847
rect 2193 833 2207 847
rect 1294 813 1308 827
rect 1333 813 1347 827
rect 1553 813 1567 827
rect 1633 813 1647 827
rect 1673 813 1687 827
rect 1773 813 1787 827
rect 1833 813 1847 827
rect 1894 813 1908 827
rect 2033 813 2047 827
rect 2073 813 2087 827
rect 973 793 987 807
rect 1173 793 1187 807
rect 1233 793 1247 807
rect 1433 793 1447 807
rect 1593 793 1607 807
rect 1653 793 1667 807
rect 1793 793 1807 807
rect 1873 793 1887 807
rect 2333 833 2347 847
rect 2833 853 2847 867
rect 2873 853 2887 867
rect 2973 853 2987 867
rect 2553 833 2567 847
rect 2592 833 2606 847
rect 2693 833 2707 847
rect 2733 833 2747 847
rect 2853 833 2867 847
rect 2933 833 2947 847
rect 2973 833 2987 847
rect 2293 813 2307 827
rect 2353 813 2367 827
rect 2533 813 2547 827
rect 2573 813 2587 827
rect 2673 813 2687 827
rect 2713 813 2727 827
rect 2953 813 2967 827
rect 4313 893 4327 907
rect 4433 893 4447 907
rect 4713 893 4727 907
rect 4852 893 4866 907
rect 3092 853 3106 867
rect 3073 833 3087 847
rect 3113 833 3127 847
rect 2953 793 2967 807
rect 2253 773 2267 787
rect 2473 773 2487 787
rect 3593 853 3607 867
rect 3713 853 3727 867
rect 3753 853 3767 867
rect 3993 853 4007 867
rect 4033 853 4047 867
rect 4113 853 4127 867
rect 4153 853 4167 867
rect 3233 833 3247 847
rect 3274 833 3288 847
rect 3333 833 3347 847
rect 3373 833 3387 847
rect 3453 833 3467 847
rect 3514 833 3528 847
rect 3553 833 3567 847
rect 3353 813 3367 827
rect 3413 813 3427 827
rect 3493 813 3507 827
rect 3534 813 3548 827
rect 3614 833 3628 847
rect 3733 833 3747 847
rect 3853 833 3867 847
rect 3893 833 3907 847
rect 4013 833 4027 847
rect 4133 833 4147 847
rect 4212 833 4226 847
rect 4254 833 4268 847
rect 3833 813 3847 827
rect 3873 813 3887 827
rect 4233 813 4247 827
rect 4273 813 4287 827
rect 4413 833 4427 847
rect 4472 833 4486 847
rect 4513 833 4527 847
rect 4633 833 4647 847
rect 4493 813 4507 827
rect 4533 813 4547 827
rect 3673 793 3687 807
rect 4313 793 4327 807
rect 4393 793 4407 807
rect 4434 793 4448 807
rect 4673 813 4687 827
rect 4733 853 4747 867
rect 4793 853 4807 867
rect 4773 833 4787 847
rect 4814 833 4828 847
rect 5014 833 5028 847
rect 5313 893 5327 907
rect 5193 853 5207 867
rect 5233 853 5247 867
rect 5273 853 5287 867
rect 5093 833 5107 847
rect 5133 833 5147 847
rect 5053 813 5067 827
rect 5113 813 5127 827
rect 5153 813 5167 827
rect 5253 833 5267 847
rect 4913 793 4927 807
rect 5013 793 5027 807
rect 5193 793 5207 807
rect 5353 833 5367 847
rect 5393 833 5407 847
rect 5372 813 5386 827
rect 5412 813 5426 827
rect 5673 873 5687 887
rect 5493 833 5507 847
rect 5533 833 5547 847
rect 5633 833 5647 847
rect 5512 813 5526 827
rect 5553 813 5567 827
rect 5613 813 5627 827
rect 5654 813 5668 827
rect 954 753 968 767
rect 3173 753 3187 767
rect 3473 753 3487 767
rect 3593 753 3607 767
rect 4573 753 4587 767
rect 4713 753 4727 767
rect 5313 753 5327 767
rect 5453 753 5467 767
rect 5113 693 5127 707
rect 553 673 567 687
rect 1393 673 1407 687
rect 2853 673 2867 687
rect 3113 673 3127 687
rect 3353 673 3367 687
rect 3733 673 3747 687
rect 4473 673 4487 687
rect 4953 673 4967 687
rect 93 653 107 667
rect 193 633 207 647
rect 233 633 247 647
rect 453 633 467 647
rect 513 633 527 647
rect 1233 653 1247 667
rect 633 633 647 647
rect 1033 633 1047 647
rect 1073 633 1087 647
rect 1133 633 1147 647
rect 1173 633 1187 647
rect 93 613 107 627
rect 173 613 187 627
rect 213 613 227 627
rect 333 613 347 627
rect 374 613 388 627
rect 433 613 447 627
rect 473 613 487 627
rect 612 613 626 627
rect 653 613 667 627
rect 753 613 767 627
rect 793 613 807 627
rect 893 613 907 627
rect 933 613 947 627
rect 972 613 986 627
rect 1013 613 1027 627
rect 1053 613 1067 627
rect 1153 613 1167 627
rect 1194 613 1208 627
rect 313 593 327 607
rect 353 593 367 607
rect 713 593 727 607
rect 773 593 787 607
rect 913 593 927 607
rect 973 573 987 587
rect 1193 573 1207 587
rect 833 553 847 567
rect 1313 633 1327 647
rect 1353 633 1367 647
rect 1673 653 1687 667
rect 1833 653 1847 667
rect 2473 653 2487 667
rect 1533 633 1547 647
rect 1614 633 1628 647
rect 1293 613 1307 627
rect 1333 613 1347 627
rect 1393 613 1407 627
rect 1453 613 1467 627
rect 1493 613 1507 627
rect 1593 613 1607 627
rect 1633 613 1647 627
rect 1733 633 1747 647
rect 1774 633 1788 647
rect 2233 633 2247 647
rect 2273 633 2287 647
rect 2392 633 2406 647
rect 2433 633 2447 647
rect 2573 633 2587 647
rect 2633 633 2647 647
rect 2673 633 2687 647
rect 2733 633 2747 647
rect 2773 633 2787 647
rect 1713 613 1727 627
rect 1753 613 1767 627
rect 1873 613 1887 627
rect 1933 613 1947 627
rect 1973 613 1987 627
rect 2113 613 2127 627
rect 2153 613 2167 627
rect 2213 613 2227 627
rect 2253 613 2267 627
rect 2372 613 2386 627
rect 2414 613 2428 627
rect 2493 613 2507 627
rect 1473 593 1487 607
rect 1673 593 1687 607
rect 1953 593 1967 607
rect 2013 593 2027 607
rect 1393 553 1407 567
rect 2133 593 2147 607
rect 2373 553 2387 567
rect 2053 533 2067 547
rect 3032 633 3046 647
rect 3073 633 3087 647
rect 2613 613 2627 627
rect 2653 613 2667 627
rect 2753 613 2767 627
rect 2793 613 2807 627
rect 2853 613 2867 627
rect 2913 613 2927 627
rect 2953 613 2967 627
rect 3013 613 3027 627
rect 3053 613 3067 627
rect 2932 593 2946 607
rect 2853 533 2867 547
rect 3273 653 3287 667
rect 3192 613 3206 627
rect 3173 593 3187 607
rect 3213 593 3227 607
rect 3473 633 3487 647
rect 3553 633 3567 647
rect 3633 633 3647 647
rect 3673 633 3687 647
rect 3413 613 3427 627
rect 3533 613 3547 627
rect 3573 613 3587 627
rect 3653 613 3667 627
rect 3693 613 3707 627
rect 4053 653 4067 667
rect 4193 653 4207 667
rect 4294 653 4308 667
rect 4412 653 4426 667
rect 3913 633 3927 647
rect 3973 633 3987 647
rect 4033 633 4047 647
rect 4073 633 4087 647
rect 4113 633 4127 647
rect 4173 633 4187 647
rect 4213 633 4227 647
rect 4273 633 4287 647
rect 4313 633 4327 647
rect 4393 633 4407 647
rect 4434 633 4448 647
rect 3813 613 3827 627
rect 3933 613 3947 627
rect 3353 593 3367 607
rect 3393 593 3407 607
rect 3733 593 3747 607
rect 3793 593 3807 607
rect 3853 593 3867 607
rect 4113 593 4127 607
rect 3253 553 3267 567
rect 3433 553 3447 567
rect 4953 653 4967 667
rect 4533 633 4547 647
rect 4513 613 4527 627
rect 4553 613 4567 627
rect 4653 633 4667 647
rect 4693 633 4707 647
rect 5013 633 5027 647
rect 5054 633 5068 647
rect 5433 653 5447 667
rect 5693 653 5707 667
rect 5313 633 5327 647
rect 5353 633 5367 647
rect 4673 613 4687 627
rect 4713 613 4727 627
rect 4812 613 4826 627
rect 4913 613 4927 627
rect 5033 613 5047 627
rect 5073 613 5087 627
rect 5113 613 5127 627
rect 5193 613 5207 627
rect 5233 613 5247 627
rect 5293 613 5307 627
rect 5333 613 5347 627
rect 5473 613 5487 627
rect 5553 613 5567 627
rect 5653 613 5667 627
rect 4793 593 4807 607
rect 4834 593 4848 607
rect 5153 593 5167 607
rect 5212 593 5226 607
rect 5533 593 5547 607
rect 5573 593 5587 607
rect 4613 573 4627 587
rect 5573 573 5587 587
rect 1233 513 1247 527
rect 2573 513 2587 527
rect 3113 513 3127 527
rect 4473 513 4487 527
rect 1173 453 1187 467
rect 1313 453 1327 467
rect 2733 453 2747 467
rect 754 433 768 447
rect 1154 393 1168 407
rect 113 373 127 387
rect 293 373 307 387
rect 493 373 507 387
rect 533 373 547 387
rect 593 373 607 387
rect 753 373 767 387
rect 913 373 927 387
rect 973 373 987 387
rect 93 353 107 367
rect 133 353 147 367
rect 192 353 206 367
rect 233 353 247 367
rect 213 333 227 347
rect 353 353 367 367
rect 393 353 407 367
rect 513 353 527 367
rect 553 353 567 367
rect 652 353 666 367
rect 693 353 707 367
rect 793 353 807 367
rect 833 353 847 367
rect 953 353 967 367
rect 993 353 1007 367
rect 1053 353 1067 367
rect 1093 353 1107 367
rect 313 333 327 347
rect 373 333 387 347
rect 593 333 607 347
rect 632 333 646 347
rect 673 333 687 347
rect 712 333 726 347
rect 813 333 827 347
rect 853 333 867 347
rect 1073 333 1087 347
rect 1213 353 1227 367
rect 1253 353 1267 367
rect 1453 433 1467 447
rect 1973 433 1987 447
rect 1333 373 1347 387
rect 1393 373 1407 387
rect 1373 353 1387 367
rect 1413 353 1427 367
rect 1173 333 1187 347
rect 1233 333 1247 347
rect 1273 333 1287 347
rect 1313 333 1327 347
rect 1753 373 1767 387
rect 1793 373 1807 387
rect 1873 373 1887 387
rect 1513 353 1527 367
rect 1554 353 1568 367
rect 1653 353 1667 367
rect 1773 353 1787 367
rect 1873 353 1887 367
rect 1913 353 1927 367
rect 1533 333 1547 347
rect 1613 333 1627 347
rect 1693 333 1707 347
rect 1893 333 1907 347
rect 2113 413 2127 427
rect 2333 413 2347 427
rect 2033 373 2047 387
rect 2153 373 2167 387
rect 2193 373 2207 387
rect 2013 353 2027 367
rect 2053 353 2067 367
rect 2173 353 2187 367
rect 2394 373 2408 387
rect 2513 373 2527 387
rect 2573 373 2587 387
rect 2653 373 2667 387
rect 2693 373 2707 387
rect 4433 433 4447 447
rect 4933 433 4947 447
rect 2873 373 2887 387
rect 3813 373 3827 387
rect 3873 373 3887 387
rect 4213 373 4227 387
rect 4253 373 4267 387
rect 4332 373 4346 387
rect 4373 373 4387 387
rect 2373 353 2387 367
rect 2413 353 2427 367
rect 2493 353 2507 367
rect 2553 353 2567 367
rect 2593 353 2607 367
rect 2673 353 2687 367
rect 2732 353 2746 367
rect 2773 353 2787 367
rect 2813 353 2827 367
rect 2093 333 2107 347
rect 2793 333 2807 347
rect 2932 353 2946 367
rect 2974 353 2988 367
rect 3353 353 3367 367
rect 3433 353 3447 367
rect 3473 353 3487 367
rect 3853 353 3867 367
rect 3893 353 3907 367
rect 3973 353 3987 367
rect 4013 353 4027 367
rect 4133 353 4147 367
rect 4233 353 4247 367
rect 4273 353 4287 367
rect 4353 353 4367 367
rect 4673 413 4687 427
rect 4473 373 4487 387
rect 4513 373 4527 387
rect 4592 373 4606 387
rect 4633 373 4647 387
rect 4753 373 4767 387
rect 5353 413 5367 427
rect 5493 413 5507 427
rect 4993 373 5007 387
rect 5033 373 5047 387
rect 4494 353 4508 367
rect 4613 353 4627 367
rect 4733 353 4747 367
rect 4773 353 4787 367
rect 4833 353 4847 367
rect 4873 353 4887 367
rect 4933 353 4947 367
rect 5013 353 5027 367
rect 2913 333 2927 347
rect 2952 333 2966 347
rect 2993 333 3007 347
rect 3053 333 3067 347
rect 3132 333 3146 347
rect 3173 333 3187 347
rect 3413 333 3427 347
rect 3453 333 3467 347
rect 3493 333 3507 347
rect 3573 333 3587 347
rect 3653 333 3667 347
rect 3713 333 3727 347
rect 3753 333 3767 347
rect 3993 333 4007 347
rect 4033 333 4047 347
rect 4433 333 4447 347
rect 4853 333 4867 347
rect 1073 313 1087 327
rect 293 293 307 307
rect 2313 313 2327 327
rect 3293 313 3307 327
rect 4093 313 4107 327
rect 4933 293 4947 307
rect 5153 373 5167 387
rect 5213 373 5227 387
rect 5293 373 5307 387
rect 5133 353 5147 367
rect 5172 353 5186 367
rect 5272 353 5286 367
rect 5313 353 5327 367
rect 5393 353 5407 367
rect 5433 353 5447 367
rect 5533 353 5547 367
rect 5573 353 5587 367
rect 5653 353 5667 367
rect 5413 333 5427 347
rect 5453 333 5467 347
rect 5493 333 5507 347
rect 5553 333 5567 347
rect 5593 333 5607 347
rect 5353 313 5367 327
rect 5693 313 5707 327
rect 33 273 47 287
rect 2092 273 2106 287
rect 5073 273 5087 287
rect 5353 213 5367 227
rect 1533 193 1547 207
rect 93 173 107 187
rect 993 173 1007 187
rect 1073 173 1087 187
rect 1453 173 1467 187
rect 333 153 347 167
rect 373 153 387 167
rect 433 153 447 167
rect 473 153 487 167
rect 93 133 107 147
rect 152 133 166 147
rect 193 133 207 147
rect 313 133 327 147
rect 353 133 367 147
rect 453 133 467 147
rect 493 133 507 147
rect 573 133 587 147
rect 613 133 627 147
rect 713 133 727 147
rect 753 133 767 147
rect 853 133 867 147
rect 893 133 907 147
rect 993 133 1007 147
rect 173 113 187 127
rect 593 113 607 127
rect 653 113 667 127
rect 733 113 747 127
rect 813 113 827 127
rect 873 113 887 127
rect 1253 153 1267 167
rect 1313 154 1327 168
rect 1393 154 1407 168
rect 1133 133 1147 147
rect 1174 133 1188 147
rect 1233 133 1247 147
rect 1273 133 1287 147
rect 1433 133 1447 147
rect 1733 173 1747 187
rect 1973 173 1987 187
rect 2653 173 2667 187
rect 2853 173 2867 187
rect 1593 153 1607 167
rect 1633 153 1647 167
rect 1873 153 1887 167
rect 1913 153 1927 167
rect 2073 153 2087 167
rect 2113 153 2127 167
rect 2373 153 2387 167
rect 2413 153 2427 167
rect 2692 153 2706 167
rect 2733 153 2747 167
rect 2953 153 2967 167
rect 2993 153 3007 167
rect 3073 153 3087 167
rect 3173 153 3187 167
rect 3213 153 3227 167
rect 1613 133 1627 147
rect 1653 133 1667 147
rect 1793 133 1807 147
rect 1853 133 1867 147
rect 1894 133 1908 147
rect 2013 133 2027 147
rect 2093 133 2107 147
rect 2133 133 2147 147
rect 2233 133 2247 147
rect 2352 133 2366 147
rect 2393 133 2407 147
rect 2513 133 2527 147
rect 2633 133 2647 147
rect 2833 133 2847 147
rect 1153 113 1167 127
rect 2213 113 2227 127
rect 2254 113 2268 127
rect 2493 113 2507 127
rect 2553 113 2567 127
rect 953 73 967 87
rect 3333 153 3347 167
rect 4353 173 4367 187
rect 4693 173 4707 187
rect 3913 153 3927 167
rect 3954 153 3968 167
rect 4033 153 4047 167
rect 4093 153 4107 167
rect 3393 133 3407 147
rect 3473 133 3487 147
rect 3533 133 3547 147
rect 3593 133 3607 147
rect 3653 133 3667 147
rect 3772 133 3786 147
rect 3814 133 3828 147
rect 3893 133 3907 147
rect 3933 133 3947 147
rect 3513 113 3527 127
rect 3553 113 3567 127
rect 3633 113 3647 127
rect 3673 113 3687 127
rect 3733 113 3747 127
rect 3794 113 3808 127
rect 4213 153 4227 167
rect 4993 153 5007 167
rect 5073 153 5087 167
rect 5113 153 5127 167
rect 5273 153 5287 167
rect 5493 193 5507 207
rect 5393 153 5407 167
rect 5433 153 5447 167
rect 5653 173 5667 187
rect 5573 153 5587 167
rect 4173 133 4187 147
rect 4293 133 4307 147
rect 4353 133 4367 147
rect 4413 133 4427 147
rect 4552 133 4566 147
rect 4594 133 4608 147
rect 4653 133 4667 147
rect 4793 133 4807 147
rect 4833 133 4847 147
rect 4913 133 4927 147
rect 5253 133 5267 147
rect 5293 133 5307 147
rect 5413 133 5427 147
rect 5453 133 5467 147
rect 5653 133 5667 147
rect 4273 113 4287 127
rect 4313 113 4327 127
rect 4393 113 4407 127
rect 4433 113 4447 127
rect 4573 113 4587 127
rect 4493 93 4507 107
rect 4813 113 4827 127
rect 4893 113 4907 127
rect 4933 113 4947 127
rect 3593 73 3607 87
rect 4113 73 4127 87
rect 4733 73 4747 87
rect 3253 53 3267 67
rect 253 33 267 47
<< metal2 >>
rect 4127 5776 4153 5783
rect 4287 5776 4793 5783
rect 4947 5776 5433 5783
rect 4027 5756 4233 5763
rect 4327 5756 4963 5763
rect 1247 5736 1513 5743
rect 1527 5736 1893 5743
rect 4956 5743 4963 5756
rect 4987 5756 5093 5763
rect 5247 5756 5553 5763
rect 4956 5736 5053 5743
rect 5287 5736 5533 5743
rect 607 5716 1313 5723
rect 4747 5713 4749 5727
rect 5027 5716 5053 5723
rect 627 5696 2113 5703
rect 2307 5696 2933 5703
rect 116 5680 313 5683
rect 113 5676 313 5680
rect 113 5667 127 5676
rect 213 5667 227 5676
rect 327 5676 833 5683
rect 887 5676 1013 5683
rect 1627 5676 1713 5683
rect 1727 5676 1773 5683
rect 2147 5676 2813 5683
rect 3747 5676 3833 5683
rect 4286 5673 4287 5680
rect 3233 5667 3247 5673
rect 4273 5667 4287 5673
rect 807 5656 913 5663
rect 927 5653 933 5667
rect 1407 5653 1413 5667
rect 1467 5653 1473 5667
rect 1500 5663 1513 5667
rect 1496 5653 1513 5663
rect 1567 5653 1573 5667
rect 1716 5660 1943 5663
rect 1713 5656 1943 5660
rect 1013 5647 1027 5653
rect 67 5636 93 5643
rect 147 5636 193 5643
rect 193 5627 207 5633
rect 327 5633 333 5647
rect 387 5633 393 5647
rect 456 5636 492 5643
rect 233 5627 247 5633
rect 347 5613 353 5627
rect 456 5623 463 5636
rect 528 5633 533 5647
rect 687 5636 753 5643
rect 767 5636 872 5643
rect 893 5633 894 5640
rect 947 5633 953 5647
rect 1067 5633 1073 5647
rect 1127 5633 1133 5647
rect 1187 5633 1193 5647
rect 1327 5636 1373 5643
rect 1496 5643 1503 5653
rect 1713 5647 1727 5656
rect 1427 5636 1503 5643
rect 1527 5636 1553 5643
rect 1607 5633 1612 5647
rect 1648 5636 1673 5643
rect 1907 5633 1913 5647
rect 1936 5643 1943 5656
rect 2407 5660 2464 5663
rect 2407 5656 2467 5660
rect 2453 5647 2467 5656
rect 2527 5656 2753 5663
rect 2653 5647 2667 5656
rect 2907 5653 2913 5667
rect 2967 5656 2993 5663
rect 3427 5653 3433 5667
rect 3487 5656 3513 5663
rect 4200 5663 4213 5667
rect 4187 5656 4213 5663
rect 4200 5653 4213 5656
rect 4286 5660 4287 5667
rect 4308 5653 4313 5667
rect 4915 5660 5073 5663
rect 4913 5656 5073 5660
rect 4913 5647 4927 5656
rect 1936 5636 1953 5643
rect 1967 5636 2033 5643
rect 2047 5636 2132 5643
rect 2168 5636 2253 5643
rect 2427 5633 2432 5647
rect 2453 5640 2454 5647
rect 2507 5636 2573 5643
rect 2587 5640 2643 5643
rect 2587 5636 2647 5640
rect 633 5627 647 5633
rect 893 5627 907 5633
rect 2293 5627 2307 5633
rect 2633 5627 2647 5636
rect 2707 5633 2713 5647
rect 2807 5633 2813 5647
rect 2867 5633 2873 5647
rect 2947 5633 2953 5647
rect 3127 5636 3173 5643
rect 3267 5636 3313 5643
rect 3467 5636 3513 5643
rect 3567 5636 3613 5643
rect 4247 5636 4293 5643
rect 4347 5633 4353 5647
rect 4847 5633 4853 5647
rect 4867 5636 4892 5643
rect 4926 5640 4927 5647
rect 4933 5633 4934 5640
rect 5167 5633 5173 5647
rect 5227 5633 5233 5647
rect 5547 5633 5553 5647
rect 427 5616 463 5623
rect 487 5613 492 5627
rect 528 5616 612 5623
rect 633 5620 634 5627
rect 653 5613 654 5620
rect 307 5596 513 5603
rect 653 5603 667 5613
rect 567 5600 667 5603
rect 693 5607 707 5613
rect 567 5596 663 5600
rect 893 5620 894 5627
rect 793 5607 807 5613
rect 993 5607 1007 5613
rect 1167 5616 1293 5623
rect 1667 5616 1693 5623
rect 1033 5603 1047 5613
rect 1033 5600 1213 5603
rect 1036 5596 1213 5600
rect 1327 5596 1433 5603
rect 1733 5603 1747 5613
rect 1987 5613 1993 5627
rect 2347 5613 2353 5627
rect 2487 5616 2513 5623
rect 2687 5613 2693 5627
rect 3067 5616 3133 5623
rect 3213 5623 3227 5633
rect 3213 5620 3413 5623
rect 3216 5616 3413 5620
rect 1933 5607 1947 5613
rect 2193 5607 2207 5613
rect 2433 5607 2447 5613
rect 1733 5600 1833 5603
rect 1736 5596 1833 5600
rect 2047 5596 2192 5603
rect 2206 5600 2207 5607
rect 2228 5596 2292 5603
rect 2328 5596 2393 5603
rect 2587 5596 2753 5603
rect 2833 5603 2847 5613
rect 2833 5600 2913 5603
rect 2836 5596 2913 5600
rect 2927 5596 3033 5603
rect 3047 5596 3153 5603
rect 3367 5596 3793 5603
rect 4136 5603 4143 5633
rect 4933 5627 4947 5633
rect 4807 5616 4893 5623
rect 5067 5613 5073 5627
rect 5087 5620 5123 5623
rect 5087 5616 5127 5620
rect 4136 5596 4213 5603
rect 5013 5603 5027 5613
rect 5113 5607 5127 5616
rect 5266 5613 5267 5620
rect 5288 5613 5293 5627
rect 5386 5613 5387 5620
rect 5408 5613 5413 5627
rect 5587 5613 5593 5627
rect 5253 5607 5267 5613
rect 5373 5607 5387 5613
rect 4867 5600 5027 5603
rect 4867 5596 5023 5600
rect 5047 5596 5073 5603
rect 5266 5600 5267 5607
rect 5386 5600 5387 5607
rect 247 5576 393 5583
rect 907 5576 1133 5583
rect 1427 5576 1653 5583
rect 1833 5583 1847 5593
rect 1833 5580 1973 5583
rect 1836 5576 1973 5580
rect 2207 5576 2333 5583
rect 2867 5576 2993 5583
rect 3007 5576 3453 5583
rect 3707 5576 3753 5583
rect 47 5556 123 5563
rect 116 5543 123 5556
rect 207 5556 333 5563
rect 347 5556 553 5563
rect 647 5556 833 5563
rect 967 5556 1073 5563
rect 1227 5556 1613 5563
rect 1627 5553 1633 5567
rect 2267 5556 2713 5563
rect 3247 5556 3513 5563
rect 3527 5556 3853 5563
rect 4127 5556 4373 5563
rect 4387 5556 4433 5563
rect 4847 5556 4973 5563
rect 116 5536 233 5543
rect 707 5536 1193 5543
rect 1487 5536 1833 5543
rect 1847 5536 2073 5543
rect 3627 5536 3913 5543
rect 4427 5536 4813 5543
rect 5067 5536 5353 5543
rect 5367 5536 5673 5543
rect 527 5516 733 5523
rect 747 5516 1513 5523
rect 1987 5516 3392 5523
rect 3428 5516 3773 5523
rect 3827 5516 4113 5523
rect 4227 5516 4773 5523
rect 5127 5516 5373 5523
rect 287 5496 473 5503
rect 487 5496 593 5503
rect 927 5496 1293 5503
rect 4156 5496 4413 5503
rect 4156 5487 4163 5496
rect 4507 5496 4733 5503
rect 4776 5503 4783 5513
rect 4776 5496 5073 5503
rect 5087 5496 5233 5503
rect 5307 5496 5573 5503
rect 67 5476 453 5483
rect 687 5476 833 5483
rect 1147 5476 1213 5483
rect 1587 5476 1853 5483
rect 3367 5476 3433 5483
rect 4147 5473 4153 5487
rect 4376 5480 4453 5483
rect 4373 5476 4453 5480
rect 4373 5467 4387 5476
rect 4467 5476 4893 5483
rect 4907 5476 5093 5483
rect 5267 5476 5413 5483
rect 5133 5467 5147 5473
rect 5513 5467 5527 5473
rect 416 5460 603 5463
rect 413 5456 603 5460
rect 413 5447 427 5456
rect 596 5447 603 5456
rect 667 5456 693 5463
rect 707 5456 753 5463
rect 1087 5456 1173 5463
rect 1567 5456 1673 5463
rect 1687 5456 2033 5463
rect 2527 5456 2573 5463
rect 2707 5456 2833 5463
rect 2987 5456 3053 5463
rect 3167 5456 3233 5463
rect 1313 5447 1327 5453
rect 47 5433 53 5447
rect 107 5433 113 5447
rect 327 5436 373 5443
rect 527 5433 532 5447
rect 568 5436 593 5443
rect 907 5433 913 5447
rect 1247 5436 1273 5443
rect 1367 5436 1453 5443
rect 1053 5427 1067 5433
rect 1673 5427 1687 5433
rect 147 5413 153 5427
rect 227 5413 233 5427
rect 287 5413 293 5427
rect 93 5407 107 5413
rect 353 5407 367 5413
rect 93 5400 113 5407
rect 96 5396 113 5400
rect 100 5393 113 5396
rect 267 5396 313 5403
rect 467 5416 493 5423
rect 393 5403 407 5413
rect 533 5403 547 5413
rect 576 5416 672 5423
rect 576 5403 583 5416
rect 708 5413 713 5427
rect 767 5413 773 5427
rect 847 5416 873 5423
rect 887 5413 893 5427
rect 947 5416 993 5423
rect 1107 5416 1153 5423
rect 1347 5413 1353 5427
rect 1407 5416 1433 5423
rect 1527 5413 1533 5427
rect 1587 5413 1593 5427
rect 1713 5427 1727 5433
rect 1853 5427 1867 5433
rect 2073 5433 2074 5440
rect 2373 5443 2387 5453
rect 3373 5447 3387 5453
rect 3887 5456 4033 5463
rect 4047 5456 4233 5463
rect 4567 5460 4623 5463
rect 4567 5456 4627 5460
rect 3413 5447 3427 5453
rect 4613 5447 4627 5456
rect 4647 5460 4764 5463
rect 4647 5456 4767 5460
rect 4753 5447 4767 5456
rect 4827 5456 4983 5463
rect 4976 5447 4983 5456
rect 5027 5456 5053 5463
rect 5227 5453 5232 5467
rect 5253 5453 5254 5460
rect 5253 5447 5267 5453
rect 5413 5447 5427 5453
rect 5593 5447 5607 5453
rect 2236 5440 2483 5443
rect 2073 5427 2087 5433
rect 2113 5427 2127 5433
rect 1947 5416 1973 5423
rect 2027 5416 2052 5423
rect 2073 5420 2074 5427
rect 2233 5436 2487 5440
rect 2233 5427 2247 5436
rect 2473 5427 2487 5436
rect 3187 5436 3352 5443
rect 3373 5440 3374 5447
rect 3366 5433 3367 5440
rect 3587 5436 3633 5443
rect 3687 5436 3792 5443
rect 3828 5436 3913 5443
rect 3927 5436 3973 5443
rect 4233 5433 4234 5440
rect 4427 5433 4432 5447
rect 4466 5433 4467 5440
rect 4488 5436 4573 5443
rect 4727 5433 4732 5447
rect 4753 5440 4754 5447
rect 4776 5440 4853 5443
rect 4773 5436 4853 5440
rect 2387 5413 2392 5427
rect 2428 5413 2433 5427
rect 2627 5416 2713 5423
rect 2767 5413 2773 5427
rect 2847 5413 2853 5427
rect 3007 5416 3113 5423
rect 1293 5407 1307 5413
rect 393 5400 583 5403
rect 396 5396 583 5400
rect 727 5393 733 5407
rect 1067 5396 1133 5403
rect 1133 5387 1147 5393
rect 367 5376 393 5383
rect 547 5376 773 5383
rect 927 5376 1093 5383
rect 1356 5403 1363 5413
rect 2893 5407 2907 5413
rect 1356 5396 1413 5403
rect 1467 5396 1493 5403
rect 1627 5396 1693 5403
rect 1887 5396 1933 5403
rect 1987 5393 1993 5407
rect 2016 5396 2093 5403
rect 1173 5387 1187 5393
rect 1553 5383 1567 5393
rect 1247 5380 1567 5383
rect 1833 5387 1847 5393
rect 1247 5376 1563 5380
rect 2016 5383 2023 5396
rect 2167 5393 2172 5407
rect 2208 5393 2213 5407
rect 2467 5396 2673 5403
rect 2727 5393 2733 5407
rect 2807 5393 2813 5407
rect 2893 5400 2894 5407
rect 2886 5393 2887 5400
rect 2253 5383 2267 5393
rect 1887 5380 2267 5383
rect 2873 5383 2887 5393
rect 2973 5387 2987 5393
rect 2873 5380 2973 5383
rect 1887 5376 2263 5380
rect 2875 5376 2973 5380
rect 3136 5403 3143 5433
rect 3353 5427 3367 5433
rect 4233 5427 4247 5433
rect 4453 5427 4467 5433
rect 4773 5427 4787 5436
rect 4976 5436 4993 5447
rect 4980 5433 4993 5436
rect 5107 5433 5113 5447
rect 5167 5433 5173 5447
rect 5367 5433 5373 5447
rect 5467 5436 5493 5443
rect 3187 5416 3233 5423
rect 3376 5416 3393 5423
rect 3136 5396 3193 5403
rect 3207 5393 3212 5407
rect 3248 5393 3253 5407
rect 3376 5403 3383 5416
rect 3407 5416 3513 5423
rect 3567 5416 3612 5423
rect 3648 5413 3653 5427
rect 3786 5413 3787 5420
rect 3773 5407 3787 5413
rect 3267 5396 3383 5403
rect 3447 5396 3493 5403
rect 3547 5396 3573 5403
rect 3766 5393 3767 5400
rect 3786 5400 3787 5407
rect 3808 5394 3813 5407
rect 3893 5407 3907 5413
rect 3808 5393 3820 5394
rect 3987 5416 4013 5423
rect 4147 5416 4193 5423
rect 4207 5413 4212 5427
rect 4233 5420 4234 5427
rect 4607 5413 4612 5427
rect 4648 5416 4673 5423
rect 4933 5427 4947 5433
rect 4887 5414 4893 5427
rect 4880 5413 4893 5414
rect 5033 5427 5047 5433
rect 5156 5423 5163 5433
rect 5553 5427 5567 5433
rect 5633 5427 5647 5433
rect 5047 5416 5163 5423
rect 5267 5416 5293 5423
rect 5566 5420 5567 5427
rect 5573 5413 5574 5420
rect 5633 5420 5634 5427
rect 5626 5413 5627 5420
rect 3933 5407 3947 5413
rect 4493 5407 4507 5413
rect 4733 5403 4747 5413
rect 5393 5407 5407 5413
rect 4733 5400 4873 5403
rect 4736 5396 4873 5400
rect 3013 5383 3027 5393
rect 3753 5387 3767 5393
rect 3013 5380 3053 5383
rect 3016 5376 3053 5380
rect 3067 5376 3173 5383
rect 3766 5380 3767 5387
rect 3827 5376 3893 5383
rect 3987 5376 4033 5383
rect 4213 5383 4227 5393
rect 5393 5400 5413 5407
rect 5396 5396 5413 5400
rect 5400 5393 5413 5396
rect 5436 5403 5443 5413
rect 5573 5403 5587 5413
rect 5436 5400 5587 5403
rect 5613 5403 5627 5413
rect 5613 5400 5673 5403
rect 5436 5396 5584 5400
rect 5615 5396 5673 5400
rect 4213 5380 4313 5383
rect 4216 5376 4313 5380
rect 4327 5376 4653 5383
rect 4747 5376 5033 5383
rect 5436 5383 5443 5396
rect 5147 5376 5443 5383
rect 5527 5376 5653 5383
rect 187 5356 413 5363
rect 1187 5356 1553 5363
rect 1787 5356 1993 5363
rect 2007 5356 2213 5363
rect 2547 5356 3073 5363
rect 3527 5356 3653 5363
rect 3987 5356 4673 5363
rect 4687 5353 4693 5367
rect 4867 5356 5213 5363
rect 827 5336 1113 5343
rect 1127 5336 1233 5343
rect 1256 5336 1393 5343
rect 887 5316 993 5323
rect 1256 5323 1263 5336
rect 1447 5336 2053 5343
rect 3147 5336 3553 5343
rect 4307 5336 4893 5343
rect 4947 5336 5593 5343
rect 1007 5316 1263 5323
rect 1307 5316 1373 5323
rect 1647 5316 1953 5323
rect 2907 5316 3053 5323
rect 3207 5316 3413 5323
rect 3427 5316 3832 5323
rect 3868 5316 4153 5323
rect 4567 5316 4853 5323
rect 5087 5313 5093 5327
rect 5447 5316 5553 5323
rect 767 5296 893 5303
rect 1227 5296 1593 5303
rect 3907 5296 3973 5303
rect 4227 5296 4592 5303
rect 4628 5296 4873 5303
rect 1507 5276 1753 5283
rect 2727 5276 3033 5283
rect 3587 5276 3873 5283
rect 4387 5276 4733 5283
rect 4747 5276 5433 5283
rect 127 5256 153 5263
rect 967 5256 1233 5263
rect 1247 5256 1773 5263
rect 2347 5256 3193 5263
rect 3867 5256 4413 5263
rect 107 5236 273 5243
rect 1147 5236 1293 5243
rect 1307 5236 1433 5243
rect 1447 5236 1933 5243
rect 2127 5236 2283 5243
rect 2276 5227 2283 5236
rect 2387 5236 2993 5243
rect 3767 5236 3933 5243
rect 3947 5236 4272 5243
rect 4308 5236 4493 5243
rect 5131 5233 5133 5247
rect 147 5216 333 5223
rect 347 5216 473 5223
rect 1347 5216 1693 5223
rect 1707 5216 2213 5223
rect 2287 5216 2353 5223
rect 2687 5216 2873 5223
rect 3387 5216 3453 5223
rect 3707 5216 3933 5223
rect 5507 5216 5533 5223
rect 287 5200 463 5203
rect 287 5196 467 5200
rect 453 5187 467 5196
rect 787 5196 973 5203
rect 1127 5196 1233 5203
rect 1567 5196 1773 5203
rect 1847 5203 1860 5207
rect 1847 5200 1862 5203
rect 1847 5193 1867 5200
rect 1887 5196 2423 5203
rect 1853 5187 1867 5193
rect 1973 5187 1987 5196
rect 87 5176 173 5183
rect 187 5173 193 5187
rect 247 5173 253 5187
rect 376 5180 453 5183
rect 333 5167 347 5173
rect 227 5156 273 5163
rect 373 5176 453 5180
rect 373 5167 387 5176
rect 527 5176 573 5183
rect 616 5180 693 5183
rect 613 5176 693 5180
rect 613 5167 627 5176
rect 773 5173 774 5180
rect 1387 5173 1393 5187
rect 1467 5173 1473 5187
rect 773 5167 787 5173
rect 1293 5167 1307 5173
rect 73 5147 87 5153
rect 433 5147 447 5153
rect 127 5133 133 5147
rect 307 5133 313 5147
rect 747 5153 752 5167
rect 773 5160 774 5167
rect 836 5156 872 5163
rect 473 5143 487 5153
rect 473 5140 573 5143
rect 476 5136 573 5140
rect 667 5133 672 5147
rect 708 5136 753 5143
rect 836 5143 843 5156
rect 906 5153 907 5160
rect 928 5156 973 5163
rect 1427 5153 1433 5167
rect 1533 5163 1547 5173
rect 1866 5180 1867 5187
rect 1873 5173 1874 5180
rect 1920 5183 1933 5187
rect 1916 5173 1933 5183
rect 2256 5180 2393 5183
rect 2253 5176 2393 5180
rect 1573 5167 1587 5173
rect 1873 5167 1887 5173
rect 1487 5160 1547 5163
rect 1487 5156 1543 5160
rect 1573 5160 1574 5167
rect 1566 5153 1567 5160
rect 1707 5153 1713 5167
rect 1787 5156 1833 5163
rect 893 5147 907 5153
rect 807 5136 843 5143
rect 353 5127 367 5133
rect 793 5127 807 5133
rect 107 5116 153 5123
rect 367 5116 433 5123
rect 906 5140 907 5147
rect 1033 5147 1047 5153
rect 1127 5133 1133 5147
rect 1186 5133 1187 5140
rect 1208 5136 1253 5143
rect 1333 5143 1347 5153
rect 1473 5147 1487 5153
rect 1333 5140 1473 5143
rect 1336 5136 1473 5140
rect 1553 5147 1567 5153
rect 1916 5147 1923 5173
rect 2253 5167 2267 5176
rect 2416 5183 2423 5196
rect 2447 5200 2843 5203
rect 2447 5196 2847 5200
rect 2833 5187 2847 5196
rect 2416 5176 2593 5183
rect 2647 5173 2653 5187
rect 2887 5200 3103 5203
rect 2887 5196 3107 5200
rect 2873 5187 2887 5193
rect 3093 5187 3107 5196
rect 3396 5196 3753 5203
rect 2927 5176 2952 5183
rect 2988 5173 2993 5187
rect 3167 5176 3193 5183
rect 3287 5173 3293 5187
rect 3396 5183 3403 5196
rect 3967 5196 4232 5203
rect 4268 5196 4333 5203
rect 4536 5196 4823 5203
rect 3316 5176 3403 5183
rect 3316 5167 3323 5176
rect 3396 5167 3403 5176
rect 3556 5180 3843 5183
rect 3513 5167 3527 5173
rect 1947 5153 1953 5167
rect 2027 5156 2073 5163
rect 2127 5153 2133 5167
rect 2200 5163 2213 5167
rect 2196 5153 2213 5163
rect 2487 5153 2493 5167
rect 2627 5153 2633 5167
rect 2687 5156 2733 5163
rect 2960 5163 2973 5167
rect 2956 5160 2973 5163
rect 1607 5136 1653 5143
rect 1747 5133 1753 5147
rect 2067 5136 2093 5143
rect 2196 5143 2203 5153
rect 2147 5136 2203 5143
rect 2227 5133 2233 5147
rect 2287 5133 2293 5147
rect 2320 5143 2332 5147
rect 2316 5140 2332 5143
rect 2313 5133 2332 5140
rect 2366 5133 2367 5140
rect 2388 5136 2433 5143
rect 2447 5133 2453 5147
rect 2476 5136 2513 5143
rect 853 5127 867 5133
rect 1073 5127 1087 5133
rect 1173 5127 1187 5133
rect 1096 5116 1152 5123
rect 1096 5103 1103 5116
rect 1173 5120 1174 5127
rect 1313 5123 1327 5133
rect 2133 5127 2147 5133
rect 1313 5120 1463 5123
rect 1316 5116 1463 5120
rect 1456 5107 1463 5116
rect 2313 5127 2327 5133
rect 2353 5127 2367 5133
rect 2366 5120 2367 5127
rect 2476 5123 2483 5136
rect 2853 5143 2867 5153
rect 2953 5153 2973 5160
rect 3047 5156 3073 5163
rect 3247 5153 3253 5167
rect 3307 5156 3323 5167
rect 3307 5153 3320 5156
rect 3347 5153 3353 5167
rect 3553 5176 3843 5180
rect 3553 5167 3567 5176
rect 3693 5167 3707 5176
rect 3627 5156 3653 5163
rect 3706 5160 3707 5167
rect 3728 5156 3813 5163
rect 3836 5163 3843 5176
rect 4193 5173 4194 5180
rect 4536 5183 4543 5196
rect 4507 5176 4543 5183
rect 4555 5180 4633 5183
rect 4553 5176 4633 5180
rect 4193 5167 4207 5173
rect 4553 5167 4567 5176
rect 4816 5167 4823 5196
rect 4876 5180 4983 5183
rect 4873 5176 4983 5180
rect 4873 5167 4887 5176
rect 4976 5167 4983 5176
rect 5033 5167 5047 5173
rect 3836 5156 3913 5163
rect 4167 5153 4172 5167
rect 4193 5160 4194 5167
rect 4236 5156 4332 5163
rect 2953 5147 2967 5153
rect 2853 5140 2913 5143
rect 2856 5136 2913 5140
rect 3113 5147 3127 5153
rect 3307 5136 3372 5143
rect 3408 5133 3413 5147
rect 3467 5136 3533 5143
rect 3587 5133 3593 5147
rect 3687 5134 3692 5147
rect 4236 5147 4243 5156
rect 4368 5153 4373 5167
rect 4566 5160 4567 5167
rect 4588 5153 4593 5167
rect 4707 5153 4713 5167
rect 4767 5156 4793 5163
rect 4816 5156 4833 5167
rect 4820 5153 4833 5156
rect 4987 5153 4993 5167
rect 5647 5153 5653 5167
rect 3687 5133 3700 5134
rect 3728 5136 3753 5143
rect 3847 5133 3853 5147
rect 4007 5133 4013 5147
rect 4067 5136 4093 5143
rect 4120 5143 4132 5147
rect 4116 5133 4132 5143
rect 4168 5133 4173 5147
rect 4227 5133 4233 5147
rect 4307 5136 4353 5143
rect 4467 5136 4533 5143
rect 2407 5116 2483 5123
rect 2607 5116 2733 5123
rect 3247 5116 3353 5123
rect 3447 5116 3613 5123
rect 807 5096 1103 5103
rect 1467 5096 1573 5103
rect 1727 5096 2133 5103
rect 2316 5103 2323 5113
rect 3707 5116 3893 5123
rect 4047 5113 4053 5127
rect 4116 5123 4123 5133
rect 4076 5116 4123 5123
rect 2316 5096 2493 5103
rect 3953 5103 3967 5113
rect 4076 5103 4083 5116
rect 4367 5116 4433 5123
rect 4573 5123 4587 5133
rect 4507 5120 4587 5123
rect 4667 5136 4693 5143
rect 4613 5123 4627 5133
rect 4733 5123 4747 5133
rect 4613 5120 4747 5123
rect 4907 5133 4913 5147
rect 4853 5127 4867 5133
rect 4853 5120 4873 5127
rect 4507 5116 4583 5120
rect 4616 5116 4743 5120
rect 4856 5116 4873 5120
rect 4860 5113 4873 5116
rect 4973 5123 4987 5133
rect 4887 5120 4987 5123
rect 5013 5127 5027 5133
rect 4887 5116 4983 5120
rect 5507 5116 5533 5123
rect 5593 5107 5607 5113
rect 3647 5100 3967 5103
rect 3647 5096 3963 5100
rect 3996 5096 4083 5103
rect 3996 5087 4003 5096
rect 4107 5096 4153 5103
rect 4267 5096 4393 5103
rect 4607 5096 4733 5103
rect 4747 5096 4773 5103
rect 5007 5096 5053 5103
rect 107 5076 233 5083
rect 687 5076 773 5083
rect 1847 5076 1913 5083
rect 1927 5076 2273 5083
rect 3367 5076 3453 5083
rect 3687 5076 3992 5083
rect 4028 5076 4483 5083
rect 427 5056 1293 5063
rect 2827 5056 3133 5063
rect 3827 5056 3893 5063
rect 3907 5056 4193 5063
rect 4287 5056 4433 5063
rect 4476 5063 4483 5076
rect 4807 5076 5013 5083
rect 5427 5076 5593 5083
rect 4476 5056 4793 5063
rect 4867 5056 5153 5063
rect 747 5036 853 5043
rect 867 5036 1393 5043
rect 2787 5036 3433 5043
rect 3947 5036 4233 5043
rect 4727 5036 4833 5043
rect 4856 5036 5093 5043
rect 167 5016 193 5023
rect 587 5016 613 5023
rect 1187 5013 1193 5027
rect 2547 5016 2653 5023
rect 2807 5016 2893 5023
rect 4027 5016 4293 5023
rect 4407 5016 4513 5023
rect 4596 5016 4633 5023
rect 327 4996 433 5003
rect 1067 4996 1133 5003
rect 1147 4996 1353 5003
rect 1367 5000 1523 5003
rect 1367 4996 1527 5000
rect 1513 4987 1527 4996
rect 2107 4996 2313 5003
rect 2233 4987 2247 4996
rect 2407 4996 2613 5003
rect 3407 4996 3753 5003
rect 4596 5003 4603 5016
rect 4856 5023 4863 5036
rect 5567 5036 5693 5043
rect 4807 5016 4863 5023
rect 5227 5016 5293 5023
rect 4107 4996 4603 5003
rect 4627 4996 4713 5003
rect 5347 4996 5713 5003
rect 3353 4987 3367 4993
rect 3953 4987 3967 4993
rect 167 4976 244 4983
rect 256 4980 423 4983
rect 187 4956 213 4963
rect 237 4947 244 4976
rect 253 4976 423 4980
rect 253 4967 267 4976
rect 267 4956 303 4963
rect 47 4936 73 4943
rect 87 4933 93 4947
rect 207 4933 212 4947
rect 296 4943 303 4956
rect 327 4953 332 4967
rect 368 4956 393 4963
rect 416 4963 423 4976
rect 867 4973 873 4987
rect 1087 4976 1173 4983
rect 1187 4976 1213 4983
rect 1227 4976 1333 4983
rect 2047 4976 2133 4983
rect 2627 4976 2693 4983
rect 2807 4980 3264 4983
rect 2807 4976 3267 4980
rect 1713 4967 1727 4973
rect 416 4956 453 4963
rect 507 4953 513 4967
rect 587 4956 633 4963
rect 987 4956 1043 4963
rect 296 4936 333 4943
rect 487 4933 493 4947
rect 547 4933 553 4947
rect 627 4933 633 4947
rect 727 4936 753 4943
rect 907 4936 952 4943
rect 986 4933 987 4940
rect 1008 4933 1013 4947
rect 1036 4943 1043 4956
rect 1247 4956 1353 4963
rect 1393 4947 1407 4953
rect 1036 4936 1113 4943
rect 1167 4936 1273 4943
rect 1493 4947 1507 4953
rect 1836 4960 1903 4963
rect 1836 4956 1907 4960
rect 1533 4947 1547 4953
rect 1647 4936 1713 4943
rect 1836 4943 1843 4956
rect 1893 4947 1907 4956
rect 2027 4956 2093 4963
rect 2187 4956 2212 4963
rect 2248 4953 2252 4967
rect 2288 4956 2372 4963
rect 2406 4953 2407 4960
rect 2473 4963 2487 4973
rect 3253 4967 3267 4976
rect 3516 4980 3593 4983
rect 3473 4967 3487 4973
rect 2428 4956 2652 4963
rect 2688 4953 2692 4967
rect 2728 4956 2773 4963
rect 2907 4956 2952 4963
rect 2988 4953 2993 4967
rect 3227 4953 3232 4967
rect 3253 4960 3254 4967
rect 3407 4956 3433 4963
rect 3513 4976 3593 4980
rect 3513 4967 3527 4976
rect 3847 4976 3893 4983
rect 4137 4980 4172 4983
rect 4133 4976 4172 4980
rect 4133 4967 4147 4976
rect 4208 4976 4233 4983
rect 4347 4976 4392 4983
rect 4406 4973 4407 4980
rect 4428 4976 4473 4983
rect 4526 4973 4527 4980
rect 4548 4976 4573 4983
rect 5336 4983 5343 4993
rect 5307 4976 5343 4983
rect 5516 4980 5553 4983
rect 5513 4976 5553 4980
rect 4393 4967 4407 4973
rect 4513 4967 4527 4973
rect 5153 4967 5167 4973
rect 5513 4967 5527 4976
rect 3536 4956 3813 4963
rect 2393 4947 2407 4953
rect 1767 4936 1843 4943
rect 1916 4936 2013 4943
rect 73 4907 87 4913
rect 187 4916 353 4923
rect 373 4923 387 4933
rect 673 4927 687 4933
rect 973 4927 987 4933
rect 1853 4927 1867 4933
rect 373 4920 593 4923
rect 376 4916 593 4920
rect 673 4920 674 4927
rect 666 4913 667 4920
rect 113 4907 127 4913
rect 653 4907 667 4913
rect 127 4896 513 4903
rect 527 4896 652 4903
rect 666 4900 667 4907
rect 733 4903 747 4913
rect 707 4900 747 4903
rect 1067 4916 1093 4923
rect 1147 4916 1173 4923
rect 773 4903 787 4913
rect 1013 4903 1027 4913
rect 773 4900 1027 4903
rect 1373 4907 1387 4913
rect 707 4896 743 4900
rect 776 4896 1023 4900
rect 1587 4916 1613 4923
rect 1767 4916 1813 4923
rect 1866 4920 1867 4927
rect 1916 4923 1923 4936
rect 2027 4936 2113 4943
rect 2627 4933 2633 4947
rect 2827 4936 2873 4943
rect 2927 4933 2933 4947
rect 2987 4936 3073 4943
rect 3087 4936 3193 4943
rect 3367 4933 3373 4947
rect 3507 4933 3513 4947
rect 3536 4943 3543 4956
rect 3736 4947 3743 4956
rect 3867 4953 3873 4967
rect 3987 4956 4013 4963
rect 4107 4953 4112 4967
rect 4133 4960 4134 4967
rect 4447 4956 4492 4963
rect 4513 4960 4514 4967
rect 4627 4956 4733 4963
rect 4807 4953 4813 4967
rect 5016 4960 5143 4963
rect 3933 4947 3947 4953
rect 4433 4947 4447 4953
rect 3527 4936 3543 4943
rect 3567 4936 3593 4943
rect 3727 4933 3743 4947
rect 3767 4933 3773 4947
rect 1888 4916 1923 4923
rect 2087 4913 2093 4927
rect 2353 4923 2367 4933
rect 2353 4920 2593 4923
rect 2356 4916 2593 4920
rect 2687 4916 2793 4923
rect 2847 4913 2853 4927
rect 1413 4907 1427 4913
rect 1653 4903 1667 4913
rect 1627 4900 1667 4903
rect 1627 4896 1663 4900
rect 1867 4896 1933 4903
rect 2133 4903 2147 4913
rect 3053 4907 3067 4913
rect 2133 4900 2373 4903
rect 2136 4896 2373 4900
rect 2387 4896 2433 4903
rect 3233 4923 3247 4933
rect 3453 4927 3467 4933
rect 3233 4920 3453 4923
rect 3236 4916 3453 4920
rect 3627 4916 3653 4923
rect 3736 4923 3743 4933
rect 4073 4927 4087 4933
rect 3736 4916 3973 4923
rect 4307 4933 4313 4947
rect 4553 4947 4567 4953
rect 4733 4947 4747 4953
rect 4687 4933 4693 4947
rect 4853 4947 4867 4953
rect 5013 4956 5147 4960
rect 5013 4947 5027 4956
rect 5133 4947 5147 4956
rect 5327 4953 5333 4967
rect 5407 4953 5413 4967
rect 5536 4960 5643 4963
rect 5533 4956 5647 4960
rect 5193 4947 5207 4953
rect 5533 4947 5547 4956
rect 5193 4940 5194 4947
rect 5186 4933 5187 4940
rect 5208 4936 5273 4943
rect 5447 4936 5472 4943
rect 5493 4933 5494 4940
rect 5633 4947 5647 4956
rect 4113 4923 4127 4933
rect 4113 4920 4233 4923
rect 4116 4916 4233 4920
rect 4647 4913 4653 4927
rect 4967 4916 4993 4923
rect 5173 4923 5187 4933
rect 5493 4927 5507 4933
rect 5047 4916 5393 4923
rect 5493 4920 5494 4927
rect 5607 4913 5613 4927
rect 3093 4907 3107 4913
rect 3573 4903 3587 4913
rect 3487 4900 3587 4903
rect 3487 4896 3583 4900
rect 3787 4896 3993 4903
rect 4127 4896 4173 4903
rect 4407 4896 4433 4903
rect 4487 4896 4613 4903
rect 207 4876 313 4883
rect 327 4876 713 4883
rect 1027 4876 1153 4883
rect 1507 4876 2233 4883
rect 2247 4876 3033 4883
rect 3767 4876 4153 4883
rect 4267 4876 4553 4883
rect 4696 4883 4703 4913
rect 5507 4896 5613 4903
rect 5653 4903 5667 4913
rect 5627 4900 5667 4903
rect 5627 4896 5663 4900
rect 5053 4887 5067 4893
rect 4567 4876 4703 4883
rect 5047 4880 5067 4887
rect 5047 4876 5063 4880
rect 5047 4873 5060 4876
rect 5107 4876 5593 4883
rect 5607 4876 5633 4883
rect 56 4856 153 4863
rect 56 4827 63 4856
rect 407 4856 433 4863
rect 447 4853 453 4867
rect 587 4856 693 4863
rect 2187 4856 2473 4863
rect 2487 4856 2793 4863
rect 2887 4856 2993 4863
rect 3007 4856 3153 4863
rect 4027 4853 4032 4867
rect 4068 4856 4473 4863
rect 5147 4856 5373 4863
rect 87 4836 153 4843
rect 167 4836 533 4843
rect 547 4836 673 4843
rect 687 4836 1733 4843
rect 2507 4836 2833 4843
rect 2887 4836 2953 4843
rect 3227 4836 3493 4843
rect 4127 4836 4493 4843
rect 4747 4836 4953 4843
rect 487 4816 613 4823
rect 627 4816 693 4823
rect 1387 4816 1573 4823
rect 2496 4823 2503 4833
rect 5387 4836 5433 4843
rect 5447 4836 5473 4843
rect 1587 4816 2503 4823
rect 2947 4816 3633 4823
rect 3647 4816 3953 4823
rect 4007 4816 4333 4823
rect 4487 4816 4653 4823
rect 4696 4816 5513 4823
rect 1967 4796 2193 4803
rect 2767 4800 2804 4803
rect 2767 4796 2807 4800
rect 2793 4787 2807 4796
rect 2927 4796 3053 4803
rect 3067 4796 3233 4803
rect 3407 4796 3573 4803
rect 3627 4796 3693 4803
rect 4087 4796 4293 4803
rect 4696 4803 4703 4816
rect 4507 4796 4703 4803
rect 4716 4796 4873 4803
rect 667 4776 1453 4783
rect 2607 4776 2653 4783
rect 2707 4776 2772 4783
rect 2793 4780 2794 4787
rect 2847 4776 3213 4783
rect 3807 4776 4093 4783
rect 4167 4776 4273 4783
rect 4716 4783 4723 4796
rect 4587 4776 4723 4783
rect 4747 4776 5033 4783
rect 367 4756 613 4763
rect 627 4756 753 4763
rect 767 4756 833 4763
rect 2687 4756 4013 4763
rect 407 4736 793 4743
rect 807 4736 933 4743
rect 1207 4736 1293 4743
rect 1607 4736 1953 4743
rect 2167 4736 2453 4743
rect 2627 4736 2933 4743
rect 3467 4736 3733 4743
rect 3967 4736 4053 4743
rect 4067 4736 4203 4743
rect 113 4707 127 4713
rect 633 4713 634 4720
rect 1636 4716 1823 4723
rect 1916 4720 2213 4723
rect 633 4707 647 4713
rect 1636 4707 1643 4716
rect 347 4700 503 4703
rect 347 4696 507 4700
rect 493 4687 507 4696
rect 633 4700 634 4707
rect 626 4693 627 4700
rect 648 4696 743 4703
rect 613 4687 627 4693
rect 736 4687 743 4696
rect 767 4693 773 4707
rect 1007 4700 1063 4703
rect 1007 4696 1067 4700
rect 1053 4687 1067 4696
rect 1187 4693 1193 4707
rect 1247 4693 1253 4707
rect 1267 4696 1313 4703
rect 1467 4696 1553 4703
rect 1606 4693 1607 4700
rect 1628 4696 1643 4707
rect 1756 4700 1793 4703
rect 1753 4696 1793 4700
rect 1628 4693 1640 4696
rect 1593 4687 1607 4693
rect 1753 4687 1767 4696
rect 1816 4703 1823 4716
rect 1913 4716 2213 4720
rect 1913 4707 1927 4716
rect 2013 4707 2027 4716
rect 2887 4716 3013 4723
rect 3207 4716 3253 4723
rect 3387 4716 3773 4723
rect 3856 4720 3933 4723
rect 3853 4716 3933 4720
rect 3293 4707 3307 4713
rect 3853 4707 3867 4716
rect 4196 4707 4203 4736
rect 1816 4696 1853 4703
rect 2026 4700 2027 4707
rect 2033 4693 2034 4700
rect 2536 4696 2573 4703
rect 2033 4687 2047 4693
rect 2536 4687 2543 4696
rect 2613 4687 2627 4693
rect 2756 4696 2873 4703
rect 67 4676 93 4683
rect 147 4673 153 4687
rect 228 4673 233 4687
rect 367 4673 372 4687
rect 408 4673 413 4687
rect 547 4673 553 4687
rect 736 4676 753 4687
rect 740 4673 753 4676
rect 767 4676 783 4683
rect 93 4667 107 4673
rect 195 4643 202 4673
rect 653 4667 667 4673
rect 287 4656 333 4663
rect 467 4653 473 4667
rect 776 4663 783 4676
rect 807 4673 812 4687
rect 848 4676 893 4683
rect 947 4673 953 4687
rect 1107 4673 1113 4687
rect 1200 4686 1213 4687
rect 1207 4673 1213 4686
rect 1287 4673 1293 4687
rect 1333 4667 1347 4673
rect 1476 4676 1523 4683
rect 776 4656 912 4663
rect 47 4636 202 4643
rect 216 4623 223 4653
rect 373 4647 387 4653
rect 513 4647 527 4653
rect 948 4656 1033 4663
rect 1407 4656 1453 4663
rect 1476 4663 1483 4676
rect 1467 4656 1483 4663
rect 1516 4663 1523 4676
rect 1647 4673 1653 4687
rect 1907 4673 1912 4687
rect 1948 4676 2033 4683
rect 2127 4673 2133 4687
rect 2407 4673 2413 4687
rect 2527 4673 2533 4687
rect 2613 4680 2614 4687
rect 2606 4673 2607 4680
rect 2667 4676 2713 4683
rect 2727 4673 2733 4687
rect 1713 4667 1727 4673
rect 2073 4667 2087 4673
rect 2353 4667 2367 4673
rect 1516 4656 1692 4663
rect 1726 4660 1727 4667
rect 1748 4653 1752 4667
rect 1788 4656 1992 4663
rect 2028 4656 2052 4663
rect 2073 4660 2074 4667
rect 2216 4656 2332 4663
rect 1073 4643 1087 4653
rect 1493 4647 1507 4653
rect 1073 4640 1333 4643
rect 1076 4636 1333 4640
rect 1493 4640 1494 4647
rect 1486 4633 1487 4640
rect 1508 4636 1713 4643
rect 1867 4636 2113 4643
rect 2127 4633 2133 4647
rect 2216 4643 2223 4656
rect 2366 4660 2367 4667
rect 2388 4653 2393 4667
rect 2447 4656 2493 4663
rect 2593 4663 2607 4673
rect 2756 4667 2763 4696
rect 2927 4696 2973 4703
rect 3127 4696 3173 4703
rect 3227 4693 3233 4707
rect 3306 4700 3307 4707
rect 3328 4696 3353 4703
rect 3407 4693 3413 4707
rect 3787 4696 3813 4703
rect 4147 4693 4153 4707
rect 4507 4693 4513 4707
rect 4567 4693 4573 4707
rect 4967 4693 4973 4707
rect 5027 4696 5073 4703
rect 5087 4696 5143 4703
rect 2787 4674 2793 4687
rect 2787 4673 2800 4674
rect 2907 4673 2913 4687
rect 3067 4676 3093 4683
rect 3167 4676 3213 4683
rect 3387 4676 3433 4683
rect 3507 4673 3513 4687
rect 3607 4673 3613 4687
rect 3627 4680 3683 4683
rect 3627 4676 3687 4680
rect 2507 4656 2583 4663
rect 2593 4660 2653 4663
rect 2596 4656 2653 4660
rect 2147 4636 2223 4643
rect 2356 4643 2363 4653
rect 2247 4636 2363 4643
rect 2576 4643 2583 4656
rect 2667 4656 2713 4663
rect 2807 4653 2813 4667
rect 2987 4653 2993 4667
rect 3096 4663 3103 4673
rect 3253 4663 3267 4673
rect 3673 4667 3687 4676
rect 3827 4673 3833 4687
rect 3960 4683 3973 4687
rect 3957 4680 3973 4683
rect 3953 4673 3973 4680
rect 4076 4680 4093 4683
rect 4073 4676 4093 4680
rect 3953 4667 3967 4673
rect 4073 4667 4087 4676
rect 4107 4676 4173 4683
rect 4547 4673 4553 4687
rect 4647 4673 4653 4687
rect 5007 4676 5113 4683
rect 5136 4683 5143 4696
rect 5136 4676 5153 4683
rect 5167 4676 5223 4683
rect 4313 4667 4327 4673
rect 4833 4667 4847 4673
rect 5216 4667 5223 4676
rect 5387 4673 5393 4687
rect 5495 4680 5553 4683
rect 5493 4676 5553 4680
rect 5493 4667 5507 4676
rect 3096 4660 3267 4663
rect 3096 4656 3263 4660
rect 3467 4653 3473 4667
rect 3727 4653 3733 4667
rect 3787 4656 3912 4663
rect 3953 4660 3954 4667
rect 3946 4653 3947 4660
rect 4007 4656 4033 4663
rect 4187 4656 4233 4663
rect 4447 4653 4453 4667
rect 4707 4653 4713 4667
rect 4907 4656 5133 4663
rect 5187 4653 5193 4667
rect 5216 4656 5233 4667
rect 5220 4653 5233 4656
rect 5287 4653 5293 4667
rect 5506 4660 5507 4667
rect 5528 4653 5533 4667
rect 5627 4653 5633 4667
rect 3933 4647 3947 4653
rect 4353 4647 4367 4653
rect 4793 4647 4807 4653
rect 2576 4636 2913 4643
rect 2987 4636 3013 4643
rect 3147 4633 3153 4647
rect 3227 4636 3413 4643
rect 3567 4633 3573 4647
rect 3596 4636 3693 4643
rect 87 4616 223 4623
rect 347 4616 413 4623
rect 567 4616 653 4623
rect 1473 4623 1487 4633
rect 1473 4620 1633 4623
rect 1476 4616 1633 4620
rect 1767 4616 2693 4623
rect 3596 4623 3603 4636
rect 3707 4636 3773 4643
rect 3946 4640 3947 4647
rect 4047 4633 4053 4647
rect 4487 4636 4613 4643
rect 4627 4633 4633 4647
rect 5107 4636 5253 4643
rect 5407 4636 5433 4643
rect 5393 4627 5407 4633
rect 3447 4616 3603 4623
rect 3667 4616 3793 4623
rect 4507 4616 4693 4623
rect 5187 4616 5313 4623
rect 627 4596 713 4603
rect 727 4596 753 4603
rect 867 4596 973 4603
rect 987 4596 1093 4603
rect 1107 4596 1233 4603
rect 1407 4596 1653 4603
rect 1907 4596 2073 4603
rect 2087 4596 2413 4603
rect 2887 4596 2933 4603
rect 3907 4596 3993 4603
rect 4547 4596 4623 4603
rect 1627 4576 1693 4583
rect 2307 4576 3373 4583
rect 4207 4576 4293 4583
rect 4367 4576 4593 4583
rect 4616 4583 4623 4596
rect 4787 4596 4833 4603
rect 5347 4596 5423 4603
rect 4616 4576 5173 4583
rect 5416 4583 5423 4596
rect 5416 4576 5513 4583
rect 527 4556 993 4563
rect 1647 4556 1753 4563
rect 2367 4556 2753 4563
rect 2987 4556 3313 4563
rect 3327 4556 3573 4563
rect 4047 4556 4533 4563
rect 4687 4556 4733 4563
rect 4807 4556 5113 4563
rect 5127 4556 5333 4563
rect 5387 4556 5553 4563
rect 107 4536 173 4543
rect 727 4536 933 4543
rect 1087 4536 1333 4543
rect 1547 4536 1733 4543
rect 1927 4536 2153 4543
rect 2347 4536 2433 4543
rect 3576 4543 3583 4553
rect 2927 4536 3563 4543
rect 3576 4536 4133 4543
rect 247 4516 283 4523
rect 276 4503 283 4516
rect 387 4516 593 4523
rect 1007 4516 1133 4523
rect 2067 4516 2613 4523
rect 2707 4516 2733 4523
rect 2747 4516 2973 4523
rect 3087 4516 3133 4523
rect 3556 4523 3563 4536
rect 4147 4536 4533 4543
rect 4707 4536 4753 4543
rect 3367 4520 3523 4523
rect 3367 4516 3527 4520
rect 3556 4516 3673 4523
rect 3513 4507 3527 4516
rect 3967 4516 4253 4523
rect 4296 4516 4433 4523
rect 276 4496 373 4503
rect 667 4496 853 4503
rect 867 4496 1073 4503
rect 1227 4496 1273 4503
rect 1507 4496 1553 4503
rect 1667 4496 2433 4503
rect 2926 4493 2927 4500
rect 2948 4496 2993 4503
rect 3016 4496 3033 4503
rect 133 4487 147 4493
rect 87 4473 93 4487
rect 267 4474 273 4487
rect 267 4473 280 4474
rect 353 4467 367 4473
rect 47 4456 73 4463
rect 127 4456 212 4463
rect 233 4453 234 4460
rect 287 4453 293 4467
rect 393 4467 407 4473
rect 493 4467 507 4473
rect 613 4467 627 4473
rect 653 4467 667 4473
rect 713 4467 727 4473
rect 753 4467 767 4473
rect 993 4467 1007 4473
rect 1133 4467 1147 4473
rect 1347 4476 1453 4483
rect 1747 4473 1753 4487
rect 1807 4473 1813 4487
rect 1866 4473 1867 4480
rect 1888 4476 2003 4483
rect 2036 4480 2113 4483
rect 1273 4467 1287 4473
rect 1853 4467 1867 4473
rect 1996 4467 2003 4476
rect 2033 4476 2113 4480
rect 2033 4467 2047 4476
rect 907 4456 933 4463
rect 947 4453 953 4467
rect 1087 4453 1093 4467
rect 1227 4453 1233 4467
rect 1407 4456 1472 4463
rect 1493 4453 1494 4460
rect 1627 4453 1632 4467
rect 1653 4453 1654 4460
rect 1707 4453 1713 4467
rect 1907 4453 1913 4467
rect 2167 4476 2253 4483
rect 2307 4473 2313 4487
rect 2913 4487 2927 4493
rect 2527 4476 2553 4483
rect 2567 4476 2593 4483
rect 2687 4473 2692 4487
rect 2728 4473 2733 4487
rect 3016 4483 3023 4496
rect 3047 4496 3333 4503
rect 3527 4496 3653 4503
rect 3987 4496 4173 4503
rect 4296 4503 4303 4516
rect 4847 4516 4973 4523
rect 5067 4516 5213 4523
rect 4227 4496 4303 4503
rect 4313 4493 4314 4500
rect 4976 4500 5153 4503
rect 4973 4496 5153 4500
rect 4313 4487 4327 4493
rect 4973 4487 4987 4496
rect 2967 4476 3023 4483
rect 3047 4473 3053 4487
rect 3107 4476 3212 4483
rect 3248 4473 3253 4487
rect 3327 4476 3373 4483
rect 3427 4476 3533 4483
rect 3547 4476 3653 4483
rect 3667 4473 3672 4487
rect 3708 4473 3713 4487
rect 3836 4480 3893 4483
rect 3833 4476 3893 4480
rect 2113 4467 2127 4473
rect 2633 4467 2647 4473
rect 3833 4467 3847 4476
rect 3947 4473 3952 4487
rect 3988 4476 4033 4483
rect 4047 4473 4053 4487
rect 4127 4476 4292 4483
rect 4313 4480 4314 4487
rect 4367 4476 4612 4483
rect 4633 4473 4634 4480
rect 4707 4473 4712 4487
rect 4748 4473 4753 4487
rect 4887 4476 4933 4483
rect 4996 4476 5083 4483
rect 4633 4467 4647 4473
rect 2246 4453 2247 4460
rect 2268 4453 2273 4467
rect 2407 4453 2413 4467
rect 2527 4453 2533 4467
rect 2646 4460 2647 4467
rect 2653 4453 2654 4460
rect 2787 4453 2793 4467
rect 3166 4453 3167 4460
rect 3188 4453 3193 4467
rect 3247 4456 3273 4463
rect 3347 4456 3393 4463
rect 3447 4453 3453 4467
rect 3567 4453 3573 4467
rect 3667 4453 3673 4467
rect 3727 4456 3793 4463
rect 4207 4456 4292 4463
rect 4328 4453 4333 4467
rect 4587 4453 4593 4467
rect 4616 4456 4633 4463
rect 233 4447 247 4453
rect 233 4443 234 4447
rect 147 4436 234 4443
rect 367 4436 433 4443
rect 447 4436 473 4443
rect 607 4436 633 4443
rect 647 4436 733 4443
rect 987 4433 993 4447
rect 1007 4436 1113 4443
rect 1167 4433 1173 4447
rect 1187 4436 1253 4443
rect 1387 4433 1392 4447
rect 1428 4436 1453 4443
rect 1493 4443 1507 4453
rect 1653 4447 1667 4453
rect 1993 4447 2007 4453
rect 2233 4447 2247 4453
rect 1467 4440 1507 4443
rect 1467 4436 1503 4440
rect 1947 4433 1953 4447
rect 2006 4440 2007 4447
rect 2013 4433 2014 4440
rect 2246 4440 2247 4447
rect 2427 4436 2453 4443
rect 2536 4443 2543 4453
rect 2653 4443 2667 4453
rect 2536 4440 2667 4443
rect 2693 4447 2707 4453
rect 3153 4447 3167 4453
rect 2536 4436 2664 4440
rect 2747 4436 2773 4443
rect 2827 4433 2833 4447
rect 3207 4436 3233 4443
rect 3393 4443 3407 4453
rect 3393 4440 3513 4443
rect 3396 4436 3513 4440
rect 3827 4433 3832 4447
rect 3853 4433 3854 4440
rect 4127 4436 4173 4443
rect 4616 4443 4623 4456
rect 4996 4463 5003 4476
rect 5076 4467 5083 4476
rect 5167 4473 5172 4487
rect 5208 4473 5213 4487
rect 5327 4473 5333 4487
rect 5487 4476 5513 4483
rect 5567 4473 5573 4487
rect 5253 4467 5267 4473
rect 4967 4456 5003 4463
rect 5047 4453 5052 4467
rect 5073 4453 5074 4460
rect 5373 4467 5387 4473
rect 5467 4456 5533 4463
rect 4913 4447 4927 4453
rect 5073 4447 5087 4453
rect 4547 4436 4623 4443
rect 4727 4436 4753 4443
rect 5027 4433 5033 4447
rect 5573 4443 5587 4453
rect 5487 4440 5587 4443
rect 5487 4436 5583 4440
rect 513 4427 527 4433
rect 267 4416 492 4423
rect 513 4420 514 4427
rect 647 4416 693 4423
rect 1613 4423 1627 4433
rect 1467 4420 1627 4423
rect 1467 4416 1623 4420
rect 2013 4423 2027 4433
rect 2093 4423 2107 4433
rect 1947 4420 2027 4423
rect 2036 4420 2107 4423
rect 1947 4416 2024 4420
rect 2036 4416 2103 4420
rect 827 4396 1073 4403
rect 2036 4403 2043 4416
rect 1927 4396 2043 4403
rect 2136 4403 2143 4433
rect 2373 4427 2387 4433
rect 2567 4416 2593 4423
rect 2736 4423 2743 4433
rect 2647 4416 3233 4423
rect 3853 4423 3867 4433
rect 3247 4416 3933 4423
rect 4213 4423 4227 4433
rect 4007 4420 4227 4423
rect 4007 4416 4223 4420
rect 4447 4416 4593 4423
rect 4927 4416 5033 4423
rect 5447 4416 5613 4423
rect 2067 4396 2143 4403
rect 2247 4396 2413 4403
rect 2707 4396 2833 4403
rect 3167 4396 3273 4403
rect 3427 4396 3833 4403
rect 3927 4396 4053 4403
rect 4067 4396 4393 4403
rect 2027 4376 2233 4383
rect 2307 4376 2333 4383
rect 2527 4376 3093 4383
rect 4347 4376 4393 4383
rect 4447 4376 4473 4383
rect 567 4356 973 4363
rect 1067 4356 1133 4363
rect 1927 4356 2633 4363
rect 2647 4356 2673 4363
rect 2687 4356 2873 4363
rect 3667 4356 3793 4363
rect 3996 4356 4493 4363
rect 1947 4336 2253 4343
rect 2427 4336 3053 4343
rect 3996 4343 4003 4356
rect 4587 4356 4693 4363
rect 4707 4356 4793 4363
rect 5427 4356 5653 4363
rect 3656 4336 4003 4343
rect 487 4316 733 4323
rect 1587 4316 2513 4323
rect 3656 4323 3663 4336
rect 4027 4336 4673 4343
rect 4716 4336 5013 4343
rect 2967 4316 3663 4323
rect 3687 4316 3753 4323
rect 4387 4316 4553 4323
rect 4716 4323 4723 4336
rect 5027 4336 5073 4343
rect 4647 4316 4723 4323
rect 4747 4316 4873 4323
rect 5047 4316 5273 4323
rect 287 4296 573 4303
rect 587 4296 1113 4303
rect 1707 4296 2073 4303
rect 2387 4303 2400 4307
rect 2387 4293 2403 4303
rect 2707 4296 2733 4303
rect 3067 4296 5253 4303
rect 5267 4296 5593 4303
rect 2396 4287 2403 4293
rect 407 4276 513 4283
rect 527 4276 613 4283
rect 627 4276 1533 4283
rect 2407 4276 3093 4283
rect 3247 4276 3413 4283
rect 3507 4276 4053 4283
rect 267 4256 853 4263
rect 1627 4256 1753 4263
rect 1847 4256 2153 4263
rect 2167 4256 2373 4263
rect 2847 4256 3153 4263
rect 3167 4256 4173 4263
rect 5227 4256 5373 4263
rect 107 4236 253 4243
rect 253 4227 267 4233
rect 187 4213 193 4227
rect 487 4240 523 4243
rect 487 4236 527 4240
rect 353 4227 367 4233
rect 513 4227 527 4236
rect 647 4236 673 4243
rect 896 4240 983 4243
rect 1215 4240 1373 4243
rect 893 4236 983 4240
rect 447 4213 453 4227
rect 893 4227 907 4236
rect 816 4220 893 4223
rect 813 4216 893 4220
rect 93 4207 107 4213
rect 393 4207 407 4213
rect 813 4207 827 4216
rect 976 4223 983 4236
rect 1213 4236 1373 4240
rect 1213 4227 1227 4236
rect 2247 4236 2413 4243
rect 2567 4236 2823 4243
rect 2033 4227 2047 4233
rect 976 4216 1153 4223
rect 933 4207 947 4213
rect 1053 4207 1067 4216
rect 1226 4220 1227 4227
rect 1248 4216 1633 4223
rect 1707 4216 1733 4223
rect 1787 4213 1792 4227
rect 1828 4213 1833 4227
rect 2127 4216 2303 4223
rect 2073 4207 2087 4213
rect 2296 4207 2303 4216
rect 2313 4213 2314 4220
rect 2633 4213 2634 4220
rect 2313 4207 2327 4213
rect 2633 4207 2647 4213
rect 147 4193 153 4207
rect 247 4203 260 4207
rect 247 4193 263 4203
rect 287 4193 293 4207
rect 316 4196 372 4203
rect 87 4176 213 4183
rect 256 4183 263 4193
rect 316 4183 323 4196
rect 393 4200 394 4207
rect 547 4196 613 4203
rect 627 4193 632 4207
rect 668 4196 713 4203
rect 867 4196 912 4203
rect 933 4200 934 4207
rect 1187 4193 1193 4207
rect 1247 4196 1293 4203
rect 1367 4196 1463 4203
rect 256 4176 323 4183
rect 493 4183 507 4193
rect 773 4187 787 4193
rect 493 4180 573 4183
rect 496 4176 573 4180
rect 126 4153 127 4160
rect 256 4163 263 4176
rect 647 4173 652 4187
rect 688 4173 693 4187
rect 747 4173 752 4187
rect 786 4180 787 4187
rect 808 4173 812 4187
rect 848 4176 933 4183
rect 947 4176 1013 4183
rect 1027 4176 1233 4183
rect 1456 4183 1463 4196
rect 1507 4193 1513 4207
rect 1567 4193 1573 4207
rect 1687 4193 1692 4207
rect 1713 4193 1714 4200
rect 1787 4193 1792 4207
rect 1828 4196 1893 4203
rect 1907 4193 1912 4207
rect 1948 4193 1953 4207
rect 2007 4196 2052 4203
rect 2073 4200 2074 4207
rect 2167 4193 2173 4207
rect 2227 4193 2233 4207
rect 2313 4200 2314 4207
rect 2306 4193 2307 4200
rect 2367 4196 2393 4203
rect 2487 4196 2573 4203
rect 2587 4193 2593 4207
rect 2633 4200 2634 4207
rect 2727 4196 2753 4203
rect 2816 4203 2823 4236
rect 3027 4236 3333 4243
rect 3136 4227 3143 4236
rect 3447 4236 3593 4243
rect 2947 4216 3013 4223
rect 3067 4216 3133 4223
rect 3207 4220 3324 4223
rect 3207 4216 3327 4220
rect 3313 4207 3327 4216
rect 3753 4227 3767 4233
rect 4647 4236 4793 4243
rect 5147 4236 5253 4243
rect 4253 4227 4267 4233
rect 5373 4227 5387 4233
rect 3587 4216 3653 4223
rect 3807 4213 3813 4227
rect 3867 4216 3893 4223
rect 3947 4213 3953 4227
rect 3967 4216 4113 4223
rect 4187 4216 4213 4223
rect 4307 4220 4402 4223
rect 4307 4216 4407 4220
rect 3413 4207 3427 4213
rect 2816 4200 2953 4203
rect 1456 4176 1533 4183
rect 1587 4173 1593 4187
rect 1713 4183 1727 4193
rect 2293 4187 2307 4193
rect 2793 4187 2807 4193
rect 1607 4180 1727 4183
rect 1607 4176 1724 4180
rect 1747 4176 1933 4183
rect 1987 4176 2112 4183
rect 2148 4176 2193 4183
rect 2247 4173 2253 4187
rect 2387 4176 2433 4183
rect 2527 4176 2553 4183
rect 2567 4173 2573 4187
rect 2600 4183 2613 4187
rect 2596 4173 2613 4183
rect 2667 4173 2672 4187
rect 2708 4176 2732 4183
rect 2768 4173 2772 4187
rect 2806 4180 2807 4187
rect 2813 4196 2953 4200
rect 2813 4187 2827 4196
rect 3007 4196 3033 4203
rect 3167 4193 3173 4207
rect 3267 4193 3272 4207
rect 3293 4193 3294 4200
rect 3313 4200 3314 4207
rect 3467 4196 3533 4203
rect 3293 4187 3307 4193
rect 3587 4196 3673 4203
rect 3693 4203 3707 4213
rect 4393 4207 4407 4216
rect 5307 4216 5333 4223
rect 5387 4216 5453 4223
rect 5467 4213 5473 4227
rect 5213 4207 5227 4213
rect 5513 4207 5527 4213
rect 3693 4200 3773 4203
rect 3696 4196 3773 4200
rect 4007 4193 4013 4207
rect 4366 4193 4367 4200
rect 4386 4193 4387 4200
rect 4406 4200 4407 4207
rect 4413 4193 4414 4200
rect 4567 4193 4573 4207
rect 5267 4196 5353 4203
rect 5487 4193 5492 4207
rect 5513 4200 5514 4207
rect 5567 4196 5593 4203
rect 5647 4193 5653 4207
rect 3913 4187 3927 4193
rect 2813 4180 2814 4187
rect 3207 4176 3233 4183
rect 3293 4180 3294 4187
rect 3387 4173 3392 4187
rect 3428 4173 3433 4187
rect 4107 4173 4113 4187
rect 4233 4183 4247 4193
rect 4353 4183 4367 4193
rect 4233 4180 4367 4183
rect 4373 4187 4387 4193
rect 4236 4176 4362 4180
rect 4413 4187 4427 4193
rect 4527 4173 4533 4187
rect 4687 4176 4712 4183
rect 4748 4176 4773 4183
rect 148 4156 263 4163
rect 1347 4153 1353 4167
rect 1447 4156 1573 4163
rect 1627 4156 1813 4163
rect 2256 4163 2263 4173
rect 2256 4156 2313 4163
rect 2333 4163 2347 4173
rect 2333 4160 2413 4163
rect 2336 4156 2413 4160
rect 2596 4163 2603 4173
rect 3333 4167 3347 4173
rect 3573 4167 3587 4173
rect 2527 4156 2603 4163
rect 2627 4156 2713 4163
rect 2887 4153 2893 4167
rect 3067 4156 3233 4163
rect 3507 4156 3573 4163
rect 3587 4156 3613 4163
rect 3927 4156 3993 4163
rect 4116 4163 4123 4173
rect 4453 4163 4467 4173
rect 4116 4160 4467 4163
rect 4873 4167 4887 4173
rect 4116 4156 4463 4160
rect 5007 4173 5012 4187
rect 5048 4176 5073 4183
rect 5147 4173 5152 4187
rect 5188 4173 5193 4187
rect 4913 4167 4927 4173
rect 5233 4167 5247 4173
rect 5573 4167 5587 4173
rect 5447 4156 5493 4163
rect 5613 4167 5627 4173
rect 5613 4160 5633 4167
rect 5616 4156 5633 4160
rect 5620 4153 5633 4156
rect 113 4143 127 4153
rect 113 4140 273 4143
rect 115 4136 273 4140
rect 647 4136 773 4143
rect 787 4136 873 4143
rect 1620 4146 1633 4147
rect 533 4123 547 4133
rect 1627 4133 1633 4146
rect 1687 4136 2133 4143
rect 2367 4136 2493 4143
rect 2567 4136 2693 4143
rect 3307 4136 3373 4143
rect 3887 4136 4013 4143
rect 4067 4136 4093 4143
rect 5407 4136 5533 4143
rect 533 4120 573 4123
rect 536 4116 573 4120
rect 727 4113 733 4127
rect 1187 4116 1513 4123
rect 1527 4116 1773 4123
rect 2147 4116 2233 4123
rect 2247 4116 2473 4123
rect 2487 4116 2953 4123
rect 3827 4116 4193 4123
rect 4347 4116 4393 4123
rect 287 4096 593 4103
rect 1367 4096 1593 4103
rect 1607 4096 1993 4103
rect 2087 4096 2113 4103
rect 2547 4096 2593 4103
rect 3247 4096 3413 4103
rect 3907 4096 4073 4103
rect 4167 4096 4193 4103
rect 4416 4103 4423 4133
rect 5467 4116 5613 4123
rect 4416 4096 4853 4103
rect 347 4076 533 4083
rect 2067 4076 2293 4083
rect 2447 4076 2613 4083
rect 2987 4076 3193 4083
rect 3207 4076 3713 4083
rect 4747 4076 5033 4083
rect 127 4056 353 4063
rect 367 4056 453 4063
rect 707 4056 853 4063
rect 1327 4056 1973 4063
rect 2107 4056 2253 4063
rect 2267 4056 2653 4063
rect 2667 4056 2793 4063
rect 3347 4056 3413 4063
rect 4307 4056 4533 4063
rect 4547 4056 4753 4063
rect 4767 4056 4913 4063
rect 4987 4056 5153 4063
rect 5227 4056 5632 4063
rect 5668 4053 5673 4067
rect 187 4036 333 4043
rect 407 4036 693 4043
rect 747 4043 760 4047
rect 747 4040 763 4043
rect 747 4033 767 4040
rect 1627 4034 1633 4047
rect 1627 4033 1640 4034
rect 2087 4036 2203 4043
rect 753 4027 767 4033
rect 127 4020 224 4023
rect 127 4016 227 4020
rect 213 4007 227 4016
rect 1147 4016 1233 4023
rect 1640 4026 1653 4027
rect 1387 4020 1522 4023
rect 1387 4016 1527 4020
rect 1513 4007 1527 4016
rect 1647 4013 1653 4026
rect 2196 4023 2203 4036
rect 2227 4036 2493 4043
rect 2996 4036 3273 4043
rect 2996 4027 3003 4036
rect 4507 4036 4553 4043
rect 4627 4036 4733 4043
rect 4807 4036 5073 4043
rect 2196 4016 2253 4023
rect 2267 4016 2473 4023
rect 2847 4016 2943 4023
rect 2173 4007 2187 4013
rect 96 4000 192 4003
rect 93 3996 192 4000
rect 93 3987 107 3996
rect 213 4000 214 4007
rect 287 3996 463 4003
rect 147 3976 173 3983
rect 187 3973 193 3987
rect 327 3973 333 3987
rect 387 3983 400 3987
rect 456 3983 463 3996
rect 487 3993 492 4007
rect 528 3993 533 4007
rect 607 4000 643 4003
rect 607 3996 647 4000
rect 633 3987 647 3996
rect 707 3996 733 4003
rect 387 3973 403 3983
rect 456 3976 493 3983
rect 633 3980 634 3987
rect 626 3973 627 3980
rect 773 3983 787 3993
rect 696 3980 787 3983
rect 1087 3996 1253 4003
rect 1327 3996 1353 4003
rect 1427 3993 1433 4007
rect 1526 4000 1527 4007
rect 1548 3993 1552 4007
rect 1588 3996 1683 4003
rect 873 3987 887 3993
rect 696 3976 783 3980
rect 67 3953 73 3967
rect 113 3947 127 3953
rect 236 3943 243 3973
rect 367 3953 373 3967
rect 396 3943 403 3973
rect 533 3967 547 3973
rect 427 3963 440 3967
rect 427 3953 443 3963
rect 613 3967 627 3973
rect 696 3967 703 3976
rect 927 3976 1013 3983
rect 1076 3983 1083 3993
rect 1076 3976 1103 3983
rect 667 3956 693 3963
rect 867 3966 880 3967
rect 867 3953 872 3966
rect 167 3936 403 3943
rect 436 3943 443 3953
rect 436 3936 533 3943
rect 696 3943 703 3953
rect 893 3953 894 3960
rect 893 3943 907 3953
rect 696 3940 907 3943
rect 993 3947 1007 3953
rect 696 3936 904 3940
rect 1096 3963 1103 3976
rect 1127 3973 1132 3987
rect 1168 3973 1173 3987
rect 1187 3976 1233 3983
rect 1273 3967 1287 3973
rect 1096 3956 1153 3963
rect 1413 3967 1427 3973
rect 1436 3963 1443 3993
rect 1467 3973 1473 3987
rect 1547 3973 1552 3987
rect 1588 3976 1653 3983
rect 1676 3983 1683 3996
rect 1887 3993 1893 4007
rect 1967 3996 2093 4003
rect 2013 3987 2027 3996
rect 2107 3996 2133 4003
rect 2347 3996 2393 4003
rect 2407 3993 2413 4007
rect 2436 3996 2513 4003
rect 1676 3976 1773 3983
rect 2127 3976 2153 3983
rect 2213 3983 2227 3993
rect 2436 3983 2443 3996
rect 2527 3993 2533 4007
rect 2807 3993 2813 4007
rect 2936 4003 2943 4016
rect 2987 4013 2993 4027
rect 3367 4013 3373 4027
rect 3687 4016 3723 4023
rect 3053 4007 3067 4013
rect 3573 4007 3587 4013
rect 3716 4007 3723 4016
rect 3847 4013 3853 4027
rect 4536 4020 4783 4023
rect 4493 4007 4507 4013
rect 2936 3996 2953 4003
rect 2967 3993 2973 4007
rect 2213 3980 2443 3983
rect 2216 3976 2443 3980
rect 2573 3987 2587 3993
rect 3093 3987 3107 3993
rect 3647 4003 3660 4007
rect 3647 3993 3663 4003
rect 3687 3993 3693 4007
rect 3716 3996 3733 4007
rect 3720 3993 3733 3996
rect 3887 3993 3893 4007
rect 3920 4003 3933 4007
rect 3916 3993 3933 4003
rect 3947 3996 3972 4003
rect 4008 3996 4173 4003
rect 4376 4000 4483 4003
rect 4373 3996 4487 4000
rect 3213 3987 3227 3993
rect 2687 3976 2733 3983
rect 2787 3976 2873 3983
rect 2927 3976 3072 3983
rect 3106 3980 3107 3987
rect 3113 3973 3114 3980
rect 3367 3976 3443 3983
rect 1913 3967 1927 3973
rect 1436 3956 1533 3963
rect 1607 3953 1613 3967
rect 1627 3956 1752 3963
rect 1788 3953 1793 3967
rect 2193 3963 2207 3973
rect 1927 3960 2207 3963
rect 1927 3956 2203 3960
rect 2227 3956 2293 3963
rect 2507 3956 2652 3963
rect 2688 3953 2693 3967
rect 2827 3956 3013 3963
rect 3113 3963 3127 3973
rect 3253 3967 3267 3973
rect 3087 3960 3127 3963
rect 3087 3956 3124 3960
rect 3187 3953 3193 3967
rect 3253 3960 3254 3967
rect 3246 3953 3247 3960
rect 3276 3956 3413 3963
rect 1033 3947 1047 3953
rect 1416 3943 1423 3953
rect 1416 3936 1653 3943
rect 1807 3936 1913 3943
rect 3233 3943 3247 3953
rect 3276 3943 3283 3956
rect 3436 3963 3443 3976
rect 3467 3973 3472 3987
rect 3508 3973 3513 3987
rect 3607 3973 3613 3987
rect 3656 3983 3663 3993
rect 3656 3976 3713 3983
rect 3833 3983 3847 3993
rect 3916 3983 3923 3993
rect 4373 3987 4387 3996
rect 3833 3980 3923 3983
rect 3836 3976 3923 3980
rect 3936 3976 3973 3983
rect 3553 3967 3567 3973
rect 3436 3956 3473 3963
rect 3487 3956 3543 3963
rect 3233 3940 3283 3943
rect 3235 3936 3283 3940
rect 3536 3943 3543 3956
rect 3753 3967 3767 3973
rect 3936 3963 3943 3976
rect 4027 3976 4053 3983
rect 4067 3976 4113 3983
rect 4473 3987 4487 3996
rect 4533 4016 4783 4020
rect 4533 4007 4547 4016
rect 4776 4007 4783 4016
rect 4867 4016 5373 4023
rect 5527 4016 5623 4023
rect 4853 4007 4867 4013
rect 5413 4007 5427 4013
rect 5616 4007 5623 4016
rect 4727 3996 4753 4003
rect 4776 3996 4793 4007
rect 4780 3993 4793 3996
rect 4807 3993 4813 4007
rect 4866 4000 4867 4007
rect 4888 3993 4893 4007
rect 5146 3993 5147 4000
rect 5168 3996 5193 4003
rect 5616 3996 5633 4007
rect 5620 3993 5633 3996
rect 5647 3993 5653 4007
rect 5133 3987 5147 3993
rect 5593 3987 5607 3993
rect 4627 3976 4733 3983
rect 4787 3976 4833 3983
rect 4847 3976 4873 3983
rect 4927 3976 5013 3983
rect 5187 3976 5273 3983
rect 5387 3973 5392 3987
rect 5428 3976 5453 3983
rect 4513 3967 4527 3973
rect 5673 3967 5687 3973
rect 3907 3956 3943 3963
rect 4307 3956 4353 3963
rect 4407 3956 4453 3963
rect 4606 3953 4607 3960
rect 4628 3953 4633 3967
rect 4647 3956 4673 3963
rect 4947 3956 4993 3963
rect 5007 3953 5012 3967
rect 5048 3956 5133 3963
rect 5247 3953 5253 3967
rect 3536 3936 3573 3943
rect 2473 3927 2487 3933
rect 3907 3936 3953 3943
rect 4593 3943 4607 3953
rect 4487 3940 4607 3943
rect 4487 3936 4602 3940
rect 5136 3943 5143 3953
rect 5293 3943 5307 3953
rect 4727 3936 5123 3943
rect 5136 3940 5307 3943
rect 5136 3936 5303 3940
rect 207 3916 273 3923
rect 707 3916 853 3923
rect 867 3916 1353 3923
rect 2007 3916 2113 3923
rect 3067 3916 4013 3923
rect 4027 3916 4233 3923
rect 4367 3916 4513 3923
rect 4847 3916 5033 3923
rect 5116 3923 5123 3936
rect 5116 3916 5253 3923
rect 487 3896 913 3903
rect 1087 3896 1393 3903
rect 1527 3896 2093 3903
rect 2467 3896 2693 3903
rect 2887 3896 3912 3903
rect 3948 3896 4373 3903
rect 4387 3896 4712 3903
rect 4748 3896 4853 3903
rect 687 3876 1113 3883
rect 1127 3876 1273 3883
rect 1347 3876 1453 3883
rect 1787 3876 1813 3883
rect 1836 3876 3053 3883
rect 1836 3863 1843 3876
rect 3867 3876 3973 3883
rect 4287 3876 4472 3883
rect 4508 3876 5213 3883
rect 5487 3876 5553 3883
rect 127 3856 1843 3863
rect 2247 3856 3033 3863
rect 3207 3856 3373 3863
rect 3467 3856 3553 3863
rect 3567 3856 3613 3863
rect 3767 3856 3993 3863
rect 4107 3856 5093 3863
rect 5107 3856 5293 3863
rect 1607 3836 1633 3843
rect 1747 3836 1953 3843
rect 2167 3836 2533 3843
rect 2587 3836 2933 3843
rect 2947 3836 3113 3843
rect 3587 3836 3813 3843
rect 4147 3836 4513 3843
rect 4627 3836 4973 3843
rect 5207 3836 5433 3843
rect 207 3816 473 3823
rect 1567 3816 1753 3823
rect 1767 3816 1992 3823
rect 2028 3816 2253 3823
rect 2747 3816 3133 3823
rect 3253 3823 3267 3833
rect 3253 3820 3753 3823
rect 3256 3816 3753 3820
rect 4107 3816 4713 3823
rect 4827 3816 5213 3823
rect 5267 3816 5313 3823
rect 247 3796 353 3803
rect 987 3796 1253 3803
rect 1667 3796 2433 3803
rect 2527 3796 2993 3803
rect 3127 3796 4133 3803
rect 3073 3787 3087 3793
rect 547 3776 853 3783
rect 1047 3776 1153 3783
rect 1167 3776 1593 3783
rect 1867 3776 1973 3783
rect 1987 3776 2072 3783
rect 2108 3773 2113 3787
rect 2667 3776 2853 3783
rect 2867 3776 2953 3783
rect 2967 3776 3013 3783
rect 3067 3780 3087 3787
rect 3067 3776 3083 3780
rect 3067 3773 3080 3776
rect 3107 3776 3253 3783
rect 3427 3776 3653 3783
rect 5107 3776 5193 3783
rect 307 3756 483 3763
rect 476 3747 483 3756
rect 1007 3756 1053 3763
rect 1067 3756 1203 3763
rect 1196 3747 1203 3756
rect 1347 3756 1733 3763
rect 1787 3756 2013 3763
rect 2967 3756 3353 3763
rect 3567 3763 3580 3767
rect 3567 3760 3583 3763
rect 3567 3753 3587 3760
rect 487 3736 813 3743
rect 867 3733 873 3747
rect 887 3736 973 3743
rect 1037 3740 1153 3743
rect 1033 3736 1153 3740
rect 233 3727 247 3733
rect -24 3703 -17 3723
rect 27 3716 153 3723
rect 167 3716 193 3723
rect 287 3716 332 3723
rect 346 3713 347 3720
rect 368 3713 373 3727
rect 387 3716 513 3723
rect 607 3716 713 3723
rect 767 3716 853 3723
rect 867 3713 872 3727
rect 893 3713 894 3720
rect 986 3713 987 3720
rect 1008 3714 1012 3727
rect 1033 3727 1047 3736
rect 1207 3736 1253 3743
rect 1327 3736 1513 3743
rect 1153 3727 1167 3733
rect 1513 3727 1527 3733
rect 1907 3736 2033 3743
rect 2047 3733 2052 3747
rect 2088 3736 2113 3743
rect 2207 3736 2253 3743
rect 2367 3736 2393 3743
rect 2407 3733 2413 3747
rect 2467 3736 2513 3743
rect 2627 3736 2653 3743
rect 2707 3734 2713 3747
rect 3573 3747 3587 3753
rect 3696 3756 3793 3763
rect 2707 3733 2720 3734
rect 2907 3733 2913 3747
rect 3007 3736 3103 3743
rect 1653 3727 1667 3733
rect 1033 3720 1034 3727
rect 1008 3713 1020 3714
rect 333 3707 347 3713
rect -24 3696 53 3703
rect 127 3693 133 3707
rect 187 3696 213 3703
rect 267 3696 292 3703
rect 328 3700 347 3707
rect 328 3696 342 3700
rect 328 3693 340 3696
rect 367 3693 372 3707
rect 480 3706 500 3707
rect 408 3696 473 3703
rect 487 3693 493 3706
rect 587 3696 673 3703
rect 893 3703 907 3713
rect 747 3700 907 3703
rect 973 3707 987 3713
rect 1193 3707 1207 3713
rect 747 3696 904 3700
rect 1013 3693 1014 3700
rect 1067 3693 1073 3707
rect 1347 3716 1393 3723
rect 1567 3713 1573 3727
rect 1707 3716 1773 3723
rect 1896 3723 1903 3733
rect 1836 3720 1903 3723
rect 1833 3716 1903 3720
rect 1293 3707 1307 3713
rect 1833 3707 1847 3716
rect 2047 3713 2053 3727
rect 2427 3713 2433 3727
rect 2456 3716 2533 3723
rect 2193 3707 2207 3713
rect 1467 3696 1533 3703
rect 1556 3696 1573 3703
rect 733 3687 747 3693
rect 1013 3687 1027 3693
rect 527 3673 533 3687
rect 747 3676 992 3683
rect 1013 3680 1014 3687
rect 1556 3683 1563 3696
rect 1587 3696 1652 3703
rect 1673 3693 1674 3700
rect 1727 3696 1753 3703
rect 1907 3693 1913 3707
rect 1967 3693 1973 3707
rect 2127 3696 2153 3703
rect 2247 3696 2313 3703
rect 2456 3703 2463 3716
rect 2687 3716 2713 3723
rect 2736 3716 2793 3723
rect 2367 3696 2463 3703
rect 2736 3703 2743 3716
rect 2807 3713 2812 3727
rect 2848 3713 2853 3727
rect 2947 3713 2953 3727
rect 2976 3716 3032 3723
rect 2667 3696 2743 3703
rect 2767 3693 2773 3707
rect 2976 3703 2983 3716
rect 3066 3713 3067 3720
rect 3053 3707 3067 3713
rect 1447 3676 1563 3683
rect 1673 3683 1687 3693
rect 1607 3680 1687 3683
rect 1607 3676 1683 3680
rect 1787 3676 1813 3683
rect 1853 3667 1867 3673
rect 387 3656 733 3663
rect 887 3656 1093 3663
rect 1307 3656 1753 3663
rect 2047 3676 2113 3683
rect 2207 3676 2333 3683
rect 2407 3676 2473 3683
rect 2547 3676 2593 3683
rect 2813 3683 2827 3693
rect 2916 3696 2983 3703
rect 2916 3687 2923 3696
rect 3007 3693 3013 3707
rect 3066 3700 3067 3707
rect 3073 3713 3074 3720
rect 3096 3723 3103 3736
rect 3147 3740 3323 3743
rect 3147 3736 3327 3740
rect 3313 3727 3327 3736
rect 3096 3716 3133 3723
rect 3427 3740 3563 3743
rect 3427 3736 3567 3740
rect 3353 3727 3367 3733
rect 3553 3727 3567 3736
rect 3627 3734 3633 3747
rect 3620 3733 3633 3734
rect 3696 3743 3703 3756
rect 4987 3760 5163 3763
rect 4987 3756 5167 3760
rect 5153 3747 5167 3756
rect 5607 3756 5713 3763
rect 3647 3736 3703 3743
rect 3727 3733 3733 3747
rect 3927 3733 3933 3747
rect 5107 3733 5113 3747
rect 3853 3727 3867 3733
rect 4173 3727 4187 3733
rect 3607 3726 3620 3727
rect 3607 3713 3613 3726
rect 3073 3707 3087 3713
rect 3667 3716 3693 3723
rect 3747 3713 3753 3727
rect 3807 3716 3832 3723
rect 3866 3720 3867 3727
rect 3873 3713 3874 3720
rect 4007 3713 4013 3727
rect 4127 3713 4133 3727
rect 4587 3713 4593 3727
rect 4987 3714 4993 3727
rect 4980 3713 4993 3714
rect 5047 3716 5133 3723
rect 5227 3716 5253 3723
rect 5627 3716 5693 3723
rect 3073 3700 3074 3707
rect 3093 3693 3094 3700
rect 3147 3696 3172 3703
rect 3208 3693 3213 3707
rect 3227 3696 3293 3703
rect 3347 3696 3413 3703
rect 3507 3696 3713 3703
rect 3873 3703 3887 3713
rect 3807 3700 3887 3703
rect 3807 3696 3884 3700
rect 3927 3696 3973 3703
rect 4047 3693 4053 3707
rect 3093 3687 3107 3693
rect 2727 3676 2913 3683
rect 3107 3676 3193 3683
rect 3453 3683 3467 3693
rect 3287 3680 3467 3683
rect 3287 3676 3463 3680
rect 3487 3676 3553 3683
rect 4113 3683 4127 3693
rect 4227 3693 4233 3707
rect 4307 3693 4313 3707
rect 4467 3693 4473 3707
rect 4547 3693 4553 3707
rect 4707 3693 4713 3707
rect 4787 3693 4792 3707
rect 4828 3693 4833 3707
rect 4967 3693 4972 3707
rect 5008 3693 5013 3707
rect 5307 3693 5313 3707
rect 5387 3693 5392 3707
rect 5428 3693 5433 3707
rect 4153 3687 4167 3693
rect 3836 3676 4143 3683
rect 1933 3663 1947 3673
rect 1933 3660 1993 3663
rect 1936 3656 1993 3660
rect 2196 3663 2203 3673
rect 2067 3656 2203 3663
rect 2247 3656 2373 3663
rect 2596 3656 2733 3663
rect 327 3636 533 3643
rect 576 3636 793 3643
rect 576 3623 583 3636
rect 1407 3636 1913 3643
rect 2596 3643 2603 3656
rect 2827 3656 3073 3663
rect 3836 3663 3843 3676
rect 3487 3656 3843 3663
rect 3867 3656 4033 3663
rect 4136 3663 4143 3676
rect 4353 3687 4367 3693
rect 4907 3676 5093 3683
rect 5507 3676 5573 3683
rect 5587 3676 5673 3683
rect 5233 3667 5247 3673
rect 4136 3656 4193 3663
rect 5047 3656 5113 3663
rect 2107 3636 2603 3643
rect 2627 3636 2933 3643
rect 3147 3636 3763 3643
rect 507 3616 583 3623
rect 1307 3616 1353 3623
rect 1447 3616 1473 3623
rect 1916 3623 1923 3633
rect 1916 3616 2333 3623
rect 2556 3616 3213 3623
rect 2556 3607 2563 3616
rect 3756 3623 3763 3636
rect 3827 3636 4133 3643
rect 4787 3636 4833 3643
rect 4927 3636 5183 3643
rect 3756 3616 3833 3623
rect 4167 3616 4353 3623
rect 4447 3616 4713 3623
rect 4727 3616 4753 3623
rect 4807 3616 4933 3623
rect 5176 3623 5183 3636
rect 5176 3616 5373 3623
rect 1387 3596 1453 3603
rect 1567 3596 1823 3603
rect 87 3576 233 3583
rect 1427 3576 1733 3583
rect 1816 3583 1823 3596
rect 1847 3596 2553 3603
rect 3067 3596 3193 3603
rect 3367 3596 3733 3603
rect 3927 3596 4473 3603
rect 4827 3596 4993 3603
rect 5067 3596 5213 3603
rect 1816 3576 2013 3583
rect 2027 3576 2413 3583
rect 2787 3576 2853 3583
rect 2927 3576 3293 3583
rect 3307 3576 3613 3583
rect 3687 3576 3753 3583
rect 4187 3576 4313 3583
rect 4327 3576 4553 3583
rect 5087 3576 5163 3583
rect 447 3556 713 3563
rect 727 3556 793 3563
rect 807 3560 1083 3563
rect 807 3556 1087 3560
rect 1073 3547 1087 3556
rect 1307 3556 1553 3563
rect 1627 3556 1813 3563
rect 2307 3556 2493 3563
rect 2716 3560 3113 3563
rect 2713 3556 3113 3560
rect 2713 3547 2727 3556
rect 3216 3556 3253 3563
rect 115 3540 173 3543
rect 113 3536 173 3540
rect 113 3527 127 3536
rect 1087 3536 1123 3543
rect 493 3527 507 3533
rect 1116 3527 1123 3536
rect 1173 3527 1187 3533
rect 1887 3536 1963 3543
rect 1733 3527 1747 3533
rect 1956 3527 1963 3536
rect 1987 3533 1992 3547
rect 2013 3533 2014 3540
rect 2156 3536 2233 3543
rect 2013 3527 2027 3533
rect 67 3513 72 3527
rect 108 3513 112 3527
rect 126 3520 127 3527
rect 148 3516 193 3523
rect 193 3507 207 3513
rect 107 3493 112 3507
rect 133 3493 134 3500
rect 347 3520 483 3523
rect 347 3516 487 3520
rect 233 3507 247 3513
rect 473 3507 487 3516
rect 567 3516 603 3523
rect 133 3483 147 3493
rect 333 3487 347 3493
rect 596 3503 603 3516
rect 627 3513 632 3527
rect 668 3513 673 3527
rect 753 3507 767 3513
rect 596 3496 633 3503
rect 927 3513 933 3527
rect 1116 3516 1133 3527
rect 1120 3513 1133 3516
rect 1227 3516 1253 3523
rect 1387 3516 1533 3523
rect 1547 3513 1552 3527
rect 1588 3516 1633 3523
rect 1647 3516 1693 3523
rect 1787 3513 1793 3527
rect 1956 3516 1973 3527
rect 1960 3513 1973 3516
rect 2127 3513 2133 3527
rect 793 3507 807 3513
rect 2156 3507 2163 3536
rect 2247 3533 2253 3547
rect 2347 3540 2483 3543
rect 2347 3536 2487 3540
rect 2287 3516 2353 3523
rect 2473 3527 2487 3536
rect 2607 3536 2653 3543
rect 2947 3534 2953 3547
rect 2940 3533 2953 3534
rect 3216 3543 3223 3556
rect 3847 3556 4433 3563
rect 5156 3563 5163 3576
rect 5156 3556 5713 3563
rect 3167 3540 3223 3543
rect 3167 3536 3227 3540
rect 2593 3523 2607 3533
rect 3213 3527 3227 3536
rect 3247 3536 3273 3543
rect 3287 3536 3333 3543
rect 3427 3536 3493 3543
rect 3453 3527 3467 3536
rect 3647 3536 3743 3543
rect 3736 3527 3743 3536
rect 4127 3536 4273 3543
rect 4747 3536 4823 3543
rect 4816 3527 4823 3536
rect 4947 3543 4960 3547
rect 4947 3540 4963 3543
rect 4947 3533 4967 3540
rect 5067 3536 5233 3543
rect 4953 3527 4967 3533
rect 2547 3520 2607 3523
rect 2547 3516 2603 3520
rect 2627 3516 2692 3523
rect 2728 3513 2733 3527
rect 2787 3516 2813 3523
rect 2867 3516 2912 3523
rect 947 3496 1033 3503
rect 1207 3496 1233 3503
rect 1247 3496 1293 3503
rect 1347 3493 1353 3507
rect 1467 3493 1473 3507
rect 1627 3496 1653 3503
rect 1667 3496 1713 3503
rect 1907 3496 2073 3503
rect 2173 3503 2187 3513
rect 2948 3520 3064 3523
rect 2948 3516 3067 3520
rect 3053 3507 3067 3516
rect 3206 3513 3207 3520
rect 3226 3520 3227 3527
rect 3233 3513 3234 3520
rect 3287 3516 3353 3523
rect 3527 3516 3713 3523
rect 3736 3516 3753 3527
rect 3740 3513 3753 3516
rect 4026 3516 4243 3523
rect 4026 3513 4027 3516
rect 3193 3507 3207 3513
rect 2173 3500 2353 3503
rect 2176 3496 2353 3500
rect 2447 3493 2453 3507
rect 2647 3496 2673 3503
rect 2827 3493 2833 3507
rect 2887 3493 2893 3507
rect 3007 3496 3032 3503
rect 3053 3500 3054 3507
rect 3107 3493 3113 3507
rect 3233 3507 3247 3513
rect 4013 3507 4027 3513
rect 4236 3507 4243 3516
rect 4267 3516 4303 3523
rect 3307 3496 3433 3503
rect 3487 3496 3572 3503
rect 3608 3493 3613 3507
rect 3727 3493 3732 3507
rect 3768 3493 3773 3507
rect 3847 3493 3853 3507
rect 4026 3500 4027 3507
rect 4048 3496 4133 3503
rect 4147 3496 4173 3503
rect 4236 3496 4253 3507
rect 4240 3493 4253 3496
rect 4296 3503 4303 3516
rect 4327 3513 4333 3527
rect 4387 3516 4433 3523
rect 4547 3516 4573 3523
rect 4647 3516 4793 3523
rect 4816 3516 4833 3527
rect 4820 3513 4833 3516
rect 4907 3513 4913 3527
rect 5113 3527 5127 3536
rect 5247 3536 5373 3543
rect 5513 3527 5527 3533
rect 5207 3516 5232 3523
rect 5268 3513 5273 3527
rect 4296 3496 4353 3503
rect 4407 3496 4493 3503
rect 4607 3493 4613 3507
rect 4667 3496 4753 3503
rect 5047 3496 5093 3503
rect 5247 3493 5253 3507
rect 5473 3503 5487 3513
rect 5427 3500 5487 3503
rect 5427 3496 5483 3500
rect 5647 3496 5693 3503
rect 373 3487 387 3493
rect 133 3480 192 3483
rect 137 3476 192 3480
rect 213 3473 214 3480
rect 287 3476 332 3483
rect 346 3480 347 3487
rect 373 3480 374 3487
rect 366 3473 367 3480
rect 513 3483 527 3493
rect 388 3480 527 3483
rect 673 3483 687 3493
rect 893 3487 907 3493
rect 673 3480 713 3483
rect 388 3476 523 3480
rect 676 3476 713 3480
rect 847 3476 883 3483
rect 213 3463 227 3473
rect 107 3460 227 3463
rect 353 3463 367 3473
rect 773 3467 787 3473
rect 353 3460 493 3463
rect 107 3456 224 3460
rect 355 3456 493 3460
rect 876 3463 883 3476
rect 1156 3467 1163 3493
rect 1287 3476 1313 3483
rect 1387 3476 1432 3483
rect 1453 3473 1454 3480
rect 1507 3476 1533 3483
rect 1556 3476 1593 3483
rect 1156 3463 1173 3467
rect 876 3456 1173 3463
rect 1160 3453 1173 3456
rect 1453 3463 1467 3473
rect 1556 3463 1563 3476
rect 1753 3483 1767 3493
rect 2113 3487 2127 3493
rect 1607 3476 1843 3483
rect 1453 3460 1563 3463
rect 1457 3456 1563 3460
rect 1836 3463 1843 3476
rect 1867 3473 1873 3487
rect 1927 3473 1933 3487
rect 2227 3476 2253 3483
rect 2267 3476 2333 3483
rect 2493 3483 2507 3493
rect 2427 3480 2507 3483
rect 2427 3476 2503 3480
rect 3087 3473 3093 3487
rect 3473 3483 3487 3493
rect 3407 3480 3487 3483
rect 3407 3476 3483 3480
rect 3507 3476 3593 3483
rect 3887 3476 4153 3483
rect 4467 3473 4473 3487
rect 4727 3473 4733 3487
rect 5133 3483 5147 3493
rect 5133 3480 5253 3483
rect 5136 3476 5253 3480
rect 5293 3483 5307 3493
rect 5493 3487 5507 3493
rect 5293 3480 5373 3483
rect 5296 3476 5373 3480
rect 5387 3476 5473 3483
rect 5487 3480 5507 3487
rect 5487 3476 5503 3480
rect 5487 3473 5500 3476
rect 5607 3473 5613 3487
rect 1836 3456 2153 3463
rect 1513 3447 1527 3456
rect 2373 3463 2387 3473
rect 2373 3460 2493 3463
rect 2376 3456 2493 3460
rect 307 3436 373 3443
rect 767 3436 893 3443
rect 1007 3436 1353 3443
rect 1526 3440 1527 3447
rect 1548 3436 1573 3443
rect 1907 3436 1993 3443
rect 2047 3436 2253 3443
rect 2376 3443 2383 3456
rect 2507 3456 2593 3463
rect 3687 3456 3873 3463
rect 4513 3463 4527 3473
rect 4267 3460 4527 3463
rect 4267 3456 4523 3460
rect 4773 3463 4787 3473
rect 4627 3460 4787 3463
rect 4627 3456 4783 3460
rect 5653 3463 5667 3473
rect 5547 3460 5667 3463
rect 5547 3456 5663 3460
rect 2307 3436 2383 3443
rect 2787 3436 2833 3443
rect 3447 3436 3893 3443
rect 3967 3436 4433 3443
rect 4487 3436 4573 3443
rect 5087 3436 5293 3443
rect 1707 3416 2212 3423
rect 2248 3416 2293 3423
rect 3167 3416 3233 3423
rect 3547 3416 3573 3423
rect 3587 3416 3772 3423
rect 3808 3416 4413 3423
rect 4487 3416 4763 3423
rect 207 3396 1013 3403
rect 1487 3396 2293 3403
rect 3087 3396 3673 3403
rect 3687 3396 3893 3403
rect 3907 3396 4033 3403
rect 4147 3396 4733 3403
rect 4756 3403 4763 3416
rect 5567 3416 5633 3423
rect 4756 3396 4973 3403
rect 5207 3396 5293 3403
rect 5627 3396 5693 3403
rect 1447 3376 1853 3383
rect 1987 3376 2253 3383
rect 2527 3376 2713 3383
rect 3427 3376 3993 3383
rect 4036 3376 4113 3383
rect 127 3356 773 3363
rect 787 3356 833 3363
rect 847 3356 913 3363
rect 1167 3356 1873 3363
rect 2007 3356 2973 3363
rect 3167 3356 3373 3363
rect 4036 3363 4043 3376
rect 4587 3376 5033 3383
rect 5047 3376 5193 3383
rect 3867 3356 4043 3363
rect 4056 3356 4233 3363
rect 1347 3336 1553 3343
rect 1747 3336 2093 3343
rect 2107 3333 2113 3347
rect 2307 3336 2713 3343
rect 2787 3336 2933 3343
rect 467 3316 703 3323
rect 487 3296 533 3303
rect 696 3303 703 3316
rect 727 3316 853 3323
rect 1247 3316 1963 3323
rect 696 3296 1133 3303
rect 1487 3296 1613 3303
rect 1676 3296 1733 3303
rect 87 3276 233 3283
rect 116 3247 123 3276
rect 396 3276 493 3283
rect 346 3253 347 3260
rect 396 3263 403 3276
rect 727 3276 1013 3283
rect 1327 3283 1340 3287
rect 1327 3273 1343 3283
rect 533 3267 547 3273
rect 368 3256 403 3263
rect 427 3256 503 3263
rect 333 3247 347 3253
rect 496 3247 503 3256
rect 893 3247 907 3253
rect 67 3233 73 3247
rect 206 3233 207 3240
rect 228 3233 232 3247
rect 268 3236 293 3243
rect 496 3236 513 3247
rect 500 3233 513 3236
rect 566 3233 567 3240
rect 588 3236 612 3243
rect 648 3233 653 3247
rect 667 3236 753 3243
rect 847 3233 853 3247
rect 1146 3253 1147 3260
rect 1168 3254 1173 3267
rect 1168 3253 1180 3254
rect 1013 3247 1027 3253
rect 1133 3247 1147 3253
rect 1336 3247 1343 3273
rect 1407 3256 1633 3263
rect 1676 3247 1683 3296
rect 1956 3303 1963 3316
rect 1987 3316 2453 3323
rect 2716 3323 2723 3333
rect 3387 3336 3453 3343
rect 4056 3343 4063 3356
rect 4387 3356 4613 3363
rect 4767 3356 4873 3363
rect 4947 3356 5533 3363
rect 3727 3336 4063 3343
rect 4087 3336 5153 3343
rect 5607 3336 5693 3343
rect 2716 3316 2813 3323
rect 4047 3316 4392 3323
rect 4428 3316 4583 3323
rect 1956 3296 2193 3303
rect 2207 3296 2433 3303
rect 2747 3296 2833 3303
rect 3187 3296 3533 3303
rect 4107 3296 4253 3303
rect 4347 3296 4373 3303
rect 4387 3296 4533 3303
rect 4576 3303 4583 3316
rect 4607 3316 4933 3323
rect 5227 3316 5253 3323
rect 4576 3296 4632 3303
rect 4668 3296 4733 3303
rect 4827 3296 4853 3303
rect 5247 3296 5573 3303
rect 1706 3273 1707 3280
rect 1728 3276 1793 3283
rect 2287 3280 2403 3283
rect 2287 3276 2407 3280
rect 1693 3267 1707 3273
rect 2193 3267 2207 3273
rect 2393 3267 2407 3276
rect 2647 3276 2793 3283
rect 2807 3276 2993 3283
rect 3047 3276 3573 3283
rect 4307 3276 4483 3283
rect 4476 3267 4483 3276
rect 4807 3276 4913 3283
rect 4987 3276 5073 3283
rect 5087 3273 5093 3287
rect 1747 3256 1773 3263
rect 1907 3253 1913 3267
rect 1967 3253 1973 3267
rect 1987 3256 2013 3263
rect 2067 3253 2073 3267
rect 2127 3256 2153 3263
rect 2267 3253 2272 3267
rect 2306 3253 2307 3260
rect 2328 3263 2340 3267
rect 2328 3253 2343 3263
rect 2467 3260 2523 3263
rect 2467 3256 2527 3260
rect 2293 3247 2307 3253
rect 2336 3247 2343 3253
rect 2513 3247 2527 3256
rect 2713 3247 2727 3253
rect 3107 3256 3213 3263
rect 3227 3253 3233 3267
rect 4107 3253 4113 3267
rect 4167 3253 4173 3267
rect 4547 3256 4573 3263
rect 4627 3256 4653 3263
rect 4680 3263 4693 3267
rect 4676 3253 4693 3263
rect 4747 3253 4753 3267
rect 5167 3256 5293 3263
rect 5307 3260 5343 3263
rect 5376 3260 5433 3263
rect 5307 3256 5347 3260
rect 3053 3247 3067 3253
rect 3533 3247 3547 3253
rect 4473 3247 4487 3253
rect 1067 3236 1093 3243
rect 1187 3233 1193 3247
rect 1287 3233 1293 3247
rect 1376 3236 1413 3243
rect 193 3227 207 3233
rect 373 3227 387 3233
rect 107 3213 112 3227
rect 148 3216 193 3223
rect 247 3216 363 3223
rect 356 3203 363 3216
rect 553 3223 567 3233
rect 1376 3227 1383 3236
rect 1727 3236 1773 3243
rect 1927 3233 1933 3247
rect 2047 3236 2113 3243
rect 2306 3240 2307 3247
rect 2347 3236 2373 3243
rect 2567 3233 2573 3247
rect 2667 3233 2673 3247
rect 2856 3240 2913 3243
rect 2853 3236 2913 3240
rect 2173 3227 2187 3233
rect 553 3220 612 3223
rect 555 3216 612 3220
rect 633 3213 634 3220
rect 847 3216 873 3223
rect 947 3216 993 3223
rect 1046 3213 1047 3220
rect 1068 3216 1313 3223
rect 1367 3216 1383 3227
rect 1456 3220 1513 3223
rect 1453 3216 1513 3220
rect 1367 3213 1380 3216
rect 356 3196 473 3203
rect 633 3203 647 3213
rect 487 3200 647 3203
rect 487 3196 644 3200
rect 807 3196 853 3203
rect 867 3196 893 3203
rect 1033 3203 1047 3213
rect 1453 3207 1467 3216
rect 1527 3216 1572 3223
rect 1608 3216 1653 3223
rect 1887 3216 1973 3223
rect 2413 3227 2427 3233
rect 2853 3227 2867 3236
rect 3007 3233 3013 3247
rect 3067 3236 3183 3243
rect 2647 3216 2693 3223
rect 2807 3213 2813 3227
rect 2867 3216 3033 3223
rect 3107 3216 3133 3223
rect 3176 3226 3183 3236
rect 3267 3236 3293 3243
rect 3427 3233 3433 3247
rect 3487 3233 3493 3247
rect 3713 3233 3714 3240
rect 3713 3227 3727 3233
rect 3953 3227 3967 3233
rect 1033 3200 1253 3203
rect 1036 3196 1253 3200
rect 1307 3196 1353 3203
rect 2167 3196 2373 3203
rect 2533 3203 2547 3213
rect 2733 3207 2747 3213
rect 3447 3213 3453 3227
rect 3476 3216 3513 3223
rect 2533 3200 2653 3203
rect 2536 3196 2653 3200
rect 2787 3196 2833 3203
rect 2907 3196 2953 3203
rect 3427 3196 3453 3203
rect 3476 3203 3483 3216
rect 3587 3213 3593 3227
rect 3687 3213 3692 3227
rect 3713 3220 3714 3227
rect 3787 3216 3833 3223
rect 3907 3213 3913 3227
rect 4220 3243 4232 3247
rect 4133 3223 4147 3233
rect 4216 3233 4232 3243
rect 4268 3233 4273 3247
rect 4387 3233 4393 3247
rect 4567 3236 4593 3243
rect 4676 3243 4683 3253
rect 4973 3247 4987 3253
rect 5333 3247 5347 3256
rect 4647 3236 4683 3243
rect 4727 3233 4733 3247
rect 4807 3233 4813 3247
rect 4867 3236 4933 3243
rect 5027 3236 5073 3243
rect 5256 3240 5333 3243
rect 5253 3236 5333 3240
rect 4216 3223 4223 3233
rect 5253 3227 5267 3236
rect 5373 3256 5433 3260
rect 5373 3247 5387 3256
rect 5513 3247 5527 3253
rect 5416 3236 5473 3243
rect 4133 3220 4223 3223
rect 4136 3216 4223 3220
rect 4247 3213 4253 3227
rect 4307 3213 4313 3227
rect 4787 3213 4793 3227
rect 4820 3223 4833 3227
rect 4816 3213 4833 3223
rect 4927 3216 4993 3223
rect 5047 3213 5053 3227
rect 5207 3213 5213 3227
rect 5307 3213 5313 3227
rect 5416 3223 5423 3236
rect 5527 3240 5624 3243
rect 5527 3236 5627 3240
rect 5613 3227 5627 3236
rect 5367 3216 5423 3223
rect 5436 3216 5493 3223
rect 3467 3196 3483 3203
rect 4367 3193 4373 3207
rect 4507 3196 4533 3203
rect 4816 3203 4823 3213
rect 4667 3196 4823 3203
rect 4873 3203 4887 3213
rect 5436 3207 5443 3216
rect 5587 3213 5592 3227
rect 5613 3220 5614 3227
rect 4873 3200 5073 3203
rect 4876 3196 5073 3200
rect 5147 3193 5153 3207
rect 5247 3196 5353 3203
rect 5427 3196 5443 3207
rect 5427 3193 5440 3196
rect 5547 3196 5633 3203
rect 1127 3176 1273 3183
rect 1813 3183 1827 3193
rect 3233 3187 3247 3193
rect 1813 3180 1833 3183
rect 1816 3176 1833 3180
rect 1847 3176 2353 3183
rect 2427 3176 2773 3183
rect 2787 3173 2793 3187
rect 3387 3176 3413 3183
rect 4327 3176 4433 3183
rect 4527 3176 4793 3183
rect 5127 3176 5163 3183
rect 1107 3156 1193 3163
rect 1267 3156 1723 3163
rect 207 3136 1393 3143
rect 1716 3143 1723 3156
rect 1927 3156 2133 3163
rect 2347 3156 2373 3163
rect 2627 3156 2853 3163
rect 2867 3156 3233 3163
rect 4307 3156 4493 3163
rect 4867 3156 5133 3163
rect 5156 3163 5163 3176
rect 5156 3156 5393 3163
rect 5527 3156 5613 3163
rect 1716 3136 2113 3143
rect 2127 3136 2313 3143
rect 2500 3143 2513 3147
rect 2496 3134 2513 3143
rect 2496 3133 2520 3134
rect 2587 3136 2893 3143
rect 2967 3136 3153 3143
rect 3527 3136 3833 3143
rect 4427 3136 4623 3143
rect 707 3116 773 3123
rect 947 3116 1053 3123
rect 1187 3116 1293 3123
rect 1767 3116 2093 3123
rect 2187 3116 2403 3123
rect 2396 3107 2403 3116
rect 2427 3116 2453 3123
rect 167 3096 273 3103
rect 287 3096 1733 3103
rect 1867 3096 1992 3103
rect 2013 3093 2014 3100
rect 2067 3096 2273 3103
rect 2396 3096 2412 3107
rect 2400 3093 2412 3096
rect 2448 3096 2473 3103
rect 2496 3103 2503 3133
rect 2527 3116 3233 3123
rect 3387 3116 3672 3123
rect 3708 3116 4073 3123
rect 4616 3123 4623 3136
rect 4747 3136 4993 3143
rect 5067 3136 5153 3143
rect 5487 3136 5553 3143
rect 4616 3116 4883 3123
rect 4876 3107 4883 3116
rect 5027 3116 5283 3123
rect 2496 3096 2643 3103
rect 2013 3087 2027 3093
rect 367 3076 613 3083
rect 1327 3076 1453 3083
rect 2013 3080 2014 3087
rect 2127 3076 2233 3083
rect 2367 3076 2433 3083
rect 2447 3076 2593 3083
rect 2636 3083 2643 3096
rect 2667 3096 2733 3103
rect 2927 3096 3473 3103
rect 3487 3096 3653 3103
rect 3847 3096 4433 3103
rect 4547 3096 4743 3103
rect 2636 3076 2723 3083
rect 293 3067 307 3073
rect 407 3056 533 3063
rect 547 3056 673 3063
rect 747 3056 903 3063
rect 896 3047 903 3056
rect 1007 3053 1012 3067
rect 1048 3060 1523 3063
rect 1048 3056 1527 3060
rect 1513 3047 1527 3056
rect 2113 3053 2114 3060
rect 2427 3056 2553 3063
rect 2616 3060 2693 3063
rect 2613 3056 2693 3060
rect 147 3033 153 3047
rect 447 3033 453 3047
rect 507 3033 512 3047
rect 533 3033 534 3040
rect 787 3036 872 3043
rect 908 3033 913 3047
rect 987 3033 993 3047
rect 1047 3036 1113 3043
rect 1256 3040 1373 3043
rect 1253 3036 1373 3040
rect 393 3027 407 3033
rect 533 3027 547 3033
rect 107 3016 183 3023
rect 176 3007 183 3016
rect 227 3013 233 3027
rect 347 3013 353 3027
rect 487 3013 493 3027
rect 627 3013 633 3027
rect 687 3016 733 3023
rect 847 3013 852 3027
rect 888 3013 893 3027
rect 913 3023 927 3033
rect 1253 3027 1267 3036
rect 1447 3036 1473 3043
rect 1567 3033 1573 3047
rect 1707 3036 1773 3043
rect 1887 3033 1893 3047
rect 1947 3036 1993 3043
rect 2066 3033 2067 3040
rect 2088 3034 2092 3047
rect 2113 3047 2127 3053
rect 2613 3047 2627 3056
rect 2716 3047 2723 3076
rect 2787 3076 2813 3083
rect 2987 3076 3373 3083
rect 3507 3076 3793 3083
rect 4246 3073 4247 3080
rect 4268 3076 4373 3083
rect 4527 3076 4592 3083
rect 4628 3076 4713 3083
rect 4736 3083 4743 3096
rect 4887 3096 5113 3103
rect 5127 3096 5253 3103
rect 5276 3103 5283 3116
rect 5467 3116 5613 3123
rect 5276 3096 5593 3103
rect 4736 3076 4913 3083
rect 4233 3067 4247 3073
rect 2753 3047 2767 3053
rect 3047 3056 3092 3063
rect 3128 3060 3283 3063
rect 3128 3056 3287 3060
rect 2893 3047 2907 3053
rect 3273 3047 3287 3056
rect 3307 3060 3423 3063
rect 3307 3056 3427 3060
rect 3413 3047 3427 3056
rect 3887 3056 3913 3063
rect 3936 3056 4013 3063
rect 2113 3040 2114 3047
rect 2088 3033 2100 3034
rect 2187 3033 2193 3047
rect 2307 3033 2313 3047
rect 2366 3033 2367 3040
rect 2388 3033 2393 3047
rect 2626 3040 2627 3047
rect 2648 3033 2653 3047
rect 2847 3033 2853 3047
rect 3147 3036 3223 3043
rect 1833 3027 1847 3033
rect 2053 3027 2067 3033
rect 2353 3027 2367 3033
rect 913 3020 1033 3023
rect 916 3016 1033 3020
rect 1056 3016 1113 3023
rect 187 2993 193 3007
rect 247 2996 272 3003
rect 308 2993 313 3007
rect 373 2983 387 2993
rect 1056 3003 1063 3016
rect 1227 3016 1253 3023
rect 1367 3013 1373 3027
rect 1487 3013 1492 3027
rect 1528 3013 1533 3027
rect 1767 3016 1793 3023
rect 1907 3013 1913 3027
rect 1967 3013 1973 3027
rect 2066 3020 2067 3027
rect 2088 3013 2093 3027
rect 2147 3016 2213 3023
rect 2487 3013 2493 3027
rect 2547 3016 2573 3023
rect 2587 3013 2593 3027
rect 2647 3013 2653 3027
rect 2707 3016 2733 3023
rect 2827 3016 2873 3023
rect 2927 3016 2993 3023
rect 3093 3023 3107 3033
rect 3047 3020 3107 3023
rect 3047 3016 3103 3020
rect 3127 3013 3132 3027
rect 3168 3016 3173 3023
rect 3187 3013 3193 3027
rect 3216 3023 3223 3036
rect 3247 3033 3252 3047
rect 3286 3040 3287 3047
rect 3293 3033 3294 3040
rect 3347 3036 3373 3043
rect 3547 3033 3552 3047
rect 3588 3033 3593 3047
rect 3767 3033 3773 3047
rect 3936 3043 3943 3056
rect 4246 3060 4247 3067
rect 4616 3060 4743 3063
rect 4093 3047 4107 3053
rect 4353 3047 4367 3053
rect 4613 3056 4747 3060
rect 3907 3036 3943 3043
rect 3293 3027 3307 3033
rect 3216 3016 3253 3023
rect 3387 3013 3393 3027
rect 3447 3013 3453 3027
rect 3707 3016 3733 3023
rect 3993 3023 4007 3033
rect 3927 3020 4007 3023
rect 4033 3027 4047 3033
rect 3927 3016 4003 3020
rect 4213 3023 4227 3033
rect 4147 3020 4227 3023
rect 4253 3027 4267 3033
rect 4447 3036 4573 3043
rect 4613 3047 4627 3056
rect 4733 3047 4747 3056
rect 4787 3056 5193 3063
rect 5207 3056 5292 3063
rect 5313 3053 5314 3060
rect 5367 3056 5473 3063
rect 5547 3053 5553 3067
rect 4773 3047 4787 3053
rect 5313 3047 5327 3053
rect 5036 3040 5233 3043
rect 5033 3036 5233 3040
rect 4313 3027 4327 3033
rect 4147 3016 4223 3020
rect 4326 3020 4327 3027
rect 4333 3013 4334 3020
rect 4387 3016 4413 3023
rect 4580 3026 4593 3027
rect 4507 3016 4563 3023
rect 987 2996 1063 3003
rect 1087 2993 1093 3007
rect 1147 2996 1253 3003
rect 1267 2993 1273 3007
rect 1293 3003 1307 3013
rect 1293 3000 1353 3003
rect 1296 2996 1353 3000
rect 1407 2996 1453 3003
rect 1516 3003 1523 3013
rect 1467 2996 1523 3003
rect 1827 2996 1993 3003
rect 2307 2996 2473 3003
rect 2527 2996 2553 3003
rect 2567 2996 2633 3003
rect 2773 3003 2787 3013
rect 3653 3007 3667 3013
rect 2773 3000 2913 3003
rect 2776 2996 2913 3000
rect 3427 2996 3552 3003
rect 3588 2996 3653 3003
rect 3727 2996 4013 3003
rect 4067 2996 4093 3003
rect 4107 2996 4173 3003
rect 4333 3003 4347 3013
rect 4247 3000 4347 3003
rect 4247 2996 4344 3000
rect 4487 2993 4492 3007
rect 4513 2993 4514 3000
rect 4556 3003 4563 3016
rect 4587 3013 4593 3026
rect 4653 3023 4667 3033
rect 5033 3027 5047 3036
rect 5326 3040 5327 3047
rect 5333 3033 5334 3040
rect 5353 3033 5354 3040
rect 5407 3036 5453 3043
rect 5507 3036 5573 3043
rect 5587 3033 5593 3047
rect 5333 3027 5347 3033
rect 4653 3020 4693 3023
rect 4656 3016 4693 3020
rect 4780 3026 4793 3027
rect 4766 3013 4767 3020
rect 4633 3003 4647 3013
rect 4753 3007 4767 3013
rect 4788 3013 4793 3026
rect 4886 3013 4887 3020
rect 4908 3016 4952 3023
rect 4988 3013 4993 3027
rect 5127 3013 5133 3027
rect 5187 3013 5193 3027
rect 5287 3013 5293 3027
rect 5346 3020 5347 3027
rect 5353 3027 5367 3033
rect 5353 3020 5354 3027
rect 4873 3007 4887 3013
rect 4556 3000 4647 3003
rect 4556 2996 4643 3000
rect 4766 3000 4767 3007
rect 4847 2993 4852 3007
rect 4873 3000 4874 3007
rect 4927 2993 4933 3007
rect 5087 2993 5093 3007
rect 5147 2993 5153 3007
rect 5433 3003 5447 3013
rect 5327 3000 5447 3003
rect 5527 3016 5613 3023
rect 5473 3007 5487 3013
rect 5327 2996 5443 3000
rect 653 2987 667 2993
rect 1353 2987 1367 2993
rect 373 2980 493 2983
rect 376 2976 493 2980
rect 667 2976 873 2983
rect 1567 2976 1873 2983
rect 2407 2976 2493 2983
rect 2847 2976 3113 2983
rect 3247 2976 3592 2983
rect 3628 2976 3733 2983
rect 3747 2976 3973 2983
rect 4047 2976 4252 2983
rect 4288 2976 4373 2983
rect 4513 2983 4527 2993
rect 4447 2980 4527 2983
rect 4447 2976 4524 2980
rect 4787 2976 4973 2983
rect 5013 2983 5027 2993
rect 5013 2980 5092 2983
rect 5016 2976 5092 2980
rect 5128 2976 5153 2983
rect 5287 2983 5300 2987
rect 5287 2973 5303 2983
rect 87 2956 273 2963
rect 287 2956 373 2963
rect 627 2956 833 2963
rect 847 2956 1193 2963
rect 1367 2956 1433 2963
rect 1447 2956 1613 2963
rect 1807 2956 1953 2963
rect 2027 2953 2033 2967
rect 2447 2956 2553 2963
rect 2827 2956 2973 2963
rect 3067 2956 3393 2963
rect 3687 2956 4093 2963
rect 4187 2956 4653 2963
rect 4767 2956 4953 2963
rect 573 2947 587 2953
rect 5167 2956 5233 2963
rect 5296 2963 5303 2973
rect 5296 2956 5553 2963
rect 267 2936 293 2943
rect 1267 2936 1473 2943
rect 1827 2936 2093 2943
rect 2107 2936 2233 2943
rect 2307 2936 2653 2943
rect 3007 2936 3193 2943
rect 3207 2936 3373 2943
rect 3547 2936 4052 2943
rect 4088 2936 4113 2943
rect 4487 2936 4553 2943
rect 4767 2936 4833 2943
rect 4927 2936 4973 2943
rect 5307 2936 5533 2943
rect 47 2916 193 2923
rect 487 2916 993 2923
rect 2327 2916 2973 2923
rect 3607 2916 3853 2923
rect 3867 2916 4013 2923
rect 4127 2916 4272 2923
rect 4308 2916 4352 2923
rect 4388 2916 4883 2923
rect 4876 2907 4883 2916
rect 4927 2916 4953 2923
rect 5007 2916 5393 2923
rect 5607 2916 5633 2923
rect 27 2896 73 2903
rect 507 2896 593 2903
rect 1667 2896 2543 2903
rect 1947 2876 2313 2883
rect 2536 2883 2543 2896
rect 2627 2896 2953 2903
rect 3047 2896 3453 2903
rect 3927 2896 4253 2903
rect 4327 2896 4473 2903
rect 4527 2896 4793 2903
rect 4887 2896 5213 2903
rect 5236 2896 5393 2903
rect 2536 2876 2713 2883
rect 2727 2876 3013 2883
rect 3127 2876 3713 2883
rect 3787 2876 3853 2883
rect 4056 2876 4132 2883
rect 847 2856 932 2863
rect 968 2856 993 2863
rect 1087 2856 1133 2863
rect 1147 2856 1613 2863
rect 1707 2856 1873 2863
rect 1887 2856 2133 2863
rect 2187 2856 2353 2863
rect 3107 2856 3312 2863
rect 3348 2856 3453 2863
rect 4056 2863 4063 2876
rect 4168 2876 4373 2883
rect 4427 2876 4993 2883
rect 5236 2883 5243 2896
rect 5087 2876 5243 2883
rect 5267 2876 5353 2883
rect 3787 2856 4063 2863
rect 4076 2856 4653 2863
rect 147 2836 213 2843
rect 887 2836 913 2843
rect 927 2836 1273 2843
rect 1987 2836 2153 2843
rect 2176 2836 2273 2843
rect 67 2816 173 2823
rect 187 2816 213 2823
rect 547 2816 793 2823
rect 816 2816 1053 2823
rect -24 2796 13 2803
rect 256 2800 293 2803
rect 213 2787 227 2793
rect 117 2780 173 2783
rect 113 2776 173 2780
rect 113 2767 127 2776
rect 253 2796 293 2800
rect 253 2787 267 2796
rect 307 2796 373 2803
rect 816 2803 823 2816
rect 1076 2816 1233 2823
rect 507 2796 823 2803
rect 1076 2787 1083 2816
rect 1247 2816 1733 2823
rect 1927 2816 2092 2823
rect 2176 2823 2183 2836
rect 2487 2836 2513 2843
rect 2687 2836 2913 2843
rect 3447 2836 3733 2843
rect 4076 2843 4083 2856
rect 4747 2856 4933 2863
rect 4947 2856 5133 2863
rect 5187 2856 5233 2863
rect 3787 2836 4083 2843
rect 4107 2836 4713 2843
rect 4727 2836 4913 2843
rect 5227 2836 5433 2843
rect 5447 2836 5693 2843
rect 2128 2816 2183 2823
rect 2267 2816 2573 2823
rect 3587 2816 3653 2823
rect 3727 2816 3813 2823
rect 4027 2816 4383 2823
rect 276 2780 373 2783
rect 273 2776 373 2780
rect 273 2767 287 2776
rect 493 2767 507 2773
rect -24 2756 13 2763
rect 67 2753 72 2767
rect 113 2760 114 2767
rect 106 2753 107 2760
rect 220 2766 233 2767
rect 93 2747 107 2753
rect 227 2753 233 2766
rect 387 2753 392 2767
rect 428 2756 453 2763
rect 776 2780 952 2783
rect 533 2767 547 2773
rect 773 2776 952 2780
rect 773 2767 787 2776
rect 607 2756 653 2763
rect 667 2756 733 2763
rect 873 2767 887 2776
rect 988 2776 1013 2783
rect 1067 2776 1083 2787
rect 1156 2800 1213 2803
rect 1113 2787 1127 2793
rect 1067 2773 1080 2776
rect 1153 2796 1213 2800
rect 1153 2787 1167 2796
rect 1956 2800 2033 2803
rect 1953 2796 2033 2800
rect 1953 2787 1967 2796
rect 2047 2796 2473 2803
rect 2867 2796 2993 2803
rect 3347 2796 3373 2803
rect 3567 2796 3613 2803
rect 3687 2796 3873 2803
rect 3947 2796 4053 2803
rect 4376 2803 4383 2816
rect 4407 2816 4533 2823
rect 4827 2816 4893 2823
rect 5007 2816 5033 2823
rect 5347 2816 5373 2823
rect 5396 2816 5553 2823
rect 4107 2796 4283 2803
rect 4376 2796 4403 2803
rect 1287 2776 1393 2783
rect 1407 2776 1673 2783
rect 1233 2767 1247 2773
rect 1553 2767 1567 2776
rect 1687 2776 1853 2783
rect 1907 2773 1913 2787
rect 2076 2780 2113 2783
rect 2073 2776 2113 2780
rect 2073 2767 2087 2776
rect 2167 2773 2172 2787
rect 2208 2776 2253 2783
rect 2387 2776 2412 2783
rect 2448 2773 2453 2787
rect 2547 2776 2593 2783
rect 2853 2767 2867 2773
rect 3436 2780 3533 2783
rect 3093 2767 3107 2773
rect 927 2753 933 2767
rect 987 2756 1032 2763
rect 1068 2756 1133 2763
rect 1246 2760 1247 2767
rect 1268 2753 1273 2767
rect 1467 2756 1513 2763
rect 1707 2756 1873 2763
rect 2007 2756 2033 2763
rect 2167 2753 2173 2767
rect 2447 2756 2533 2763
rect 2767 2756 2813 2763
rect 2947 2753 2953 2767
rect 3007 2756 3033 2763
rect 3433 2776 3533 2780
rect 3433 2767 3447 2776
rect 3907 2776 3933 2783
rect 3593 2767 3607 2773
rect 3487 2756 3572 2763
rect 3593 2760 3594 2767
rect 3947 2753 3953 2767
rect 3973 2763 3987 2773
rect 4053 2767 4067 2773
rect 4276 2783 4283 2796
rect 4396 2783 4403 2796
rect 4467 2796 4513 2803
rect 4687 2796 4963 2803
rect 4276 2776 4383 2783
rect 4396 2776 4493 2783
rect 4253 2767 4267 2773
rect 3973 2760 4013 2763
rect 3976 2756 4013 2760
rect 4107 2753 4113 2767
rect 4207 2753 4213 2767
rect 4347 2753 4353 2767
rect 1653 2747 1667 2753
rect 1933 2747 1947 2753
rect 2313 2747 2327 2753
rect 2573 2747 2587 2753
rect 27 2733 33 2747
rect 106 2740 107 2747
rect 147 2733 152 2747
rect 188 2736 293 2743
rect 307 2736 333 2743
rect 387 2733 393 2747
rect 447 2736 513 2743
rect 553 2727 567 2733
rect 747 2733 753 2747
rect 807 2736 853 2743
rect 867 2733 872 2747
rect 893 2733 894 2740
rect 1367 2736 1433 2743
rect 1447 2736 1492 2743
rect 1528 2733 1533 2747
rect 1680 2743 1693 2747
rect 1676 2733 1693 2743
rect 1827 2733 1833 2747
rect 2007 2736 2053 2743
rect 2107 2733 2113 2747
rect 2367 2733 2373 2747
rect 2547 2733 2552 2747
rect 2573 2740 2574 2747
rect 2787 2733 2793 2747
rect 2907 2736 2933 2743
rect 2987 2733 2993 2747
rect 653 2727 667 2733
rect 893 2723 907 2733
rect 676 2720 907 2723
rect 676 2716 903 2720
rect 247 2696 453 2703
rect 676 2703 683 2716
rect 987 2716 1012 2723
rect 1048 2716 1113 2723
rect 1127 2716 1333 2723
rect 1573 2723 1587 2733
rect 1573 2720 1613 2723
rect 1576 2716 1613 2720
rect 1676 2723 1683 2733
rect 1773 2727 1787 2733
rect 2733 2727 2747 2733
rect 1627 2716 1713 2723
rect 1887 2716 1953 2723
rect 467 2696 683 2703
rect 2007 2696 2193 2703
rect 2287 2696 2393 2703
rect 2647 2696 2773 2703
rect 2836 2703 2843 2733
rect 3233 2727 3247 2733
rect 2867 2716 3113 2723
rect 3127 2716 3153 2723
rect 3347 2736 3453 2743
rect 3733 2747 3747 2753
rect 4013 2747 4027 2753
rect 4376 2747 4383 2776
rect 4547 2776 4573 2783
rect 4956 2783 4963 2796
rect 4987 2796 5123 2803
rect 4956 2776 5032 2783
rect 5068 2773 5073 2787
rect 5116 2783 5123 2796
rect 5396 2803 5403 2816
rect 5727 2816 5783 2823
rect 5207 2796 5403 2803
rect 5427 2800 5483 2803
rect 5427 2796 5487 2800
rect 5473 2787 5487 2796
rect 5116 2776 5293 2783
rect 5307 2773 5313 2787
rect 5367 2773 5373 2787
rect 5707 2796 5763 2803
rect 5513 2787 5527 2793
rect 4873 2767 4887 2773
rect 4407 2756 4513 2763
rect 4626 2753 4627 2760
rect 4648 2753 4653 2767
rect 4707 2756 4753 2763
rect 4807 2753 4813 2767
rect 4947 2756 5032 2763
rect 5068 2756 5172 2763
rect 5208 2753 5213 2767
rect 5407 2753 5413 2767
rect 5467 2756 5492 2763
rect 5528 2756 5633 2763
rect 5647 2753 5653 2767
rect 5727 2756 5763 2763
rect 4613 2747 4627 2753
rect 3667 2736 3693 2743
rect 3787 2733 3793 2747
rect 3847 2733 3853 2747
rect 4013 2740 4032 2747
rect 4016 2736 4032 2740
rect 4020 2733 4032 2736
rect 4068 2733 4073 2747
rect 4187 2733 4193 2747
rect 4220 2743 4233 2747
rect 4216 2733 4233 2743
rect 3273 2727 3287 2733
rect 3667 2716 3713 2723
rect 4216 2723 4223 2733
rect 4147 2716 4223 2723
rect 4273 2727 4287 2733
rect 4547 2736 4592 2743
rect 4626 2740 4627 2747
rect 4648 2736 4673 2743
rect 4747 2736 4773 2743
rect 4827 2736 4872 2743
rect 4893 2733 4894 2740
rect 4967 2733 4973 2747
rect 5027 2736 5153 2743
rect 5167 2736 5193 2743
rect 5287 2736 5353 2743
rect 5567 2736 5593 2743
rect 5776 2743 5783 2816
rect 5756 2736 5783 2743
rect 4333 2723 4347 2733
rect 4333 2720 4413 2723
rect 4336 2716 4413 2720
rect 4536 2723 4543 2733
rect 4536 2716 4693 2723
rect 4893 2723 4907 2733
rect 4807 2720 4907 2723
rect 4807 2716 4904 2720
rect 5647 2716 5673 2723
rect 2836 2696 2953 2703
rect 3427 2696 3773 2703
rect 3947 2696 4173 2703
rect 4727 2693 4733 2707
rect 4867 2696 4993 2703
rect 5007 2696 5093 2703
rect 5207 2696 5233 2703
rect 27 2676 2653 2683
rect 2747 2676 2853 2683
rect 2947 2676 3053 2683
rect 3407 2676 3833 2683
rect 4067 2676 4252 2683
rect 4288 2676 4593 2683
rect 4647 2676 4793 2683
rect 5007 2676 5332 2683
rect 5368 2676 5453 2683
rect 5687 2673 5693 2687
rect 47 2656 1073 2663
rect 1667 2656 1813 2663
rect 1867 2656 2313 2663
rect 2587 2656 3293 2663
rect 3447 2656 3773 2663
rect 4207 2656 4313 2663
rect 4327 2656 4693 2663
rect 4767 2656 4873 2663
rect 4967 2656 5152 2663
rect 5188 2656 5253 2663
rect 5327 2656 5713 2663
rect 336 2640 633 2643
rect 333 2636 633 2640
rect 333 2627 347 2636
rect 727 2636 833 2643
rect 1027 2636 1453 2643
rect 1467 2636 1693 2643
rect 1787 2636 2493 2643
rect 2927 2636 3033 2643
rect 3087 2636 3233 2643
rect 3287 2636 3333 2643
rect 3356 2636 3413 2643
rect 447 2616 573 2623
rect 807 2616 973 2623
rect 1207 2613 1213 2627
rect 1407 2616 1513 2623
rect 1627 2616 2153 2623
rect 2367 2613 2373 2627
rect 2467 2616 2793 2623
rect 2847 2616 2873 2623
rect 3356 2623 3363 2636
rect 3547 2636 4293 2643
rect 4447 2636 4573 2643
rect 4587 2636 4853 2643
rect 5407 2636 5473 2643
rect 3227 2616 3363 2623
rect 3387 2616 3433 2623
rect 3587 2616 3633 2623
rect 3947 2616 4052 2623
rect 4088 2616 4393 2623
rect 4607 2616 5073 2623
rect 5756 2623 5763 2736
rect 5707 2616 5763 2623
rect 147 2596 173 2603
rect 507 2596 583 2603
rect 107 2576 203 2583
rect 196 2567 203 2576
rect 307 2573 312 2587
rect 348 2576 523 2583
rect 516 2567 523 2576
rect 576 2567 583 2596
rect 867 2593 873 2607
rect 1416 2600 1693 2603
rect 1413 2596 1693 2600
rect 1413 2587 1427 2596
rect 1707 2596 1773 2603
rect 1887 2596 1973 2603
rect 2147 2596 2233 2603
rect 2447 2596 2553 2603
rect 3367 2596 3453 2603
rect 3527 2596 3633 2603
rect 4187 2596 4573 2603
rect 4936 2600 5353 2603
rect 4933 2596 5353 2600
rect 696 2580 753 2583
rect 693 2576 753 2580
rect 693 2567 707 2576
rect 807 2573 813 2587
rect 947 2576 1153 2583
rect 1387 2576 1413 2583
rect 1527 2573 1533 2587
rect 1927 2573 1933 2587
rect 1947 2576 2063 2583
rect 2156 2580 2193 2583
rect 1773 2567 1787 2573
rect 93 2547 107 2553
rect 206 2553 207 2560
rect 133 2547 147 2553
rect 193 2547 207 2553
rect 147 2536 172 2543
rect 206 2540 207 2547
rect 213 2553 214 2560
rect 287 2556 312 2563
rect 348 2560 383 2563
rect 348 2556 387 2560
rect 213 2547 227 2553
rect 373 2547 387 2556
rect 407 2556 473 2563
rect 487 2553 493 2567
rect 516 2556 533 2567
rect 520 2553 533 2556
rect 627 2553 633 2567
rect 1147 2553 1152 2567
rect 1188 2556 1313 2563
rect 1656 2560 1733 2563
rect 1033 2547 1047 2553
rect 1613 2547 1627 2553
rect 213 2540 214 2547
rect 248 2536 333 2543
rect 427 2533 433 2547
rect 447 2536 513 2543
rect 553 2527 567 2533
rect 47 2513 53 2527
rect 127 2516 213 2523
rect 227 2516 333 2523
rect 673 2527 687 2533
rect 867 2536 913 2543
rect 1087 2536 1133 2543
rect 1207 2536 1293 2543
rect 1427 2533 1433 2547
rect 1507 2533 1513 2547
rect 1653 2556 1733 2560
rect 1653 2547 1667 2556
rect 1747 2553 1752 2567
rect 1773 2560 1774 2567
rect 1827 2553 1833 2567
rect 2056 2547 2063 2576
rect 2153 2576 2193 2580
rect 2153 2567 2167 2576
rect 2287 2576 2313 2583
rect 2513 2567 2527 2573
rect 2107 2553 2113 2567
rect 2166 2560 2167 2567
rect 2173 2553 2174 2560
rect 2188 2556 2253 2563
rect 2347 2553 2353 2567
rect 2367 2556 2413 2563
rect 2716 2580 2753 2583
rect 2573 2567 2587 2573
rect 2713 2576 2753 2580
rect 2713 2567 2727 2576
rect 2767 2576 3003 2583
rect 2996 2567 3003 2576
rect 3396 2576 3533 2583
rect 2926 2553 2927 2560
rect 2967 2553 2973 2567
rect 2996 2556 3013 2567
rect 3000 2553 3013 2556
rect 3087 2553 3093 2567
rect 3306 2553 3307 2560
rect 3396 2563 3403 2576
rect 3593 2567 3607 2573
rect 3328 2556 3403 2563
rect 3427 2553 3433 2567
rect 4087 2580 4122 2583
rect 4296 2580 4413 2583
rect 4087 2576 4127 2580
rect 3633 2567 3647 2573
rect 4113 2567 4127 2576
rect 4293 2576 4413 2580
rect 4293 2567 4307 2576
rect 4933 2587 4947 2596
rect 5416 2596 5453 2603
rect 4467 2576 4523 2583
rect 4516 2567 4523 2576
rect 4807 2573 4813 2587
rect 5056 2576 5273 2583
rect 3687 2556 3733 2563
rect 3847 2553 3853 2567
rect 3907 2553 3913 2567
rect 3956 2556 4053 2563
rect 2173 2547 2187 2553
rect 2453 2547 2467 2553
rect 1747 2533 1753 2547
rect 1807 2533 1813 2547
rect 2007 2533 2013 2547
rect 2147 2533 2152 2547
rect 2173 2540 2174 2547
rect 2307 2533 2313 2547
rect 2567 2536 2593 2543
rect 2873 2543 2887 2553
rect 2913 2547 2927 2553
rect 3133 2547 3147 2553
rect 2827 2540 2887 2543
rect 2827 2536 2883 2540
rect 2906 2533 2907 2540
rect 2926 2540 2927 2547
rect 2948 2536 2993 2543
rect 3293 2547 3307 2553
rect 3956 2547 3963 2556
rect 4067 2556 4092 2563
rect 4126 2560 4127 2567
rect 4146 2553 4147 2560
rect 4168 2556 4212 2563
rect 4248 2553 4253 2567
rect 4347 2556 4393 2563
rect 4133 2547 4147 2553
rect 4467 2560 4503 2563
rect 4467 2556 4507 2560
rect 4516 2556 4533 2567
rect 4493 2547 4507 2556
rect 4520 2553 4533 2556
rect 4707 2556 4733 2563
rect 5056 2563 5063 2576
rect 5416 2583 5423 2596
rect 5527 2596 5553 2603
rect 5647 2596 5673 2603
rect 5347 2576 5423 2583
rect 5376 2567 5383 2576
rect 5433 2567 5447 2573
rect 5567 2576 5693 2583
rect 5027 2556 5063 2563
rect 5087 2556 5113 2563
rect 5227 2556 5293 2563
rect 5347 2553 5353 2567
rect 5376 2556 5393 2567
rect 5380 2553 5393 2556
rect 5487 2563 5500 2567
rect 5487 2553 5503 2563
rect 5527 2556 5653 2563
rect 3387 2536 3412 2543
rect 3448 2533 3453 2547
rect 3547 2536 3573 2543
rect 3667 2536 3713 2543
rect 3767 2536 3793 2543
rect 3887 2536 3923 2543
rect 713 2527 727 2533
rect 807 2516 833 2523
rect 887 2513 893 2527
rect 1027 2516 1053 2523
rect 1267 2513 1273 2527
rect 1567 2513 1573 2527
rect 1736 2523 1743 2533
rect 1647 2516 1743 2523
rect 1787 2516 1873 2523
rect 1927 2516 1973 2523
rect 2047 2513 2053 2527
rect 2687 2516 2873 2523
rect 2893 2523 2907 2533
rect 2887 2520 2907 2523
rect 2887 2516 2902 2520
rect 3333 2523 3347 2533
rect 3267 2520 3347 2523
rect 3267 2516 3343 2520
rect 3367 2516 3452 2523
rect 3488 2516 3553 2523
rect 3613 2523 3627 2533
rect 3613 2520 3673 2523
rect 3616 2516 3673 2520
rect 3916 2523 3923 2536
rect 3947 2536 3963 2547
rect 3947 2533 3960 2536
rect 4007 2533 4013 2547
rect 4187 2533 4193 2547
rect 4287 2533 4292 2547
rect 4313 2533 4314 2540
rect 4427 2536 4453 2543
rect 4587 2536 4713 2543
rect 4787 2533 4793 2547
rect 4887 2536 4913 2543
rect 5167 2536 5273 2543
rect 4313 2527 4327 2533
rect 3916 2516 3993 2523
rect 4047 2516 4073 2523
rect 4313 2520 4314 2527
rect 4396 2516 4473 2523
rect 393 2507 407 2513
rect 687 2496 913 2503
rect 933 2503 947 2513
rect 1313 2507 1327 2513
rect 933 2500 1033 2503
rect 936 2496 1033 2500
rect 1047 2496 1193 2503
rect 1547 2496 1893 2503
rect 1967 2496 2093 2503
rect 2167 2496 2293 2503
rect 2316 2496 2633 2503
rect 313 2487 327 2493
rect 507 2476 753 2483
rect 907 2476 993 2483
rect 2316 2483 2323 2496
rect 3247 2496 3433 2503
rect 3447 2496 3693 2503
rect 4147 2496 4183 2503
rect 1087 2476 2323 2483
rect 2467 2476 2813 2483
rect 3267 2476 3413 2483
rect 4107 2476 4153 2483
rect 4176 2483 4183 2496
rect 4396 2503 4403 2516
rect 4627 2516 4673 2523
rect 4687 2513 4693 2527
rect 4747 2516 4853 2523
rect 5146 2513 5147 2520
rect 5168 2513 5173 2527
rect 5313 2523 5327 2533
rect 5467 2533 5473 2547
rect 5496 2543 5503 2553
rect 5496 2536 5573 2543
rect 5313 2520 5393 2523
rect 5316 2516 5393 2520
rect 5413 2523 5427 2533
rect 5413 2520 5513 2523
rect 5416 2516 5513 2520
rect 5607 2516 5633 2523
rect 5647 2516 5673 2523
rect 4287 2496 4403 2503
rect 4427 2496 4473 2503
rect 4487 2496 4553 2503
rect 4727 2496 4753 2503
rect 4907 2496 4973 2503
rect 5133 2503 5147 2513
rect 5107 2500 5147 2503
rect 5553 2503 5567 2513
rect 5553 2500 5613 2503
rect 5107 2496 5142 2500
rect 5556 2496 5613 2500
rect 5627 2496 5693 2503
rect 4176 2476 4433 2483
rect 4507 2476 4633 2483
rect 4747 2476 5633 2483
rect 1267 2456 1433 2463
rect 1747 2456 1853 2463
rect 2047 2456 2193 2463
rect 2820 2466 2833 2467
rect 2827 2453 2833 2466
rect 3327 2456 3373 2463
rect 3827 2456 4013 2463
rect 4027 2456 4873 2463
rect 5076 2456 5153 2463
rect 107 2436 173 2443
rect 767 2433 773 2447
rect 887 2436 973 2443
rect 1207 2433 1213 2447
rect 1427 2436 1953 2443
rect 2487 2436 2733 2443
rect 2913 2443 2927 2453
rect 2913 2440 3133 2443
rect 2916 2436 3133 2440
rect 3227 2436 3513 2443
rect 3747 2436 3813 2443
rect 4187 2436 4213 2443
rect 4327 2436 4513 2443
rect 4647 2436 4673 2443
rect 5076 2443 5083 2456
rect 5327 2456 5473 2463
rect 5527 2453 5533 2467
rect 5707 2453 5713 2467
rect 4887 2436 5083 2443
rect 5256 2436 5333 2443
rect 507 2416 833 2423
rect 847 2416 973 2423
rect 2507 2416 3393 2423
rect 3507 2416 3753 2423
rect 4267 2416 4713 2423
rect 5256 2423 5263 2436
rect 4787 2416 5263 2423
rect 5287 2416 5633 2423
rect 267 2396 453 2403
rect 667 2396 913 2403
rect 1607 2396 1673 2403
rect 2887 2396 2913 2403
rect 3107 2396 3712 2403
rect 3748 2396 3913 2403
rect 4287 2396 4533 2403
rect 4707 2396 5053 2403
rect 5096 2396 5213 2403
rect 547 2376 693 2383
rect 707 2376 903 2383
rect 896 2367 903 2376
rect 1167 2376 1673 2383
rect 1767 2376 1813 2383
rect 1893 2383 1907 2393
rect 1893 2380 2673 2383
rect 1896 2376 2673 2380
rect 3327 2376 3653 2383
rect 3827 2376 3853 2383
rect 4007 2376 4053 2383
rect 4307 2376 4373 2383
rect 5096 2383 5103 2396
rect 5507 2396 5713 2403
rect 4627 2376 5103 2383
rect 5167 2376 5313 2383
rect 5387 2376 5453 2383
rect 5647 2376 5673 2383
rect 447 2356 553 2363
rect 567 2356 793 2363
rect 907 2356 1393 2363
rect 2356 2356 2513 2363
rect 2356 2348 2363 2356
rect 2567 2356 2593 2363
rect 2887 2356 3173 2363
rect 3687 2356 3773 2363
rect 3907 2356 3993 2363
rect 4007 2356 4093 2363
rect 4147 2356 4333 2363
rect 4427 2356 4613 2363
rect 4847 2356 4933 2363
rect 5436 2356 5713 2363
rect 527 2336 573 2343
rect 587 2336 853 2343
rect 1247 2336 1653 2343
rect 2007 2336 2133 2343
rect 2187 2336 2353 2343
rect 2927 2336 3053 2343
rect 3067 2336 3313 2343
rect 3447 2336 3973 2343
rect 3987 2336 4153 2343
rect 4227 2336 4353 2343
rect 4447 2336 4553 2343
rect 4567 2336 4673 2343
rect 4727 2336 5043 2343
rect 5036 2327 5043 2336
rect 5207 2336 5353 2343
rect 5436 2343 5443 2356
rect 5367 2336 5443 2343
rect 5467 2336 5552 2343
rect 5588 2336 5673 2343
rect 167 2316 404 2323
rect 67 2293 72 2307
rect 108 2294 113 2307
rect 100 2293 113 2294
rect 147 2273 153 2287
rect 207 2274 213 2287
rect 200 2273 213 2274
rect 267 2276 313 2283
rect 397 2287 404 2316
rect 627 2316 772 2323
rect 786 2313 787 2320
rect 808 2323 820 2327
rect 960 2323 973 2327
rect 808 2320 823 2323
rect 808 2313 827 2320
rect 773 2307 787 2313
rect 507 2296 533 2303
rect 556 2300 713 2303
rect 553 2296 713 2300
rect 553 2287 567 2296
rect 727 2303 740 2307
rect 727 2293 743 2303
rect 813 2307 827 2313
rect 956 2313 973 2323
rect 1047 2316 1173 2323
rect 1196 2316 1233 2323
rect 913 2293 914 2300
rect 327 2276 352 2283
rect 386 2273 387 2280
rect 500 2286 513 2287
rect 93 2267 107 2273
rect 373 2267 387 2273
rect 507 2273 513 2286
rect 627 2273 632 2287
rect 736 2287 743 2293
rect 913 2287 927 2293
rect 956 2287 963 2313
rect 1007 2296 1033 2303
rect 1196 2303 1203 2316
rect 1107 2296 1203 2303
rect 1233 2307 1247 2313
rect 1327 2316 1513 2323
rect 1567 2316 1773 2323
rect 1836 2316 1903 2323
rect 1313 2307 1327 2313
rect 1367 2293 1373 2307
rect 1507 2296 1613 2303
rect 1836 2303 1843 2316
rect 1627 2296 1843 2303
rect 1493 2287 1507 2293
rect 1753 2287 1767 2296
rect 1896 2287 1903 2316
rect 1976 2316 2353 2323
rect 1976 2307 1983 2316
rect 2407 2316 2433 2323
rect 2527 2320 2603 2323
rect 2527 2316 2607 2320
rect 1917 2296 1972 2303
rect 668 2274 672 2287
rect 660 2273 672 2274
rect 693 2273 694 2280
rect 736 2276 753 2287
rect 740 2273 753 2276
rect 913 2280 914 2287
rect 906 2273 907 2280
rect 1047 2276 1073 2283
rect 1127 2273 1133 2287
rect 1187 2276 1213 2283
rect 1347 2273 1353 2287
rect 1447 2273 1453 2287
rect 1707 2273 1713 2287
rect 1827 2276 1853 2283
rect 693 2267 707 2273
rect 207 2256 233 2263
rect 320 2266 333 2267
rect 287 2256 313 2263
rect 327 2253 333 2266
rect 386 2260 387 2267
rect 667 2253 672 2267
rect 693 2260 694 2267
rect 793 2263 807 2273
rect 893 2267 907 2273
rect 1253 2267 1267 2273
rect 1613 2267 1627 2273
rect 1853 2267 1867 2273
rect 1917 2267 1924 2296
rect 1993 2293 1994 2300
rect 2067 2296 2133 2303
rect 2187 2294 2193 2307
rect 2593 2307 2607 2316
rect 2747 2316 2933 2323
rect 3387 2316 3563 2323
rect 2187 2293 2200 2294
rect 2447 2296 2493 2303
rect 2587 2293 2593 2307
rect 2667 2293 2673 2307
rect 3136 2300 3233 2303
rect 3133 2296 3233 2300
rect 1993 2287 2007 2293
rect 3133 2287 3147 2296
rect 3287 2296 3433 2303
rect 3520 2303 3533 2307
rect 3517 2293 3533 2303
rect 3556 2303 3563 2316
rect 3667 2316 3733 2323
rect 3906 2313 3907 2320
rect 3928 2316 4073 2323
rect 4087 2316 4113 2323
rect 4207 2316 4233 2323
rect 3893 2307 3907 2313
rect 4413 2307 4427 2313
rect 4767 2316 4833 2323
rect 5047 2316 5173 2323
rect 5187 2316 5373 2323
rect 5447 2316 5633 2323
rect 4613 2307 4627 2313
rect 3556 2296 3613 2303
rect 1947 2276 1993 2283
rect 2047 2276 2153 2283
rect 2167 2276 2193 2283
rect 2387 2276 2413 2283
rect 2607 2273 2613 2287
rect 2827 2273 2833 2287
rect 2987 2276 3093 2283
rect 2273 2267 2287 2273
rect 793 2260 853 2263
rect 796 2256 853 2260
rect 920 2263 933 2267
rect 916 2253 933 2263
rect 1527 2256 1553 2263
rect 1567 2253 1573 2267
rect 1667 2256 1733 2263
rect 1866 2260 1867 2267
rect 1888 2253 1892 2267
rect 1967 2253 1973 2267
rect 2000 2263 2013 2267
rect 1996 2253 2013 2263
rect 2273 2263 2292 2267
rect 2067 2256 2292 2263
rect 2280 2253 2292 2256
rect 2328 2253 2333 2267
rect 2493 2263 2507 2273
rect 2713 2267 2727 2273
rect 3493 2267 3507 2273
rect 3517 2267 3524 2293
rect 3853 2287 3867 2293
rect 3973 2287 3987 2293
rect 4127 2296 4313 2303
rect 4367 2293 4373 2307
rect 4113 2287 4127 2293
rect 4513 2287 4527 2293
rect 3607 2276 3712 2283
rect 3748 2273 3753 2287
rect 3866 2280 3867 2287
rect 3888 2273 3893 2287
rect 4167 2273 4173 2287
rect 4187 2280 4242 2283
rect 4187 2276 4247 2280
rect 2347 2260 2507 2263
rect 2347 2256 2503 2260
rect 2787 2256 2853 2263
rect 2927 2256 2953 2263
rect 3047 2256 3072 2263
rect 3108 2253 3113 2267
rect 3167 2253 3173 2267
rect 3287 2256 3372 2263
rect 3408 2256 3433 2263
rect 3506 2260 3507 2267
rect 3533 2263 3547 2273
rect 3533 2260 3693 2263
rect 3536 2256 3693 2260
rect 3747 2256 3813 2263
rect 3927 2256 3953 2263
rect 3980 2263 3993 2267
rect 3976 2253 3993 2263
rect 4013 2263 4027 2273
rect 4233 2267 4247 2276
rect 4407 2280 4502 2283
rect 4407 2276 4507 2280
rect 4493 2267 4507 2276
rect 4636 2296 4713 2303
rect 4553 2287 4567 2293
rect 4636 2267 4643 2296
rect 4867 2293 4873 2307
rect 4987 2296 5213 2303
rect 4667 2274 4672 2287
rect 4813 2287 4827 2293
rect 5073 2287 5087 2296
rect 5275 2300 5313 2303
rect 5273 2296 5313 2300
rect 5273 2287 5287 2296
rect 5427 2303 5440 2307
rect 5427 2300 5443 2303
rect 5427 2293 5447 2300
rect 5547 2300 5583 2303
rect 5547 2296 5587 2300
rect 5433 2287 5447 2293
rect 5573 2287 5587 2296
rect 4667 2273 4680 2274
rect 4708 2276 4773 2283
rect 4826 2280 4827 2287
rect 4848 2273 4853 2287
rect 4927 2276 4953 2283
rect 5127 2276 5153 2283
rect 5247 2273 5252 2287
rect 5286 2280 5287 2287
rect 5308 2276 5393 2283
rect 5507 2283 5520 2287
rect 5507 2280 5522 2283
rect 5507 2273 5527 2280
rect 4013 2260 4073 2263
rect 4016 2256 4073 2260
rect 4087 2256 4133 2263
rect 4246 2260 4247 2267
rect 4266 2253 4267 2260
rect 4288 2256 4313 2263
rect 4506 2260 4507 2267
rect 4520 2266 4533 2267
rect 916 2243 923 2253
rect 847 2236 923 2243
rect 1067 2236 1153 2243
rect 1473 2243 1487 2253
rect 1773 2247 1787 2253
rect 1367 2240 1487 2243
rect 1367 2236 1483 2240
rect 1527 2236 1593 2243
rect 1996 2243 2003 2253
rect 1827 2236 2003 2243
rect 2513 2247 2527 2253
rect 2967 2233 2973 2247
rect 2993 2243 3007 2253
rect 2993 2240 3053 2243
rect 2996 2236 3053 2240
rect 3693 2247 3707 2253
rect 3247 2234 3253 2247
rect 3240 2233 3253 2234
rect 3387 2236 3413 2243
rect 3507 2236 3533 2243
rect 3620 2243 3633 2247
rect 3616 2233 3633 2243
rect 3976 2243 3983 2253
rect 3867 2236 3983 2243
rect 4047 2236 4093 2243
rect 807 2216 1413 2223
rect 2887 2216 3233 2223
rect 2553 2207 2567 2213
rect 3616 2223 3623 2233
rect 4176 2227 4183 2253
rect 4253 2247 4267 2253
rect 4528 2253 4533 2266
rect 4727 2256 4753 2263
rect 4827 2256 4913 2263
rect 4987 2253 4993 2267
rect 5007 2253 5012 2267
rect 5048 2253 5052 2267
rect 5513 2267 5527 2273
rect 5533 2267 5547 2273
rect 5088 2254 5093 2267
rect 5080 2253 5093 2254
rect 5187 2256 5213 2263
rect 5307 2253 5313 2267
rect 5367 2256 5413 2263
rect 5467 2253 5473 2267
rect 5526 2260 5527 2267
rect 5546 2260 5547 2267
rect 5568 2253 5573 2267
rect 4266 2240 4267 2247
rect 4573 2247 4587 2253
rect 4673 2247 4687 2253
rect 4847 2236 4953 2243
rect 5133 2243 5147 2253
rect 5253 2247 5267 2253
rect 5087 2240 5147 2243
rect 5087 2236 5143 2240
rect 5247 2240 5267 2247
rect 5247 2236 5263 2240
rect 5247 2233 5260 2236
rect 5347 2236 5453 2243
rect 5516 2243 5523 2253
rect 5516 2236 5563 2243
rect 3447 2216 3623 2223
rect 3647 2216 3933 2223
rect 4176 2216 4193 2227
rect 4180 2213 4193 2216
rect 4347 2216 4553 2223
rect 4667 2216 4913 2223
rect 5047 2216 5173 2223
rect 5487 2216 5533 2223
rect 4073 2207 4087 2213
rect 327 2196 453 2203
rect 767 2196 1573 2203
rect 1867 2196 2213 2203
rect 2227 2193 2233 2207
rect 2767 2196 2833 2203
rect 3207 2196 3473 2203
rect 3487 2196 3833 2203
rect 4047 2193 4052 2207
rect 4073 2200 4074 2207
rect 4507 2196 4773 2203
rect 4787 2196 5133 2203
rect 5267 2196 5353 2203
rect 5556 2203 5563 2236
rect 5407 2196 5563 2203
rect 5613 2187 5627 2193
rect 1267 2176 1433 2183
rect 1447 2176 2373 2183
rect 2487 2176 2513 2183
rect 2927 2176 2953 2183
rect 2967 2176 3413 2183
rect 3527 2176 3703 2183
rect 1213 2167 1227 2173
rect 1213 2160 1233 2167
rect 1216 2156 1233 2160
rect 1220 2153 1233 2156
rect 1287 2156 1353 2163
rect 1987 2156 2073 2163
rect 2476 2163 2483 2173
rect 3696 2167 3703 2176
rect 3767 2176 4113 2183
rect 4167 2176 4993 2183
rect 5247 2176 5413 2183
rect 2087 2156 2483 2163
rect 3387 2156 3653 2163
rect 3707 2156 3913 2163
rect 3987 2156 4013 2163
rect 4067 2156 4453 2163
rect 4567 2156 4673 2163
rect 4687 2156 4852 2163
rect 4888 2156 4913 2163
rect 4956 2156 5133 2163
rect 3313 2147 3327 2153
rect 47 2136 113 2143
rect 447 2133 453 2147
rect 1667 2136 1893 2143
rect 2027 2136 2813 2143
rect 3107 2136 3273 2143
rect 3607 2136 4153 2143
rect 4287 2133 4293 2147
rect 2933 2127 2947 2133
rect 4467 2136 4613 2143
rect 4667 2133 4673 2147
rect 4956 2143 4963 2156
rect 4827 2136 4963 2143
rect 4976 2136 5303 2143
rect 87 2116 153 2123
rect 247 2116 373 2123
rect 427 2116 713 2123
rect 727 2116 953 2123
rect 1167 2116 1273 2123
rect 1507 2116 1713 2123
rect 2107 2116 2253 2123
rect 2447 2116 2513 2123
rect 3227 2116 3333 2123
rect 3727 2116 3813 2123
rect 3986 2113 3987 2120
rect 4008 2116 4223 2123
rect 113 2093 114 2100
rect 236 2103 243 2113
rect 187 2096 243 2103
rect 696 2100 793 2103
rect 693 2096 793 2100
rect 113 2087 127 2093
rect 87 2073 92 2087
rect 113 2080 114 2087
rect 128 2080 204 2083
rect 128 2076 207 2080
rect 193 2067 207 2076
rect 287 2076 333 2083
rect 407 2074 413 2087
rect 693 2087 707 2096
rect 867 2096 993 2103
rect 1127 2096 1183 2103
rect 407 2073 420 2074
rect 467 2076 513 2083
rect 567 2073 573 2087
rect 1176 2083 1183 2096
rect 1347 2096 1433 2103
rect 1447 2093 1453 2107
rect 1596 2100 1653 2103
rect 1553 2087 1567 2093
rect 1176 2076 1383 2083
rect 233 2067 247 2073
rect 1153 2067 1167 2073
rect 47 2056 93 2063
rect 147 2056 172 2063
rect 193 2060 194 2067
rect 307 2056 372 2063
rect 408 2053 413 2067
rect 287 2036 473 2043
rect 493 2043 507 2053
rect 487 2040 507 2043
rect 666 2053 667 2060
rect 688 2056 773 2063
rect 847 2056 893 2063
rect 967 2056 1033 2063
rect 1193 2067 1207 2076
rect 1376 2067 1383 2076
rect 1507 2073 1513 2087
rect 1593 2096 1653 2100
rect 1593 2087 1607 2096
rect 1667 2096 1693 2103
rect 1827 2103 1840 2107
rect 1827 2100 1843 2103
rect 1827 2093 1847 2100
rect 1887 2096 1983 2103
rect 1833 2087 1847 2093
rect 1727 2076 1793 2083
rect 1887 2073 1893 2087
rect 1976 2067 1983 2096
rect 2073 2087 2087 2093
rect 2256 2103 2263 2113
rect 3973 2107 3987 2113
rect 2256 2096 2503 2103
rect 2113 2087 2127 2093
rect 2467 2073 2473 2087
rect 2496 2067 2503 2096
rect 2767 2096 2813 2103
rect 3027 2096 3133 2103
rect 3147 2096 3363 2103
rect 2527 2073 2533 2087
rect 2587 2076 2613 2083
rect 2687 2073 2693 2087
rect 3047 2076 3093 2083
rect 3107 2074 3112 2087
rect 3356 2087 3363 2096
rect 3600 2103 3613 2107
rect 3447 2096 3613 2103
rect 3596 2093 3613 2096
rect 3667 2093 3673 2107
rect 4027 2096 4053 2103
rect 3107 2073 3120 2074
rect 3148 2076 3343 2083
rect 3356 2076 3373 2087
rect 3336 2067 3343 2076
rect 3360 2073 3373 2076
rect 3507 2073 3512 2087
rect 3548 2073 3553 2087
rect 3596 2083 3603 2093
rect 3596 2076 3633 2083
rect 3647 2076 3792 2083
rect 3828 2076 3953 2083
rect 4187 2073 4193 2087
rect 4216 2067 4223 2116
rect 4976 2127 4983 2136
rect 4447 2116 4493 2123
rect 4587 2116 4713 2123
rect 4736 2116 4973 2123
rect 4296 2096 4433 2103
rect 4247 2073 4253 2087
rect 4296 2067 4303 2096
rect 4736 2103 4743 2116
rect 5107 2116 5233 2123
rect 5296 2123 5303 2136
rect 5327 2136 5373 2143
rect 5473 2143 5487 2153
rect 5473 2140 5613 2143
rect 5476 2136 5613 2140
rect 5296 2116 5332 2123
rect 5368 2116 5453 2123
rect 5527 2116 5593 2123
rect 4536 2096 4743 2103
rect 4536 2087 4543 2096
rect 4767 2096 4813 2103
rect 5036 2100 5123 2103
rect 5033 2096 5123 2100
rect 5033 2087 5047 2096
rect 5116 2087 5123 2096
rect 5567 2096 5713 2103
rect 4327 2073 4333 2087
rect 4387 2076 4413 2083
rect 4487 2076 4513 2083
rect 4527 2076 4543 2087
rect 4527 2073 4540 2076
rect 4567 2073 4573 2087
rect 4627 2076 4713 2083
rect 4827 2073 4833 2087
rect 4967 2076 4993 2083
rect 5080 2083 5093 2087
rect 5076 2073 5093 2083
rect 5116 2076 5133 2087
rect 5120 2073 5133 2076
rect 5187 2076 5232 2083
rect 5268 2073 5272 2087
rect 5293 2073 5294 2080
rect 5347 2076 5453 2083
rect 5467 2076 5513 2083
rect 1287 2053 1293 2067
rect 1347 2053 1353 2067
rect 1376 2056 1393 2067
rect 1380 2053 1393 2056
rect 1487 2056 1513 2063
rect 1527 2053 1533 2067
rect 1687 2053 1693 2067
rect 1767 2056 1813 2063
rect 1827 2053 1832 2067
rect 1853 2053 1854 2060
rect 2027 2053 2033 2067
rect 533 2047 547 2053
rect 487 2036 503 2040
rect 653 2043 667 2053
rect 653 2040 733 2043
rect 655 2036 733 2040
rect 747 2033 753 2047
rect 807 2033 813 2047
rect 867 2033 873 2047
rect 213 2023 227 2033
rect 47 2020 227 2023
rect 913 2027 927 2033
rect 47 2016 223 2020
rect 1067 2033 1073 2047
rect 1100 2043 1113 2047
rect 1096 2033 1113 2043
rect 1187 2036 1313 2043
rect 1327 2046 1340 2047
rect 1327 2033 1333 2046
rect 1013 2023 1027 2033
rect 1096 2023 1103 2033
rect 1573 2043 1587 2053
rect 1573 2040 1633 2043
rect 1576 2036 1633 2040
rect 1647 2036 1672 2043
rect 1708 2033 1713 2047
rect 1853 2043 1867 2053
rect 2093 2047 2107 2053
rect 1853 2040 1893 2043
rect 1857 2036 1893 2040
rect 1967 2033 1972 2047
rect 2008 2043 2020 2047
rect 2008 2033 2023 2043
rect 2267 2056 2373 2063
rect 2427 2053 2433 2067
rect 2547 2056 2593 2063
rect 2647 2053 2653 2067
rect 2727 2056 2792 2063
rect 2828 2056 2873 2063
rect 2947 2056 2993 2063
rect 3100 2066 3113 2067
rect 2133 2047 2147 2053
rect 3107 2053 3113 2066
rect 3167 2056 3252 2063
rect 3273 2053 3274 2060
rect 3336 2056 3353 2067
rect 3340 2053 3353 2056
rect 3407 2053 3413 2067
rect 3273 2047 3287 2053
rect 2227 2033 2233 2047
rect 2407 2036 2733 2043
rect 2867 2036 2973 2043
rect 2987 2033 2993 2047
rect 3227 2033 3233 2047
rect 3513 2047 3527 2053
rect 3607 2056 3793 2063
rect 3847 2053 3853 2067
rect 3906 2053 3907 2060
rect 3928 2053 3933 2067
rect 4047 2053 4052 2067
rect 4088 2053 4093 2067
rect 4107 2056 4173 2063
rect 4296 2056 4313 2067
rect 4300 2053 4313 2056
rect 4367 2056 4413 2063
rect 4487 2053 4493 2067
rect 4547 2056 4593 2063
rect 4647 2056 4733 2063
rect 4887 2056 4973 2063
rect 5027 2056 5053 2063
rect 3553 2043 3567 2053
rect 3893 2047 3907 2053
rect 3553 2040 3593 2043
rect 3556 2036 3593 2040
rect 1013 2020 1103 2023
rect 1016 2016 1103 2020
rect 2016 2023 2023 2033
rect 2016 2016 2112 2023
rect 2148 2016 2273 2023
rect 2787 2016 3013 2023
rect 3247 2016 3373 2023
rect 3556 2020 3563 2036
rect 3747 2033 3753 2047
rect 3827 2046 3840 2047
rect 3827 2033 3833 2046
rect 4047 2043 4060 2047
rect 4047 2033 4063 2043
rect 4087 2036 4153 2043
rect 4207 2036 4373 2043
rect 4687 2036 4713 2043
rect 4767 2036 4792 2043
rect 4828 2036 4852 2043
rect 4888 2033 4892 2047
rect 5076 2043 5083 2073
rect 5293 2067 5307 2073
rect 5553 2067 5567 2073
rect 5127 2053 5132 2067
rect 5153 2053 5154 2060
rect 5367 2056 5413 2063
rect 5567 2053 5573 2067
rect 4928 2036 5083 2043
rect 5153 2043 5167 2053
rect 5253 2043 5267 2053
rect 5673 2047 5687 2053
rect 5153 2040 5203 2043
rect 5253 2040 5333 2043
rect 5157 2036 5203 2040
rect 5256 2036 5333 2040
rect 587 1996 833 2003
rect 927 1996 1233 2003
rect 1587 1996 1673 2003
rect 1907 1996 1993 2003
rect 2276 2003 2283 2013
rect 3553 2007 3567 2020
rect 3588 2016 3633 2023
rect 2276 1996 2673 2003
rect 2827 1996 2853 2003
rect 2867 1993 2873 2007
rect 3936 2003 3943 2033
rect 3973 2027 3987 2033
rect 4056 2023 4063 2033
rect 4056 2016 4253 2023
rect 4347 2016 4573 2023
rect 4667 2016 4813 2023
rect 4867 2016 5173 2023
rect 5196 2023 5203 2036
rect 5347 2033 5353 2047
rect 5547 2036 5633 2043
rect 5196 2016 5293 2023
rect 5307 2016 5613 2023
rect 5667 2016 5693 2023
rect 3936 1996 4033 2003
rect 4187 1996 4313 2003
rect 4487 1996 4593 2003
rect 4687 1993 4693 2007
rect 5147 1993 5152 2007
rect 1896 1983 1903 1993
rect 5188 1996 5213 2003
rect 5227 1996 5353 2003
rect 5647 1996 5693 2003
rect 1527 1976 1903 1983
rect 2487 1976 2513 1983
rect 2867 1976 3113 1983
rect 3167 1976 3313 1983
rect 3727 1976 3993 1983
rect 4127 1976 4173 1983
rect 4287 1973 4293 1987
rect 4547 1976 4803 1983
rect 387 1956 453 1963
rect 567 1956 593 1963
rect 1707 1956 2073 1963
rect 2087 1956 2313 1963
rect 2507 1956 2813 1963
rect 2947 1956 3133 1963
rect 3187 1956 3313 1963
rect 3467 1956 3673 1963
rect 3847 1956 4113 1963
rect 4287 1956 4393 1963
rect 4433 1963 4447 1973
rect 4796 1967 4803 1976
rect 4867 1976 5033 1983
rect 5567 1976 5613 1983
rect 5667 1973 5673 1987
rect 4433 1960 4783 1963
rect 4436 1956 4783 1960
rect 247 1936 673 1943
rect 700 1943 713 1947
rect 696 1940 713 1943
rect 693 1933 713 1940
rect 1807 1936 2233 1943
rect 2707 1936 2913 1943
rect 3007 1936 3233 1943
rect 3287 1936 4013 1943
rect 4056 1936 4413 1943
rect 693 1927 707 1933
rect 107 1916 333 1923
rect 347 1916 533 1923
rect 587 1916 653 1923
rect 747 1916 1553 1923
rect 2067 1916 2113 1923
rect 2127 1916 2933 1923
rect 3047 1916 3353 1923
rect 4056 1923 4063 1936
rect 4776 1943 4783 1956
rect 4807 1956 5633 1963
rect 5680 1966 5693 1967
rect 5687 1953 5693 1966
rect 4776 1936 4893 1943
rect 4987 1936 5293 1943
rect 3427 1916 4063 1923
rect 4567 1916 4772 1923
rect 4808 1916 5073 1923
rect 5447 1916 5613 1923
rect 307 1896 413 1903
rect 427 1896 633 1903
rect 647 1896 753 1903
rect 1207 1896 1293 1903
rect 1947 1896 2053 1903
rect 2167 1896 2253 1903
rect 2307 1896 2353 1903
rect 3067 1896 3193 1903
rect 3247 1896 3513 1903
rect 3567 1893 3573 1907
rect 3727 1893 3733 1907
rect 3907 1896 4813 1903
rect 4907 1896 5133 1903
rect 5347 1896 5693 1903
rect 487 1876 653 1883
rect 667 1876 793 1883
rect 907 1876 1133 1883
rect 1747 1876 1953 1883
rect 2007 1876 2773 1883
rect 3147 1876 3413 1883
rect 3487 1876 3533 1883
rect 3687 1876 3713 1883
rect 4047 1876 4153 1883
rect 4427 1876 4673 1883
rect 4687 1876 4912 1883
rect 4948 1876 5113 1883
rect 5287 1873 5293 1887
rect 5487 1876 5512 1883
rect 5548 1873 5553 1887
rect 107 1856 293 1863
rect 307 1856 493 1863
rect 616 1856 913 1863
rect 87 1836 153 1843
rect 347 1836 433 1843
rect 616 1843 623 1856
rect 1527 1856 1752 1863
rect 1788 1856 1813 1863
rect 2167 1856 2413 1863
rect 2427 1856 2593 1863
rect 2847 1856 3113 1863
rect 3127 1856 3273 1863
rect 3407 1856 3773 1863
rect 4647 1856 4693 1863
rect 4787 1856 5193 1863
rect 5207 1856 5533 1863
rect 5547 1856 5713 1863
rect 487 1836 623 1843
rect 927 1836 1033 1843
rect 913 1827 927 1833
rect 1693 1827 1707 1833
rect 135 1820 193 1823
rect 133 1816 193 1820
rect 133 1807 147 1816
rect 207 1813 213 1827
rect 307 1820 364 1823
rect 307 1816 367 1820
rect 353 1807 367 1816
rect 627 1813 633 1827
rect 707 1816 743 1823
rect 493 1807 507 1813
rect 736 1807 743 1816
rect 767 1813 773 1827
rect 987 1813 993 1827
rect 1596 1820 1693 1823
rect 1593 1816 1693 1820
rect 1593 1807 1607 1816
rect 2347 1840 2603 1843
rect 2347 1836 2607 1840
rect 1733 1827 1747 1833
rect 2593 1827 2607 1836
rect 2947 1836 3153 1843
rect 3647 1836 3693 1843
rect 3716 1836 3892 1843
rect 3273 1827 3287 1833
rect 1887 1816 1953 1823
rect 2487 1816 2553 1823
rect 2647 1813 2653 1827
rect 2667 1816 2833 1823
rect 2887 1816 2913 1823
rect 3007 1816 3053 1823
rect 3206 1813 3207 1820
rect 3228 1813 3233 1827
rect 3347 1816 3433 1823
rect 3507 1816 3573 1823
rect 3587 1820 3662 1823
rect 3587 1816 3667 1820
rect 1993 1807 2007 1813
rect 107 1793 112 1807
rect 146 1800 147 1807
rect 168 1796 193 1803
rect 353 1800 354 1807
rect 346 1793 347 1800
rect 407 1793 413 1807
rect 547 1796 593 1803
rect 607 1793 613 1807
rect 667 1793 673 1807
rect 736 1803 753 1807
rect 696 1796 753 1803
rect 87 1773 92 1787
rect 126 1773 127 1780
rect 148 1776 193 1783
rect 233 1783 247 1793
rect 207 1780 247 1783
rect 333 1787 347 1793
rect 207 1776 243 1780
rect 447 1776 473 1783
rect 696 1783 703 1796
rect 740 1793 753 1796
rect 587 1776 703 1783
rect 793 1787 807 1793
rect 893 1787 907 1793
rect 1027 1793 1033 1807
rect 1167 1796 1193 1803
rect 1247 1796 1313 1803
rect 1340 1803 1353 1807
rect 1336 1793 1353 1803
rect 1407 1796 1453 1803
rect 1647 1796 1713 1803
rect 1807 1793 1813 1807
rect 1947 1796 1972 1803
rect 1993 1800 1994 1807
rect 2087 1793 2093 1807
rect 2147 1796 2193 1803
rect 2307 1796 2353 1803
rect 2407 1793 2413 1807
rect 2607 1793 2613 1807
rect 2807 1796 2852 1803
rect 2888 1796 2953 1803
rect 2967 1793 2973 1807
rect 3027 1793 3033 1807
rect 3153 1807 3167 1813
rect 3107 1794 3113 1807
rect 3100 1793 3113 1794
rect 3193 1803 3207 1813
rect 3653 1807 3667 1816
rect 3716 1823 3723 1836
rect 4107 1836 4273 1843
rect 4587 1836 4793 1843
rect 4927 1836 5013 1843
rect 3687 1816 3723 1823
rect 3827 1816 3873 1823
rect 3895 1807 3902 1833
rect 4056 1820 4133 1823
rect 4053 1816 4133 1820
rect 4053 1807 4067 1816
rect 4196 1820 4233 1823
rect 4193 1816 4233 1820
rect 4193 1807 4207 1816
rect 4507 1820 4583 1823
rect 4507 1816 4587 1820
rect 4573 1807 4587 1816
rect 4607 1816 4793 1823
rect 4653 1807 4667 1816
rect 4947 1816 5013 1823
rect 5053 1807 5067 1813
rect 3193 1800 3223 1803
rect 3195 1796 3223 1800
rect 933 1787 947 1793
rect 1073 1787 1087 1793
rect 1007 1776 1052 1783
rect 1073 1780 1074 1787
rect 1127 1773 1133 1787
rect 1227 1776 1263 1783
rect 113 1763 127 1773
rect 87 1760 127 1763
rect 373 1763 387 1773
rect 513 1767 527 1773
rect 1173 1767 1187 1773
rect 373 1760 473 1763
rect 87 1756 122 1760
rect 376 1756 473 1760
rect 887 1756 933 1763
rect 947 1756 1073 1763
rect 1256 1763 1263 1776
rect 1336 1783 1343 1793
rect 2233 1787 2247 1793
rect 2513 1787 2527 1793
rect 1287 1776 1343 1783
rect 1367 1773 1373 1787
rect 1547 1773 1553 1787
rect 1647 1776 1733 1783
rect 2007 1776 2113 1783
rect 2167 1773 2173 1787
rect 2287 1776 2313 1783
rect 2327 1776 2352 1783
rect 2386 1773 2387 1780
rect 2408 1776 2473 1783
rect 2733 1783 2747 1793
rect 2567 1780 2747 1783
rect 2567 1776 2743 1780
rect 2907 1773 2913 1787
rect 2967 1773 2973 1787
rect 3067 1776 3093 1783
rect 3120 1783 3133 1787
rect 1873 1767 1887 1773
rect 1256 1756 1293 1763
rect 1507 1756 1533 1763
rect 1886 1760 1887 1767
rect 1996 1763 2003 1773
rect 2373 1767 2387 1773
rect 3116 1773 3133 1783
rect 3187 1773 3193 1787
rect 1908 1756 2003 1763
rect 2016 1756 2253 1763
rect 427 1736 573 1743
rect 727 1736 893 1743
rect 907 1736 992 1743
rect 1028 1736 1133 1743
rect 1747 1736 1773 1743
rect 2016 1743 2023 1756
rect 2507 1756 2593 1763
rect 2767 1756 2793 1763
rect 2867 1756 2933 1763
rect 3007 1753 3012 1767
rect 3116 1763 3123 1773
rect 3048 1756 3123 1763
rect 3216 1763 3223 1796
rect 3247 1793 3253 1807
rect 3356 1800 3433 1803
rect 3353 1796 3433 1800
rect 3353 1787 3367 1796
rect 3587 1796 3613 1803
rect 3666 1800 3667 1807
rect 3673 1793 3674 1800
rect 3727 1796 3772 1803
rect 3808 1793 3813 1807
rect 3928 1793 3933 1807
rect 4115 1800 4193 1803
rect 3407 1774 3413 1787
rect 3436 1787 3443 1793
rect 3673 1787 3687 1793
rect 4093 1787 4107 1793
rect 4113 1796 4193 1800
rect 4113 1787 4127 1796
rect 4347 1793 4353 1807
rect 4407 1793 4413 1807
rect 4527 1793 4533 1807
rect 4587 1796 4643 1803
rect 4233 1787 4247 1793
rect 3407 1773 3420 1774
rect 3436 1773 3453 1787
rect 3647 1783 3660 1787
rect 3647 1773 3663 1783
rect 3747 1773 3752 1787
rect 3788 1773 3793 1787
rect 3907 1773 3913 1787
rect 3987 1776 4023 1783
rect 3436 1767 3443 1773
rect 3216 1756 3373 1763
rect 3420 1766 3443 1767
rect 3427 1756 3443 1766
rect 3427 1753 3440 1756
rect 3467 1756 3493 1763
rect 3656 1763 3663 1773
rect 3833 1767 3847 1773
rect 3656 1756 3823 1763
rect 1887 1736 2023 1743
rect 2747 1736 2793 1743
rect 3447 1746 3460 1747
rect 3447 1733 3453 1746
rect 3587 1736 3713 1743
rect 3816 1743 3823 1756
rect 4016 1763 4023 1776
rect 4047 1776 4072 1783
rect 4106 1780 4107 1787
rect 4126 1780 4127 1787
rect 4148 1776 4212 1783
rect 4246 1780 4247 1787
rect 4268 1776 4373 1783
rect 4447 1776 4472 1783
rect 4508 1776 4553 1783
rect 4607 1773 4613 1787
rect 4636 1783 4643 1796
rect 4666 1800 4667 1807
rect 4688 1793 4693 1807
rect 4927 1793 4933 1807
rect 4987 1793 4993 1807
rect 5147 1814 5153 1827
rect 5140 1813 5153 1814
rect 5247 1816 5272 1823
rect 5308 1820 5583 1823
rect 5308 1816 5587 1820
rect 5093 1807 5107 1813
rect 5573 1807 5587 1816
rect 5607 1823 5620 1827
rect 5607 1816 5673 1823
rect 5607 1813 5627 1816
rect 5147 1800 5243 1803
rect 5147 1796 5247 1800
rect 5233 1787 5247 1796
rect 5613 1807 5627 1813
rect 5727 1796 5763 1803
rect 4636 1776 4673 1783
rect 4747 1773 4752 1787
rect 4788 1773 4792 1787
rect 4828 1773 4833 1787
rect 4967 1776 5003 1783
rect 4913 1767 4927 1773
rect 4016 1756 4093 1763
rect 4107 1756 4233 1763
rect 4247 1756 4313 1763
rect 4367 1756 4413 1763
rect 4647 1756 4673 1763
rect 4996 1763 5003 1776
rect 5027 1776 5072 1783
rect 5100 1786 5113 1787
rect 5108 1773 5113 1786
rect 5207 1773 5212 1787
rect 5233 1780 5234 1787
rect 5307 1776 5333 1783
rect 5387 1776 5433 1783
rect 5507 1776 5533 1783
rect 5593 1767 5607 1773
rect 4996 1756 5073 1763
rect 5633 1767 5647 1773
rect 5673 1767 5687 1773
rect 3816 1736 3933 1743
rect 4527 1736 4623 1743
rect 387 1716 693 1723
rect 867 1716 923 1723
rect 427 1696 573 1703
rect 916 1703 923 1716
rect 1187 1716 1493 1723
rect 1507 1716 1533 1723
rect 1547 1716 1933 1723
rect 2067 1713 2073 1727
rect 3067 1716 3513 1723
rect 3567 1716 3933 1723
rect 4007 1716 4133 1723
rect 4547 1716 4593 1723
rect 4616 1723 4623 1736
rect 5067 1736 5132 1743
rect 5353 1747 5367 1753
rect 5168 1736 5273 1743
rect 5427 1736 5453 1743
rect 5547 1736 5693 1743
rect 4616 1716 4663 1723
rect 916 1696 1053 1703
rect 1207 1696 1233 1703
rect 1387 1696 1633 1703
rect 2447 1696 2913 1703
rect 3367 1696 3543 1703
rect 367 1676 553 1683
rect 987 1676 1353 1683
rect 1367 1676 1613 1683
rect 1627 1676 1893 1683
rect 2067 1676 2693 1683
rect 2767 1676 2913 1683
rect 2967 1676 3233 1683
rect 3536 1683 3543 1696
rect 3787 1696 4033 1703
rect 4387 1696 4613 1703
rect 4656 1703 4663 1716
rect 4727 1716 4773 1723
rect 5160 1726 5173 1727
rect 4967 1716 5023 1723
rect 4656 1696 4713 1703
rect 4727 1696 4993 1703
rect 5016 1703 5023 1716
rect 5167 1713 5173 1726
rect 5227 1716 5272 1723
rect 5308 1713 5313 1727
rect 5547 1713 5553 1727
rect 5687 1726 5700 1727
rect 5687 1713 5693 1726
rect 5016 1696 5353 1703
rect 5367 1696 5412 1703
rect 5448 1696 5513 1703
rect 5527 1696 5633 1703
rect 3536 1676 3653 1683
rect 3807 1676 3953 1683
rect 4507 1676 4633 1683
rect 4807 1676 5033 1683
rect 5047 1680 5203 1683
rect 5047 1676 5207 1680
rect 5193 1667 5207 1676
rect 5287 1676 5433 1683
rect 5567 1676 5663 1683
rect 5656 1667 5663 1676
rect 5687 1676 5713 1683
rect 187 1653 193 1667
rect 547 1656 993 1663
rect 1287 1656 1313 1663
rect 1327 1656 1653 1663
rect 1667 1656 1913 1663
rect 2467 1656 2773 1663
rect 2787 1656 3133 1663
rect 3376 1656 3493 1663
rect 127 1636 503 1643
rect 327 1616 473 1623
rect 376 1607 383 1616
rect 496 1623 503 1636
rect 667 1636 833 1643
rect 1067 1636 1133 1643
rect 1567 1634 1573 1647
rect 1567 1633 1580 1634
rect 1707 1636 1753 1643
rect 2127 1636 2293 1643
rect 2307 1640 2623 1643
rect 2307 1636 2627 1640
rect 2613 1627 2627 1636
rect 3376 1643 3383 1656
rect 3507 1656 3893 1663
rect 4347 1656 4533 1663
rect 4547 1656 4632 1663
rect 4668 1656 4713 1663
rect 4867 1656 4953 1663
rect 5347 1656 5473 1663
rect 5607 1653 5613 1667
rect 5656 1656 5673 1667
rect 5660 1653 5673 1656
rect 2907 1636 3383 1643
rect 3407 1636 3433 1643
rect 4227 1634 4233 1647
rect 4220 1633 4233 1634
rect 4927 1636 5153 1643
rect 5176 1636 5293 1643
rect 496 1616 683 1623
rect 47 1596 93 1603
rect 147 1596 193 1603
rect 207 1596 232 1603
rect 268 1596 353 1603
rect 376 1596 393 1607
rect 380 1593 393 1596
rect 516 1600 573 1603
rect 473 1587 487 1593
rect 127 1573 133 1587
rect 287 1576 333 1583
rect 427 1573 433 1587
rect 513 1596 573 1600
rect 513 1587 527 1596
rect 676 1603 683 1616
rect 747 1620 903 1623
rect 747 1616 907 1620
rect 893 1607 907 1616
rect 676 1596 752 1603
rect 788 1596 812 1603
rect 833 1593 834 1600
rect 1147 1616 1273 1623
rect 1287 1616 1443 1623
rect 933 1607 947 1613
rect 1313 1607 1327 1616
rect 1436 1607 1443 1616
rect 1467 1616 1573 1623
rect 1887 1616 1933 1623
rect 2147 1616 2193 1623
rect 2627 1620 2823 1623
rect 2627 1616 2827 1620
rect 2813 1607 2827 1616
rect 2853 1607 2867 1613
rect 2907 1616 3033 1623
rect 3196 1620 3233 1623
rect 3193 1616 3233 1620
rect 3193 1607 3207 1616
rect 3247 1616 3263 1623
rect 3376 1620 3483 1623
rect 976 1596 1012 1603
rect 653 1587 667 1593
rect 833 1587 847 1593
rect 976 1587 983 1596
rect 1048 1593 1053 1607
rect 1127 1596 1153 1603
rect 1167 1596 1263 1603
rect 707 1576 793 1583
rect 967 1576 983 1587
rect 967 1573 980 1576
rect 1007 1576 1033 1583
rect 1147 1576 1173 1583
rect 1227 1573 1233 1587
rect 1256 1583 1263 1596
rect 1367 1596 1413 1603
rect 1436 1596 1452 1607
rect 1440 1593 1452 1596
rect 1488 1593 1493 1607
rect 1707 1596 1753 1603
rect 1873 1587 1887 1593
rect 1256 1576 1333 1583
rect 1467 1573 1473 1587
rect 1527 1576 1573 1583
rect 1587 1573 1592 1587
rect 1626 1573 1627 1580
rect 1648 1573 1653 1587
rect 1727 1573 1733 1587
rect 2027 1593 2033 1607
rect 2267 1596 2293 1603
rect 2367 1596 2423 1603
rect 1913 1587 1927 1593
rect 2416 1587 2423 1596
rect 2707 1593 2713 1607
rect 2767 1593 2773 1607
rect 2866 1600 2867 1607
rect 2888 1596 3033 1603
rect 2473 1587 2487 1593
rect 1987 1576 2013 1583
rect 2067 1576 2133 1583
rect 2147 1573 2153 1587
rect 2207 1573 2213 1587
rect 2307 1576 2333 1583
rect 2387 1573 2393 1587
rect 2416 1573 2433 1587
rect 2627 1576 2693 1583
rect 2776 1583 2783 1593
rect 3056 1600 3163 1603
rect 3053 1596 3163 1600
rect 3053 1587 3067 1596
rect 3113 1587 3127 1596
rect 2776 1576 2833 1583
rect 2947 1576 2973 1583
rect 3106 1573 3107 1580
rect 3126 1580 3127 1587
rect 3133 1573 3134 1580
rect 3156 1583 3163 1596
rect 3256 1603 3263 1616
rect 3373 1616 3487 1620
rect 3373 1607 3387 1616
rect 3256 1596 3333 1603
rect 3473 1607 3487 1616
rect 3767 1613 3773 1627
rect 3787 1613 3793 1627
rect 3887 1620 3923 1623
rect 3887 1616 3927 1620
rect 3513 1607 3527 1613
rect 3913 1607 3927 1616
rect 4147 1616 4173 1623
rect 4187 1616 4213 1623
rect 4033 1607 4047 1613
rect 4267 1616 4313 1623
rect 4407 1616 4453 1623
rect 4787 1620 4824 1623
rect 4787 1616 4827 1620
rect 4533 1607 4547 1613
rect 4813 1607 4827 1616
rect 4847 1623 4860 1627
rect 4847 1620 4863 1623
rect 4847 1613 4867 1620
rect 4966 1613 4967 1620
rect 4853 1607 4867 1613
rect 4953 1607 4967 1613
rect 5133 1607 5147 1613
rect 3587 1600 3763 1603
rect 3587 1596 3767 1600
rect 3753 1587 3767 1596
rect 3987 1593 3993 1607
rect 4207 1600 4523 1603
rect 4207 1596 4527 1600
rect 4513 1587 4527 1596
rect 4607 1596 4713 1603
rect 4767 1596 4792 1603
rect 4813 1593 4814 1607
rect 4966 1600 4967 1607
rect 4988 1593 4993 1607
rect 5047 1596 5093 1603
rect 4813 1587 4827 1593
rect 5176 1587 5183 1636
rect 5627 1636 5673 1643
rect 5347 1616 5393 1623
rect 5647 1616 5713 1623
rect 5207 1596 5253 1603
rect 5447 1596 5483 1603
rect 3156 1576 3233 1583
rect 3247 1576 3353 1583
rect 3407 1573 3413 1587
rect 3487 1573 3493 1587
rect 3547 1576 3633 1583
rect 3827 1573 3833 1587
rect 4147 1576 4192 1583
rect 4228 1576 4292 1583
rect 4313 1573 4314 1580
rect 4367 1576 4433 1583
rect 4447 1573 4453 1587
rect 4536 1576 4573 1583
rect 73 1567 87 1573
rect 233 1563 247 1573
rect 373 1567 387 1573
rect 127 1556 313 1563
rect 436 1563 443 1573
rect 436 1556 492 1563
rect 528 1553 533 1567
rect 687 1553 693 1567
rect 707 1556 773 1563
rect 793 1563 807 1573
rect 913 1567 927 1573
rect 1073 1567 1087 1573
rect 793 1560 892 1563
rect 796 1556 892 1560
rect 913 1560 914 1567
rect 1373 1563 1387 1573
rect 1613 1567 1627 1573
rect 1373 1560 1493 1563
rect 1376 1556 1493 1560
rect 1773 1567 1787 1573
rect 1967 1556 2033 1563
rect 2047 1556 2173 1563
rect 2416 1563 2423 1573
rect 2733 1567 2747 1573
rect 2247 1556 2423 1563
rect 2727 1560 2747 1567
rect 2873 1567 2887 1573
rect 3093 1567 3107 1573
rect 2727 1556 2743 1560
rect 2727 1553 2740 1556
rect 2966 1553 2967 1560
rect 2988 1553 2993 1567
rect 3133 1567 3147 1573
rect 4313 1567 4327 1573
rect 3387 1556 3553 1563
rect 3607 1556 3653 1563
rect 3667 1553 3673 1567
rect 4326 1560 4327 1567
rect 4348 1556 4413 1563
rect 4467 1553 4473 1567
rect 4536 1563 4543 1576
rect 4647 1576 4693 1583
rect 4747 1576 4773 1583
rect 4826 1580 4827 1587
rect 4833 1573 4834 1580
rect 4887 1576 4952 1583
rect 4973 1573 4974 1580
rect 5027 1576 5053 1583
rect 5167 1576 5183 1587
rect 5167 1573 5180 1576
rect 5207 1576 5233 1583
rect 5476 1583 5483 1596
rect 5507 1593 5513 1607
rect 5567 1596 5613 1603
rect 5520 1586 5532 1587
rect 5476 1576 5513 1583
rect 4487 1556 4543 1563
rect 4596 1556 4673 1563
rect 407 1536 573 1543
rect 1193 1543 1207 1553
rect 1893 1547 1907 1553
rect 1007 1540 1207 1543
rect 1007 1536 1203 1540
rect 1347 1536 1453 1543
rect 2453 1543 2467 1553
rect 2453 1540 2693 1543
rect 2456 1536 2693 1540
rect 2953 1543 2967 1553
rect 2867 1540 2967 1543
rect 2867 1536 2962 1540
rect 3307 1536 3493 1543
rect 4107 1536 4153 1543
rect 4273 1543 4287 1553
rect 4227 1536 4353 1543
rect 4596 1543 4603 1556
rect 4833 1563 4847 1573
rect 4973 1563 4987 1573
rect 4747 1560 4987 1563
rect 5113 1563 5127 1573
rect 5273 1567 5287 1573
rect 5113 1560 5173 1563
rect 4747 1556 4984 1560
rect 5116 1556 5173 1560
rect 4507 1536 4603 1543
rect 4827 1536 5053 1543
rect 5416 1543 5423 1573
rect 5453 1563 5467 1573
rect 5527 1573 5532 1586
rect 5568 1573 5573 1587
rect 5453 1560 5493 1563
rect 5456 1556 5493 1560
rect 5607 1556 5693 1563
rect 5127 1536 5403 1543
rect 5416 1536 5613 1543
rect 1087 1516 1213 1523
rect 1427 1516 1713 1523
rect 1847 1516 2753 1523
rect 2807 1516 3093 1523
rect 4667 1516 4772 1523
rect 4808 1516 5353 1523
rect 5396 1523 5403 1536
rect 5396 1516 5493 1523
rect 5548 1516 5653 1523
rect 87 1496 313 1503
rect 327 1496 593 1503
rect 1567 1493 1573 1507
rect 1867 1496 2053 1503
rect 2327 1496 2713 1503
rect 2727 1496 2873 1503
rect 3227 1496 3333 1503
rect 3447 1496 3533 1503
rect 4167 1496 4273 1503
rect 4447 1496 4673 1503
rect 5147 1496 5273 1503
rect 5333 1493 5334 1500
rect 5587 1496 5613 1503
rect 5333 1487 5347 1493
rect 1487 1476 1973 1483
rect 1987 1476 2213 1483
rect 2547 1476 2993 1483
rect 3147 1476 3503 1483
rect 1127 1456 1213 1463
rect 1227 1456 1793 1463
rect 2567 1456 3113 1463
rect 3167 1456 3393 1463
rect 3496 1463 3503 1476
rect 3807 1476 4133 1483
rect 4247 1476 4313 1483
rect 4407 1476 4713 1483
rect 4927 1473 4933 1487
rect 4947 1476 5053 1483
rect 5167 1476 5312 1483
rect 5333 1480 5334 1487
rect 5356 1476 5633 1483
rect 3496 1456 4353 1463
rect 4667 1456 4953 1463
rect 5356 1463 5363 1476
rect 5687 1473 5693 1487
rect 5247 1456 5363 1463
rect 5376 1456 5453 1463
rect 616 1436 853 1443
rect 616 1423 623 1436
rect 1207 1436 1413 1443
rect 1427 1436 2332 1443
rect 2368 1436 2793 1443
rect 3327 1436 3413 1443
rect 3467 1436 3993 1443
rect 4047 1436 4173 1443
rect 4287 1436 4333 1443
rect 4607 1436 4693 1443
rect 4927 1436 5113 1443
rect 5376 1443 5383 1456
rect 5327 1436 5383 1443
rect 5427 1436 5553 1443
rect 467 1416 623 1423
rect 707 1416 913 1423
rect 927 1416 1232 1423
rect 1268 1416 1533 1423
rect 2407 1416 2453 1423
rect 2467 1413 2473 1427
rect 2947 1416 3413 1423
rect 3427 1416 3633 1423
rect 4107 1416 4373 1423
rect 4607 1416 4852 1423
rect 4888 1416 4933 1423
rect 5027 1416 5273 1423
rect 5407 1416 5613 1423
rect 647 1396 933 1403
rect 1287 1396 1513 1403
rect 2347 1396 2433 1403
rect 4147 1396 4473 1403
rect 4567 1396 4833 1403
rect 4967 1396 5113 1403
rect 5407 1396 5433 1403
rect 5527 1396 5713 1403
rect 247 1376 343 1383
rect 336 1367 343 1376
rect 587 1376 1013 1383
rect 1747 1376 1833 1383
rect 2047 1376 2393 1383
rect 2627 1376 2953 1383
rect 3967 1376 4013 1383
rect 4647 1376 4793 1383
rect 4907 1376 4973 1383
rect 5107 1376 5173 1383
rect 5507 1376 5583 1383
rect 217 1360 312 1363
rect 213 1356 312 1360
rect 213 1347 227 1356
rect 348 1363 360 1367
rect 348 1356 513 1363
rect 348 1353 367 1356
rect 807 1360 923 1363
rect 807 1356 927 1360
rect 353 1347 367 1353
rect 913 1347 927 1356
rect 1173 1347 1187 1353
rect 76 1340 192 1343
rect 73 1336 192 1340
rect 73 1327 87 1336
rect 213 1340 214 1347
rect 206 1333 207 1340
rect 287 1333 293 1347
rect 427 1336 493 1343
rect 987 1333 993 1347
rect 1467 1356 2113 1363
rect 2127 1356 2213 1363
rect 2227 1356 2333 1363
rect 2467 1360 2543 1363
rect 2467 1356 2547 1360
rect 1213 1347 1227 1353
rect 1287 1336 1313 1343
rect 1367 1336 1393 1343
rect 1407 1333 1413 1347
rect 1547 1333 1553 1347
rect 1607 1336 1753 1343
rect 1995 1340 2073 1343
rect 1993 1336 2073 1340
rect 193 1327 207 1333
rect 633 1327 647 1333
rect 1993 1327 2007 1336
rect 2267 1333 2273 1347
rect 2533 1347 2547 1356
rect 3047 1356 3193 1363
rect 3207 1356 3273 1363
rect 3627 1356 3893 1363
rect 3987 1356 4273 1363
rect 4296 1360 4833 1363
rect 4293 1356 4833 1360
rect 4293 1347 4307 1356
rect 4847 1356 4873 1363
rect 4967 1353 4973 1367
rect 5087 1356 5253 1363
rect 5296 1360 5453 1363
rect 5293 1356 5453 1360
rect 5293 1347 5307 1356
rect 5540 1363 5553 1367
rect 5536 1360 5553 1363
rect 5533 1353 5553 1360
rect 5533 1347 5547 1353
rect 5576 1347 5583 1376
rect 2367 1336 2412 1343
rect 2448 1336 2493 1343
rect 2616 1340 2742 1343
rect 2777 1340 2893 1343
rect 2616 1336 2747 1340
rect 2616 1327 2623 1336
rect 2733 1327 2747 1336
rect 2773 1336 2893 1340
rect 2773 1327 2787 1336
rect 2920 1343 2933 1347
rect 2916 1340 2933 1343
rect 2913 1333 2933 1340
rect 4227 1333 4233 1347
rect 4367 1333 4373 1347
rect 4427 1336 4453 1343
rect 4540 1343 4553 1347
rect 4536 1333 4553 1343
rect 4987 1336 5013 1343
rect 5056 1340 5093 1343
rect 5053 1336 5093 1340
rect 2913 1327 2927 1333
rect 4133 1327 4147 1333
rect 247 1313 253 1327
rect 327 1313 332 1327
rect 368 1313 373 1327
rect 447 1316 512 1323
rect 548 1313 553 1327
rect 787 1313 792 1327
rect 828 1313 833 1327
rect 887 1313 893 1327
rect 1087 1316 1172 1323
rect 1208 1313 1212 1327
rect 1248 1316 1333 1323
rect 1447 1316 1513 1323
rect 1587 1316 1633 1323
rect 1727 1316 1793 1323
rect 1927 1320 1983 1323
rect 1927 1316 1987 1320
rect 113 1307 127 1313
rect 673 1307 687 1313
rect 106 1293 107 1300
rect 126 1300 127 1307
rect 148 1293 153 1307
rect 666 1293 667 1300
rect 686 1300 687 1307
rect 708 1296 753 1303
rect 847 1293 853 1307
rect 933 1303 947 1313
rect 1973 1307 1987 1316
rect 2006 1320 2007 1327
rect 2028 1313 2033 1327
rect 2167 1316 2213 1323
rect 2227 1316 2353 1323
rect 2407 1313 2413 1327
rect 2467 1313 2473 1327
rect 2513 1307 2527 1313
rect 933 1300 1033 1303
rect 936 1296 1033 1300
rect 1127 1293 1133 1307
rect 1680 1306 1700 1307
rect 93 1287 107 1293
rect 533 1283 547 1293
rect 533 1280 633 1283
rect 536 1276 633 1280
rect 653 1283 667 1293
rect 793 1283 807 1293
rect 1687 1293 1693 1306
rect 653 1280 783 1283
rect 793 1280 1073 1283
rect 656 1276 783 1280
rect 796 1276 1073 1280
rect 227 1256 553 1263
rect 776 1263 783 1276
rect 1746 1273 1747 1280
rect 1768 1276 1873 1283
rect 2013 1283 2027 1293
rect 2307 1293 2313 1307
rect 2613 1307 2627 1313
rect 2746 1320 2747 1327
rect 2773 1320 2774 1327
rect 2766 1313 2767 1320
rect 2936 1316 3013 1323
rect 2653 1307 2667 1313
rect 2753 1307 2767 1313
rect 2667 1296 2713 1303
rect 2766 1300 2767 1307
rect 2936 1303 2943 1316
rect 3166 1313 3167 1320
rect 3188 1313 3193 1327
rect 3216 1316 3253 1323
rect 2907 1296 2943 1303
rect 2967 1293 2973 1307
rect 3027 1296 3053 1303
rect 3107 1293 3113 1307
rect 2233 1287 2247 1293
rect 2793 1287 2807 1293
rect 2013 1280 2073 1283
rect 2016 1276 2073 1280
rect 2167 1273 2173 1287
rect 2647 1276 2743 1283
rect 776 1256 1033 1263
rect 1247 1253 1253 1267
rect 1733 1263 1747 1273
rect 1687 1260 1747 1263
rect 1687 1256 1742 1260
rect 1947 1256 2233 1263
rect 2247 1256 2493 1263
rect 2736 1263 2743 1276
rect 3135 1283 3142 1313
rect 3153 1307 3167 1313
rect 3216 1307 3223 1316
rect 3647 1316 3733 1323
rect 3787 1313 3792 1327
rect 3828 1316 3853 1323
rect 3907 1313 3913 1327
rect 4227 1316 4273 1323
rect 4356 1323 4363 1333
rect 4327 1316 4363 1323
rect 4407 1316 4473 1323
rect 4536 1307 4543 1333
rect 4633 1327 4647 1333
rect 4687 1316 4713 1323
rect 4787 1314 4792 1327
rect 5053 1327 5067 1336
rect 5175 1336 5243 1343
rect 4787 1313 4800 1314
rect 4828 1313 4833 1327
rect 4947 1313 4953 1327
rect 4967 1316 5013 1323
rect 3166 1300 3167 1307
rect 3207 1296 3223 1307
rect 3207 1293 3220 1296
rect 3427 1293 3432 1307
rect 3453 1293 3454 1300
rect 3707 1293 3713 1307
rect 3867 1293 3873 1307
rect 3987 1293 3993 1307
rect 4047 1296 4133 1303
rect 4187 1296 4273 1303
rect 4427 1296 4493 1303
rect 4607 1293 4612 1307
rect 4648 1293 4653 1307
rect 4716 1303 4723 1313
rect 5175 1307 5182 1336
rect 5236 1323 5243 1336
rect 5347 1336 5413 1343
rect 5236 1316 5313 1323
rect 5356 1316 5432 1323
rect 4716 1296 4753 1303
rect 4807 1293 4813 1307
rect 4947 1296 4993 1303
rect 5087 1296 5152 1303
rect 5208 1293 5213 1307
rect 5356 1303 5363 1316
rect 5468 1313 5473 1327
rect 5487 1316 5553 1323
rect 5596 1316 5653 1323
rect 5327 1296 5363 1303
rect 5387 1293 5392 1307
rect 5428 1296 5453 1303
rect 5596 1303 5603 1316
rect 5467 1296 5603 1303
rect 3135 1276 3233 1283
rect 3307 1273 3313 1287
rect 3333 1283 3347 1293
rect 3327 1280 3347 1283
rect 3327 1276 3343 1280
rect 3453 1283 3467 1293
rect 3407 1280 3467 1283
rect 3753 1287 3767 1293
rect 3407 1276 3464 1280
rect 3767 1276 3813 1283
rect 3913 1283 3927 1293
rect 4893 1287 4907 1293
rect 3913 1280 4013 1283
rect 3916 1276 4013 1280
rect 4327 1276 4373 1283
rect 4527 1273 4532 1287
rect 4568 1276 4613 1283
rect 4667 1276 4833 1283
rect 5033 1283 5047 1293
rect 5033 1280 5133 1283
rect 5036 1276 5133 1280
rect 5207 1276 5443 1283
rect 2736 1256 2853 1263
rect 2993 1263 3007 1273
rect 2993 1260 3053 1263
rect 2996 1256 3053 1260
rect 3647 1256 3693 1263
rect 3707 1256 4033 1263
rect 4587 1256 4913 1263
rect 5027 1256 5093 1263
rect 5107 1256 5193 1263
rect 5207 1256 5293 1263
rect 5436 1263 5443 1276
rect 5667 1276 5693 1283
rect 5436 1256 5473 1263
rect 47 1236 353 1243
rect 556 1243 563 1253
rect 556 1236 893 1243
rect 1087 1236 1733 1243
rect 1747 1236 1792 1243
rect 1828 1236 2253 1243
rect 2307 1236 2372 1243
rect 2408 1236 2653 1243
rect 2767 1236 2953 1243
rect 3927 1236 4073 1243
rect 4087 1236 4573 1243
rect 4767 1236 4893 1243
rect 4967 1236 5013 1243
rect 5647 1236 5673 1243
rect 687 1216 832 1223
rect 868 1216 1213 1223
rect 1307 1216 1973 1223
rect 2367 1216 2553 1223
rect 2727 1216 2903 1223
rect 107 1196 553 1203
rect 1267 1196 1573 1203
rect 2896 1207 2903 1216
rect 3387 1216 3453 1223
rect 3467 1216 3703 1223
rect 2347 1196 2753 1203
rect 2907 1196 3113 1203
rect 3327 1196 3443 1203
rect 127 1176 173 1183
rect 447 1176 753 1183
rect 1147 1176 1373 1183
rect 1587 1176 1853 1183
rect 2307 1176 2353 1183
rect 3227 1176 3333 1183
rect 3436 1183 3443 1196
rect 3467 1196 3513 1203
rect 3696 1203 3703 1216
rect 3727 1216 4213 1223
rect 4627 1216 4933 1223
rect 5007 1216 5233 1223
rect 5347 1216 5513 1223
rect 3696 1196 3753 1203
rect 4967 1196 5313 1203
rect 5607 1196 5693 1203
rect 3436 1176 3473 1183
rect 4687 1176 4853 1183
rect 5147 1176 5233 1183
rect 5507 1176 5573 1183
rect 5653 1167 5667 1173
rect 107 1156 173 1163
rect 187 1156 293 1163
rect 587 1156 673 1163
rect 687 1156 713 1163
rect 807 1156 933 1163
rect 1007 1156 1193 1163
rect 1207 1156 1353 1163
rect 1447 1156 1673 1163
rect 1687 1153 1693 1167
rect 1827 1153 1833 1167
rect 2527 1156 2793 1163
rect 2807 1160 2923 1163
rect 2807 1156 2927 1160
rect 2913 1147 2927 1156
rect 3047 1156 3273 1163
rect 3287 1156 3513 1163
rect 3587 1156 3613 1163
rect 4167 1156 4293 1163
rect 4547 1156 4993 1163
rect 5167 1156 5253 1163
rect 5276 1156 5373 1163
rect 5093 1147 5107 1153
rect 93 1127 107 1133
rect 133 1127 147 1133
rect 507 1136 613 1143
rect 916 1136 1013 1143
rect 493 1127 507 1133
rect 160 1123 173 1127
rect 156 1113 173 1123
rect 287 1116 353 1123
rect 427 1113 433 1127
rect 536 1116 683 1123
rect 47 1096 73 1103
rect 156 1103 163 1113
rect 273 1107 287 1113
rect 536 1107 543 1116
rect 676 1107 683 1116
rect 747 1113 753 1127
rect 916 1123 923 1136
rect 1367 1136 1453 1143
rect 1707 1136 1793 1143
rect 1807 1136 1853 1143
rect 1867 1133 1873 1147
rect 2307 1136 2413 1143
rect 2827 1133 2833 1147
rect 2927 1136 3013 1143
rect 3056 1140 3093 1143
rect 3053 1136 3093 1140
rect 1353 1127 1367 1133
rect 3053 1127 3067 1136
rect 3107 1140 3183 1143
rect 3107 1136 3187 1140
rect 3173 1127 3187 1136
rect 3267 1136 3312 1143
rect 3333 1133 3334 1140
rect 3427 1136 3483 1143
rect 3333 1127 3347 1133
rect 3476 1127 3483 1136
rect 3647 1143 3660 1147
rect 3647 1133 3663 1143
rect 3987 1133 3993 1147
rect 4047 1133 4053 1147
rect 4367 1136 4453 1143
rect 4667 1136 4733 1143
rect 4807 1136 4873 1143
rect 5027 1133 5033 1147
rect 3656 1127 3663 1133
rect 4593 1127 4607 1133
rect 5173 1127 5187 1133
rect 5276 1127 5283 1156
rect 5387 1156 5553 1163
rect 5427 1133 5433 1147
rect 5313 1127 5327 1133
rect 5516 1127 5523 1156
rect 5547 1136 5573 1143
rect 807 1116 923 1123
rect 1047 1113 1052 1127
rect 1088 1113 1092 1127
rect 1128 1113 1133 1127
rect 1556 1120 1643 1123
rect 1556 1116 1647 1120
rect 933 1107 947 1113
rect 127 1096 163 1103
rect 187 1096 233 1103
rect 286 1100 287 1107
rect 308 1096 333 1103
rect 227 1073 232 1087
rect 268 1076 313 1083
rect 373 1083 387 1093
rect 327 1080 387 1083
rect 527 1096 543 1107
rect 527 1093 540 1096
rect 607 1093 613 1107
rect 667 1093 673 1107
rect 727 1096 773 1103
rect 827 1096 853 1103
rect 867 1096 893 1103
rect 473 1083 487 1093
rect 473 1080 553 1083
rect 327 1076 383 1080
rect 476 1076 553 1080
rect 567 1076 633 1083
rect 707 1076 793 1083
rect 907 1073 913 1087
rect 1073 1083 1087 1093
rect 987 1080 1087 1083
rect 1187 1093 1192 1107
rect 1228 1093 1233 1107
rect 1327 1093 1333 1107
rect 1556 1103 1563 1116
rect 1633 1107 1647 1116
rect 1727 1113 1733 1127
rect 1787 1116 1933 1123
rect 1987 1116 2133 1123
rect 2207 1123 2220 1127
rect 2207 1113 2223 1123
rect 2247 1113 2253 1127
rect 2307 1116 2333 1123
rect 2380 1123 2393 1127
rect 2376 1113 2393 1123
rect 2447 1116 2473 1123
rect 2727 1116 2793 1123
rect 2847 1113 2853 1127
rect 3107 1113 3113 1127
rect 3247 1116 3292 1123
rect 3333 1120 3334 1127
rect 3326 1113 3327 1120
rect 3407 1116 3453 1123
rect 3476 1116 3493 1127
rect 3480 1113 3493 1116
rect 3547 1123 3560 1127
rect 3547 1113 3563 1123
rect 3656 1123 3673 1127
rect 3627 1116 3673 1123
rect 3660 1113 3673 1116
rect 3747 1113 3753 1127
rect 3867 1116 3952 1123
rect 3988 1113 3993 1127
rect 4087 1113 4093 1127
rect 4540 1123 4553 1127
rect 4536 1113 4553 1123
rect 4615 1120 4913 1123
rect 4613 1116 4913 1120
rect 1973 1107 1987 1113
rect 1507 1096 1563 1103
rect 1113 1083 1127 1093
rect 1373 1087 1387 1093
rect 1593 1087 1607 1093
rect 1113 1080 1153 1083
rect 987 1076 1083 1080
rect 1116 1076 1153 1080
rect 1287 1073 1293 1087
rect 1467 1073 1473 1087
rect 1606 1080 1607 1087
rect 1613 1073 1614 1080
rect 1753 1083 1767 1093
rect 1707 1080 1767 1083
rect 1927 1096 1963 1103
rect 1793 1087 1807 1093
rect 1707 1076 1763 1080
rect 1956 1083 1963 1096
rect 2027 1093 2033 1107
rect 2047 1096 2113 1103
rect 2216 1103 2223 1113
rect 2216 1096 2273 1103
rect 2287 1093 2292 1107
rect 2313 1093 2314 1100
rect 2376 1103 2383 1113
rect 3313 1107 3327 1113
rect 2328 1096 2383 1103
rect 2407 1093 2413 1107
rect 2507 1096 2532 1103
rect 2568 1093 2573 1107
rect 2627 1096 2693 1103
rect 2716 1100 2753 1103
rect 2713 1096 2753 1100
rect 1956 1076 1993 1083
rect 2153 1083 2167 1093
rect 2007 1080 2167 1083
rect 2007 1076 2163 1080
rect 2187 1076 2233 1083
rect 2313 1083 2327 1093
rect 2247 1080 2327 1083
rect 2453 1083 2467 1093
rect 2713 1087 2727 1096
rect 2887 1096 2913 1103
rect 3027 1093 3033 1107
rect 2453 1080 2553 1083
rect 2247 1076 2324 1080
rect 2456 1076 2553 1080
rect 2627 1076 2673 1083
rect 3073 1087 3087 1093
rect 3153 1087 3167 1093
rect 3447 1096 3472 1103
rect 3508 1093 3513 1107
rect 3556 1103 3563 1113
rect 3556 1096 3593 1103
rect 3193 1087 3207 1093
rect 3353 1083 3367 1093
rect 3793 1103 3807 1113
rect 3767 1100 3807 1103
rect 3767 1096 3803 1100
rect 4127 1093 4133 1107
rect 4227 1093 4233 1107
rect 4347 1093 4353 1107
rect 4536 1103 4543 1113
rect 4613 1107 4627 1116
rect 4856 1107 4863 1116
rect 4967 1113 4973 1127
rect 5127 1113 5133 1127
rect 5387 1116 5413 1123
rect 5467 1113 5473 1127
rect 5516 1116 5533 1127
rect 5520 1113 5533 1116
rect 5587 1116 5613 1123
rect 5627 1113 5633 1127
rect 4507 1096 4543 1103
rect 4567 1093 4573 1107
rect 4626 1100 4627 1107
rect 4648 1096 4693 1103
rect 4847 1096 4863 1107
rect 4847 1093 4860 1096
rect 4887 1093 4893 1107
rect 4947 1096 5033 1103
rect 5147 1093 5153 1107
rect 5207 1093 5213 1107
rect 5267 1096 5293 1103
rect 5527 1096 5553 1103
rect 4273 1087 4287 1093
rect 3307 1076 3653 1083
rect 3987 1076 4073 1083
rect 4187 1073 4193 1087
rect 4247 1073 4252 1087
rect 4273 1080 4274 1087
rect 4327 1073 4333 1087
rect 4387 1076 4593 1083
rect 4707 1076 4833 1083
rect 5127 1076 5273 1083
rect 5333 1083 5347 1093
rect 5287 1080 5347 1083
rect 5593 1087 5607 1093
rect 5287 1076 5343 1080
rect 687 1056 973 1063
rect 1213 1063 1227 1073
rect 1027 1056 1313 1063
rect 1513 1063 1527 1073
rect 1327 1060 1527 1063
rect 1327 1056 1523 1060
rect 1613 1063 1627 1073
rect 1567 1060 1627 1063
rect 1653 1063 1667 1073
rect 1653 1060 2033 1063
rect 1567 1056 1624 1060
rect 1656 1056 2033 1060
rect 2553 1063 2567 1073
rect 2087 1060 2567 1063
rect 2087 1056 2563 1060
rect 3067 1056 3193 1063
rect 3407 1056 3573 1063
rect 4287 1056 4373 1063
rect 4727 1056 5093 1063
rect 5207 1056 5313 1063
rect 5447 1056 5633 1063
rect 1127 1036 1593 1043
rect 2707 1036 2733 1043
rect 2867 1036 3073 1043
rect 4167 1033 4173 1047
rect 4247 1036 4313 1043
rect 4487 1036 4873 1043
rect 5007 1036 5033 1043
rect 5467 1036 5493 1043
rect 287 1016 1213 1023
rect 1227 1016 1373 1023
rect 2227 1016 3333 1023
rect 5027 1016 5073 1023
rect 5387 1016 5553 1023
rect 1833 1007 1847 1013
rect 2447 996 2593 1003
rect 2747 996 3253 1003
rect 3427 996 3603 1003
rect 3596 983 3603 996
rect 3627 996 3652 1003
rect 3688 996 4033 1003
rect 4507 996 5113 1003
rect 5247 996 5593 1003
rect 3596 976 3753 983
rect 4087 976 4153 983
rect 4327 976 4373 983
rect 5007 976 5093 983
rect 5507 976 5533 983
rect 5653 983 5667 993
rect 5607 980 5667 983
rect 5607 976 5663 980
rect 2667 956 3173 963
rect 3807 956 4033 963
rect 4047 956 4333 963
rect 4427 956 4793 963
rect 4847 956 5133 963
rect 267 936 373 943
rect 707 936 973 943
rect 1027 936 1153 943
rect 1167 936 1553 943
rect 3047 936 3233 943
rect 3567 936 3833 943
rect 4127 936 4373 943
rect 4687 936 5053 943
rect 5307 936 5393 943
rect 5467 933 5473 947
rect 5567 936 5633 943
rect 347 916 593 923
rect 607 916 693 923
rect 1327 916 1833 923
rect 2007 916 2313 923
rect 2647 916 3273 923
rect 3547 916 3733 923
rect 4107 916 4173 923
rect 4527 916 4813 923
rect 4867 916 4973 923
rect 5067 916 5173 923
rect 5247 916 5693 923
rect 107 896 253 903
rect 267 896 713 903
rect 727 896 813 903
rect 1827 896 2053 903
rect 2867 896 3113 903
rect 3127 896 3153 903
rect 3927 896 4243 903
rect 167 876 233 883
rect 616 876 693 883
rect 327 853 333 867
rect 387 853 393 867
rect 616 863 623 876
rect 707 876 724 883
rect 527 856 623 863
rect 193 847 207 853
rect 453 847 467 853
rect 107 836 153 843
rect 247 836 293 843
rect 427 833 432 847
rect 453 840 454 847
rect 473 833 474 840
rect 607 834 612 847
rect 717 847 724 876
rect 1207 876 1573 883
rect 1587 876 1693 883
rect 1887 876 2013 883
rect 2027 876 2273 883
rect 2296 876 2413 883
rect 747 853 753 867
rect 807 856 853 863
rect 896 860 1233 863
rect 893 856 1233 860
rect 893 847 907 856
rect 1327 856 1353 863
rect 1647 856 1773 863
rect 1787 856 1913 863
rect 1927 856 1993 863
rect 2096 860 2173 863
rect 2093 856 2173 860
rect 1313 847 1327 853
rect 2093 847 2107 856
rect 2296 863 2303 876
rect 4236 887 4243 896
rect 4327 896 4433 903
rect 4727 893 4733 907
rect 4807 896 4852 903
rect 4888 896 5033 903
rect 5207 896 5273 903
rect 5327 893 5333 907
rect 5407 896 5433 903
rect 2927 876 2973 883
rect 3106 873 3107 880
rect 2873 867 2887 873
rect 3093 867 3107 873
rect 3993 867 4007 873
rect 2187 856 2303 863
rect 2487 856 2573 863
rect 2595 860 2633 863
rect 2593 856 2633 860
rect 607 833 620 834
rect 648 836 692 843
rect 827 836 853 843
rect 876 836 893 843
rect 333 823 347 833
rect 473 823 487 833
rect 333 820 573 823
rect 336 816 573 820
rect 627 813 632 827
rect 653 813 654 820
rect 753 823 767 833
rect 876 823 883 836
rect 947 836 1013 843
rect 1157 840 1252 843
rect 1053 827 1067 833
rect 1153 836 1252 840
rect 1153 827 1167 836
rect 1273 833 1274 840
rect 1447 833 1452 847
rect 1488 833 1493 847
rect 1947 833 1953 847
rect 2047 833 2053 847
rect 2207 833 2213 847
rect 2327 833 2333 847
rect 2593 847 2607 856
rect 2827 853 2833 867
rect 2927 856 2973 863
rect 3106 860 3107 867
rect 3113 853 3114 860
rect 3280 863 3292 867
rect 3277 860 3292 863
rect 3273 853 3292 860
rect 3328 856 3373 863
rect 3427 860 3524 863
rect 3427 856 3527 860
rect 3113 847 3127 853
rect 3273 847 3287 853
rect 2547 834 2553 847
rect 2540 833 2553 834
rect 2606 840 2607 847
rect 2628 836 2693 843
rect 2747 836 2773 843
rect 2867 833 2873 847
rect 2987 836 3013 843
rect 3067 833 3073 847
rect 3187 836 3233 843
rect 3247 833 3252 847
rect 3273 840 3274 847
rect 3387 836 3453 843
rect 3467 836 3492 843
rect 3513 847 3527 856
rect 3587 853 3593 867
rect 3707 853 3713 867
rect 3767 856 3873 863
rect 4033 867 4047 873
rect 4247 876 4953 883
rect 4976 876 5173 883
rect 4113 867 4127 873
rect 4167 853 4173 867
rect 4636 860 4733 863
rect 4633 856 4733 860
rect 4633 847 4647 856
rect 4787 853 4793 867
rect 4976 863 4983 876
rect 5367 876 5473 883
rect 5547 876 5673 883
rect 5233 867 5247 873
rect 4927 856 4983 863
rect 5136 860 5193 863
rect 5133 856 5193 860
rect 5133 847 5147 856
rect 5287 853 5293 867
rect 5396 860 5433 863
rect 5353 847 5367 853
rect 3513 840 3514 847
rect 3567 836 3592 843
rect 3613 833 3614 840
rect 3747 836 3853 843
rect 3907 833 3913 847
rect 4027 836 4053 843
rect 4207 833 4212 847
rect 4246 833 4247 840
rect 4268 836 4353 843
rect 4407 833 4413 847
rect 4467 833 4472 847
rect 4508 833 4513 847
rect 4787 846 4800 847
rect 4787 833 4792 846
rect 1273 827 1287 833
rect 753 820 883 823
rect 756 816 883 820
rect 987 816 1032 823
rect 1066 820 1067 827
rect 1088 816 1132 823
rect 1153 820 1154 827
rect 1207 813 1213 827
rect 1286 820 1287 827
rect 1293 813 1294 820
rect 1567 813 1573 827
rect 1687 813 1693 827
rect 1767 813 1773 827
rect 1847 816 1872 823
rect 1886 813 1887 820
rect 1908 813 1913 827
rect 2087 813 2093 827
rect 2153 823 2167 833
rect 2107 820 2167 823
rect 2107 816 2163 820
rect 2287 813 2293 827
rect 2367 816 2413 823
rect 2527 813 2533 827
rect 2667 813 2673 827
rect 2933 823 2947 833
rect 2727 820 2947 823
rect 2727 816 2943 820
rect 2967 816 2993 823
rect 3333 823 3347 833
rect 3167 820 3347 823
rect 3167 816 3343 820
rect 3427 813 3433 827
rect 3507 813 3512 827
rect 3613 823 3627 833
rect 3548 820 3627 823
rect 3548 816 3623 820
rect 3807 816 3833 823
rect 3887 816 3953 823
rect 173 807 187 813
rect 107 793 113 807
rect 247 796 433 803
rect 653 803 667 813
rect 653 800 813 803
rect 657 796 813 800
rect 887 796 973 803
rect 996 796 1173 803
rect 227 776 693 783
rect 996 783 1003 796
rect 1293 803 1307 813
rect 1333 807 1347 813
rect 1247 800 1307 803
rect 1247 796 1303 800
rect 1327 803 1347 807
rect 1327 796 1433 803
rect 1327 793 1340 796
rect 1447 796 1513 803
rect 1633 803 1647 813
rect 1873 807 1887 813
rect 1607 800 1647 803
rect 1607 796 1643 800
rect 1807 793 1813 807
rect 2033 803 2047 813
rect 2573 807 2587 813
rect 3353 807 3367 813
rect 2033 800 2133 803
rect 2036 796 2133 800
rect 2827 796 2953 803
rect 3366 800 3367 807
rect 3388 796 3453 803
rect 3687 796 4033 803
rect 4136 803 4143 833
rect 4233 827 4247 833
rect 4828 833 4833 847
rect 4847 836 4992 843
rect 5028 836 5093 843
rect 5187 836 5253 843
rect 5393 856 5433 860
rect 5393 847 5407 856
rect 5536 860 5593 863
rect 5533 856 5593 860
rect 5533 847 5547 856
rect 5607 856 5643 863
rect 5636 847 5643 856
rect 5487 833 5493 847
rect 5647 836 5673 843
rect 4287 813 4293 827
rect 4456 816 4493 823
rect 4456 807 4463 816
rect 4687 813 4693 827
rect 5067 816 5113 823
rect 5167 816 5372 823
rect 5408 813 5412 827
rect 5448 816 5512 823
rect 5548 813 5553 827
rect 5627 813 5632 827
rect 5653 813 5654 820
rect 4047 796 4143 803
rect 4167 796 4313 803
rect 4367 796 4393 803
rect 4407 793 4412 807
rect 4448 796 4463 807
rect 4533 803 4547 813
rect 4533 800 4633 803
rect 4536 796 4633 800
rect 4448 793 4460 796
rect 5007 793 5013 807
rect 5207 796 5353 803
rect 5653 803 5667 813
rect 5507 800 5667 803
rect 5507 796 5663 800
rect 707 776 1003 783
rect 1287 776 1503 783
rect 1496 767 1503 776
rect 1653 783 1667 793
rect 1607 776 1793 783
rect 1967 776 2213 783
rect 2267 776 2433 783
rect 2487 776 2673 783
rect 2747 776 2833 783
rect 3007 776 3553 783
rect 4467 776 4593 783
rect 4913 783 4927 793
rect 4913 780 5153 783
rect 4916 776 5153 780
rect 187 756 453 763
rect 627 756 733 763
rect 747 756 813 763
rect 867 756 932 763
rect 968 756 1053 763
rect 1067 756 1153 763
rect 1507 756 1973 763
rect 2047 756 2533 763
rect 2807 756 2913 763
rect 3187 756 3213 763
rect 3467 753 3473 767
rect 3527 756 3593 763
rect 3887 756 4573 763
rect 4727 756 4893 763
rect 5007 756 5313 763
rect 5467 756 5613 763
rect 367 736 493 743
rect 507 736 1553 743
rect 1576 736 1933 743
rect 927 716 1013 723
rect 1576 723 1583 736
rect 2067 736 2403 743
rect 1327 716 1583 723
rect 2396 723 2403 736
rect 2587 736 3153 743
rect 3247 736 3313 743
rect 3367 736 3493 743
rect 3967 736 4433 743
rect 4487 736 4533 743
rect 4947 736 5413 743
rect 2396 716 2733 723
rect 2787 716 3413 723
rect 3947 716 3993 723
rect 4387 716 4753 723
rect 4887 716 5273 723
rect 5347 716 5653 723
rect 107 696 333 703
rect 767 696 993 703
rect 1007 696 1233 703
rect 1467 696 1633 703
rect 1767 696 2153 703
rect 2227 696 2613 703
rect 2667 696 2693 703
rect 2856 696 3013 703
rect 2856 687 2863 696
rect 3347 696 3393 703
rect 3847 696 4173 703
rect 4287 696 4513 703
rect 4527 696 4673 703
rect 4807 696 4853 703
rect 5047 696 5113 703
rect 5327 696 5393 703
rect 327 676 553 683
rect 607 676 1073 683
rect 1147 676 1213 683
rect 1407 676 1593 683
rect 2447 676 2853 683
rect 2987 676 3113 683
rect 3287 676 3353 683
rect 3367 676 3593 683
rect 3607 676 3733 683
rect 3987 676 4083 683
rect 93 667 107 673
rect 1833 667 1847 673
rect 240 663 253 667
rect 236 660 253 663
rect 193 647 207 653
rect 233 653 253 660
rect 636 660 753 663
rect 633 656 753 660
rect 233 647 247 653
rect 633 647 647 656
rect 1176 660 1233 663
rect 1073 647 1087 653
rect 1173 656 1233 660
rect 1173 647 1187 656
rect 1547 656 1673 663
rect 1353 647 1367 653
rect 1613 647 1627 656
rect 2167 660 2243 663
rect 2167 656 2247 660
rect 2233 647 2247 656
rect 2387 656 2453 663
rect 2467 653 2473 667
rect 2776 660 2913 663
rect 387 636 453 643
rect 527 636 593 643
rect 607 640 622 643
rect 607 636 627 640
rect 107 616 173 623
rect 227 613 233 627
rect 347 614 352 627
rect 373 627 387 633
rect 613 627 627 636
rect 687 636 1033 643
rect 1087 636 1133 643
rect 1267 636 1313 643
rect 1456 640 1493 643
rect 1453 636 1493 640
rect 1453 627 1467 636
rect 1547 633 1553 647
rect 1613 640 1614 647
rect 1606 633 1607 640
rect 1747 633 1752 647
rect 1788 636 1833 643
rect 1593 627 1607 633
rect 1933 627 1947 633
rect 373 620 374 627
rect 347 613 360 614
rect 487 613 493 627
rect 626 620 627 627
rect 648 613 653 627
rect 747 613 753 627
rect 807 616 853 623
rect 947 616 972 623
rect 1008 613 1013 627
rect 1167 613 1172 627
rect 1208 613 1213 627
rect 1347 616 1393 623
rect 1507 616 1533 623
rect 1647 613 1653 627
rect 1667 616 1713 623
rect 1767 616 1793 623
rect 1887 616 1923 623
rect 327 603 340 607
rect 327 593 343 603
rect 367 593 373 607
rect 433 603 447 613
rect 387 600 447 603
rect 387 596 443 600
rect 707 593 713 607
rect 893 603 907 613
rect 207 576 313 583
rect 336 583 343 593
rect 336 576 633 583
rect 773 583 787 593
rect 836 600 907 603
rect 836 596 903 600
rect 836 583 843 596
rect 1053 603 1067 613
rect 1156 603 1163 613
rect 1053 600 1163 603
rect 1056 596 1163 600
rect 1293 607 1307 613
rect 1487 593 1493 607
rect 1916 603 1923 616
rect 1973 627 1987 633
rect 2136 640 2223 643
rect 2136 636 2227 640
rect 2056 616 2113 623
rect 1687 596 1953 603
rect 2056 603 2063 616
rect 2136 623 2143 636
rect 2213 627 2227 636
rect 2287 633 2293 647
rect 2406 633 2407 640
rect 2447 636 2473 643
rect 2673 647 2687 653
rect 2773 656 2913 660
rect 2587 636 2633 643
rect 2773 647 2787 656
rect 2927 656 2983 663
rect 2727 634 2733 647
rect 2720 633 2733 634
rect 2976 643 2983 656
rect 3227 656 3273 663
rect 3347 656 3473 663
rect 3553 647 3567 653
rect 3747 660 3923 663
rect 3747 656 3927 660
rect 3673 647 3687 653
rect 2976 636 3032 643
rect 3068 633 3073 647
rect 3487 633 3493 647
rect 3607 636 3633 643
rect 3913 647 3927 656
rect 3967 656 4053 663
rect 4076 663 4083 676
rect 4327 676 4473 683
rect 4607 676 4953 683
rect 5147 676 5553 683
rect 4076 656 4193 663
rect 4286 653 4287 660
rect 4308 666 4320 667
rect 4308 653 4313 666
rect 4273 647 4287 653
rect 4336 656 4412 663
rect 4336 647 4343 656
rect 4433 653 4434 660
rect 4448 656 4513 663
rect 4433 647 4447 653
rect 3696 640 3823 643
rect 3693 636 3827 640
rect 2353 627 2367 633
rect 2393 627 2407 633
rect 2953 627 2967 633
rect 3693 627 3707 636
rect 2127 616 2143 623
rect 2167 613 2173 627
rect 2353 620 2372 627
rect 2356 616 2372 620
rect 2360 613 2372 616
rect 2406 620 2407 627
rect 2480 626 2493 627
rect 2428 616 2473 623
rect 2027 596 2063 603
rect 2127 593 2133 607
rect 2253 603 2267 613
rect 2487 613 2493 626
rect 2607 613 2613 627
rect 2653 607 2667 613
rect 2727 616 2753 623
rect 2867 616 2913 623
rect 3007 613 3013 627
rect 3147 616 3192 623
rect 3213 613 3214 620
rect 3427 613 3432 627
rect 3468 616 3533 623
rect 3647 613 3653 627
rect 3813 627 3827 636
rect 3987 633 3993 647
rect 4087 636 4113 643
rect 4167 633 4173 647
rect 4327 636 4343 647
rect 4327 633 4340 636
rect 4407 633 4412 647
rect 4433 640 4434 647
rect 4496 636 4533 643
rect 4033 627 4047 633
rect 4213 627 4227 633
rect 3947 613 3953 627
rect 4033 620 4053 627
rect 4036 616 4053 620
rect 4040 613 4053 616
rect 4396 623 4403 633
rect 4496 623 4503 636
rect 4647 633 4653 647
rect 4707 633 4713 647
rect 4953 643 4967 653
rect 5076 656 5193 663
rect 5076 647 5083 656
rect 5407 656 5433 663
rect 5447 653 5452 667
rect 5488 656 5693 663
rect 4953 640 5013 643
rect 4956 636 5013 640
rect 5027 633 5032 647
rect 5068 633 5073 647
rect 5096 636 5273 643
rect 4396 616 4503 623
rect 4636 623 4643 633
rect 5096 627 5103 636
rect 5287 636 5313 643
rect 5367 633 5373 647
rect 5416 640 5563 643
rect 5416 636 5567 640
rect 4567 616 4643 623
rect 4667 613 4673 627
rect 4767 616 4812 623
rect 4848 616 4913 623
rect 4967 616 4993 623
rect 5087 616 5103 627
rect 5087 613 5100 616
rect 5127 613 5133 627
rect 5187 613 5193 627
rect 5280 626 5293 627
rect 2147 600 2267 603
rect 2147 596 2263 600
rect 2427 596 2652 603
rect 2666 600 2667 607
rect 2793 603 2807 613
rect 2688 600 2807 603
rect 2688 596 2803 600
rect 2927 593 2932 607
rect 3053 603 3067 613
rect 3213 607 3227 613
rect 3573 607 3587 613
rect 4513 607 4527 613
rect 2968 600 3067 603
rect 2968 596 3063 600
rect 3087 596 3173 603
rect 3367 596 3393 603
rect 3586 600 3587 607
rect 3608 596 3653 603
rect 3747 596 3793 603
rect 3867 596 4113 603
rect 4127 596 4313 603
rect 4713 603 4727 613
rect 4713 600 4793 603
rect 4716 596 4793 600
rect 4807 593 4812 607
rect 4833 593 4834 600
rect 5033 603 5047 613
rect 5233 607 5247 613
rect 5287 613 5293 626
rect 5416 623 5423 636
rect 5553 627 5567 636
rect 5347 616 5423 623
rect 5487 620 5543 623
rect 5487 616 5547 620
rect 5533 607 5547 616
rect 5596 616 5653 623
rect 5596 607 5603 616
rect 4848 600 5047 603
rect 4848 596 5043 600
rect 5056 596 5153 603
rect 647 576 843 583
rect 913 583 927 593
rect 867 580 927 583
rect 867 576 923 580
rect 987 576 1193 583
rect 2187 576 2393 583
rect 2667 576 2713 583
rect 3587 576 3673 583
rect 4833 583 4847 593
rect 4627 580 4847 583
rect 4627 576 4844 580
rect 5056 583 5063 596
rect 5233 600 5234 607
rect 5226 593 5227 600
rect 5587 596 5603 607
rect 5587 593 5600 596
rect 5213 587 5227 593
rect 4867 576 5063 583
rect 5226 580 5227 587
rect 5248 576 5573 583
rect 287 556 353 563
rect 567 556 833 563
rect 1067 556 1393 563
rect 1667 556 2373 563
rect 2627 556 2833 563
rect 2847 556 3253 563
rect 3447 556 4013 563
rect 5236 563 5243 573
rect 5047 556 5243 563
rect 5387 556 5673 563
rect 627 536 1093 543
rect 1147 536 1403 543
rect 187 516 1233 523
rect 1396 523 1403 536
rect 1487 536 2053 543
rect 2407 536 2853 543
rect 4827 536 5293 543
rect 1396 516 2573 523
rect 3027 516 3113 523
rect 4487 516 4553 523
rect 4927 516 5353 523
rect 807 496 1293 503
rect 1847 496 3092 503
rect 3128 496 3233 503
rect 4607 496 4993 503
rect 5007 496 5073 503
rect 5167 496 5213 503
rect 5227 496 5533 503
rect 907 476 1193 483
rect 1207 476 2173 483
rect 2887 476 3793 483
rect 4687 476 5233 483
rect 647 456 673 463
rect 1187 456 1253 463
rect 1327 456 1513 463
rect 1527 456 2273 463
rect 2747 456 3072 463
rect 3108 456 3633 463
rect 3767 456 3893 463
rect 4487 456 4653 463
rect 4727 456 4813 463
rect 4936 456 5473 463
rect 4936 447 4943 456
rect 227 436 732 443
rect 768 436 1453 443
rect 1987 436 2033 443
rect 2127 436 2193 443
rect 4187 436 4433 443
rect 4567 436 4633 443
rect 4647 436 4933 443
rect 4987 436 5413 443
rect 267 416 693 423
rect 847 416 1163 423
rect 1156 407 1163 416
rect 2233 423 2247 433
rect 2127 420 2247 423
rect 2127 416 2243 420
rect 2347 416 2432 423
rect 2468 416 2693 423
rect 3727 416 3893 423
rect 4335 416 4673 423
rect 116 400 183 403
rect 113 396 183 400
rect 113 387 127 396
rect 176 387 183 396
rect 533 387 547 393
rect 1036 396 1093 403
rect 187 383 200 387
rect 187 380 202 383
rect 187 373 207 380
rect 307 380 363 383
rect 307 376 367 380
rect 193 367 207 373
rect 353 367 367 376
rect 487 373 493 387
rect 607 376 753 383
rect 807 376 913 383
rect 1036 383 1043 396
rect 1107 396 1132 403
rect 1168 396 1253 403
rect 1396 400 1473 403
rect 1393 396 1473 400
rect 1393 387 1407 396
rect 1647 400 1763 403
rect 1647 396 1767 400
rect 987 376 1043 383
rect 793 367 807 373
rect 1053 367 1067 373
rect 93 347 107 353
rect 206 360 207 367
rect 228 353 233 367
rect 407 353 413 367
rect 567 353 573 367
rect 587 356 652 363
rect 688 353 693 367
rect 715 360 793 363
rect 713 356 793 360
rect 133 343 147 353
rect 313 347 327 353
rect 133 340 213 343
rect 136 336 213 340
rect 227 336 253 343
rect 367 333 373 347
rect 513 343 527 353
rect 713 347 727 356
rect 847 353 853 367
rect 1007 353 1013 367
rect 1036 356 1053 363
rect 513 340 593 343
rect 516 336 593 340
rect 646 333 647 340
rect 668 333 673 347
rect 726 340 727 347
rect 748 336 813 343
rect 867 336 893 343
rect 953 343 967 353
rect 1036 343 1043 356
rect 1307 383 1320 387
rect 1307 373 1323 383
rect 1347 373 1353 387
rect 1753 387 1767 396
rect 2247 396 2394 403
rect 2393 393 2394 396
rect 2796 396 2913 403
rect 2033 387 2047 393
rect 2393 387 2407 393
rect 2796 387 2803 396
rect 3427 396 3453 403
rect 3876 400 4213 403
rect 3873 396 4213 400
rect 3873 387 3887 396
rect 4213 387 4227 393
rect 4335 387 4342 416
rect 4767 416 5033 423
rect 5107 416 5353 423
rect 5507 416 5633 423
rect 4606 393 4607 400
rect 4593 387 4607 393
rect 4927 396 4953 403
rect 4753 387 4767 393
rect 1807 373 1813 387
rect 1867 373 1873 387
rect 1887 376 2003 383
rect 1093 367 1107 373
rect 1207 353 1213 367
rect 1267 353 1273 367
rect 1316 363 1323 373
rect 1996 367 2003 376
rect 2127 376 2153 383
rect 2207 376 2372 383
rect 2393 380 2394 387
rect 2386 373 2387 380
rect 2507 373 2513 387
rect 2567 373 2573 387
rect 2587 376 2653 383
rect 2707 373 2713 387
rect 2807 383 2820 387
rect 2807 380 2823 383
rect 2807 373 2827 380
rect 2887 380 2984 383
rect 2887 376 2987 380
rect 2373 367 2387 373
rect 2813 367 2827 373
rect 2973 367 2987 376
rect 3807 373 3813 387
rect 4027 376 4173 383
rect 4267 376 4312 383
rect 4368 373 4373 387
rect 4447 376 4473 383
rect 4527 376 4553 383
rect 4606 380 4607 387
rect 4628 373 4633 387
rect 4993 387 5007 393
rect 5327 396 5673 403
rect 5153 387 5167 393
rect 5047 373 5053 387
rect 5227 373 5233 387
rect 5307 376 5393 383
rect 3473 367 3487 373
rect 4013 367 4027 373
rect 1316 356 1373 363
rect 1527 353 1532 367
rect 1553 353 1554 360
rect 1667 353 1673 367
rect 1787 356 1833 363
rect 1927 356 1953 363
rect 1996 356 2013 367
rect 2000 353 2013 356
rect 1413 347 1427 353
rect 953 340 1043 343
rect 956 336 1043 340
rect 1087 336 1173 343
rect 1227 333 1233 347
rect 1287 336 1313 343
rect 1487 336 1533 343
rect 1553 343 1567 353
rect 1553 340 1613 343
rect 1556 336 1613 340
rect 633 327 647 333
rect 107 316 213 323
rect 547 316 632 323
rect 646 320 647 327
rect 1007 316 1073 323
rect 1556 323 1563 336
rect 1873 343 1887 353
rect 1827 340 1887 343
rect 1827 336 1883 340
rect 1956 343 1963 353
rect 2053 343 2067 353
rect 2427 353 2433 367
rect 2507 356 2553 363
rect 2607 353 2613 367
rect 2687 356 2732 363
rect 2768 353 2773 367
rect 2927 353 2932 367
rect 2973 360 2974 367
rect 2966 353 2967 360
rect 3367 356 3403 363
rect 1956 340 2067 343
rect 1956 336 2063 340
rect 2173 343 2187 353
rect 2107 340 2187 343
rect 2556 343 2563 353
rect 2953 347 2967 353
rect 3396 347 3403 356
rect 3427 353 3433 367
rect 3847 353 3853 367
rect 3907 353 3913 367
rect 3927 356 3973 363
rect 4147 356 4233 363
rect 4336 363 4343 373
rect 4287 356 4343 363
rect 4373 363 4387 373
rect 5393 367 5407 373
rect 4373 360 4472 363
rect 4376 356 4472 360
rect 4493 353 4494 360
rect 4547 356 4613 363
rect 4707 356 4733 363
rect 4827 353 4833 367
rect 4887 356 4933 363
rect 2107 336 2183 340
rect 2556 336 2713 343
rect 2807 333 2813 347
rect 2966 340 2967 347
rect 3007 333 3012 347
rect 3048 333 3053 347
rect 3127 333 3132 347
rect 3168 333 3173 347
rect 3396 336 3413 347
rect 3400 333 3413 336
rect 3507 333 3513 347
rect 3587 333 3593 347
rect 3647 333 3653 347
rect 3707 333 3713 347
rect 3967 336 3993 343
rect 4353 343 4367 353
rect 4187 340 4367 343
rect 4187 336 4363 340
rect 4493 343 4507 353
rect 4447 340 4507 343
rect 4773 343 4787 353
rect 4773 340 4833 343
rect 4447 336 4504 340
rect 4776 336 4833 340
rect 4847 333 4853 347
rect 5013 343 5027 353
rect 5147 353 5152 367
rect 5186 353 5187 360
rect 5208 356 5272 363
rect 5308 353 5313 367
rect 5433 367 5447 373
rect 5580 383 5593 387
rect 5576 380 5593 383
rect 5533 367 5547 373
rect 5573 373 5593 380
rect 5573 367 5587 373
rect 5596 360 5633 363
rect 5593 356 5633 360
rect 5133 343 5147 353
rect 5013 340 5147 343
rect 5173 343 5187 353
rect 5296 343 5303 353
rect 5593 347 5607 356
rect 5647 353 5653 367
rect 5173 340 5303 343
rect 5016 336 5143 340
rect 5175 336 5303 340
rect 5316 336 5413 343
rect 1427 316 1563 323
rect 1693 327 1707 333
rect 1896 323 1903 333
rect 1896 316 2033 323
rect 307 296 453 303
rect 1896 303 1903 316
rect 2913 323 2927 333
rect 3453 327 3467 333
rect 2707 320 2927 323
rect 2707 316 2923 320
rect 3016 316 3053 323
rect 807 296 1903 303
rect 1927 296 2073 303
rect 2313 303 2327 313
rect 3016 303 3023 316
rect 3247 316 3293 323
rect 3753 327 3767 333
rect 4033 327 4047 333
rect 4047 316 4093 323
rect 5027 316 5053 323
rect 5316 323 5323 336
rect 5467 336 5493 343
rect 5516 336 5553 343
rect 5107 316 5323 323
rect 5367 316 5393 323
rect 5516 323 5523 336
rect 5447 316 5523 323
rect 5687 313 5693 327
rect 2087 296 3023 303
rect 4627 296 4673 303
rect 4947 296 5453 303
rect 5467 296 5593 303
rect 47 276 173 283
rect 187 276 393 283
rect 407 276 613 283
rect 707 276 1333 283
rect 1696 276 2092 283
rect 1696 267 1703 276
rect 2128 276 2573 283
rect 2827 276 3033 283
rect 4567 276 4833 283
rect 4847 276 5073 283
rect 5127 276 5593 283
rect 527 256 1693 263
rect 2167 256 2473 263
rect 2967 256 3173 263
rect 4447 256 4793 263
rect 4807 256 5093 263
rect 5187 256 5713 263
rect 867 236 913 243
rect 1867 236 1973 243
rect 1987 236 2233 243
rect 2287 236 3133 243
rect 4667 236 5273 243
rect 5407 236 5453 243
rect 1167 216 1213 223
rect 1447 216 1653 223
rect 1667 216 2223 223
rect 2216 207 2223 216
rect 2407 216 2773 223
rect 5367 213 5373 227
rect 5396 216 5553 223
rect 96 200 313 203
rect 93 196 313 200
rect 93 187 107 196
rect 327 196 513 203
rect 1427 196 1453 203
rect 1467 196 1473 203
rect 1547 196 1952 203
rect 1453 187 1467 193
rect 1733 187 1747 196
rect 1973 193 1974 200
rect 2027 196 2153 203
rect 2227 196 2493 203
rect 3407 196 4953 203
rect 5396 203 5403 216
rect 5327 196 5403 203
rect 5427 196 5493 203
rect 5607 196 5643 203
rect 1973 187 1987 193
rect 5636 187 5643 196
rect 147 176 293 183
rect 436 180 653 183
rect 333 167 347 173
rect 433 176 653 180
rect 433 167 447 176
rect 727 176 993 183
rect 1007 176 1073 183
rect 1156 176 1213 183
rect 387 156 433 163
rect 487 156 553 163
rect 713 147 727 153
rect 107 136 133 143
rect 147 133 152 147
rect 188 133 193 147
rect 307 133 313 147
rect 447 133 453 147
rect 507 133 513 147
rect 527 136 573 143
rect 627 133 633 147
rect 1156 163 1163 176
rect 1256 180 1333 183
rect 1253 176 1333 180
rect 1253 167 1267 176
rect 1807 180 1883 183
rect 1807 176 1887 180
rect 887 156 1163 163
rect 1177 160 1253 163
rect 1173 156 1253 160
rect 753 147 767 153
rect 847 133 853 147
rect 907 133 913 147
rect 956 143 963 156
rect 956 136 993 143
rect 1127 133 1133 147
rect 1147 134 1152 147
rect 1173 147 1187 156
rect 1327 157 1373 164
rect 1387 154 1393 167
rect 1633 167 1647 173
rect 1387 153 1400 154
rect 1587 153 1593 167
rect 1873 167 1887 176
rect 2073 167 2087 173
rect 1927 156 2013 163
rect 2380 183 2393 187
rect 2376 180 2393 183
rect 2113 167 2127 173
rect 2373 173 2393 180
rect 2667 176 2813 183
rect 2373 167 2387 173
rect 2693 167 2707 176
rect 2867 173 2873 187
rect 3076 180 3243 183
rect 3073 176 3243 180
rect 3073 167 3087 176
rect 3236 167 3243 176
rect 3607 176 3633 183
rect 3957 180 4353 183
rect 3953 176 4353 180
rect 3333 167 3347 173
rect 3953 167 3967 176
rect 4407 176 4613 183
rect 4707 176 4773 183
rect 4787 176 4933 183
rect 5367 176 5423 183
rect 5636 176 5653 187
rect 5273 167 5287 173
rect 5416 167 5423 176
rect 5640 173 5653 176
rect 2427 156 2453 163
rect 2706 160 2707 167
rect 2728 153 2733 167
rect 2953 147 2967 153
rect 1173 140 1174 147
rect 1147 133 1160 134
rect 1227 133 1233 147
rect 1287 136 1313 143
rect 1447 133 1453 147
rect 1667 133 1673 147
rect 1787 133 1793 147
rect 1867 133 1872 147
rect 1908 133 1913 147
rect 2027 136 2093 143
rect 2147 133 2153 147
rect 2247 136 2332 143
rect 2366 133 2367 140
rect 2388 133 2393 147
rect 2416 136 2513 143
rect 353 123 367 133
rect 436 123 443 133
rect 353 120 443 123
rect 356 116 443 120
rect 507 116 593 123
rect 667 116 733 123
rect 807 113 813 127
rect 887 113 893 127
rect 1167 113 1173 127
rect 1307 116 1413 123
rect 1613 123 1627 133
rect 1427 120 1627 123
rect 1427 116 1623 120
rect 2227 113 2232 127
rect 2268 113 2273 127
rect 2353 123 2367 133
rect 2416 123 2423 136
rect 2647 136 2693 143
rect 3167 153 3173 167
rect 3227 153 3233 167
rect 3676 156 3913 163
rect 2993 147 3007 153
rect 3387 133 3393 147
rect 3487 136 3533 143
rect 3607 136 3653 143
rect 2353 120 2423 123
rect 2355 116 2423 120
rect 2467 116 2493 123
rect 2833 123 2847 133
rect 3676 127 3683 156
rect 3927 153 3932 167
rect 3953 160 3954 167
rect 4027 153 4033 167
rect 4107 153 4113 167
rect 4267 160 4303 163
rect 4267 156 4307 160
rect 4213 147 4227 153
rect 3786 133 3787 140
rect 3806 133 3807 140
rect 3828 136 3873 143
rect 3887 133 3893 147
rect 3947 133 3953 147
rect 4293 147 4307 156
rect 4587 156 4643 163
rect 4636 147 4643 156
rect 4967 156 4993 163
rect 5067 153 5073 167
rect 5327 156 5393 163
rect 5416 156 5433 167
rect 5420 153 5433 156
rect 5527 156 5573 163
rect 4793 147 4807 153
rect 5113 147 5127 153
rect 4367 136 4413 143
rect 4547 133 4552 147
rect 4586 133 4587 140
rect 4608 133 4613 147
rect 4636 136 4653 147
rect 4640 133 4653 136
rect 4847 133 4853 147
rect 4927 133 4933 147
rect 5187 136 5253 143
rect 5347 136 5413 143
rect 5567 136 5653 143
rect 3773 127 3787 133
rect 2567 120 2847 123
rect 2567 116 2843 120
rect 173 103 187 113
rect 496 103 503 113
rect 3513 107 3527 113
rect 173 100 503 103
rect 176 96 503 100
rect 1127 96 1213 103
rect 1327 96 1793 103
rect 3627 113 3633 127
rect 3696 116 3733 123
rect 3553 103 3567 113
rect 3696 103 3703 116
rect 3786 120 3787 127
rect 3793 127 3807 133
rect 4173 127 4187 133
rect 3793 120 3794 127
rect 4227 116 4273 123
rect 4273 107 4287 113
rect 4387 113 4393 127
rect 4536 123 4543 133
rect 4447 116 4543 123
rect 4573 127 4587 133
rect 5293 127 5307 133
rect 4787 116 4813 123
rect 4887 113 4893 127
rect 5453 127 5467 133
rect 4313 107 4327 113
rect 3553 100 3703 103
rect 3556 96 3703 100
rect 3787 96 4252 103
rect 4273 100 4274 107
rect 4327 96 4493 103
rect 4933 103 4947 113
rect 4933 100 4973 103
rect 4936 96 4973 100
rect 5307 96 5613 103
rect 347 76 753 83
rect 967 76 1813 83
rect 3527 76 3593 83
rect 3647 76 4113 83
rect 4287 76 4733 83
rect 5247 76 5513 83
rect 567 56 913 63
rect 1167 56 1313 63
rect 1387 56 1593 63
rect 3267 56 3633 63
rect 4187 56 4313 63
rect 267 36 853 43
rect 2967 36 3453 43
rect 4087 36 5113 43
rect 5167 36 5693 43
rect 3007 16 3093 23
rect 4547 16 5433 23
<< m3contact >>
rect 4113 5773 4127 5787
rect 4153 5773 4167 5787
rect 4273 5773 4287 5787
rect 4793 5773 4807 5787
rect 4933 5773 4947 5787
rect 5433 5773 5447 5787
rect 4013 5753 4027 5767
rect 4233 5753 4247 5767
rect 4313 5753 4327 5767
rect 1513 5733 1527 5747
rect 1893 5733 1907 5747
rect 4973 5753 4987 5767
rect 5093 5753 5107 5767
rect 5233 5753 5247 5767
rect 5553 5753 5567 5767
rect 5053 5734 5067 5748
rect 5273 5733 5287 5747
rect 5533 5733 5547 5747
rect 593 5713 607 5727
rect 1313 5713 1327 5727
rect 4733 5713 4747 5727
rect 5013 5713 5027 5727
rect 5053 5712 5067 5726
rect 613 5693 627 5707
rect 2113 5693 2127 5707
rect 2293 5693 2307 5707
rect 2933 5693 2947 5707
rect 313 5673 327 5687
rect 873 5673 887 5687
rect 1013 5673 1027 5687
rect 1613 5673 1627 5687
rect 1713 5673 1727 5687
rect 2133 5673 2147 5687
rect 2813 5673 2827 5687
rect 3233 5673 3247 5687
rect 3833 5673 3847 5687
rect 4272 5673 4286 5687
rect 793 5653 807 5667
rect 933 5653 947 5667
rect 1013 5653 1027 5667
rect 1413 5653 1427 5667
rect 1473 5653 1487 5667
rect 1553 5653 1567 5667
rect 53 5633 67 5647
rect 193 5613 207 5627
rect 313 5633 327 5647
rect 393 5633 407 5647
rect 233 5613 247 5627
rect 333 5613 347 5627
rect 514 5633 528 5647
rect 872 5633 886 5647
rect 953 5633 967 5647
rect 1073 5633 1087 5647
rect 1113 5633 1127 5647
rect 1193 5633 1207 5647
rect 1513 5633 1527 5647
rect 1612 5633 1626 5647
rect 1893 5633 1907 5647
rect 2393 5653 2407 5667
rect 2893 5653 2907 5667
rect 3413 5653 3427 5667
rect 4294 5653 4308 5667
rect 4773 5653 4787 5667
rect 5073 5653 5087 5667
rect 2132 5633 2146 5647
rect 2253 5633 2267 5647
rect 2293 5633 2307 5647
rect 2432 5633 2446 5647
rect 2493 5633 2507 5647
rect 2713 5633 2727 5647
rect 2793 5633 2807 5647
rect 2873 5633 2887 5647
rect 2953 5633 2967 5647
rect 3173 5633 3187 5647
rect 3513 5633 3527 5647
rect 3613 5633 3627 5647
rect 3753 5633 3767 5647
rect 3833 5633 3847 5647
rect 4233 5633 4247 5647
rect 4333 5633 4347 5647
rect 4433 5633 4447 5647
rect 4733 5633 4747 5647
rect 4853 5633 4867 5647
rect 4892 5633 4906 5647
rect 4934 5633 4948 5647
rect 5153 5633 5167 5647
rect 5213 5633 5227 5647
rect 5533 5633 5547 5647
rect 492 5613 506 5627
rect 612 5613 626 5627
rect 634 5613 648 5627
rect 513 5593 527 5607
rect 553 5593 567 5607
rect 693 5593 707 5607
rect 793 5613 807 5627
rect 894 5613 908 5627
rect 993 5593 1007 5607
rect 1293 5613 1307 5627
rect 1653 5613 1667 5627
rect 1213 5593 1227 5607
rect 1433 5593 1447 5607
rect 1993 5613 2007 5627
rect 2353 5613 2367 5627
rect 2513 5613 2527 5627
rect 2693 5613 2707 5627
rect 3133 5613 3147 5627
rect 3413 5613 3427 5627
rect 1933 5593 1947 5607
rect 2033 5593 2047 5607
rect 2192 5593 2206 5607
rect 2292 5593 2306 5607
rect 2393 5593 2407 5607
rect 2433 5593 2447 5607
rect 2753 5593 2767 5607
rect 2913 5593 2927 5607
rect 3793 5593 3807 5607
rect 4013 5593 4027 5607
rect 4793 5613 4807 5627
rect 5053 5613 5067 5627
rect 4213 5593 4227 5607
rect 4613 5593 4627 5607
rect 4853 5593 4867 5607
rect 5252 5613 5266 5627
rect 5274 5613 5288 5627
rect 5394 5613 5408 5627
rect 5593 5613 5607 5627
rect 5073 5593 5087 5607
rect 5372 5593 5386 5607
rect 233 5573 247 5587
rect 393 5573 407 5587
rect 893 5573 907 5587
rect 1133 5573 1147 5587
rect 1413 5573 1427 5587
rect 1653 5573 1667 5587
rect 1973 5573 1987 5587
rect 2193 5573 2207 5587
rect 2333 5573 2347 5587
rect 2853 5573 2867 5587
rect 3453 5573 3467 5587
rect 3693 5573 3707 5587
rect 3753 5573 3767 5587
rect 193 5553 207 5567
rect 333 5553 347 5567
rect 553 5553 567 5567
rect 633 5553 647 5567
rect 833 5553 847 5567
rect 953 5553 967 5567
rect 1073 5553 1087 5567
rect 1213 5553 1227 5567
rect 1613 5553 1627 5567
rect 2253 5553 2267 5567
rect 2713 5553 2727 5567
rect 3233 5553 3247 5567
rect 3853 5553 3867 5567
rect 4113 5553 4127 5567
rect 4373 5553 4387 5567
rect 4433 5553 4447 5567
rect 4833 5553 4847 5567
rect 4973 5553 4987 5567
rect 233 5533 247 5547
rect 693 5533 707 5547
rect 1193 5533 1207 5547
rect 1473 5533 1487 5547
rect 1833 5533 1847 5547
rect 2073 5533 2087 5547
rect 3613 5533 3627 5547
rect 3913 5533 3927 5547
rect 4413 5533 4427 5547
rect 4813 5533 4827 5547
rect 5053 5533 5067 5547
rect 5353 5533 5367 5547
rect 5673 5533 5687 5547
rect 513 5513 527 5527
rect 733 5513 747 5527
rect 1513 5513 1527 5527
rect 1973 5513 1987 5527
rect 3392 5513 3406 5527
rect 3414 5513 3428 5527
rect 3773 5513 3787 5527
rect 3813 5513 3827 5527
rect 4113 5513 4127 5527
rect 4213 5513 4227 5527
rect 4773 5513 4787 5527
rect 5113 5513 5127 5527
rect 5373 5513 5387 5527
rect 273 5493 287 5507
rect 473 5493 487 5507
rect 913 5493 927 5507
rect 1293 5493 1307 5507
rect 4413 5493 4427 5507
rect 4493 5493 4507 5507
rect 4733 5493 4747 5507
rect 5233 5493 5247 5507
rect 5293 5493 5307 5507
rect 5573 5493 5587 5507
rect 53 5473 67 5487
rect 673 5473 687 5487
rect 1133 5473 1147 5487
rect 1213 5473 1227 5487
rect 1573 5473 1587 5487
rect 1853 5473 1867 5487
rect 3353 5473 3367 5487
rect 3433 5473 3447 5487
rect 4153 5473 4167 5487
rect 4453 5473 4467 5487
rect 4893 5473 4907 5487
rect 5093 5473 5107 5487
rect 5133 5473 5147 5487
rect 5253 5473 5267 5487
rect 5413 5473 5427 5487
rect 5513 5473 5527 5487
rect 693 5453 707 5467
rect 753 5453 767 5467
rect 1173 5453 1187 5467
rect 1313 5453 1327 5467
rect 1553 5453 1567 5467
rect 1673 5453 1687 5467
rect 2033 5453 2047 5467
rect 2513 5453 2527 5467
rect 2693 5453 2707 5467
rect 2833 5453 2847 5467
rect 2973 5453 2987 5467
rect 3233 5453 3247 5467
rect 3373 5453 3387 5467
rect 53 5433 67 5447
rect 93 5433 107 5447
rect 532 5433 546 5447
rect 593 5433 607 5447
rect 893 5433 907 5447
rect 1233 5433 1247 5447
rect 1453 5433 1467 5447
rect 1673 5433 1687 5447
rect 153 5413 167 5427
rect 213 5413 227 5427
rect 293 5413 307 5427
rect 113 5393 127 5407
rect 353 5393 367 5407
rect 672 5413 686 5427
rect 694 5413 708 5427
rect 773 5413 787 5427
rect 833 5413 847 5427
rect 873 5413 887 5427
rect 1053 5413 1067 5427
rect 1093 5413 1107 5427
rect 1353 5413 1367 5427
rect 1393 5413 1407 5427
rect 1513 5413 1527 5427
rect 1593 5413 1607 5427
rect 1713 5433 1727 5447
rect 1853 5433 1867 5447
rect 2074 5433 2088 5447
rect 2113 5433 2127 5447
rect 3413 5453 3427 5467
rect 3873 5453 3887 5467
rect 4233 5453 4247 5467
rect 4553 5453 4567 5467
rect 4633 5453 4647 5467
rect 4813 5453 4827 5467
rect 5053 5453 5067 5467
rect 5213 5453 5227 5467
rect 5254 5453 5268 5467
rect 5413 5453 5427 5467
rect 5593 5453 5607 5467
rect 1933 5413 1947 5427
rect 2052 5413 2066 5427
rect 3173 5433 3187 5447
rect 3352 5433 3366 5447
rect 3792 5433 3806 5447
rect 3814 5433 3828 5447
rect 4234 5433 4248 5447
rect 4413 5433 4427 5447
rect 4452 5433 4466 5447
rect 4732 5433 4746 5447
rect 2373 5413 2387 5427
rect 2414 5413 2428 5427
rect 2773 5413 2787 5427
rect 2833 5413 2847 5427
rect 3113 5413 3127 5427
rect 713 5393 727 5407
rect 1053 5393 1067 5407
rect 353 5373 367 5387
rect 393 5373 407 5387
rect 533 5373 547 5387
rect 773 5373 787 5387
rect 913 5373 927 5387
rect 1093 5373 1107 5387
rect 1133 5373 1147 5387
rect 1293 5393 1307 5407
rect 1453 5393 1467 5407
rect 1493 5393 1507 5407
rect 1613 5393 1627 5407
rect 1973 5393 1987 5407
rect 1173 5373 1187 5387
rect 1833 5373 1847 5387
rect 2153 5393 2167 5407
rect 2194 5393 2208 5407
rect 2673 5393 2687 5407
rect 2713 5393 2727 5407
rect 2813 5393 2827 5407
rect 2894 5393 2908 5407
rect 2973 5373 2987 5387
rect 5093 5433 5107 5447
rect 5173 5433 5187 5447
rect 5353 5433 5367 5447
rect 5493 5433 5507 5447
rect 3193 5393 3207 5407
rect 3234 5393 3248 5407
rect 3553 5413 3567 5427
rect 3634 5413 3648 5427
rect 3433 5393 3447 5407
rect 3772 5393 3786 5407
rect 3813 5394 3827 5408
rect 3893 5393 3907 5407
rect 3973 5413 3987 5427
rect 4212 5413 4226 5427
rect 4612 5413 4626 5427
rect 4873 5414 4887 5428
rect 4933 5413 4947 5427
rect 5033 5413 5047 5427
rect 5253 5413 5267 5427
rect 5552 5413 5566 5427
rect 5634 5413 5648 5427
rect 3933 5393 3947 5407
rect 4493 5393 4507 5407
rect 3752 5373 3766 5387
rect 3813 5372 3827 5386
rect 3893 5373 3907 5387
rect 4033 5373 4047 5387
rect 4873 5392 4887 5406
rect 5413 5393 5427 5407
rect 4653 5373 4667 5387
rect 4733 5373 4747 5387
rect 5033 5373 5047 5387
rect 5133 5373 5147 5387
rect 5673 5393 5687 5407
rect 5653 5373 5667 5387
rect 413 5353 427 5367
rect 1173 5353 1187 5367
rect 1553 5353 1567 5367
rect 1993 5353 2007 5367
rect 2213 5353 2227 5367
rect 3073 5353 3087 5367
rect 3513 5353 3527 5367
rect 3653 5353 3667 5367
rect 3973 5353 3987 5367
rect 4693 5353 4707 5367
rect 4853 5353 4867 5367
rect 5213 5353 5227 5367
rect 1113 5333 1127 5347
rect 873 5313 887 5327
rect 993 5313 1007 5327
rect 1393 5333 1407 5347
rect 1433 5333 1447 5347
rect 2053 5333 2067 5347
rect 3133 5333 3147 5347
rect 3553 5333 3567 5347
rect 4893 5333 4907 5347
rect 4933 5333 4947 5347
rect 5593 5333 5607 5347
rect 1293 5313 1307 5327
rect 1373 5313 1387 5327
rect 1953 5313 1967 5327
rect 2893 5313 2907 5327
rect 3193 5313 3207 5327
rect 3413 5313 3427 5327
rect 3854 5313 3868 5327
rect 4153 5313 4167 5327
rect 4553 5313 4567 5327
rect 4853 5313 4867 5327
rect 5093 5313 5107 5327
rect 5433 5313 5447 5327
rect 5553 5313 5567 5327
rect 753 5293 767 5307
rect 893 5293 907 5307
rect 1213 5293 1227 5307
rect 1593 5293 1607 5307
rect 3893 5293 3907 5307
rect 3973 5293 3987 5307
rect 4213 5293 4227 5307
rect 4592 5293 4606 5307
rect 4614 5293 4628 5307
rect 4873 5293 4887 5307
rect 1493 5273 1507 5287
rect 1753 5273 1767 5287
rect 2713 5273 2727 5287
rect 3033 5273 3047 5287
rect 3573 5273 3587 5287
rect 3873 5273 3887 5287
rect 4373 5273 4387 5287
rect 4733 5273 4747 5287
rect 5433 5273 5447 5287
rect 113 5253 127 5267
rect 953 5253 967 5267
rect 1233 5253 1247 5267
rect 2333 5253 2347 5267
rect 3853 5253 3867 5267
rect 93 5233 107 5247
rect 1133 5233 1147 5247
rect 1293 5233 1307 5247
rect 1433 5233 1447 5247
rect 1933 5233 1947 5247
rect 2113 5233 2127 5247
rect 2373 5233 2387 5247
rect 2993 5233 3007 5247
rect 3753 5233 3767 5247
rect 3933 5234 3947 5248
rect 4294 5233 4308 5247
rect 5133 5233 5147 5247
rect 133 5213 147 5227
rect 333 5213 347 5227
rect 473 5213 487 5227
rect 1333 5213 1347 5227
rect 1693 5213 1707 5227
rect 2213 5213 2227 5227
rect 2273 5213 2287 5227
rect 2353 5213 2367 5227
rect 2673 5213 2687 5227
rect 2873 5213 2887 5227
rect 3373 5213 3387 5227
rect 3693 5213 3707 5227
rect 3933 5212 3947 5226
rect 5493 5213 5507 5227
rect 773 5193 787 5207
rect 1113 5193 1127 5207
rect 1233 5193 1247 5207
rect 1553 5193 1567 5207
rect 1773 5193 1787 5207
rect 1833 5193 1847 5207
rect 1873 5193 1887 5207
rect 73 5173 87 5187
rect 173 5173 187 5187
rect 253 5173 267 5187
rect 333 5173 347 5187
rect 73 5153 87 5167
rect 573 5173 587 5187
rect 774 5173 788 5187
rect 1293 5173 1307 5187
rect 1373 5173 1387 5187
rect 1473 5173 1487 5187
rect 133 5133 147 5147
rect 293 5133 307 5147
rect 433 5133 447 5147
rect 473 5153 487 5167
rect 613 5153 627 5167
rect 752 5153 766 5167
rect 672 5133 686 5147
rect 892 5153 906 5167
rect 973 5153 987 5167
rect 1413 5153 1427 5167
rect 1874 5173 1888 5187
rect 1574 5153 1588 5167
rect 1713 5153 1727 5167
rect 1773 5153 1787 5167
rect 153 5113 167 5127
rect 353 5113 367 5127
rect 433 5113 447 5127
rect 793 5113 807 5127
rect 1033 5133 1047 5147
rect 1113 5133 1127 5147
rect 1194 5133 1208 5147
rect 1473 5133 1487 5147
rect 2393 5173 2407 5187
rect 2433 5193 2447 5207
rect 2633 5173 2647 5187
rect 2873 5193 2887 5207
rect 2974 5173 2988 5187
rect 3193 5173 3207 5187
rect 3293 5173 3307 5187
rect 3953 5193 3967 5207
rect 4232 5193 4246 5207
rect 4333 5193 4347 5207
rect 3513 5173 3527 5187
rect 1933 5153 1947 5167
rect 2013 5153 2027 5167
rect 2133 5153 2147 5167
rect 2473 5153 2487 5167
rect 2613 5153 2627 5167
rect 1553 5133 1567 5147
rect 1593 5133 1607 5147
rect 1753 5133 1767 5147
rect 1913 5133 1927 5147
rect 2053 5133 2067 5147
rect 2213 5133 2227 5147
rect 2293 5133 2307 5147
rect 2352 5133 2366 5147
rect 2433 5133 2447 5147
rect 853 5113 867 5127
rect 1073 5113 1087 5127
rect 793 5093 807 5107
rect 1174 5113 1188 5127
rect 2133 5113 2147 5127
rect 2313 5113 2327 5127
rect 2393 5113 2407 5127
rect 3033 5153 3047 5167
rect 3233 5153 3247 5167
rect 3333 5153 3347 5167
rect 3714 5153 3728 5167
rect 4194 5173 4208 5187
rect 4493 5173 4507 5187
rect 4633 5173 4647 5187
rect 5033 5173 5047 5187
rect 5093 5173 5107 5187
rect 4172 5153 4186 5167
rect 2953 5133 2967 5147
rect 3113 5133 3127 5147
rect 3293 5133 3307 5147
rect 3394 5133 3408 5147
rect 3453 5133 3467 5147
rect 3593 5133 3607 5147
rect 3692 5134 3706 5148
rect 4354 5153 4368 5167
rect 4574 5153 4588 5167
rect 4693 5153 4707 5167
rect 4793 5153 4807 5167
rect 4973 5153 4987 5167
rect 5133 5153 5147 5167
rect 5433 5153 5447 5167
rect 5513 5153 5527 5167
rect 5633 5153 5647 5167
rect 3753 5133 3767 5147
rect 3833 5133 3847 5147
rect 3993 5133 4007 5147
rect 4093 5133 4107 5147
rect 4154 5133 4168 5147
rect 4233 5133 4247 5147
rect 4293 5133 4307 5147
rect 4453 5133 4467 5147
rect 2593 5113 2607 5127
rect 3233 5113 3247 5127
rect 3353 5113 3367 5127
rect 3433 5113 3447 5127
rect 1453 5093 1467 5107
rect 1573 5093 1587 5107
rect 1713 5093 1727 5107
rect 2133 5093 2147 5107
rect 3693 5112 3707 5126
rect 3893 5113 3907 5127
rect 4053 5113 4067 5127
rect 2493 5093 2507 5107
rect 3633 5093 3647 5107
rect 4653 5133 4667 5147
rect 4913 5133 4927 5147
rect 4873 5113 4887 5127
rect 5013 5113 5027 5127
rect 5253 5113 5267 5127
rect 5493 5113 5507 5127
rect 4093 5093 4107 5107
rect 4153 5093 4167 5107
rect 4393 5093 4407 5107
rect 4593 5093 4607 5107
rect 4733 5093 4747 5107
rect 4773 5093 4787 5107
rect 4993 5093 5007 5107
rect 5053 5093 5067 5107
rect 5593 5093 5607 5107
rect 93 5073 107 5087
rect 233 5073 247 5087
rect 673 5073 687 5087
rect 773 5073 787 5087
rect 1833 5073 1847 5087
rect 1913 5073 1927 5087
rect 2273 5073 2287 5087
rect 3353 5073 3367 5087
rect 3673 5073 3687 5087
rect 3992 5073 4006 5087
rect 4014 5073 4028 5087
rect 413 5053 427 5067
rect 1293 5053 1307 5067
rect 2813 5053 2827 5067
rect 3133 5053 3147 5067
rect 3813 5053 3827 5067
rect 3893 5053 3907 5067
rect 4193 5053 4207 5067
rect 4273 5053 4287 5067
rect 4433 5053 4447 5067
rect 4793 5074 4807 5088
rect 5013 5073 5027 5087
rect 5413 5073 5427 5087
rect 5593 5073 5607 5087
rect 4793 5052 4807 5066
rect 4853 5053 4867 5067
rect 5153 5053 5167 5067
rect 733 5033 747 5047
rect 853 5033 867 5047
rect 1393 5033 1407 5047
rect 2773 5033 2787 5047
rect 3433 5033 3447 5047
rect 3933 5033 3947 5047
rect 4233 5033 4247 5047
rect 4713 5033 4727 5047
rect 4833 5033 4847 5047
rect 193 5013 207 5027
rect 613 5013 627 5027
rect 1173 5013 1187 5027
rect 2653 5013 2667 5027
rect 2793 5013 2807 5027
rect 2893 5013 2907 5027
rect 4293 5013 4307 5027
rect 4393 5013 4407 5027
rect 4513 5013 4527 5027
rect 313 4993 327 5007
rect 1053 4993 1067 5007
rect 1133 4993 1147 5007
rect 2093 4993 2107 5007
rect 2313 4993 2327 5007
rect 2393 4993 2407 5007
rect 3353 4993 3367 5007
rect 3393 4993 3407 5007
rect 3753 4993 3767 5007
rect 3953 4993 3967 5007
rect 4093 4993 4107 5007
rect 4633 5013 4647 5027
rect 4793 5013 4807 5027
rect 5093 5033 5107 5047
rect 5553 5033 5567 5047
rect 5693 5033 5707 5047
rect 5213 5013 5227 5027
rect 5293 5013 5307 5027
rect 4613 4993 4627 5007
rect 4713 4993 4727 5007
rect 5333 4993 5347 5007
rect 5713 4993 5727 5007
rect 153 4973 167 4987
rect 173 4953 187 4967
rect 33 4933 47 4947
rect 73 4933 87 4947
rect 212 4933 226 4947
rect 332 4953 346 4967
rect 393 4953 407 4967
rect 873 4973 887 4987
rect 1073 4973 1087 4987
rect 1333 4973 1347 4987
rect 2133 4973 2147 4987
rect 2793 4973 2807 4987
rect 493 4953 507 4967
rect 573 4953 587 4967
rect 633 4953 647 4967
rect 973 4953 987 4967
rect 373 4933 387 4947
rect 473 4933 487 4947
rect 553 4933 567 4947
rect 613 4933 627 4947
rect 713 4933 727 4947
rect 972 4933 986 4947
rect 1013 4933 1027 4947
rect 1393 4953 1407 4967
rect 1153 4933 1167 4947
rect 1493 4933 1507 4947
rect 1713 4953 1727 4967
rect 1533 4933 1547 4947
rect 1713 4933 1727 4947
rect 2093 4953 2107 4967
rect 2173 4953 2187 4967
rect 2234 4953 2248 4967
rect 2274 4953 2288 4967
rect 2392 4953 2406 4967
rect 3473 4973 3487 4987
rect 2652 4953 2666 4967
rect 2692 4953 2706 4967
rect 2773 4953 2787 4967
rect 2893 4953 2907 4967
rect 2974 4953 2988 4967
rect 3232 4953 3246 4967
rect 3393 4953 3407 4967
rect 3593 4973 3607 4987
rect 3893 4973 3907 4987
rect 4172 4973 4186 4987
rect 4233 4973 4247 4987
rect 4392 4973 4406 4987
rect 4473 4973 4487 4987
rect 4512 4973 4526 4987
rect 4573 4973 4587 4987
rect 5153 4973 5167 4987
rect 5553 4973 5567 4987
rect 73 4893 87 4907
rect 173 4913 187 4927
rect 353 4913 367 4927
rect 674 4913 688 4927
rect 113 4893 127 4907
rect 513 4893 527 4907
rect 652 4893 666 4907
rect 773 4913 787 4927
rect 1053 4913 1067 4927
rect 1373 4893 1387 4907
rect 1573 4913 1587 4927
rect 1753 4913 1767 4927
rect 1852 4913 1866 4927
rect 2013 4933 2027 4947
rect 2613 4933 2627 4947
rect 2913 4933 2927 4947
rect 3353 4933 3367 4947
rect 3513 4933 3527 4947
rect 3873 4953 3887 4967
rect 4112 4953 4126 4967
rect 4492 4953 4506 4967
rect 4793 4953 4807 4967
rect 3553 4933 3567 4947
rect 3753 4933 3767 4947
rect 3933 4933 3947 4947
rect 2073 4913 2087 4927
rect 2133 4913 2147 4927
rect 2593 4913 2607 4927
rect 2673 4913 2687 4927
rect 2853 4913 2867 4927
rect 1413 4893 1427 4907
rect 1613 4893 1627 4907
rect 1853 4893 1867 4907
rect 2373 4893 2387 4907
rect 2433 4893 2447 4907
rect 3053 4893 3067 4907
rect 3453 4913 3467 4927
rect 3653 4913 3667 4927
rect 3973 4913 3987 4927
rect 4073 4913 4087 4927
rect 4293 4933 4307 4947
rect 4433 4933 4447 4947
rect 4553 4933 4567 4947
rect 4693 4933 4707 4947
rect 4733 4933 4747 4947
rect 4853 4933 4867 4947
rect 5313 4953 5327 4967
rect 5413 4953 5427 4967
rect 5194 4933 5208 4947
rect 5433 4933 5447 4947
rect 5472 4933 5486 4947
rect 4233 4913 4247 4927
rect 4633 4913 4647 4927
rect 5393 4913 5407 4927
rect 5494 4913 5508 4927
rect 5593 4913 5607 4927
rect 3093 4893 3107 4907
rect 3473 4893 3487 4907
rect 3773 4893 3787 4907
rect 3993 4893 4007 4907
rect 4113 4893 4127 4907
rect 4173 4893 4187 4907
rect 4393 4893 4407 4907
rect 4433 4893 4447 4907
rect 193 4873 207 4887
rect 313 4873 327 4887
rect 713 4873 727 4887
rect 1013 4873 1027 4887
rect 1153 4873 1167 4887
rect 1493 4873 1507 4887
rect 2233 4873 2247 4887
rect 3033 4873 3047 4887
rect 3753 4873 3767 4887
rect 4153 4873 4167 4887
rect 4553 4873 4567 4887
rect 5053 4893 5067 4907
rect 5493 4893 5507 4907
rect 5613 4893 5627 4907
rect 5033 4873 5047 4887
rect 5093 4873 5107 4887
rect 5593 4873 5607 4887
rect 5633 4873 5647 4887
rect 393 4853 407 4867
rect 453 4853 467 4867
rect 2173 4853 2187 4867
rect 2473 4853 2487 4867
rect 2793 4853 2807 4867
rect 2993 4853 3007 4867
rect 3153 4853 3167 4867
rect 4032 4853 4046 4867
rect 4054 4853 4068 4867
rect 5133 4853 5147 4867
rect 5373 4854 5387 4868
rect 73 4833 87 4847
rect 153 4833 167 4847
rect 533 4833 547 4847
rect 673 4833 687 4847
rect 1733 4833 1747 4847
rect 2493 4833 2507 4847
rect 2833 4833 2847 4847
rect 2873 4833 2887 4847
rect 2953 4833 2967 4847
rect 3213 4833 3227 4847
rect 3493 4833 3507 4847
rect 4113 4833 4127 4847
rect 4493 4833 4507 4847
rect 4733 4833 4747 4847
rect 53 4813 67 4827
rect 473 4813 487 4827
rect 613 4813 627 4827
rect 693 4813 707 4827
rect 1373 4813 1387 4827
rect 1573 4813 1587 4827
rect 5373 4832 5387 4846
rect 5473 4833 5487 4847
rect 2933 4813 2947 4827
rect 3633 4813 3647 4827
rect 3953 4813 3967 4827
rect 3993 4813 4007 4827
rect 4333 4813 4347 4827
rect 4473 4813 4487 4827
rect 4653 4813 4667 4827
rect 1953 4793 1967 4807
rect 2193 4793 2207 4807
rect 2753 4793 2767 4807
rect 2913 4793 2927 4807
rect 3053 4793 3067 4807
rect 3233 4793 3247 4807
rect 3393 4793 3407 4807
rect 3573 4793 3587 4807
rect 3613 4793 3627 4807
rect 3693 4793 3707 4807
rect 4073 4793 4087 4807
rect 4293 4793 4307 4807
rect 4493 4793 4507 4807
rect 5513 4813 5527 4827
rect 653 4773 667 4787
rect 1453 4773 1467 4787
rect 2593 4773 2607 4787
rect 2693 4773 2707 4787
rect 2772 4773 2786 4787
rect 2794 4773 2808 4787
rect 2833 4773 2847 4787
rect 3213 4773 3227 4787
rect 3793 4773 3807 4787
rect 4093 4773 4107 4787
rect 4153 4773 4167 4787
rect 4273 4773 4287 4787
rect 4573 4773 4587 4787
rect 4873 4793 4887 4807
rect 4733 4773 4747 4787
rect 5033 4773 5047 4787
rect 353 4753 367 4767
rect 613 4753 627 4767
rect 753 4753 767 4767
rect 833 4753 847 4767
rect 2673 4753 2687 4767
rect 4013 4753 4027 4767
rect 793 4733 807 4747
rect 933 4733 947 4747
rect 1193 4733 1207 4747
rect 1293 4733 1307 4747
rect 1593 4733 1607 4747
rect 1953 4733 1967 4747
rect 2153 4733 2167 4747
rect 2453 4733 2467 4747
rect 2933 4733 2947 4747
rect 3453 4733 3467 4747
rect 3733 4733 3747 4747
rect 3953 4733 3967 4747
rect 4053 4733 4067 4747
rect 113 4713 127 4727
rect 634 4713 648 4727
rect 333 4693 347 4707
rect 612 4693 626 4707
rect 753 4693 767 4707
rect 1173 4693 1187 4707
rect 1253 4693 1267 4707
rect 1453 4693 1467 4707
rect 1592 4693 1606 4707
rect 1793 4693 1807 4707
rect 3013 4713 3027 4727
rect 3193 4713 3207 4727
rect 3253 4713 3267 4727
rect 3293 4713 3307 4727
rect 3373 4713 3387 4727
rect 3933 4713 3947 4727
rect 2012 4693 2026 4707
rect 2034 4693 2048 4707
rect 53 4673 67 4687
rect 153 4673 167 4687
rect 214 4673 228 4687
rect 372 4673 386 4687
rect 413 4673 427 4687
rect 553 4673 567 4687
rect 93 4653 107 4667
rect 333 4653 347 4667
rect 453 4653 467 4667
rect 653 4653 667 4667
rect 812 4673 826 4687
rect 834 4673 848 4687
rect 953 4673 967 4687
rect 1113 4673 1127 4687
rect 1193 4672 1207 4686
rect 1273 4673 1287 4687
rect 73 4613 87 4627
rect 373 4633 387 4647
rect 934 4652 948 4666
rect 1333 4653 1347 4667
rect 1393 4653 1407 4667
rect 1653 4673 1667 4687
rect 1912 4673 1926 4687
rect 2113 4673 2127 4687
rect 2413 4673 2427 4687
rect 2533 4673 2547 4687
rect 2614 4673 2628 4687
rect 2653 4673 2667 4687
rect 2713 4673 2727 4687
rect 1712 4653 1726 4667
rect 1752 4653 1766 4667
rect 2014 4653 2028 4667
rect 2074 4653 2088 4667
rect 513 4633 527 4647
rect 1333 4633 1347 4647
rect 1494 4633 1508 4647
rect 1713 4633 1727 4647
rect 1853 4633 1867 4647
rect 2113 4633 2127 4647
rect 2352 4653 2366 4667
rect 2393 4653 2407 4667
rect 2433 4653 2447 4667
rect 2973 4693 2987 4707
rect 3113 4693 3127 4707
rect 3173 4693 3187 4707
rect 3213 4693 3227 4707
rect 3314 4693 3328 4707
rect 3413 4693 3427 4707
rect 3773 4693 3787 4707
rect 4133 4693 4147 4707
rect 4493 4693 4507 4707
rect 4573 4693 4587 4707
rect 4953 4693 4967 4707
rect 5073 4693 5087 4707
rect 2793 4674 2807 4688
rect 2913 4673 2927 4687
rect 3093 4673 3107 4687
rect 3433 4673 3447 4687
rect 3493 4673 3507 4687
rect 3593 4673 3607 4687
rect 2813 4653 2827 4667
rect 2973 4653 2987 4667
rect 3813 4673 3827 4687
rect 3973 4673 3987 4687
rect 4093 4673 4107 4687
rect 4313 4673 4327 4687
rect 4553 4673 4567 4687
rect 4633 4673 4647 4687
rect 4833 4673 4847 4687
rect 5393 4673 5407 4687
rect 5553 4673 5567 4687
rect 3453 4653 3467 4667
rect 3733 4653 3747 4667
rect 3932 4653 3946 4667
rect 4173 4653 4187 4667
rect 4233 4653 4247 4667
rect 4453 4653 4467 4667
rect 4693 4653 4707 4667
rect 4893 4653 4907 4667
rect 5173 4653 5187 4667
rect 5273 4653 5287 4667
rect 5514 4653 5528 4667
rect 5633 4653 5647 4667
rect 2913 4633 2927 4647
rect 3013 4633 3027 4647
rect 3133 4633 3147 4647
rect 3213 4633 3227 4647
rect 3413 4633 3427 4647
rect 3553 4633 3567 4647
rect 333 4613 347 4627
rect 413 4613 427 4627
rect 553 4613 567 4627
rect 653 4613 667 4627
rect 1633 4613 1647 4627
rect 1753 4613 1767 4627
rect 2693 4613 2707 4627
rect 3433 4613 3447 4627
rect 3773 4633 3787 4647
rect 4033 4633 4047 4647
rect 4353 4633 4367 4647
rect 4473 4633 4487 4647
rect 4613 4633 4627 4647
rect 4793 4633 4807 4647
rect 5093 4633 5107 4647
rect 5253 4633 5267 4647
rect 5433 4633 5447 4647
rect 3653 4613 3667 4627
rect 3793 4613 3807 4627
rect 4493 4613 4507 4627
rect 4693 4613 4707 4627
rect 5173 4613 5187 4627
rect 5313 4613 5327 4627
rect 5393 4613 5407 4627
rect 613 4593 627 4607
rect 753 4593 767 4607
rect 973 4593 987 4607
rect 1093 4593 1107 4607
rect 1233 4593 1247 4607
rect 1653 4593 1667 4607
rect 1893 4593 1907 4607
rect 2073 4593 2087 4607
rect 2413 4593 2427 4607
rect 2873 4593 2887 4607
rect 2933 4593 2947 4607
rect 3893 4593 3907 4607
rect 4533 4593 4547 4607
rect 1613 4573 1627 4587
rect 1693 4573 1707 4587
rect 2293 4573 2307 4587
rect 3373 4573 3387 4587
rect 4193 4573 4207 4587
rect 4293 4573 4307 4587
rect 4353 4573 4367 4587
rect 4593 4573 4607 4587
rect 4773 4593 4787 4607
rect 4833 4593 4847 4607
rect 5333 4593 5347 4607
rect 5173 4573 5187 4587
rect 5513 4573 5527 4587
rect 513 4553 527 4567
rect 993 4553 1007 4567
rect 1633 4553 1647 4567
rect 1753 4553 1767 4567
rect 2353 4553 2367 4567
rect 2753 4553 2767 4567
rect 2973 4553 2987 4567
rect 3313 4553 3327 4567
rect 3573 4553 3587 4567
rect 4033 4553 4047 4567
rect 4533 4554 4547 4568
rect 4673 4553 4687 4567
rect 4733 4553 4747 4567
rect 4793 4553 4807 4567
rect 5113 4553 5127 4567
rect 5333 4553 5347 4567
rect 5373 4553 5387 4567
rect 5553 4553 5567 4567
rect 93 4533 107 4547
rect 713 4533 727 4547
rect 933 4533 947 4547
rect 1073 4533 1087 4547
rect 1333 4533 1347 4547
rect 1533 4533 1547 4547
rect 1733 4533 1747 4547
rect 1913 4533 1927 4547
rect 2433 4533 2447 4547
rect 2913 4533 2927 4547
rect 233 4513 247 4527
rect 133 4493 147 4507
rect 373 4513 387 4527
rect 593 4513 607 4527
rect 993 4513 1007 4527
rect 1133 4513 1147 4527
rect 2053 4513 2067 4527
rect 2613 4513 2627 4527
rect 2693 4513 2707 4527
rect 2733 4513 2747 4527
rect 2973 4513 2987 4527
rect 3073 4513 3087 4527
rect 3133 4513 3147 4527
rect 3353 4513 3367 4527
rect 4133 4533 4147 4547
rect 4533 4532 4547 4546
rect 4693 4533 4707 4547
rect 4753 4533 4767 4547
rect 3673 4513 3687 4527
rect 3953 4513 3967 4527
rect 4253 4513 4267 4527
rect 653 4493 667 4507
rect 1073 4493 1087 4507
rect 1213 4493 1227 4507
rect 1273 4493 1287 4507
rect 1493 4493 1507 4507
rect 1553 4493 1567 4507
rect 1653 4493 1667 4507
rect 2433 4493 2447 4507
rect 2912 4493 2926 4507
rect 2993 4493 3007 4507
rect 73 4473 87 4487
rect 273 4474 287 4488
rect 33 4453 47 4467
rect 212 4453 226 4467
rect 293 4453 307 4467
rect 353 4453 367 4467
rect 393 4453 407 4467
rect 493 4473 507 4487
rect 613 4473 627 4487
rect 653 4473 667 4487
rect 713 4473 727 4487
rect 753 4473 767 4487
rect 993 4473 1007 4487
rect 1133 4473 1147 4487
rect 1273 4473 1287 4487
rect 1753 4473 1767 4487
rect 1793 4473 1807 4487
rect 1852 4473 1866 4487
rect 933 4453 947 4467
rect 1073 4453 1087 4467
rect 1213 4453 1227 4467
rect 1472 4453 1486 4467
rect 1613 4453 1627 4467
rect 1654 4453 1668 4467
rect 1693 4453 1707 4467
rect 1913 4453 1927 4467
rect 2113 4473 2127 4487
rect 2313 4473 2327 4487
rect 2513 4474 2527 4488
rect 2593 4473 2607 4487
rect 2692 4473 2706 4487
rect 2733 4473 2747 4487
rect 3033 4493 3047 4507
rect 3333 4493 3347 4507
rect 3653 4493 3667 4507
rect 3973 4493 3987 4507
rect 4173 4493 4187 4507
rect 4213 4493 4227 4507
rect 4433 4513 4447 4527
rect 4833 4513 4847 4527
rect 4973 4513 4987 4527
rect 5053 4513 5067 4527
rect 5213 4513 5227 4527
rect 4314 4493 4328 4507
rect 5153 4493 5167 4507
rect 3053 4473 3067 4487
rect 3093 4473 3107 4487
rect 3212 4473 3226 4487
rect 3253 4473 3267 4487
rect 3373 4473 3387 4487
rect 3672 4473 3686 4487
rect 3713 4473 3727 4487
rect 3893 4473 3907 4487
rect 3952 4473 3966 4487
rect 4053 4473 4067 4487
rect 4292 4473 4306 4487
rect 4612 4473 4626 4487
rect 4693 4473 4707 4487
rect 4734 4473 4748 4487
rect 4873 4473 4887 4487
rect 2254 4453 2268 4467
rect 2413 4453 2427 4467
rect 2533 4453 2547 4467
rect 2632 4453 2646 4467
rect 2773 4453 2787 4467
rect 3152 4453 3166 4467
rect 3193 4453 3207 4467
rect 3233 4453 3247 4467
rect 3333 4453 3347 4467
rect 3453 4453 3467 4467
rect 3553 4453 3567 4467
rect 3653 4453 3667 4467
rect 3793 4453 3807 4467
rect 4314 4453 4328 4467
rect 4593 4453 4607 4467
rect 133 4433 147 4447
rect 234 4433 248 4447
rect 353 4433 367 4447
rect 433 4433 447 4447
rect 593 4433 607 4447
rect 993 4433 1007 4447
rect 1153 4433 1167 4447
rect 1392 4433 1406 4447
rect 1453 4433 1467 4447
rect 1953 4433 1967 4447
rect 1992 4433 2006 4447
rect 2232 4433 2246 4447
rect 2693 4433 2707 4447
rect 2733 4433 2747 4447
rect 2833 4433 2847 4447
rect 3513 4433 3527 4447
rect 3832 4433 3846 4447
rect 4213 4433 4227 4447
rect 4533 4433 4547 4447
rect 4633 4453 4647 4467
rect 5172 4473 5186 4487
rect 5194 4473 5208 4487
rect 5313 4473 5327 4487
rect 5473 4473 5487 4487
rect 5573 4473 5587 4487
rect 5033 4453 5047 4467
rect 5074 4453 5088 4467
rect 5253 4453 5267 4467
rect 5373 4453 5387 4467
rect 5453 4453 5467 4467
rect 4713 4433 4727 4447
rect 4753 4433 4767 4447
rect 4913 4433 4927 4447
rect 5013 4433 5027 4447
rect 5473 4433 5487 4447
rect 253 4413 267 4427
rect 492 4413 506 4427
rect 514 4413 528 4427
rect 633 4413 647 4427
rect 693 4413 707 4427
rect 1933 4413 1947 4427
rect 1073 4393 1087 4407
rect 1913 4393 1927 4407
rect 2053 4393 2067 4407
rect 2373 4413 2387 4427
rect 2553 4413 2567 4427
rect 2593 4413 2607 4427
rect 2633 4413 2647 4427
rect 3233 4413 3247 4427
rect 3933 4413 3947 4427
rect 3993 4413 4007 4427
rect 4433 4413 4447 4427
rect 4593 4413 4607 4427
rect 4913 4413 4927 4427
rect 5033 4413 5047 4427
rect 5433 4413 5447 4427
rect 5613 4413 5627 4427
rect 2233 4394 2247 4408
rect 2693 4393 2707 4407
rect 2833 4393 2847 4407
rect 3273 4393 3287 4407
rect 3413 4393 3427 4407
rect 3833 4393 3847 4407
rect 3913 4393 3927 4407
rect 4053 4393 4067 4407
rect 2013 4373 2027 4387
rect 2233 4372 2247 4386
rect 2293 4373 2307 4387
rect 2513 4373 2527 4387
rect 3093 4373 3107 4387
rect 4333 4373 4347 4387
rect 4393 4373 4407 4387
rect 4433 4373 4447 4387
rect 4473 4373 4487 4387
rect 973 4353 987 4367
rect 1133 4353 1147 4367
rect 1913 4353 1927 4367
rect 2633 4353 2647 4367
rect 2673 4353 2687 4367
rect 2873 4353 2887 4367
rect 3653 4353 3667 4367
rect 3793 4353 3807 4367
rect 1933 4333 1947 4347
rect 2253 4333 2267 4347
rect 2413 4333 2427 4347
rect 3053 4333 3067 4347
rect 4493 4353 4507 4367
rect 4573 4353 4587 4367
rect 4693 4353 4707 4367
rect 4793 4353 4807 4367
rect 5413 4353 5427 4367
rect 5653 4353 5667 4367
rect 473 4313 487 4327
rect 733 4313 747 4327
rect 1573 4313 1587 4327
rect 2513 4313 2527 4327
rect 2953 4313 2967 4327
rect 4013 4333 4027 4347
rect 4673 4333 4687 4347
rect 3673 4313 3687 4327
rect 3753 4313 3767 4327
rect 4373 4313 4387 4327
rect 4553 4313 4567 4327
rect 4633 4313 4647 4327
rect 5013 4333 5027 4347
rect 5073 4333 5087 4347
rect 4733 4313 4747 4327
rect 4873 4313 4887 4327
rect 5033 4313 5047 4327
rect 5273 4313 5287 4327
rect 273 4293 287 4307
rect 1693 4293 1707 4307
rect 2073 4293 2087 4307
rect 2373 4293 2387 4307
rect 2733 4293 2747 4307
rect 3053 4293 3067 4307
rect 5253 4293 5267 4307
rect 5593 4293 5607 4307
rect 393 4273 407 4287
rect 513 4273 527 4287
rect 613 4273 627 4287
rect 1533 4273 1547 4287
rect 3413 4273 3427 4287
rect 3493 4273 3507 4287
rect 253 4253 267 4267
rect 853 4253 867 4267
rect 1753 4253 1767 4267
rect 1833 4253 1847 4267
rect 2153 4253 2167 4267
rect 2373 4253 2387 4267
rect 2833 4253 2847 4267
rect 3153 4253 3167 4267
rect 5213 4253 5227 4267
rect 5373 4253 5387 4267
rect 93 4233 107 4247
rect 253 4233 267 4247
rect 93 4213 107 4227
rect 173 4213 187 4227
rect 353 4233 367 4247
rect 473 4233 487 4247
rect 633 4233 647 4247
rect 673 4233 687 4247
rect 453 4213 467 4227
rect 2033 4233 2047 4247
rect 2233 4233 2247 4247
rect 2553 4233 2567 4247
rect 1234 4213 1248 4227
rect 1733 4213 1747 4227
rect 1792 4213 1806 4227
rect 1833 4213 1847 4227
rect 2113 4213 2127 4227
rect 2314 4213 2328 4227
rect 2634 4213 2648 4227
rect 153 4193 167 4207
rect 293 4193 307 4207
rect 213 4173 227 4187
rect 394 4193 408 4207
rect 632 4193 646 4207
rect 853 4193 867 4207
rect 934 4193 948 4207
rect 1173 4193 1187 4207
rect 1353 4193 1367 4207
rect 134 4153 148 4167
rect 652 4173 666 4187
rect 693 4173 707 4187
rect 733 4173 747 4187
rect 772 4173 786 4187
rect 812 4173 826 4187
rect 933 4173 947 4187
rect 1233 4173 1247 4187
rect 1493 4193 1507 4207
rect 1573 4193 1587 4207
rect 1692 4193 1706 4207
rect 1773 4193 1787 4207
rect 1814 4193 1828 4207
rect 1893 4193 1907 4207
rect 1934 4193 1948 4207
rect 1993 4193 2007 4207
rect 2074 4193 2088 4207
rect 2153 4193 2167 4207
rect 2233 4193 2247 4207
rect 2292 4193 2306 4207
rect 2573 4193 2587 4207
rect 2713 4193 2727 4207
rect 3013 4233 3027 4247
rect 3333 4233 3347 4247
rect 3433 4233 3447 4247
rect 3593 4233 3607 4247
rect 3753 4233 3767 4247
rect 2933 4213 2947 4227
rect 3133 4213 3147 4227
rect 3193 4213 3207 4227
rect 3413 4213 3427 4227
rect 3573 4214 3587 4228
rect 4253 4233 4267 4247
rect 4633 4233 4647 4247
rect 4793 4233 4807 4247
rect 5133 4233 5147 4247
rect 5253 4233 5267 4247
rect 5373 4233 5387 4247
rect 3813 4213 3827 4227
rect 3853 4213 3867 4227
rect 3953 4213 3967 4227
rect 4113 4213 4127 4227
rect 4293 4213 4307 4227
rect 1593 4173 1607 4187
rect 1733 4173 1747 4187
rect 1973 4173 1987 4187
rect 2112 4173 2126 4187
rect 2253 4173 2267 4187
rect 2373 4173 2387 4187
rect 2553 4173 2567 4187
rect 2672 4173 2686 4187
rect 2754 4173 2768 4187
rect 2792 4173 2806 4187
rect 2953 4193 2967 4207
rect 2993 4193 3007 4207
rect 3173 4193 3187 4207
rect 3253 4193 3267 4207
rect 3294 4193 3308 4207
rect 3573 4192 3587 4206
rect 5213 4213 5227 4227
rect 5293 4213 5307 4227
rect 5453 4213 5467 4227
rect 3993 4193 4007 4207
rect 4372 4193 4386 4207
rect 4414 4193 4428 4207
rect 4553 4193 4567 4207
rect 5473 4193 5487 4207
rect 5514 4193 5528 4207
rect 5553 4193 5567 4207
rect 5653 4193 5667 4207
rect 3233 4173 3247 4187
rect 3373 4173 3387 4187
rect 3414 4173 3428 4187
rect 3573 4173 3587 4187
rect 3913 4173 3927 4187
rect 4113 4173 4127 4187
rect 4513 4173 4527 4187
rect 4673 4173 4687 4187
rect 4734 4173 4748 4187
rect 1353 4153 1367 4167
rect 1573 4153 1587 4167
rect 1613 4154 1627 4168
rect 1813 4153 1827 4167
rect 2313 4153 2327 4167
rect 2513 4153 2527 4167
rect 2613 4153 2627 4167
rect 2713 4153 2727 4167
rect 2873 4153 2887 4167
rect 3053 4153 3067 4167
rect 3333 4153 3347 4167
rect 3493 4153 3507 4167
rect 3613 4153 3627 4167
rect 3913 4153 3927 4167
rect 4873 4153 4887 4167
rect 5012 4173 5026 4187
rect 5034 4173 5048 4187
rect 5133 4173 5147 4187
rect 5174 4173 5188 4187
rect 4913 4153 4927 4167
rect 5233 4153 5247 4167
rect 5433 4153 5447 4167
rect 5493 4153 5507 4167
rect 5573 4153 5587 4167
rect 5633 4153 5647 4167
rect 273 4133 287 4147
rect 533 4133 547 4147
rect 633 4133 647 4147
rect 773 4133 787 4147
rect 873 4133 887 4147
rect 1613 4132 1627 4146
rect 1673 4133 1687 4147
rect 2353 4133 2367 4147
rect 2493 4133 2507 4147
rect 2553 4133 2567 4147
rect 3293 4133 3307 4147
rect 3373 4133 3387 4147
rect 3873 4133 3887 4147
rect 4013 4133 4027 4147
rect 4093 4133 4107 4147
rect 4413 4133 4427 4147
rect 5393 4133 5407 4147
rect 5533 4133 5547 4147
rect 573 4113 587 4127
rect 733 4113 747 4127
rect 1173 4113 1187 4127
rect 1513 4113 1527 4127
rect 1773 4113 1787 4127
rect 2133 4113 2147 4127
rect 2233 4113 2247 4127
rect 2473 4113 2487 4127
rect 3813 4113 3827 4127
rect 4193 4114 4207 4128
rect 4333 4113 4347 4127
rect 4393 4113 4407 4127
rect 273 4093 287 4107
rect 593 4093 607 4107
rect 1353 4093 1367 4107
rect 1593 4093 1607 4107
rect 1993 4093 2007 4107
rect 2073 4093 2087 4107
rect 2113 4093 2127 4107
rect 2533 4093 2547 4107
rect 2593 4093 2607 4107
rect 3233 4093 3247 4107
rect 3413 4093 3427 4107
rect 3893 4093 3907 4107
rect 4073 4093 4087 4107
rect 4153 4093 4167 4107
rect 4193 4092 4207 4106
rect 5453 4113 5467 4127
rect 5613 4113 5627 4127
rect 4853 4093 4867 4107
rect 333 4073 347 4087
rect 533 4073 547 4087
rect 2053 4073 2067 4087
rect 2293 4073 2307 4087
rect 2433 4073 2447 4087
rect 2613 4073 2627 4087
rect 2973 4073 2987 4087
rect 3193 4073 3207 4087
rect 3713 4073 3727 4087
rect 4733 4073 4747 4087
rect 5033 4073 5047 4087
rect 113 4053 127 4067
rect 353 4053 367 4067
rect 453 4053 467 4067
rect 693 4053 707 4067
rect 853 4053 867 4067
rect 1313 4053 1327 4067
rect 1973 4053 1987 4067
rect 2093 4053 2107 4067
rect 2653 4053 2667 4067
rect 2793 4053 2807 4067
rect 3333 4053 3347 4067
rect 3413 4053 3427 4067
rect 4533 4053 4547 4067
rect 4753 4053 4767 4067
rect 4913 4053 4927 4067
rect 4973 4053 4987 4067
rect 5153 4053 5167 4067
rect 5632 4053 5646 4067
rect 5654 4053 5668 4067
rect 173 4033 187 4047
rect 333 4033 347 4047
rect 393 4033 407 4047
rect 733 4033 747 4047
rect 1633 4034 1647 4048
rect 113 4013 127 4027
rect 1133 4013 1147 4027
rect 1233 4013 1247 4027
rect 1373 4013 1387 4027
rect 1633 4012 1647 4026
rect 2173 4013 2187 4027
rect 2213 4033 2227 4047
rect 3273 4033 3287 4047
rect 4493 4033 4507 4047
rect 4553 4033 4567 4047
rect 4613 4033 4627 4047
rect 4733 4033 4747 4047
rect 4793 4033 4807 4047
rect 2253 4013 2267 4027
rect 2473 4013 2487 4027
rect 192 3993 206 4007
rect 173 3973 187 3987
rect 313 3973 327 3987
rect 492 3993 506 4007
rect 533 3993 547 4007
rect 593 3993 607 4007
rect 612 3973 626 3987
rect 873 3993 887 4007
rect 1073 3993 1087 4007
rect 1353 3993 1367 4007
rect 1413 3993 1427 4007
rect 1534 3993 1548 4007
rect 1574 3993 1588 4007
rect 53 3953 67 3967
rect 113 3933 127 3947
rect 153 3933 167 3947
rect 373 3953 387 3967
rect 533 3953 547 3967
rect 913 3973 927 3987
rect 693 3953 707 3967
rect 533 3933 547 3947
rect 872 3952 886 3966
rect 993 3933 1007 3947
rect 1113 3973 1127 3987
rect 1154 3973 1168 3987
rect 1273 3953 1287 3967
rect 1413 3953 1427 3967
rect 1473 3973 1487 3987
rect 1552 3973 1566 3987
rect 1873 3993 1887 4007
rect 2093 3993 2107 4007
rect 2413 3993 2427 4007
rect 2113 3973 2127 3987
rect 2533 3993 2547 4007
rect 2793 3993 2807 4007
rect 2993 4013 3007 4027
rect 3053 4013 3067 4027
rect 3373 4013 3387 4027
rect 3573 4013 3587 4027
rect 3673 4013 3687 4027
rect 3833 4013 3847 4027
rect 4493 4013 4507 4027
rect 2973 3993 2987 4007
rect 3213 3993 3227 4007
rect 3693 3993 3707 4007
rect 3893 3993 3907 4007
rect 3972 3993 3986 4007
rect 4173 3993 4187 4007
rect 2573 3973 2587 3987
rect 2733 3973 2747 3987
rect 2873 3973 2887 3987
rect 3092 3973 3106 3987
rect 1533 3953 1547 3967
rect 1593 3953 1607 3967
rect 1774 3953 1788 3967
rect 1913 3953 1927 3967
rect 2213 3953 2227 3967
rect 2293 3953 2307 3967
rect 2652 3953 2666 3967
rect 2674 3953 2688 3967
rect 2813 3953 2827 3967
rect 3013 3953 3027 3967
rect 3073 3953 3087 3967
rect 3173 3953 3187 3967
rect 3254 3953 3268 3967
rect 1033 3933 1047 3947
rect 1653 3933 1667 3947
rect 1793 3933 1807 3947
rect 1913 3933 1927 3947
rect 3472 3973 3486 3987
rect 3513 3973 3527 3987
rect 3613 3973 3627 3987
rect 3553 3953 3567 3967
rect 3753 3953 3767 3967
rect 3893 3954 3907 3968
rect 4013 3973 4027 3987
rect 4053 3973 4067 3987
rect 4853 4013 4867 4027
rect 5373 4013 5387 4027
rect 5513 4013 5527 4027
rect 4713 3993 4727 4007
rect 4813 3993 4827 4007
rect 4874 3993 4888 4007
rect 5132 3993 5146 4007
rect 5193 3993 5207 4007
rect 5413 3993 5427 4007
rect 5653 3993 5667 4007
rect 4833 3973 4847 3987
rect 5373 3973 5387 3987
rect 5414 3973 5428 3987
rect 5593 3973 5607 3987
rect 4293 3953 4307 3967
rect 4453 3953 4467 3967
rect 4513 3953 4527 3967
rect 4614 3953 4628 3967
rect 4673 3953 4687 3967
rect 4933 3953 4947 3967
rect 5012 3953 5026 3967
rect 5133 3953 5147 3967
rect 5233 3953 5247 3967
rect 5673 3953 5687 3967
rect 3573 3933 3587 3947
rect 3893 3932 3907 3946
rect 3953 3933 3967 3947
rect 4473 3933 4487 3947
rect 193 3913 207 3927
rect 273 3913 287 3927
rect 853 3913 867 3927
rect 1993 3913 2007 3927
rect 2113 3913 2127 3927
rect 2473 3913 2487 3927
rect 3053 3913 3067 3927
rect 4233 3913 4247 3927
rect 4513 3913 4527 3927
rect 4833 3913 4847 3927
rect 5253 3913 5267 3927
rect 473 3893 487 3907
rect 913 3893 927 3907
rect 1393 3893 1407 3907
rect 1513 3893 1527 3907
rect 2093 3893 2107 3907
rect 2453 3893 2467 3907
rect 2693 3893 2707 3907
rect 2873 3893 2887 3907
rect 3912 3893 3926 3907
rect 3934 3893 3948 3907
rect 4373 3893 4387 3907
rect 4734 3893 4748 3907
rect 4853 3893 4867 3907
rect 673 3873 687 3887
rect 1113 3873 1127 3887
rect 1273 3873 1287 3887
rect 1333 3873 1347 3887
rect 1453 3873 1467 3887
rect 1773 3873 1787 3887
rect 1813 3873 1827 3887
rect 113 3853 127 3867
rect 3053 3873 3067 3887
rect 3853 3873 3867 3887
rect 3973 3873 3987 3887
rect 4273 3873 4287 3887
rect 4472 3873 4486 3887
rect 4494 3873 4508 3887
rect 5473 3873 5487 3887
rect 2233 3853 2247 3867
rect 3033 3853 3047 3867
rect 3193 3853 3207 3867
rect 3373 3853 3387 3867
rect 3453 3853 3467 3867
rect 3553 3853 3567 3867
rect 3613 3853 3627 3867
rect 3753 3853 3767 3867
rect 3993 3853 4007 3867
rect 4093 3853 4107 3867
rect 5093 3853 5107 3867
rect 5293 3853 5307 3867
rect 1593 3833 1607 3847
rect 1633 3833 1647 3847
rect 1733 3833 1747 3847
rect 1953 3833 1967 3847
rect 2153 3833 2167 3847
rect 2533 3833 2547 3847
rect 2573 3833 2587 3847
rect 2933 3833 2947 3847
rect 3113 3833 3127 3847
rect 3253 3833 3267 3847
rect 3573 3833 3587 3847
rect 3813 3833 3827 3847
rect 4133 3833 4147 3847
rect 4513 3833 4527 3847
rect 4613 3833 4627 3847
rect 4973 3833 4987 3847
rect 5193 3833 5207 3847
rect 5433 3833 5447 3847
rect 193 3813 207 3827
rect 473 3813 487 3827
rect 1553 3813 1567 3827
rect 1753 3813 1767 3827
rect 2014 3813 2028 3827
rect 2733 3813 2747 3827
rect 3133 3813 3147 3827
rect 3753 3813 3767 3827
rect 4093 3813 4107 3827
rect 4713 3813 4727 3827
rect 4813 3813 4827 3827
rect 5213 3813 5227 3827
rect 5253 3813 5267 3827
rect 5313 3813 5327 3827
rect 233 3793 247 3807
rect 353 3793 367 3807
rect 973 3793 987 3807
rect 1253 3793 1267 3807
rect 1653 3793 1667 3807
rect 2433 3793 2447 3807
rect 2513 3793 2527 3807
rect 3073 3793 3087 3807
rect 3113 3793 3127 3807
rect 4133 3793 4147 3807
rect 533 3773 547 3787
rect 853 3773 867 3787
rect 1033 3773 1047 3787
rect 1153 3773 1167 3787
rect 1593 3773 1607 3787
rect 1853 3773 1867 3787
rect 1973 3773 1987 3787
rect 2094 3773 2108 3787
rect 2653 3773 2667 3787
rect 2853 3773 2867 3787
rect 3013 3773 3027 3787
rect 3053 3773 3067 3787
rect 3093 3773 3107 3787
rect 3253 3773 3267 3787
rect 3413 3773 3427 3787
rect 3653 3773 3667 3787
rect 5093 3773 5107 3787
rect 5193 3773 5207 3787
rect 993 3753 1007 3767
rect 1053 3753 1067 3767
rect 1333 3753 1347 3767
rect 1733 3753 1747 3767
rect 1773 3753 1787 3767
rect 2013 3753 2027 3767
rect 2953 3753 2967 3767
rect 3353 3753 3367 3767
rect 3553 3753 3567 3767
rect 233 3733 247 3747
rect 473 3733 487 3747
rect 813 3733 827 3747
rect 853 3733 867 3747
rect 973 3733 987 3747
rect 13 3713 27 3727
rect 153 3713 167 3727
rect 273 3713 287 3727
rect 354 3713 368 3727
rect 872 3713 886 3727
rect 972 3713 986 3727
rect 1012 3714 1026 3728
rect 1153 3733 1167 3747
rect 1193 3733 1207 3747
rect 1513 3733 1527 3747
rect 1653 3733 1667 3747
rect 1893 3733 1907 3747
rect 2052 3733 2066 3747
rect 2113 3733 2127 3747
rect 2193 3733 2207 3747
rect 2253 3733 2267 3747
rect 2353 3733 2367 3747
rect 2393 3733 2407 3747
rect 2513 3733 2527 3747
rect 2613 3733 2627 3747
rect 2713 3734 2727 3748
rect 2893 3733 2907 3747
rect 1193 3713 1207 3727
rect 133 3693 147 3707
rect 173 3693 187 3707
rect 314 3693 328 3707
rect 372 3693 386 3707
rect 493 3692 507 3706
rect 573 3693 587 3707
rect 1073 3693 1087 3707
rect 1573 3713 1587 3727
rect 1773 3713 1787 3727
rect 2033 3713 2047 3727
rect 2413 3713 2427 3727
rect 1293 3693 1307 3707
rect 1453 3693 1467 3707
rect 513 3673 527 3687
rect 733 3673 747 3687
rect 992 3673 1006 3687
rect 1014 3673 1028 3687
rect 1652 3693 1666 3707
rect 1753 3693 1767 3707
rect 1893 3693 1907 3707
rect 1973 3693 1987 3707
rect 2113 3693 2127 3707
rect 2193 3693 2207 3707
rect 2233 3693 2247 3707
rect 2353 3693 2367 3707
rect 2713 3712 2727 3726
rect 2653 3693 2667 3707
rect 2812 3713 2826 3727
rect 2853 3713 2867 3727
rect 2953 3713 2967 3727
rect 2753 3693 2767 3707
rect 3052 3713 3066 3727
rect 1593 3673 1607 3687
rect 1773 3673 1787 3687
rect 1813 3673 1827 3687
rect 373 3653 387 3667
rect 733 3653 747 3667
rect 873 3653 887 3667
rect 1293 3653 1307 3667
rect 1853 3653 1867 3667
rect 2033 3673 2047 3687
rect 2193 3673 2207 3687
rect 2393 3673 2407 3687
rect 2473 3673 2487 3687
rect 2593 3673 2607 3687
rect 2713 3673 2727 3687
rect 2993 3693 3007 3707
rect 3133 3733 3147 3747
rect 3353 3733 3367 3747
rect 3413 3733 3427 3747
rect 3613 3734 3627 3748
rect 3793 3753 3807 3767
rect 4973 3753 4987 3767
rect 5593 3753 5607 3767
rect 5713 3753 5727 3767
rect 3733 3733 3747 3747
rect 3933 3733 3947 3747
rect 4173 3733 4187 3747
rect 5093 3733 5107 3747
rect 3613 3712 3627 3726
rect 3653 3713 3667 3727
rect 3753 3713 3767 3727
rect 3793 3713 3807 3727
rect 3852 3713 3866 3727
rect 3993 3713 4007 3727
rect 4113 3713 4127 3727
rect 4573 3713 4587 3727
rect 4973 3714 4987 3728
rect 5213 3713 5227 3727
rect 5693 3713 5707 3727
rect 3074 3693 3088 3707
rect 3133 3693 3147 3707
rect 3194 3693 3208 3707
rect 3413 3693 3427 3707
rect 3713 3693 3727 3707
rect 3913 3693 3927 3707
rect 4053 3693 4067 3707
rect 2913 3673 2927 3687
rect 3093 3673 3107 3687
rect 3273 3673 3287 3687
rect 3553 3673 3567 3687
rect 4213 3693 4227 3707
rect 4293 3693 4307 3707
rect 4453 3693 4467 3707
rect 4533 3693 4547 3707
rect 4693 3693 4707 3707
rect 4773 3693 4787 3707
rect 4814 3693 4828 3707
rect 4953 3693 4967 3707
rect 4994 3693 5008 3707
rect 5293 3693 5307 3707
rect 5373 3693 5387 3707
rect 5414 3693 5428 3707
rect 2053 3653 2067 3667
rect 2233 3653 2247 3667
rect 2373 3653 2387 3667
rect 313 3633 327 3647
rect 533 3633 547 3647
rect 493 3613 507 3627
rect 1393 3633 1407 3647
rect 1913 3633 1927 3647
rect 2093 3633 2107 3647
rect 2733 3653 2747 3667
rect 2813 3653 2827 3667
rect 3073 3653 3087 3667
rect 3473 3653 3487 3667
rect 3853 3653 3867 3667
rect 4033 3653 4047 3667
rect 4153 3673 4167 3687
rect 4353 3673 4367 3687
rect 4893 3673 4907 3687
rect 5093 3673 5107 3687
rect 5493 3673 5507 3687
rect 5673 3673 5687 3687
rect 4193 3653 4207 3667
rect 5033 3653 5047 3667
rect 5113 3653 5127 3667
rect 5233 3653 5247 3667
rect 2613 3633 2627 3647
rect 2933 3633 2947 3647
rect 1293 3613 1307 3627
rect 1353 3613 1367 3627
rect 1433 3613 1447 3627
rect 1473 3613 1487 3627
rect 2333 3613 2347 3627
rect 3213 3613 3227 3627
rect 3813 3633 3827 3647
rect 4133 3633 4147 3647
rect 4773 3633 4787 3647
rect 4833 3633 4847 3647
rect 4913 3633 4927 3647
rect 3833 3613 3847 3627
rect 4153 3613 4167 3627
rect 4353 3613 4367 3627
rect 4433 3613 4447 3627
rect 4713 3613 4727 3627
rect 4753 3613 4767 3627
rect 4793 3613 4807 3627
rect 4933 3613 4947 3627
rect 5373 3613 5387 3627
rect 1373 3593 1387 3607
rect 1453 3593 1467 3607
rect 1553 3593 1567 3607
rect 73 3573 87 3587
rect 233 3573 247 3587
rect 1413 3573 1427 3587
rect 1733 3573 1747 3587
rect 1833 3593 1847 3607
rect 2553 3593 2567 3607
rect 3053 3593 3067 3607
rect 3193 3593 3207 3607
rect 3353 3593 3367 3607
rect 3733 3593 3747 3607
rect 3913 3593 3927 3607
rect 4473 3593 4487 3607
rect 4813 3593 4827 3607
rect 4993 3593 5007 3607
rect 5053 3593 5067 3607
rect 5213 3593 5227 3607
rect 2013 3573 2027 3587
rect 2413 3573 2427 3587
rect 2773 3573 2787 3587
rect 2853 3573 2867 3587
rect 2913 3573 2927 3587
rect 3613 3573 3627 3587
rect 3753 3573 3767 3587
rect 4173 3573 4187 3587
rect 4313 3573 4327 3587
rect 4553 3573 4567 3587
rect 5073 3573 5087 3587
rect 713 3553 727 3567
rect 793 3553 807 3567
rect 1293 3553 1307 3567
rect 1553 3553 1567 3567
rect 1613 3553 1627 3567
rect 1813 3553 1827 3567
rect 2493 3553 2507 3567
rect 3113 3553 3127 3567
rect 173 3533 187 3547
rect 493 3533 507 3547
rect 1173 3533 1187 3547
rect 1733 3533 1747 3547
rect 1873 3533 1887 3547
rect 1973 3533 1987 3547
rect 2014 3533 2028 3547
rect 53 3513 67 3527
rect 94 3513 108 3527
rect 134 3513 148 3527
rect 193 3513 207 3527
rect 112 3493 126 3507
rect 233 3513 247 3527
rect 333 3513 347 3527
rect 632 3513 646 3527
rect 673 3513 687 3527
rect 753 3513 767 3527
rect 793 3513 807 3527
rect 933 3513 947 3527
rect 1253 3513 1267 3527
rect 1373 3513 1387 3527
rect 1533 3513 1547 3527
rect 1574 3513 1588 3527
rect 1773 3513 1787 3527
rect 2113 3513 2127 3527
rect 2253 3533 2267 3547
rect 2333 3533 2347 3547
rect 2273 3513 2287 3527
rect 2353 3514 2367 3528
rect 2653 3533 2667 3547
rect 2933 3534 2947 3548
rect 3253 3553 3267 3567
rect 3833 3553 3847 3567
rect 4433 3553 4447 3567
rect 5713 3553 5727 3567
rect 3233 3533 3247 3547
rect 3273 3533 3287 3547
rect 3413 3533 3427 3547
rect 3493 3533 3507 3547
rect 3633 3533 3647 3547
rect 4113 3533 4127 3547
rect 4273 3533 4287 3547
rect 4733 3533 4747 3547
rect 4933 3533 4947 3547
rect 5053 3533 5067 3547
rect 2613 3513 2627 3527
rect 2714 3513 2728 3527
rect 2912 3513 2926 3527
rect 1233 3493 1247 3507
rect 1353 3493 1367 3507
rect 1453 3493 1467 3507
rect 1613 3493 1627 3507
rect 1653 3493 1667 3507
rect 2073 3493 2087 3507
rect 2934 3512 2948 3526
rect 3192 3513 3206 3527
rect 3234 3513 3248 3527
rect 3353 3513 3367 3527
rect 4012 3513 4026 3527
rect 2353 3493 2367 3506
rect 2433 3493 2447 3507
rect 2673 3493 2687 3507
rect 2813 3493 2827 3507
rect 2893 3493 2907 3507
rect 3032 3493 3046 3507
rect 3113 3493 3127 3507
rect 4253 3513 4267 3527
rect 3594 3493 3608 3507
rect 3713 3493 3727 3507
rect 3754 3493 3768 3507
rect 3833 3493 3847 3507
rect 4034 3493 4048 3507
rect 4173 3493 4187 3507
rect 4313 3513 4327 3527
rect 4533 3513 4547 3527
rect 4793 3513 4807 3527
rect 4893 3513 4907 3527
rect 5233 3533 5247 3547
rect 5513 3533 5527 3547
rect 5193 3513 5207 3527
rect 5254 3513 5268 3527
rect 4593 3493 4607 3507
rect 5033 3493 5047 3507
rect 5233 3493 5247 3507
rect 192 3473 206 3487
rect 332 3473 346 3487
rect 374 3473 388 3487
rect 713 3473 727 3487
rect 93 3453 107 3467
rect 493 3453 507 3467
rect 773 3453 787 3467
rect 893 3473 907 3487
rect 1273 3473 1287 3487
rect 1432 3473 1446 3487
rect 1173 3453 1187 3467
rect 2353 3492 2367 3493
rect 1853 3473 1867 3487
rect 1933 3473 1947 3487
rect 2113 3473 2127 3487
rect 2213 3473 2227 3487
rect 2253 3473 2267 3487
rect 2413 3473 2427 3487
rect 3093 3473 3107 3487
rect 3493 3473 3507 3487
rect 3873 3474 3887 3488
rect 4153 3473 4167 3487
rect 4453 3473 4467 3487
rect 4713 3473 4727 3487
rect 5253 3473 5267 3487
rect 5373 3473 5387 3487
rect 5473 3473 5487 3487
rect 5593 3473 5607 3487
rect 2153 3453 2167 3467
rect 293 3433 307 3447
rect 373 3433 387 3447
rect 753 3433 767 3447
rect 893 3433 907 3447
rect 1353 3433 1367 3447
rect 1512 3433 1526 3447
rect 1573 3433 1587 3447
rect 1893 3433 1907 3447
rect 1993 3433 2007 3447
rect 2033 3433 2047 3447
rect 2253 3433 2267 3447
rect 2293 3433 2307 3447
rect 2493 3453 2507 3467
rect 2593 3453 2607 3467
rect 3673 3453 3687 3467
rect 3873 3452 3887 3466
rect 4253 3453 4267 3467
rect 4613 3453 4627 3467
rect 5533 3453 5547 3467
rect 2833 3433 2847 3447
rect 3433 3433 3447 3447
rect 3893 3433 3907 3447
rect 3953 3433 3967 3447
rect 4473 3434 4487 3448
rect 4573 3433 4587 3447
rect 5073 3433 5087 3447
rect 1693 3413 1707 3427
rect 2234 3413 2248 3427
rect 3153 3413 3167 3427
rect 3233 3413 3247 3427
rect 3533 3413 3547 3427
rect 3573 3413 3587 3427
rect 3772 3413 3786 3427
rect 3794 3413 3808 3427
rect 4413 3413 4427 3427
rect 4473 3412 4487 3426
rect 193 3393 207 3407
rect 1013 3393 1027 3407
rect 1473 3393 1487 3407
rect 2293 3393 2307 3407
rect 3073 3393 3087 3407
rect 3673 3393 3687 3407
rect 3893 3393 3907 3407
rect 4033 3393 4047 3407
rect 4133 3393 4147 3407
rect 4733 3393 4747 3407
rect 5553 3413 5567 3427
rect 5633 3413 5647 3427
rect 4973 3393 4987 3407
rect 5293 3393 5307 3407
rect 5613 3393 5627 3407
rect 1433 3373 1447 3387
rect 1853 3373 1867 3387
rect 1973 3373 1987 3387
rect 2253 3373 2267 3387
rect 2513 3373 2527 3387
rect 2713 3373 2727 3387
rect 3413 3373 3427 3387
rect 3993 3373 4007 3387
rect 113 3353 127 3367
rect 773 3353 787 3367
rect 833 3353 847 3367
rect 913 3353 927 3367
rect 1153 3353 1167 3367
rect 1873 3353 1887 3367
rect 1993 3353 2007 3367
rect 2973 3353 2987 3367
rect 3153 3353 3167 3367
rect 3373 3354 3387 3368
rect 3853 3353 3867 3367
rect 4113 3373 4127 3387
rect 4573 3373 4587 3387
rect 5033 3373 5047 3387
rect 5193 3373 5207 3387
rect 1333 3333 1347 3347
rect 1553 3333 1567 3347
rect 1733 3333 1747 3347
rect 2113 3333 2127 3347
rect 2293 3333 2307 3347
rect 2713 3333 2727 3347
rect 2933 3333 2947 3347
rect 473 3293 487 3307
rect 533 3293 547 3307
rect 713 3313 727 3327
rect 853 3313 867 3327
rect 1133 3293 1147 3307
rect 1473 3293 1487 3307
rect 1613 3293 1627 3307
rect 73 3273 87 3287
rect 233 3273 247 3287
rect 332 3253 346 3267
rect 493 3273 507 3287
rect 533 3273 547 3287
rect 1013 3273 1027 3287
rect 1313 3273 1327 3287
rect 893 3253 907 3267
rect 53 3233 67 3247
rect 192 3233 206 3247
rect 232 3233 246 3247
rect 293 3233 307 3247
rect 513 3233 527 3247
rect 574 3233 588 3247
rect 634 3233 648 3247
rect 853 3233 867 3247
rect 1013 3253 1027 3267
rect 1132 3253 1146 3267
rect 1173 3254 1187 3268
rect 1393 3253 1407 3267
rect 1733 3293 1747 3307
rect 1973 3313 1987 3327
rect 2453 3313 2467 3327
rect 3373 3332 3387 3346
rect 3453 3333 3467 3347
rect 3713 3333 3727 3347
rect 4233 3353 4247 3367
rect 4373 3353 4387 3367
rect 4613 3353 4627 3367
rect 4753 3353 4767 3367
rect 4873 3353 4887 3367
rect 4933 3353 4947 3367
rect 5533 3353 5547 3367
rect 4073 3333 4087 3347
rect 5153 3333 5167 3347
rect 5593 3333 5607 3347
rect 2813 3313 2827 3327
rect 4033 3313 4047 3327
rect 4392 3313 4406 3327
rect 4414 3313 4428 3327
rect 2193 3293 2207 3307
rect 2433 3293 2447 3307
rect 2733 3293 2747 3307
rect 2833 3293 2847 3307
rect 3173 3293 3187 3307
rect 3533 3293 3547 3307
rect 4093 3293 4107 3307
rect 4253 3293 4267 3307
rect 4333 3293 4347 3307
rect 4373 3293 4387 3307
rect 4533 3293 4547 3307
rect 4593 3313 4607 3327
rect 4933 3313 4947 3327
rect 5213 3313 5227 3327
rect 5253 3313 5267 3327
rect 4632 3293 4646 3307
rect 4733 3293 4747 3307
rect 4813 3293 4827 3307
rect 4853 3293 4867 3307
rect 5233 3293 5247 3307
rect 5573 3293 5587 3307
rect 1692 3273 1706 3287
rect 1714 3273 1728 3287
rect 1793 3273 1807 3287
rect 2193 3273 2207 3287
rect 2793 3273 2807 3287
rect 2993 3273 3007 3287
rect 3033 3273 3047 3287
rect 3573 3273 3587 3287
rect 4293 3273 4307 3287
rect 4793 3273 4807 3287
rect 4973 3273 4987 3287
rect 5093 3273 5107 3287
rect 1733 3253 1747 3267
rect 1773 3253 1787 3267
rect 1893 3253 1907 3267
rect 1953 3253 1967 3267
rect 2073 3253 2087 3267
rect 2113 3253 2127 3267
rect 2253 3253 2267 3267
rect 2292 3253 2306 3267
rect 2713 3253 2727 3267
rect 3053 3253 3067 3267
rect 3093 3253 3107 3267
rect 3233 3253 3247 3267
rect 3533 3253 3547 3267
rect 4093 3253 4107 3267
rect 4173 3253 4187 3267
rect 4473 3253 4487 3267
rect 4533 3253 4547 3267
rect 4753 3253 4767 3267
rect 4973 3253 4987 3267
rect 5153 3253 5167 3267
rect 5293 3253 5307 3267
rect 1093 3233 1107 3247
rect 1193 3233 1207 3247
rect 1273 3233 1287 3247
rect 112 3213 126 3227
rect 373 3213 387 3227
rect 1933 3233 1947 3247
rect 2333 3233 2347 3247
rect 2573 3233 2587 3247
rect 2653 3233 2667 3247
rect 612 3213 626 3227
rect 833 3213 847 3227
rect 1054 3213 1068 3227
rect 473 3193 487 3207
rect 853 3193 867 3207
rect 893 3193 907 3207
rect 1572 3213 1586 3227
rect 1653 3213 1667 3227
rect 1973 3213 1987 3227
rect 2173 3213 2187 3227
rect 2993 3233 3007 3247
rect 2413 3213 2427 3227
rect 2793 3213 2807 3227
rect 3133 3213 3147 3227
rect 3253 3233 3267 3247
rect 3413 3233 3427 3247
rect 3473 3233 3487 3247
rect 1293 3193 1307 3207
rect 1353 3193 1367 3207
rect 2153 3193 2167 3207
rect 2373 3193 2387 3207
rect 3433 3213 3447 3227
rect 2653 3193 2667 3207
rect 2733 3193 2747 3207
rect 2773 3193 2787 3207
rect 2893 3193 2907 3207
rect 3453 3193 3467 3207
rect 3573 3213 3587 3227
rect 3692 3213 3706 3227
rect 3714 3213 3728 3227
rect 3773 3213 3787 3227
rect 3893 3213 3907 3227
rect 3953 3213 3967 3227
rect 4254 3233 4268 3247
rect 4393 3233 4407 3247
rect 4553 3233 4567 3247
rect 4633 3233 4647 3247
rect 4733 3233 4747 3247
rect 4793 3233 4807 3247
rect 4933 3233 4947 3247
rect 5073 3233 5087 3247
rect 5333 3233 5347 3247
rect 5433 3253 5447 3267
rect 5513 3253 5527 3267
rect 4233 3213 4247 3227
rect 4313 3213 4327 3227
rect 4773 3213 4787 3227
rect 5053 3213 5067 3227
rect 5193 3213 5207 3227
rect 5293 3213 5307 3227
rect 5473 3233 5487 3247
rect 4373 3193 4387 3207
rect 4533 3193 4547 3207
rect 4653 3193 4667 3207
rect 5592 3213 5606 3227
rect 5073 3193 5087 3207
rect 5153 3193 5167 3207
rect 5353 3193 5367 3207
rect 5413 3193 5427 3207
rect 5533 3193 5547 3207
rect 1113 3173 1127 3187
rect 1273 3173 1287 3187
rect 1833 3173 1847 3187
rect 2353 3173 2367 3187
rect 2413 3173 2427 3187
rect 2793 3173 2807 3187
rect 3233 3173 3247 3187
rect 3373 3173 3387 3187
rect 3413 3173 3427 3187
rect 4313 3173 4327 3187
rect 4433 3173 4447 3187
rect 4513 3173 4527 3187
rect 4793 3173 4807 3187
rect 5113 3173 5127 3187
rect 1093 3153 1107 3167
rect 1193 3153 1207 3167
rect 193 3133 207 3147
rect 1393 3133 1407 3147
rect 1913 3153 1927 3167
rect 2133 3153 2147 3167
rect 2333 3153 2347 3167
rect 2373 3153 2387 3167
rect 2853 3153 2867 3167
rect 3233 3153 3247 3167
rect 4293 3153 4307 3167
rect 4493 3153 4507 3167
rect 4853 3153 4867 3167
rect 5133 3153 5147 3167
rect 5393 3153 5407 3167
rect 5513 3153 5527 3167
rect 5613 3153 5627 3167
rect 2113 3133 2127 3147
rect 2313 3133 2327 3147
rect 2513 3134 2527 3148
rect 2573 3133 2587 3147
rect 2893 3133 2907 3147
rect 2953 3133 2967 3147
rect 3153 3133 3167 3147
rect 3513 3133 3527 3147
rect 3833 3133 3847 3147
rect 4413 3133 4427 3147
rect 693 3113 707 3127
rect 773 3113 787 3127
rect 933 3113 947 3127
rect 1053 3113 1067 3127
rect 1173 3113 1187 3127
rect 1293 3113 1307 3127
rect 1753 3113 1767 3127
rect 2093 3113 2107 3127
rect 2173 3113 2187 3127
rect 2413 3113 2427 3127
rect 2453 3113 2467 3127
rect 153 3093 167 3107
rect 1853 3093 1867 3107
rect 1992 3093 2006 3107
rect 2014 3093 2028 3107
rect 2053 3093 2067 3107
rect 2473 3093 2487 3107
rect 2513 3112 2527 3126
rect 3233 3113 3247 3127
rect 3373 3113 3387 3127
rect 3672 3113 3686 3127
rect 3694 3113 3708 3127
rect 4073 3113 4087 3127
rect 4733 3133 4747 3147
rect 4993 3133 5007 3147
rect 5053 3133 5067 3147
rect 5153 3133 5167 3147
rect 5473 3133 5487 3147
rect 5553 3133 5567 3147
rect 5013 3113 5027 3127
rect 293 3073 307 3087
rect 353 3073 367 3087
rect 613 3073 627 3087
rect 1313 3073 1327 3087
rect 1453 3073 1467 3087
rect 2113 3073 2127 3087
rect 2233 3073 2247 3087
rect 2353 3073 2367 3087
rect 2433 3073 2447 3087
rect 2593 3073 2607 3087
rect 2653 3093 2667 3107
rect 2733 3093 2747 3107
rect 2913 3093 2927 3107
rect 3473 3093 3487 3107
rect 3653 3093 3667 3107
rect 4433 3093 4447 3107
rect 4533 3093 4547 3107
rect 393 3053 407 3067
rect 533 3053 547 3067
rect 673 3053 687 3067
rect 993 3053 1007 3067
rect 1034 3053 1048 3067
rect 2114 3053 2128 3067
rect 153 3033 167 3047
rect 393 3033 407 3047
rect 433 3033 447 3047
rect 493 3033 507 3047
rect 534 3033 548 3047
rect 773 3033 787 3047
rect 894 3033 908 3047
rect 973 3033 987 3047
rect 1113 3033 1127 3047
rect 233 3013 247 3027
rect 333 3013 347 3027
rect 473 3013 487 3027
rect 613 3013 627 3027
rect 673 3013 687 3027
rect 833 3013 847 3027
rect 874 3013 888 3027
rect 1373 3033 1387 3047
rect 1573 3033 1587 3047
rect 1773 3033 1787 3047
rect 1833 3033 1847 3047
rect 1873 3033 1887 3047
rect 2052 3033 2066 3047
rect 2092 3034 2106 3048
rect 2693 3053 2707 3067
rect 2773 3073 2787 3087
rect 3373 3073 3387 3087
rect 3493 3073 3507 3087
rect 3793 3073 3807 3087
rect 4232 3073 4246 3087
rect 4254 3073 4268 3087
rect 4373 3073 4387 3087
rect 4513 3073 4527 3087
rect 4592 3073 4606 3087
rect 4614 3073 4628 3087
rect 4713 3073 4727 3087
rect 4873 3093 4887 3107
rect 5113 3093 5127 3107
rect 5253 3093 5267 3107
rect 5453 3113 5467 3127
rect 5613 3113 5627 3127
rect 5593 3093 5607 3107
rect 4913 3073 4927 3087
rect 2753 3053 2767 3067
rect 2893 3053 2907 3067
rect 3092 3053 3106 3067
rect 3114 3053 3128 3067
rect 3293 3053 3307 3067
rect 3913 3053 3927 3067
rect 2193 3033 2207 3047
rect 2293 3033 2307 3047
rect 2352 3033 2366 3047
rect 2393 3033 2407 3047
rect 2634 3033 2648 3047
rect 2833 3033 2847 3047
rect 1033 3013 1047 3027
rect 173 2993 187 3007
rect 294 2993 308 3007
rect 973 2993 987 3007
rect 1213 3013 1227 3027
rect 1353 3013 1367 3027
rect 1473 3013 1487 3027
rect 1514 3013 1528 3027
rect 1753 3013 1767 3027
rect 1893 3013 1907 3027
rect 1973 3013 1987 3027
rect 2074 3013 2088 3027
rect 2133 3013 2147 3027
rect 2473 3013 2487 3027
rect 2533 3013 2547 3027
rect 2573 3013 2587 3027
rect 2653 3013 2667 3027
rect 2693 3013 2707 3027
rect 2993 3013 3007 3027
rect 3132 3013 3146 3027
rect 3173 3013 3187 3027
rect 3252 3033 3266 3047
rect 3294 3033 3308 3047
rect 3333 3033 3347 3047
rect 3552 3033 3566 3047
rect 3593 3033 3607 3047
rect 3773 3033 3787 3047
rect 3893 3033 3907 3047
rect 4353 3053 4367 3067
rect 4573 3047 4587 3048
rect 3373 3013 3387 3027
rect 3453 3013 3467 3027
rect 3733 3013 3747 3027
rect 4093 3033 4107 3047
rect 4033 3013 4047 3027
rect 4433 3033 4447 3047
rect 4573 3034 4587 3047
rect 4773 3053 4787 3067
rect 5193 3053 5207 3067
rect 5292 3053 5306 3067
rect 5314 3053 5328 3067
rect 5353 3053 5367 3067
rect 5473 3053 5487 3067
rect 5533 3053 5547 3067
rect 4253 3013 4267 3027
rect 4312 3013 4326 3027
rect 4413 3013 4427 3027
rect 1073 2993 1087 3007
rect 1253 2993 1267 3007
rect 1453 2993 1467 3007
rect 2293 2993 2307 3007
rect 2633 2993 2647 3007
rect 3413 2993 3427 3007
rect 3552 2993 3566 3007
rect 3574 2993 3588 3007
rect 3653 2993 3667 3007
rect 3713 2993 3727 3007
rect 4013 2993 4027 3007
rect 4093 2993 4107 3007
rect 4173 2993 4187 3007
rect 4233 2993 4247 3007
rect 4492 2993 4506 3007
rect 4573 3012 4587 3026
rect 5334 3033 5348 3047
rect 5593 3033 5607 3047
rect 4693 3013 4707 3027
rect 4774 3012 4788 3026
rect 4872 3013 4886 3027
rect 4974 3013 4988 3027
rect 5113 3013 5127 3027
rect 5193 3013 5207 3027
rect 5273 3013 5287 3027
rect 5354 3013 5368 3027
rect 5433 3013 5447 3027
rect 4752 2993 4766 3007
rect 4852 2993 4866 3007
rect 4933 2993 4947 3007
rect 5073 2993 5087 3007
rect 5133 2993 5147 3007
rect 5313 2993 5327 3007
rect 5513 3013 5527 3027
rect 5473 2993 5487 3007
rect 493 2973 507 2987
rect 653 2973 667 2987
rect 873 2973 887 2987
rect 1353 2973 1367 2987
rect 1553 2973 1567 2987
rect 1873 2973 1887 2987
rect 2393 2973 2407 2987
rect 2493 2973 2507 2987
rect 2833 2973 2847 2987
rect 3113 2973 3127 2987
rect 3233 2973 3247 2987
rect 3614 2973 3628 2987
rect 3733 2973 3747 2987
rect 3973 2973 3987 2987
rect 4033 2973 4047 2987
rect 4252 2973 4266 2987
rect 4433 2973 4447 2987
rect 4773 2973 4787 2987
rect 4973 2973 4987 2987
rect 5092 2973 5106 2987
rect 5114 2973 5128 2987
rect 5153 2974 5167 2988
rect 5273 2973 5287 2987
rect 73 2953 87 2967
rect 273 2953 287 2967
rect 373 2953 387 2967
rect 613 2953 627 2967
rect 833 2953 847 2967
rect 1353 2953 1367 2967
rect 1793 2953 1807 2967
rect 2033 2953 2047 2967
rect 2553 2953 2567 2967
rect 2813 2953 2827 2967
rect 2973 2953 2987 2967
rect 3053 2953 3067 2967
rect 3393 2953 3407 2967
rect 3673 2953 3687 2967
rect 4093 2953 4107 2967
rect 4173 2953 4187 2967
rect 4653 2953 4667 2967
rect 4753 2954 4767 2968
rect 5153 2952 5167 2966
rect 5233 2953 5247 2967
rect 5553 2953 5567 2967
rect 253 2933 267 2947
rect 573 2933 587 2947
rect 1253 2933 1267 2947
rect 1473 2933 1487 2947
rect 1813 2933 1827 2947
rect 2093 2933 2107 2947
rect 2233 2933 2247 2947
rect 2293 2933 2307 2947
rect 2653 2933 2667 2947
rect 2993 2933 3007 2947
rect 3373 2933 3387 2947
rect 3533 2933 3547 2947
rect 4074 2933 4088 2947
rect 4113 2934 4127 2948
rect 4473 2933 4487 2947
rect 4553 2933 4567 2947
rect 4753 2932 4767 2946
rect 4913 2934 4927 2948
rect 4973 2933 4987 2947
rect 5293 2933 5307 2947
rect 5533 2933 5547 2947
rect 193 2913 207 2927
rect 473 2913 487 2927
rect 993 2913 1007 2927
rect 2313 2913 2327 2927
rect 3853 2913 3867 2927
rect 4013 2913 4027 2927
rect 4113 2912 4127 2926
rect 4294 2913 4308 2927
rect 4352 2913 4366 2927
rect 4374 2913 4388 2927
rect 4913 2912 4927 2926
rect 4953 2913 4967 2927
rect 4993 2913 5007 2927
rect 5593 2913 5607 2927
rect 5633 2913 5647 2927
rect 13 2893 27 2907
rect 73 2893 87 2907
rect 493 2893 507 2907
rect 593 2893 607 2907
rect 1653 2893 1667 2907
rect 1933 2873 1947 2887
rect 2313 2873 2327 2887
rect 2613 2893 2627 2907
rect 2953 2893 2967 2907
rect 3033 2893 3047 2907
rect 3453 2893 3467 2907
rect 3913 2893 3927 2907
rect 4253 2893 4267 2907
rect 4313 2893 4327 2907
rect 4473 2893 4487 2907
rect 4513 2893 4527 2907
rect 4793 2893 4807 2907
rect 4873 2893 4887 2907
rect 5213 2893 5227 2907
rect 2713 2873 2727 2887
rect 3013 2873 3027 2887
rect 3113 2873 3127 2887
rect 3713 2873 3727 2887
rect 3773 2873 3787 2887
rect 3853 2873 3867 2887
rect 833 2853 847 2867
rect 932 2853 946 2867
rect 954 2853 968 2867
rect 993 2853 1007 2867
rect 1073 2853 1087 2867
rect 1133 2853 1147 2867
rect 1693 2853 1707 2867
rect 2133 2853 2147 2867
rect 2173 2853 2187 2867
rect 2353 2853 2367 2867
rect 3093 2853 3107 2867
rect 3312 2853 3326 2867
rect 3334 2853 3348 2867
rect 3453 2853 3467 2867
rect 4132 2873 4146 2887
rect 4154 2873 4168 2887
rect 4373 2873 4387 2887
rect 4413 2873 4427 2887
rect 4993 2873 5007 2887
rect 5073 2873 5087 2887
rect 5393 2893 5407 2907
rect 5253 2873 5267 2887
rect 5353 2873 5367 2887
rect 133 2833 147 2847
rect 213 2834 227 2848
rect 873 2833 887 2847
rect 913 2833 927 2847
rect 1273 2833 1287 2847
rect 1973 2833 1987 2847
rect 2153 2833 2167 2847
rect 53 2813 67 2827
rect 173 2813 187 2827
rect 213 2812 227 2826
rect 533 2813 547 2827
rect 793 2813 807 2827
rect 213 2793 227 2807
rect 293 2793 307 2807
rect 373 2793 387 2807
rect 493 2793 507 2807
rect 1053 2813 1067 2827
rect 1733 2813 1747 2827
rect 1913 2813 1927 2827
rect 2092 2813 2106 2827
rect 2273 2833 2287 2847
rect 2473 2833 2487 2847
rect 2513 2833 2527 2847
rect 2673 2833 2687 2847
rect 2913 2833 2927 2847
rect 3433 2833 3447 2847
rect 3733 2833 3747 2847
rect 3773 2833 3787 2847
rect 4653 2853 4667 2867
rect 4733 2853 4747 2867
rect 4933 2853 4947 2867
rect 5133 2853 5147 2867
rect 5173 2853 5187 2867
rect 4093 2833 4107 2847
rect 4913 2833 4927 2847
rect 5213 2833 5227 2847
rect 2253 2813 2267 2827
rect 2573 2813 2587 2827
rect 3573 2813 3587 2827
rect 3653 2813 3667 2827
rect 3713 2813 3727 2827
rect 3813 2813 3827 2827
rect 4013 2813 4027 2827
rect 493 2773 507 2787
rect 13 2753 27 2767
rect 53 2753 67 2767
rect 92 2753 106 2767
rect 213 2752 227 2766
rect 392 2753 406 2767
rect 453 2753 467 2767
rect 533 2773 547 2787
rect 593 2753 607 2767
rect 952 2773 966 2787
rect 1113 2793 1127 2807
rect 1213 2793 1227 2807
rect 2033 2793 2047 2807
rect 2473 2793 2487 2807
rect 2853 2793 2867 2807
rect 2993 2793 3007 2807
rect 3333 2793 3347 2807
rect 3613 2793 3627 2807
rect 3673 2793 3687 2807
rect 3873 2793 3887 2807
rect 4053 2793 4067 2807
rect 4093 2793 4107 2807
rect 4393 2813 4407 2827
rect 4813 2813 4827 2827
rect 4893 2813 4907 2827
rect 5033 2813 5047 2827
rect 5373 2813 5387 2827
rect 1673 2773 1687 2787
rect 1853 2773 1867 2787
rect 1893 2773 1907 2787
rect 2172 2773 2186 2787
rect 2194 2773 2208 2787
rect 2373 2773 2387 2787
rect 2434 2773 2448 2787
rect 2593 2773 2607 2787
rect 2853 2773 2867 2787
rect 3093 2773 3107 2787
rect 933 2753 947 2767
rect 973 2753 987 2767
rect 1054 2753 1068 2767
rect 1232 2753 1246 2767
rect 1273 2753 1287 2767
rect 1453 2753 1467 2767
rect 1653 2753 1667 2767
rect 1693 2753 1707 2767
rect 2153 2753 2167 2767
rect 2753 2753 2767 2767
rect 2933 2753 2947 2767
rect 3033 2753 3047 2767
rect 3893 2773 3907 2787
rect 3594 2753 3608 2767
rect 3733 2753 3747 2767
rect 3933 2753 3947 2767
rect 4053 2773 4067 2787
rect 4253 2773 4267 2787
rect 4453 2793 4467 2807
rect 4513 2793 4527 2807
rect 4673 2793 4687 2807
rect 4013 2753 4027 2767
rect 4113 2753 4127 2767
rect 4193 2753 4207 2767
rect 4333 2753 4347 2767
rect 33 2733 47 2747
rect 152 2733 166 2747
rect 293 2733 307 2747
rect 373 2733 387 2747
rect 433 2733 447 2747
rect 553 2713 567 2727
rect 653 2733 667 2747
rect 733 2733 747 2747
rect 872 2733 886 2747
rect 1353 2733 1367 2747
rect 1514 2733 1528 2747
rect 1833 2733 1847 2747
rect 1933 2733 1947 2747
rect 1993 2733 2007 2747
rect 2113 2733 2127 2747
rect 2313 2733 2327 2747
rect 2373 2733 2387 2747
rect 2533 2733 2547 2747
rect 2574 2733 2588 2747
rect 2773 2733 2787 2747
rect 2893 2733 2907 2747
rect 2993 2733 3007 2747
rect 233 2693 247 2707
rect 453 2693 467 2707
rect 1012 2713 1026 2727
rect 1034 2713 1048 2727
rect 1113 2713 1127 2727
rect 1713 2713 1727 2727
rect 1773 2713 1787 2727
rect 1873 2713 1887 2727
rect 1953 2713 1967 2727
rect 2733 2713 2747 2727
rect 2193 2693 2207 2707
rect 2273 2693 2287 2707
rect 2393 2693 2407 2707
rect 2773 2693 2787 2707
rect 2853 2713 2867 2727
rect 3233 2713 3247 2727
rect 3333 2733 3347 2747
rect 3653 2734 3667 2748
rect 4573 2773 4587 2787
rect 4873 2773 4887 2787
rect 4973 2793 4987 2807
rect 5054 2773 5068 2787
rect 5193 2793 5207 2807
rect 5713 2813 5727 2827
rect 5413 2793 5427 2807
rect 5313 2773 5327 2787
rect 5353 2773 5367 2787
rect 5513 2793 5527 2807
rect 4634 2753 4648 2767
rect 4813 2753 4827 2767
rect 5032 2753 5046 2767
rect 5172 2753 5186 2767
rect 5213 2753 5227 2767
rect 5413 2753 5427 2767
rect 5453 2753 5467 2767
rect 5514 2753 5528 2767
rect 5653 2753 5667 2767
rect 5713 2753 5727 2767
rect 3773 2733 3787 2747
rect 3833 2733 3847 2747
rect 4054 2733 4068 2747
rect 4173 2733 4187 2747
rect 3273 2713 3287 2727
rect 3653 2712 3667 2726
rect 4133 2713 4147 2727
rect 4273 2713 4287 2727
rect 4533 2733 4547 2747
rect 4612 2733 4626 2747
rect 4673 2733 4687 2747
rect 4733 2733 4747 2747
rect 4872 2733 4886 2747
rect 4973 2733 4987 2747
rect 5013 2733 5027 2747
rect 5193 2733 5207 2747
rect 5353 2733 5367 2747
rect 4413 2713 4427 2727
rect 4793 2713 4807 2727
rect 5633 2713 5647 2727
rect 5673 2713 5687 2727
rect 2953 2693 2967 2707
rect 3413 2693 3427 2707
rect 3933 2693 3947 2707
rect 4173 2693 4187 2707
rect 4733 2693 4747 2707
rect 4853 2693 4867 2707
rect 5093 2693 5107 2707
rect 5193 2693 5207 2707
rect 13 2673 27 2687
rect 2733 2673 2747 2687
rect 2853 2673 2867 2687
rect 2933 2673 2947 2687
rect 3053 2673 3067 2687
rect 3393 2673 3407 2687
rect 3833 2673 3847 2687
rect 4053 2673 4067 2687
rect 4252 2673 4266 2687
rect 4274 2673 4288 2687
rect 4593 2673 4607 2687
rect 4633 2673 4647 2687
rect 4793 2673 4807 2687
rect 4993 2673 5007 2687
rect 5354 2673 5368 2687
rect 5453 2673 5467 2687
rect 5673 2673 5687 2687
rect 33 2653 47 2667
rect 1073 2653 1087 2667
rect 1653 2653 1667 2667
rect 1813 2653 1827 2667
rect 1853 2653 1867 2667
rect 2313 2653 2327 2667
rect 2573 2653 2587 2667
rect 3293 2653 3307 2667
rect 3433 2653 3447 2667
rect 3773 2653 3787 2667
rect 4193 2653 4207 2667
rect 4313 2653 4327 2667
rect 4693 2653 4707 2667
rect 4753 2653 4767 2667
rect 4873 2653 4887 2667
rect 4953 2653 4967 2667
rect 5152 2653 5166 2667
rect 5174 2653 5188 2667
rect 5253 2653 5267 2667
rect 5313 2653 5327 2667
rect 5713 2653 5727 2667
rect 633 2633 647 2647
rect 713 2633 727 2647
rect 833 2633 847 2647
rect 1013 2633 1027 2647
rect 1453 2633 1467 2647
rect 1693 2633 1707 2647
rect 1773 2633 1787 2647
rect 2493 2633 2507 2647
rect 2913 2633 2927 2647
rect 3033 2633 3047 2647
rect 3073 2633 3087 2647
rect 3233 2633 3247 2647
rect 3273 2633 3287 2647
rect 3333 2633 3347 2647
rect 433 2613 447 2627
rect 573 2613 587 2627
rect 793 2613 807 2627
rect 973 2613 987 2627
rect 1193 2613 1207 2627
rect 1393 2613 1407 2627
rect 1513 2613 1527 2627
rect 1613 2613 1627 2627
rect 2153 2613 2167 2627
rect 2353 2613 2367 2627
rect 2453 2613 2467 2627
rect 2793 2613 2807 2627
rect 2873 2613 2887 2627
rect 3213 2613 3227 2627
rect 3413 2633 3427 2647
rect 3533 2633 3547 2647
rect 4293 2633 4307 2647
rect 4433 2633 4447 2647
rect 4573 2633 4587 2647
rect 4853 2633 4867 2647
rect 5393 2633 5407 2647
rect 5473 2633 5487 2647
rect 3433 2613 3447 2627
rect 3573 2613 3587 2627
rect 3633 2614 3647 2628
rect 3933 2613 3947 2627
rect 4052 2613 4066 2627
rect 4393 2613 4407 2627
rect 4593 2613 4607 2627
rect 5073 2613 5087 2627
rect 133 2593 147 2607
rect 173 2593 187 2607
rect 493 2593 507 2607
rect 93 2573 107 2587
rect 293 2573 307 2587
rect 334 2573 348 2587
rect 853 2593 867 2607
rect 1693 2593 1707 2607
rect 1773 2593 1787 2607
rect 1873 2593 1887 2607
rect 1973 2593 1987 2607
rect 2133 2593 2147 2607
rect 2233 2593 2247 2607
rect 2433 2593 2447 2607
rect 2553 2593 2567 2607
rect 3353 2593 3367 2607
rect 3453 2593 3467 2607
rect 3633 2592 3647 2606
rect 4173 2593 4187 2607
rect 4573 2593 4587 2607
rect 793 2573 807 2587
rect 933 2573 947 2587
rect 1373 2573 1387 2587
rect 1533 2573 1547 2587
rect 1773 2573 1787 2587
rect 1933 2573 1947 2587
rect 93 2553 107 2567
rect 133 2553 147 2567
rect 192 2553 206 2567
rect 172 2533 186 2547
rect 312 2553 326 2567
rect 393 2553 407 2567
rect 473 2553 487 2567
rect 573 2553 587 2567
rect 633 2553 647 2567
rect 1033 2553 1047 2567
rect 1152 2553 1166 2567
rect 1313 2553 1327 2567
rect 1613 2553 1627 2567
rect 214 2533 228 2547
rect 333 2533 347 2547
rect 433 2533 447 2547
rect 33 2513 47 2527
rect 113 2513 127 2527
rect 213 2513 227 2527
rect 553 2513 567 2527
rect 673 2513 687 2527
rect 1133 2533 1147 2547
rect 1193 2533 1207 2547
rect 1433 2533 1447 2547
rect 1513 2533 1527 2547
rect 1752 2553 1766 2567
rect 1833 2553 1847 2567
rect 2193 2573 2207 2587
rect 2273 2573 2287 2587
rect 2313 2573 2327 2587
rect 2513 2573 2527 2587
rect 2093 2553 2107 2567
rect 2174 2553 2188 2567
rect 2353 2553 2367 2567
rect 2413 2553 2427 2567
rect 2573 2573 2587 2587
rect 2973 2553 2987 2567
rect 3073 2553 3087 2567
rect 3292 2553 3306 2567
rect 3593 2573 3607 2587
rect 3413 2553 3427 2567
rect 3633 2573 3647 2587
rect 4073 2573 4087 2587
rect 4413 2573 4427 2587
rect 4453 2574 4467 2588
rect 5353 2593 5367 2607
rect 4813 2573 4827 2587
rect 3833 2553 3847 2567
rect 3893 2553 3907 2567
rect 1733 2533 1747 2547
rect 1813 2533 1827 2547
rect 1993 2533 2007 2547
rect 2152 2533 2166 2547
rect 2313 2533 2327 2547
rect 2453 2533 2467 2547
rect 2593 2533 2607 2547
rect 2912 2533 2926 2547
rect 2993 2533 3007 2547
rect 3133 2533 3147 2547
rect 4053 2553 4067 2567
rect 4092 2553 4106 2567
rect 4132 2553 4146 2567
rect 4234 2553 4248 2567
rect 4453 2552 4467 2566
rect 4693 2553 4707 2567
rect 4733 2553 4747 2567
rect 5273 2573 5287 2587
rect 5333 2574 5347 2588
rect 5453 2593 5467 2607
rect 5553 2594 5567 2608
rect 5673 2593 5687 2607
rect 5433 2573 5447 2587
rect 5553 2572 5567 2586
rect 5693 2573 5707 2587
rect 5113 2553 5127 2567
rect 5213 2553 5227 2567
rect 5353 2553 5367 2567
rect 5513 2553 5527 2567
rect 5653 2553 5667 2567
rect 3434 2533 3448 2547
rect 3653 2533 3667 2547
rect 3793 2533 3807 2547
rect 713 2513 727 2527
rect 793 2513 807 2527
rect 833 2513 847 2527
rect 893 2513 907 2527
rect 1013 2513 1027 2527
rect 1253 2513 1267 2527
rect 1573 2513 1587 2527
rect 1773 2513 1787 2527
rect 1873 2513 1887 2527
rect 1913 2513 1927 2527
rect 1973 2513 1987 2527
rect 2053 2513 2067 2527
rect 2673 2513 2687 2527
rect 2873 2513 2887 2527
rect 3253 2513 3267 2527
rect 3353 2513 3367 2527
rect 3452 2513 3466 2527
rect 3474 2513 3488 2527
rect 3553 2513 3567 2527
rect 3993 2533 4007 2547
rect 4193 2533 4207 2547
rect 4292 2533 4306 2547
rect 4413 2533 4427 2547
rect 4573 2533 4587 2547
rect 4773 2533 4787 2547
rect 4314 2513 4328 2527
rect 393 2493 407 2507
rect 673 2493 687 2507
rect 913 2493 927 2507
rect 1033 2493 1047 2507
rect 1193 2493 1207 2507
rect 1313 2493 1327 2507
rect 1533 2493 1547 2507
rect 1893 2493 1907 2507
rect 1953 2493 1967 2507
rect 2093 2493 2107 2507
rect 2153 2493 2167 2507
rect 2293 2493 2307 2507
rect 313 2473 327 2487
rect 493 2473 507 2487
rect 753 2473 767 2487
rect 893 2473 907 2487
rect 993 2473 1007 2487
rect 1073 2473 1087 2487
rect 3433 2493 3447 2507
rect 3693 2493 3707 2507
rect 4133 2493 4147 2507
rect 2453 2473 2467 2487
rect 2813 2474 2827 2488
rect 3253 2473 3267 2487
rect 3413 2473 3427 2487
rect 4093 2473 4107 2487
rect 4153 2473 4167 2487
rect 4273 2493 4287 2507
rect 4613 2513 4627 2527
rect 4693 2513 4707 2527
rect 4853 2513 4867 2527
rect 5154 2513 5168 2527
rect 5473 2533 5487 2547
rect 5393 2513 5407 2527
rect 5513 2513 5527 2527
rect 5673 2513 5687 2527
rect 4413 2493 4427 2507
rect 4473 2493 4487 2507
rect 4553 2493 4567 2507
rect 4713 2493 4727 2507
rect 4753 2493 4767 2507
rect 4893 2493 4907 2507
rect 4973 2493 4987 2507
rect 5093 2493 5107 2507
rect 5613 2493 5627 2507
rect 5693 2493 5707 2507
rect 4433 2473 4447 2487
rect 4493 2473 4507 2487
rect 4633 2473 4647 2487
rect 4733 2473 4747 2487
rect 5633 2473 5647 2487
rect 1253 2453 1267 2467
rect 1433 2453 1447 2467
rect 1733 2453 1747 2467
rect 2033 2453 2047 2467
rect 2193 2453 2207 2467
rect 2813 2452 2827 2466
rect 2913 2453 2927 2467
rect 3313 2453 3327 2467
rect 4013 2453 4027 2467
rect 93 2433 107 2447
rect 173 2433 187 2447
rect 773 2433 787 2447
rect 873 2433 887 2447
rect 1193 2433 1207 2447
rect 1413 2433 1427 2447
rect 2473 2433 2487 2447
rect 2733 2433 2747 2447
rect 3133 2433 3147 2447
rect 3213 2433 3227 2447
rect 3513 2433 3527 2447
rect 3733 2433 3747 2447
rect 3813 2433 3827 2447
rect 4173 2433 4187 2447
rect 4313 2433 4327 2447
rect 4513 2433 4527 2447
rect 4673 2433 4687 2447
rect 4873 2433 4887 2447
rect 5153 2453 5167 2467
rect 5313 2453 5327 2467
rect 5473 2453 5487 2467
rect 5533 2453 5547 2467
rect 5713 2453 5727 2467
rect 493 2413 507 2427
rect 833 2413 847 2427
rect 973 2413 987 2427
rect 2493 2413 2507 2427
rect 3393 2413 3407 2427
rect 3493 2413 3507 2427
rect 3753 2413 3767 2427
rect 4253 2413 4267 2427
rect 4713 2413 4727 2427
rect 4773 2413 4787 2427
rect 5333 2433 5347 2447
rect 5273 2413 5287 2427
rect 5633 2413 5647 2427
rect 253 2393 267 2407
rect 453 2393 467 2407
rect 653 2393 667 2407
rect 913 2393 927 2407
rect 1593 2393 1607 2407
rect 1673 2394 1687 2408
rect 1893 2393 1907 2407
rect 2873 2393 2887 2407
rect 2913 2393 2927 2407
rect 3093 2393 3107 2407
rect 3712 2393 3726 2407
rect 3734 2393 3748 2407
rect 3913 2393 3927 2407
rect 4273 2393 4287 2407
rect 4533 2393 4547 2407
rect 4693 2393 4707 2407
rect 5053 2393 5067 2407
rect 533 2373 547 2387
rect 693 2373 707 2387
rect 1153 2373 1167 2387
rect 1673 2372 1687 2386
rect 1753 2373 1767 2387
rect 3653 2373 3667 2387
rect 3853 2373 3867 2387
rect 3993 2374 4007 2388
rect 4293 2373 4307 2387
rect 4373 2373 4387 2387
rect 5213 2393 5227 2407
rect 5493 2393 5507 2407
rect 5713 2393 5727 2407
rect 5153 2373 5167 2387
rect 5313 2373 5327 2387
rect 5373 2373 5387 2387
rect 5453 2373 5467 2387
rect 5673 2373 5687 2387
rect 433 2353 447 2367
rect 553 2353 567 2367
rect 793 2353 807 2367
rect 893 2353 907 2367
rect 1393 2353 1407 2367
rect 2513 2353 2527 2367
rect 2593 2353 2607 2367
rect 2873 2353 2887 2367
rect 3173 2353 3187 2367
rect 3673 2353 3687 2367
rect 3773 2353 3787 2367
rect 3893 2353 3907 2367
rect 3993 2352 4007 2366
rect 4093 2353 4107 2367
rect 4133 2353 4147 2367
rect 4413 2353 4427 2367
rect 4613 2353 4627 2367
rect 4833 2353 4847 2367
rect 4933 2353 4947 2367
rect 513 2333 527 2347
rect 573 2333 587 2347
rect 853 2333 867 2347
rect 1233 2333 1247 2347
rect 1993 2333 2007 2347
rect 2133 2333 2147 2347
rect 2173 2333 2187 2347
rect 2353 2334 2367 2348
rect 3053 2333 3067 2347
rect 3973 2333 3987 2347
rect 4153 2333 4167 2347
rect 4213 2333 4227 2347
rect 4353 2333 4367 2347
rect 4433 2333 4447 2347
rect 4553 2333 4567 2347
rect 4673 2333 4687 2347
rect 4713 2333 4727 2347
rect 5193 2333 5207 2347
rect 5713 2353 5727 2367
rect 5453 2333 5467 2347
rect 5552 2333 5566 2347
rect 5574 2333 5588 2347
rect 5673 2333 5687 2347
rect 153 2313 167 2327
rect 53 2293 67 2307
rect 94 2294 108 2308
rect 153 2273 167 2287
rect 193 2274 207 2288
rect 313 2274 327 2288
rect 613 2313 627 2327
rect 772 2313 786 2327
rect 794 2313 808 2327
rect 493 2294 507 2308
rect 713 2293 727 2307
rect 973 2313 987 2327
rect 1033 2313 1047 2327
rect 1173 2313 1187 2327
rect 914 2293 928 2307
rect 372 2273 386 2287
rect 493 2272 507 2286
rect 613 2273 627 2287
rect 654 2274 668 2288
rect 993 2293 1007 2307
rect 1233 2313 1247 2327
rect 1313 2313 1327 2327
rect 1513 2313 1527 2327
rect 1553 2313 1567 2327
rect 1773 2313 1787 2327
rect 1373 2293 1387 2307
rect 1493 2293 1507 2307
rect 1613 2293 1627 2307
rect 2353 2312 2367 2326
rect 2433 2313 2447 2327
rect 2513 2313 2527 2327
rect 694 2273 708 2287
rect 892 2273 906 2287
rect 1033 2273 1047 2287
rect 1133 2273 1147 2287
rect 1173 2273 1187 2287
rect 1353 2273 1367 2287
rect 1433 2273 1447 2287
rect 1613 2273 1627 2287
rect 1693 2273 1707 2287
rect 1813 2273 1827 2287
rect 93 2253 107 2267
rect 193 2252 207 2266
rect 313 2252 327 2266
rect 672 2253 686 2267
rect 1972 2293 1986 2307
rect 1994 2293 2008 2307
rect 2053 2293 2067 2307
rect 2193 2294 2207 2308
rect 2733 2313 2747 2327
rect 2933 2313 2947 2327
rect 3373 2313 3387 2327
rect 2493 2293 2507 2307
rect 2573 2293 2587 2307
rect 2653 2293 2667 2307
rect 3233 2293 3247 2307
rect 3273 2293 3287 2307
rect 3433 2293 3447 2307
rect 3533 2293 3547 2307
rect 3733 2313 3747 2327
rect 3892 2313 3906 2327
rect 3914 2313 3928 2327
rect 4073 2313 4087 2327
rect 4113 2313 4127 2327
rect 4193 2313 4207 2327
rect 4233 2313 4247 2327
rect 4413 2313 4427 2327
rect 4833 2313 4847 2327
rect 5033 2313 5047 2327
rect 5373 2313 5387 2327
rect 5433 2313 5447 2327
rect 3613 2293 3627 2307
rect 3973 2293 3987 2307
rect 1933 2273 1947 2287
rect 2193 2272 2207 2286
rect 2373 2273 2387 2287
rect 2593 2273 2607 2287
rect 2713 2273 2727 2287
rect 2813 2273 2827 2287
rect 2973 2273 2987 2287
rect 853 2253 867 2267
rect 1253 2253 1267 2267
rect 1553 2253 1567 2267
rect 1852 2253 1866 2267
rect 1892 2253 1906 2267
rect 1953 2253 1967 2267
rect 2053 2253 2067 2267
rect 2292 2253 2306 2267
rect 2333 2253 2347 2267
rect 4113 2293 4127 2307
rect 4313 2293 4327 2307
rect 4353 2293 4367 2307
rect 4513 2293 4527 2307
rect 3593 2273 3607 2287
rect 3734 2273 3748 2287
rect 3852 2273 3866 2287
rect 3893 2273 3907 2287
rect 4173 2273 4187 2287
rect 2853 2253 2867 2267
rect 3033 2253 3047 2267
rect 3094 2253 3108 2267
rect 3173 2253 3187 2267
rect 3372 2253 3386 2267
rect 3433 2253 3447 2267
rect 3492 2253 3506 2267
rect 3913 2253 3927 2267
rect 4553 2293 4567 2307
rect 4613 2293 4627 2307
rect 4713 2293 4727 2307
rect 4873 2293 4887 2307
rect 4973 2293 4987 2307
rect 4672 2274 4686 2288
rect 5213 2293 5227 2307
rect 5313 2293 5327 2307
rect 5413 2293 5427 2307
rect 5533 2293 5547 2307
rect 4812 2273 4826 2287
rect 4853 2273 4867 2287
rect 4913 2273 4927 2287
rect 5153 2273 5167 2287
rect 5252 2273 5266 2287
rect 5294 2273 5308 2287
rect 5493 2273 5507 2287
rect 4252 2253 4266 2267
rect 4313 2253 4327 2267
rect 833 2233 847 2247
rect 1053 2233 1067 2247
rect 1353 2233 1367 2247
rect 1513 2233 1527 2247
rect 1773 2233 1787 2247
rect 2513 2233 2527 2247
rect 2953 2233 2967 2247
rect 3053 2233 3067 2247
rect 3233 2234 3247 2248
rect 3413 2233 3427 2247
rect 3493 2233 3507 2247
rect 3533 2233 3547 2247
rect 3693 2233 3707 2247
rect 3853 2233 3867 2247
rect 4033 2233 4047 2247
rect 4093 2233 4107 2247
rect 793 2213 807 2227
rect 1413 2213 1427 2227
rect 3233 2212 3247 2226
rect 4514 2252 4528 2266
rect 4813 2253 4827 2267
rect 4973 2253 4987 2267
rect 5012 2253 5026 2267
rect 5034 2253 5048 2267
rect 5074 2254 5088 2268
rect 5313 2253 5327 2267
rect 5353 2253 5367 2267
rect 5473 2253 5487 2267
rect 5532 2253 5546 2267
rect 5573 2253 5587 2267
rect 4573 2233 4587 2247
rect 4673 2233 4687 2247
rect 4833 2233 4847 2247
rect 4953 2233 4967 2247
rect 5073 2232 5087 2246
rect 5233 2233 5247 2247
rect 5333 2233 5347 2247
rect 5453 2233 5467 2247
rect 3633 2213 3647 2227
rect 3933 2213 3947 2227
rect 4073 2213 4087 2227
rect 4193 2213 4207 2227
rect 4553 2213 4567 2227
rect 4653 2213 4667 2227
rect 4913 2213 4927 2227
rect 5033 2213 5047 2227
rect 5173 2213 5187 2227
rect 5473 2213 5487 2227
rect 5533 2213 5547 2227
rect 313 2193 327 2207
rect 753 2193 767 2207
rect 1573 2193 1587 2207
rect 1853 2193 1867 2207
rect 2233 2193 2247 2207
rect 2553 2193 2567 2207
rect 2753 2193 2767 2207
rect 2833 2193 2847 2207
rect 3473 2193 3487 2207
rect 3833 2193 3847 2207
rect 4033 2193 4047 2207
rect 4493 2193 4507 2207
rect 5133 2193 5147 2207
rect 5253 2193 5267 2207
rect 5393 2193 5407 2207
rect 1213 2173 1227 2187
rect 1253 2173 1267 2187
rect 1433 2173 1447 2187
rect 2373 2173 2387 2187
rect 2473 2173 2487 2187
rect 2513 2173 2527 2187
rect 2913 2173 2927 2187
rect 2953 2173 2967 2187
rect 3413 2173 3427 2187
rect 3513 2173 3527 2187
rect 1233 2153 1247 2167
rect 1273 2153 1287 2167
rect 1353 2153 1367 2167
rect 1973 2153 1987 2167
rect 2073 2153 2087 2167
rect 3753 2173 3767 2187
rect 4113 2173 4127 2187
rect 4153 2173 4167 2187
rect 4993 2173 5007 2187
rect 5233 2173 5247 2187
rect 5413 2173 5427 2187
rect 5613 2173 5627 2187
rect 3313 2153 3327 2167
rect 3373 2153 3387 2167
rect 3653 2153 3667 2167
rect 3693 2153 3707 2167
rect 3913 2153 3927 2167
rect 3973 2153 3987 2167
rect 4013 2153 4027 2167
rect 4053 2153 4067 2167
rect 4453 2154 4467 2168
rect 4553 2153 4567 2167
rect 4673 2153 4687 2167
rect 4852 2153 4866 2167
rect 4874 2153 4888 2167
rect 4913 2153 4927 2167
rect 33 2133 47 2147
rect 113 2133 127 2147
rect 433 2133 447 2147
rect 1653 2133 1667 2147
rect 1893 2133 1907 2147
rect 2013 2133 2027 2147
rect 2813 2133 2827 2147
rect 2933 2133 2947 2147
rect 3093 2133 3107 2147
rect 3273 2133 3287 2147
rect 3593 2133 3607 2147
rect 4153 2133 4167 2147
rect 4293 2133 4307 2147
rect 4453 2132 4467 2146
rect 4613 2133 4627 2147
rect 4653 2133 4667 2147
rect 4813 2133 4827 2147
rect 5133 2153 5147 2167
rect 5473 2153 5487 2167
rect 73 2113 87 2127
rect 153 2113 167 2127
rect 233 2113 247 2127
rect 373 2113 387 2127
rect 413 2113 427 2127
rect 713 2113 727 2127
rect 953 2113 967 2127
rect 1153 2113 1167 2127
rect 1273 2113 1287 2127
rect 1493 2113 1507 2127
rect 1713 2113 1727 2127
rect 2093 2113 2107 2127
rect 2253 2113 2267 2127
rect 2433 2113 2447 2127
rect 2513 2113 2527 2127
rect 3213 2113 3227 2127
rect 3333 2113 3347 2127
rect 3713 2113 3727 2127
rect 3813 2113 3827 2127
rect 3972 2113 3986 2127
rect 3994 2113 4008 2127
rect 114 2093 128 2107
rect 173 2093 187 2107
rect 92 2073 106 2087
rect 233 2073 247 2087
rect 273 2073 287 2087
rect 413 2074 427 2088
rect 793 2093 807 2107
rect 853 2093 867 2107
rect 993 2093 1007 2107
rect 1113 2093 1127 2107
rect 453 2073 467 2087
rect 573 2073 587 2087
rect 1153 2073 1167 2087
rect 1333 2093 1347 2107
rect 1453 2093 1467 2107
rect 1553 2093 1567 2107
rect 33 2053 47 2067
rect 172 2053 186 2067
rect 293 2053 307 2067
rect 394 2053 408 2067
rect 473 2033 487 2047
rect 674 2053 688 2067
rect 953 2053 967 2067
rect 1493 2073 1507 2087
rect 1653 2093 1667 2107
rect 1693 2093 1707 2107
rect 1813 2093 1827 2107
rect 1873 2093 1887 2107
rect 1713 2073 1727 2087
rect 1893 2073 1907 2087
rect 2073 2093 2087 2107
rect 2113 2093 2127 2107
rect 2453 2073 2467 2087
rect 2813 2093 2827 2107
rect 3013 2093 3027 2107
rect 3133 2093 3147 2107
rect 2533 2073 2547 2087
rect 2573 2074 2587 2088
rect 2693 2073 2707 2087
rect 3033 2073 3047 2087
rect 3112 2074 3126 2088
rect 3433 2093 3447 2107
rect 3613 2093 3627 2107
rect 3673 2093 3687 2107
rect 4013 2093 4027 2107
rect 4053 2093 4067 2107
rect 3512 2073 3526 2087
rect 3553 2073 3567 2087
rect 3792 2073 3806 2087
rect 3814 2073 3828 2087
rect 3953 2073 3967 2087
rect 4173 2073 4187 2087
rect 4433 2114 4447 2128
rect 4493 2113 4507 2127
rect 4573 2113 4587 2127
rect 4713 2113 4727 2127
rect 4253 2073 4267 2087
rect 4433 2092 4447 2106
rect 4973 2113 4987 2127
rect 5093 2113 5107 2127
rect 5233 2113 5247 2127
rect 5313 2133 5327 2147
rect 5373 2133 5387 2147
rect 5354 2113 5368 2127
rect 5453 2113 5467 2127
rect 5513 2113 5527 2127
rect 5593 2113 5607 2127
rect 4753 2093 4767 2107
rect 4813 2093 4827 2107
rect 5553 2093 5567 2107
rect 5713 2093 5727 2107
rect 4313 2073 4327 2087
rect 4413 2073 4427 2087
rect 4473 2073 4487 2087
rect 4553 2073 4567 2087
rect 4713 2073 4727 2087
rect 4833 2073 4847 2087
rect 4953 2073 4967 2087
rect 5173 2073 5187 2087
rect 5254 2073 5268 2087
rect 5294 2073 5308 2087
rect 5553 2073 5567 2087
rect 1273 2053 1287 2067
rect 1353 2053 1367 2067
rect 1473 2053 1487 2067
rect 1513 2053 1527 2067
rect 1673 2053 1687 2067
rect 1753 2053 1767 2067
rect 1832 2053 1846 2067
rect 2033 2053 2047 2067
rect 533 2033 547 2047
rect 733 2033 747 2047
rect 813 2033 827 2047
rect 853 2033 867 2047
rect 33 2013 47 2027
rect 913 2013 927 2027
rect 1073 2033 1087 2047
rect 1333 2032 1347 2046
rect 1633 2033 1647 2047
rect 1694 2033 1708 2047
rect 1972 2033 1986 2047
rect 2093 2033 2107 2047
rect 2433 2053 2447 2067
rect 2593 2053 2607 2067
rect 2633 2053 2647 2067
rect 2713 2053 2727 2067
rect 2792 2053 2806 2067
rect 2814 2053 2828 2067
rect 2933 2053 2947 2067
rect 3093 2052 3107 2066
rect 3274 2053 3288 2067
rect 3413 2053 3427 2067
rect 2133 2033 2147 2047
rect 2213 2033 2227 2047
rect 2853 2033 2867 2047
rect 2993 2033 3007 2047
rect 3213 2033 3227 2047
rect 3513 2033 3527 2047
rect 3593 2053 3607 2067
rect 3853 2053 3867 2067
rect 3892 2053 3906 2067
rect 3933 2053 3947 2067
rect 4033 2053 4047 2067
rect 4074 2053 4088 2067
rect 4353 2053 4367 2067
rect 4493 2053 4507 2067
rect 4533 2053 4547 2067
rect 5053 2053 5067 2067
rect 2112 2013 2126 2027
rect 2134 2013 2148 2027
rect 2773 2013 2787 2027
rect 3373 2013 3387 2027
rect 3733 2033 3747 2047
rect 3833 2032 3847 2046
rect 4153 2033 4167 2047
rect 4193 2033 4207 2047
rect 4373 2033 4387 2047
rect 4673 2033 4687 2047
rect 4814 2033 4828 2047
rect 4874 2033 4888 2047
rect 4914 2033 4928 2047
rect 5132 2053 5146 2067
rect 5353 2053 5367 2067
rect 5573 2053 5587 2067
rect 5673 2053 5687 2067
rect 573 1993 587 2007
rect 913 1993 927 2007
rect 1573 1993 1587 2007
rect 1673 1993 1687 2007
rect 1993 1993 2007 2007
rect 3574 2013 3588 2027
rect 3633 2013 3647 2027
rect 2673 1993 2687 2007
rect 2813 1993 2827 2007
rect 2873 1993 2887 2007
rect 3553 1993 3567 2007
rect 3973 2013 3987 2027
rect 4253 2013 4267 2027
rect 4333 2013 4347 2027
rect 4573 2013 4587 2027
rect 4653 2013 4667 2027
rect 5173 2014 5187 2028
rect 5333 2033 5347 2047
rect 5533 2033 5547 2047
rect 5633 2033 5647 2047
rect 5293 2013 5307 2027
rect 5613 2013 5627 2027
rect 5653 2013 5667 2027
rect 4033 1993 4047 2007
rect 4173 1994 4187 2008
rect 4313 1993 4327 2007
rect 4473 1993 4487 2007
rect 4593 1993 4607 2007
rect 4673 1993 4687 2007
rect 5133 1993 5147 2007
rect 1513 1973 1527 1987
rect 5174 1992 5188 2006
rect 5213 1993 5227 2007
rect 5353 1993 5367 2007
rect 5633 1993 5647 2007
rect 5693 1993 5707 2007
rect 2473 1973 2487 1987
rect 2513 1973 2527 1987
rect 2853 1973 2867 1987
rect 3113 1973 3127 1987
rect 3153 1973 3167 1987
rect 3313 1973 3327 1987
rect 3993 1973 4007 1987
rect 4113 1974 4127 1988
rect 4173 1972 4187 1986
rect 4293 1973 4307 1987
rect 4433 1973 4447 1987
rect 4533 1973 4547 1987
rect 373 1953 387 1967
rect 553 1953 567 1967
rect 1693 1953 1707 1967
rect 2073 1953 2087 1967
rect 2493 1953 2507 1967
rect 2813 1953 2827 1967
rect 3133 1953 3147 1967
rect 3173 1953 3187 1967
rect 3673 1953 3687 1967
rect 3833 1953 3847 1967
rect 4113 1952 4127 1966
rect 4273 1953 4287 1967
rect 4393 1953 4407 1967
rect 4853 1973 4867 1987
rect 5033 1973 5047 1987
rect 5553 1973 5567 1987
rect 5653 1973 5667 1987
rect 233 1933 247 1947
rect 673 1933 687 1947
rect 713 1933 727 1947
rect 1793 1933 1807 1947
rect 2233 1933 2247 1947
rect 2693 1933 2707 1947
rect 2913 1933 2927 1947
rect 2993 1933 3007 1947
rect 3233 1933 3247 1947
rect 3273 1933 3287 1947
rect 4013 1933 4027 1947
rect 93 1913 107 1927
rect 333 1913 347 1927
rect 533 1913 547 1927
rect 573 1913 587 1927
rect 653 1913 667 1927
rect 693 1913 707 1927
rect 733 1913 747 1927
rect 1553 1913 1567 1927
rect 2053 1913 2067 1927
rect 2113 1913 2127 1927
rect 2933 1913 2947 1927
rect 3033 1913 3047 1927
rect 3353 1913 3367 1927
rect 3413 1913 3427 1927
rect 4413 1933 4427 1947
rect 5633 1953 5647 1967
rect 5693 1953 5707 1967
rect 4893 1933 4907 1947
rect 4973 1933 4987 1947
rect 5293 1933 5307 1947
rect 4553 1913 4567 1927
rect 4772 1913 4786 1927
rect 4794 1913 4808 1927
rect 5073 1913 5087 1927
rect 5433 1913 5447 1927
rect 5613 1913 5627 1927
rect 413 1893 427 1907
rect 633 1893 647 1907
rect 753 1893 767 1907
rect 1193 1893 1207 1907
rect 1933 1893 1947 1907
rect 2153 1893 2167 1907
rect 2253 1893 2267 1907
rect 2293 1893 2307 1907
rect 2353 1893 2367 1907
rect 3053 1893 3067 1907
rect 3233 1893 3247 1907
rect 3513 1893 3527 1907
rect 3553 1893 3567 1907
rect 3733 1893 3747 1907
rect 3893 1893 3907 1907
rect 4813 1893 4827 1907
rect 4893 1893 4907 1907
rect 5133 1893 5147 1907
rect 5333 1893 5347 1907
rect 473 1873 487 1887
rect 653 1873 667 1887
rect 793 1873 807 1887
rect 893 1873 907 1887
rect 1733 1873 1747 1887
rect 1953 1873 1967 1887
rect 1993 1873 2007 1887
rect 2773 1873 2787 1887
rect 3133 1873 3147 1887
rect 3413 1873 3427 1887
rect 3473 1873 3487 1887
rect 3533 1873 3547 1887
rect 3673 1873 3687 1887
rect 3713 1873 3727 1887
rect 4033 1873 4047 1887
rect 4153 1873 4167 1887
rect 4413 1873 4427 1887
rect 4673 1873 4687 1887
rect 4912 1873 4926 1887
rect 4934 1873 4948 1887
rect 5113 1873 5127 1887
rect 5273 1873 5287 1887
rect 5473 1873 5487 1887
rect 5512 1873 5526 1887
rect 5553 1873 5567 1887
rect 93 1853 107 1867
rect 293 1853 307 1867
rect 493 1853 507 1867
rect 73 1833 87 1847
rect 153 1833 167 1847
rect 333 1833 347 1847
rect 473 1833 487 1847
rect 913 1853 927 1867
rect 1513 1853 1527 1867
rect 1752 1853 1766 1867
rect 1813 1853 1827 1867
rect 2153 1853 2167 1867
rect 2413 1853 2427 1867
rect 2593 1853 2607 1867
rect 3113 1853 3127 1867
rect 3273 1853 3287 1867
rect 3393 1853 3407 1867
rect 3773 1853 3787 1867
rect 4633 1853 4647 1867
rect 4693 1853 4707 1867
rect 4773 1853 4787 1867
rect 5193 1853 5207 1867
rect 5533 1853 5547 1867
rect 5713 1853 5727 1867
rect 913 1833 927 1847
rect 1033 1833 1047 1847
rect 1693 1833 1707 1847
rect 193 1813 207 1827
rect 293 1813 307 1827
rect 493 1813 507 1827
rect 613 1813 627 1827
rect 693 1813 707 1827
rect 753 1813 767 1827
rect 973 1813 987 1827
rect 1733 1833 1747 1847
rect 2333 1833 2347 1847
rect 2933 1833 2947 1847
rect 3153 1833 3167 1847
rect 3273 1833 3287 1847
rect 3633 1833 3647 1847
rect 3693 1833 3707 1847
rect 1873 1813 1887 1827
rect 2473 1813 2487 1827
rect 2653 1813 2667 1827
rect 2993 1813 3007 1827
rect 3153 1813 3167 1827
rect 3214 1813 3228 1827
rect 3333 1813 3347 1827
rect 3493 1813 3507 1827
rect 3573 1813 3587 1827
rect 112 1793 126 1807
rect 154 1793 168 1807
rect 332 1793 346 1807
rect 413 1793 427 1807
rect 593 1793 607 1807
rect 673 1793 687 1807
rect 92 1773 106 1787
rect 134 1773 148 1787
rect 193 1773 207 1787
rect 793 1773 807 1787
rect 893 1773 907 1787
rect 1013 1793 1027 1807
rect 1153 1793 1167 1807
rect 1313 1793 1327 1807
rect 1453 1793 1467 1807
rect 1633 1793 1647 1807
rect 1793 1793 1807 1807
rect 1933 1793 1947 1807
rect 1994 1793 2008 1807
rect 2073 1793 2087 1807
rect 2193 1793 2207 1807
rect 2233 1793 2247 1807
rect 2293 1793 2307 1807
rect 2413 1793 2427 1807
rect 2513 1793 2527 1807
rect 2593 1793 2607 1807
rect 2874 1793 2888 1807
rect 2953 1793 2967 1807
rect 3033 1793 3047 1807
rect 3093 1794 3107 1808
rect 3673 1813 3687 1827
rect 3892 1833 3906 1847
rect 4093 1833 4107 1847
rect 4273 1833 4287 1847
rect 4573 1833 4587 1847
rect 4793 1834 4807 1848
rect 4913 1833 4927 1847
rect 3813 1813 3827 1827
rect 3873 1813 3887 1827
rect 4133 1813 4147 1827
rect 4233 1813 4247 1827
rect 4493 1813 4507 1827
rect 4593 1813 4607 1827
rect 4793 1812 4807 1826
rect 4933 1813 4947 1827
rect 5013 1813 5027 1827
rect 5053 1813 5067 1827
rect 933 1773 947 1787
rect 993 1773 1007 1787
rect 1074 1773 1088 1787
rect 1133 1773 1147 1787
rect 73 1753 87 1767
rect 473 1753 487 1767
rect 513 1753 527 1767
rect 873 1753 887 1767
rect 933 1753 947 1767
rect 1073 1753 1087 1767
rect 1173 1753 1187 1767
rect 1273 1773 1287 1787
rect 1353 1773 1367 1787
rect 1533 1773 1547 1787
rect 1733 1773 1747 1787
rect 1993 1773 2007 1787
rect 2173 1773 2187 1787
rect 2352 1773 2366 1787
rect 2394 1773 2408 1787
rect 2473 1773 2487 1787
rect 2893 1773 2907 1787
rect 2973 1773 2987 1787
rect 3093 1773 3107 1786
rect 1293 1753 1307 1767
rect 1872 1753 1886 1767
rect 3093 1772 3107 1773
rect 3193 1773 3207 1787
rect 413 1733 427 1747
rect 893 1733 907 1747
rect 992 1733 1006 1747
rect 1014 1733 1028 1747
rect 1733 1733 1747 1747
rect 1873 1733 1887 1747
rect 2373 1753 2387 1767
rect 2593 1753 2607 1767
rect 2793 1753 2807 1767
rect 2853 1753 2867 1767
rect 2933 1753 2947 1767
rect 3012 1753 3026 1767
rect 3034 1753 3048 1767
rect 3233 1793 3247 1807
rect 3433 1793 3447 1807
rect 3674 1793 3688 1807
rect 3713 1793 3727 1807
rect 3794 1793 3808 1807
rect 3914 1793 3928 1807
rect 3413 1774 3427 1788
rect 4193 1793 4207 1807
rect 4353 1793 4367 1807
rect 4413 1793 4427 1807
rect 4513 1793 4527 1807
rect 3733 1773 3747 1787
rect 3774 1773 3788 1787
rect 3893 1773 3907 1787
rect 3413 1752 3427 1766
rect 3453 1754 3467 1768
rect 2733 1733 2747 1747
rect 3453 1732 3467 1746
rect 3573 1733 3587 1747
rect 3833 1753 3847 1767
rect 4033 1773 4047 1787
rect 4092 1773 4106 1787
rect 4134 1773 4148 1787
rect 4232 1773 4246 1787
rect 4373 1773 4387 1787
rect 4433 1773 4447 1787
rect 4472 1773 4486 1787
rect 4494 1773 4508 1787
rect 4613 1773 4627 1787
rect 4674 1793 4688 1807
rect 4913 1793 4927 1807
rect 4993 1793 5007 1807
rect 5093 1813 5107 1827
rect 5133 1814 5147 1828
rect 5233 1813 5247 1827
rect 5294 1813 5308 1827
rect 5593 1813 5607 1827
rect 5133 1792 5147 1806
rect 5573 1793 5587 1807
rect 5713 1793 5727 1807
rect 4733 1773 4747 1787
rect 4774 1773 4788 1787
rect 4814 1773 4828 1787
rect 4093 1753 4107 1767
rect 4233 1753 4247 1767
rect 4353 1753 4367 1767
rect 4633 1753 4647 1767
rect 4673 1753 4687 1767
rect 4913 1753 4927 1767
rect 5094 1772 5108 1786
rect 5212 1773 5226 1787
rect 5293 1773 5307 1787
rect 5433 1773 5447 1787
rect 5533 1773 5547 1787
rect 5073 1753 5087 1767
rect 5593 1753 5607 1767
rect 5633 1753 5647 1767
rect 5673 1753 5687 1767
rect 3933 1734 3947 1748
rect 4513 1733 4527 1747
rect 373 1713 387 1727
rect 693 1713 707 1727
rect 413 1693 427 1707
rect 573 1693 587 1707
rect 1173 1713 1187 1727
rect 1493 1713 1507 1727
rect 1933 1713 1947 1727
rect 2073 1713 2087 1727
rect 3053 1713 3067 1727
rect 3513 1713 3527 1727
rect 3933 1712 3947 1726
rect 3993 1713 4007 1727
rect 4133 1713 4147 1727
rect 4533 1713 4547 1727
rect 4593 1713 4607 1727
rect 5053 1733 5067 1747
rect 5132 1733 5146 1747
rect 5154 1734 5168 1748
rect 5273 1733 5287 1747
rect 5353 1733 5367 1747
rect 5413 1733 5427 1747
rect 5453 1733 5467 1747
rect 5533 1733 5547 1747
rect 5693 1734 5707 1748
rect 1053 1693 1067 1707
rect 1193 1693 1207 1707
rect 1233 1693 1247 1707
rect 1373 1693 1387 1707
rect 1633 1693 1647 1707
rect 2433 1693 2447 1707
rect 2913 1694 2927 1708
rect 3353 1693 3367 1707
rect 353 1673 367 1687
rect 553 1673 567 1687
rect 973 1673 987 1687
rect 1353 1673 1367 1687
rect 1613 1673 1627 1687
rect 1893 1673 1907 1687
rect 2053 1673 2067 1687
rect 2693 1673 2707 1687
rect 2753 1673 2767 1687
rect 2913 1672 2927 1686
rect 2953 1673 2967 1687
rect 3233 1673 3247 1687
rect 3773 1693 3787 1707
rect 4033 1693 4047 1707
rect 4373 1693 4387 1707
rect 4613 1693 4627 1707
rect 4713 1714 4727 1728
rect 4773 1713 4787 1727
rect 4953 1713 4967 1727
rect 4713 1692 4727 1706
rect 4993 1693 5007 1707
rect 5153 1712 5167 1726
rect 5213 1713 5227 1727
rect 5313 1713 5327 1727
rect 5553 1713 5567 1727
rect 5693 1712 5707 1726
rect 5353 1693 5367 1707
rect 5412 1693 5426 1707
rect 5434 1694 5448 1708
rect 5513 1693 5527 1707
rect 5633 1693 5647 1707
rect 3653 1673 3667 1687
rect 3793 1673 3807 1687
rect 3953 1673 3967 1687
rect 4493 1673 4507 1687
rect 4633 1674 4647 1688
rect 4793 1673 4807 1687
rect 5033 1673 5047 1687
rect 5273 1673 5287 1687
rect 5433 1672 5447 1686
rect 5553 1673 5567 1687
rect 5673 1673 5687 1687
rect 5713 1673 5727 1687
rect 193 1653 207 1667
rect 533 1653 547 1667
rect 1313 1653 1327 1667
rect 1653 1653 1667 1667
rect 1913 1653 1927 1667
rect 2453 1653 2467 1667
rect 2773 1653 2787 1667
rect 3133 1653 3147 1667
rect 113 1633 127 1647
rect 313 1613 327 1627
rect 473 1613 487 1627
rect 653 1633 667 1647
rect 833 1633 847 1647
rect 1053 1633 1067 1647
rect 1573 1634 1587 1648
rect 1693 1633 1707 1647
rect 1753 1633 1767 1647
rect 2293 1633 2307 1647
rect 2893 1634 2907 1648
rect 3493 1653 3507 1667
rect 3893 1653 3907 1667
rect 4333 1653 4347 1667
rect 4533 1653 4547 1667
rect 4632 1652 4646 1666
rect 4713 1653 4727 1667
rect 4853 1653 4867 1667
rect 4953 1653 4967 1667
rect 5473 1653 5487 1667
rect 5593 1653 5607 1667
rect 3393 1633 3407 1647
rect 4213 1634 4227 1648
rect 5153 1633 5167 1647
rect 33 1593 47 1607
rect 193 1593 207 1607
rect 232 1593 246 1607
rect 353 1593 367 1607
rect 473 1593 487 1607
rect 133 1573 147 1587
rect 333 1573 347 1587
rect 433 1573 447 1587
rect 573 1593 587 1607
rect 653 1593 667 1607
rect 733 1613 747 1627
rect 774 1593 788 1607
rect 834 1593 848 1607
rect 933 1613 947 1627
rect 1133 1613 1147 1627
rect 1273 1613 1287 1627
rect 1453 1613 1467 1627
rect 1573 1612 1587 1626
rect 1873 1613 1887 1627
rect 1933 1613 1947 1627
rect 2133 1613 2147 1627
rect 2193 1613 2207 1627
rect 2853 1613 2867 1627
rect 2893 1612 2907 1626
rect 3033 1614 3047 1628
rect 3233 1613 3247 1627
rect 1012 1593 1026 1607
rect 1034 1593 1048 1607
rect 1153 1593 1167 1607
rect 1233 1573 1247 1587
rect 1413 1593 1427 1607
rect 1474 1593 1488 1607
rect 1873 1593 1887 1607
rect 1333 1573 1347 1587
rect 1453 1573 1467 1587
rect 1573 1573 1587 1587
rect 1612 1573 1626 1587
rect 1653 1573 1667 1587
rect 1713 1573 1727 1587
rect 1913 1593 1927 1607
rect 2013 1593 2027 1607
rect 2253 1593 2267 1607
rect 2473 1593 2487 1607
rect 2693 1593 2707 1607
rect 2773 1593 2787 1607
rect 2874 1593 2888 1607
rect 1973 1573 1987 1587
rect 2133 1573 2147 1587
rect 2213 1573 2227 1587
rect 2293 1573 2307 1587
rect 2393 1573 2407 1587
rect 3033 1592 3047 1606
rect 2933 1573 2947 1587
rect 3053 1573 3067 1587
rect 3092 1573 3106 1587
rect 3134 1573 3148 1587
rect 3513 1613 3527 1627
rect 3753 1613 3767 1627
rect 3793 1613 3807 1627
rect 3873 1613 3887 1627
rect 4033 1613 4047 1627
rect 4213 1612 4227 1626
rect 4253 1613 4267 1627
rect 4313 1613 4327 1627
rect 4393 1613 4407 1627
rect 4453 1613 4467 1627
rect 4533 1613 4547 1627
rect 4773 1613 4787 1627
rect 4833 1613 4847 1627
rect 4952 1613 4966 1627
rect 5133 1613 5147 1627
rect 3973 1593 3987 1607
rect 4193 1593 4207 1607
rect 4792 1593 4806 1607
rect 4974 1593 4988 1607
rect 5033 1593 5047 1607
rect 5293 1633 5307 1647
rect 5613 1633 5627 1647
rect 5673 1633 5687 1647
rect 5333 1613 5347 1627
rect 5393 1613 5407 1627
rect 5633 1613 5647 1627
rect 5713 1613 5727 1627
rect 5193 1593 5207 1607
rect 3413 1573 3427 1587
rect 3473 1573 3487 1587
rect 3833 1573 3847 1587
rect 4133 1573 4147 1587
rect 4214 1573 4228 1587
rect 4314 1573 4328 1587
rect 4453 1573 4467 1587
rect 73 1553 87 1567
rect 113 1552 127 1566
rect 373 1553 387 1567
rect 514 1553 528 1567
rect 693 1553 707 1567
rect 773 1553 787 1567
rect 892 1553 906 1567
rect 914 1553 928 1567
rect 1073 1553 1087 1567
rect 1493 1553 1507 1567
rect 1773 1553 1787 1567
rect 2033 1553 2047 1567
rect 2713 1553 2727 1567
rect 2873 1553 2887 1567
rect 2974 1553 2988 1567
rect 3373 1553 3387 1567
rect 3553 1553 3567 1567
rect 3593 1553 3607 1567
rect 3673 1553 3687 1567
rect 4334 1553 4348 1567
rect 4473 1553 4487 1567
rect 4633 1573 4647 1587
rect 4773 1573 4787 1587
rect 4812 1573 4826 1587
rect 4952 1573 4966 1587
rect 5493 1593 5507 1607
rect 5613 1593 5627 1607
rect 393 1533 407 1547
rect 573 1533 587 1547
rect 1333 1533 1347 1547
rect 1453 1533 1467 1547
rect 1893 1533 1907 1547
rect 2853 1533 2867 1547
rect 3493 1533 3507 1547
rect 4093 1533 4107 1547
rect 4153 1533 4167 1547
rect 4213 1533 4227 1547
rect 4493 1533 4507 1547
rect 4673 1553 4687 1567
rect 4733 1553 4747 1567
rect 5173 1553 5187 1567
rect 5273 1553 5287 1567
rect 4813 1533 4827 1547
rect 5113 1533 5127 1547
rect 5513 1572 5527 1586
rect 5554 1573 5568 1587
rect 5493 1553 5507 1567
rect 5593 1553 5607 1567
rect 5693 1553 5707 1567
rect 1073 1513 1087 1527
rect 1213 1513 1227 1527
rect 1413 1513 1427 1527
rect 1713 1513 1727 1527
rect 2753 1513 2767 1527
rect 2793 1513 2807 1527
rect 4772 1513 4786 1527
rect 4794 1513 4808 1527
rect 5613 1533 5627 1547
rect 5493 1513 5507 1527
rect 5534 1513 5548 1527
rect 5653 1513 5667 1527
rect 73 1493 87 1507
rect 313 1493 327 1507
rect 1573 1493 1587 1507
rect 1853 1493 1867 1507
rect 2053 1493 2067 1507
rect 2313 1493 2327 1507
rect 2713 1493 2727 1507
rect 2873 1493 2887 1507
rect 3213 1493 3227 1507
rect 3333 1493 3347 1507
rect 3533 1493 3547 1507
rect 4153 1493 4167 1507
rect 4273 1493 4287 1507
rect 4433 1493 4447 1507
rect 4673 1493 4687 1507
rect 5133 1493 5147 1507
rect 5273 1493 5287 1507
rect 5573 1493 5587 1507
rect 1473 1473 1487 1487
rect 1973 1473 1987 1487
rect 2213 1473 2227 1487
rect 2993 1473 3007 1487
rect 3133 1473 3147 1487
rect 1113 1453 1127 1467
rect 1213 1453 1227 1467
rect 1793 1453 1807 1467
rect 2553 1453 2567 1467
rect 3113 1453 3127 1467
rect 3153 1453 3167 1467
rect 3393 1453 3407 1467
rect 3793 1473 3807 1487
rect 4313 1473 4327 1487
rect 4393 1473 4407 1487
rect 4713 1473 4727 1487
rect 4933 1473 4947 1487
rect 5053 1473 5067 1487
rect 5153 1473 5167 1487
rect 5312 1473 5326 1487
rect 5334 1473 5348 1487
rect 4353 1453 4367 1467
rect 4653 1453 4667 1467
rect 4953 1453 4967 1467
rect 5233 1453 5247 1467
rect 5633 1473 5647 1487
rect 5693 1473 5707 1487
rect 853 1433 867 1447
rect 1193 1433 1207 1447
rect 1413 1433 1427 1447
rect 2332 1433 2346 1447
rect 2354 1433 2368 1447
rect 2793 1433 2807 1447
rect 3313 1433 3327 1447
rect 3413 1434 3427 1448
rect 3453 1433 3467 1447
rect 3993 1433 4007 1447
rect 4033 1433 4047 1447
rect 4173 1433 4187 1447
rect 4273 1433 4287 1447
rect 4333 1433 4347 1447
rect 4593 1434 4607 1448
rect 4693 1433 4707 1447
rect 4913 1433 4927 1447
rect 5113 1433 5127 1447
rect 5313 1433 5327 1447
rect 5453 1453 5467 1467
rect 5413 1433 5427 1447
rect 5553 1433 5567 1447
rect 693 1413 707 1427
rect 913 1413 927 1427
rect 1232 1413 1246 1427
rect 1533 1413 1547 1427
rect 2393 1413 2407 1427
rect 2473 1413 2487 1427
rect 2933 1413 2947 1427
rect 3413 1412 3427 1426
rect 3633 1413 3647 1427
rect 4093 1413 4107 1427
rect 4373 1413 4387 1427
rect 4593 1412 4607 1426
rect 4852 1413 4866 1427
rect 4933 1413 4947 1427
rect 5013 1413 5027 1427
rect 5273 1413 5287 1427
rect 5393 1414 5407 1428
rect 5613 1413 5627 1427
rect 633 1393 647 1407
rect 933 1393 947 1407
rect 1273 1393 1287 1407
rect 1513 1393 1527 1407
rect 2333 1393 2347 1407
rect 2433 1393 2447 1407
rect 4133 1393 4147 1407
rect 4473 1393 4487 1407
rect 4953 1393 4967 1407
rect 5113 1393 5127 1407
rect 5393 1392 5407 1406
rect 5433 1393 5447 1407
rect 5513 1393 5527 1407
rect 5713 1393 5727 1407
rect 233 1373 247 1387
rect 573 1373 587 1387
rect 1013 1373 1027 1387
rect 1733 1373 1747 1387
rect 1833 1373 1847 1387
rect 2393 1373 2407 1387
rect 2613 1373 2627 1387
rect 2953 1373 2967 1387
rect 3953 1373 3967 1387
rect 4013 1373 4027 1387
rect 4633 1373 4647 1387
rect 4793 1373 4807 1387
rect 4893 1373 4907 1387
rect 5173 1373 5187 1387
rect 5493 1373 5507 1387
rect 312 1353 326 1367
rect 334 1353 348 1367
rect 513 1353 527 1367
rect 793 1353 807 1367
rect 1173 1353 1187 1367
rect 192 1333 206 1347
rect 273 1333 287 1347
rect 493 1333 507 1347
rect 633 1333 647 1347
rect 993 1333 1007 1347
rect 1213 1353 1227 1367
rect 2113 1353 2127 1367
rect 2213 1353 2227 1367
rect 2453 1353 2467 1367
rect 1273 1333 1287 1347
rect 1413 1333 1427 1347
rect 1533 1333 1547 1347
rect 1753 1333 1767 1347
rect 2073 1333 2087 1347
rect 2273 1333 2287 1347
rect 2353 1334 2367 1348
rect 3033 1353 3047 1367
rect 3193 1353 3207 1367
rect 3273 1353 3287 1367
rect 3613 1353 3627 1367
rect 3893 1353 3907 1367
rect 3973 1353 3987 1367
rect 4273 1353 4287 1367
rect 4833 1353 4847 1367
rect 4873 1353 4887 1367
rect 4973 1353 4987 1367
rect 5073 1353 5087 1367
rect 5253 1353 5267 1367
rect 5453 1353 5467 1367
rect 5553 1353 5567 1367
rect 2434 1333 2448 1347
rect 2893 1333 2907 1347
rect 2933 1333 2947 1347
rect 4133 1333 4147 1347
rect 4233 1333 4247 1347
rect 4353 1333 4367 1347
rect 4453 1333 4467 1347
rect 4633 1333 4647 1347
rect 5013 1333 5027 1347
rect 253 1313 267 1327
rect 313 1313 327 1327
rect 354 1313 368 1327
rect 433 1313 447 1327
rect 534 1313 548 1327
rect 792 1313 806 1327
rect 833 1313 847 1327
rect 873 1313 887 1327
rect 933 1313 947 1327
rect 1172 1313 1186 1327
rect 1212 1313 1226 1327
rect 1234 1313 1248 1327
rect 1513 1313 1527 1327
rect 1633 1313 1647 1327
rect 1793 1313 1807 1327
rect 112 1293 126 1307
rect 153 1293 167 1307
rect 672 1293 686 1307
rect 753 1293 767 1307
rect 853 1293 867 1307
rect 2014 1313 2028 1327
rect 2353 1312 2367 1326
rect 2413 1313 2427 1327
rect 2473 1313 2487 1327
rect 1133 1293 1147 1307
rect 93 1273 107 1287
rect 633 1273 647 1287
rect 1693 1292 1707 1306
rect 213 1253 227 1267
rect 553 1253 567 1267
rect 1073 1273 1087 1287
rect 1754 1273 1768 1287
rect 2313 1293 2327 1307
rect 2513 1293 2527 1307
rect 2613 1313 2627 1327
rect 2653 1313 2667 1327
rect 2752 1313 2766 1327
rect 3013 1313 3027 1327
rect 3152 1313 3166 1327
rect 3193 1313 3207 1327
rect 2953 1293 2967 1307
rect 3053 1293 3067 1307
rect 3093 1293 3107 1307
rect 2073 1273 2087 1287
rect 2173 1273 2187 1287
rect 2233 1273 2247 1287
rect 1033 1253 1047 1267
rect 1233 1253 1247 1267
rect 1673 1253 1687 1267
rect 1933 1253 1947 1267
rect 2233 1253 2247 1267
rect 2493 1253 2507 1267
rect 2793 1273 2807 1287
rect 3792 1313 3806 1327
rect 3913 1313 3927 1327
rect 4213 1313 4227 1327
rect 4473 1313 4487 1327
rect 4713 1313 4727 1327
rect 4792 1314 4806 1328
rect 4833 1313 4847 1327
rect 4953 1313 4967 1327
rect 3432 1293 3446 1307
rect 3693 1293 3707 1307
rect 3853 1293 3867 1307
rect 3973 1293 3987 1307
rect 4133 1293 4147 1307
rect 4273 1293 4287 1307
rect 4413 1293 4427 1307
rect 4593 1293 4607 1307
rect 4634 1293 4648 1307
rect 5413 1333 5427 1347
rect 4813 1293 4827 1307
rect 4893 1293 4907 1307
rect 4933 1293 4947 1307
rect 5152 1293 5166 1307
rect 5194 1293 5208 1307
rect 5313 1293 5327 1307
rect 5454 1313 5468 1327
rect 5373 1293 5387 1307
rect 5414 1293 5428 1307
rect 3233 1273 3247 1287
rect 3313 1273 3327 1287
rect 3393 1273 3407 1287
rect 3753 1273 3767 1287
rect 4313 1273 4327 1287
rect 4373 1273 4387 1287
rect 4532 1273 4546 1287
rect 4554 1273 4568 1287
rect 4613 1273 4627 1287
rect 4653 1273 4667 1287
rect 4833 1273 4847 1287
rect 5133 1273 5147 1287
rect 2853 1253 2867 1267
rect 3053 1253 3067 1267
rect 3693 1253 3707 1267
rect 4033 1253 4047 1267
rect 4573 1254 4587 1268
rect 4913 1253 4927 1267
rect 5013 1254 5027 1268
rect 5093 1253 5107 1267
rect 5193 1253 5207 1267
rect 5293 1253 5307 1267
rect 5653 1273 5667 1287
rect 5473 1253 5487 1267
rect 33 1233 47 1247
rect 353 1233 367 1247
rect 893 1233 907 1247
rect 1073 1233 1087 1247
rect 1733 1233 1747 1247
rect 1792 1233 1806 1247
rect 2253 1233 2267 1247
rect 2293 1233 2307 1247
rect 2372 1233 2386 1247
rect 2394 1233 2408 1247
rect 2653 1233 2667 1247
rect 2753 1233 2767 1247
rect 2953 1233 2967 1247
rect 3913 1233 3927 1247
rect 4573 1232 4587 1246
rect 4753 1233 4767 1247
rect 4893 1233 4907 1247
rect 5013 1232 5027 1246
rect 5633 1233 5647 1247
rect 5673 1233 5687 1247
rect 673 1213 687 1227
rect 832 1213 846 1227
rect 854 1213 868 1227
rect 1213 1213 1227 1227
rect 1293 1213 1307 1227
rect 1973 1213 1987 1227
rect 2353 1213 2367 1227
rect 2553 1213 2567 1227
rect 2713 1213 2727 1227
rect 93 1193 107 1207
rect 553 1193 567 1207
rect 1253 1193 1267 1207
rect 1573 1194 1587 1208
rect 3373 1213 3387 1227
rect 3453 1214 3467 1228
rect 2333 1193 2347 1207
rect 2753 1193 2767 1207
rect 2893 1193 2907 1207
rect 3113 1193 3127 1207
rect 3313 1193 3327 1207
rect 113 1173 127 1187
rect 433 1173 447 1187
rect 753 1173 767 1187
rect 1133 1173 1147 1187
rect 1373 1173 1387 1187
rect 1573 1172 1587 1186
rect 1853 1173 1867 1187
rect 2293 1173 2307 1187
rect 2353 1173 2367 1187
rect 3213 1173 3227 1187
rect 3333 1173 3347 1187
rect 3453 1192 3467 1206
rect 3513 1193 3527 1207
rect 3713 1213 3727 1227
rect 4213 1213 4227 1227
rect 4613 1213 4627 1227
rect 4933 1213 4947 1227
rect 4993 1213 5007 1227
rect 5233 1213 5247 1227
rect 5333 1213 5347 1227
rect 5513 1213 5527 1227
rect 3753 1193 3767 1207
rect 4953 1193 4967 1207
rect 5313 1193 5327 1207
rect 5593 1193 5607 1207
rect 5693 1193 5707 1207
rect 3473 1173 3487 1187
rect 4673 1173 4687 1187
rect 4853 1173 4867 1187
rect 5133 1173 5147 1187
rect 5573 1173 5587 1187
rect 5653 1173 5667 1187
rect 93 1153 107 1167
rect 173 1153 187 1167
rect 293 1153 307 1167
rect 673 1153 687 1167
rect 793 1153 807 1167
rect 933 1153 947 1167
rect 993 1153 1007 1167
rect 1193 1153 1207 1167
rect 1353 1153 1367 1167
rect 1673 1153 1687 1167
rect 1813 1153 1827 1167
rect 2513 1153 2527 1167
rect 2793 1153 2807 1167
rect 3033 1153 3047 1167
rect 3273 1153 3287 1167
rect 3513 1153 3527 1167
rect 3613 1153 3627 1167
rect 4293 1153 4307 1167
rect 4533 1153 4547 1167
rect 4993 1153 5007 1167
rect 5093 1153 5107 1167
rect 5153 1153 5167 1167
rect 5253 1153 5267 1167
rect 93 1133 107 1147
rect 133 1133 147 1147
rect 493 1133 507 1147
rect 613 1133 627 1147
rect 273 1113 287 1127
rect 433 1113 447 1127
rect 33 1093 47 1107
rect 733 1113 747 1127
rect 1013 1133 1027 1147
rect 1353 1133 1367 1147
rect 1453 1133 1467 1147
rect 1693 1133 1707 1147
rect 1793 1133 1807 1147
rect 1853 1133 1867 1147
rect 2293 1133 2307 1147
rect 2413 1133 2427 1147
rect 2833 1133 2847 1147
rect 3013 1133 3027 1147
rect 3093 1133 3107 1147
rect 3312 1133 3326 1147
rect 3334 1133 3348 1147
rect 3993 1133 4007 1147
rect 4033 1133 4047 1147
rect 4353 1133 4367 1147
rect 4593 1133 4607 1147
rect 4653 1133 4667 1147
rect 4873 1133 4887 1147
rect 5013 1133 5027 1147
rect 5173 1133 5187 1147
rect 5313 1133 5327 1147
rect 5413 1133 5427 1147
rect 5553 1153 5567 1167
rect 5533 1133 5547 1147
rect 5573 1133 5587 1147
rect 933 1113 947 1127
rect 1033 1113 1047 1127
rect 1074 1113 1088 1127
rect 1114 1113 1128 1127
rect 173 1093 187 1107
rect 294 1093 308 1107
rect 232 1073 246 1087
rect 313 1073 327 1087
rect 593 1093 607 1107
rect 673 1093 687 1107
rect 853 1093 867 1107
rect 553 1073 567 1087
rect 793 1073 807 1087
rect 893 1073 907 1087
rect 1173 1093 1187 1107
rect 1214 1093 1228 1107
rect 1313 1093 1327 1107
rect 1713 1113 1727 1127
rect 1933 1113 1947 1127
rect 1973 1113 1987 1127
rect 2133 1113 2147 1127
rect 2233 1113 2247 1127
rect 2333 1113 2347 1127
rect 2473 1113 2487 1127
rect 2713 1113 2727 1127
rect 2853 1113 2867 1127
rect 3113 1113 3127 1127
rect 3312 1113 3326 1127
rect 3613 1113 3627 1127
rect 3733 1113 3747 1127
rect 3853 1113 3867 1127
rect 3974 1113 3988 1127
rect 4093 1113 4107 1127
rect 1153 1073 1167 1087
rect 1293 1073 1307 1087
rect 1373 1073 1387 1087
rect 1453 1073 1467 1087
rect 1592 1073 1606 1087
rect 1793 1073 1807 1087
rect 2033 1093 2047 1107
rect 2292 1093 2306 1107
rect 2393 1093 2407 1107
rect 2493 1093 2507 1107
rect 2554 1093 2568 1107
rect 2613 1093 2627 1107
rect 2173 1073 2187 1087
rect 2233 1073 2247 1087
rect 2753 1093 2767 1107
rect 2873 1093 2887 1107
rect 3013 1093 3027 1107
rect 3073 1073 3087 1087
rect 3153 1073 3167 1087
rect 3433 1093 3447 1107
rect 3494 1093 3508 1107
rect 3193 1073 3207 1087
rect 3293 1073 3307 1087
rect 3753 1092 3767 1106
rect 4133 1093 4147 1107
rect 4213 1093 4227 1107
rect 4333 1093 4347 1107
rect 4973 1113 4987 1127
rect 5113 1113 5127 1127
rect 5373 1113 5387 1127
rect 5473 1113 5487 1127
rect 5613 1113 5627 1127
rect 4553 1093 4567 1107
rect 4634 1093 4648 1107
rect 4873 1093 4887 1107
rect 5133 1093 5147 1107
rect 5213 1093 5227 1107
rect 5253 1093 5267 1107
rect 5513 1093 5527 1107
rect 3653 1073 3667 1087
rect 3973 1073 3987 1087
rect 4073 1073 4087 1087
rect 4193 1073 4207 1087
rect 4233 1073 4247 1087
rect 4274 1073 4288 1087
rect 4313 1073 4327 1087
rect 4593 1073 4607 1087
rect 4693 1073 4707 1087
rect 4833 1073 4847 1087
rect 5113 1073 5127 1087
rect 5273 1073 5287 1087
rect 5593 1073 5607 1087
rect 673 1053 687 1067
rect 973 1053 987 1067
rect 1013 1053 1027 1067
rect 1313 1053 1327 1067
rect 1553 1053 1567 1067
rect 2033 1053 2047 1067
rect 3053 1053 3067 1067
rect 3193 1053 3207 1067
rect 4273 1053 4287 1067
rect 4713 1053 4727 1067
rect 5193 1053 5207 1067
rect 5313 1053 5327 1067
rect 5433 1053 5447 1067
rect 1113 1033 1127 1047
rect 1593 1033 1607 1047
rect 2693 1033 2707 1047
rect 2733 1033 2747 1047
rect 2853 1033 2867 1047
rect 3073 1033 3087 1047
rect 4173 1033 4187 1047
rect 4233 1033 4247 1047
rect 4313 1033 4327 1047
rect 4473 1033 4487 1047
rect 4873 1033 4887 1047
rect 4993 1033 5007 1047
rect 5033 1033 5047 1047
rect 5453 1033 5467 1047
rect 273 1013 287 1027
rect 1213 1013 1227 1027
rect 1373 1013 1387 1027
rect 2213 1013 2227 1027
rect 3333 1013 3347 1027
rect 5013 1013 5027 1027
rect 5073 1013 5087 1027
rect 5553 1013 5567 1027
rect 1833 993 1847 1007
rect 2433 993 2447 1007
rect 2593 993 2607 1007
rect 2733 993 2747 1007
rect 3613 993 3627 1007
rect 3652 993 3666 1007
rect 3674 993 3688 1007
rect 4033 993 4047 1007
rect 4493 993 4507 1007
rect 5113 993 5127 1007
rect 5593 994 5607 1008
rect 3753 973 3767 987
rect 4073 973 4087 987
rect 4153 973 4167 987
rect 4313 973 4327 987
rect 4373 973 4387 987
rect 4993 973 5007 987
rect 5093 973 5107 987
rect 5493 973 5507 987
rect 5533 973 5547 987
rect 5593 972 5607 986
rect 2653 953 2667 967
rect 3173 953 3187 967
rect 3793 953 3807 967
rect 4033 953 4047 967
rect 4333 953 4347 967
rect 4413 953 4427 967
rect 4793 953 4807 967
rect 4833 953 4847 967
rect 5133 953 5147 967
rect 373 933 387 947
rect 1013 933 1027 947
rect 1153 933 1167 947
rect 1553 933 1567 947
rect 3233 933 3247 947
rect 3553 933 3567 947
rect 3833 933 3847 947
rect 4113 933 4127 947
rect 4373 933 4387 947
rect 4673 933 4687 947
rect 5293 933 5307 947
rect 5393 933 5407 947
rect 5473 933 5487 947
rect 5553 933 5567 947
rect 5633 933 5647 947
rect 333 913 347 927
rect 593 913 607 927
rect 693 913 707 927
rect 1313 913 1327 927
rect 1833 913 1847 927
rect 1993 913 2007 927
rect 2313 913 2327 927
rect 2633 913 2647 927
rect 3273 913 3287 927
rect 3533 913 3547 927
rect 3733 913 3747 927
rect 4093 913 4107 927
rect 4173 913 4187 927
rect 4513 913 4527 927
rect 4813 913 4827 927
rect 4853 913 4867 927
rect 4973 913 4987 927
rect 5053 913 5067 927
rect 5173 913 5187 927
rect 5233 913 5247 927
rect 5693 913 5707 927
rect 93 893 107 907
rect 253 893 267 907
rect 713 893 727 907
rect 1813 893 1827 907
rect 2053 893 2067 907
rect 2853 893 2867 907
rect 3113 893 3127 907
rect 3153 893 3167 907
rect 3913 893 3927 907
rect 153 873 167 887
rect 233 873 247 887
rect 193 853 207 867
rect 333 853 347 867
rect 373 853 387 867
rect 153 833 167 847
rect 233 833 247 847
rect 413 833 427 847
rect 454 833 468 847
rect 612 834 626 848
rect 1193 873 1207 887
rect 1573 873 1587 887
rect 1693 873 1707 887
rect 1873 873 1887 887
rect 2013 873 2027 887
rect 2273 873 2287 887
rect 753 853 767 867
rect 853 853 867 867
rect 1313 853 1327 867
rect 1353 853 1367 867
rect 1633 853 1647 867
rect 1773 853 1787 867
rect 1913 853 1927 867
rect 1993 853 2007 867
rect 2873 873 2887 887
rect 2913 874 2927 888
rect 4733 893 4747 907
rect 4793 893 4807 907
rect 4874 893 4888 907
rect 5033 893 5047 907
rect 5193 893 5207 907
rect 5273 893 5287 907
rect 5333 893 5347 907
rect 5393 893 5407 907
rect 5433 893 5447 907
rect 2973 873 2987 887
rect 3092 873 3106 887
rect 3993 873 4007 887
rect 2473 853 2487 867
rect 2573 853 2587 867
rect 692 833 706 847
rect 813 833 827 847
rect 573 813 587 827
rect 632 813 646 827
rect 933 833 947 847
rect 1252 833 1266 847
rect 1452 833 1466 847
rect 1493 833 1507 847
rect 1953 833 1967 847
rect 2033 833 2047 847
rect 2213 833 2227 847
rect 2313 833 2327 847
rect 2533 834 2547 848
rect 2633 853 2647 867
rect 2813 853 2827 867
rect 2913 852 2927 866
rect 3114 853 3128 867
rect 3292 853 3306 867
rect 3314 853 3328 867
rect 3373 853 3387 867
rect 3413 853 3427 867
rect 2614 833 2628 847
rect 2773 833 2787 847
rect 2873 833 2887 847
rect 3013 833 3027 847
rect 3053 833 3067 847
rect 3173 833 3187 847
rect 3252 833 3266 847
rect 3492 834 3506 848
rect 3573 853 3587 867
rect 3693 853 3707 867
rect 3873 853 3887 867
rect 4033 873 4047 887
rect 4113 873 4127 887
rect 4233 873 4247 887
rect 4953 873 4967 887
rect 4173 853 4187 867
rect 4773 853 4787 867
rect 4913 853 4927 867
rect 5173 873 5187 887
rect 5233 873 5247 887
rect 5353 873 5367 887
rect 5473 873 5487 887
rect 5533 873 5547 887
rect 5293 853 5307 867
rect 5353 853 5367 867
rect 3592 833 3606 847
rect 3913 833 3927 847
rect 4053 833 4067 847
rect 4193 833 4207 847
rect 4232 833 4246 847
rect 4353 833 4367 847
rect 4393 833 4407 847
rect 4453 833 4467 847
rect 4494 833 4508 847
rect 973 813 987 827
rect 1052 813 1066 827
rect 1132 813 1146 827
rect 1213 813 1227 827
rect 1272 813 1286 827
rect 1573 813 1587 827
rect 1633 813 1647 827
rect 1693 813 1707 827
rect 1753 813 1767 827
rect 1872 813 1886 827
rect 1913 813 1927 827
rect 2093 813 2107 827
rect 2273 813 2287 827
rect 2413 813 2427 827
rect 2513 813 2527 827
rect 2653 813 2667 827
rect 2993 813 3007 827
rect 3153 813 3167 827
rect 3433 813 3447 827
rect 3512 813 3526 827
rect 3793 813 3807 827
rect 3953 813 3967 827
rect 113 793 127 807
rect 173 793 187 807
rect 233 793 247 807
rect 433 793 447 807
rect 213 773 227 787
rect 693 773 707 787
rect 1313 793 1327 807
rect 1513 793 1527 807
rect 1813 793 1827 807
rect 2133 793 2147 807
rect 2573 793 2587 807
rect 2813 793 2827 807
rect 3352 793 3366 807
rect 3374 793 3388 807
rect 3453 793 3467 807
rect 4033 793 4047 807
rect 4792 832 4806 846
rect 4833 833 4847 847
rect 4992 833 5006 847
rect 5173 833 5187 847
rect 5433 853 5447 867
rect 5593 853 5607 867
rect 5473 833 5487 847
rect 5673 833 5687 847
rect 4293 813 4307 827
rect 4693 813 4707 827
rect 5153 813 5167 827
rect 5394 813 5408 827
rect 5434 813 5448 827
rect 5534 813 5548 827
rect 5632 813 5646 827
rect 4153 793 4167 807
rect 4353 793 4367 807
rect 4412 793 4426 807
rect 4633 793 4647 807
rect 4993 793 5007 807
rect 5353 793 5367 807
rect 5493 793 5507 807
rect 1273 773 1287 787
rect 1593 773 1607 787
rect 1793 773 1807 787
rect 1953 773 1967 787
rect 2213 773 2227 787
rect 2433 773 2447 787
rect 2673 773 2687 787
rect 2733 773 2747 787
rect 2833 773 2847 787
rect 2993 773 3007 787
rect 3553 773 3567 787
rect 4453 773 4467 787
rect 4593 773 4607 787
rect 5153 773 5167 787
rect 173 753 187 767
rect 453 753 467 767
rect 613 753 627 767
rect 733 753 747 767
rect 813 753 827 767
rect 853 753 867 767
rect 932 753 946 767
rect 1053 753 1067 767
rect 1153 753 1167 767
rect 1493 753 1507 767
rect 1973 753 1987 767
rect 2033 753 2047 767
rect 2533 753 2547 767
rect 2793 753 2807 767
rect 2913 753 2927 767
rect 3213 753 3227 767
rect 3453 753 3467 767
rect 3513 753 3527 767
rect 3873 753 3887 767
rect 4893 753 4907 767
rect 4993 753 5007 767
rect 5613 753 5627 767
rect 353 733 367 747
rect 493 733 507 747
rect 1553 733 1567 747
rect 913 713 927 727
rect 1013 713 1027 727
rect 1313 713 1327 727
rect 1933 733 1947 747
rect 2053 733 2067 747
rect 2573 733 2587 747
rect 3153 733 3167 747
rect 3233 733 3247 747
rect 3313 733 3327 747
rect 3353 733 3367 747
rect 3493 733 3507 747
rect 3953 733 3967 747
rect 4433 733 4447 747
rect 4473 733 4487 747
rect 4533 733 4547 747
rect 4933 733 4947 747
rect 5413 733 5427 747
rect 2733 713 2747 727
rect 2773 713 2787 727
rect 3413 713 3427 727
rect 3933 713 3947 727
rect 3993 713 4007 727
rect 4373 713 4387 727
rect 4753 713 4767 727
rect 4873 713 4887 727
rect 5273 713 5287 727
rect 5333 713 5347 727
rect 5653 713 5667 727
rect 93 693 107 707
rect 333 693 347 707
rect 753 693 767 707
rect 993 693 1007 707
rect 1233 693 1247 707
rect 1453 693 1467 707
rect 1633 693 1647 707
rect 1753 693 1767 707
rect 2153 693 2167 707
rect 2213 693 2227 707
rect 2613 693 2627 707
rect 2653 693 2667 707
rect 2693 693 2707 707
rect 3013 693 3027 707
rect 3333 693 3347 707
rect 3393 693 3407 707
rect 3833 693 3847 707
rect 4173 693 4187 707
rect 4273 693 4287 707
rect 4513 693 4527 707
rect 4673 693 4687 707
rect 4793 693 4807 707
rect 4853 693 4867 707
rect 5033 693 5047 707
rect 5313 693 5327 707
rect 5393 693 5407 707
rect 93 673 107 687
rect 313 673 327 687
rect 593 673 607 687
rect 1073 673 1087 687
rect 1133 673 1147 687
rect 1213 673 1227 687
rect 1593 673 1607 687
rect 1833 673 1847 687
rect 2433 673 2447 687
rect 2973 673 2987 687
rect 3273 673 3287 687
rect 3593 673 3607 687
rect 3973 673 3987 687
rect 193 653 207 667
rect 253 653 267 667
rect 753 653 767 667
rect 1073 653 1087 667
rect 1353 653 1367 667
rect 1533 653 1547 667
rect 2153 653 2167 667
rect 2373 653 2387 667
rect 2453 653 2467 667
rect 2673 653 2687 667
rect 373 633 387 647
rect 593 633 607 647
rect 173 613 187 627
rect 233 613 247 627
rect 352 614 366 628
rect 673 633 687 647
rect 1253 633 1267 647
rect 1493 633 1507 647
rect 1553 633 1567 647
rect 1592 633 1606 647
rect 1752 633 1766 647
rect 1833 633 1847 647
rect 1933 633 1947 647
rect 493 613 507 627
rect 634 613 648 627
rect 733 613 747 627
rect 853 613 867 627
rect 994 613 1008 627
rect 1172 613 1186 627
rect 1213 613 1227 627
rect 1533 613 1547 627
rect 1653 613 1667 627
rect 1793 613 1807 627
rect 373 593 387 607
rect 693 593 707 607
rect 193 573 207 587
rect 313 573 327 587
rect 633 573 647 587
rect 1293 593 1307 607
rect 1493 593 1507 607
rect 1973 633 1987 647
rect 2293 633 2307 647
rect 2353 633 2367 647
rect 2473 634 2487 648
rect 2713 634 2727 648
rect 2913 653 2927 667
rect 2953 633 2967 647
rect 3213 653 3227 667
rect 3333 653 3347 667
rect 3473 653 3487 667
rect 3553 653 3567 667
rect 3673 653 3687 667
rect 3733 653 3747 667
rect 3054 633 3068 647
rect 3493 633 3507 647
rect 3593 633 3607 647
rect 3953 653 3967 667
rect 4313 674 4327 688
rect 4593 673 4607 687
rect 5133 673 5147 687
rect 5553 673 5567 687
rect 4272 653 4286 667
rect 4313 652 4327 666
rect 4434 653 4448 667
rect 4513 653 4527 667
rect 2173 613 2187 627
rect 2392 613 2406 627
rect 2113 593 2127 607
rect 2473 612 2487 626
rect 2593 613 2607 627
rect 2713 612 2727 626
rect 2993 613 3007 627
rect 3133 613 3147 627
rect 3214 613 3228 627
rect 3432 613 3446 627
rect 3454 613 3468 627
rect 3633 613 3647 627
rect 3993 633 4007 647
rect 4153 633 4167 647
rect 4412 633 4426 647
rect 3953 613 3967 627
rect 4053 613 4067 627
rect 4213 613 4227 627
rect 4633 633 4647 647
rect 4713 633 4727 647
rect 5193 653 5207 667
rect 5393 653 5407 667
rect 5452 653 5466 667
rect 5474 653 5488 667
rect 5032 633 5046 647
rect 5073 633 5087 647
rect 5273 634 5287 648
rect 5373 633 5387 647
rect 4653 613 4667 627
rect 4753 613 4767 627
rect 4834 613 4848 627
rect 4953 613 4967 627
rect 4993 613 5007 627
rect 5133 613 5147 627
rect 5173 613 5187 627
rect 2413 593 2427 607
rect 2652 593 2666 607
rect 2674 593 2688 607
rect 2913 593 2927 607
rect 2954 593 2968 607
rect 3073 593 3087 607
rect 3572 593 3586 607
rect 3594 593 3608 607
rect 3653 593 3667 607
rect 4313 593 4327 607
rect 4513 593 4527 607
rect 4812 593 4826 607
rect 5273 612 5287 626
rect 853 573 867 587
rect 2173 573 2187 587
rect 2393 573 2407 587
rect 2653 573 2667 587
rect 2713 573 2727 587
rect 3573 573 3587 587
rect 3673 573 3687 587
rect 4853 573 4867 587
rect 5234 593 5248 607
rect 5533 593 5547 607
rect 5212 573 5226 587
rect 5234 573 5248 587
rect 273 553 287 567
rect 353 553 367 567
rect 553 553 567 567
rect 1053 553 1067 567
rect 1653 553 1667 567
rect 2613 553 2627 567
rect 2833 553 2847 567
rect 4013 553 4027 567
rect 5033 553 5047 567
rect 5373 553 5387 567
rect 5673 553 5687 567
rect 613 533 627 547
rect 1093 533 1107 547
rect 1133 533 1147 547
rect 173 513 187 527
rect 1473 533 1487 547
rect 2393 533 2407 547
rect 4813 533 4827 547
rect 5293 533 5307 547
rect 3013 513 3027 527
rect 4553 513 4567 527
rect 4913 513 4927 527
rect 5353 513 5367 527
rect 793 493 807 507
rect 1293 493 1307 507
rect 1833 493 1847 507
rect 3092 493 3106 507
rect 3114 493 3128 507
rect 3233 493 3247 507
rect 4593 493 4607 507
rect 4993 493 5007 507
rect 5073 493 5087 507
rect 5153 493 5167 507
rect 5213 493 5227 507
rect 5533 493 5547 507
rect 893 473 907 487
rect 1193 473 1207 487
rect 2173 473 2187 487
rect 2873 473 2887 487
rect 3793 473 3807 487
rect 4673 473 4687 487
rect 5233 473 5247 487
rect 633 453 647 467
rect 673 453 687 467
rect 1253 453 1267 467
rect 1513 453 1527 467
rect 2273 453 2287 467
rect 3072 453 3086 467
rect 3094 453 3108 467
rect 3633 453 3647 467
rect 3753 453 3767 467
rect 3893 453 3907 467
rect 4473 453 4487 467
rect 4653 453 4667 467
rect 4713 453 4727 467
rect 4813 453 4827 467
rect 5473 453 5487 467
rect 213 433 227 447
rect 732 433 746 447
rect 2033 433 2047 447
rect 2113 433 2127 447
rect 2193 433 2207 447
rect 2233 433 2247 447
rect 4173 433 4187 447
rect 4553 433 4567 447
rect 4633 433 4647 447
rect 4973 433 4987 447
rect 5413 433 5427 447
rect 253 413 267 427
rect 693 413 707 427
rect 833 413 847 427
rect 2432 413 2446 427
rect 2454 413 2468 427
rect 2693 413 2707 427
rect 3713 413 3727 427
rect 3893 413 3907 427
rect 533 393 547 407
rect 173 373 187 387
rect 473 373 487 387
rect 793 373 807 387
rect 1093 393 1107 407
rect 1132 393 1146 407
rect 1253 393 1267 407
rect 1473 393 1487 407
rect 1633 393 1647 407
rect 1053 373 1067 387
rect 93 333 107 347
rect 214 353 228 367
rect 313 353 327 367
rect 413 353 427 367
rect 573 353 587 367
rect 674 353 688 367
rect 253 333 267 347
rect 353 333 367 347
rect 853 353 867 367
rect 1013 353 1027 367
rect 654 333 668 347
rect 734 333 748 347
rect 893 333 907 347
rect 1093 373 1107 387
rect 1293 373 1307 387
rect 1353 373 1367 387
rect 2033 393 2047 407
rect 2233 393 2247 407
rect 2394 393 2408 407
rect 2913 393 2927 407
rect 3413 393 3427 407
rect 3453 393 3467 407
rect 4213 393 4227 407
rect 4753 413 4767 427
rect 5033 413 5047 427
rect 5093 413 5107 427
rect 5633 413 5647 427
rect 4592 393 4606 407
rect 4753 393 4767 407
rect 4913 393 4927 407
rect 4953 393 4967 407
rect 4993 393 5007 407
rect 1813 373 1827 387
rect 1853 373 1867 387
rect 1193 353 1207 367
rect 1273 353 1287 367
rect 2113 373 2127 387
rect 2372 373 2386 387
rect 2493 373 2507 387
rect 2553 373 2567 387
rect 2713 373 2727 387
rect 2793 373 2807 387
rect 3473 373 3487 387
rect 3793 373 3807 387
rect 4013 373 4027 387
rect 4173 373 4187 387
rect 4312 373 4326 387
rect 4354 373 4368 387
rect 4433 373 4447 387
rect 4553 373 4567 387
rect 4614 373 4628 387
rect 5153 393 5167 407
rect 5313 393 5327 407
rect 5673 393 5687 407
rect 5053 373 5067 387
rect 5233 373 5247 387
rect 5393 373 5407 387
rect 1532 353 1546 367
rect 1673 353 1687 367
rect 1833 353 1847 367
rect 1953 353 1967 367
rect 1213 333 1227 347
rect 1413 333 1427 347
rect 1473 333 1487 347
rect 93 313 107 327
rect 213 313 227 327
rect 533 313 547 327
rect 632 313 646 327
rect 993 313 1007 327
rect 1413 313 1427 327
rect 1813 333 1827 347
rect 2433 353 2447 367
rect 2613 353 2627 367
rect 2754 353 2768 367
rect 2913 353 2927 367
rect 2952 353 2966 367
rect 3413 353 3427 367
rect 3833 353 3847 367
rect 3913 353 3927 367
rect 4472 353 4486 367
rect 4533 353 4547 367
rect 4693 353 4707 367
rect 4813 353 4827 367
rect 2713 333 2727 347
rect 2813 333 2827 347
rect 3012 333 3026 347
rect 3034 333 3048 347
rect 3113 333 3127 347
rect 3154 333 3168 347
rect 3513 333 3527 347
rect 3593 333 3607 347
rect 3633 333 3647 347
rect 3693 333 3707 347
rect 3953 333 3967 347
rect 4173 333 4187 347
rect 4833 333 4847 347
rect 5152 353 5166 367
rect 5194 353 5208 367
rect 5294 353 5308 367
rect 5433 373 5447 387
rect 5533 373 5547 387
rect 5593 373 5607 387
rect 5633 353 5647 367
rect 1693 313 1707 327
rect 453 293 467 307
rect 793 293 807 307
rect 2033 313 2047 327
rect 2693 313 2707 327
rect 1913 293 1927 307
rect 2073 293 2087 307
rect 3053 313 3067 327
rect 3233 313 3247 327
rect 3453 313 3467 327
rect 3753 313 3767 327
rect 4033 313 4047 327
rect 5013 313 5027 327
rect 5053 313 5067 327
rect 5093 313 5107 327
rect 5393 313 5407 327
rect 5433 313 5447 327
rect 5673 313 5687 327
rect 4613 293 4627 307
rect 4673 293 4687 307
rect 5453 293 5467 307
rect 5593 294 5607 308
rect 173 273 187 287
rect 393 273 407 287
rect 613 273 627 287
rect 693 273 707 287
rect 1333 273 1347 287
rect 2114 273 2128 287
rect 2573 273 2587 287
rect 2813 273 2827 287
rect 3033 273 3047 287
rect 4553 273 4567 287
rect 4833 273 4847 287
rect 5113 273 5127 287
rect 5593 272 5607 286
rect 513 253 527 267
rect 1693 253 1707 267
rect 2153 253 2167 267
rect 2473 253 2487 267
rect 2953 253 2967 267
rect 3173 253 3187 267
rect 4433 253 4447 267
rect 4793 253 4807 267
rect 5093 253 5107 267
rect 5173 253 5187 267
rect 5713 253 5727 267
rect 853 233 867 247
rect 913 233 927 247
rect 1853 233 1867 247
rect 1973 233 1987 247
rect 2233 233 2247 247
rect 2273 233 2287 247
rect 3133 233 3147 247
rect 4653 233 4667 247
rect 5273 233 5287 247
rect 5393 233 5407 247
rect 5453 233 5467 247
rect 1153 213 1167 227
rect 1213 213 1227 227
rect 1433 213 1447 227
rect 1653 213 1667 227
rect 2393 213 2407 227
rect 2773 213 2787 227
rect 5373 213 5387 227
rect 313 193 327 207
rect 513 193 527 207
rect 1413 193 1427 207
rect 1453 193 1467 207
rect 1473 193 1487 207
rect 1952 193 1966 207
rect 1974 193 1988 207
rect 2013 193 2027 207
rect 2153 193 2167 207
rect 2213 193 2227 207
rect 2493 193 2507 207
rect 3393 193 3407 207
rect 4953 193 4967 207
rect 5313 193 5327 207
rect 5553 213 5567 227
rect 5413 193 5427 207
rect 5593 193 5607 207
rect 133 173 147 187
rect 293 173 307 187
rect 333 173 347 187
rect 653 173 667 187
rect 713 173 727 187
rect 553 153 567 167
rect 713 153 727 167
rect 133 133 147 147
rect 174 133 188 147
rect 293 133 307 147
rect 433 133 447 147
rect 513 133 527 147
rect 633 133 647 147
rect 753 153 767 167
rect 873 153 887 167
rect 1213 173 1227 187
rect 1333 173 1347 187
rect 1633 173 1647 187
rect 1793 173 1807 187
rect 833 133 847 147
rect 913 133 927 147
rect 1113 133 1127 147
rect 1152 134 1166 148
rect 1373 153 1387 167
rect 1573 153 1587 167
rect 2073 173 2087 187
rect 2013 153 2027 167
rect 2113 173 2127 187
rect 2393 173 2407 187
rect 2813 173 2827 187
rect 2873 173 2887 187
rect 3333 173 3347 187
rect 3593 173 3607 187
rect 3633 173 3647 187
rect 4393 173 4407 187
rect 4613 173 4627 187
rect 4773 173 4787 187
rect 4933 173 4947 187
rect 5273 173 5287 187
rect 5353 173 5367 187
rect 2453 153 2467 167
rect 2714 153 2728 167
rect 1213 133 1227 147
rect 1313 133 1327 147
rect 1453 133 1467 147
rect 1673 133 1687 147
rect 1773 133 1787 147
rect 1872 133 1886 147
rect 1913 133 1927 147
rect 2153 133 2167 147
rect 2332 133 2346 147
rect 2374 133 2388 147
rect 493 113 507 127
rect 793 113 807 127
rect 893 113 907 127
rect 1173 113 1187 127
rect 1293 113 1307 127
rect 1413 113 1427 127
rect 2232 113 2246 127
rect 2273 113 2287 127
rect 2693 133 2707 147
rect 2953 133 2967 147
rect 3153 153 3167 167
rect 3233 153 3247 167
rect 2993 133 3007 147
rect 3373 133 3387 147
rect 2453 113 2467 127
rect 3932 153 3946 167
rect 4013 153 4027 167
rect 4113 153 4127 167
rect 4253 153 4267 167
rect 3792 133 3806 147
rect 3873 133 3887 147
rect 3953 133 3967 147
rect 4213 133 4227 147
rect 4573 153 4587 167
rect 4793 153 4807 167
rect 4953 153 4967 167
rect 5053 153 5067 167
rect 5313 153 5327 167
rect 5513 153 5527 167
rect 4533 133 4547 147
rect 4572 133 4586 147
rect 4613 133 4627 147
rect 4853 133 4867 147
rect 4933 133 4947 147
rect 5113 133 5127 147
rect 5173 133 5187 147
rect 5333 133 5347 147
rect 5553 133 5567 147
rect 1113 93 1127 107
rect 1213 93 1227 107
rect 1313 93 1327 107
rect 1793 93 1807 107
rect 3513 93 3527 107
rect 3613 113 3627 127
rect 3772 113 3786 127
rect 4173 113 4187 127
rect 4213 113 4227 127
rect 4373 113 4387 127
rect 4773 113 4787 127
rect 4873 113 4887 127
rect 5293 113 5307 127
rect 5453 113 5467 127
rect 3773 93 3787 107
rect 4252 93 4266 107
rect 4274 93 4288 107
rect 4313 93 4327 107
rect 4973 93 4987 107
rect 5293 93 5307 107
rect 5613 93 5627 107
rect 333 73 347 87
rect 753 73 767 87
rect 1813 73 1827 87
rect 3513 73 3527 87
rect 3633 74 3647 88
rect 4273 73 4287 87
rect 5233 73 5247 87
rect 5513 73 5527 87
rect 553 53 567 67
rect 913 53 927 67
rect 1153 53 1167 67
rect 1313 53 1327 67
rect 1373 53 1387 67
rect 1593 53 1607 67
rect 3633 52 3647 66
rect 4173 53 4187 67
rect 4313 53 4327 67
rect 853 33 867 47
rect 2953 33 2967 47
rect 3453 33 3467 47
rect 4073 33 4087 47
rect 5113 33 5127 47
rect 5153 33 5167 47
rect 5693 33 5707 47
rect 2993 13 3007 27
rect 3093 13 3107 27
rect 4533 13 4547 27
rect 5433 13 5447 27
<< metal3 >>
rect 316 5647 324 5673
rect 56 5487 64 5633
rect 196 5567 204 5613
rect 236 5587 244 5613
rect 336 5567 344 5613
rect 396 5587 404 5633
rect 480 5624 492 5627
rect 476 5613 492 5624
rect 56 5447 64 5473
rect 96 5247 104 5433
rect 236 5427 244 5533
rect 140 5424 153 5427
rect 136 5413 153 5424
rect 227 5416 244 5427
rect 276 5427 284 5493
rect 276 5416 293 5427
rect 227 5413 240 5416
rect 280 5413 293 5416
rect 116 5267 124 5393
rect 136 5227 144 5413
rect 353 5387 367 5393
rect 396 5387 404 5573
rect 476 5507 484 5613
rect 516 5607 524 5633
rect 516 5527 524 5593
rect 556 5567 564 5593
rect 596 5447 604 5713
rect 616 5627 624 5693
rect 796 5627 804 5653
rect 876 5647 884 5673
rect 1013 5667 1027 5673
rect 920 5664 933 5667
rect 916 5653 933 5664
rect 636 5567 644 5613
rect 696 5547 704 5593
rect 896 5587 904 5613
rect 536 5387 544 5433
rect 676 5427 684 5473
rect 696 5427 704 5453
rect 736 5407 744 5513
rect 727 5396 744 5407
rect 727 5393 740 5396
rect 336 5187 344 5213
rect 187 5184 200 5187
rect 240 5184 253 5187
rect 187 5173 204 5184
rect 73 5167 87 5173
rect 96 5136 133 5144
rect 96 5087 104 5136
rect 96 4947 104 5073
rect 156 4987 164 5113
rect 196 5027 204 5173
rect 236 5173 253 5184
rect 236 5087 244 5173
rect 307 5144 320 5147
rect 307 5133 324 5144
rect 356 5140 384 5144
rect 316 5007 324 5133
rect 353 5136 384 5140
rect 353 5127 367 5136
rect 320 4964 332 4967
rect 316 4953 332 4964
rect 87 4936 104 4947
rect 87 4933 100 4936
rect 36 4467 44 4933
rect 176 4927 184 4953
rect 200 4944 212 4947
rect 196 4933 212 4944
rect 76 4847 84 4893
rect 56 4687 64 4813
rect 116 4727 124 4893
rect 196 4887 204 4933
rect 156 4687 164 4833
rect 216 4687 224 4933
rect 316 4887 324 4953
rect 376 4947 384 5136
rect 396 4967 404 5373
rect 416 5067 424 5353
rect 756 5307 764 5453
rect 836 5427 844 5553
rect 916 5507 924 5653
rect 1127 5644 1140 5647
rect 1127 5633 1144 5644
rect 956 5567 964 5633
rect 907 5444 920 5447
rect 907 5433 924 5444
rect 776 5387 784 5413
rect 876 5327 884 5413
rect 916 5387 924 5433
rect 476 5167 484 5213
rect 773 5187 787 5193
rect 773 5180 774 5187
rect 433 5127 447 5133
rect 576 4967 584 5173
rect 896 5167 904 5293
rect 956 5267 964 5553
rect 996 5327 1004 5593
rect 1076 5567 1084 5633
rect 1136 5587 1144 5633
rect 1136 5487 1144 5573
rect 1196 5547 1204 5633
rect 1216 5567 1224 5593
rect 1053 5407 1067 5413
rect 1096 5387 1104 5413
rect 1176 5387 1184 5453
rect 1116 5207 1124 5333
rect 1136 5247 1144 5373
rect 1173 5367 1187 5373
rect 740 5164 752 5167
rect 736 5153 752 5164
rect 906 5153 907 5160
rect 616 5027 624 5153
rect 676 5087 684 5133
rect 736 5047 744 5153
rect 893 5140 907 5153
rect 896 5136 904 5140
rect 793 5107 807 5113
rect 507 4964 520 4967
rect 507 4953 524 4964
rect 356 4767 364 4913
rect 336 4667 344 4693
rect 396 4687 404 4853
rect 386 4676 404 4687
rect 386 4673 400 4676
rect 76 4487 84 4613
rect 96 4547 104 4653
rect 136 4447 144 4493
rect 93 4227 107 4233
rect 140 4204 153 4207
rect 136 4193 153 4204
rect 136 4167 144 4193
rect 116 4027 124 4053
rect 176 4047 184 4213
rect 216 4187 224 4453
rect 236 4447 244 4513
rect 260 4485 273 4487
rect 256 4474 273 4485
rect 256 4473 280 4474
rect 256 4427 264 4473
rect 280 4464 293 4467
rect 276 4453 293 4464
rect 276 4307 284 4453
rect 253 4247 267 4253
rect 280 4204 293 4207
rect 276 4193 293 4204
rect 227 4176 244 4184
rect 67 3964 80 3967
rect 67 3953 84 3964
rect 16 2907 24 3713
rect 76 3587 84 3953
rect 116 3947 124 4013
rect 176 3987 184 4033
rect 116 3707 124 3853
rect 156 3727 164 3933
rect 196 3927 204 3993
rect 116 3696 133 3707
rect 120 3693 133 3696
rect 176 3547 184 3693
rect 196 3527 204 3813
rect 236 3807 244 4176
rect 276 4147 284 4193
rect 276 4107 284 4133
rect 336 4087 344 4613
rect 376 4527 384 4633
rect 416 4627 424 4673
rect 456 4667 464 4853
rect 476 4827 484 4933
rect 516 4907 524 4953
rect 540 4944 553 4947
rect 536 4933 553 4944
rect 536 4847 544 4933
rect 616 4827 624 4933
rect 616 4707 624 4753
rect 636 4727 644 4953
rect 656 4787 664 4893
rect 676 4847 684 4913
rect 716 4887 724 4933
rect 776 4927 784 5073
rect 856 5047 864 5113
rect 856 4987 864 5033
rect 856 4976 873 4987
rect 860 4973 873 4976
rect 976 4967 984 5153
rect 1196 5147 1204 5533
rect 1296 5507 1304 5613
rect 1216 5307 1224 5473
rect 1236 5267 1244 5433
rect 1296 5407 1304 5493
rect 1316 5467 1324 5713
rect 1416 5587 1424 5653
rect 1340 5424 1353 5427
rect 1336 5413 1353 5424
rect 1296 5327 1304 5393
rect 1127 5144 1140 5147
rect 1127 5133 1144 5144
rect 1036 5004 1044 5133
rect 1036 4996 1053 5004
rect 973 4947 987 4953
rect 986 4940 987 4947
rect 1016 4887 1024 4933
rect 1056 4927 1064 4993
rect 1076 4987 1084 5113
rect 1136 5007 1144 5133
rect 1176 5027 1184 5113
rect 1156 4887 1164 4933
rect 516 4660 524 4664
rect 513 4647 527 4660
rect 516 4567 524 4633
rect 556 4627 564 4673
rect 656 4627 664 4653
rect 353 4447 367 4453
rect 356 4247 364 4433
rect 396 4287 404 4453
rect 336 3987 344 4033
rect 327 3976 344 3987
rect 327 3973 340 3976
rect 356 3967 364 4053
rect 396 4047 404 4193
rect 356 3956 373 3967
rect 360 3953 373 3956
rect 236 3747 244 3793
rect 276 3727 284 3913
rect 356 3727 364 3793
rect 316 3647 324 3693
rect 376 3667 384 3693
rect 236 3527 244 3573
rect 67 3524 80 3527
rect 67 3513 84 3524
rect 133 3513 134 3520
rect 76 3287 84 3513
rect 96 3467 104 3513
rect 133 3507 147 3513
rect 126 3500 147 3507
rect 126 3496 144 3500
rect 126 3493 140 3496
rect 236 3484 244 3513
rect 206 3476 244 3484
rect 67 3244 80 3247
rect 67 3233 84 3244
rect 76 2967 84 3233
rect 116 3227 124 3353
rect 196 3247 204 3393
rect 236 3247 244 3273
rect 296 3247 304 3433
rect 156 3047 164 3093
rect 196 3007 204 3133
rect 296 3087 304 3233
rect 220 3024 233 3027
rect 187 2996 204 3007
rect 216 3013 233 3024
rect 187 2993 200 2996
rect 76 2864 84 2893
rect 76 2856 104 2864
rect 56 2767 64 2813
rect 96 2767 104 2856
rect 106 2753 107 2760
rect 16 2687 24 2753
rect 93 2740 107 2753
rect 136 2747 144 2833
rect 96 2736 104 2740
rect 136 2736 152 2747
rect 140 2733 152 2736
rect 36 2667 44 2733
rect 93 2567 107 2573
rect 136 2567 144 2593
rect 36 2147 44 2513
rect 96 2308 104 2433
rect 67 2304 80 2307
rect 67 2293 84 2304
rect 76 2127 84 2293
rect 116 2284 124 2513
rect 156 2327 164 2733
rect 176 2607 184 2813
rect 196 2567 204 2913
rect 216 2848 224 3013
rect 216 2807 224 2812
rect 213 2780 227 2793
rect 216 2776 224 2780
rect 220 2766 240 2767
rect 227 2763 240 2766
rect 227 2753 244 2763
rect 236 2707 244 2753
rect 176 2447 184 2533
rect 156 2287 164 2313
rect 196 2288 204 2553
rect 213 2533 214 2540
rect 213 2527 227 2533
rect 256 2407 264 2933
rect 96 2280 124 2284
rect 93 2276 124 2280
rect 93 2267 107 2276
rect 116 2107 124 2133
rect 36 2027 44 2053
rect 36 1607 44 2013
rect 96 1927 104 2073
rect 76 1767 84 1833
rect 96 1787 104 1853
rect 156 1847 164 2113
rect 176 2067 184 2093
rect 156 1807 164 1833
rect 196 1827 204 2252
rect 236 2087 244 2113
rect 276 2087 284 2953
rect 296 2807 304 2993
rect 296 2587 304 2733
rect 316 2567 324 3633
rect 336 3487 344 3513
rect 336 3267 344 3473
rect 376 3447 384 3473
rect 356 3027 364 3073
rect 347 3016 364 3027
rect 347 3013 360 3016
rect 376 2967 384 3213
rect 393 3047 407 3053
rect 436 3047 444 4433
rect 496 4427 504 4473
rect 476 4416 492 4424
rect 476 4327 484 4416
rect 476 4247 484 4313
rect 516 4287 524 4413
rect 556 4264 564 4613
rect 596 4447 604 4513
rect 616 4487 624 4593
rect 653 4487 667 4493
rect 696 4427 704 4813
rect 756 4707 764 4753
rect 796 4687 804 4733
rect 836 4687 844 4753
rect 936 4687 944 4733
rect 1196 4707 1204 4733
rect 1187 4696 1204 4707
rect 1236 4707 1244 5193
rect 1296 5187 1304 5233
rect 1336 5227 1344 5413
rect 1396 5347 1404 5413
rect 1436 5347 1444 5593
rect 1476 5547 1484 5653
rect 1516 5647 1524 5733
rect 1456 5407 1464 5433
rect 1516 5427 1524 5513
rect 1556 5467 1564 5653
rect 1616 5647 1624 5673
rect 1656 5587 1664 5613
rect 1576 5427 1584 5473
rect 1576 5416 1593 5427
rect 1580 5413 1593 5416
rect 1616 5407 1624 5553
rect 1673 5447 1687 5453
rect 1716 5447 1724 5673
rect 1896 5647 1904 5733
rect 1980 5624 1993 5627
rect 1936 5620 1944 5624
rect 1933 5607 1947 5620
rect 1976 5613 1993 5624
rect 1376 5187 1384 5313
rect 1496 5287 1504 5393
rect 1836 5387 1844 5533
rect 1856 5447 1864 5473
rect 1853 5420 1867 5433
rect 1936 5427 1944 5593
rect 1976 5587 1984 5613
rect 1976 5527 1984 5573
rect 2036 5467 2044 5593
rect 2076 5447 2084 5533
rect 2116 5447 2124 5693
rect 2136 5647 2144 5673
rect 2296 5647 2304 5693
rect 2206 5593 2207 5600
rect 2193 5587 2207 5593
rect 2256 5567 2264 5633
rect 2296 5607 2304 5633
rect 2340 5624 2353 5627
rect 2336 5613 2353 5624
rect 2336 5587 2344 5613
rect 2396 5607 2404 5653
rect 2816 5647 2824 5673
rect 2907 5664 2920 5667
rect 2907 5653 2924 5664
rect 2446 5636 2493 5644
rect 2807 5636 2824 5647
rect 2860 5644 2873 5647
rect 2807 5633 2820 5636
rect 2856 5633 2873 5644
rect 1856 5416 1864 5420
rect 1987 5404 2000 5407
rect 1987 5393 2004 5404
rect 1996 5367 2004 5393
rect 1436 5167 1444 5233
rect 1556 5207 1564 5353
rect 2056 5347 2064 5413
rect 2208 5404 2220 5407
rect 2208 5393 2224 5404
rect 1460 5184 1473 5187
rect 1427 5156 1444 5167
rect 1456 5173 1473 5184
rect 1427 5153 1440 5156
rect 1456 5107 1464 5173
rect 1556 5147 1564 5193
rect 1296 4747 1304 5053
rect 1336 4804 1344 4973
rect 1396 4967 1404 5033
rect 1393 4940 1407 4953
rect 1396 4936 1404 4940
rect 1376 4827 1384 4893
rect 1336 4796 1364 4804
rect 1236 4696 1253 4707
rect 1187 4693 1200 4696
rect 1240 4693 1253 4696
rect 1296 4687 1304 4733
rect 796 4676 812 4687
rect 800 4673 812 4676
rect 936 4676 953 4687
rect 940 4673 953 4676
rect 1100 4684 1113 4687
rect 1096 4673 1113 4684
rect 1200 4686 1220 4687
rect 716 4487 724 4533
rect 756 4487 764 4593
rect 936 4547 944 4652
rect 1096 4607 1104 4673
rect 1207 4684 1220 4686
rect 1207 4673 1224 4684
rect 1287 4676 1304 4687
rect 1287 4673 1300 4676
rect 936 4467 944 4533
rect 976 4447 984 4593
rect 996 4527 1004 4553
rect 996 4487 1004 4513
rect 1076 4507 1084 4533
rect 1076 4467 1084 4493
rect 1136 4487 1144 4513
rect 1216 4507 1224 4673
rect 1333 4647 1347 4653
rect 1236 4467 1244 4593
rect 1273 4487 1287 4493
rect 1227 4456 1244 4467
rect 1227 4453 1240 4456
rect 976 4436 993 4447
rect 980 4433 993 4436
rect 536 4256 564 4264
rect 456 4067 464 4213
rect 536 4147 544 4256
rect 536 4007 544 4073
rect 480 4004 492 4007
rect 476 3993 492 4004
rect 476 3907 484 3993
rect 533 3947 547 3953
rect 476 3827 484 3893
rect 536 3787 544 3933
rect 476 3707 484 3733
rect 576 3707 584 4113
rect 596 4007 604 4093
rect 616 3987 624 4273
rect 636 4247 644 4413
rect 636 4147 644 4193
rect 676 4187 684 4233
rect 736 4187 744 4313
rect 856 4207 864 4253
rect 933 4193 934 4200
rect 666 4176 684 4187
rect 666 4173 680 4176
rect 696 4067 704 4173
rect 776 4147 784 4173
rect 736 4047 744 4113
rect 476 3706 500 3707
rect 476 3696 493 3706
rect 480 3693 493 3696
rect 527 3684 540 3687
rect 527 3673 544 3684
rect 536 3647 544 3673
rect 496 3547 504 3613
rect 496 3467 504 3533
rect 676 3527 684 3873
rect 476 3207 484 3293
rect 496 3287 504 3453
rect 533 3287 547 3293
rect 636 3247 644 3513
rect 527 3236 574 3244
rect 636 3227 644 3233
rect 626 3216 644 3227
rect 626 3213 640 3216
rect 696 3127 704 3953
rect 816 3747 824 4173
rect 856 4067 864 4193
rect 933 4187 947 4193
rect 876 4007 884 4133
rect 873 3980 887 3993
rect 876 3976 884 3980
rect 860 3966 880 3967
rect 860 3964 872 3966
rect 856 3953 872 3964
rect 856 3927 864 3953
rect 916 3907 924 3973
rect 976 3807 984 4353
rect 1076 4007 1084 4393
rect 1136 4027 1144 4353
rect 1156 3987 1164 4433
rect 1176 4127 1184 4193
rect 1236 4187 1244 4213
rect 856 3747 864 3773
rect 996 3767 1004 3933
rect 1036 3787 1044 3933
rect 1116 3887 1124 3973
rect 973 3727 987 3733
rect 986 3720 987 3727
rect 1000 3724 1012 3727
rect 996 3714 1012 3724
rect 996 3713 1020 3714
rect 733 3667 747 3673
rect 876 3667 884 3713
rect 996 3687 1004 3713
rect 1056 3707 1064 3753
rect 1156 3747 1164 3773
rect 1193 3727 1207 3733
rect 1016 3700 1024 3704
rect 1013 3687 1027 3700
rect 1056 3696 1073 3707
rect 1060 3693 1073 3696
rect 1013 3680 1014 3687
rect 716 3487 724 3553
rect 796 3527 804 3553
rect 920 3524 933 3527
rect 916 3513 933 3524
rect 716 3327 724 3473
rect 756 3447 764 3513
rect 776 3367 784 3453
rect 896 3447 904 3473
rect 836 3227 844 3353
rect 856 3247 864 3313
rect 896 3267 904 3433
rect 916 3367 924 3513
rect 1016 3407 1024 3673
rect 1176 3484 1184 3533
rect 1236 3507 1244 4013
rect 1276 3887 1284 3953
rect 1256 3527 1264 3793
rect 1296 3667 1304 3693
rect 1296 3567 1304 3613
rect 1267 3516 1284 3524
rect 1276 3487 1284 3516
rect 1156 3476 1184 3484
rect 1156 3367 1164 3476
rect 1013 3267 1027 3273
rect 1136 3267 1144 3293
rect 1176 3268 1184 3453
rect 1316 3287 1324 4053
rect 1336 3887 1344 4533
rect 1356 4207 1364 4796
rect 1396 4447 1404 4653
rect 1416 4564 1424 4893
rect 1456 4787 1464 5093
rect 1456 4707 1464 4773
rect 1416 4556 1444 4564
rect 1406 4444 1420 4447
rect 1406 4433 1424 4444
rect 1356 4107 1364 4153
rect 1336 3347 1344 3753
rect 1356 3627 1364 3993
rect 1376 3607 1384 4013
rect 1416 4007 1424 4433
rect 1396 3647 1404 3893
rect 1416 3587 1424 3953
rect 1436 3627 1444 4556
rect 1476 4467 1484 5133
rect 1576 5107 1584 5153
rect 1596 5147 1604 5293
rect 1696 5167 1704 5213
rect 1696 5156 1713 5167
rect 1700 5153 1713 5156
rect 1756 5147 1764 5273
rect 1776 5167 1784 5193
rect 1716 4967 1724 5093
rect 1713 4947 1727 4953
rect 1496 4887 1504 4933
rect 1496 4507 1504 4633
rect 1536 4547 1544 4933
rect 1756 4927 1764 5133
rect 1836 5087 1844 5193
rect 1873 5187 1887 5193
rect 1873 5180 1874 5187
rect 1936 5167 1944 5233
rect 1916 5087 1924 5133
rect 1866 4913 1867 4920
rect 1576 4827 1584 4913
rect 1853 4907 1867 4913
rect 1596 4707 1604 4733
rect 1616 4587 1624 4893
rect 1640 4684 1653 4687
rect 1636 4673 1653 4684
rect 1636 4627 1644 4673
rect 1736 4667 1744 4833
rect 1956 4807 1964 5313
rect 2016 4947 2024 5153
rect 2056 5147 2064 5333
rect 2116 5167 2124 5233
rect 2116 5156 2133 5167
rect 2120 5153 2133 5156
rect 2133 5107 2147 5113
rect 2096 4967 2104 4993
rect 2096 4927 2104 4953
rect 2136 4927 2144 4973
rect 2087 4916 2104 4927
rect 2087 4913 2100 4916
rect 2156 4747 2164 5393
rect 2216 5367 2224 5393
rect 2336 5267 2344 5573
rect 2436 5427 2444 5593
rect 2516 5467 2524 5613
rect 2696 5467 2704 5613
rect 2716 5567 2724 5633
rect 2428 5413 2444 5427
rect 2376 5247 2384 5413
rect 2216 5147 2224 5213
rect 2276 5147 2284 5213
rect 2356 5147 2364 5213
rect 2436 5207 2444 5413
rect 2716 5407 2724 5553
rect 2756 5424 2764 5593
rect 2856 5587 2864 5633
rect 2916 5607 2924 5653
rect 2936 5647 2944 5693
rect 2936 5636 2953 5647
rect 2940 5633 2953 5636
rect 2836 5427 2844 5453
rect 2756 5416 2773 5424
rect 2676 5227 2684 5393
rect 2716 5287 2724 5393
rect 2776 5384 2784 5413
rect 2776 5376 2804 5384
rect 2647 5184 2660 5187
rect 2647 5173 2664 5184
rect 2276 5136 2293 5147
rect 2280 5133 2293 5136
rect 2366 5133 2367 5140
rect 2353 5120 2367 5133
rect 2396 5127 2404 5173
rect 2487 5164 2500 5167
rect 2487 5153 2504 5164
rect 2356 5116 2364 5120
rect 2276 4967 2284 5073
rect 2316 5007 2324 5113
rect 2396 4967 2404 4993
rect 2176 4867 2184 4953
rect 2236 4887 2244 4953
rect 2436 4907 2444 5133
rect 2496 5107 2504 5153
rect 2596 4927 2604 5113
rect 2616 4947 2624 5153
rect 2656 5027 2664 5173
rect 2776 4967 2784 5033
rect 2796 5027 2804 5376
rect 2816 5067 2824 5393
rect 2896 5327 2904 5393
rect 2976 5387 2984 5453
rect 2873 5207 2887 5213
rect 2996 5187 3004 5233
rect 2988 5176 3004 5187
rect 2988 5173 3000 5176
rect 3036 5167 3044 5273
rect 2756 4956 2773 4964
rect 1726 4653 1727 4660
rect 1736 4656 1752 4667
rect 1740 4653 1752 4656
rect 1713 4647 1727 4653
rect 1456 3987 1464 4433
rect 1507 4204 1520 4207
rect 1507 4193 1524 4204
rect 1516 4127 1524 4193
rect 1536 4007 1544 4273
rect 1556 3987 1564 4493
rect 1576 4207 1584 4313
rect 1576 4167 1584 4193
rect 1596 4107 1604 4173
rect 1616 4168 1624 4453
rect 1573 3993 1574 4000
rect 1573 3987 1587 3993
rect 1456 3976 1473 3987
rect 1460 3973 1473 3976
rect 1566 3980 1587 3987
rect 1566 3976 1584 3980
rect 1566 3973 1580 3976
rect 1456 3707 1464 3873
rect 1516 3747 1524 3893
rect 1356 3447 1364 3493
rect 896 3207 904 3253
rect 1180 3244 1193 3247
rect 1176 3233 1193 3244
rect 1287 3244 1300 3247
rect 1287 3233 1304 3244
rect 533 3047 547 3053
rect 533 3040 534 3047
rect 476 2927 484 3013
rect 496 2987 504 3033
rect 616 3027 624 3073
rect 676 3027 684 3053
rect 776 3047 784 3113
rect 496 2907 504 2973
rect 616 2967 624 3013
rect 376 2747 384 2793
rect 493 2787 507 2793
rect 536 2787 544 2813
rect 406 2764 420 2767
rect 406 2753 424 2764
rect 416 2747 424 2753
rect 416 2736 433 2747
rect 420 2733 433 2736
rect 456 2707 464 2753
rect 336 2547 344 2573
rect 316 2288 324 2473
rect 336 2267 344 2533
rect 396 2507 404 2553
rect 436 2547 444 2613
rect 496 2607 504 2773
rect 556 2604 564 2713
rect 576 2627 584 2933
rect 596 2767 604 2893
rect 656 2747 664 2973
rect 836 2967 844 3013
rect 747 2744 760 2747
rect 747 2733 764 2744
rect 536 2596 564 2604
rect 487 2564 500 2567
rect 487 2553 504 2564
rect 496 2487 504 2553
rect 320 2266 344 2267
rect 327 2255 344 2266
rect 327 2253 340 2255
rect 126 1804 140 1807
rect 126 1800 144 1804
rect 126 1793 147 1800
rect 133 1787 147 1793
rect 133 1780 134 1787
rect 196 1667 204 1773
rect 116 1587 124 1633
rect 236 1607 244 1933
rect 296 1867 304 2053
rect 296 1827 304 1853
rect 316 1627 324 2193
rect 376 2127 384 2273
rect 436 2147 444 2353
rect 416 2088 424 2113
rect 456 2087 464 2393
rect 496 2308 504 2413
rect 536 2387 544 2596
rect 636 2567 644 2633
rect 556 2367 564 2513
rect 576 2347 584 2553
rect 716 2527 724 2633
rect 673 2507 687 2513
rect 516 2287 524 2333
rect 616 2287 624 2313
rect 656 2288 664 2393
rect 500 2286 524 2287
rect 507 2275 524 2286
rect 507 2273 520 2275
rect 696 2287 704 2373
rect 716 2307 724 2513
rect 756 2487 764 2733
rect 796 2627 804 2813
rect 836 2647 844 2853
rect 796 2587 804 2613
rect 856 2607 864 3193
rect 1056 3127 1064 3213
rect 1096 3167 1104 3233
rect 876 2987 884 3013
rect 876 2847 884 2973
rect 896 2747 904 3033
rect 936 2867 944 3113
rect 976 3007 984 3033
rect 996 2927 1004 3053
rect 1036 3027 1044 3053
rect 1116 3047 1124 3173
rect 1176 3127 1184 3233
rect 1276 3187 1284 3233
rect 1296 3207 1304 3233
rect 996 2867 1004 2913
rect 1076 2867 1084 2993
rect 916 2767 924 2833
rect 956 2787 964 2853
rect 1056 2767 1064 2813
rect 916 2756 933 2767
rect 920 2753 933 2756
rect 886 2736 904 2747
rect 886 2733 900 2736
rect 976 2627 984 2753
rect 1116 2727 1124 2793
rect 1016 2647 1024 2713
rect 796 2527 804 2573
rect 936 2544 944 2573
rect 916 2536 944 2544
rect 776 2327 784 2433
rect 836 2427 844 2513
rect 896 2487 904 2513
rect 916 2507 924 2536
rect 1016 2527 1024 2633
rect 1036 2567 1044 2713
rect 796 2327 804 2353
rect 856 2267 864 2333
rect 660 2264 672 2267
rect 656 2253 672 2264
rect 408 2064 420 2067
rect 408 2053 424 2064
rect 336 1847 344 1913
rect 336 1807 344 1833
rect 376 1727 384 1953
rect 416 1907 424 2053
rect 476 1887 484 2033
rect 536 1927 544 2033
rect 576 2007 584 2073
rect 587 1996 604 2004
rect 416 1747 424 1793
rect 476 1767 484 1833
rect 496 1827 504 1853
rect 516 1780 524 1784
rect 513 1767 527 1780
rect 356 1607 364 1673
rect 116 1576 133 1587
rect 120 1573 133 1576
rect 76 1507 84 1553
rect 116 1307 124 1552
rect 136 1307 144 1573
rect 196 1347 204 1593
rect 236 1327 244 1373
rect 316 1367 324 1493
rect 336 1367 344 1573
rect 236 1316 253 1327
rect 240 1313 253 1316
rect 96 1300 104 1304
rect 93 1287 107 1300
rect 136 1293 153 1307
rect 36 1107 44 1233
rect 96 1207 104 1273
rect 116 1187 124 1293
rect 96 1147 104 1153
rect 136 1147 144 1293
rect 93 1120 107 1133
rect 96 1116 104 1120
rect 176 1107 184 1153
rect 216 1087 224 1253
rect 276 1127 284 1333
rect 316 1327 324 1353
rect 356 1327 364 1593
rect 416 1587 424 1693
rect 516 1684 524 1753
rect 556 1687 564 1953
rect 576 1707 584 1913
rect 596 1807 604 1996
rect 656 1927 664 2253
rect 676 1947 684 2053
rect 716 1947 724 2113
rect 756 2047 764 2193
rect 796 2107 804 2213
rect 747 2036 764 2047
rect 796 2047 804 2093
rect 796 2036 813 2047
rect 747 2033 760 2036
rect 800 2033 813 2036
rect 636 1827 644 1893
rect 627 1816 644 1827
rect 627 1813 640 1816
rect 656 1807 664 1873
rect 696 1827 704 1913
rect 656 1796 673 1807
rect 660 1793 673 1796
rect 516 1680 544 1684
rect 516 1676 547 1680
rect 533 1667 547 1676
rect 473 1607 487 1613
rect 656 1607 664 1633
rect 376 1580 404 1584
rect 373 1576 404 1580
rect 416 1576 433 1587
rect 373 1567 387 1576
rect 396 1547 404 1576
rect 420 1573 433 1576
rect 356 1247 364 1313
rect 296 1107 304 1153
rect 216 1076 232 1087
rect 220 1073 232 1076
rect 96 807 104 893
rect 156 847 164 873
rect 193 844 207 853
rect 236 847 244 873
rect 193 840 224 844
rect 196 836 224 840
rect 96 796 113 807
rect 100 793 113 796
rect 176 767 184 793
rect 216 787 224 836
rect 236 807 244 833
rect 93 687 107 693
rect 176 627 184 753
rect 196 587 204 653
rect 216 627 224 773
rect 256 667 264 893
rect 216 616 233 627
rect 220 613 233 616
rect 276 567 284 1013
rect 316 687 324 1073
rect 396 1024 404 1533
rect 516 1367 524 1553
rect 576 1547 584 1593
rect 696 1567 704 1713
rect 736 1627 744 1913
rect 756 1827 764 1893
rect 796 1787 804 1873
rect 836 1647 844 2233
rect 856 2047 864 2093
rect 876 2064 884 2433
rect 916 2407 924 2493
rect 896 2287 904 2353
rect 916 2307 924 2393
rect 976 2327 984 2413
rect 996 2307 1004 2473
rect 1036 2327 1044 2493
rect 1076 2487 1084 2653
rect 1136 2547 1144 2853
rect 1196 2627 1204 3153
rect 1216 2807 1224 3013
rect 1256 2947 1264 2993
rect 1276 2767 1284 2833
rect 1156 2387 1164 2553
rect 1236 2544 1244 2753
rect 1216 2536 1244 2544
rect 1196 2507 1204 2533
rect 1216 2504 1224 2536
rect 1216 2496 1244 2504
rect 956 2067 964 2113
rect 996 2107 1004 2293
rect 1036 2287 1044 2313
rect 1176 2287 1184 2313
rect 1120 2284 1133 2287
rect 1116 2273 1133 2284
rect 876 2056 904 2064
rect 896 1887 904 2056
rect 1056 2047 1064 2233
rect 1116 2107 1124 2273
rect 1156 2087 1164 2113
rect 1056 2036 1073 2047
rect 1060 2033 1073 2036
rect 913 2007 927 2013
rect 1196 1907 1204 2433
rect 1236 2424 1244 2496
rect 1256 2467 1264 2513
rect 1216 2416 1244 2424
rect 1216 2187 1224 2416
rect 1233 2327 1247 2333
rect 1256 2187 1264 2253
rect 913 1847 927 1853
rect 716 1616 733 1624
rect 436 1187 444 1313
rect 436 1127 444 1173
rect 496 1147 504 1333
rect 548 1324 560 1327
rect 548 1313 564 1324
rect 556 1267 564 1313
rect 556 1087 564 1193
rect 376 1016 404 1024
rect 376 947 384 1016
rect 336 867 344 913
rect 336 707 344 853
rect 356 628 364 733
rect 376 647 384 853
rect 427 844 440 847
rect 427 833 444 844
rect 436 807 444 833
rect 456 767 464 833
rect 576 827 584 1373
rect 636 1347 644 1393
rect 636 1287 644 1333
rect 676 1227 684 1293
rect 676 1167 684 1213
rect 616 1107 624 1133
rect 607 1096 624 1107
rect 607 1093 620 1096
rect 676 1067 684 1093
rect 696 927 704 1413
rect 596 847 604 913
rect 716 907 724 1616
rect 836 1607 844 1633
rect 776 1567 784 1593
rect 876 1584 884 1753
rect 896 1747 904 1773
rect 933 1767 947 1773
rect 976 1687 984 1813
rect 1036 1807 1044 1833
rect 1027 1796 1044 1807
rect 1027 1793 1040 1796
rect 1073 1773 1074 1780
rect 996 1747 1004 1773
rect 1073 1767 1087 1773
rect 933 1604 947 1613
rect 1016 1607 1024 1733
rect 1056 1647 1064 1693
rect 1056 1607 1064 1633
rect 1136 1627 1144 1773
rect 1156 1607 1164 1793
rect 1176 1727 1184 1753
rect 916 1600 947 1604
rect 916 1596 944 1600
rect 916 1584 924 1596
rect 1048 1596 1064 1607
rect 1048 1593 1060 1596
rect 856 1576 884 1584
rect 896 1580 924 1584
rect 893 1576 924 1580
rect 856 1447 864 1576
rect 893 1567 907 1576
rect 906 1560 907 1567
rect 916 1427 924 1553
rect 796 1327 804 1353
rect 936 1327 944 1393
rect 1016 1387 1024 1593
rect 1076 1527 1084 1553
rect 887 1324 900 1327
rect 887 1313 904 1324
rect 756 1187 764 1293
rect 756 1127 764 1173
rect 796 1167 804 1313
rect 836 1227 844 1313
rect 856 1227 864 1293
rect 896 1247 904 1313
rect 747 1116 764 1127
rect 747 1113 760 1116
rect 796 1087 804 1153
rect 856 1107 864 1213
rect 896 1087 904 1233
rect 996 1167 1004 1333
rect 1076 1287 1084 1513
rect 1116 1307 1124 1453
rect 1176 1367 1184 1713
rect 1236 1707 1244 2153
rect 1276 2127 1284 2153
rect 1276 2067 1284 2113
rect 1196 1447 1204 1693
rect 1276 1627 1284 1773
rect 1296 1767 1304 3113
rect 1316 2567 1324 3073
rect 1356 3027 1364 3193
rect 1376 3047 1384 3513
rect 1456 3507 1464 3593
rect 1436 3387 1444 3473
rect 1396 3147 1404 3253
rect 1456 3087 1464 3493
rect 1476 3407 1484 3613
rect 1536 3527 1544 3953
rect 1596 3847 1604 3953
rect 1556 3727 1564 3813
rect 1556 3716 1573 3727
rect 1560 3713 1573 3716
rect 1596 3687 1604 3773
rect 1556 3567 1564 3593
rect 1616 3567 1624 4132
rect 1636 4048 1644 4553
rect 1656 4507 1664 4593
rect 1656 4467 1664 4493
rect 1696 4467 1704 4573
rect 1756 4567 1764 4613
rect 1736 4487 1744 4533
rect 1796 4487 1804 4693
rect 1900 4684 1912 4687
rect 1896 4673 1912 4684
rect 1856 4487 1864 4633
rect 1896 4607 1904 4673
rect 1736 4476 1753 4487
rect 1740 4473 1753 4476
rect 1696 4307 1704 4453
rect 1756 4267 1764 4473
rect 1916 4467 1924 4533
rect 1927 4456 1944 4464
rect 1936 4427 1944 4456
rect 1956 4447 1964 4733
rect 2033 4693 2034 4700
rect 2016 4667 2024 4693
rect 2033 4684 2047 4693
rect 2033 4680 2113 4684
rect 2036 4676 2113 4680
rect 2076 4607 2084 4653
rect 1996 4460 2024 4464
rect 1993 4456 2024 4460
rect 1993 4447 2007 4456
rect 2006 4440 2007 4447
rect 1916 4367 1924 4393
rect 2016 4387 2024 4456
rect 2056 4407 2064 4513
rect 2116 4487 2124 4633
rect 2113 4460 2127 4473
rect 2116 4456 2124 4460
rect 1836 4227 1844 4253
rect 1806 4224 1820 4227
rect 1806 4220 1824 4224
rect 1806 4213 1827 4220
rect 1680 4204 1692 4207
rect 1676 4193 1692 4204
rect 1676 4147 1684 4193
rect 1736 4187 1744 4213
rect 1813 4207 1827 4213
rect 1813 4200 1814 4207
rect 1776 4127 1784 4193
rect 1640 4026 1660 4027
rect 1647 4023 1660 4026
rect 1647 4013 1664 4023
rect 1656 3947 1664 4013
rect 1776 3887 1784 3953
rect 1636 3684 1644 3833
rect 1656 3747 1664 3793
rect 1736 3767 1744 3833
rect 1656 3707 1664 3733
rect 1756 3707 1764 3813
rect 1776 3727 1784 3753
rect 1636 3676 1664 3684
rect 1576 3447 1584 3513
rect 1656 3507 1664 3676
rect 1736 3547 1744 3573
rect 1733 3520 1747 3533
rect 1776 3527 1784 3673
rect 1736 3516 1744 3520
rect 1476 3027 1484 3293
rect 1516 3027 1524 3433
rect 1353 2967 1367 2973
rect 1356 2747 1364 2953
rect 1456 2767 1464 2993
rect 1476 2947 1484 3013
rect 1556 2987 1564 3333
rect 1576 3227 1584 3433
rect 1616 3307 1624 3493
rect 1696 3287 1704 3413
rect 1736 3307 1744 3333
rect 1713 3273 1714 3280
rect 1713 3264 1727 3273
rect 1776 3267 1784 3513
rect 1796 3287 1804 3933
rect 1816 3904 1824 4153
rect 1896 4007 1904 4193
rect 1887 3996 1904 4007
rect 1887 3993 1900 3996
rect 1916 3967 1924 4353
rect 1936 4264 1944 4333
rect 1936 4256 1964 4264
rect 1956 4207 1964 4256
rect 2033 4224 2047 4233
rect 2056 4224 2064 4393
rect 2033 4220 2064 4224
rect 2036 4216 2064 4220
rect 1948 4193 1964 4207
rect 1913 3947 1927 3953
rect 1816 3896 1844 3904
rect 1816 3687 1824 3873
rect 1836 3607 1844 3896
rect 1956 3847 1964 4193
rect 1976 4067 1984 4173
rect 1996 4107 2004 4193
rect 2056 4087 2064 4216
rect 2076 4207 2084 4293
rect 2076 4107 2084 4193
rect 2116 4187 2124 4213
rect 2156 4207 2164 4253
rect 2096 4007 2104 4053
rect 2116 3987 2124 4093
rect 2116 3927 2124 3973
rect 1856 3667 1864 3773
rect 1896 3707 1904 3733
rect 1976 3707 1984 3773
rect 1696 3260 1727 3264
rect 1696 3256 1724 3260
rect 1576 3047 1584 3213
rect 1656 2907 1664 3213
rect 1656 2767 1664 2893
rect 1696 2867 1704 3256
rect 1736 2827 1744 3253
rect 1756 3027 1764 3113
rect 1316 2327 1324 2493
rect 1376 2307 1384 2573
rect 1396 2367 1404 2613
rect 1436 2467 1444 2533
rect 1340 2284 1353 2287
rect 1336 2273 1353 2284
rect 1336 2124 1344 2273
rect 1356 2167 1364 2233
rect 1416 2227 1424 2433
rect 1436 2287 1444 2453
rect 1316 2116 1344 2124
rect 1316 2047 1324 2116
rect 1436 2107 1444 2173
rect 1456 2164 1464 2633
rect 1516 2627 1524 2733
rect 1500 2544 1513 2547
rect 1496 2533 1513 2544
rect 1496 2307 1504 2533
rect 1536 2507 1544 2573
rect 1616 2567 1624 2613
rect 1516 2247 1524 2313
rect 1556 2267 1564 2313
rect 1576 2207 1584 2513
rect 1596 2244 1604 2393
rect 1613 2287 1627 2293
rect 1596 2236 1624 2244
rect 1456 2156 1484 2164
rect 1436 2096 1453 2107
rect 1440 2093 1453 2096
rect 1336 2067 1344 2093
rect 1476 2067 1484 2156
rect 1616 2124 1624 2236
rect 1656 2147 1664 2653
rect 1676 2408 1684 2773
rect 1696 2647 1704 2753
rect 1776 2727 1784 3033
rect 1616 2116 1644 2124
rect 1496 2087 1504 2113
rect 1336 2056 1353 2067
rect 1340 2053 1353 2056
rect 1316 2046 1340 2047
rect 1316 2035 1333 2046
rect 1320 2033 1333 2035
rect 1516 1987 1524 2053
rect 1556 1927 1564 2093
rect 1636 2047 1644 2116
rect 1656 2107 1664 2133
rect 1676 2067 1684 2372
rect 1696 2287 1704 2593
rect 1716 2127 1724 2713
rect 1776 2647 1784 2713
rect 1776 2587 1784 2593
rect 1773 2560 1787 2573
rect 1776 2556 1784 2560
rect 1736 2467 1744 2533
rect 1756 2387 1764 2553
rect 1796 2547 1804 2953
rect 1816 2947 1824 3553
rect 1856 3387 1864 3473
rect 1876 3367 1884 3533
rect 1916 3487 1924 3633
rect 1916 3476 1933 3487
rect 1920 3473 1933 3476
rect 1896 3267 1904 3433
rect 1976 3387 1984 3533
rect 1996 3447 2004 3913
rect 2016 3767 2024 3813
rect 2096 3787 2104 3893
rect 2036 3687 2044 3713
rect 2056 3667 2064 3733
rect 2116 3707 2124 3733
rect 2096 3604 2104 3633
rect 2076 3596 2104 3604
rect 2016 3547 2024 3573
rect 2076 3507 2084 3596
rect 2116 3527 2124 3693
rect 1836 3047 1844 3173
rect 1856 2787 1864 3093
rect 1876 2987 1884 3033
rect 1916 3027 1924 3153
rect 1907 3016 1924 3027
rect 1907 3013 1920 3016
rect 1820 2744 1833 2747
rect 1816 2733 1833 2744
rect 1816 2667 1824 2733
rect 1876 2727 1884 2973
rect 1936 2887 1944 3233
rect 1956 3027 1964 3253
rect 1976 3227 1984 3313
rect 1996 3107 2004 3353
rect 2036 3344 2044 3433
rect 2116 3347 2124 3473
rect 2016 3336 2044 3344
rect 2016 3107 2024 3336
rect 2060 3264 2073 3267
rect 2056 3253 2073 3264
rect 2056 3107 2064 3253
rect 2116 3147 2124 3253
rect 2136 3167 2144 4113
rect 2196 4047 2204 4793
rect 2376 4667 2384 4893
rect 2376 4656 2393 4667
rect 2380 4653 2393 4656
rect 2296 4487 2304 4573
rect 2356 4567 2364 4653
rect 2416 4607 2424 4673
rect 2296 4476 2313 4487
rect 2300 4473 2313 4476
rect 2416 4467 2424 4593
rect 2436 4547 2444 4653
rect 2236 4408 2244 4433
rect 2236 4247 2244 4372
rect 2256 4347 2264 4453
rect 2296 4207 2304 4373
rect 2376 4307 2384 4413
rect 2236 4127 2244 4193
rect 2196 4036 2213 4047
rect 2200 4033 2213 4036
rect 2256 4027 2264 4173
rect 2316 4167 2324 4213
rect 2376 4187 2384 4253
rect 2176 3884 2184 4013
rect 2296 3967 2304 4073
rect 2176 3876 2204 3884
rect 2156 3467 2164 3833
rect 2196 3747 2204 3876
rect 2193 3687 2207 3693
rect 2216 3487 2224 3953
rect 2236 3707 2244 3853
rect 2356 3747 2364 4133
rect 2416 4007 2424 4333
rect 2436 4087 2444 4493
rect 2456 3907 2464 4733
rect 2476 4127 2484 4853
rect 2496 4147 2504 4833
rect 2596 4787 2604 4913
rect 2656 4687 2664 4953
rect 2676 4767 2684 4913
rect 2696 4787 2704 4953
rect 2756 4807 2764 4956
rect 2796 4867 2804 4973
rect 2896 4967 2904 5013
rect 2840 4924 2853 4927
rect 2836 4913 2853 4924
rect 2836 4847 2844 4913
rect 2836 4787 2844 4833
rect 2520 4684 2533 4687
rect 2516 4673 2533 4684
rect 2516 4488 2524 4673
rect 2616 4527 2624 4673
rect 2520 4464 2533 4467
rect 2516 4453 2533 4464
rect 2516 4387 2524 4453
rect 2596 4427 2604 4473
rect 2636 4427 2644 4453
rect 2516 4167 2524 4313
rect 2556 4247 2564 4413
rect 2676 4367 2684 4753
rect 2696 4527 2704 4613
rect 2716 4504 2724 4673
rect 2776 4664 2784 4773
rect 2796 4688 2804 4773
rect 2800 4664 2813 4667
rect 2776 4656 2813 4664
rect 2796 4653 2813 4656
rect 2696 4500 2724 4504
rect 2693 4496 2724 4500
rect 2693 4487 2707 4496
rect 2736 4487 2744 4513
rect 2706 4480 2707 4487
rect 2696 4407 2704 4433
rect 2556 4187 2564 4233
rect 2636 4227 2644 4353
rect 2736 4307 2744 4433
rect 2587 4204 2600 4207
rect 2587 4196 2624 4204
rect 2587 4193 2604 4196
rect 2476 3964 2484 4013
rect 2536 4007 2544 4093
rect 2556 3984 2564 4133
rect 2596 4107 2604 4193
rect 2616 4167 2624 4196
rect 2660 4184 2672 4187
rect 2656 4173 2672 4184
rect 2536 3976 2564 3984
rect 2476 3956 2504 3964
rect 2236 3667 2244 3693
rect 2256 3547 2264 3733
rect 2336 3547 2344 3613
rect 2356 3528 2364 3693
rect 2396 3687 2404 3733
rect 2436 3727 2444 3793
rect 2427 3716 2444 3727
rect 2427 3713 2440 3716
rect 2476 3704 2484 3913
rect 2456 3696 2484 3704
rect 2256 3447 2264 3473
rect 2193 3287 2207 3293
rect 2176 3240 2184 3244
rect 2173 3227 2187 3240
rect 2056 3047 2064 3093
rect 2096 3048 2104 3113
rect 2113 3067 2127 3073
rect 2113 3060 2114 3067
rect 1956 3016 1973 3027
rect 1960 3013 1973 3016
rect 2088 3024 2100 3027
rect 2088 3013 2104 3024
rect 1796 2536 1813 2547
rect 1800 2533 1813 2536
rect 1836 2524 1844 2553
rect 1816 2516 1844 2524
rect 1776 2327 1784 2513
rect 1776 2247 1784 2313
rect 1816 2287 1824 2516
rect 1856 2504 1864 2653
rect 1876 2527 1884 2593
rect 1896 2507 1904 2773
rect 1916 2527 1924 2813
rect 1936 2760 1944 2764
rect 1933 2747 1947 2760
rect 1936 2587 1944 2733
rect 1956 2507 1964 2713
rect 1976 2607 1984 2833
rect 2036 2807 2044 2953
rect 2096 2947 2104 3013
rect 2116 2844 2124 3053
rect 2136 2867 2144 3013
rect 2156 2847 2164 3193
rect 2176 3127 2184 3213
rect 2236 3087 2244 3413
rect 2256 3267 2264 3373
rect 2180 3044 2193 3047
rect 2176 3033 2193 3044
rect 2176 2867 2184 3033
rect 2096 2836 2124 2844
rect 2096 2827 2104 2836
rect 2096 2747 2104 2813
rect 2096 2736 2113 2747
rect 2100 2733 2113 2736
rect 1996 2547 2004 2733
rect 2156 2627 2164 2753
rect 2040 2524 2053 2527
rect 2036 2513 2053 2524
rect 1836 2496 1864 2504
rect 1676 2007 1684 2053
rect 1696 2047 1704 2093
rect 1716 2087 1724 2113
rect 1776 2084 1784 2233
rect 1776 2076 1804 2084
rect 1708 2036 1724 2044
rect 1316 1667 1324 1793
rect 1356 1687 1364 1773
rect 1220 1584 1233 1587
rect 1216 1573 1233 1584
rect 1216 1527 1224 1573
rect 1336 1547 1344 1573
rect 1216 1367 1224 1453
rect 1176 1327 1184 1353
rect 1236 1327 1244 1413
rect 1276 1347 1284 1393
rect 1116 1296 1133 1307
rect 1120 1293 1133 1296
rect 936 1127 944 1153
rect 1016 1067 1024 1133
rect 1036 1127 1044 1253
rect 1076 1127 1084 1233
rect 1216 1227 1224 1313
rect 740 864 753 867
rect 736 853 753 864
rect 596 836 612 847
rect 600 834 612 836
rect 600 833 620 834
rect 620 824 632 827
rect 616 813 632 824
rect 616 767 624 813
rect 696 787 704 833
rect 736 767 744 853
rect 816 767 824 833
rect 856 767 864 853
rect 936 767 944 833
rect 976 827 984 1053
rect 1116 1047 1124 1113
rect 1116 1004 1124 1033
rect 1096 996 1124 1004
rect 496 627 504 733
rect 596 647 604 673
rect 756 667 764 693
rect 316 600 373 604
rect 313 596 373 600
rect 313 587 327 596
rect 636 587 644 613
rect 176 387 184 513
rect 216 367 224 433
rect 93 327 107 333
rect 216 327 224 353
rect 256 347 264 413
rect 136 147 144 173
rect 176 147 184 273
rect 316 207 324 353
rect 356 347 364 553
rect 487 384 500 387
rect 487 373 504 384
rect 400 364 413 367
rect 396 353 413 364
rect 396 287 404 353
rect 296 147 304 173
rect 336 87 344 173
rect 456 147 464 293
rect 447 136 464 147
rect 447 133 460 136
rect 496 127 504 373
rect 536 327 544 393
rect 556 367 564 553
rect 556 356 573 367
rect 560 353 573 356
rect 616 287 624 533
rect 676 467 684 633
rect 756 627 764 653
rect 856 627 864 753
rect 1016 727 1024 933
rect 1056 767 1064 813
rect 747 616 764 627
rect 747 613 760 616
rect 636 327 644 453
rect 696 427 704 593
rect 856 587 864 613
rect 688 364 700 367
rect 688 353 704 364
rect 516 207 524 253
rect 516 147 524 193
rect 556 67 564 153
rect 616 147 624 273
rect 656 187 664 333
rect 696 287 704 353
rect 736 347 744 433
rect 796 387 804 493
rect 836 367 844 413
rect 836 356 853 367
rect 840 353 853 356
rect 896 347 904 473
rect 713 167 727 173
rect 616 136 633 147
rect 620 133 633 136
rect 756 87 764 153
rect 796 127 804 293
rect 916 247 924 713
rect 996 627 1004 693
rect 1073 667 1087 673
rect 1056 387 1064 553
rect 1096 547 1104 996
rect 1136 827 1144 1173
rect 1196 1107 1204 1153
rect 1187 1096 1204 1107
rect 1187 1093 1200 1096
rect 1156 947 1164 1073
rect 1216 1027 1224 1093
rect 1196 827 1204 873
rect 1196 816 1213 827
rect 1200 813 1213 816
rect 1136 687 1144 813
rect 1156 627 1164 753
rect 1236 707 1244 1253
rect 1256 847 1264 1193
rect 1296 1087 1304 1213
rect 1376 1187 1384 1693
rect 1456 1627 1464 1793
rect 1416 1527 1424 1593
rect 1456 1547 1464 1573
rect 1476 1487 1484 1593
rect 1496 1567 1504 1713
rect 1416 1347 1424 1433
rect 1516 1407 1524 1853
rect 1536 1427 1544 1773
rect 1576 1648 1584 1993
rect 1696 1847 1704 1953
rect 1636 1707 1644 1793
rect 1716 1724 1724 2036
rect 1736 1847 1744 1873
rect 1756 1867 1764 2053
rect 1796 1947 1804 2076
rect 1816 1867 1824 2093
rect 1836 2067 1844 2496
rect 1896 2407 1904 2493
rect 1976 2307 1984 2513
rect 2036 2467 2044 2513
rect 2096 2507 2104 2553
rect 2136 2547 2144 2593
rect 2176 2567 2184 2773
rect 2196 2707 2204 2773
rect 2236 2607 2244 2933
rect 2256 2827 2264 3253
rect 2276 2847 2284 3513
rect 2296 3407 2304 3433
rect 2296 3267 2304 3333
rect 2306 3253 2307 3260
rect 2293 3240 2307 3253
rect 2296 3236 2304 3240
rect 2336 3167 2344 3233
rect 2356 3187 2364 3492
rect 2376 3207 2384 3653
rect 2416 3487 2424 3573
rect 2436 3307 2444 3493
rect 2456 3327 2464 3696
rect 2416 3187 2424 3213
rect 2316 3047 2324 3133
rect 2356 3047 2364 3073
rect 2376 3047 2384 3153
rect 2307 3036 2324 3047
rect 2307 3033 2320 3036
rect 2376 3033 2393 3047
rect 2296 2947 2304 2993
rect 2276 2724 2284 2833
rect 2256 2716 2284 2724
rect 2136 2533 2152 2547
rect 1996 2307 2004 2333
rect 1880 2264 1892 2267
rect 1876 2253 1892 2264
rect 1856 2207 1864 2253
rect 1876 2107 1884 2253
rect 1896 2087 1904 2133
rect 1936 1907 1944 2273
rect 2056 2267 2064 2293
rect 1967 2264 1980 2267
rect 1967 2253 1984 2264
rect 1976 2167 1984 2253
rect 2016 2067 2024 2133
rect 2016 2056 2033 2067
rect 2020 2053 2033 2056
rect 1960 2044 1972 2047
rect 1956 2033 1972 2044
rect 1956 1887 1964 2033
rect 1996 1887 2004 1993
rect 2056 1927 2064 2253
rect 2096 2244 2104 2493
rect 2136 2347 2144 2533
rect 2076 2236 2104 2244
rect 2076 2167 2084 2236
rect 2076 2107 2084 2153
rect 2096 2047 2104 2113
rect 2116 2027 2124 2093
rect 2133 2027 2147 2033
rect 2133 2020 2134 2027
rect 1736 1787 1744 1833
rect 1696 1716 1724 1724
rect 1576 1587 1584 1612
rect 1616 1587 1624 1673
rect 1656 1587 1664 1653
rect 1696 1647 1704 1716
rect 1716 1527 1724 1573
rect 1516 1384 1524 1393
rect 1516 1376 1544 1384
rect 1536 1347 1544 1376
rect 1353 1147 1367 1153
rect 1316 1067 1324 1093
rect 1456 1087 1464 1133
rect 1376 1027 1384 1073
rect 1316 867 1324 913
rect 1276 787 1284 813
rect 1316 727 1324 793
rect 1216 627 1224 673
rect 1156 616 1172 627
rect 1160 613 1172 616
rect 1136 407 1144 533
rect 1093 387 1107 393
rect 1196 367 1204 473
rect 1256 467 1264 633
rect 1316 624 1324 713
rect 1356 667 1364 853
rect 1456 707 1464 833
rect 1496 767 1504 833
rect 1516 807 1524 1313
rect 1576 1208 1584 1493
rect 1736 1387 1744 1733
rect 1756 1347 1764 1633
rect 1556 947 1564 1053
rect 1576 887 1584 1172
rect 1596 1047 1604 1073
rect 1576 827 1584 873
rect 1636 867 1644 1313
rect 1676 1167 1684 1253
rect 1696 1147 1704 1292
rect 1756 1287 1764 1333
rect 1776 1324 1784 1553
rect 1796 1467 1804 1793
rect 1876 1767 1884 1813
rect 2076 1807 2084 1953
rect 1993 1793 1994 1800
rect 1886 1753 1887 1760
rect 1873 1747 1887 1753
rect 1936 1727 1944 1793
rect 1993 1787 2007 1793
rect 1873 1607 1887 1613
rect 1896 1547 1904 1673
rect 1916 1607 1924 1653
rect 1936 1627 1944 1713
rect 2027 1604 2040 1607
rect 2027 1593 2044 1604
rect 1776 1316 1793 1324
rect 1796 1247 1804 1313
rect 1736 1127 1744 1233
rect 1836 1167 1844 1373
rect 1856 1187 1864 1493
rect 1976 1487 1984 1573
rect 2036 1567 2044 1593
rect 2056 1507 2064 1673
rect 2076 1347 2084 1713
rect 2116 1367 2124 1913
rect 2136 1627 2144 2013
rect 2156 1907 2164 2493
rect 2196 2467 2204 2573
rect 2176 2307 2184 2333
rect 2176 2297 2193 2307
rect 2180 2294 2193 2297
rect 2180 2293 2200 2294
rect 2156 1787 2164 1853
rect 2196 1807 2204 2272
rect 2236 2047 2244 2193
rect 2256 2127 2264 2716
rect 2276 2587 2284 2693
rect 2296 2507 2304 2933
rect 2316 2887 2324 2913
rect 2316 2747 2324 2873
rect 2356 2747 2364 2853
rect 2376 2787 2384 3033
rect 2356 2733 2373 2747
rect 2316 2667 2324 2733
rect 2356 2627 2364 2733
rect 2396 2707 2404 2973
rect 2336 2616 2353 2624
rect 2316 2547 2324 2573
rect 2316 2424 2324 2533
rect 2296 2416 2324 2424
rect 2296 2267 2304 2416
rect 2336 2267 2344 2616
rect 2416 2567 2424 3113
rect 2436 3087 2444 3293
rect 2456 3127 2464 3313
rect 2476 3107 2484 3673
rect 2496 3567 2504 3956
rect 2536 3847 2544 3976
rect 2576 3847 2584 3973
rect 2516 3747 2524 3793
rect 2616 3747 2624 4073
rect 2656 4067 2664 4173
rect 2716 4167 2724 4193
rect 2756 4187 2764 4553
rect 2796 4467 2804 4653
rect 2876 4607 2884 4833
rect 2916 4807 2924 4933
rect 2956 4847 2964 5133
rect 2988 4964 3000 4967
rect 2988 4953 3004 4964
rect 2996 4867 3004 4953
rect 2916 4687 2924 4793
rect 2936 4747 2944 4813
rect 2976 4667 2984 4693
rect 2987 4664 3000 4667
rect 2987 4653 3004 4664
rect 2916 4547 2924 4633
rect 2916 4507 2924 4533
rect 2787 4456 2804 4467
rect 2787 4453 2800 4456
rect 2836 4407 2844 4433
rect 2836 4267 2844 4393
rect 2796 4067 2804 4173
rect 2876 4167 2884 4353
rect 2936 4227 2944 4593
rect 2976 4527 2984 4553
rect 2996 4507 3004 4653
rect 3016 4647 3024 4713
rect 3036 4507 3044 4873
rect 3056 4807 3064 4893
rect 3076 4527 3084 5353
rect 3116 5147 3124 5413
rect 3136 5347 3144 5613
rect 3176 5447 3184 5633
rect 3236 5567 3244 5673
rect 3416 5627 3424 5653
rect 3616 5647 3624 5824
rect 4116 5787 4124 5824
rect 3836 5647 3844 5673
rect 3416 5527 3424 5613
rect 3236 5407 3244 5453
rect 3356 5447 3364 5473
rect 3196 5327 3204 5393
rect 3376 5227 3384 5453
rect 3096 4687 3104 4893
rect 3136 4884 3144 5053
rect 3116 4876 3144 4884
rect 3116 4707 3124 4876
rect 3156 4647 3164 4853
rect 3196 4727 3204 5173
rect 3236 5127 3244 5153
rect 3296 5147 3304 5173
rect 3347 5164 3360 5167
rect 3347 5153 3364 5164
rect 3236 4967 3244 5113
rect 3216 4787 3224 4833
rect 3236 4707 3244 4793
rect 3296 4727 3304 5133
rect 3356 5127 3364 5153
rect 3396 5147 3404 5513
rect 3416 5327 3424 5453
rect 3436 5407 3444 5473
rect 3456 5147 3464 5573
rect 3516 5367 3524 5633
rect 3616 5547 3624 5633
rect 3756 5587 3764 5633
rect 3648 5424 3660 5427
rect 3648 5413 3664 5424
rect 3516 5187 3524 5353
rect 3556 5347 3564 5413
rect 3656 5367 3664 5413
rect 3356 5007 3364 5073
rect 3436 5047 3444 5113
rect 3396 4967 3404 4993
rect 3227 4696 3244 4707
rect 3227 4693 3240 4696
rect 3147 4636 3164 4647
rect 3147 4633 3160 4636
rect 2956 4207 2964 4313
rect 2807 4004 2820 4007
rect 2807 3993 2824 4004
rect 2688 3964 2700 3967
rect 2688 3953 2704 3964
rect 2656 3787 2664 3953
rect 2696 3907 2704 3953
rect 2707 3896 2724 3904
rect 2716 3748 2724 3896
rect 2736 3827 2744 3973
rect 2816 3967 2824 3993
rect 2956 3984 2964 4193
rect 2976 4007 2984 4073
rect 2996 4027 3004 4193
rect 2956 3976 2984 3984
rect 2876 3907 2884 3973
rect 2496 3127 2504 3453
rect 2516 3148 2524 3373
rect 2556 3247 2564 3593
rect 2596 3467 2604 3673
rect 2616 3647 2624 3733
rect 2856 3727 2864 3773
rect 2907 3744 2920 3747
rect 2907 3733 2924 3744
rect 2656 3547 2664 3693
rect 2716 3687 2724 3712
rect 2767 3704 2780 3707
rect 2767 3693 2784 3704
rect 2736 3527 2744 3653
rect 2776 3587 2784 3693
rect 2816 3667 2824 3713
rect 2916 3687 2924 3733
rect 2936 3664 2944 3833
rect 2956 3727 2964 3753
rect 2936 3656 2964 3664
rect 2728 3516 2744 3527
rect 2728 3513 2740 3516
rect 2556 3236 2573 3247
rect 2560 3233 2573 3236
rect 2576 3147 2584 3233
rect 2496 3126 2520 3127
rect 2496 3113 2513 3126
rect 2476 2847 2484 3013
rect 2496 2987 2504 3113
rect 2596 3027 2604 3073
rect 2587 3016 2604 3027
rect 2587 3013 2600 3016
rect 2448 2784 2460 2787
rect 2448 2773 2464 2784
rect 2456 2627 2464 2773
rect 2356 2348 2364 2553
rect 2436 2327 2444 2593
rect 2456 2487 2464 2533
rect 2476 2447 2484 2793
rect 2496 2427 2504 2633
rect 2516 2587 2524 2833
rect 2536 2747 2544 3013
rect 2616 3004 2624 3513
rect 2676 3247 2684 3493
rect 2716 3387 2724 3513
rect 2856 3504 2864 3573
rect 2916 3527 2924 3573
rect 2936 3548 2944 3633
rect 2856 3496 2893 3504
rect 2716 3267 2724 3333
rect 2816 3327 2824 3493
rect 2836 3307 2844 3433
rect 2936 3347 2944 3512
rect 2667 3236 2684 3247
rect 2667 3233 2680 3236
rect 2656 3207 2664 3233
rect 2736 3207 2744 3293
rect 2796 3227 2804 3273
rect 2736 3107 2744 3193
rect 2636 3007 2644 3033
rect 2656 3027 2664 3093
rect 2776 3087 2784 3193
rect 2696 3027 2704 3053
rect 2616 2996 2633 3004
rect 2556 2607 2564 2953
rect 2656 2947 2664 3013
rect 2576 2747 2584 2813
rect 2576 2587 2584 2653
rect 2573 2560 2587 2573
rect 2576 2556 2584 2560
rect 2596 2547 2604 2773
rect 2616 2424 2624 2893
rect 2676 2527 2684 2833
rect 2596 2416 2624 2424
rect 2596 2367 2604 2416
rect 2516 2327 2524 2353
rect 2227 2036 2244 2047
rect 2227 2033 2240 2036
rect 2236 1807 2244 1933
rect 2156 1776 2173 1787
rect 2160 1773 2173 1776
rect 1827 1156 1844 1167
rect 1827 1153 1840 1156
rect 1727 1116 1744 1127
rect 1727 1113 1740 1116
rect 1796 1087 1804 1133
rect 1836 927 1844 993
rect 1636 827 1644 853
rect 1696 827 1704 873
rect 1776 827 1784 853
rect 1767 816 1784 827
rect 1767 813 1780 816
rect 1816 807 1824 893
rect 1296 620 1324 624
rect 1293 616 1324 620
rect 1293 607 1307 616
rect 1456 604 1464 693
rect 1496 647 1504 753
rect 1536 627 1544 653
rect 1556 647 1564 733
rect 1596 687 1604 773
rect 1596 647 1604 673
rect 1636 627 1644 693
rect 1756 647 1764 693
rect 1796 627 1804 773
rect 1836 687 1844 913
rect 1836 647 1844 673
rect 1636 616 1653 627
rect 1640 613 1653 616
rect 1456 596 1493 604
rect 1256 367 1264 393
rect 1296 387 1304 493
rect 1476 407 1484 533
rect 1340 384 1353 387
rect 1336 373 1353 384
rect 1000 364 1013 367
rect 996 353 1013 364
rect 1256 356 1273 367
rect 1260 353 1273 356
rect 996 327 1004 353
rect 856 147 864 233
rect 1216 227 1224 333
rect 1336 287 1344 373
rect 1476 347 1484 393
rect 1516 367 1524 453
rect 1516 356 1532 367
rect 1520 353 1532 356
rect 1413 327 1427 333
rect 847 133 864 147
rect 856 47 864 133
rect 876 127 884 153
rect 1156 148 1164 213
rect 1336 187 1344 273
rect 1213 164 1227 173
rect 1213 160 1244 164
rect 1216 156 1244 160
rect 876 116 893 127
rect 880 113 893 116
rect 916 67 924 133
rect 1116 107 1124 133
rect 1160 124 1173 127
rect 1156 113 1173 124
rect 1156 67 1164 113
rect 1216 107 1224 133
rect 1236 124 1244 156
rect 1236 116 1293 124
rect 1316 107 1324 133
rect 1316 67 1324 93
rect 1376 67 1384 153
rect 1416 127 1424 193
rect 1436 147 1444 213
rect 1467 193 1473 207
rect 1636 187 1644 393
rect 1656 367 1664 553
rect 1776 376 1813 384
rect 1656 356 1673 367
rect 1660 353 1673 356
rect 1696 267 1704 313
rect 1587 164 1600 167
rect 1587 153 1604 164
rect 1633 160 1647 173
rect 1636 156 1644 160
rect 1436 136 1453 147
rect 1440 133 1453 136
rect 1596 67 1604 153
rect 1656 147 1664 213
rect 1776 147 1784 376
rect 1836 367 1844 493
rect 1856 387 1864 1133
rect 1936 1127 1944 1253
rect 1976 1127 1984 1213
rect 1876 827 1884 873
rect 1996 867 2004 913
rect 2016 887 2024 1313
rect 2036 1067 2044 1093
rect 1916 827 1924 853
rect 2056 847 2064 893
rect 2047 833 2064 847
rect 1956 787 1964 833
rect 1936 647 1944 733
rect 1976 647 1984 753
rect 2036 447 2044 753
rect 2056 747 2064 833
rect 2076 827 2084 1273
rect 2136 1127 2144 1573
rect 2176 1087 2184 1273
rect 2076 816 2093 827
rect 2080 813 2093 816
rect 2136 607 2144 793
rect 2156 667 2164 693
rect 2156 627 2164 653
rect 2156 616 2173 627
rect 2160 613 2173 616
rect 2127 596 2144 607
rect 2127 593 2140 596
rect 2176 487 2184 573
rect 2196 447 2204 1613
rect 2256 1607 2264 1893
rect 2296 1807 2304 1893
rect 2336 1847 2344 2253
rect 2356 1907 2364 2312
rect 2376 2187 2384 2273
rect 2436 2067 2444 2113
rect 2476 2087 2484 2173
rect 2467 2073 2484 2087
rect 2476 1987 2484 2073
rect 2496 1967 2504 2293
rect 2516 2187 2524 2233
rect 2516 2087 2524 2113
rect 2516 2076 2533 2087
rect 2520 2073 2533 2076
rect 2416 1807 2424 1853
rect 2476 1787 2484 1813
rect 2516 1807 2524 1973
rect 2366 1776 2394 1784
rect 2296 1587 2304 1633
rect 2216 1487 2224 1573
rect 2216 1027 2224 1353
rect 2260 1344 2273 1347
rect 2256 1333 2273 1344
rect 2233 1267 2247 1273
rect 2256 1247 2264 1333
rect 2316 1307 2324 1493
rect 2336 1407 2344 1433
rect 2356 1348 2364 1433
rect 2256 1127 2264 1233
rect 2296 1187 2304 1233
rect 2356 1227 2364 1312
rect 2376 1247 2384 1753
rect 2396 1427 2404 1573
rect 2436 1407 2444 1693
rect 2396 1327 2404 1373
rect 2436 1347 2444 1393
rect 2456 1367 2464 1653
rect 2476 1427 2484 1593
rect 2556 1467 2564 2193
rect 2576 2088 2584 2293
rect 2596 2067 2604 2273
rect 2656 2067 2664 2293
rect 2716 2287 2724 2873
rect 2756 2767 2764 3053
rect 2736 2687 2744 2713
rect 2776 2707 2784 2733
rect 2796 2627 2804 3173
rect 2856 3047 2864 3153
rect 2896 3147 2904 3193
rect 2956 3164 2964 3656
rect 2976 3367 2984 3976
rect 3016 3967 3024 4233
rect 3036 3867 3044 4493
rect 3056 4347 3064 4473
rect 3096 4387 3104 4473
rect 3056 4307 3064 4333
rect 3136 4227 3144 4513
rect 3176 4484 3184 4693
rect 3216 4487 3224 4633
rect 3256 4487 3264 4713
rect 3316 4567 3324 4693
rect 3356 4527 3364 4933
rect 3396 4924 3404 4953
rect 3376 4916 3404 4924
rect 3376 4727 3384 4916
rect 3376 4587 3384 4713
rect 3156 4480 3184 4484
rect 3153 4476 3184 4480
rect 3153 4467 3167 4476
rect 3336 4467 3344 4493
rect 3376 4487 3384 4573
rect 3166 4460 3167 4467
rect 3156 4207 3164 4253
rect 3196 4227 3204 4453
rect 3236 4427 3244 4453
rect 3156 4196 3173 4207
rect 3160 4193 3173 4196
rect 3056 4027 3064 4153
rect 3196 4087 3204 4213
rect 3236 4187 3244 4413
rect 3276 4207 3284 4393
rect 3267 4196 3284 4207
rect 3267 4193 3280 4196
rect 3296 4147 3304 4193
rect 3336 4167 3344 4233
rect 3053 4000 3067 4013
rect 3056 3996 3064 4000
rect 3213 3984 3227 3993
rect 3236 3984 3244 4093
rect 3336 4067 3344 4153
rect 3376 4147 3384 4173
rect 3213 3980 3244 3984
rect 3216 3976 3244 3980
rect 3056 3887 3064 3913
rect 3076 3807 3084 3953
rect 3096 3787 3104 3973
rect 3187 3964 3200 3967
rect 3187 3953 3204 3964
rect 3196 3867 3204 3953
rect 3256 3847 3264 3953
rect 3116 3807 3124 3833
rect 3016 3707 3024 3773
rect 3056 3727 3064 3773
rect 3136 3747 3144 3813
rect 3007 3696 3024 3707
rect 3007 3693 3020 3696
rect 3056 3607 3064 3713
rect 3136 3707 3144 3733
rect 3208 3704 3220 3707
rect 3208 3693 3224 3704
rect 3076 3667 3084 3693
rect 3036 3304 3044 3493
rect 3096 3487 3104 3673
rect 3116 3507 3124 3553
rect 3136 3524 3144 3693
rect 3216 3627 3224 3693
rect 3196 3527 3204 3593
rect 3256 3567 3264 3773
rect 3276 3687 3284 4033
rect 3376 4027 3384 4133
rect 3353 3747 3367 3753
rect 3276 3547 3284 3673
rect 3233 3527 3247 3533
rect 3356 3527 3364 3593
rect 3136 3516 3164 3524
rect 3156 3427 3164 3516
rect 3233 3520 3234 3527
rect 3036 3296 3064 3304
rect 3020 3284 3033 3287
rect 3016 3273 3033 3284
rect 2996 3247 3004 3273
rect 2956 3156 2984 3164
rect 2847 3036 2864 3047
rect 2847 3033 2860 3036
rect 2736 2327 2744 2433
rect 2680 2084 2693 2087
rect 2576 2056 2593 2064
rect 2396 1313 2413 1327
rect 2516 1320 2524 1324
rect 2396 1247 2404 1313
rect 2247 1116 2264 1127
rect 2247 1113 2260 1116
rect 2296 1107 2304 1133
rect 2336 1127 2344 1193
rect 2216 787 2224 833
rect 2216 707 2224 773
rect 2236 447 2244 1073
rect 2276 827 2284 873
rect 2316 847 2324 913
rect 2356 647 2364 1173
rect 2416 1107 2424 1133
rect 2476 1127 2484 1313
rect 2513 1307 2527 1320
rect 2496 1107 2504 1253
rect 2516 1167 2524 1293
rect 2556 1107 2564 1213
rect 2407 1096 2424 1107
rect 2407 1093 2420 1096
rect 2436 844 2444 993
rect 2556 904 2564 1093
rect 2536 896 2564 904
rect 2436 836 2464 844
rect 2280 644 2293 647
rect 2276 633 2293 644
rect 2276 467 2284 633
rect 1656 136 1673 147
rect 1660 133 1673 136
rect 1796 107 1804 173
rect 1816 87 1824 333
rect 1856 147 1864 233
rect 1916 147 1924 293
rect 1956 207 1964 353
rect 2036 327 2044 393
rect 2116 387 2124 433
rect 1976 207 1984 233
rect 2016 167 2024 193
rect 2076 187 2084 293
rect 2116 187 2124 273
rect 2156 207 2164 253
rect 2236 247 2244 393
rect 2376 387 2384 653
rect 2396 640 2404 644
rect 2393 627 2407 640
rect 2406 620 2407 627
rect 2396 587 2404 613
rect 2416 607 2424 813
rect 2436 687 2444 773
rect 2456 667 2464 836
rect 2476 648 2484 853
rect 2536 848 2544 896
rect 2576 867 2584 2056
rect 2647 2056 2664 2067
rect 2676 2073 2693 2084
rect 2647 2053 2660 2056
rect 2596 1807 2604 1853
rect 2636 1827 2644 2053
rect 2676 2007 2684 2073
rect 2636 1816 2653 1827
rect 2640 1813 2653 1816
rect 2596 1007 2604 1753
rect 2696 1687 2704 1933
rect 2716 1607 2724 2053
rect 2707 1596 2724 1607
rect 2707 1593 2720 1596
rect 2716 1507 2724 1553
rect 2616 1327 2624 1373
rect 2656 1247 2664 1313
rect 2716 1127 2724 1213
rect 2616 847 2624 1093
rect 2736 1047 2744 1733
rect 2756 1687 2764 2193
rect 2796 2067 2804 2613
rect 2816 2488 2824 2953
rect 2816 2287 2824 2452
rect 2836 2207 2844 2973
rect 2853 2787 2867 2793
rect 2896 2764 2904 3053
rect 2916 2847 2924 3093
rect 2956 2907 2964 3133
rect 2976 2967 2984 3156
rect 2996 2947 3004 3013
rect 3016 2887 3024 3273
rect 3056 3267 3064 3296
rect 2896 2756 2924 2764
rect 2856 2687 2864 2713
rect 2896 2664 2904 2733
rect 2876 2656 2904 2664
rect 2876 2627 2884 2656
rect 2916 2647 2924 2756
rect 2936 2687 2944 2753
rect 2996 2747 3004 2793
rect 3036 2767 3044 2893
rect 2956 2567 2964 2693
rect 3056 2687 3064 2953
rect 2916 2560 2924 2564
rect 2913 2547 2927 2560
rect 2956 2556 2973 2567
rect 2960 2553 2973 2556
rect 2926 2540 2927 2547
rect 2876 2407 2884 2513
rect 2916 2467 2924 2533
rect 2816 2107 2824 2133
rect 2816 2067 2824 2093
rect 2856 2047 2864 2253
rect 2776 1887 2784 2013
rect 2876 2007 2884 2353
rect 2916 2187 2924 2393
rect 2936 2147 2944 2313
rect 2976 2247 2984 2273
rect 2967 2236 2984 2247
rect 2967 2233 2980 2236
rect 2996 2224 3004 2533
rect 3036 2267 3044 2633
rect 3056 2347 3064 2673
rect 3076 2647 3084 3393
rect 3096 3067 3104 3253
rect 3116 2987 3124 3053
rect 3136 3027 3144 3213
rect 3156 3147 3164 3353
rect 3176 3027 3184 3293
rect 3236 3267 3244 3413
rect 3376 3368 3384 3853
rect 3233 3167 3247 3173
rect 3236 2987 3244 3113
rect 3256 3047 3264 3233
rect 3376 3187 3384 3332
rect 3376 3087 3384 3113
rect 3293 3047 3307 3053
rect 3293 3040 3294 3047
rect 3096 2787 3104 2853
rect 3076 2567 3084 2633
rect 3096 2267 3104 2393
rect 3116 2324 3124 2873
rect 3336 2867 3344 3033
rect 3396 3027 3404 4793
rect 3416 4647 3424 4693
rect 3436 4687 3444 5033
rect 3456 4747 3464 4913
rect 3476 4907 3484 4973
rect 3556 4947 3564 5333
rect 3456 4667 3464 4733
rect 3496 4687 3504 4833
rect 3476 4676 3493 4684
rect 3416 4407 3424 4633
rect 3436 4467 3444 4613
rect 3436 4456 3453 4467
rect 3440 4453 3453 4456
rect 3476 4304 3484 4676
rect 3516 4447 3524 4933
rect 3576 4807 3584 5273
rect 3696 5227 3704 5573
rect 3776 5407 3784 5513
rect 3796 5447 3804 5593
rect 3836 5584 3844 5633
rect 4016 5607 4024 5753
rect 3816 5576 3844 5584
rect 3816 5527 3824 5576
rect 3756 5247 3764 5373
rect 3700 5164 3714 5167
rect 3696 5160 3714 5164
rect 3693 5153 3714 5160
rect 3693 5148 3707 5153
rect 3706 5140 3707 5148
rect 3596 4987 3604 5133
rect 3596 4687 3604 4973
rect 3636 4827 3644 5093
rect 3567 4644 3580 4647
rect 3567 4633 3584 4644
rect 3576 4567 3584 4633
rect 3616 4544 3624 4793
rect 3656 4627 3664 4913
rect 3596 4536 3624 4544
rect 3567 4464 3580 4467
rect 3567 4453 3584 4464
rect 3476 4300 3504 4304
rect 3476 4296 3507 4300
rect 3493 4287 3507 4296
rect 3416 4227 3424 4273
rect 3416 4107 3424 4173
rect 3416 3787 3424 4053
rect 3416 3707 3424 3733
rect 3416 3547 3424 3693
rect 3436 3524 3444 4233
rect 3576 4228 3584 4453
rect 3596 4247 3604 4536
rect 3676 4527 3684 5073
rect 3696 4807 3704 5112
rect 3756 5007 3764 5133
rect 3767 4944 3780 4947
rect 3767 4933 3784 4944
rect 3776 4907 3784 4933
rect 3756 4744 3764 4873
rect 3796 4787 3804 5433
rect 3816 5408 3824 5433
rect 3816 5067 3824 5372
rect 3856 5327 3864 5553
rect 3876 5287 3884 5453
rect 3893 5387 3907 5393
rect 3856 5147 3864 5253
rect 3847 5133 3864 5147
rect 3856 4967 3864 5133
rect 3896 5127 3904 5293
rect 3896 4987 3904 5053
rect 3856 4956 3873 4967
rect 3860 4953 3873 4956
rect 3747 4736 3764 4744
rect 3736 4667 3744 4733
rect 3776 4647 3784 4693
rect 3816 4624 3824 4673
rect 3807 4616 3824 4624
rect 3656 4467 3664 4493
rect 3656 4367 3664 4453
rect 3676 4327 3684 4473
rect 3573 4187 3587 4192
rect 3496 3987 3504 4153
rect 3460 3984 3472 3987
rect 3456 3973 3472 3984
rect 3496 3976 3513 3987
rect 3500 3973 3513 3976
rect 3456 3867 3464 3973
rect 3556 3867 3564 3953
rect 3576 3947 3584 4013
rect 3616 3987 3624 4153
rect 3716 4124 3724 4473
rect 3796 4467 3804 4613
rect 3896 4487 3904 4593
rect 3836 4407 3844 4433
rect 3916 4407 3924 5533
rect 4116 5527 4124 5553
rect 4156 5487 4164 5773
rect 4236 5647 4244 5753
rect 4276 5687 4284 5773
rect 4216 5527 4224 5593
rect 4233 5447 4247 5453
rect 4233 5440 4234 5447
rect 3936 5248 3944 5393
rect 3976 5367 3984 5413
rect 3976 5307 3984 5353
rect 3936 5047 3944 5212
rect 3956 5007 3964 5193
rect 3996 5087 4004 5133
rect 4036 5127 4044 5373
rect 4156 5147 4164 5313
rect 4216 5307 4224 5413
rect 4296 5247 4304 5653
rect 4036 5116 4053 5127
rect 4040 5113 4053 5116
rect 4096 5107 4104 5133
rect 4176 5104 4184 5153
rect 4167 5096 4184 5104
rect 3953 4980 3967 4993
rect 3956 4976 3964 4980
rect 3936 4727 3944 4933
rect 3956 4747 3964 4813
rect 3936 4667 3944 4713
rect 3976 4687 3984 4913
rect 3996 4827 4004 4893
rect 3946 4653 3947 4660
rect 3933 4640 3947 4653
rect 3936 4636 3944 4640
rect 3956 4487 3964 4513
rect 3756 4247 3764 4313
rect 3796 4227 3804 4353
rect 3796 4216 3813 4227
rect 3800 4213 3813 4216
rect 3696 4116 3724 4124
rect 3556 3687 3564 3753
rect 3436 3516 3464 3524
rect 3416 3247 3424 3373
rect 3436 3227 3444 3433
rect 3456 3347 3464 3516
rect 3476 3247 3484 3653
rect 3496 3487 3504 3533
rect 3576 3427 3584 3833
rect 3616 3748 3624 3853
rect 3656 3727 3664 3773
rect 3616 3587 3624 3712
rect 3616 3507 3624 3573
rect 3608 3496 3624 3507
rect 3608 3493 3620 3496
rect 3536 3307 3544 3413
rect 3536 3267 3544 3293
rect 3387 3013 3404 3027
rect 3396 2967 3404 3013
rect 3416 3007 3424 3173
rect 3316 2807 3324 2853
rect 3316 2796 3333 2807
rect 3320 2793 3333 2796
rect 3236 2647 3244 2713
rect 3276 2647 3284 2713
rect 3176 2616 3213 2624
rect 3136 2447 3144 2533
rect 3176 2367 3184 2616
rect 3296 2567 3304 2653
rect 3336 2647 3344 2733
rect 3356 2527 3364 2593
rect 3256 2487 3264 2513
rect 3116 2316 3144 2324
rect 2976 2216 3004 2224
rect 2816 1967 2824 1993
rect 2816 1864 2824 1953
rect 2796 1856 2824 1864
rect 2796 1767 2804 1856
rect 2856 1767 2864 1973
rect 2936 1964 2944 2053
rect 2916 1960 2944 1964
rect 2913 1956 2944 1960
rect 2913 1947 2927 1956
rect 2936 1847 2944 1913
rect 2956 1807 2964 2173
rect 2776 1756 2793 1764
rect 2776 1667 2784 1756
rect 2760 1604 2773 1607
rect 2756 1593 2773 1604
rect 2756 1527 2764 1593
rect 2856 1547 2864 1613
rect 2876 1607 2884 1793
rect 2976 1787 2984 2216
rect 2996 1947 3004 2033
rect 2996 1827 3004 1933
rect 2907 1784 2920 1787
rect 2907 1773 2924 1784
rect 2896 1648 2904 1773
rect 2916 1708 2924 1773
rect 3016 1767 3024 2093
rect 3036 1927 3044 2073
rect 3056 1907 3064 2233
rect 3096 2087 3104 2133
rect 3136 2107 3144 2316
rect 3160 2264 3173 2267
rect 3156 2253 3173 2264
rect 3096 2076 3112 2087
rect 3100 2074 3112 2076
rect 3100 2073 3120 2074
rect 3100 2066 3120 2067
rect 3107 2063 3120 2066
rect 3107 2053 3124 2063
rect 3116 1987 3124 2053
rect 3156 1987 3164 2253
rect 3216 2127 3224 2433
rect 3236 2248 3244 2293
rect 3236 2047 3244 2212
rect 3276 2147 3284 2293
rect 3316 2167 3324 2453
rect 3376 2327 3384 2933
rect 3436 2847 3444 3213
rect 3456 3027 3464 3193
rect 3476 3107 3484 3233
rect 3576 3227 3584 3273
rect 3587 3216 3604 3224
rect 3456 2907 3464 3013
rect 3396 2427 3404 2673
rect 3416 2647 3424 2693
rect 3416 2567 3424 2633
rect 3436 2627 3444 2653
rect 3456 2607 3464 2853
rect 3436 2507 3444 2533
rect 3376 2167 3384 2253
rect 3416 2247 3424 2473
rect 3436 2307 3444 2493
rect 3276 2067 3284 2133
rect 3227 2036 3244 2047
rect 3227 2033 3240 2036
rect 3136 1887 3144 1953
rect 3047 1804 3060 1807
rect 3047 1793 3064 1804
rect 3116 1807 3124 1853
rect 3153 1827 3167 1833
rect 3107 1797 3124 1807
rect 3107 1794 3120 1797
rect 3100 1793 3120 1794
rect 2796 1447 2804 1513
rect 2876 1507 2884 1553
rect 2896 1347 2904 1612
rect 2756 1247 2764 1313
rect 2756 1107 2764 1193
rect 2796 1167 2804 1273
rect 2636 867 2644 913
rect 2656 827 2664 953
rect 2527 824 2540 827
rect 2527 813 2544 824
rect 2576 820 2584 824
rect 2536 767 2544 813
rect 2573 807 2587 820
rect 2576 747 2584 793
rect 2656 707 2664 813
rect 2696 784 2704 1033
rect 2736 787 2744 993
rect 2836 867 2844 1133
rect 2856 1127 2864 1253
rect 2896 1207 2904 1333
rect 2856 1047 2864 1113
rect 2827 856 2844 867
rect 2827 853 2840 856
rect 2856 847 2864 893
rect 2876 887 2884 1093
rect 2916 888 2924 1672
rect 2936 1587 2944 1753
rect 2936 1347 2944 1413
rect 2956 1387 2964 1673
rect 2988 1564 3000 1567
rect 2988 1553 3004 1564
rect 2996 1487 3004 1553
rect 2956 1307 2964 1373
rect 3016 1327 3024 1753
rect 3036 1628 3044 1753
rect 3056 1727 3064 1793
rect 3176 1787 3184 1953
rect 3236 1907 3244 1933
rect 3276 1867 3284 1933
rect 3273 1847 3287 1853
rect 3176 1776 3193 1787
rect 3180 1773 3193 1776
rect 3216 1784 3224 1813
rect 3207 1776 3224 1784
rect 3036 1367 3044 1592
rect 3096 1587 3104 1772
rect 3236 1687 3244 1793
rect 3316 1684 3324 1973
rect 3336 1827 3344 2113
rect 3416 2067 3424 2173
rect 3436 2164 3444 2253
rect 3456 2184 3464 2513
rect 3476 2207 3484 2513
rect 3496 2427 3504 3073
rect 3516 2447 3524 3133
rect 3596 3047 3604 3216
rect 3540 3044 3552 3047
rect 3536 3033 3552 3044
rect 3536 2947 3544 3033
rect 3536 2647 3544 2933
rect 3536 2307 3544 2633
rect 3556 2527 3564 2993
rect 3576 2827 3584 2993
rect 3616 2807 3624 2973
rect 3506 2253 3507 2260
rect 3493 2247 3507 2253
rect 3456 2176 3484 2184
rect 3436 2156 3464 2164
rect 3396 2056 3413 2064
rect 3356 1707 3364 1913
rect 3316 1676 3344 1684
rect 3136 1587 3144 1653
rect 3236 1627 3244 1673
rect 2996 1316 3013 1324
rect 2856 836 2873 847
rect 2860 833 2873 836
rect 2687 776 2704 784
rect 2616 627 2624 693
rect 2676 667 2684 773
rect 2776 727 2784 833
rect 2607 616 2624 627
rect 2607 613 2620 616
rect 2396 407 2404 533
rect 2436 367 2444 413
rect 2113 160 2127 173
rect 2116 156 2124 160
rect 2156 147 2164 193
rect 1856 136 1872 147
rect 1860 133 1872 136
rect 2216 127 2224 193
rect 2276 127 2284 233
rect 2396 187 2404 213
rect 2456 167 2464 413
rect 2476 267 2484 612
rect 2676 607 2684 653
rect 2666 593 2667 600
rect 2653 587 2667 593
rect 2567 384 2580 387
rect 2567 373 2584 384
rect 2496 207 2504 373
rect 2576 287 2584 373
rect 2616 367 2624 553
rect 2696 427 2704 693
rect 2736 647 2744 713
rect 2727 637 2744 647
rect 2727 634 2740 637
rect 2720 633 2740 634
rect 2716 587 2724 612
rect 2796 387 2804 753
rect 2716 347 2724 373
rect 2768 364 2780 367
rect 2768 353 2784 364
rect 2346 136 2374 144
rect 2456 127 2464 153
rect 2696 147 2704 313
rect 2776 227 2784 353
rect 2816 347 2824 793
rect 2836 567 2844 773
rect 2916 767 2924 852
rect 2916 607 2924 653
rect 2956 647 2964 1233
rect 2976 687 2984 873
rect 2996 827 3004 1316
rect 3056 1307 3064 1573
rect 3136 1487 3144 1573
rect 3336 1507 3344 1676
rect 3376 1567 3384 2013
rect 3396 1867 3404 2056
rect 3416 1887 3424 1913
rect 3436 1807 3444 2093
rect 3400 1784 3413 1787
rect 3396 1774 3413 1784
rect 3396 1773 3420 1774
rect 3396 1647 3404 1773
rect 3456 1768 3464 2156
rect 3476 1887 3484 2176
rect 3516 2087 3524 2173
rect 3536 2087 3544 2233
rect 3536 2076 3553 2087
rect 3540 2073 3553 2076
rect 3576 2067 3584 2613
rect 3596 2587 3604 2753
rect 3636 2628 3644 3533
rect 3676 3467 3684 4013
rect 3696 4007 3704 4116
rect 3716 3747 3724 4073
rect 3756 3867 3764 3953
rect 3756 3827 3764 3853
rect 3816 3847 3824 4113
rect 3856 4027 3864 4213
rect 3916 4200 3924 4204
rect 3913 4187 3927 4200
rect 3916 4167 3924 4173
rect 3847 4013 3864 4027
rect 3856 3887 3864 4013
rect 3716 3733 3733 3747
rect 3716 3707 3724 3733
rect 3796 3727 3804 3753
rect 3736 3507 3744 3593
rect 3756 3587 3764 3713
rect 3856 3667 3864 3713
rect 3727 3496 3744 3507
rect 3727 3493 3740 3496
rect 3768 3504 3780 3507
rect 3768 3493 3784 3504
rect 3776 3427 3784 3493
rect 3676 3227 3684 3393
rect 3716 3227 3724 3333
rect 3676 3216 3692 3227
rect 3680 3213 3692 3216
rect 3656 3007 3664 3093
rect 3676 2967 3684 3113
rect 3656 2748 3664 2813
rect 3633 2587 3647 2592
rect 3593 2560 3607 2573
rect 3596 2556 3604 2560
rect 3656 2547 3664 2712
rect 3656 2387 3664 2533
rect 3676 2367 3684 2793
rect 3696 2507 3704 3113
rect 3776 3047 3784 3213
rect 3796 3087 3804 3413
rect 3716 2887 3724 2993
rect 3736 2987 3744 3013
rect 3776 2887 3784 3033
rect 3716 2407 3724 2813
rect 3736 2767 3744 2833
rect 3736 2447 3744 2753
rect 3776 2747 3784 2833
rect 3816 2827 3824 3633
rect 3836 3567 3844 3613
rect 3836 3147 3844 3493
rect 3876 3488 3884 4133
rect 3896 4007 3904 4093
rect 3896 3968 3904 3993
rect 3856 2927 3864 3353
rect 3856 2747 3864 2873
rect 3876 2807 3884 3452
rect 3896 3447 3904 3932
rect 3936 3907 3944 4413
rect 3956 3947 3964 4213
rect 3976 4007 3984 4493
rect 3996 4427 4004 4813
rect 4016 4767 4024 5073
rect 4096 4967 4104 4993
rect 4096 4956 4112 4967
rect 4100 4953 4112 4956
rect 4036 4647 4044 4853
rect 4056 4747 4064 4853
rect 4076 4807 4084 4913
rect 4116 4847 4124 4893
rect 4156 4887 4164 5093
rect 4196 5067 4204 5173
rect 4236 5147 4244 5193
rect 4236 4987 4244 5033
rect 4176 4907 4184 4973
rect 4236 4927 4244 4973
rect 4036 4487 4044 4553
rect 4036 4476 4053 4487
rect 4040 4473 4053 4476
rect 4016 4207 4024 4333
rect 4007 4193 4024 4207
rect 4016 4147 4024 4193
rect 4056 3987 4064 4393
rect 4076 4107 4084 4793
rect 4096 4687 4104 4773
rect 4116 4227 4124 4833
rect 4136 4547 4144 4693
rect 4116 4144 4124 4173
rect 4116 4136 4144 4144
rect 3916 3707 3924 3893
rect 3896 3227 3904 3393
rect 3916 3067 3924 3593
rect 3896 2787 3904 3033
rect 3916 2907 3924 3053
rect 3936 2804 3944 3733
rect 3956 3227 3964 3433
rect 3976 2987 3984 3873
rect 3996 3727 4004 3853
rect 3996 3387 4004 3713
rect 4016 3527 4024 3973
rect 4096 3867 4104 4133
rect 4136 3847 4144 4136
rect 4156 4107 4164 4773
rect 4236 4667 4244 4913
rect 4276 4787 4284 5053
rect 4296 5027 4304 5133
rect 4296 4807 4304 4933
rect 4316 4784 4324 5753
rect 4736 5647 4744 5713
rect 4336 5207 4344 5633
rect 4436 5567 4444 5633
rect 4376 5287 4384 5553
rect 4416 5507 4424 5533
rect 4416 5447 4424 5493
rect 4456 5447 4464 5473
rect 4496 5407 4504 5493
rect 4616 5467 4624 5593
rect 4776 5527 4784 5653
rect 4796 5627 4804 5773
rect 4856 5647 4864 5824
rect 4936 5647 4944 5773
rect 4616 5456 4633 5467
rect 4620 5453 4633 5456
rect 4556 5327 4564 5453
rect 4736 5447 4744 5493
rect 4816 5467 4824 5533
rect 4616 5307 4624 5413
rect 4736 5387 4744 5433
rect 4340 5164 4354 5167
rect 4336 5153 4354 5164
rect 4336 4827 4344 5153
rect 4453 5124 4467 5133
rect 4436 5120 4467 5124
rect 4436 5116 4464 5120
rect 4396 5027 4404 5093
rect 4436 5067 4444 5116
rect 4396 4987 4404 5013
rect 4436 4907 4444 4933
rect 4296 4776 4324 4784
rect 4176 4507 4184 4653
rect 4296 4587 4304 4776
rect 4196 4128 4204 4573
rect 4216 4447 4224 4493
rect 4256 4247 4264 4513
rect 4316 4507 4324 4673
rect 4356 4587 4364 4633
rect 4306 4473 4307 4480
rect 4293 4467 4307 4473
rect 4293 4460 4314 4467
rect 4296 4453 4314 4460
rect 4040 3704 4053 3707
rect 4036 3693 4053 3704
rect 4036 3667 4044 3693
rect 4036 3407 4044 3493
rect 4020 3324 4033 3327
rect 4016 3313 4033 3324
rect 4016 3007 4024 3313
rect 4076 3127 4084 3333
rect 4096 3324 4104 3813
rect 4136 3807 4144 3833
rect 4176 3747 4184 3993
rect 4127 3724 4140 3727
rect 4127 3713 4144 3724
rect 4136 3647 4144 3713
rect 4156 3700 4164 3704
rect 4153 3687 4167 3700
rect 4156 3627 4164 3673
rect 4196 3667 4204 4092
rect 4236 3707 4244 3913
rect 4227 3696 4244 3707
rect 4227 3693 4240 3696
rect 4116 3387 4124 3533
rect 4176 3507 4184 3573
rect 4256 3527 4264 4233
rect 4296 4227 4304 4453
rect 4396 4387 4404 4893
rect 4476 4827 4484 4973
rect 4496 4967 4504 5173
rect 4596 5167 4604 5293
rect 4588 5156 4604 5167
rect 4588 5153 4600 5156
rect 4516 4987 4524 5013
rect 4556 4887 4564 4933
rect 4496 4807 4504 4833
rect 4496 4707 4504 4793
rect 4576 4787 4584 4973
rect 4576 4707 4584 4773
rect 4540 4684 4553 4687
rect 4536 4673 4553 4684
rect 4440 4664 4453 4667
rect 4436 4653 4453 4664
rect 4436 4527 4444 4653
rect 4436 4427 4444 4513
rect 4476 4387 4484 4633
rect 4296 3967 4304 4213
rect 4336 4127 4344 4373
rect 4376 4207 4384 4313
rect 4416 4147 4424 4193
rect 4276 3547 4284 3873
rect 4307 3704 4320 3707
rect 4307 3693 4324 3704
rect 4316 3587 4324 3693
rect 4356 3627 4364 3673
rect 4327 3524 4340 3527
rect 4327 3513 4344 3524
rect 4096 3316 4124 3324
rect 4096 3267 4104 3293
rect 4036 2987 4044 3013
rect 4096 3007 4104 3033
rect 4016 2827 4024 2913
rect 4076 2824 4084 2933
rect 4096 2847 4104 2953
rect 4116 2948 4124 3316
rect 4036 2816 4084 2824
rect 3936 2796 3964 2804
rect 3847 2736 3864 2747
rect 3847 2733 3860 2736
rect 3776 2667 3784 2733
rect 3836 2687 3844 2733
rect 3936 2707 3944 2753
rect 3847 2564 3860 2567
rect 3847 2553 3864 2564
rect 3907 2564 3920 2567
rect 3907 2553 3924 2564
rect 3736 2327 3744 2393
rect 3596 2147 3604 2273
rect 3616 2107 3624 2293
rect 3736 2287 3744 2313
rect 3576 2056 3593 2067
rect 3580 2053 3593 2056
rect 3516 1907 3524 2033
rect 3636 2027 3644 2213
rect 3696 2167 3704 2233
rect 3756 2187 3764 2413
rect 3656 2107 3664 2153
rect 3656 2096 3673 2107
rect 3660 2093 3673 2096
rect 3556 1907 3564 1993
rect 3416 1587 3424 1752
rect 3116 1307 3124 1453
rect 3156 1327 3164 1453
rect 3196 1327 3204 1353
rect 3166 1313 3167 1320
rect 3107 1296 3124 1307
rect 3153 1300 3167 1313
rect 3156 1296 3164 1300
rect 3107 1293 3120 1296
rect 3016 1107 3024 1133
rect 3036 984 3044 1153
rect 3056 1067 3064 1253
rect 3016 976 3044 984
rect 3016 847 3024 976
rect 3056 847 3064 1053
rect 3076 1047 3084 1073
rect 3096 887 3104 1133
rect 3116 1127 3124 1193
rect 3216 1187 3224 1493
rect 3156 907 3164 1073
rect 3193 1067 3207 1073
rect 3116 867 3124 893
rect 3176 847 3184 953
rect 3236 947 3244 1273
rect 3276 1167 3284 1353
rect 3316 1304 3324 1433
rect 3296 1296 3324 1304
rect 3296 1087 3304 1296
rect 3396 1287 3404 1453
rect 3416 1448 3424 1573
rect 3456 1447 3464 1732
rect 3496 1667 3504 1813
rect 3516 1627 3524 1713
rect 3513 1600 3527 1613
rect 3516 1596 3524 1600
rect 3487 1584 3500 1587
rect 3536 1584 3544 1873
rect 3576 1827 3584 2013
rect 3676 1887 3684 1953
rect 3716 1904 3724 2113
rect 3736 1907 3744 2033
rect 3696 1896 3724 1904
rect 3696 1847 3704 1896
rect 3776 1884 3784 2353
rect 3796 2087 3804 2533
rect 3816 2127 3824 2433
rect 3856 2387 3864 2553
rect 3916 2407 3924 2553
rect 3896 2327 3904 2353
rect 3856 2247 3864 2273
rect 3756 1876 3784 1884
rect 3487 1573 3504 1584
rect 3496 1547 3504 1573
rect 3516 1576 3544 1584
rect 3316 1207 3324 1273
rect 3336 1147 3344 1173
rect 3326 1133 3327 1140
rect 3313 1127 3327 1133
rect 3326 1120 3327 1127
rect 3333 1133 3334 1140
rect 3333 1120 3347 1133
rect 3336 1116 3344 1120
rect 3276 1076 3293 1084
rect 3276 927 3284 1076
rect 3276 904 3284 913
rect 3276 896 3304 904
rect 3296 867 3304 896
rect 3266 833 3267 840
rect 3253 824 3267 833
rect 3253 820 3284 824
rect 3256 816 3284 820
rect 2996 787 3004 813
rect 3156 747 3164 813
rect 2956 607 2964 633
rect 3016 627 3024 693
rect 3216 667 3224 753
rect 3007 616 3024 627
rect 3007 613 3020 616
rect 2816 187 2824 273
rect 2876 187 2884 473
rect 2916 367 2924 393
rect 2956 267 2964 353
rect 3016 347 3024 513
rect 3036 287 3044 333
rect 3056 327 3064 633
rect 3216 627 3224 653
rect 3076 467 3084 593
rect 3096 467 3104 493
rect 3116 347 3124 493
rect 2216 116 2232 127
rect 2220 113 2232 116
rect 2716 -24 2724 153
rect 2956 47 2964 133
rect 2996 27 3004 133
rect 3116 44 3124 333
rect 3136 247 3144 613
rect 3236 507 3244 733
rect 3276 687 3284 816
rect 3316 747 3324 853
rect 3336 707 3344 1013
rect 3376 867 3384 1213
rect 3416 867 3424 1412
rect 3456 1307 3464 1433
rect 3446 1293 3464 1307
rect 3456 1228 3464 1293
rect 3516 1207 3524 1576
rect 3436 827 3444 1093
rect 3456 807 3464 1192
rect 3356 747 3364 793
rect 3168 344 3180 347
rect 3168 333 3184 344
rect 3176 267 3184 333
rect 3236 167 3244 313
rect 3336 187 3344 653
rect 3167 164 3180 167
rect 3167 153 3184 164
rect 3096 40 3124 44
rect 3093 36 3124 40
rect 3093 27 3107 36
rect 3176 -24 3184 153
rect 3376 147 3384 793
rect 3396 207 3404 693
rect 3416 627 3424 713
rect 3456 627 3464 753
rect 3476 667 3484 1173
rect 3516 1107 3524 1153
rect 3508 1096 3524 1107
rect 3508 1093 3520 1096
rect 3496 848 3504 1093
rect 3536 927 3544 1493
rect 3556 947 3564 1553
rect 3576 867 3584 1733
rect 3596 847 3604 1553
rect 3636 1427 3644 1833
rect 3673 1807 3687 1813
rect 3716 1807 3724 1873
rect 3673 1800 3674 1807
rect 3756 1804 3764 1876
rect 3736 1800 3764 1804
rect 3733 1796 3764 1800
rect 3776 1807 3784 1853
rect 3816 1827 3824 2073
rect 3836 2067 3844 2193
rect 3896 2067 3904 2273
rect 3916 2267 3924 2313
rect 3936 2227 3944 2613
rect 3836 2056 3853 2067
rect 3840 2053 3853 2056
rect 3836 1967 3844 2032
rect 3916 1904 3924 2153
rect 3956 2087 3964 2796
rect 4016 2767 4024 2813
rect 3996 2388 4004 2533
rect 3976 2307 3984 2333
rect 3976 2127 3984 2153
rect 3996 2127 4004 2352
rect 4016 2167 4024 2453
rect 4036 2247 4044 2816
rect 4053 2787 4067 2793
rect 4068 2744 4080 2747
rect 4068 2733 4084 2744
rect 4056 2627 4064 2673
rect 4076 2587 4084 2733
rect 4096 2567 4104 2793
rect 4116 2767 4124 2912
rect 4136 2887 4144 3393
rect 4156 2887 4164 3473
rect 4256 3467 4264 3513
rect 4176 3007 4184 3253
rect 4236 3227 4244 3353
rect 4256 3307 4264 3453
rect 4336 3307 4344 3513
rect 4376 3367 4384 3893
rect 4396 3327 4404 4113
rect 4436 4104 4444 4373
rect 4496 4367 4504 4613
rect 4536 4607 4544 4673
rect 4536 4568 4544 4593
rect 4596 4587 4604 5093
rect 4636 5027 4644 5173
rect 4656 5147 4664 5373
rect 4696 5167 4704 5353
rect 4736 5107 4744 5273
rect 4716 5007 4724 5033
rect 4616 4647 4624 4993
rect 4776 4967 4784 5093
rect 4796 5088 4804 5153
rect 4796 5027 4804 5052
rect 4836 5047 4844 5553
rect 4856 5404 4864 5593
rect 4896 5487 4904 5633
rect 4976 5567 4984 5753
rect 5016 5727 5024 5824
rect 5056 5748 5064 5824
rect 5096 5767 5104 5824
rect 5236 5724 5244 5753
rect 5276 5747 5284 5824
rect 5276 5724 5284 5733
rect 5236 5716 5264 5724
rect 5276 5716 5324 5724
rect 5056 5627 5064 5712
rect 5076 5607 5084 5653
rect 5227 5644 5240 5647
rect 5227 5633 5244 5644
rect 5056 5467 5064 5533
rect 5096 5447 5104 5473
rect 4887 5425 4900 5427
rect 4887 5414 4904 5425
rect 4880 5413 4904 5414
rect 4856 5396 4873 5404
rect 4856 5327 4864 5353
rect 4876 5307 4884 5392
rect 4896 5347 4904 5413
rect 4936 5347 4944 5413
rect 5036 5387 5044 5413
rect 4876 5224 4884 5293
rect 4876 5216 4904 5224
rect 4896 5147 4904 5216
rect 5036 5187 5044 5373
rect 5096 5187 5104 5313
rect 4987 5164 5000 5167
rect 4987 5153 5004 5164
rect 4896 5136 4913 5147
rect 4900 5133 4913 5136
rect 4776 4956 4793 4967
rect 4780 4953 4793 4956
rect 4856 4947 4864 5053
rect 4647 4924 4660 4927
rect 4693 4924 4707 4933
rect 4647 4913 4664 4924
rect 4693 4920 4724 4924
rect 4696 4916 4724 4920
rect 4656 4827 4664 4913
rect 4636 4564 4644 4673
rect 4696 4627 4704 4653
rect 4616 4556 4644 4564
rect 4536 4447 4544 4532
rect 4616 4487 4624 4556
rect 4580 4464 4593 4467
rect 4576 4453 4593 4464
rect 4576 4367 4584 4453
rect 4556 4207 4564 4313
rect 4527 4184 4540 4187
rect 4596 4184 4604 4413
rect 4616 4304 4624 4473
rect 4636 4327 4644 4453
rect 4676 4347 4684 4553
rect 4696 4547 4704 4613
rect 4696 4367 4704 4473
rect 4716 4447 4724 4916
rect 4736 4847 4744 4933
rect 4876 4807 4884 5113
rect 4996 5107 5004 5153
rect 5016 5140 5024 5144
rect 5013 5127 5027 5140
rect 5016 5087 5024 5113
rect 5056 4907 5064 5093
rect 5096 4887 5104 5033
rect 5036 4787 5044 4873
rect 4736 4567 4744 4773
rect 4967 4704 4980 4707
rect 4967 4693 4984 4704
rect 4833 4664 4847 4673
rect 4833 4660 4893 4664
rect 4836 4656 4893 4660
rect 4760 4604 4773 4607
rect 4756 4593 4773 4604
rect 4756 4547 4764 4593
rect 4796 4567 4804 4633
rect 4736 4327 4744 4473
rect 4616 4296 4644 4304
rect 4636 4247 4644 4296
rect 4527 4173 4544 4184
rect 4596 4176 4624 4184
rect 4416 4096 4444 4104
rect 4416 3427 4424 4096
rect 4536 4067 4544 4173
rect 4616 4047 4624 4176
rect 4756 4184 4764 4433
rect 4796 4367 4804 4553
rect 4836 4527 4844 4593
rect 4976 4527 4984 4693
rect 4876 4327 4884 4473
rect 4913 4427 4927 4433
rect 4748 4176 4764 4184
rect 4493 4027 4507 4033
rect 4553 4024 4567 4033
rect 4553 4020 4584 4024
rect 4556 4016 4584 4020
rect 4456 3707 4464 3953
rect 4476 3887 4484 3933
rect 4516 3927 4524 3953
rect 4467 3704 4480 3707
rect 4467 3693 4484 3704
rect 4436 3567 4444 3613
rect 4476 3607 4484 3693
rect 4256 3247 4264 3293
rect 4296 3227 4304 3273
rect 4376 3247 4384 3293
rect 4376 3236 4393 3247
rect 4380 3233 4393 3236
rect 4296 3216 4313 3227
rect 4300 3213 4313 3216
rect 4416 3224 4424 3313
rect 4396 3216 4424 3224
rect 4236 3007 4244 3073
rect 4256 3027 4264 3073
rect 4256 2987 4264 3013
rect 4176 2784 4184 2953
rect 4296 2927 4304 3153
rect 4316 3027 4324 3173
rect 4376 3087 4384 3193
rect 4316 2907 4324 3013
rect 4356 2944 4364 3053
rect 4336 2936 4364 2944
rect 4256 2787 4264 2893
rect 4156 2776 4184 2784
rect 4136 2567 4144 2713
rect 4056 2424 4064 2553
rect 4056 2416 4084 2424
rect 4076 2327 4084 2416
rect 4096 2367 4104 2473
rect 4136 2367 4144 2493
rect 4156 2487 4164 2776
rect 4176 2707 4184 2733
rect 4196 2667 4204 2753
rect 4256 2687 4264 2773
rect 4336 2767 4344 2936
rect 4376 2927 4384 3073
rect 4276 2687 4284 2713
rect 4276 2604 4284 2673
rect 4256 2596 4284 2604
rect 4176 2547 4184 2593
rect 4256 2567 4264 2596
rect 4248 2553 4264 2567
rect 4176 2536 4193 2547
rect 4180 2533 4193 2536
rect 4176 2364 4184 2433
rect 4256 2427 4264 2553
rect 4296 2547 4304 2633
rect 4276 2536 4292 2544
rect 4276 2507 4284 2536
rect 4316 2527 4324 2653
rect 4316 2447 4324 2513
rect 4176 2356 4204 2364
rect 4113 2307 4127 2313
rect 4156 2287 4164 2333
rect 4196 2327 4204 2356
rect 4156 2276 4173 2287
rect 4160 2273 4173 2276
rect 3933 2044 3947 2053
rect 3933 2040 3964 2044
rect 3936 2036 3964 2040
rect 3907 1896 3924 1904
rect 3896 1847 3904 1893
rect 3776 1796 3794 1807
rect 3733 1787 3747 1796
rect 3780 1793 3794 1796
rect 3776 1707 3784 1773
rect 3656 1567 3664 1673
rect 3796 1627 3804 1673
rect 3656 1556 3673 1567
rect 3660 1553 3673 1556
rect 3616 1167 3624 1353
rect 3707 1304 3720 1307
rect 3707 1293 3724 1304
rect 3616 1007 3624 1113
rect 3656 1024 3664 1073
rect 3656 1020 3684 1024
rect 3656 1016 3687 1020
rect 3673 1007 3687 1016
rect 3673 1000 3674 1007
rect 3500 824 3512 827
rect 3496 813 3512 824
rect 3496 747 3504 813
rect 3416 616 3432 627
rect 3420 613 3432 616
rect 3456 407 3464 613
rect 3416 367 3424 393
rect 3473 364 3487 373
rect 3496 364 3504 633
rect 3473 360 3504 364
rect 3476 356 3504 360
rect 3516 347 3524 753
rect 3556 667 3564 773
rect 3596 687 3604 833
rect 3596 647 3604 673
rect 3586 593 3587 600
rect 3573 587 3587 593
rect 3596 347 3604 593
rect 3636 467 3644 613
rect 3656 607 3664 993
rect 3696 867 3704 1253
rect 3716 1227 3724 1293
rect 3756 1287 3764 1613
rect 3836 1587 3844 1753
rect 3876 1644 3884 1813
rect 3928 1804 3940 1807
rect 3928 1793 3944 1804
rect 3896 1667 3904 1773
rect 3936 1748 3944 1793
rect 3876 1636 3904 1644
rect 3796 1327 3804 1473
rect 3756 1127 3764 1193
rect 3856 1127 3864 1293
rect 3876 1144 3884 1613
rect 3896 1367 3904 1636
rect 3916 1247 3924 1313
rect 3876 1136 3904 1144
rect 3747 1116 3764 1127
rect 3747 1113 3760 1116
rect 3867 1116 3884 1124
rect 3756 987 3764 1092
rect 3696 684 3704 853
rect 3696 676 3724 684
rect 3676 587 3684 653
rect 3716 427 3724 676
rect 3736 667 3744 913
rect 3796 827 3804 953
rect 3796 487 3804 813
rect 3836 707 3844 933
rect 3876 867 3884 1116
rect 3456 340 3464 344
rect 3453 327 3467 340
rect 3707 344 3720 347
rect 3707 333 3724 344
rect 3456 47 3464 313
rect 3636 187 3644 333
rect 3513 87 3527 93
rect 3596 -24 3604 173
rect 3627 124 3640 127
rect 3627 113 3644 124
rect 3636 88 3644 113
rect 3636 -24 3644 52
rect 3716 -24 3724 333
rect 3756 327 3764 453
rect 3796 147 3804 373
rect 3836 367 3844 693
rect 3876 147 3884 753
rect 3896 467 3904 1136
rect 3936 1104 3944 1712
rect 3956 1687 3964 2036
rect 3976 1704 3984 2013
rect 3996 1727 4004 1973
rect 4016 1947 4024 2093
rect 4036 2067 4044 2193
rect 4056 2107 4064 2153
rect 4076 2067 4084 2213
rect 4036 2007 4044 2053
rect 4036 1787 4044 1873
rect 4096 1847 4104 2233
rect 4116 1988 4124 2173
rect 4156 2147 4164 2173
rect 4106 1773 4107 1780
rect 4093 1767 4107 1773
rect 3976 1696 4004 1704
rect 3996 1644 4004 1696
rect 3956 1636 4004 1644
rect 3956 1387 3964 1636
rect 4036 1627 4044 1693
rect 3987 1604 4000 1607
rect 3987 1593 4004 1604
rect 3996 1447 4004 1593
rect 3976 1307 3984 1353
rect 4016 1284 4024 1373
rect 3996 1276 4024 1284
rect 3996 1204 4004 1276
rect 4036 1267 4044 1433
rect 4096 1427 4104 1533
rect 3976 1196 4004 1204
rect 3976 1127 3984 1196
rect 3936 1096 3964 1104
rect 3916 847 3924 893
rect 3956 827 3964 1096
rect 3976 844 3984 1073
rect 3996 887 4004 1133
rect 4036 1007 4044 1133
rect 4080 1124 4093 1127
rect 4076 1113 4093 1124
rect 4076 1087 4084 1113
rect 4116 1107 4124 1952
rect 4156 1887 4164 2033
rect 4176 2008 4184 2073
rect 4196 2047 4204 2213
rect 4136 1787 4144 1813
rect 4148 1776 4164 1784
rect 4136 1587 4144 1713
rect 4156 1547 4164 1776
rect 4136 1347 4144 1393
rect 4136 1307 4144 1333
rect 4116 1096 4133 1107
rect 4120 1093 4133 1096
rect 4156 987 4164 1493
rect 4176 1447 4184 1972
rect 4196 1607 4204 1793
rect 4216 1648 4224 2333
rect 4236 1827 4244 2313
rect 4256 2087 4264 2253
rect 4246 1773 4247 1780
rect 4233 1767 4247 1773
rect 4256 1627 4264 2013
rect 4276 1967 4284 2393
rect 4296 2147 4304 2373
rect 4356 2347 4364 2913
rect 4376 2387 4384 2873
rect 4396 2827 4404 3216
rect 4436 3187 4444 3553
rect 4467 3484 4480 3487
rect 4467 3473 4484 3484
rect 4476 3448 4484 3473
rect 4476 3267 4484 3412
rect 4496 3167 4504 3873
rect 4516 3187 4524 3833
rect 4576 3727 4584 4016
rect 4676 3967 4684 4173
rect 4736 4087 4744 4173
rect 4616 3847 4624 3953
rect 4547 3704 4560 3707
rect 4547 3693 4564 3704
rect 4556 3587 4564 3693
rect 4536 3307 4544 3513
rect 4616 3507 4624 3833
rect 4716 3827 4724 3993
rect 4736 3907 4744 4033
rect 4756 3707 4764 4053
rect 4796 4047 4804 4233
rect 4856 4027 4864 4093
rect 4876 4007 4884 4153
rect 4916 4067 4924 4153
rect 4976 4067 4984 4513
rect 5016 4347 5024 4433
rect 5036 4427 5044 4453
rect 5036 4187 5044 4313
rect 4816 3827 4824 3993
rect 4836 3927 4844 3973
rect 4707 3704 4720 3707
rect 4707 3693 4724 3704
rect 4756 3696 4773 3707
rect 4760 3693 4773 3696
rect 4716 3627 4724 3693
rect 4776 3647 4784 3693
rect 4607 3493 4624 3507
rect 4616 3467 4624 3493
rect 4736 3487 4744 3533
rect 4727 3473 4744 3487
rect 4576 3387 4584 3433
rect 4736 3407 4744 3473
rect 4536 3207 4544 3253
rect 4416 3027 4424 3133
rect 4536 3107 4544 3193
rect 4436 3047 4444 3093
rect 4436 2987 4444 3033
rect 4480 3004 4492 3007
rect 4476 2993 4492 3004
rect 4476 2947 4484 2993
rect 4516 2924 4524 3073
rect 4556 3027 4564 3233
rect 4576 3048 4584 3373
rect 4596 3087 4604 3313
rect 4616 3087 4624 3353
rect 4736 3307 4744 3393
rect 4756 3367 4764 3613
rect 4796 3527 4804 3613
rect 4816 3607 4824 3693
rect 4636 3247 4644 3293
rect 4756 3267 4764 3353
rect 4796 3247 4804 3273
rect 4556 3026 4580 3027
rect 4556 3015 4573 3026
rect 4560 3013 4573 3015
rect 4656 2967 4664 3193
rect 4736 3147 4744 3233
rect 4496 2916 4524 2924
rect 4416 2744 4424 2873
rect 4396 2736 4424 2744
rect 4396 2627 4404 2736
rect 4416 2587 4424 2713
rect 4416 2507 4424 2533
rect 4436 2487 4444 2633
rect 4456 2588 4464 2793
rect 4476 2564 4484 2893
rect 4467 2556 4484 2564
rect 4416 2327 4424 2353
rect 4316 2267 4324 2293
rect 4327 2084 4340 2087
rect 4327 2073 4344 2084
rect 4336 2027 4344 2073
rect 4356 2067 4364 2293
rect 4416 2087 4424 2313
rect 4436 2128 4444 2333
rect 4456 2168 4464 2552
rect 4216 1587 4224 1612
rect 4216 1327 4224 1533
rect 4276 1507 4284 1833
rect 4276 1367 4284 1433
rect 4216 1107 4224 1213
rect 4236 1087 4244 1333
rect 4276 1307 4284 1353
rect 4296 1167 4304 1973
rect 4316 1644 4324 1993
rect 4340 1804 4353 1807
rect 4336 1793 4353 1804
rect 4336 1667 4344 1793
rect 4376 1787 4384 2033
rect 4436 1987 4444 2092
rect 4396 1804 4404 1953
rect 4416 1887 4424 1933
rect 4396 1796 4413 1804
rect 4316 1636 4344 1644
rect 4316 1587 4324 1613
rect 4336 1567 4344 1636
rect 4316 1287 4324 1473
rect 4336 1447 4344 1553
rect 4356 1467 4364 1753
rect 4376 1707 4384 1773
rect 4396 1487 4404 1613
rect 4376 1347 4384 1413
rect 4367 1336 4384 1347
rect 4367 1333 4380 1336
rect 4356 1147 4364 1333
rect 4416 1307 4424 1793
rect 4436 1507 4444 1773
rect 4456 1627 4464 2132
rect 4476 2087 4484 2493
rect 4496 2487 4504 2916
rect 4516 2807 4524 2893
rect 4516 2307 4524 2433
rect 4536 2407 4544 2733
rect 4556 2507 4564 2933
rect 4576 2647 4584 2773
rect 4656 2767 4664 2853
rect 4648 2756 4664 2767
rect 4648 2753 4660 2756
rect 4616 2704 4624 2733
rect 4596 2700 4624 2704
rect 4593 2696 4624 2700
rect 4593 2687 4607 2696
rect 4636 2687 4644 2753
rect 4676 2747 4684 2793
rect 4696 2667 4704 3013
rect 4576 2547 4584 2593
rect 4556 2307 4564 2333
rect 4513 2284 4527 2293
rect 4496 2280 4527 2284
rect 4496 2276 4524 2280
rect 4496 2207 4504 2276
rect 4520 2266 4540 2267
rect 4528 2264 4540 2266
rect 4528 2253 4544 2264
rect 4496 2067 4504 2113
rect 4536 2067 4544 2253
rect 4556 2167 4564 2213
rect 4576 2127 4584 2233
rect 4567 2084 4580 2087
rect 4567 2073 4584 2084
rect 4476 1787 4484 1993
rect 4496 1827 4504 2053
rect 4576 2027 4584 2073
rect 4596 2007 4604 2613
rect 4696 2527 4704 2553
rect 4616 2367 4624 2513
rect 4716 2507 4724 3073
rect 4776 3067 4784 3213
rect 4773 3040 4787 3053
rect 4776 3036 4784 3040
rect 4756 2968 4764 2993
rect 4776 2987 4784 3012
rect 4736 2747 4744 2853
rect 4736 2567 4744 2693
rect 4756 2667 4764 2932
rect 4796 2907 4804 3173
rect 4816 2827 4824 3293
rect 4800 2764 4813 2767
rect 4796 2753 4813 2764
rect 4796 2727 4804 2753
rect 4776 2716 4793 2724
rect 4776 2547 4784 2716
rect 4796 2587 4804 2673
rect 4796 2576 4813 2587
rect 4800 2573 4813 2576
rect 4616 2147 4624 2293
rect 4496 1687 4504 1773
rect 4516 1747 4524 1793
rect 4536 1727 4544 1973
rect 4536 1627 4544 1653
rect 4456 1347 4464 1573
rect 4476 1407 4484 1553
rect 4273 1073 4274 1080
rect 4036 887 4044 953
rect 3976 836 4004 844
rect 3956 747 3964 813
rect 3996 727 4004 836
rect 3896 367 3904 413
rect 3896 356 3913 367
rect 3900 353 3913 356
rect 3936 167 3944 713
rect 3956 627 3964 653
rect 3976 647 3984 673
rect 3976 636 3993 647
rect 3980 633 3993 636
rect 4016 387 4024 553
rect 3956 147 3964 333
rect 4036 327 4044 793
rect 4056 627 4064 833
rect 4027 164 4040 167
rect 4027 153 4044 164
rect 3786 113 3787 120
rect 3773 107 3787 113
rect 4036 -24 4044 153
rect 4076 47 4084 973
rect 4096 167 4104 913
rect 4116 887 4124 933
rect 4176 927 4184 1033
rect 4160 864 4173 867
rect 4156 853 4173 864
rect 4156 807 4164 853
rect 4196 847 4204 1073
rect 4236 1047 4244 1073
rect 4273 1067 4287 1073
rect 4316 1047 4324 1073
rect 4236 847 4244 873
rect 4280 824 4293 827
rect 4276 813 4293 824
rect 4276 707 4284 813
rect 4176 647 4184 693
rect 4276 667 4284 693
rect 4316 688 4324 973
rect 4336 967 4344 1093
rect 4376 987 4384 1273
rect 4476 1047 4484 1313
rect 4496 1007 4504 1533
rect 4556 1287 4564 1913
rect 4636 1867 4644 2473
rect 4676 2347 4684 2433
rect 4660 2284 4672 2287
rect 4656 2274 4672 2284
rect 4656 2273 4680 2274
rect 4656 2227 4664 2273
rect 4696 2264 4704 2393
rect 4716 2347 4724 2413
rect 4716 2307 4724 2333
rect 4676 2260 4704 2264
rect 4673 2256 4704 2260
rect 4673 2247 4687 2256
rect 4656 2147 4664 2213
rect 4676 2047 4684 2153
rect 4716 2127 4724 2293
rect 4736 2084 4744 2473
rect 4756 2107 4764 2493
rect 4736 2076 4764 2084
rect 4520 1284 4532 1287
rect 4516 1273 4532 1284
rect 4356 807 4364 833
rect 4376 727 4384 933
rect 4167 633 4184 647
rect 4176 447 4184 633
rect 4216 407 4224 613
rect 4316 607 4324 652
rect 4396 647 4404 833
rect 4416 807 4424 953
rect 4516 927 4524 1273
rect 4576 1268 4584 1833
rect 4596 1787 4604 1813
rect 4596 1776 4613 1787
rect 4600 1773 4613 1776
rect 4596 1448 4604 1713
rect 4616 1424 4624 1693
rect 4636 1688 4644 1753
rect 4636 1587 4644 1652
rect 4656 1467 4664 2013
rect 4676 1887 4684 1993
rect 4676 1767 4684 1793
rect 4696 1704 4704 1853
rect 4716 1728 4724 2073
rect 4676 1696 4704 1704
rect 4676 1567 4684 1696
rect 4716 1667 4724 1692
rect 4736 1567 4744 1773
rect 4607 1416 4624 1424
rect 4596 1307 4604 1412
rect 4636 1347 4644 1373
rect 4648 1304 4660 1307
rect 4648 1293 4664 1304
rect 4656 1287 4664 1293
rect 4508 844 4520 847
rect 4508 833 4524 844
rect 4456 787 4464 833
rect 4436 667 4444 733
rect 4396 636 4412 647
rect 4400 633 4412 636
rect 4476 467 4484 733
rect 4516 707 4524 833
rect 4536 747 4544 1153
rect 4576 1107 4584 1232
rect 4616 1227 4624 1273
rect 4656 1147 4664 1273
rect 4676 1187 4684 1493
rect 4567 1096 4584 1107
rect 4567 1093 4580 1096
rect 4596 1087 4604 1133
rect 4636 807 4644 1093
rect 4696 1087 4704 1433
rect 4716 1327 4724 1473
rect 4756 1247 4764 2076
rect 4776 1927 4784 2413
rect 4836 2367 4844 3633
rect 4856 3307 4864 3893
rect 4880 3684 4893 3687
rect 4876 3673 4893 3684
rect 4876 3367 4884 3673
rect 4916 3647 4924 4053
rect 5016 3967 5024 4173
rect 5036 4087 5044 4173
rect 4936 3684 4944 3953
rect 4976 3767 4984 3833
rect 4976 3728 4984 3753
rect 4967 3704 4980 3707
rect 4967 3693 4984 3704
rect 4936 3676 4964 3684
rect 4916 3527 4924 3633
rect 4936 3547 4944 3613
rect 4907 3516 4924 3527
rect 4907 3513 4920 3516
rect 4936 3327 4944 3353
rect 4936 3247 4944 3313
rect 4856 3007 4864 3153
rect 4876 3027 4884 3093
rect 4916 2948 4924 3073
rect 4876 2787 4884 2893
rect 4916 2847 4924 2912
rect 4936 2867 4944 2993
rect 4956 2927 4964 3676
rect 4976 3407 4984 3693
rect 4996 3607 5004 3693
rect 5036 3667 5044 4073
rect 5056 3607 5064 4513
rect 5076 4467 5084 4693
rect 5076 3587 5084 4333
rect 5096 3867 5104 4633
rect 5116 4567 5124 5513
rect 5136 5387 5144 5473
rect 5156 5447 5164 5633
rect 5236 5507 5244 5633
rect 5256 5627 5264 5716
rect 5266 5613 5267 5620
rect 5253 5600 5267 5613
rect 5256 5596 5264 5600
rect 5253 5467 5267 5473
rect 5253 5460 5254 5467
rect 5156 5436 5173 5447
rect 5160 5433 5173 5436
rect 5216 5367 5224 5453
rect 5136 5167 5144 5233
rect 5256 5127 5264 5413
rect 5276 5104 5284 5613
rect 5316 5604 5324 5716
rect 5316 5596 5344 5604
rect 5256 5096 5284 5104
rect 5156 4987 5164 5053
rect 5136 4247 5144 4853
rect 5196 4667 5204 4933
rect 5187 4656 5204 4667
rect 5187 4653 5200 4656
rect 5176 4587 5184 4613
rect 5156 4464 5164 4493
rect 5176 4487 5184 4573
rect 5216 4527 5224 5013
rect 5256 4647 5264 5096
rect 5296 5027 5304 5493
rect 5336 5007 5344 5596
rect 5356 5447 5364 5533
rect 5376 5527 5384 5593
rect 5396 4984 5404 5613
rect 5416 5467 5424 5473
rect 5413 5440 5427 5453
rect 5416 5436 5424 5440
rect 5416 5087 5424 5393
rect 5436 5327 5444 5773
rect 5436 5167 5444 5273
rect 5376 4976 5404 4984
rect 5208 4484 5220 4487
rect 5208 4473 5224 4484
rect 5156 4456 5184 4464
rect 5176 4187 5184 4456
rect 5216 4267 5224 4473
rect 5256 4307 5264 4453
rect 5276 4327 5284 4653
rect 5316 4627 5324 4953
rect 5376 4868 5384 4976
rect 5416 4967 5424 5073
rect 5400 4964 5413 4967
rect 5396 4953 5413 4964
rect 5396 4927 5404 4953
rect 5476 4947 5484 5824
rect 5516 5487 5524 5824
rect 5556 5767 5564 5824
rect 5536 5647 5544 5733
rect 5580 5624 5593 5627
rect 5576 5613 5593 5624
rect 5576 5507 5584 5613
rect 5496 5227 5504 5433
rect 5556 5327 5564 5413
rect 5596 5347 5604 5453
rect 5376 4687 5384 4832
rect 5376 4676 5393 4687
rect 5380 4673 5393 4676
rect 5436 4647 5444 4933
rect 5496 4927 5504 5113
rect 5493 4913 5494 4920
rect 5493 4907 5507 4913
rect 5336 4567 5344 4593
rect 5336 4487 5344 4553
rect 5327 4476 5344 4487
rect 5327 4473 5340 4476
rect 5376 4467 5384 4553
rect 5216 4227 5224 4253
rect 5373 4247 5387 4253
rect 5256 4184 5264 4233
rect 5236 4180 5264 4184
rect 5233 4176 5264 4180
rect 5136 4007 5144 4173
rect 5136 3967 5144 3993
rect 5096 3787 5104 3853
rect 5096 3687 5104 3733
rect 5156 3664 5164 4053
rect 5136 3656 5164 3664
rect 5036 3387 5044 3493
rect 4973 3267 4987 3273
rect 5056 3227 5064 3533
rect 5076 3247 5084 3433
rect 5056 3147 5064 3213
rect 4996 3027 5004 3133
rect 4988 3016 5004 3027
rect 4988 3013 5000 3016
rect 4976 2987 4984 3013
rect 5016 2984 5024 3113
rect 5076 3007 5084 3193
rect 5096 2987 5104 3273
rect 5116 3187 5124 3653
rect 5136 3167 5144 3656
rect 5176 3644 5184 4173
rect 5233 4167 5247 4176
rect 5196 3847 5204 3993
rect 5247 3964 5260 3967
rect 5247 3953 5264 3964
rect 5256 3927 5264 3953
rect 5256 3827 5264 3913
rect 5296 3867 5304 4213
rect 5396 4147 5404 4613
rect 5476 4487 5484 4833
rect 5516 4827 5524 5153
rect 5556 5047 5564 5313
rect 5636 5167 5644 5413
rect 5676 5407 5684 5533
rect 5593 5087 5607 5093
rect 5556 4687 5564 4973
rect 5596 4887 5604 4913
rect 5516 4587 5524 4653
rect 5556 4487 5564 4553
rect 5556 4476 5573 4487
rect 5560 4473 5573 4476
rect 5376 3987 5384 4013
rect 5416 4007 5424 4353
rect 5436 4167 5444 4413
rect 5456 4227 5464 4453
rect 5476 4207 5484 4433
rect 5616 4427 5624 4893
rect 5636 4667 5644 4873
rect 5413 3987 5427 3993
rect 5413 3980 5414 3987
rect 5156 3636 5184 3644
rect 5156 3347 5164 3636
rect 5196 3544 5204 3773
rect 5216 3727 5224 3813
rect 5316 3707 5324 3813
rect 5436 3707 5444 3833
rect 5307 3696 5324 3707
rect 5307 3693 5320 3696
rect 5428 3696 5444 3707
rect 5428 3693 5440 3696
rect 5176 3536 5204 3544
rect 5156 3207 5164 3253
rect 5116 3027 5124 3093
rect 5016 2976 5044 2984
rect 4876 2747 4884 2773
rect 4856 2647 4864 2693
rect 4856 2527 4864 2633
rect 4876 2447 4884 2653
rect 4896 2507 4904 2813
rect 4976 2807 4984 2933
rect 4996 2887 5004 2913
rect 5036 2827 5044 2976
rect 4976 2747 4984 2793
rect 5053 2773 5054 2780
rect 5053 2767 5067 2773
rect 5046 2760 5067 2767
rect 5046 2756 5064 2760
rect 5046 2753 5060 2756
rect 4836 2287 4844 2313
rect 4876 2307 4884 2433
rect 4826 2273 4827 2280
rect 4836 2276 4853 2287
rect 4840 2273 4853 2276
rect 4813 2267 4827 2273
rect 4816 2147 4824 2253
rect 4816 2047 4824 2093
rect 4836 2087 4844 2233
rect 4876 2167 4884 2293
rect 4916 2227 4924 2273
rect 4866 2153 4867 2160
rect 4853 2144 4867 2153
rect 4853 2140 4884 2144
rect 4856 2136 4884 2140
rect 4876 2047 4884 2136
rect 4916 2047 4924 2153
rect 4776 1787 4784 1853
rect 4796 1848 4804 1913
rect 4776 1627 4784 1713
rect 4796 1687 4804 1812
rect 4816 1787 4824 1893
rect 4796 1607 4804 1673
rect 4856 1667 4864 1973
rect 4896 1907 4904 1933
rect 4936 1887 4944 2353
rect 4956 2247 4964 2653
rect 4976 2307 4984 2493
rect 4976 2127 4984 2253
rect 4996 2187 5004 2673
rect 5016 2267 5024 2733
rect 5076 2627 5084 2873
rect 5096 2507 5104 2693
rect 5116 2567 5124 2973
rect 5136 2867 5144 2993
rect 5156 2988 5164 3133
rect 5156 2667 5164 2952
rect 5176 2867 5184 3536
rect 5196 3387 5204 3513
rect 5216 3327 5224 3593
rect 5236 3547 5244 3653
rect 5376 3627 5384 3693
rect 5236 3507 5244 3533
rect 5256 3487 5264 3513
rect 5196 3067 5204 3213
rect 5196 2844 5204 3013
rect 5236 2967 5244 3293
rect 5256 3107 5264 3313
rect 5296 3267 5304 3393
rect 5256 3004 5264 3093
rect 5296 3067 5304 3213
rect 5296 3027 5304 3053
rect 5287 3016 5304 3027
rect 5287 3013 5300 3016
rect 5316 3007 5324 3053
rect 5336 3047 5344 3233
rect 5356 3067 5364 3193
rect 5256 3000 5284 3004
rect 5256 2996 5287 3000
rect 5273 2987 5287 2996
rect 5216 2847 5224 2893
rect 5176 2836 5204 2844
rect 5176 2767 5184 2836
rect 5196 2747 5204 2793
rect 5216 2767 5224 2833
rect 5156 2467 5164 2513
rect 5036 2267 5044 2313
rect 4916 1847 4924 1873
rect 4956 1844 4964 2073
rect 4996 2004 5004 2173
rect 4976 1996 5004 2004
rect 4976 1947 4984 1996
rect 5036 1987 5044 2213
rect 5056 2067 5064 2393
rect 5156 2287 5164 2373
rect 5136 2276 5153 2284
rect 5088 2264 5100 2267
rect 5088 2254 5104 2264
rect 5080 2253 5104 2254
rect 4936 1840 4964 1844
rect 4933 1836 4964 1840
rect 4916 1807 4924 1833
rect 4933 1827 4947 1836
rect 4976 1807 4984 1933
rect 5076 1927 5084 2232
rect 5096 2127 5104 2253
rect 5136 2207 5144 2276
rect 5176 2227 5184 2653
rect 5196 2347 5204 2693
rect 5256 2667 5264 2873
rect 5216 2407 5224 2553
rect 5276 2427 5284 2573
rect 5136 2067 5144 2153
rect 5176 2028 5184 2073
rect 5156 2016 5173 2024
rect 5136 1907 5144 1993
rect 4976 1796 4993 1807
rect 4980 1793 4993 1796
rect 4776 1527 4784 1573
rect 4816 1547 4824 1573
rect 4796 1387 4804 1513
rect 4796 1328 4804 1373
rect 4836 1367 4844 1613
rect 4856 1427 4864 1653
rect 4916 1447 4924 1753
rect 4956 1667 4964 1713
rect 4996 1707 5004 1793
rect 4956 1627 4964 1653
rect 4973 1593 4974 1600
rect 4973 1587 4987 1593
rect 4966 1580 4987 1587
rect 4966 1573 4984 1580
rect 4936 1427 4944 1473
rect 4800 1304 4813 1307
rect 4796 1293 4813 1304
rect 4676 827 4684 933
rect 4716 907 4724 1053
rect 4796 967 4804 1293
rect 4836 1287 4844 1313
rect 4836 967 4844 1073
rect 4856 927 4864 1173
rect 4876 1147 4884 1353
rect 4896 1307 4904 1373
rect 4936 1307 4944 1413
rect 4956 1407 4964 1453
rect 4976 1367 4984 1573
rect 5016 1427 5024 1813
rect 5056 1747 5064 1813
rect 5093 1804 5107 1813
rect 5076 1800 5107 1804
rect 5076 1796 5104 1800
rect 5076 1767 5084 1796
rect 5036 1736 5053 1744
rect 5036 1687 5044 1736
rect 5036 1607 5044 1673
rect 5096 1584 5104 1772
rect 5076 1576 5104 1584
rect 5056 1384 5064 1473
rect 5036 1376 5064 1384
rect 4876 1047 4884 1093
rect 4896 1024 4904 1233
rect 4876 1016 4904 1024
rect 4716 896 4733 907
rect 4720 893 4733 896
rect 4796 867 4804 893
rect 4787 856 4804 867
rect 4787 853 4800 856
rect 4816 847 4824 913
rect 4876 907 4884 1016
rect 4916 867 4924 1253
rect 4816 836 4833 847
rect 4820 833 4833 836
rect 4936 844 4944 1213
rect 4956 1207 4964 1313
rect 5016 1268 5024 1333
rect 4996 1167 5004 1213
rect 5016 1147 5024 1232
rect 4960 1124 4973 1127
rect 4956 1113 4973 1124
rect 4956 887 4964 1113
rect 5036 1047 5044 1376
rect 5076 1367 5084 1576
rect 5116 1564 5124 1873
rect 5136 1828 5144 1893
rect 5136 1747 5144 1792
rect 5156 1748 5164 2016
rect 5216 2007 5224 2293
rect 5296 2287 5304 2933
rect 5356 2887 5364 3013
rect 5376 2827 5384 3473
rect 5396 2907 5404 3153
rect 5416 2807 5424 3193
rect 5436 3027 5444 3253
rect 5456 3127 5464 4113
rect 5476 3487 5484 3873
rect 5496 3687 5504 4153
rect 5516 4027 5524 4193
rect 5516 3267 5524 3533
rect 5536 3467 5544 4133
rect 5556 3427 5564 4193
rect 5476 3147 5484 3233
rect 5536 3207 5544 3353
rect 5576 3307 5584 4153
rect 5596 3987 5604 4293
rect 5636 4184 5644 4653
rect 5656 4367 5664 5373
rect 5616 4176 5644 4184
rect 5616 4127 5624 4176
rect 5636 4067 5644 4153
rect 5656 4067 5664 4193
rect 5596 3487 5604 3753
rect 5596 3347 5604 3473
rect 5596 3227 5604 3333
rect 5476 3007 5484 3053
rect 5516 3044 5524 3153
rect 5556 3067 5564 3133
rect 5596 3107 5604 3213
rect 5616 3167 5624 3393
rect 5547 3056 5564 3067
rect 5547 3053 5560 3056
rect 5516 3036 5544 3044
rect 5516 2807 5524 3013
rect 5536 2947 5544 3036
rect 5316 2667 5324 2773
rect 5356 2747 5364 2773
rect 5400 2764 5413 2767
rect 5396 2753 5413 2764
rect 5356 2704 5364 2733
rect 5336 2696 5364 2704
rect 5336 2588 5344 2696
rect 5356 2607 5364 2673
rect 5396 2647 5404 2753
rect 5456 2687 5464 2753
rect 5340 2564 5353 2567
rect 5336 2553 5353 2564
rect 5316 2387 5324 2453
rect 5336 2447 5344 2553
rect 5436 2544 5444 2573
rect 5416 2536 5444 2544
rect 5416 2527 5424 2536
rect 5407 2516 5424 2527
rect 5407 2513 5420 2516
rect 5456 2387 5464 2593
rect 5476 2547 5484 2633
rect 5516 2567 5524 2753
rect 5556 2608 5564 2953
rect 5596 2944 5604 3033
rect 5576 2936 5604 2944
rect 5476 2467 5484 2533
rect 5516 2527 5524 2553
rect 5316 2307 5324 2373
rect 5376 2327 5384 2373
rect 5236 2187 5244 2233
rect 5256 2207 5264 2273
rect 5316 2147 5324 2253
rect 5336 2124 5344 2233
rect 5356 2127 5364 2253
rect 5316 2116 5344 2124
rect 5156 1647 5164 1712
rect 5096 1556 5124 1564
rect 5096 1284 5104 1556
rect 5116 1447 5124 1533
rect 5136 1507 5144 1613
rect 5176 1607 5184 1992
rect 5196 1787 5204 1853
rect 5236 1827 5244 2113
rect 5268 2084 5280 2087
rect 5268 2073 5284 2084
rect 5276 1887 5284 2073
rect 5296 2027 5304 2073
rect 5296 1827 5304 1933
rect 5296 1787 5304 1813
rect 5196 1776 5212 1787
rect 5200 1773 5212 1776
rect 5176 1593 5193 1607
rect 5176 1567 5184 1593
rect 5216 1504 5224 1713
rect 5276 1687 5284 1733
rect 5296 1647 5304 1773
rect 5316 1744 5324 2116
rect 5336 1907 5344 2033
rect 5356 2007 5364 2053
rect 5316 1736 5344 1744
rect 5276 1507 5284 1553
rect 5196 1496 5224 1504
rect 5076 1276 5104 1284
rect 5116 1284 5124 1393
rect 5156 1307 5164 1473
rect 5196 1464 5204 1496
rect 5316 1487 5324 1713
rect 5336 1627 5344 1736
rect 5356 1707 5364 1733
rect 5376 1684 5384 2133
rect 5396 1824 5404 2193
rect 5416 2187 5424 2293
rect 5436 1927 5444 2313
rect 5456 2247 5464 2333
rect 5496 2287 5504 2393
rect 5536 2307 5544 2453
rect 5556 2347 5564 2572
rect 5576 2347 5584 2936
rect 5560 2264 5573 2267
rect 5546 2253 5547 2260
rect 5476 2227 5484 2253
rect 5533 2244 5547 2253
rect 5496 2240 5547 2244
rect 5556 2253 5573 2264
rect 5496 2236 5544 2240
rect 5496 2204 5504 2236
rect 5556 2227 5564 2253
rect 5547 2216 5564 2227
rect 5547 2213 5560 2216
rect 5476 2196 5504 2204
rect 5476 2167 5484 2196
rect 5596 2127 5604 2913
rect 5616 2507 5624 3113
rect 5636 2927 5644 3413
rect 5656 2767 5664 3993
rect 5676 3704 5684 3953
rect 5696 3727 5704 5033
rect 5716 3767 5724 4993
rect 5676 3696 5704 3704
rect 5676 2727 5684 3673
rect 5636 2487 5644 2713
rect 5676 2607 5684 2673
rect 5696 2587 5704 3696
rect 5716 2827 5724 3553
rect 5716 2667 5724 2753
rect 5456 1964 5464 2113
rect 5456 1956 5484 1964
rect 5476 1904 5484 1956
rect 5476 1896 5504 1904
rect 5396 1816 5424 1824
rect 5416 1747 5424 1816
rect 5436 1708 5444 1773
rect 5356 1676 5384 1684
rect 5176 1456 5204 1464
rect 5176 1387 5184 1456
rect 5116 1276 5133 1284
rect 4996 987 5004 1033
rect 5076 1027 5084 1276
rect 5096 1167 5104 1253
rect 5136 1187 5144 1273
rect 5196 1267 5204 1293
rect 5236 1227 5244 1453
rect 5256 1167 5264 1353
rect 5116 1087 5124 1113
rect 5156 1107 5164 1153
rect 5147 1096 5164 1107
rect 5147 1093 5160 1096
rect 4916 836 4944 844
rect 4676 816 4693 827
rect 4680 813 4693 816
rect 4596 687 4604 773
rect 4516 607 4524 653
rect 4636 647 4644 793
rect 4676 627 4684 693
rect 4667 616 4684 627
rect 4667 613 4680 616
rect 4556 447 4564 513
rect 4596 407 4604 493
rect 4636 387 4644 433
rect 4326 376 4354 384
rect 4628 376 4644 387
rect 4628 373 4640 376
rect 4176 347 4184 373
rect 4436 267 4444 373
rect 4486 356 4533 364
rect 4556 287 4564 373
rect 4616 187 4624 293
rect 4656 247 4664 453
rect 4676 307 4684 473
rect 4716 467 4724 633
rect 4756 627 4764 713
rect 4796 707 4804 832
rect 4833 613 4834 620
rect 4833 607 4847 613
rect 4826 600 4847 607
rect 4826 596 4844 600
rect 4826 593 4840 596
rect 4856 587 4864 693
rect 4816 467 4824 533
rect 4716 404 4724 453
rect 4696 396 4724 404
rect 4753 407 4767 413
rect 4696 367 4704 396
rect 4816 367 4824 453
rect 4876 344 4884 713
rect 4847 336 4884 344
rect 4096 156 4113 167
rect 4100 153 4113 156
rect 4213 127 4227 133
rect 4176 67 4184 113
rect 4256 107 4264 153
rect 4396 127 4404 173
rect 4573 147 4587 153
rect 4616 147 4624 173
rect 4586 140 4587 147
rect 4387 116 4404 127
rect 4387 113 4400 116
rect 4273 93 4274 100
rect 4273 87 4287 93
rect 4316 67 4324 93
rect 4536 27 4544 133
rect 4776 127 4784 173
rect 4796 167 4804 253
rect 4836 147 4844 273
rect 4836 136 4853 147
rect 4840 133 4853 136
rect 4896 127 4904 753
rect 4916 527 4924 836
rect 4916 147 4924 393
rect 4936 187 4944 733
rect 4956 407 4964 613
rect 4976 447 4984 913
rect 4996 807 5004 833
rect 4996 627 5004 753
rect 4996 407 5004 493
rect 5016 327 5024 1013
rect 5036 707 5044 893
rect 5056 647 5064 913
rect 5046 636 5064 647
rect 5046 633 5060 636
rect 5036 427 5044 553
rect 5076 507 5084 633
rect 5096 427 5104 973
rect 5036 387 5044 413
rect 5036 376 5053 387
rect 5040 373 5053 376
rect 4956 167 4964 193
rect 5056 167 5064 313
rect 5096 267 5104 313
rect 5116 287 5124 993
rect 5136 687 5144 953
rect 5176 927 5184 1133
rect 5256 1107 5264 1153
rect 5200 1104 5213 1107
rect 5196 1093 5213 1104
rect 5196 1067 5204 1093
rect 5276 1087 5284 1413
rect 5316 1324 5324 1433
rect 5296 1316 5324 1324
rect 5296 1267 5304 1316
rect 5316 1207 5324 1293
rect 5336 1227 5344 1473
rect 5356 1204 5364 1676
rect 5396 1428 5404 1613
rect 5416 1447 5424 1693
rect 5436 1407 5444 1672
rect 5456 1467 5464 1733
rect 5476 1667 5484 1873
rect 5496 1624 5504 1896
rect 5516 1887 5524 2113
rect 5553 2087 5567 2093
rect 5536 1867 5544 2033
rect 5556 1887 5564 1973
rect 5576 1904 5584 2053
rect 5616 2027 5624 2173
rect 5636 2047 5644 2413
rect 5656 2027 5664 2553
rect 5676 2387 5684 2513
rect 5676 2067 5684 2333
rect 5696 2007 5704 2493
rect 5716 2407 5724 2453
rect 5716 2107 5724 2353
rect 5636 1967 5644 1993
rect 5576 1896 5604 1904
rect 5536 1787 5544 1853
rect 5596 1827 5604 1896
rect 5476 1616 5504 1624
rect 5476 1424 5484 1616
rect 5516 1607 5524 1693
rect 5507 1596 5524 1607
rect 5507 1593 5520 1596
rect 5496 1567 5504 1593
rect 5536 1587 5544 1733
rect 5556 1687 5564 1713
rect 5576 1587 5584 1793
rect 5596 1780 5604 1784
rect 5593 1767 5607 1780
rect 5596 1667 5604 1753
rect 5616 1647 5624 1913
rect 5636 1707 5644 1753
rect 5520 1586 5544 1587
rect 5527 1575 5544 1586
rect 5527 1573 5540 1575
rect 5568 1576 5584 1587
rect 5568 1573 5580 1576
rect 5496 1527 5504 1553
rect 5507 1516 5524 1524
rect 5476 1416 5504 1424
rect 5336 1196 5364 1204
rect 5316 1067 5324 1133
rect 5196 907 5204 1053
rect 5236 887 5244 913
rect 5176 847 5184 873
rect 5156 787 5164 813
rect 5276 727 5284 893
rect 5296 867 5304 933
rect 5336 907 5344 1196
rect 5376 1127 5384 1293
rect 5396 947 5404 1392
rect 5496 1387 5504 1416
rect 5516 1407 5524 1516
rect 5416 1307 5424 1333
rect 5456 1327 5464 1353
rect 5353 867 5367 873
rect 5396 827 5404 893
rect 5196 627 5204 653
rect 5276 648 5284 713
rect 5187 616 5204 627
rect 5280 626 5300 627
rect 5187 613 5200 616
rect 5136 324 5144 613
rect 5287 623 5300 626
rect 5287 613 5304 623
rect 5233 593 5234 600
rect 5233 587 5247 593
rect 5233 580 5234 587
rect 5216 507 5224 573
rect 5296 547 5304 613
rect 5156 407 5164 493
rect 5236 387 5244 473
rect 5316 407 5324 693
rect 5316 367 5324 393
rect 5166 356 5194 364
rect 5308 356 5324 367
rect 5308 353 5320 356
rect 5136 316 5244 324
rect 5176 147 5184 253
rect 4916 136 4933 147
rect 4920 133 4933 136
rect 4887 116 4904 127
rect 4887 113 4900 116
rect 4987 96 5084 104
rect 5076 24 5084 96
rect 5116 47 5124 133
rect 5236 87 5244 316
rect 5276 187 5284 233
rect 5316 167 5324 193
rect 5336 147 5344 713
rect 5356 647 5364 793
rect 5396 707 5404 813
rect 5416 747 5424 1133
rect 5476 1127 5484 1253
rect 5436 907 5444 1053
rect 5456 947 5464 1033
rect 5496 987 5504 1373
rect 5516 1107 5524 1213
rect 5536 1147 5544 1513
rect 5556 1367 5564 1433
rect 5556 1167 5564 1353
rect 5576 1187 5584 1493
rect 5596 1207 5604 1553
rect 5616 1547 5624 1593
rect 5636 1487 5644 1613
rect 5656 1527 5664 1973
rect 5676 1687 5684 1753
rect 5696 1748 5704 1953
rect 5716 1807 5724 1853
rect 5456 936 5473 947
rect 5460 933 5473 936
rect 5536 887 5544 973
rect 5556 947 5564 1013
rect 5436 827 5444 853
rect 5476 847 5484 873
rect 5487 844 5500 847
rect 5487 833 5504 844
rect 5436 667 5444 813
rect 5496 807 5504 833
rect 5536 827 5544 873
rect 5436 656 5452 667
rect 5440 653 5452 656
rect 5356 636 5373 647
rect 5360 633 5373 636
rect 5356 187 5364 513
rect 5376 227 5384 553
rect 5396 387 5404 653
rect 5476 467 5484 653
rect 5536 507 5544 593
rect 5396 247 5404 313
rect 5416 207 5424 433
rect 5536 387 5544 493
rect 5433 364 5447 373
rect 5433 360 5464 364
rect 5436 356 5464 360
rect 5293 107 5307 113
rect 5153 24 5167 33
rect 5436 27 5444 313
rect 5456 307 5464 356
rect 5456 127 5464 233
rect 5556 227 5564 673
rect 5576 204 5584 1133
rect 5616 1127 5624 1413
rect 5596 1008 5604 1073
rect 5596 867 5604 972
rect 5636 964 5644 1233
rect 5656 1187 5664 1273
rect 5676 1247 5684 1633
rect 5696 1567 5704 1712
rect 5716 1627 5724 1673
rect 5696 1224 5704 1473
rect 5676 1216 5704 1224
rect 5636 956 5664 964
rect 5636 827 5644 933
rect 5596 308 5604 373
rect 5596 207 5604 272
rect 5556 196 5584 204
rect 5516 87 5524 153
rect 5556 147 5564 196
rect 5616 107 5624 753
rect 5656 727 5664 956
rect 5676 864 5684 1216
rect 5696 927 5704 1193
rect 5676 856 5704 864
rect 5676 567 5684 833
rect 5636 367 5644 413
rect 5676 327 5684 393
rect 5696 47 5704 856
rect 5716 267 5724 1393
rect 5076 20 5167 24
rect 5076 16 5164 20
use INVX1  _927_
timestamp 0
transform -1 0 4350 0 -1 5050
box -6 -8 66 248
use NOR2X1  _928_
timestamp 0
transform 1 0 3830 0 -1 4090
box -6 -8 86 248
use NAND2X1  _929_
timestamp 0
transform -1 0 3950 0 1 4090
box -6 -8 86 248
use INVX1  _930_
timestamp 0
transform 1 0 3990 0 1 4090
box -6 -8 66 248
use INVX1  _931_
timestamp 0
transform 1 0 4190 0 -1 5050
box -6 -8 66 248
use INVX2  _932_
timestamp 0
transform -1 0 2930 0 1 1210
box -6 -8 66 248
use NOR2X1  _933_
timestamp 0
transform 1 0 4390 0 -1 5050
box -6 -8 86 248
use NAND2X1  _934_
timestamp 0
transform -1 0 4710 0 -1 5050
box -6 -8 86 248
use INVX1  _935_
timestamp 0
transform 1 0 5570 0 1 3610
box -6 -8 66 248
use NOR2X1  _936_
timestamp 0
transform 1 0 4510 0 -1 5050
box -6 -8 86 248
use AOI21X1  _937_
timestamp 0
transform 1 0 4830 0 1 5050
box -6 -8 106 248
use NOR2X1  _938_
timestamp 0
transform -1 0 5070 0 1 5530
box -6 -8 86 248
use OAI21X1  _939_
timestamp 0
transform -1 0 4950 0 1 5530
box -6 -8 106 248
use INVX1  _940_
timestamp 0
transform -1 0 4150 0 -1 5530
box -6 -8 66 248
use INVX4  _941_
timestamp 0
transform -1 0 3710 0 -1 3130
box -6 -8 86 248
use OAI21X1  _942_
timestamp 0
transform -1 0 4150 0 -1 5050
box -6 -8 106 248
use INVX1  _943_
timestamp 0
transform -1 0 4390 0 -1 5530
box -6 -8 66 248
use NOR2X1  _944_
timestamp 0
transform -1 0 3750 0 1 2650
box -6 -8 86 248
use INVX1  _945_
timestamp 0
transform -1 0 4050 0 -1 5530
box -6 -8 66 248
use INVX1  _946_
timestamp 0
transform 1 0 5110 0 1 5530
box -6 -8 66 248
use OAI21X1  _947_
timestamp 0
transform 1 0 4970 0 1 5050
box -6 -8 106 248
use OAI21X1  _948_
timestamp 0
transform 1 0 4690 0 1 5050
box -6 -8 106 248
use AOI22X1  _949_
timestamp 0
transform 1 0 4530 0 1 5050
box -6 -8 126 248
use NAND2X1  _950_
timestamp 0
transform -1 0 4330 0 1 5530
box -6 -8 86 248
use OAI21X1  _951_
timestamp 0
transform 1 0 4430 0 -1 5530
box -6 -8 106 248
use OAI21X1  _952_
timestamp 0
transform 1 0 4570 0 -1 5530
box -6 -8 106 248
use NAND2X1  _953_
timestamp 0
transform 1 0 4510 0 1 4570
box -6 -8 86 248
use NOR2X1  _954_
timestamp 0
transform 1 0 4990 0 -1 5530
box -6 -8 86 248
use NOR2X1  _955_
timestamp 0
transform 1 0 5110 0 -1 5530
box -6 -8 86 248
use OAI22X1  _956_
timestamp 0
transform 1 0 5370 0 -1 5530
box -6 -8 126 248
use OR2X2  _957_
timestamp 0
transform 1 0 5230 0 -1 5530
box -6 -8 106 248
use INVX1  _958_
timestamp 0
transform 1 0 5590 0 1 5050
box -6 -8 66 248
use AOI22X1  _959_
timestamp 0
transform -1 0 5650 0 -1 5530
box -6 -8 126 248
use NAND3X1  _960_
timestamp 0
transform 1 0 4190 0 -1 5530
box -6 -8 106 248
use AND2X2  _961_
timestamp 0
transform -1 0 4950 0 -1 5530
box -6 -8 106 248
use OAI21X1  _962_
timestamp 0
transform 1 0 4710 0 -1 5530
box -6 -8 106 248
use INVX1  _963_
timestamp 0
transform -1 0 5270 0 1 5530
box -6 -8 66 248
use INVX1  _964_
timestamp 0
transform 1 0 4350 0 1 3130
box -6 -8 66 248
use NAND2X1  _965_
timestamp 0
transform 1 0 4470 0 -1 3610
box -6 -8 86 248
use OAI21X1  _966_
timestamp 0
transform 1 0 4330 0 -1 3610
box -6 -8 106 248
use INVX1  _967_
timestamp 0
transform -1 0 4510 0 1 3130
box -6 -8 66 248
use NAND2X1  _968_
timestamp 0
transform -1 0 4170 0 1 3130
box -6 -8 86 248
use OAI21X1  _969_
timestamp 0
transform -1 0 4310 0 1 3130
box -6 -8 106 248
use INVX1  _970_
timestamp 0
transform 1 0 5230 0 1 3610
box -6 -8 66 248
use NAND2X1  _971_
timestamp 0
transform -1 0 4410 0 -1 4090
box -6 -8 86 248
use OAI21X1  _972_
timestamp 0
transform -1 0 4550 0 -1 4090
box -6 -8 106 248
use INVX1  _973_
timestamp 0
transform -1 0 5430 0 -1 4090
box -6 -8 66 248
use NAND2X1  _974_
timestamp 0
transform 1 0 4210 0 1 4090
box -6 -8 86 248
use OAI21X1  _975_
timestamp 0
transform -1 0 4430 0 1 4090
box -6 -8 106 248
use INVX1  _976_
timestamp 0
transform -1 0 5410 0 1 4570
box -6 -8 66 248
use NAND2X1  _977_
timestamp 0
transform -1 0 5530 0 1 4090
box -6 -8 86 248
use OAI21X1  _978_
timestamp 0
transform 1 0 5510 0 -1 4570
box -6 -8 106 248
use INVX1  _979_
timestamp 0
transform -1 0 5310 0 -1 5050
box -6 -8 66 248
use NAND2X1  _980_
timestamp 0
transform 1 0 4990 0 -1 5050
box -6 -8 86 248
use OAI21X1  _981_
timestamp 0
transform -1 0 5210 0 -1 5050
box -6 -8 106 248
use INVX1  _982_
timestamp 0
transform 1 0 4630 0 1 4570
box -6 -8 66 248
use NAND2X1  _983_
timestamp 0
transform -1 0 4230 0 -1 4570
box -6 -8 86 248
use OAI21X1  _984_
timestamp 0
transform -1 0 4370 0 -1 4570
box -6 -8 106 248
use INVX4  _985_
timestamp 0
transform -1 0 3290 0 1 730
box -6 -8 86 248
use NAND2X1  _986_
timestamp 0
transform 1 0 5330 0 1 4090
box -6 -8 86 248
use OAI21X1  _987_
timestamp 0
transform 1 0 5190 0 1 4090
box -6 -8 106 248
use INVX1  _988_
timestamp 0
transform -1 0 3130 0 1 2650
box -6 -8 66 248
use INVX1  _989_
timestamp 0
transform -1 0 2770 0 1 1690
box -6 -8 66 248
use INVX2  _990_
timestamp 0
transform 1 0 2490 0 1 2170
box -6 -8 66 248
use NOR2X1  _991_
timestamp 0
transform 1 0 2470 0 1 1690
box -6 -8 86 248
use AND2X2  _992_
timestamp 0
transform 1 0 2610 0 -1 2170
box -6 -8 106 248
use NAND2X1  _993_
timestamp 0
transform 1 0 2150 0 1 250
box -6 -8 86 248
use NAND2X1  _994_
timestamp 0
transform -1 0 2430 0 1 1210
box -6 -8 86 248
use NAND2X1  _995_
timestamp 0
transform -1 0 1610 0 1 1210
box -6 -8 86 248
use OR2X2  _996_
timestamp 0
transform 1 0 1870 0 1 730
box -6 -8 106 248
use NAND2X1  _997_
timestamp 0
transform -1 0 2890 0 1 1690
box -6 -8 86 248
use AND2X2  _998_
timestamp 0
transform 1 0 2290 0 1 730
box -6 -8 106 248
use OAI21X1  _999_
timestamp 0
transform -1 0 2690 0 -1 730
box -6 -8 106 248
use NAND2X1  _1000_
timestamp 0
transform 1 0 1410 0 1 1210
box -6 -8 86 248
use INVX1  _1001_
timestamp 0
transform -1 0 1450 0 1 730
box -6 -8 66 248
use NAND2X1  _1002_
timestamp 0
transform 1 0 2970 0 -1 2170
box -6 -8 86 248
use OR2X2  _1003_
timestamp 0
transform -1 0 1590 0 1 730
box -6 -8 106 248
use AOI22X1  _1004_
timestamp 0
transform -1 0 1890 0 -1 2170
box -6 -8 126 248
use INVX1  _1005_
timestamp 0
transform 1 0 1830 0 -1 730
box -6 -8 66 248
use NAND3X1  _1006_
timestamp 0
transform -1 0 1510 0 -1 730
box -6 -8 106 248
use NOR2X1  _1007_
timestamp 0
transform 1 0 1630 0 1 730
box -6 -8 86 248
use OAI21X1  _1008_
timestamp 0
transform -1 0 1370 0 -1 730
box -6 -8 106 248
use NAND3X1  _1009_
timestamp 0
transform -1 0 1010 0 1 250
box -6 -8 106 248
use INVX1  _1010_
timestamp 0
transform 1 0 2490 0 -1 730
box -6 -8 66 248
use NAND2X1  _1011_
timestamp 0
transform 1 0 2590 0 1 2170
box -6 -8 86 248
use INVX2  _1012_
timestamp 0
transform 1 0 2010 0 -1 4090
box -6 -8 66 248
use NAND2X1  _1013_
timestamp 0
transform 1 0 2590 0 1 1690
box -6 -8 86 248
use OAI21X1  _1014_
timestamp 0
transform 1 0 2330 0 1 1690
box -6 -8 106 248
use OAI21X1  _1015_
timestamp 0
transform -1 0 2450 0 -1 730
box -6 -8 106 248
use AOI21X1  _1016_
timestamp 0
transform 1 0 1050 0 1 250
box -6 -8 106 248
use OAI21X1  _1017_
timestamp 0
transform -1 0 870 0 1 250
box -6 -8 106 248
use OAI21X1  _1018_
timestamp 0
transform -1 0 1350 0 1 730
box -6 -8 106 248
use AND2X2  _1019_
timestamp 0
transform -1 0 1450 0 1 2650
box -6 -8 106 248
use NAND3X1  _1020_
timestamp 0
transform -1 0 1090 0 -1 2650
box -6 -8 106 248
use AOI22X1  _1021_
timestamp 0
transform -1 0 1610 0 -1 2170
box -6 -8 126 248
use INVX1  _1022_
timestamp 0
transform -1 0 110 0 1 730
box -6 -8 66 248
use NAND2X1  _1023_
timestamp 0
transform -1 0 1370 0 1 1210
box -6 -8 86 248
use INVX1  _1024_
timestamp 0
transform -1 0 110 0 -1 730
box -6 -8 66 248
use NAND3X1  _1025_
timestamp 0
transform 1 0 430 0 1 730
box -6 -8 106 248
use NAND2X1  _1026_
timestamp 0
transform -1 0 1730 0 -1 2170
box -6 -8 86 248
use NOR2X1  _1027_
timestamp 0
transform -1 0 1210 0 1 730
box -6 -8 86 248
use OAI21X1  _1028_
timestamp 0
transform -1 0 670 0 1 730
box -6 -8 106 248
use NAND3X1  _1029_
timestamp 0
transform 1 0 710 0 1 730
box -6 -8 106 248
use AOI21X1  _1030_
timestamp 0
transform -1 0 1650 0 -1 730
box -6 -8 106 248
use OAI21X1  _1031_
timestamp 0
transform -1 0 250 0 -1 730
box -6 -8 106 248
use NAND3X1  _1032_
timestamp 0
transform 1 0 290 0 1 730
box -6 -8 106 248
use NAND3X1  _1033_
timestamp 0
transform -1 0 390 0 -1 730
box -6 -8 106 248
use NAND2X1  _1034_
timestamp 0
transform 1 0 2850 0 -1 2170
box -6 -8 86 248
use INVX1  _1035_
timestamp 0
transform 1 0 2750 0 -1 2170
box -6 -8 66 248
use AND2X2  _1036_
timestamp 0
transform -1 0 2330 0 1 2170
box -6 -8 106 248
use NAND2X1  _1037_
timestamp 0
transform -1 0 2290 0 -1 2170
box -6 -8 86 248
use INVX1  _1038_
timestamp 0
transform 1 0 2530 0 1 3610
box -6 -8 66 248
use OAI21X1  _1039_
timestamp 0
transform 1 0 2470 0 -1 2170
box -6 -8 106 248
use NAND3X1  _1040_
timestamp 0
transform -1 0 2430 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1041_
timestamp 0
transform 1 0 2070 0 -1 2170
box -6 -8 106 248
use INVX1  _1042_
timestamp 0
transform -1 0 1530 0 -1 2650
box -6 -8 66 248
use OAI21X1  _1043_
timestamp 0
transform -1 0 1930 0 1 2170
box -6 -8 106 248
use NAND3X1  _1044_
timestamp 0
transform -1 0 2030 0 -1 2170
box -6 -8 106 248
use AND2X2  _1045_
timestamp 0
transform -1 0 1650 0 1 1690
box -6 -8 106 248
use NAND3X1  _1046_
timestamp 0
transform -1 0 810 0 -1 730
box -6 -8 106 248
use AOI21X1  _1047_
timestamp 0
transform 1 0 430 0 -1 730
box -6 -8 106 248
use AOI21X1  _1048_
timestamp 0
transform 1 0 850 0 1 730
box -6 -8 106 248
use NAND2X1  _1049_
timestamp 0
transform 1 0 1690 0 1 1690
box -6 -8 86 248
use OAI21X1  _1050_
timestamp 0
transform 1 0 1130 0 -1 730
box -6 -8 106 248
use NAND3X1  _1051_
timestamp 0
transform -1 0 150 0 1 250
box -6 -8 106 248
use AOI21X1  _1052_
timestamp 0
transform 1 0 190 0 1 250
box -6 -8 106 248
use OAI21X1  _1053_
timestamp 0
transform 1 0 330 0 1 250
box -6 -8 106 248
use AOI21X1  _1054_
timestamp 0
transform -1 0 670 0 -1 730
box -6 -8 106 248
use OAI21X1  _1055_
timestamp 0
transform 1 0 890 0 -1 1690
box -6 -8 106 248
use AND2X2  _1056_
timestamp 0
transform -1 0 1650 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1057_
timestamp 0
transform 1 0 1110 0 1 2650
box -6 -8 86 248
use INVX1  _1058_
timestamp 0
transform -1 0 1470 0 1 3130
box -6 -8 66 248
use INVX2  _1059_
timestamp 0
transform -1 0 2530 0 1 4570
box -6 -8 66 248
use NAND2X1  _1060_
timestamp 0
transform 1 0 1350 0 -1 3130
box -6 -8 86 248
use OAI21X1  _1061_
timestamp 0
transform -1 0 1370 0 1 3130
box -6 -8 106 248
use NAND2X1  _1062_
timestamp 0
transform -1 0 1070 0 1 2650
box -6 -8 86 248
use INVX1  _1063_
timestamp 0
transform -1 0 830 0 -1 2650
box -6 -8 66 248
use NAND3X1  _1064_
timestamp 0
transform 1 0 750 0 1 2170
box -6 -8 106 248
use NAND2X1  _1065_
timestamp 0
transform -1 0 1510 0 -1 3610
box -6 -8 86 248
use NOR2X1  _1066_
timestamp 0
transform 1 0 1130 0 -1 2650
box -6 -8 86 248
use AOI22X1  _1067_
timestamp 0
transform 1 0 1490 0 1 2650
box -6 -8 126 248
use OAI21X1  _1068_
timestamp 0
transform 1 0 890 0 1 2170
box -6 -8 106 248
use AOI21X1  _1069_
timestamp 0
transform -1 0 850 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1070_
timestamp 0
transform 1 0 150 0 1 730
box -6 -8 106 248
use OAI21X1  _1071_
timestamp 0
transform -1 0 710 0 1 2170
box -6 -8 106 248
use NAND3X1  _1072_
timestamp 0
transform -1 0 570 0 1 2170
box -6 -8 106 248
use AOI21X1  _1073_
timestamp 0
transform -1 0 430 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1074_
timestamp 0
transform -1 0 1970 0 1 2650
box -6 -8 86 248
use INVX1  _1075_
timestamp 0
transform -1 0 1930 0 -1 2650
box -6 -8 66 248
use AND2X2  _1076_
timestamp 0
transform -1 0 2350 0 -1 2650
box -6 -8 106 248
use AND2X2  _1077_
timestamp 0
transform -1 0 2370 0 1 2650
box -6 -8 106 248
use NAND2X1  _1078_
timestamp 0
transform 1 0 2150 0 1 2650
box -6 -8 86 248
use INVX2  _1079_
timestamp 0
transform 1 0 1710 0 -1 4570
box -6 -8 66 248
use NAND2X1  _1080_
timestamp 0
transform -1 0 2190 0 1 2170
box -6 -8 86 248
use OAI21X1  _1081_
timestamp 0
transform 1 0 1970 0 1 2170
box -6 -8 106 248
use NAND3X1  _1082_
timestamp 0
transform -1 0 1670 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1083_
timestamp 0
transform 1 0 2110 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1084_
timestamp 0
transform -1 0 2110 0 1 2650
box -6 -8 106 248
use NAND3X1  _1085_
timestamp 0
transform -1 0 2070 0 -1 2650
box -6 -8 106 248
use AND2X2  _1086_
timestamp 0
transform -1 0 710 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1087_
timestamp 0
transform -1 0 150 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1088_
timestamp 0
transform 1 0 470 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1089_
timestamp 0
transform -1 0 710 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1090_
timestamp 0
transform 1 0 750 0 -1 2170
box -6 -8 86 248
use NAND3X1  _1091_
timestamp 0
transform 1 0 190 0 1 1210
box -6 -8 106 248
use NAND3X1  _1092_
timestamp 0
transform -1 0 290 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1093_
timestamp 0
transform -1 0 1090 0 1 730
box -6 -8 106 248
use NAND3X1  _1094_
timestamp 0
transform 1 0 330 0 1 1210
box -6 -8 106 248
use OAI21X1  _1095_
timestamp 0
transform -1 0 150 0 1 1210
box -6 -8 106 248
use NAND3X1  _1096_
timestamp 0
transform 1 0 610 0 -1 1210
box -6 -8 106 248
use INVX4  _1097_
timestamp 0
transform -1 0 3770 0 -1 5050
box -6 -8 86 248
use NOR2X1  _1098_
timestamp 0
transform -1 0 2290 0 1 1690
box -6 -8 86 248
use OAI21X1  _1099_
timestamp 0
transform -1 0 2170 0 1 1690
box -6 -8 106 248
use NAND2X1  _1100_
timestamp 0
transform 1 0 1950 0 1 1690
box -6 -8 86 248
use OR2X2  _1101_
timestamp 0
transform -1 0 1910 0 1 1690
box -6 -8 106 248
use AND2X2  _1102_
timestamp 0
transform -1 0 1130 0 1 1210
box -6 -8 106 248
use NAND3X1  _1103_
timestamp 0
transform 1 0 890 0 1 1210
box -6 -8 106 248
use AOI21X1  _1104_
timestamp 0
transform 1 0 470 0 -1 1210
box -6 -8 106 248
use AOI21X1  _1105_
timestamp 0
transform 1 0 330 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1106_
timestamp 0
transform 1 0 1170 0 1 1210
box -6 -8 86 248
use OAI21X1  _1107_
timestamp 0
transform 1 0 750 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1108_
timestamp 0
transform 1 0 1190 0 -1 1210
box -6 -8 106 248
use INVX1  _1109_
timestamp 0
transform -1 0 1510 0 1 1690
box -6 -8 66 248
use OAI21X1  _1110_
timestamp 0
transform -1 0 850 0 1 1210
box -6 -8 106 248
use AOI21X1  _1111_
timestamp 0
transform -1 0 290 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1112_
timestamp 0
transform -1 0 570 0 1 2650
box -6 -8 106 248
use NAND3X1  _1113_
timestamp 0
transform -1 0 1310 0 -1 3130
box -6 -8 106 248
use AOI22X1  _1114_
timestamp 0
transform 1 0 1470 0 -1 3130
box -6 -8 126 248
use INVX1  _1115_
timestamp 0
transform 1 0 730 0 -1 3130
box -6 -8 66 248
use NAND2X1  _1116_
timestamp 0
transform 1 0 1230 0 1 2650
box -6 -8 86 248
use INVX1  _1117_
timestamp 0
transform -1 0 670 0 1 2650
box -6 -8 66 248
use NAND3X1  _1118_
timestamp 0
transform -1 0 410 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1119_
timestamp 0
transform 1 0 1090 0 -1 3130
box -6 -8 86 248
use NOR2X1  _1120_
timestamp 0
transform -1 0 1050 0 -1 3130
box -6 -8 86 248
use OAI21X1  _1121_
timestamp 0
transform 1 0 850 0 1 2650
box -6 -8 106 248
use AOI21X1  _1122_
timestamp 0
transform -1 0 430 0 1 2650
box -6 -8 106 248
use OAI21X1  _1123_
timestamp 0
transform -1 0 810 0 1 2650
box -6 -8 106 248
use NAND3X1  _1124_
timestamp 0
transform -1 0 690 0 -1 3130
box -6 -8 106 248
use AOI22X1  _1125_
timestamp 0
transform -1 0 590 0 -1 2650
box -6 -8 126 248
use NAND2X1  _1126_
timestamp 0
transform 1 0 2330 0 -1 3610
box -6 -8 86 248
use INVX1  _1127_
timestamp 0
transform -1 0 1830 0 1 3130
box -6 -8 66 248
use AND2X2  _1128_
timestamp 0
transform 1 0 1870 0 1 3130
box -6 -8 106 248
use AND2X2  _1129_
timestamp 0
transform 1 0 2170 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1130_
timestamp 0
transform 1 0 2010 0 1 3130
box -6 -8 86 248
use AOI22X1  _1131_
timestamp 0
transform -1 0 2230 0 -1 4090
box -6 -8 126 248
use INVX1  _1132_
timestamp 0
transform 1 0 2230 0 -1 3610
box -6 -8 66 248
use NAND3X1  _1133_
timestamp 0
transform -1 0 1730 0 1 3130
box -6 -8 106 248
use INVX1  _1134_
timestamp 0
transform 1 0 2890 0 1 4090
box -6 -8 66 248
use OAI21X1  _1135_
timestamp 0
transform 1 0 1890 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1136_
timestamp 0
transform -1 0 2130 0 -1 3130
box -6 -8 106 248
use NAND3X1  _1137_
timestamp 0
transform -1 0 1850 0 -1 3130
box -6 -8 106 248
use AND2X2  _1138_
timestamp 0
transform -1 0 150 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1139_
timestamp 0
transform -1 0 290 0 1 2170
box -6 -8 106 248
use AOI21X1  _1140_
timestamp 0
transform -1 0 730 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1141_
timestamp 0
transform -1 0 430 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1142_
timestamp 0
transform -1 0 290 0 1 2650
box -6 -8 106 248
use NAND2X1  _1143_
timestamp 0
transform 1 0 190 0 -1 3130
box -6 -8 86 248
use NAND3X1  _1144_
timestamp 0
transform -1 0 150 0 1 2170
box -6 -8 106 248
use NAND3X1  _1145_
timestamp 0
transform 1 0 190 0 1 1690
box -6 -8 106 248
use OAI21X1  _1146_
timestamp 0
transform -1 0 150 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1147_
timestamp 0
transform -1 0 150 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1148_
timestamp 0
transform 1 0 330 0 1 2170
box -6 -8 106 248
use NAND3X1  _1149_
timestamp 0
transform 1 0 190 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1150_
timestamp 0
transform -1 0 2450 0 1 2170
box -6 -8 86 248
use INVX1  _1151_
timestamp 0
transform -1 0 1450 0 -1 2170
box -6 -8 66 248
use AOI22X1  _1152_
timestamp 0
transform -1 0 1830 0 -1 2650
box -6 -8 126 248
use INVX1  _1153_
timestamp 0
transform -1 0 1430 0 -1 2650
box -6 -8 66 248
use OAI21X1  _1154_
timestamp 0
transform -1 0 1530 0 1 2170
box -6 -8 106 248
use NOR2X1  _1155_
timestamp 0
transform 1 0 1570 0 1 2170
box -6 -8 86 248
use NAND2X1  _1156_
timestamp 0
transform 1 0 1310 0 1 2170
box -6 -8 86 248
use NAND3X1  _1157_
timestamp 0
transform -1 0 1210 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1158_
timestamp 0
transform -1 0 1330 0 -1 2650
box -6 -8 86 248
use OAI21X1  _1159_
timestamp 0
transform -1 0 1790 0 1 2170
box -6 -8 106 248
use NAND3X1  _1160_
timestamp 0
transform -1 0 1270 0 1 2170
box -6 -8 106 248
use NAND2X1  _1161_
timestamp 0
transform -1 0 1070 0 -1 2170
box -6 -8 86 248
use NAND3X1  _1162_
timestamp 0
transform 1 0 750 0 1 1690
box -6 -8 106 248
use AOI21X1  _1163_
timestamp 0
transform -1 0 150 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1164_
timestamp 0
transform -1 0 150 0 1 1690
box -6 -8 106 248
use NAND3X1  _1165_
timestamp 0
transform -1 0 1130 0 1 2170
box -6 -8 106 248
use NAND3X1  _1166_
timestamp 0
transform -1 0 1350 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1167_
timestamp 0
transform 1 0 870 0 -1 2170
box -6 -8 86 248
use OAI21X1  _1168_
timestamp 0
transform 1 0 470 0 1 1690
box -6 -8 106 248
use AOI21X1  _1169_
timestamp 0
transform 1 0 1030 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1170_
timestamp 0
transform -1 0 570 0 1 1210
box -6 -8 106 248
use OAI21X1  _1171_
timestamp 0
transform 1 0 330 0 1 1690
box -6 -8 106 248
use NAND3X1  _1172_
timestamp 0
transform 1 0 610 0 1 1690
box -6 -8 106 248
use AOI21X1  _1173_
timestamp 0
transform 1 0 1030 0 1 1690
box -6 -8 106 248
use OAI21X1  _1174_
timestamp 0
transform 1 0 1450 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1175_
timestamp 0
transform 1 0 890 0 1 1690
box -6 -8 106 248
use NAND3X1  _1176_
timestamp 0
transform 1 0 1170 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1177_
timestamp 0
transform 1 0 1870 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1178_
timestamp 0
transform 1 0 2010 0 -1 1690
box -6 -8 106 248
use INVX1  _1179_
timestamp 0
transform -1 0 2630 0 -1 1690
box -6 -8 66 248
use INVX1  _1180_
timestamp 0
transform -1 0 110 0 -1 250
box -6 -8 66 248
use NOR2X1  _1181_
timestamp 0
transform -1 0 1830 0 1 730
box -6 -8 86 248
use INVX1  _1182_
timestamp 0
transform -1 0 2490 0 1 730
box -6 -8 66 248
use INVX1  _1183_
timestamp 0
transform 1 0 1870 0 1 1210
box -6 -8 66 248
use OAI21X1  _1184_
timestamp 0
transform 1 0 1970 0 1 1210
box -6 -8 106 248
use AOI21X1  _1185_
timestamp 0
transform -1 0 2110 0 1 730
box -6 -8 106 248
use OAI21X1  _1186_
timestamp 0
transform -1 0 1790 0 -1 730
box -6 -8 106 248
use NAND3X1  _1187_
timestamp 0
transform 1 0 1930 0 -1 730
box -6 -8 106 248
use AOI21X1  _1188_
timestamp 0
transform 1 0 2210 0 -1 730
box -6 -8 106 248
use AND2X2  _1189_
timestamp 0
transform -1 0 1710 0 1 250
box -6 -8 106 248
use NAND3X1  _1190_
timestamp 0
transform -1 0 2170 0 -1 730
box -6 -8 106 248
use AOI21X1  _1191_
timestamp 0
transform -1 0 1570 0 1 250
box -6 -8 106 248
use OAI21X1  _1192_
timestamp 0
transform -1 0 1090 0 -1 730
box -6 -8 106 248
use NAND3X1  _1193_
timestamp 0
transform -1 0 950 0 -1 730
box -6 -8 106 248
use NAND3X1  _1194_
timestamp 0
transform -1 0 570 0 1 250
box -6 -8 106 248
use NAND3X1  _1195_
timestamp 0
transform 1 0 150 0 -1 250
box -6 -8 106 248
use OAI21X1  _1196_
timestamp 0
transform -1 0 710 0 1 1210
box -6 -8 106 248
use NAND3X1  _1197_
timestamp 0
transform 1 0 890 0 -1 1210
box -6 -8 106 248
use AOI22X1  _1198_
timestamp 0
transform -1 0 1150 0 -1 1210
box -6 -8 126 248
use NAND3X1  _1199_
timestamp 0
transform 1 0 1590 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1200_
timestamp 0
transform 1 0 1310 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1201_
timestamp 0
transform 1 0 1730 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1202_
timestamp 0
transform -1 0 1430 0 1 250
box -6 -8 106 248
use NAND3X1  _1203_
timestamp 0
transform 1 0 2150 0 1 730
box -6 -8 106 248
use NAND2X1  _1204_
timestamp 0
transform 1 0 3230 0 1 1690
box -6 -8 86 248
use NAND2X1  _1205_
timestamp 0
transform -1 0 2550 0 1 1210
box -6 -8 86 248
use AOI22X1  _1206_
timestamp 0
transform -1 0 3190 0 1 1690
box -6 -8 126 248
use OAI22X1  _1207_
timestamp 0
transform 1 0 2710 0 1 1210
box -6 -8 126 248
use OAI21X1  _1208_
timestamp 0
transform 1 0 2730 0 -1 730
box -6 -8 106 248
use NAND3X1  _1209_
timestamp 0
transform -1 0 2970 0 -1 730
box -6 -8 106 248
use AOI21X1  _1210_
timestamp 0
transform 1 0 3010 0 -1 730
box -6 -8 106 248
use OAI21X1  _1211_
timestamp 0
transform -1 0 1930 0 -1 250
box -6 -8 106 248
use OAI21X1  _1212_
timestamp 0
transform -1 0 1290 0 1 250
box -6 -8 106 248
use NAND3X1  _1213_
timestamp 0
transform -1 0 1190 0 -1 250
box -6 -8 106 248
use INVX1  _1214_
timestamp 0
transform 1 0 990 0 -1 250
box -6 -8 66 248
use AOI22X1  _1215_
timestamp 0
transform -1 0 730 0 1 250
box -6 -8 126 248
use OAI21X1  _1216_
timestamp 0
transform 1 0 430 0 -1 250
box -6 -8 106 248
use NAND3X1  _1217_
timestamp 0
transform 1 0 850 0 -1 250
box -6 -8 106 248
use AOI21X1  _1218_
timestamp 0
transform 1 0 1330 0 -1 1210
box -6 -8 106 248
use NOR3X1  _1219_
timestamp 0
transform 1 0 1650 0 1 1210
box -6 -8 186 248
use INVX1  _1220_
timestamp 0
transform -1 0 2330 0 1 250
box -6 -8 66 248
use NAND3X1  _1221_
timestamp 0
transform 1 0 2370 0 1 250
box -6 -8 106 248
use INVX1  _1222_
timestamp 0
transform 1 0 2910 0 -1 1210
box -6 -8 66 248
use NOR2X1  _1223_
timestamp 0
transform -1 0 2670 0 1 1210
box -6 -8 86 248
use NOR2X1  _1224_
timestamp 0
transform 1 0 2790 0 -1 1210
box -6 -8 86 248
use NAND2X1  _1225_
timestamp 0
transform -1 0 2890 0 1 730
box -6 -8 86 248
use NAND2X1  _1226_
timestamp 0
transform -1 0 3150 0 -1 1690
box -6 -8 86 248
use NOR2X1  _1227_
timestamp 0
transform 1 0 2970 0 1 1210
box -6 -8 86 248
use OAI21X1  _1228_
timestamp 0
transform -1 0 3110 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1229_
timestamp 0
transform 1 0 3070 0 1 730
box -6 -8 106 248
use INVX1  _1230_
timestamp 0
transform 1 0 3270 0 -1 730
box -6 -8 66 248
use INVX1  _1231_
timestamp 0
transform 1 0 1970 0 -1 250
box -6 -8 66 248
use OAI21X1  _1232_
timestamp 0
transform 1 0 2070 0 -1 250
box -6 -8 106 248
use NAND3X1  _1233_
timestamp 0
transform -1 0 2610 0 1 250
box -6 -8 106 248
use AOI21X1  _1234_
timestamp 0
transform 1 0 1230 0 -1 250
box -6 -8 106 248
use NOR3X1  _1235_
timestamp 0
transform 1 0 1370 0 -1 250
box -6 -8 186 248
use OAI21X1  _1236_
timestamp 0
transform -1 0 390 0 -1 250
box -6 -8 106 248
use NAND3X1  _1237_
timestamp 0
transform 1 0 570 0 -1 250
box -6 -8 106 248
use NAND3X1  _1238_
timestamp 0
transform 1 0 710 0 -1 250
box -6 -8 106 248
use NAND3X1  _1239_
timestamp 0
transform 1 0 2010 0 1 250
box -6 -8 106 248
use INVX1  _1240_
timestamp 0
transform -1 0 2170 0 1 1210
box -6 -8 66 248
use OAI21X1  _1241_
timestamp 0
transform 1 0 1730 0 -1 1210
box -6 -8 106 248
use AOI21X1  _1242_
timestamp 0
transform 1 0 2210 0 1 1210
box -6 -8 106 248
use OAI21X1  _1243_
timestamp 0
transform -1 0 2770 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1244_
timestamp 0
transform -1 0 1410 0 1 1690
box -6 -8 106 248
use NAND2X1  _1245_
timestamp 0
transform -1 0 950 0 -1 2650
box -6 -8 86 248
use OAI21X1  _1246_
timestamp 0
transform -1 0 570 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1247_
timestamp 0
transform 1 0 2410 0 1 3610
box -6 -8 86 248
use INVX1  _1248_
timestamp 0
transform -1 0 1450 0 1 3610
box -6 -8 66 248
use NOR2X1  _1249_
timestamp 0
transform -1 0 2370 0 1 3610
box -6 -8 86 248
use OAI21X1  _1250_
timestamp 0
transform -1 0 2190 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1251_
timestamp 0
transform 1 0 2030 0 1 3610
box -6 -8 86 248
use OR2X2  _1252_
timestamp 0
transform -1 0 1870 0 1 3610
box -6 -8 106 248
use NAND3X1  _1253_
timestamp 0
transform -1 0 1350 0 1 3610
box -6 -8 106 248
use AND2X2  _1254_
timestamp 0
transform 1 0 2150 0 1 3610
box -6 -8 106 248
use NOR2X1  _1255_
timestamp 0
transform 1 0 1910 0 1 3610
box -6 -8 86 248
use OAI21X1  _1256_
timestamp 0
transform -1 0 1730 0 1 3610
box -6 -8 106 248
use NAND2X1  _1257_
timestamp 0
transform -1 0 1050 0 -1 4090
box -6 -8 86 248
use AOI21X1  _1258_
timestamp 0
transform 1 0 190 0 -1 2650
box -6 -8 106 248
use NAND2X1  _1259_
timestamp 0
transform 1 0 2030 0 1 4090
box -6 -8 86 248
use AND2X2  _1260_
timestamp 0
transform -1 0 1970 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1261_
timestamp 0
transform -1 0 1990 0 1 4090
box -6 -8 106 248
use AND2X2  _1262_
timestamp 0
transform -1 0 2530 0 1 4090
box -6 -8 106 248
use OAI21X1  _1263_
timestamp 0
transform -1 0 2250 0 1 4090
box -6 -8 106 248
use NAND3X1  _1264_
timestamp 0
transform -1 0 1730 0 1 4090
box -6 -8 106 248
use INVX1  _1265_
timestamp 0
transform -1 0 1350 0 1 4090
box -6 -8 66 248
use NAND2X1  _1266_
timestamp 0
transform 1 0 1770 0 1 4090
box -6 -8 86 248
use AOI22X1  _1267_
timestamp 0
transform 1 0 2570 0 1 4090
box -6 -8 126 248
use INVX1  _1268_
timestamp 0
transform -1 0 1450 0 1 4090
box -6 -8 66 248
use NAND3X1  _1269_
timestamp 0
transform -1 0 1250 0 1 4090
box -6 -8 106 248
use NAND2X1  _1270_
timestamp 0
transform 1 0 890 0 1 4090
box -6 -8 86 248
use AOI21X1  _1271_
timestamp 0
transform -1 0 550 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1272_
timestamp 0
transform 1 0 1750 0 -1 4090
box -6 -8 86 248
use INVX1  _1273_
timestamp 0
transform 1 0 1490 0 -1 4570
box -6 -8 66 248
use AOI22X1  _1274_
timestamp 0
transform 1 0 1690 0 -1 3610
box -6 -8 126 248
use AOI21X1  _1275_
timestamp 0
transform -1 0 1470 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1276_
timestamp 0
transform -1 0 410 0 1 4090
box -6 -8 86 248
use OAI21X1  _1277_
timestamp 0
transform -1 0 930 0 -1 3130
box -6 -8 106 248
use INVX1  _1278_
timestamp 0
transform 1 0 1650 0 -1 4090
box -6 -8 66 248
use OAI21X1  _1279_
timestamp 0
transform 1 0 1510 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1280_
timestamp 0
transform 1 0 610 0 -1 4090
box -6 -8 86 248
use NAND3X1  _1281_
timestamp 0
transform -1 0 290 0 1 4090
box -6 -8 106 248
use AND2X2  _1282_
timestamp 0
transform 1 0 1010 0 1 4090
box -6 -8 106 248
use NAND2X1  _1283_
timestamp 0
transform 1 0 850 0 -1 4090
box -6 -8 86 248
use NAND2X1  _1284_
timestamp 0
transform -1 0 530 0 -1 4570
box -6 -8 86 248
use NAND3X1  _1285_
timestamp 0
transform -1 0 550 0 1 4090
box -6 -8 106 248
use NAND3X1  _1286_
timestamp 0
transform -1 0 150 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1287_
timestamp 0
transform -1 0 150 0 1 2650
box -6 -8 106 248
use AOI22X1  _1288_
timestamp 0
transform -1 0 850 0 1 4090
box -6 -8 126 248
use AOI21X1  _1289_
timestamp 0
transform -1 0 150 0 1 4090
box -6 -8 106 248
use OAI21X1  _1290_
timestamp 0
transform -1 0 270 0 1 3610
box -6 -8 106 248
use NAND3X1  _1291_
timestamp 0
transform 1 0 190 0 -1 3610
box -6 -8 106 248
use AND2X2  _1292_
timestamp 0
transform -1 0 1210 0 1 3610
box -6 -8 106 248
use NAND3X1  _1293_
timestamp 0
transform 1 0 330 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1294_
timestamp 0
transform -1 0 410 0 1 3610
box -6 -8 106 248
use NAND3X1  _1295_
timestamp 0
transform -1 0 910 0 1 3610
box -6 -8 106 248
use NAND3X1  _1296_
timestamp 0
transform 1 0 330 0 -1 3610
box -6 -8 106 248
use AOI21X1  _1297_
timestamp 0
transform -1 0 430 0 -1 2170
box -6 -8 106 248
use AOI22X1  _1298_
timestamp 0
transform -1 0 1070 0 1 3610
box -6 -8 126 248
use AOI21X1  _1299_
timestamp 0
transform -1 0 150 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1300_
timestamp 0
transform -1 0 150 0 1 3130
box -6 -8 106 248
use AOI21X1  _1301_
timestamp 0
transform 1 0 850 0 1 3130
box -6 -8 106 248
use INVX1  _1302_
timestamp 0
transform -1 0 810 0 1 3130
box -6 -8 66 248
use NAND3X1  _1303_
timestamp 0
transform 1 0 330 0 1 3130
box -6 -8 106 248
use OAI21X1  _1304_
timestamp 0
transform 1 0 190 0 1 3130
box -6 -8 106 248
use AOI21X1  _1305_
timestamp 0
transform 1 0 610 0 1 3130
box -6 -8 106 248
use OAI21X1  _1306_
timestamp 0
transform 1 0 990 0 1 3130
box -6 -8 106 248
use OAI21X1  _1307_
timestamp 0
transform 1 0 1170 0 1 1690
box -6 -8 106 248
use NAND3X1  _1308_
timestamp 0
transform -1 0 570 0 1 3130
box -6 -8 106 248
use NAND3X1  _1309_
timestamp 0
transform 1 0 750 0 -1 3610
box -6 -8 106 248
use NAND3X1  _1310_
timestamp 0
transform 1 0 1130 0 1 3130
box -6 -8 106 248
use AND2X2  _1311_
timestamp 0
transform 1 0 2310 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1312_
timestamp 0
transform 1 0 2410 0 1 2650
box -6 -8 86 248
use NAND3X1  _1313_
timestamp 0
transform 1 0 2150 0 -1 1690
box -6 -8 106 248
use INVX1  _1314_
timestamp 0
transform 1 0 1870 0 -1 1210
box -6 -8 66 248
use NAND2X1  _1315_
timestamp 0
transform 1 0 1470 0 -1 1210
box -6 -8 86 248
use NAND3X1  _1316_
timestamp 0
transform 1 0 1590 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1317_
timestamp 0
transform 1 0 1970 0 -1 1210
box -6 -8 106 248
use AOI21X1  _1318_
timestamp 0
transform 1 0 2110 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1319_
timestamp 0
transform 1 0 2390 0 -1 1210
box -6 -8 106 248
use AOI21X1  _1320_
timestamp 0
transform -1 0 2390 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1321_
timestamp 0
transform -1 0 2210 0 1 3130
box -6 -8 86 248
use NAND2X1  _1322_
timestamp 0
transform -1 0 2530 0 -1 3130
box -6 -8 86 248
use AND2X2  _1323_
timestamp 0
transform 1 0 2510 0 -1 2650
box -6 -8 106 248
use NOR2X1  _1324_
timestamp 0
transform 1 0 3470 0 1 1690
box -6 -8 86 248
use NOR2X1  _1325_
timestamp 0
transform -1 0 3410 0 1 2170
box -6 -8 86 248
use OAI21X1  _1326_
timestamp 0
transform 1 0 3270 0 -1 2650
box -6 -8 106 248
use AOI21X1  _1327_
timestamp 0
transform 1 0 3410 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1328_
timestamp 0
transform -1 0 3790 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1329_
timestamp 0
transform -1 0 3650 0 -1 2650
box -6 -8 106 248
use NAND2X1  _1330_
timestamp 0
transform 1 0 3550 0 1 2650
box -6 -8 86 248
use OAI21X1  _1331_
timestamp 0
transform 1 0 3410 0 1 2650
box -6 -8 106 248
use INVX1  _1332_
timestamp 0
transform 1 0 2770 0 -1 2650
box -6 -8 66 248
use INVX1  _1333_
timestamp 0
transform -1 0 2890 0 1 2170
box -6 -8 66 248
use OAI21X1  _1334_
timestamp 0
transform 1 0 3470 0 1 3130
box -6 -8 106 248
use OAI21X1  _1335_
timestamp 0
transform 1 0 2930 0 1 2650
box -6 -8 106 248
use AOI21X1  _1336_
timestamp 0
transform 1 0 470 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1337_
timestamp 0
transform 1 0 610 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1338_
timestamp 0
transform -1 0 1590 0 1 3610
box -6 -8 106 248
use AOI21X1  _1339_
timestamp 0
transform 1 0 190 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1340_
timestamp 0
transform 1 0 470 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1341_
timestamp 0
transform -1 0 1430 0 -1 5050
box -6 -8 86 248
use INVX1  _1342_
timestamp 0
transform 1 0 850 0 -1 5050
box -6 -8 66 248
use NOR2X1  _1343_
timestamp 0
transform -1 0 1550 0 -1 5050
box -6 -8 86 248
use OAI21X1  _1344_
timestamp 0
transform -1 0 1590 0 1 4090
box -6 -8 106 248
use NAND2X1  _1345_
timestamp 0
transform 1 0 1090 0 -1 5050
box -6 -8 86 248
use OR2X2  _1346_
timestamp 0
transform 1 0 1210 0 -1 5050
box -6 -8 106 248
use NAND3X1  _1347_
timestamp 0
transform 1 0 950 0 -1 5050
box -6 -8 106 248
use AND2X2  _1348_
timestamp 0
transform -1 0 1090 0 1 5050
box -6 -8 106 248
use NOR2X1  _1349_
timestamp 0
transform 1 0 1130 0 1 5050
box -6 -8 86 248
use OAI21X1  _1350_
timestamp 0
transform -1 0 810 0 1 5050
box -6 -8 106 248
use NAND2X1  _1351_
timestamp 0
transform 1 0 730 0 -1 5050
box -6 -8 86 248
use NOR2X1  _1352_
timestamp 0
transform -1 0 410 0 -1 4570
box -6 -8 86 248
use AOI21X1  _1353_
timestamp 0
transform -1 0 290 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1354_
timestamp 0
transform 1 0 2090 0 -1 4570
box -6 -8 86 248
use INVX1  _1355_
timestamp 0
transform 1 0 2130 0 1 4570
box -6 -8 66 248
use AND2X2  _1356_
timestamp 0
transform -1 0 2570 0 -1 4570
box -6 -8 106 248
use AND2X2  _1357_
timestamp 0
transform -1 0 3210 0 1 4090
box -6 -8 106 248
use NAND2X1  _1358_
timestamp 0
transform -1 0 2430 0 -1 4570
box -6 -8 86 248
use AOI22X1  _1359_
timestamp 0
transform 1 0 2730 0 1 4090
box -6 -8 126 248
use INVX1  _1360_
timestamp 0
transform 1 0 2230 0 1 4570
box -6 -8 66 248
use AOI21X1  _1361_
timestamp 0
transform -1 0 2090 0 1 4570
box -6 -8 106 248
use INVX2  _1362_
timestamp 0
transform 1 0 3270 0 -1 4570
box -6 -8 66 248
use OAI21X1  _1363_
timestamp 0
transform -1 0 2310 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1364_
timestamp 0
transform 1 0 2290 0 1 4090
box -6 -8 106 248
use AOI21X1  _1365_
timestamp 0
transform -1 0 1910 0 -1 4570
box -6 -8 106 248
use OAI22X1  _1366_
timestamp 0
transform 1 0 1690 0 1 4570
box -6 -8 126 248
use NAND3X1  _1367_
timestamp 0
transform -1 0 2050 0 -1 4570
box -6 -8 106 248
use NAND3X1  _1368_
timestamp 0
transform -1 0 1950 0 1 4570
box -6 -8 106 248
use NOR2X1  _1369_
timestamp 0
transform -1 0 1510 0 1 4570
box -6 -8 86 248
use NAND3X1  _1370_
timestamp 0
transform -1 0 1650 0 1 4570
box -6 -8 106 248
use NAND2X1  _1371_
timestamp 0
transform -1 0 130 0 -1 5050
box -6 -8 86 248
use NOR2X1  _1372_
timestamp 0
transform -1 0 130 0 1 5050
box -6 -8 86 248
use NOR2X1  _1373_
timestamp 0
transform 1 0 730 0 -1 4090
box -6 -8 86 248
use OAI21X1  _1374_
timestamp 0
transform -1 0 690 0 1 4090
box -6 -8 106 248
use AOI21X1  _1375_
timestamp 0
transform -1 0 550 0 -1 5050
box -6 -8 106 248
use OAI21X1  _1376_
timestamp 0
transform -1 0 270 0 -1 5050
box -6 -8 106 248
use AND2X2  _1377_
timestamp 0
transform -1 0 670 0 1 5050
box -6 -8 106 248
use NAND3X1  _1378_
timestamp 0
transform -1 0 690 0 -1 5050
box -6 -8 106 248
use NAND2X1  _1379_
timestamp 0
transform -1 0 250 0 1 5050
box -6 -8 86 248
use NAND3X1  _1380_
timestamp 0
transform 1 0 430 0 1 5050
box -6 -8 106 248
use NAND3X1  _1381_
timestamp 0
transform 1 0 750 0 1 4570
box -6 -8 106 248
use NOR3X1  _1382_
timestamp 0
transform 1 0 450 0 1 3610
box -6 -8 186 248
use AOI21X1  _1383_
timestamp 0
transform -1 0 770 0 1 3610
box -6 -8 106 248
use AOI21X1  _1384_
timestamp 0
transform -1 0 390 0 1 5050
box -6 -8 106 248
use NAND3X1  _1385_
timestamp 0
transform -1 0 150 0 1 4570
box -6 -8 106 248
use OAI21X1  _1386_
timestamp 0
transform -1 0 150 0 -1 4570
box -6 -8 106 248
use AOI21X1  _1387_
timestamp 0
transform 1 0 190 0 1 4570
box -6 -8 106 248
use OAI21X1  _1388_
timestamp 0
transform 1 0 470 0 1 4570
box -6 -8 106 248
use NAND3X1  _1389_
timestamp 0
transform 1 0 1090 0 -1 4570
box -6 -8 106 248
use INVX1  _1390_
timestamp 0
transform 1 0 850 0 -1 4570
box -6 -8 66 248
use NAND3X1  _1391_
timestamp 0
transform 1 0 610 0 1 4570
box -6 -8 106 248
use OAI21X1  _1392_
timestamp 0
transform 1 0 330 0 1 4570
box -6 -8 106 248
use NAND3X1  _1393_
timestamp 0
transform 1 0 710 0 -1 4570
box -6 -8 106 248
use AOI21X1  _1394_
timestamp 0
transform 1 0 1230 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1395_
timestamp 0
transform 1 0 950 0 -1 4570
box -6 -8 106 248
use NAND3X1  _1396_
timestamp 0
transform -1 0 670 0 -1 4570
box -6 -8 106 248
use AOI22X1  _1397_
timestamp 0
transform 1 0 1130 0 -1 3610
box -6 -8 126 248
use NOR2X1  _1398_
timestamp 0
transform 1 0 1970 0 -1 3610
box -6 -8 86 248
use AOI21X1  _1399_
timestamp 0
transform 1 0 2530 0 1 2650
box -6 -8 106 248
use OAI21X1  _1400_
timestamp 0
transform -1 0 2670 0 -1 3130
box -6 -8 106 248
use INVX1  _1401_
timestamp 0
transform -1 0 1090 0 -1 3610
box -6 -8 66 248
use AOI21X1  _1402_
timestamp 0
transform 1 0 890 0 -1 3610
box -6 -8 106 248
use NAND3X1  _1403_
timestamp 0
transform 1 0 1290 0 -1 3610
box -6 -8 106 248
use NAND3X1  _1404_
timestamp 0
transform -1 0 1190 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1405_
timestamp 0
transform -1 0 1930 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1406_
timestamp 0
transform 1 0 2710 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1407_
timestamp 0
transform 1 0 2790 0 1 2650
box -6 -8 106 248
use AND2X2  _1408_
timestamp 0
transform 1 0 3190 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1409_
timestamp 0
transform 1 0 3610 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1410_
timestamp 0
transform 1 0 3330 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1411_
timestamp 0
transform 1 0 3470 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1412_
timestamp 0
transform -1 0 3030 0 1 1690
box -6 -8 106 248
use AOI22X1  _1413_
timestamp 0
transform 1 0 2870 0 -1 2650
box -6 -8 126 248
use OAI21X1  _1414_
timestamp 0
transform 1 0 3950 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1415_
timestamp 0
transform 1 0 2370 0 1 3130
box -6 -8 106 248
use AOI21X1  _1416_
timestamp 0
transform 1 0 2450 0 -1 3610
box -6 -8 106 248
use INVX1  _1417_
timestamp 0
transform 1 0 2590 0 -1 3610
box -6 -8 66 248
use OAI21X1  _1418_
timestamp 0
transform 1 0 850 0 1 5050
box -6 -8 106 248
use INVX1  _1419_
timestamp 0
transform -1 0 670 0 -1 5530
box -6 -8 66 248
use AOI21X1  _1420_
timestamp 0
transform -1 0 150 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1421_
timestamp 0
transform -1 0 1670 0 -1 5050
box -6 -8 86 248
use INVX1  _1422_
timestamp 0
transform 1 0 1710 0 -1 5050
box -6 -8 66 248
use NOR2X1  _1423_
timestamp 0
transform 1 0 2210 0 -1 5050
box -6 -8 86 248
use OAI21X1  _1424_
timestamp 0
transform 1 0 2330 0 1 4570
box -6 -8 106 248
use NAND2X1  _1425_
timestamp 0
transform 1 0 2090 0 -1 5050
box -6 -8 86 248
use OR2X2  _1426_
timestamp 0
transform -1 0 2050 0 -1 5050
box -6 -8 106 248
use NAND3X1  _1427_
timestamp 0
transform -1 0 1910 0 -1 5050
box -6 -8 106 248
use AND2X2  _1428_
timestamp 0
transform 1 0 2450 0 1 5050
box -6 -8 106 248
use NOR2X1  _1429_
timestamp 0
transform 1 0 2330 0 1 5050
box -6 -8 86 248
use OAI21X1  _1430_
timestamp 0
transform -1 0 2290 0 1 5050
box -6 -8 106 248
use NAND2X1  _1431_
timestamp 0
transform 1 0 1410 0 -1 5530
box -6 -8 86 248
use NAND2X1  _1432_
timestamp 0
transform 1 0 1370 0 -1 4570
box -6 -8 86 248
use NAND2X1  _1433_
timestamp 0
transform 1 0 2570 0 1 4570
box -6 -8 86 248
use INVX1  _1434_
timestamp 0
transform 1 0 2730 0 1 5050
box -6 -8 66 248
use NAND2X1  _1435_
timestamp 0
transform 1 0 2770 0 -1 4570
box -6 -8 86 248
use NAND2X1  _1436_
timestamp 0
transform 1 0 3350 0 1 4570
box -6 -8 86 248
use NOR2X1  _1437_
timestamp 0
transform 1 0 2670 0 -1 5050
box -6 -8 86 248
use INVX1  _1438_
timestamp 0
transform -1 0 2630 0 -1 5050
box -6 -8 66 248
use AOI22X1  _1439_
timestamp 0
transform -1 0 2730 0 -1 4570
box -6 -8 126 248
use INVX1  _1440_
timestamp 0
transform 1 0 2470 0 -1 5050
box -6 -8 66 248
use NAND3X1  _1441_
timestamp 0
transform -1 0 2690 0 1 5050
box -6 -8 106 248
use OAI21X1  _1442_
timestamp 0
transform -1 0 2430 0 -1 5050
box -6 -8 106 248
use NAND2X1  _1443_
timestamp 0
transform 1 0 1930 0 1 5050
box -6 -8 86 248
use AOI21X1  _1444_
timestamp 0
transform -1 0 1350 0 1 5050
box -6 -8 106 248
use NAND3X1  _1445_
timestamp 0
transform -1 0 1490 0 1 5050
box -6 -8 106 248
use INVX1  _1446_
timestamp 0
transform -1 0 810 0 1 5530
box -6 -8 66 248
use OAI21X1  _1447_
timestamp 0
transform -1 0 710 0 1 5530
box -6 -8 106 248
use AND2X2  _1448_
timestamp 0
transform -1 0 1750 0 1 5050
box -6 -8 106 248
use NAND2X1  _1449_
timestamp 0
transform 1 0 1530 0 1 5050
box -6 -8 86 248
use NAND3X1  _1450_
timestamp 0
transform -1 0 1890 0 1 5050
box -6 -8 106 248
use NAND3X1  _1451_
timestamp 0
transform -1 0 950 0 1 5530
box -6 -8 106 248
use NAND3X1  _1452_
timestamp 0
transform -1 0 150 0 1 5530
box -6 -8 106 248
use OAI21X1  _1453_
timestamp 0
transform 1 0 310 0 -1 5050
box -6 -8 106 248
use AOI22X1  _1454_
timestamp 0
transform -1 0 1370 0 -1 5530
box -6 -8 126 248
use OR2X2  _1455_
timestamp 0
transform -1 0 1090 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1456_
timestamp 0
transform 1 0 1130 0 -1 5530
box -6 -8 86 248
use AOI21X1  _1457_
timestamp 0
transform -1 0 950 0 -1 5530
box -6 -8 106 248
use OAI21X1  _1458_
timestamp 0
transform -1 0 430 0 -1 5530
box -6 -8 106 248
use NAND3X1  _1459_
timestamp 0
transform -1 0 290 0 -1 5530
box -6 -8 106 248
use NAND3X1  _1460_
timestamp 0
transform 1 0 190 0 1 5530
box -6 -8 106 248
use OAI21X1  _1461_
timestamp 0
transform -1 0 570 0 -1 5530
box -6 -8 106 248
use NAND3X1  _1462_
timestamp 0
transform 1 0 710 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1463_
timestamp 0
transform -1 0 1250 0 1 4570
box -6 -8 86 248
use NAND3X1  _1464_
timestamp 0
transform 1 0 1230 0 -1 4570
box -6 -8 106 248
use AOI21X1  _1465_
timestamp 0
transform 1 0 890 0 1 4570
box -6 -8 106 248
use OAI21X1  _1466_
timestamp 0
transform 1 0 1030 0 1 4570
box -6 -8 106 248
use NAND3X1  _1467_
timestamp 0
transform 1 0 1290 0 1 4570
box -6 -8 106 248
use NAND2X1  _1468_
timestamp 0
transform -1 0 1670 0 -1 4570
box -6 -8 86 248
use AOI21X1  _1469_
timestamp 0
transform 1 0 2510 0 1 3130
box -6 -8 106 248
use NAND2X1  _1470_
timestamp 0
transform -1 0 2330 0 1 3130
box -6 -8 86 248
use OAI21X1  _1471_
timestamp 0
transform -1 0 2750 0 1 3130
box -6 -8 106 248
use INVX1  _1472_
timestamp 0
transform -1 0 2970 0 1 3130
box -6 -8 66 248
use NOR2X1  _1473_
timestamp 0
transform -1 0 2870 0 1 3130
box -6 -8 86 248
use OAI21X1  _1474_
timestamp 0
transform 1 0 2850 0 -1 3130
box -6 -8 106 248
use NOR2X1  _1475_
timestamp 0
transform 1 0 3350 0 1 1690
box -6 -8 86 248
use NOR2X1  _1476_
timestamp 0
transform -1 0 3010 0 1 2170
box -6 -8 86 248
use AOI21X1  _1477_
timestamp 0
transform 1 0 3150 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1478_
timestamp 0
transform 1 0 3290 0 -1 1210
box -6 -8 106 248
use NOR2X1  _1479_
timestamp 0
transform 1 0 3630 0 -1 2170
box -6 -8 86 248
use NOR2X1  _1480_
timestamp 0
transform -1 0 3290 0 1 2170
box -6 -8 86 248
use AOI22X1  _1481_
timestamp 0
transform -1 0 3170 0 1 2170
box -6 -8 126 248
use OAI21X1  _1482_
timestamp 0
transform 1 0 4110 0 1 3610
box -6 -8 106 248
use INVX1  _1483_
timestamp 0
transform -1 0 2650 0 -1 250
box -6 -8 66 248
use INVX1  _1484_
timestamp 0
transform -1 0 3450 0 -1 250
box -6 -8 66 248
use OAI21X1  _1485_
timestamp 0
transform 1 0 3370 0 -1 3130
box -6 -8 106 248
use INVX1  _1486_
timestamp 0
transform 1 0 2950 0 -1 3610
box -6 -8 66 248
use OAI21X1  _1487_
timestamp 0
transform -1 0 2150 0 1 5050
box -6 -8 106 248
use INVX1  _1488_
timestamp 0
transform -1 0 1330 0 1 5530
box -6 -8 66 248
use AOI21X1  _1489_
timestamp 0
transform 1 0 1130 0 1 5530
box -6 -8 106 248
use NAND2X1  _1490_
timestamp 0
transform 1 0 2790 0 -1 5050
box -6 -8 86 248
use INVX1  _1491_
timestamp 0
transform -1 0 3170 0 1 4570
box -6 -8 66 248
use NOR2X1  _1492_
timestamp 0
transform 1 0 2910 0 -1 4570
box -6 -8 86 248
use OAI22X1  _1493_
timestamp 0
transform -1 0 2810 0 1 4570
box -6 -8 126 248
use NAND2X1  _1494_
timestamp 0
transform -1 0 2930 0 1 4570
box -6 -8 86 248
use OR2X2  _1495_
timestamp 0
transform 1 0 2970 0 1 4570
box -6 -8 106 248
use NAND3X1  _1496_
timestamp 0
transform 1 0 3210 0 1 4570
box -6 -8 106 248
use INVX2  _1497_
timestamp 0
transform -1 0 3530 0 1 4570
box -6 -8 66 248
use NAND2X1  _1498_
timestamp 0
transform 1 0 3050 0 -1 5050
box -6 -8 86 248
use OAI21X1  _1499_
timestamp 0
transform -1 0 3270 0 -1 5050
box -6 -8 106 248
use NAND2X1  _1500_
timestamp 0
transform -1 0 3870 0 -1 4570
box -6 -8 86 248
use NAND2X1  _1501_
timestamp 0
transform 1 0 4150 0 1 4570
box -6 -8 86 248
use NOR2X1  _1502_
timestamp 0
transform 1 0 4030 0 1 4570
box -6 -8 86 248
use INVX1  _1503_
timestamp 0
transform 1 0 4430 0 1 5050
box -6 -8 66 248
use INVX1  _1504_
timestamp 0
transform -1 0 3970 0 1 5050
box -6 -8 66 248
use OAI21X1  _1505_
timestamp 0
transform -1 0 3730 0 1 5050
box -6 -8 106 248
use AND2X2  _1506_
timestamp 0
transform -1 0 3870 0 1 5050
box -6 -8 106 248
use AOI21X1  _1507_
timestamp 0
transform 1 0 3350 0 1 5050
box -6 -8 106 248
use INVX1  _1508_
timestamp 0
transform -1 0 1850 0 1 5530
box -6 -8 66 248
use NAND3X1  _1509_
timestamp 0
transform -1 0 3310 0 1 5050
box -6 -8 106 248
use NAND3X1  _1510_
timestamp 0
transform -1 0 1610 0 1 5530
box -6 -8 106 248
use OAI21X1  _1511_
timestamp 0
transform 1 0 990 0 1 5530
box -6 -8 106 248
use INVX1  _1512_
timestamp 0
transform 1 0 2030 0 1 5530
box -6 -8 66 248
use OAI21X1  _1513_
timestamp 0
transform -1 0 1750 0 1 5530
box -6 -8 106 248
use NAND3X1  _1514_
timestamp 0
transform 1 0 1370 0 1 5530
box -6 -8 106 248
use NAND3X1  _1515_
timestamp 0
transform 1 0 1670 0 -1 5530
box -6 -8 106 248
use OAI21X1  _1516_
timestamp 0
transform -1 0 1990 0 1 5530
box -6 -8 106 248
use NAND3X1  _1517_
timestamp 0
transform -1 0 2030 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1518_
timestamp 0
transform -1 0 1890 0 -1 5530
box -6 -8 86 248
use NAND3X1  _1519_
timestamp 0
transform 1 0 1530 0 -1 5530
box -6 -8 106 248
use AOI21X1  _1520_
timestamp 0
transform 1 0 330 0 1 5530
box -6 -8 106 248
use OAI21X1  _1521_
timestamp 0
transform 1 0 470 0 1 5530
box -6 -8 106 248
use NAND3X1  _1522_
timestamp 0
transform 1 0 2070 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1523_
timestamp 0
transform -1 0 2710 0 -1 4090
box -6 -8 86 248
use NOR3X1  _1524_
timestamp 0
transform 1 0 3150 0 1 3130
box -6 -8 186 248
use AOI21X1  _1525_
timestamp 0
transform 1 0 3010 0 1 3130
box -6 -8 106 248
use INVX1  _1526_
timestamp 0
transform -1 0 3050 0 -1 3130
box -6 -8 66 248
use OAI21X1  _1527_
timestamp 0
transform 1 0 3090 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1528_
timestamp 0
transform 1 0 3230 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1529_
timestamp 0
transform 1 0 2650 0 1 250
box -6 -8 86 248
use NAND2X1  _1530_
timestamp 0
transform -1 0 3230 0 -1 730
box -6 -8 86 248
use NAND2X1  _1531_
timestamp 0
transform 1 0 2210 0 -1 250
box -6 -8 86 248
use NAND2X1  _1532_
timestamp 0
transform -1 0 2550 0 -1 250
box -6 -8 86 248
use OAI21X1  _1533_
timestamp 0
transform -1 0 2430 0 -1 250
box -6 -8 106 248
use AOI21X1  _1534_
timestamp 0
transform 1 0 2770 0 1 250
box -6 -8 106 248
use AOI22X1  _1535_
timestamp 0
transform 1 0 2910 0 1 250
box -6 -8 126 248
use INVX1  _1536_
timestamp 0
transform 1 0 3310 0 1 250
box -6 -8 66 248
use NAND2X1  _1537_
timestamp 0
transform 1 0 2210 0 -1 5530
box -6 -8 86 248
use INVX1  _1538_
timestamp 0
transform -1 0 2390 0 -1 5530
box -6 -8 66 248
use OAI21X1  _1539_
timestamp 0
transform -1 0 3010 0 -1 5050
box -6 -8 106 248
use INVX1  _1540_
timestamp 0
transform -1 0 2590 0 1 5530
box -6 -8 66 248
use INVX1  _1541_
timestamp 0
transform 1 0 3570 0 1 4570
box -6 -8 66 248
use NOR2X1  _1542_
timestamp 0
transform 1 0 4010 0 1 5050
box -6 -8 86 248
use NOR2X1  _1543_
timestamp 0
transform 1 0 3910 0 1 4570
box -6 -8 86 248
use NOR2X1  _1544_
timestamp 0
transform 1 0 3930 0 -1 5050
box -6 -8 86 248
use AOI21X1  _1545_
timestamp 0
transform -1 0 4390 0 1 5050
box -6 -8 106 248
use NAND2X1  _1546_
timestamp 0
transform -1 0 3810 0 -1 5530
box -6 -8 86 248
use NOR2X1  _1547_
timestamp 0
transform 1 0 3810 0 -1 5050
box -6 -8 86 248
use OAI22X1  _1548_
timestamp 0
transform 1 0 4130 0 1 5050
box -6 -8 126 248
use NAND2X1  _1549_
timestamp 0
transform -1 0 3490 0 1 5530
box -6 -8 86 248
use OAI21X1  _1550_
timestamp 0
transform -1 0 3590 0 1 5050
box -6 -8 106 248
use INVX1  _1551_
timestamp 0
transform -1 0 3370 0 1 5530
box -6 -8 66 248
use NAND3X1  _1552_
timestamp 0
transform -1 0 3270 0 1 5530
box -6 -8 106 248
use NAND2X1  _1553_
timestamp 0
transform 1 0 2910 0 1 5530
box -6 -8 86 248
use NOR2X1  _1554_
timestamp 0
transform -1 0 2350 0 1 5530
box -6 -8 86 248
use AOI21X1  _1555_
timestamp 0
transform -1 0 2870 0 1 5530
box -6 -8 106 248
use OAI21X1  _1556_
timestamp 0
transform -1 0 2490 0 1 5530
box -6 -8 106 248
use OR2X2  _1557_
timestamp 0
transform -1 0 2230 0 1 5530
box -6 -8 106 248
use INVX1  _1558_
timestamp 0
transform 1 0 2570 0 -1 5530
box -6 -8 66 248
use NAND3X1  _1559_
timestamp 0
transform -1 0 2770 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1560_
timestamp 0
transform 1 0 2830 0 1 5050
box -6 -8 86 248
use NAND2X1  _1561_
timestamp 0
transform 1 0 2950 0 1 5050
box -6 -8 86 248
use NAND3X1  _1562_
timestamp 0
transform 1 0 2430 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1563_
timestamp 0
transform -1 0 3070 0 1 4090
box -6 -8 86 248
use NOR2X1  _1564_
timestamp 0
transform 1 0 2690 0 -1 3610
box -6 -8 86 248
use NOR2X1  _1565_
timestamp 0
transform 1 0 3170 0 1 3610
box -6 -8 86 248
use NAND3X1  _1566_
timestamp 0
transform 1 0 3050 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1567_
timestamp 0
transform -1 0 2710 0 1 3610
box -6 -8 86 248
use AOI22X1  _1568_
timestamp 0
transform 1 0 3010 0 1 3610
box -6 -8 126 248
use AOI21X1  _1569_
timestamp 0
transform 1 0 3190 0 -1 3610
box -6 -8 106 248
use INVX1  _1570_
timestamp 0
transform 1 0 3330 0 -1 3610
box -6 -8 66 248
use NAND2X1  _1571_
timestamp 0
transform -1 0 2970 0 1 3610
box -6 -8 86 248
use OAI21X1  _1572_
timestamp 0
transform 1 0 3290 0 1 3610
box -6 -8 106 248
use AOI21X1  _1573_
timestamp 0
transform -1 0 2850 0 1 3610
box -6 -8 106 248
use OAI21X1  _1574_
timestamp 0
transform 1 0 2810 0 -1 3610
box -6 -8 106 248
use AOI21X1  _1575_
timestamp 0
transform 1 0 3430 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1576_
timestamp 0
transform 1 0 3710 0 -1 3610
box -6 -8 106 248
use OR2X2  _1577_
timestamp 0
transform 1 0 4050 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1578_
timestamp 0
transform -1 0 3850 0 -1 2170
box -6 -8 106 248
use INVX1  _1579_
timestamp 0
transform 1 0 1730 0 -1 250
box -6 -8 66 248
use OAI21X1  _1580_
timestamp 0
transform 1 0 1590 0 -1 250
box -6 -8 106 248
use NAND2X1  _1581_
timestamp 0
transform 1 0 1750 0 1 250
box -6 -8 86 248
use NAND2X1  _1582_
timestamp 0
transform -1 0 3850 0 -1 730
box -6 -8 86 248
use OAI21X1  _1583_
timestamp 0
transform 1 0 3630 0 -1 730
box -6 -8 106 248
use AOI21X1  _1584_
timestamp 0
transform -1 0 3590 0 -1 730
box -6 -8 106 248
use AOI22X1  _1585_
timestamp 0
transform 1 0 3410 0 1 250
box -6 -8 126 248
use INVX1  _1586_
timestamp 0
transform -1 0 3650 0 -1 1210
box -6 -8 66 248
use AOI21X1  _1587_
timestamp 0
transform -1 0 3950 0 -1 5530
box -6 -8 106 248
use NOR2X1  _1588_
timestamp 0
transform 1 0 3670 0 1 4570
box -6 -8 86 248
use NAND2X1  _1589_
timestamp 0
transform -1 0 3870 0 1 4570
box -6 -8 86 248
use OAI22X1  _1590_
timestamp 0
transform -1 0 3530 0 -1 5050
box -6 -8 126 248
use NAND2X1  _1591_
timestamp 0
transform 1 0 3570 0 -1 5050
box -6 -8 86 248
use OR2X2  _1592_
timestamp 0
transform 1 0 3030 0 1 5530
box -6 -8 106 248
use OAI21X1  _1593_
timestamp 0
transform -1 0 3690 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1594_
timestamp 0
transform -1 0 3550 0 -1 5530
box -6 -8 86 248
use NAND2X1  _1595_
timestamp 0
transform 1 0 3210 0 -1 5530
box -6 -8 86 248
use OR2X2  _1596_
timestamp 0
transform -1 0 3170 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1597_
timestamp 0
transform -1 0 3030 0 -1 5530
box -6 -8 86 248
use NAND3X1  _1598_
timestamp 0
transform 1 0 3070 0 1 5050
box -6 -8 106 248
use OAI21X1  _1599_
timestamp 0
transform 1 0 2630 0 1 5530
box -6 -8 106 248
use NAND3X1  _1600_
timestamp 0
transform -1 0 2910 0 -1 5530
box -6 -8 106 248
use NAND2X1  _1601_
timestamp 0
transform 1 0 3150 0 -1 4570
box -6 -8 86 248
use NOR2X1  _1602_
timestamp 0
transform -1 0 3510 0 1 3610
box -6 -8 86 248
use NAND3X1  _1603_
timestamp 0
transform 1 0 3550 0 1 3610
box -6 -8 106 248
use NAND3X1  _1604_
timestamp 0
transform 1 0 3570 0 -1 3610
box -6 -8 106 248
use NAND3X1  _1605_
timestamp 0
transform 1 0 3690 0 1 3610
box -6 -8 106 248
use INVX1  _1606_
timestamp 0
transform -1 0 3430 0 1 3130
box -6 -8 66 248
use OR2X2  _1607_
timestamp 0
transform -1 0 2850 0 -1 4090
box -6 -8 106 248
use AND2X2  _1608_
timestamp 0
transform 1 0 3970 0 1 3610
box -6 -8 106 248
use NAND3X1  _1609_
timestamp 0
transform 1 0 3830 0 1 3610
box -6 -8 106 248
use AOI21X1  _1610_
timestamp 0
transform 1 0 1870 0 1 250
box -6 -8 106 248
use OAI21X1  _1611_
timestamp 0
transform 1 0 2530 0 1 730
box -6 -8 106 248
use INVX1  _1612_
timestamp 0
transform -1 0 3670 0 1 730
box -6 -8 66 248
use AOI21X1  _1613_
timestamp 0
transform -1 0 3570 0 1 730
box -6 -8 106 248
use AOI21X1  _1614_
timestamp 0
transform 1 0 3330 0 1 730
box -6 -8 106 248
use AOI22X1  _1615_
timestamp 0
transform -1 0 3550 0 -1 1210
box -6 -8 126 248
use INVX1  _1616_
timestamp 0
transform -1 0 3310 0 1 1210
box -6 -8 66 248
use OAI21X1  _1617_
timestamp 0
transform -1 0 3350 0 1 4090
box -6 -8 106 248
use INVX1  _1618_
timestamp 0
transform -1 0 3370 0 -1 4090
box -6 -8 66 248
use OAI21X1  _1619_
timestamp 0
transform -1 0 3430 0 -1 5530
box -6 -8 106 248
use INVX1  _1620_
timestamp 0
transform -1 0 3370 0 -1 5050
box -6 -8 66 248
use OAI21X1  _1621_
timestamp 0
transform 1 0 3370 0 -1 4570
box -6 -8 106 248
use OR2X2  _1622_
timestamp 0
transform 1 0 3510 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1623_
timestamp 0
transform 1 0 3750 0 1 4090
box -6 -8 86 248
use NAND2X1  _1624_
timestamp 0
transform -1 0 3710 0 1 4090
box -6 -8 86 248
use NAND3X1  _1625_
timestamp 0
transform -1 0 3510 0 -1 4090
box -6 -8 106 248
use OR2X2  _1626_
timestamp 0
transform -1 0 2990 0 -1 4090
box -6 -8 106 248
use AOI21X1  _1627_
timestamp 0
transform -1 0 3130 0 -1 4090
box -6 -8 106 248
use INVX1  _1628_
timestamp 0
transform -1 0 3590 0 1 4090
box -6 -8 66 248
use OAI21X1  _1629_
timestamp 0
transform 1 0 3390 0 1 4090
box -6 -8 106 248
use NAND3X1  _1630_
timestamp 0
transform -1 0 3270 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1631_
timestamp 0
transform 1 0 2530 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1632_
timestamp 0
transform 1 0 2250 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1633_
timestamp 0
transform 1 0 2670 0 -1 1210
box -6 -8 86 248
use NAND2X1  _1634_
timestamp 0
transform -1 0 3450 0 -1 730
box -6 -8 86 248
use OAI21X1  _1635_
timestamp 0
transform 1 0 2670 0 1 730
box -6 -8 106 248
use AOI21X1  _1636_
timestamp 0
transform 1 0 2930 0 1 730
box -6 -8 106 248
use AOI22X1  _1637_
timestamp 0
transform -1 0 3210 0 1 1210
box -6 -8 126 248
use INVX1  _1638_
timestamp 0
transform -1 0 3890 0 -1 1690
box -6 -8 66 248
use AOI21X1  _1639_
timestamp 0
transform 1 0 3550 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1640_
timestamp 0
transform 1 0 3650 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1641_
timestamp 0
transform 1 0 3690 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1642_
timestamp 0
transform 1 0 2430 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1643_
timestamp 0
transform 1 0 2810 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1644_
timestamp 0
transform 1 0 2950 0 -1 1690
box -6 -8 86 248
use NAND2X1  _1645_
timestamp 0
transform 1 0 3230 0 -1 2170
box -6 -8 86 248
use OAI21X1  _1646_
timestamp 0
transform 1 0 3090 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1647_
timestamp 0
transform 1 0 3350 0 -1 2170
box -6 -8 106 248
use AOI22X1  _1648_
timestamp 0
transform -1 0 3850 0 1 1690
box -6 -8 126 248
use NAND2X1  _1649_
timestamp 0
transform 1 0 4730 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1650_
timestamp 0
transform 1 0 4590 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1651_
timestamp 0
transform 1 0 5110 0 1 3610
box -6 -8 86 248
use OAI21X1  _1652_
timestamp 0
transform 1 0 4970 0 1 3610
box -6 -8 106 248
use NAND2X1  _1653_
timestamp 0
transform 1 0 4590 0 -1 4090
box -6 -8 86 248
use OAI21X1  _1654_
timestamp 0
transform -1 0 4810 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1655_
timestamp 0
transform 1 0 4990 0 -1 4090
box -6 -8 86 248
use OAI21X1  _1656_
timestamp 0
transform 1 0 4850 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1657_
timestamp 0
transform 1 0 5610 0 -1 5050
box -6 -8 86 248
use OAI21X1  _1658_
timestamp 0
transform 1 0 5470 0 -1 5050
box -6 -8 106 248
use NAND2X1  _1659_
timestamp 0
transform 1 0 4970 0 1 4570
box -6 -8 86 248
use OAI21X1  _1660_
timestamp 0
transform -1 0 5190 0 1 4570
box -6 -8 106 248
use NAND2X1  _1661_
timestamp 0
transform 1 0 5250 0 -1 4090
box -6 -8 86 248
use OAI21X1  _1662_
timestamp 0
transform 1 0 5110 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1663_
timestamp 0
transform 1 0 5030 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1664_
timestamp 0
transform -1 0 4990 0 -1 4570
box -6 -8 106 248
use DFFPOSX1  _1665_
timestamp 0
transform -1 0 4050 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _1666_
timestamp 0
transform -1 0 3810 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _1667_
timestamp 0
transform -1 0 4690 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _1668_
timestamp 0
transform -1 0 4670 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _1669_
timestamp 0
transform -1 0 5470 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _1670_
timestamp 0
transform -1 0 4950 0 -1 5050
box -6 -8 246 248
use DFFPOSX1  _1671_
timestamp 0
transform 1 0 4230 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _1672_
timestamp 0
transform -1 0 5510 0 1 5530
box -6 -8 246 248
use DFFPOSX1  _1673_
timestamp 0
transform -1 0 3370 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _1674_
timestamp 0
transform -1 0 3230 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _1675_
timestamp 0
transform -1 0 4450 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _1676_
timestamp 0
transform -1 0 3270 0 1 250
box -6 -8 246 248
use DFFPOSX1  _1677_
timestamp 0
transform 1 0 2870 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _1678_
timestamp 0
transform -1 0 3890 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _1679_
timestamp 0
transform -1 0 3550 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _1680_
timestamp 0
transform -1 0 4130 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _1681_
timestamp 0
transform -1 0 5050 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1682_
timestamp 0
transform -1 0 4930 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _1683_
timestamp 0
transform -1 0 5210 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _1684_
timestamp 0
transform 1 0 4790 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _1685_
timestamp 0
transform 1 0 5410 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _1686_
timestamp 0
transform -1 0 4930 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _1687_
timestamp 0
transform -1 0 5530 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _1688_
timestamp 0
transform -1 0 4850 0 -1 4570
box -6 -8 246 248
use DFFSR  _1689_
timestamp 0
transform -1 0 4210 0 1 5530
box -6 -8 486 248
use DFFSR  _1690_
timestamp 0
transform 1 0 5070 0 1 5050
box -6 -8 486 248
use DFFSR  _1691_
timestamp 0
transform -1 0 4810 0 1 5530
box -6 -8 486 248
use INVX1  _1692_
timestamp 0
transform 1 0 5370 0 -1 3610
box -6 -8 66 248
use INVX4  _1693_
timestamp 0
transform 1 0 5470 0 -1 4090
box -6 -8 86 248
use OAI21X1  _1694_
timestamp 0
transform 1 0 5470 0 -1 3610
box -6 -8 106 248
use NOR2X1  _1695_
timestamp 0
transform -1 0 5670 0 1 3130
box -6 -8 86 248
use INVX1  _1696_
timestamp 0
transform 1 0 5650 0 -1 250
box -6 -8 66 248
use INVX2  _1697_
timestamp 0
transform -1 0 5310 0 1 2650
box -6 -8 66 248
use NAND2X1  _1698_
timestamp 0
transform -1 0 5430 0 1 2650
box -6 -8 86 248
use INVX2  _1699_
timestamp 0
transform -1 0 5210 0 1 2650
box -6 -8 66 248
use NAND2X1  _1700_
timestamp 0
transform -1 0 4530 0 -1 3130
box -6 -8 86 248
use NAND2X1  _1701_
timestamp 0
transform -1 0 4630 0 1 3130
box -6 -8 86 248
use AOI22X1  _1702_
timestamp 0
transform 1 0 4570 0 -1 3130
box -6 -8 126 248
use INVX2  _1703_
timestamp 0
transform 1 0 5550 0 1 5530
box -6 -8 66 248
use INVX1  _1704_
timestamp 0
transform 1 0 4790 0 -1 2650
box -6 -8 66 248
use INVX1  _1705_
timestamp 0
transform 1 0 4410 0 1 1690
box -6 -8 66 248
use OAI21X1  _1706_
timestamp 0
transform -1 0 4830 0 1 2650
box -6 -8 106 248
use NAND2X1  _1707_
timestamp 0
transform 1 0 4870 0 -1 3130
box -6 -8 86 248
use NAND2X1  _1708_
timestamp 0
transform -1 0 4750 0 1 3130
box -6 -8 86 248
use OAI21X1  _1709_
timestamp 0
transform 1 0 4730 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1710_
timestamp 0
transform 1 0 5230 0 -1 3610
box -6 -8 106 248
use AOI21X1  _1711_
timestamp 0
transform 1 0 5090 0 -1 3610
box -6 -8 106 248
use NOR2X1  _1712_
timestamp 0
transform -1 0 5390 0 1 1690
box -6 -8 86 248
use OAI21X1  _1713_
timestamp 0
transform -1 0 5370 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1714_
timestamp 0
transform 1 0 5310 0 1 3130
box -6 -8 106 248
use OR2X2  _1715_
timestamp 0
transform 1 0 5550 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1716_
timestamp 0
transform -1 0 5550 0 1 3130
box -6 -8 106 248
use NAND2X1  _1717_
timestamp 0
transform 1 0 5470 0 1 2650
box -6 -8 86 248
use INVX1  _1718_
timestamp 0
transform -1 0 4950 0 -1 2650
box -6 -8 66 248
use NOR2X1  _1719_
timestamp 0
transform -1 0 5270 0 1 3130
box -6 -8 86 248
use OAI21X1  _1720_
timestamp 0
transform -1 0 5510 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1721_
timestamp 0
transform -1 0 4550 0 1 2650
box -6 -8 86 248
use NAND3X1  _1722_
timestamp 0
transform -1 0 4510 0 -1 2650
box -6 -8 106 248
use AOI22X1  _1723_
timestamp 0
transform 1 0 4250 0 -1 2650
box -6 -8 126 248
use INVX1  _1724_
timestamp 0
transform 1 0 4090 0 -1 3130
box -6 -8 66 248
use NOR2X1  _1725_
timestamp 0
transform -1 0 4270 0 -1 3130
box -6 -8 86 248
use OAI21X1  _1726_
timestamp 0
transform 1 0 4310 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1727_
timestamp 0
transform 1 0 4330 0 1 2650
box -6 -8 106 248
use OAI21X1  _1728_
timestamp 0
transform 1 0 3490 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1729_
timestamp 0
transform -1 0 3550 0 1 2170
box -6 -8 106 248
use INVX1  _1730_
timestamp 0
transform -1 0 3650 0 1 2170
box -6 -8 66 248
use OAI21X1  _1731_
timestamp 0
transform 1 0 3690 0 1 2170
box -6 -8 106 248
use MUX2X1  _1732_
timestamp 0
transform -1 0 3950 0 -1 2650
box -6 -8 126 248
use NAND2X1  _1733_
timestamp 0
transform 1 0 3990 0 -1 2650
box -6 -8 86 248
use INVX1  _1734_
timestamp 0
transform -1 0 5150 0 1 3130
box -6 -8 66 248
use OAI21X1  _1735_
timestamp 0
transform -1 0 5050 0 1 3130
box -6 -8 106 248
use MUX2X1  _1736_
timestamp 0
transform 1 0 4870 0 1 2650
box -6 -8 126 248
use OAI21X1  _1737_
timestamp 0
transform 1 0 4590 0 1 2650
box -6 -8 106 248
use NAND2X1  _1738_
timestamp 0
transform 1 0 5030 0 1 2650
box -6 -8 86 248
use NAND3X1  _1739_
timestamp 0
transform 1 0 5130 0 -1 3130
box -6 -8 106 248
use NAND3X1  _1740_
timestamp 0
transform 1 0 4990 0 -1 3130
box -6 -8 106 248
use AOI22X1  _1741_
timestamp 0
transform 1 0 4790 0 1 3130
box -6 -8 126 248
use OAI21X1  _1742_
timestamp 0
transform -1 0 4190 0 1 2170
box -6 -8 106 248
use OAI21X1  _1743_
timestamp 0
transform 1 0 3950 0 1 2170
box -6 -8 106 248
use NAND2X1  _1744_
timestamp 0
transform -1 0 3910 0 1 2170
box -6 -8 86 248
use NAND2X1  _1745_
timestamp 0
transform 1 0 3890 0 -1 2170
box -6 -8 86 248
use INVX1  _1746_
timestamp 0
transform -1 0 3790 0 -1 1690
box -6 -8 66 248
use NOR2X1  _1747_
timestamp 0
transform 1 0 4230 0 1 2170
box -6 -8 86 248
use OAI21X1  _1748_
timestamp 0
transform -1 0 4250 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1749_
timestamp 0
transform -1 0 4750 0 -1 2650
box -6 -8 86 248
use INVX1  _1750_
timestamp 0
transform 1 0 3870 0 -1 3130
box -6 -8 66 248
use NOR2X1  _1751_
timestamp 0
transform -1 0 4050 0 -1 3130
box -6 -8 86 248
use NAND2X1  _1752_
timestamp 0
transform -1 0 3990 0 1 2650
box -6 -8 86 248
use AOI22X1  _1753_
timestamp 0
transform -1 0 4290 0 1 2650
box -6 -8 126 248
use OAI21X1  _1754_
timestamp 0
transform 1 0 4030 0 1 2650
box -6 -8 106 248
use OAI21X1  _1755_
timestamp 0
transform 1 0 4110 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1756_
timestamp 0
transform -1 0 3690 0 1 1690
box -6 -8 106 248
use AOI21X1  _1757_
timestamp 0
transform 1 0 3890 0 1 1690
box -6 -8 106 248
use INVX1  _1758_
timestamp 0
transform 1 0 4310 0 1 1690
box -6 -8 66 248
use OAI21X1  _1759_
timestamp 0
transform -1 0 4770 0 -1 1690
box -6 -8 106 248
use MUX2X1  _1760_
timestamp 0
transform 1 0 4510 0 -1 1690
box -6 -8 126 248
use NAND2X1  _1761_
timestamp 0
transform -1 0 4470 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1762_
timestamp 0
transform -1 0 4270 0 1 1690
box -6 -8 106 248
use OAI21X1  _1763_
timestamp 0
transform -1 0 4130 0 1 1690
box -6 -8 106 248
use NAND3X1  _1764_
timestamp 0
transform -1 0 4110 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1765_
timestamp 0
transform 1 0 4270 0 -1 1690
box -6 -8 86 248
use INVX1  _1766_
timestamp 0
transform 1 0 4170 0 -1 1690
box -6 -8 66 248
use INVX1  _1767_
timestamp 0
transform 1 0 4450 0 -1 1210
box -6 -8 66 248
use AND2X2  _1768_
timestamp 0
transform -1 0 4190 0 1 1210
box -6 -8 106 248
use NAND2X1  _1769_
timestamp 0
transform 1 0 4710 0 -1 2170
box -6 -8 86 248
use AND2X2  _1770_
timestamp 0
transform -1 0 4530 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1771_
timestamp 0
transform -1 0 4430 0 1 2170
box -6 -8 86 248
use AOI22X1  _1772_
timestamp 0
transform -1 0 4590 0 1 2170
box -6 -8 126 248
use OAI21X1  _1773_
timestamp 0
transform -1 0 4390 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1774_
timestamp 0
transform 1 0 4570 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1775_
timestamp 0
transform -1 0 4610 0 1 1690
box -6 -8 106 248
use AOI21X1  _1776_
timestamp 0
transform 1 0 4650 0 1 1690
box -6 -8 106 248
use OAI21X1  _1777_
timestamp 0
transform 1 0 4950 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1778_
timestamp 0
transform 1 0 4810 0 -1 1690
box -6 -8 106 248
use INVX1  _1779_
timestamp 0
transform 1 0 4790 0 -1 1210
box -6 -8 66 248
use OAI21X1  _1780_
timestamp 0
transform 1 0 4550 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1781_
timestamp 0
transform -1 0 4330 0 1 1210
box -6 -8 106 248
use NAND2X1  _1782_
timestamp 0
transform 1 0 4330 0 -1 1210
box -6 -8 86 248
use INVX1  _1783_
timestamp 0
transform -1 0 2870 0 -1 250
box -6 -8 66 248
use INVX1  _1784_
timestamp 0
transform -1 0 3650 0 1 1210
box -6 -8 66 248
use AOI21X1  _1785_
timestamp 0
transform -1 0 3790 0 1 1210
box -6 -8 106 248
use NAND3X1  _1786_
timestamp 0
transform -1 0 4290 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1787_
timestamp 0
transform 1 0 4370 0 1 1210
box -6 -8 86 248
use INVX1  _1788_
timestamp 0
transform 1 0 5030 0 -1 1210
box -6 -8 66 248
use AOI21X1  _1789_
timestamp 0
transform 1 0 4890 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1790_
timestamp 0
transform 1 0 5130 0 -1 2650
box -6 -8 86 248
use AND2X2  _1791_
timestamp 0
transform 1 0 5590 0 1 2650
box -6 -8 106 248
use NAND2X1  _1792_
timestamp 0
transform 1 0 5550 0 -1 2650
box -6 -8 86 248
use AOI22X1  _1793_
timestamp 0
transform 1 0 5390 0 -1 2650
box -6 -8 126 248
use OAI21X1  _1794_
timestamp 0
transform 1 0 5390 0 -1 250
box -6 -8 106 248
use OAI21X1  _1795_
timestamp 0
transform -1 0 5350 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1796_
timestamp 0
transform 1 0 5510 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1797_
timestamp 0
transform -1 0 5470 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1798_
timestamp 0
transform 1 0 4610 0 1 1210
box -6 -8 106 248
use OAI21X1  _1799_
timestamp 0
transform 1 0 4750 0 1 1210
box -6 -8 106 248
use AOI21X1  _1800_
timestamp 0
transform 1 0 4210 0 1 730
box -6 -8 106 248
use NOR2X1  _1801_
timestamp 0
transform -1 0 4050 0 1 1210
box -6 -8 86 248
use OAI21X1  _1802_
timestamp 0
transform -1 0 3930 0 1 1210
box -6 -8 106 248
use NAND2X1  _1803_
timestamp 0
transform 1 0 3710 0 1 730
box -6 -8 86 248
use OAI21X1  _1804_
timestamp 0
transform 1 0 3830 0 1 730
box -6 -8 106 248
use INVX1  _1805_
timestamp 0
transform -1 0 4410 0 1 730
box -6 -8 66 248
use NOR2X1  _1806_
timestamp 0
transform 1 0 4390 0 -1 730
box -6 -8 86 248
use NOR2X1  _1807_
timestamp 0
transform 1 0 4270 0 -1 730
box -6 -8 86 248
use INVX1  _1808_
timestamp 0
transform -1 0 4750 0 -1 1210
box -6 -8 66 248
use NAND2X1  _1809_
timestamp 0
transform -1 0 4910 0 -1 2170
box -6 -8 86 248
use AND2X2  _1810_
timestamp 0
transform -1 0 5010 0 1 2170
box -6 -8 106 248
use NAND2X1  _1811_
timestamp 0
transform -1 0 4870 0 1 2170
box -6 -8 86 248
use AOI22X1  _1812_
timestamp 0
transform 1 0 4630 0 1 2170
box -6 -8 126 248
use OAI21X1  _1813_
timestamp 0
transform 1 0 5090 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1814_
timestamp 0
transform -1 0 5050 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1815_
timestamp 0
transform 1 0 4910 0 1 1690
box -6 -8 106 248
use AOI21X1  _1816_
timestamp 0
transform 1 0 5050 0 1 1690
box -6 -8 106 248
use OAI21X1  _1817_
timestamp 0
transform 1 0 5270 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1818_
timestamp 0
transform 1 0 5130 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1819_
timestamp 0
transform -1 0 4550 0 1 730
box -6 -8 106 248
use AOI21X1  _1820_
timestamp 0
transform 1 0 4510 0 -1 730
box -6 -8 106 248
use INVX1  _1821_
timestamp 0
transform -1 0 4970 0 -1 730
box -6 -8 66 248
use NAND2X1  _1822_
timestamp 0
transform 1 0 4790 0 -1 730
box -6 -8 86 248
use NAND2X1  _1823_
timestamp 0
transform -1 0 4170 0 1 730
box -6 -8 86 248
use OAI21X1  _1824_
timestamp 0
transform 1 0 5010 0 -1 730
box -6 -8 106 248
use INVX1  _1825_
timestamp 0
transform 1 0 4890 0 1 1210
box -6 -8 66 248
use AND2X2  _1826_
timestamp 0
transform -1 0 5470 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1827_
timestamp 0
transform -1 0 5290 0 1 730
box -6 -8 86 248
use AOI22X1  _1828_
timestamp 0
transform 1 0 5050 0 1 2170
box -6 -8 126 248
use OAI21X1  _1829_
timestamp 0
transform 1 0 5230 0 -1 2170
box -6 -8 106 248
use OAI22X1  _1830_
timestamp 0
transform 1 0 4990 0 1 1210
box -6 -8 126 248
use OAI21X1  _1831_
timestamp 0
transform 1 0 5090 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1832_
timestamp 0
transform 1 0 5230 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1833_
timestamp 0
transform 1 0 5530 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1834_
timestamp 0
transform 1 0 5570 0 1 4090
box -6 -8 106 248
use NAND2X1  _1835_
timestamp 0
transform -1 0 4650 0 1 250
box -6 -8 86 248
use OAI21X1  _1836_
timestamp 0
transform 1 0 4650 0 -1 730
box -6 -8 106 248
use INVX1  _1837_
timestamp 0
transform -1 0 5710 0 -1 730
box -6 -8 66 248
use NAND3X1  _1838_
timestamp 0
transform -1 0 4790 0 1 250
box -6 -8 106 248
use NAND2X1  _1839_
timestamp 0
transform 1 0 4330 0 1 250
box -6 -8 86 248
use INVX1  _1840_
timestamp 0
transform -1 0 5710 0 1 250
box -6 -8 66 248
use AOI21X1  _1841_
timestamp 0
transform 1 0 4830 0 1 250
box -6 -8 106 248
use NAND2X1  _1842_
timestamp 0
transform 1 0 5610 0 -1 3610
box -6 -8 86 248
use AND2X2  _1843_
timestamp 0
transform 1 0 5510 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1844_
timestamp 0
transform 1 0 4890 0 -1 250
box -6 -8 86 248
use AOI22X1  _1845_
timestamp 0
transform 1 0 5210 0 1 2170
box -6 -8 126 248
use OAI21X1  _1846_
timestamp 0
transform 1 0 5510 0 1 2170
box -6 -8 106 248
use OAI21X1  _1847_
timestamp 0
transform -1 0 5470 0 1 2170
box -6 -8 106 248
use OAI21X1  _1848_
timestamp 0
transform -1 0 5650 0 1 1690
box -6 -8 106 248
use AOI21X1  _1849_
timestamp 0
transform 1 0 5250 0 -1 250
box -6 -8 106 248
use OAI21X1  _1850_
timestamp 0
transform 1 0 5610 0 1 730
box -6 -8 106 248
use OAI21X1  _1851_
timestamp 0
transform -1 0 5570 0 1 730
box -6 -8 106 248
use OAI21X1  _1852_
timestamp 0
transform -1 0 5470 0 1 250
box -6 -8 106 248
use NAND2X1  _1853_
timestamp 0
transform -1 0 5050 0 1 250
box -6 -8 86 248
use INVX1  _1854_
timestamp 0
transform 1 0 5430 0 -1 730
box -6 -8 66 248
use NAND3X1  _1855_
timestamp 0
transform -1 0 5190 0 1 250
box -6 -8 106 248
use NAND2X1  _1856_
timestamp 0
transform -1 0 4530 0 1 250
box -6 -8 86 248
use NOR2X1  _1857_
timestamp 0
transform -1 0 4010 0 -1 1210
box -6 -8 86 248
use NAND2X1  _1858_
timestamp 0
transform -1 0 4050 0 1 730
box -6 -8 86 248
use NOR2X1  _1859_
timestamp 0
transform 1 0 4030 0 -1 730
box -6 -8 86 248
use INVX1  _1860_
timestamp 0
transform 1 0 4090 0 1 250
box -6 -8 66 248
use NAND3X1  _1861_
timestamp 0
transform -1 0 4290 0 1 250
box -6 -8 106 248
use NOR2X1  _1862_
timestamp 0
transform -1 0 4230 0 -1 730
box -6 -8 86 248
use AND2X2  _1863_
timestamp 0
transform -1 0 3990 0 -1 730
box -6 -8 106 248
use NAND3X1  _1864_
timestamp 0
transform -1 0 5330 0 1 250
box -6 -8 106 248
use OAI21X1  _1865_
timestamp 0
transform -1 0 5610 0 1 250
box -6 -8 106 248
use NAND2X1  _1866_
timestamp 0
transform 1 0 4390 0 -1 250
box -6 -8 86 248
use OAI21X1  _1867_
timestamp 0
transform -1 0 4050 0 1 250
box -6 -8 106 248
use NOR2X1  _1868_
timestamp 0
transform 1 0 4490 0 1 1210
box -6 -8 86 248
use OAI21X1  _1869_
timestamp 0
transform -1 0 5430 0 1 730
box -6 -8 106 248
use INVX1  _1870_
timestamp 0
transform -1 0 4930 0 1 730
box -6 -8 66 248
use NAND3X1  _1871_
timestamp 0
transform -1 0 5250 0 -1 730
box -6 -8 106 248
use NAND3X1  _1872_
timestamp 0
transform -1 0 4830 0 1 730
box -6 -8 106 248
use INVX1  _1873_
timestamp 0
transform -1 0 5030 0 1 730
box -6 -8 66 248
use NAND2X1  _1874_
timestamp 0
transform 1 0 5530 0 -1 730
box -6 -8 86 248
use AOI21X1  _1875_
timestamp 0
transform 1 0 5290 0 -1 730
box -6 -8 106 248
use OAI21X1  _1876_
timestamp 0
transform -1 0 5170 0 1 730
box -6 -8 106 248
use AND2X2  _1877_
timestamp 0
transform -1 0 4690 0 1 730
box -6 -8 106 248
use OAI21X1  _1878_
timestamp 0
transform -1 0 3970 0 -1 250
box -6 -8 106 248
use NAND3X1  _1879_
timestamp 0
transform -1 0 3910 0 1 250
box -6 -8 106 248
use INVX1  _1880_
timestamp 0
transform -1 0 5710 0 1 1210
box -6 -8 66 248
use NAND2X1  _1881_
timestamp 0
transform 1 0 5530 0 1 1210
box -6 -8 86 248
use AOI21X1  _1882_
timestamp 0
transform -1 0 5490 0 1 1210
box -6 -8 106 248
use NAND2X1  _1883_
timestamp 0
transform -1 0 5350 0 1 1210
box -6 -8 86 248
use NOR2X1  _1884_
timestamp 0
transform -1 0 5230 0 1 1210
box -6 -8 86 248
use NOR2X1  _1885_
timestamp 0
transform 1 0 5410 0 -1 1210
box -6 -8 86 248
use NAND3X1  _1886_
timestamp 0
transform -1 0 4850 0 -1 250
box -6 -8 106 248
use INVX1  _1887_
timestamp 0
transform -1 0 4710 0 -1 250
box -6 -8 66 248
use NAND3X1  _1888_
timestamp 0
transform -1 0 4610 0 -1 250
box -6 -8 106 248
use NAND2X1  _1889_
timestamp 0
transform 1 0 4270 0 -1 250
box -6 -8 86 248
use NAND3X1  _1890_
timestamp 0
transform -1 0 3830 0 -1 250
box -6 -8 106 248
use AND2X2  _1891_
timestamp 0
transform -1 0 4230 0 -1 250
box -6 -8 106 248
use NAND2X1  _1892_
timestamp 0
transform -1 0 3690 0 -1 250
box -6 -8 86 248
use NAND2X1  _1893_
timestamp 0
transform -1 0 3570 0 -1 250
box -6 -8 86 248
use BUFX2  _1894_
timestamp 0
transform -1 0 2750 0 1 2650
box -6 -8 86 248
use BUFX2  _1895_
timestamp 0
transform -1 0 2730 0 -1 2650
box -6 -8 86 248
use BUFX2  _1896_
timestamp 0
transform -1 0 130 0 1 3610
box -6 -8 86 248
use BUFX2  _1897_
timestamp 0
transform 1 0 2690 0 -1 250
box -6 -8 86 248
use BUFX2  _1898_
timestamp 0
transform -1 0 3230 0 -1 250
box -6 -8 86 248
use BUFX2  _1899_
timestamp 0
transform 1 0 3570 0 1 250
box -6 -8 86 248
use BUFX2  _1900_
timestamp 0
transform -1 0 3350 0 -1 250
box -6 -8 86 248
use BUFX2  _1901_
timestamp 0
transform -1 0 3770 0 1 250
box -6 -8 86 248
use BUFX2  _1902_
timestamp 0
transform -1 0 4090 0 -1 250
box -6 -8 86 248
use BUFX2  BUFX2_insert0
timestamp 0
transform -1 0 2470 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert1
timestamp 0
transform -1 0 2590 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert2
timestamp 0
transform 1 0 4090 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert3
timestamp 0
transform 1 0 4550 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert4
timestamp 0
transform -1 0 3870 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert5
timestamp 0
transform 1 0 1770 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert6
timestamp 0
transform -1 0 1710 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert7
timestamp 0
transform 1 0 3750 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert8
timestamp 0
transform -1 0 4790 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert9
timestamp 0
transform 1 0 5070 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert10
timestamp 0
transform -1 0 5310 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert11
timestamp 0
transform 1 0 5530 0 -1 250
box -6 -8 86 248
use BUFX2  BUFX2_insert17
timestamp 0
transform -1 0 3990 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert18
timestamp 0
transform 1 0 4030 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert19
timestamp 0
transform 1 0 5150 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert20
timestamp 0
transform 1 0 5350 0 -1 5050
box -6 -8 86 248
use BUFX2  BUFX2_insert21
timestamp 0
transform 1 0 2390 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert22
timestamp 0
transform 1 0 5590 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert23
timestamp 0
transform -1 0 2350 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert24
timestamp 0
transform 1 0 3030 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert25
timestamp 0
transform 1 0 2710 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert26
timestamp 0
transform 1 0 1650 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert27
timestamp 0
transform -1 0 3590 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert28
timestamp 0
transform -1 0 1590 0 1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert29
timestamp 0
transform -1 0 5510 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert30
timestamp 0
transform 1 0 5190 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert31
timestamp 0
transform 1 0 4790 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert32
timestamp 0
transform 1 0 5010 0 -1 2650
box -6 -8 86 248
use CLKBUF1  CLKBUF1_insert12
timestamp 0
transform 1 0 4090 0 -1 4090
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert13
timestamp 0
transform -1 0 4290 0 -1 3610
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert14
timestamp 0
transform 1 0 3530 0 1 5530
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert15
timestamp 0
transform -1 0 4050 0 -1 3610
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert16
timestamp 0
transform 1 0 4410 0 -1 4570
box -6 -8 206 248
use FILL  FILL84150x21750
timestamp 0
transform -1 0 5630 0 -1 1690
box -6 -8 26 248
use FILL  FILL84150x28950
timestamp 0
transform -1 0 5630 0 -1 2170
box -6 -8 26 248
use FILL  FILL84150x32550
timestamp 0
transform 1 0 5610 0 1 2170
box -6 -8 26 248
use FILL  FILL84150x64950
timestamp 0
transform -1 0 5630 0 -1 4570
box -6 -8 26 248
use FILL  FILL84150x82950
timestamp 0
transform 1 0 5610 0 1 5530
box -6 -8 26 248
use FILL  FILL84450x14550
timestamp 0
transform -1 0 5650 0 -1 1210
box -6 -8 26 248
use FILL  FILL84450x21750
timestamp 0
transform -1 0 5650 0 -1 1690
box -6 -8 26 248
use FILL  FILL84450x28950
timestamp 0
transform -1 0 5650 0 -1 2170
box -6 -8 26 248
use FILL  FILL84450x32550
timestamp 0
transform 1 0 5630 0 1 2170
box -6 -8 26 248
use FILL  FILL84450x36150
timestamp 0
transform -1 0 5650 0 -1 2650
box -6 -8 26 248
use FILL  FILL84450x54150
timestamp 0
transform 1 0 5630 0 1 3610
box -6 -8 26 248
use FILL  FILL84450x64950
timestamp 0
transform -1 0 5650 0 -1 4570
box -6 -8 26 248
use FILL  FILL84450x82950
timestamp 0
transform 1 0 5630 0 1 5530
box -6 -8 26 248
use FILL  FILL84750x14550
timestamp 0
transform -1 0 5670 0 -1 1210
box -6 -8 26 248
use FILL  FILL84750x21750
timestamp 0
transform -1 0 5670 0 -1 1690
box -6 -8 26 248
use FILL  FILL84750x25350
timestamp 0
transform 1 0 5650 0 1 1690
box -6 -8 26 248
use FILL  FILL84750x28950
timestamp 0
transform -1 0 5670 0 -1 2170
box -6 -8 26 248
use FILL  FILL84750x32550
timestamp 0
transform 1 0 5650 0 1 2170
box -6 -8 26 248
use FILL  FILL84750x36150
timestamp 0
transform -1 0 5670 0 -1 2650
box -6 -8 26 248
use FILL  FILL84750x43350
timestamp 0
transform -1 0 5670 0 -1 3130
box -6 -8 26 248
use FILL  FILL84750x54150
timestamp 0
transform 1 0 5650 0 1 3610
box -6 -8 26 248
use FILL  FILL84750x64950
timestamp 0
transform -1 0 5670 0 -1 4570
box -6 -8 26 248
use FILL  FILL84750x68550
timestamp 0
transform 1 0 5650 0 1 4570
box -6 -8 26 248
use FILL  FILL84750x75750
timestamp 0
transform 1 0 5650 0 1 5050
box -6 -8 26 248
use FILL  FILL84750x79350
timestamp 0
transform -1 0 5670 0 -1 5530
box -6 -8 26 248
use FILL  FILL84750x82950
timestamp 0
transform 1 0 5650 0 1 5530
box -6 -8 26 248
use FILL  FILL85050x14550
timestamp 0
transform -1 0 5690 0 -1 1210
box -6 -8 26 248
use FILL  FILL85050x21750
timestamp 0
transform -1 0 5690 0 -1 1690
box -6 -8 26 248
use FILL  FILL85050x25350
timestamp 0
transform 1 0 5670 0 1 1690
box -6 -8 26 248
use FILL  FILL85050x28950
timestamp 0
transform -1 0 5690 0 -1 2170
box -6 -8 26 248
use FILL  FILL85050x32550
timestamp 0
transform 1 0 5670 0 1 2170
box -6 -8 26 248
use FILL  FILL85050x36150
timestamp 0
transform -1 0 5690 0 -1 2650
box -6 -8 26 248
use FILL  FILL85050x43350
timestamp 0
transform -1 0 5690 0 -1 3130
box -6 -8 26 248
use FILL  FILL85050x46950
timestamp 0
transform 1 0 5670 0 1 3130
box -6 -8 26 248
use FILL  FILL85050x54150
timestamp 0
transform 1 0 5670 0 1 3610
box -6 -8 26 248
use FILL  FILL85050x57750
timestamp 0
transform -1 0 5690 0 -1 4090
box -6 -8 26 248
use FILL  FILL85050x61350
timestamp 0
transform 1 0 5670 0 1 4090
box -6 -8 26 248
use FILL  FILL85050x64950
timestamp 0
transform -1 0 5690 0 -1 4570
box -6 -8 26 248
use FILL  FILL85050x68550
timestamp 0
transform 1 0 5670 0 1 4570
box -6 -8 26 248
use FILL  FILL85050x75750
timestamp 0
transform 1 0 5670 0 1 5050
box -6 -8 26 248
use FILL  FILL85050x79350
timestamp 0
transform -1 0 5690 0 -1 5530
box -6 -8 26 248
use FILL  FILL85050x82950
timestamp 0
transform 1 0 5670 0 1 5530
box -6 -8 26 248
use FILL  FILL85350x14550
timestamp 0
transform -1 0 5710 0 -1 1210
box -6 -8 26 248
use FILL  FILL85350x21750
timestamp 0
transform -1 0 5710 0 -1 1690
box -6 -8 26 248
use FILL  FILL85350x25350
timestamp 0
transform 1 0 5690 0 1 1690
box -6 -8 26 248
use FILL  FILL85350x28950
timestamp 0
transform -1 0 5710 0 -1 2170
box -6 -8 26 248
use FILL  FILL85350x32550
timestamp 0
transform 1 0 5690 0 1 2170
box -6 -8 26 248
use FILL  FILL85350x36150
timestamp 0
transform -1 0 5710 0 -1 2650
box -6 -8 26 248
use FILL  FILL85350x39750
timestamp 0
transform 1 0 5690 0 1 2650
box -6 -8 26 248
use FILL  FILL85350x43350
timestamp 0
transform -1 0 5710 0 -1 3130
box -6 -8 26 248
use FILL  FILL85350x46950
timestamp 0
transform 1 0 5690 0 1 3130
box -6 -8 26 248
use FILL  FILL85350x50550
timestamp 0
transform -1 0 5710 0 -1 3610
box -6 -8 26 248
use FILL  FILL85350x54150
timestamp 0
transform 1 0 5690 0 1 3610
box -6 -8 26 248
use FILL  FILL85350x57750
timestamp 0
transform -1 0 5710 0 -1 4090
box -6 -8 26 248
use FILL  FILL85350x61350
timestamp 0
transform 1 0 5690 0 1 4090
box -6 -8 26 248
use FILL  FILL85350x64950
timestamp 0
transform -1 0 5710 0 -1 4570
box -6 -8 26 248
use FILL  FILL85350x68550
timestamp 0
transform 1 0 5690 0 1 4570
box -6 -8 26 248
use FILL  FILL85350x72150
timestamp 0
transform -1 0 5710 0 -1 5050
box -6 -8 26 248
use FILL  FILL85350x75750
timestamp 0
transform 1 0 5690 0 1 5050
box -6 -8 26 248
use FILL  FILL85350x79350
timestamp 0
transform -1 0 5710 0 -1 5530
box -6 -8 26 248
use FILL  FILL85350x82950
timestamp 0
transform 1 0 5690 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__927_
timestamp 0
transform -1 0 4270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__928_
timestamp 0
transform 1 0 3790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__929_
timestamp 0
transform -1 0 3850 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__930_
timestamp 0
transform 1 0 3950 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__931_
timestamp 0
transform 1 0 4150 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__932_
timestamp 0
transform -1 0 2850 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__933_
timestamp 0
transform 1 0 4350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__934_
timestamp 0
transform -1 0 4610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__935_
timestamp 0
transform 1 0 5530 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__936_
timestamp 0
transform 1 0 4470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__937_
timestamp 0
transform 1 0 4790 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__938_
timestamp 0
transform -1 0 4970 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__939_
timestamp 0
transform -1 0 4830 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__940_
timestamp 0
transform -1 0 4070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__941_
timestamp 0
transform -1 0 3610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__942_
timestamp 0
transform -1 0 4030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__943_
timestamp 0
transform -1 0 4310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__944_
timestamp 0
transform -1 0 3650 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__945_
timestamp 0
transform -1 0 3970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__946_
timestamp 0
transform 1 0 5070 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__947_
timestamp 0
transform 1 0 4930 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__948_
timestamp 0
transform 1 0 4650 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__949_
timestamp 0
transform 1 0 4490 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__950_
timestamp 0
transform -1 0 4230 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__951_
timestamp 0
transform 1 0 4390 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__952_
timestamp 0
transform 1 0 4530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__953_
timestamp 0
transform 1 0 4470 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__954_
timestamp 0
transform 1 0 4950 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__955_
timestamp 0
transform 1 0 5070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__956_
timestamp 0
transform 1 0 5330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__957_
timestamp 0
transform 1 0 5190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__958_
timestamp 0
transform 1 0 5550 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__959_
timestamp 0
transform -1 0 5510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__960_
timestamp 0
transform 1 0 4150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__961_
timestamp 0
transform -1 0 4830 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__962_
timestamp 0
transform 1 0 4670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__963_
timestamp 0
transform -1 0 5190 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__964_
timestamp 0
transform 1 0 4310 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__965_
timestamp 0
transform 1 0 4430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__966_
timestamp 0
transform 1 0 4290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__967_
timestamp 0
transform -1 0 4430 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__968_
timestamp 0
transform -1 0 4070 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__969_
timestamp 0
transform -1 0 4190 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__970_
timestamp 0
transform 1 0 5190 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__971_
timestamp 0
transform -1 0 4310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__972_
timestamp 0
transform -1 0 4430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__973_
timestamp 0
transform -1 0 5350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__974_
timestamp 0
transform 1 0 4170 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__975_
timestamp 0
transform -1 0 4310 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__976_
timestamp 0
transform -1 0 5330 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__977_
timestamp 0
transform -1 0 5430 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__978_
timestamp 0
transform 1 0 5470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__979_
timestamp 0
transform -1 0 5230 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__980_
timestamp 0
transform 1 0 4950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__981_
timestamp 0
transform -1 0 5090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__982_
timestamp 0
transform 1 0 4590 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__983_
timestamp 0
transform -1 0 4130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__984_
timestamp 0
transform -1 0 4250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__985_
timestamp 0
transform -1 0 3190 0 1 730
box -6 -8 26 248
use FILL  FILL_0__986_
timestamp 0
transform 1 0 5290 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__987_
timestamp 0
transform 1 0 5150 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__988_
timestamp 0
transform -1 0 3050 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__989_
timestamp 0
transform -1 0 2690 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__990_
timestamp 0
transform 1 0 2450 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__991_
timestamp 0
transform 1 0 2430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__992_
timestamp 0
transform 1 0 2570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__993_
timestamp 0
transform 1 0 2110 0 1 250
box -6 -8 26 248
use FILL  FILL_0__994_
timestamp 0
transform -1 0 2330 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__995_
timestamp 0
transform -1 0 1510 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__996_
timestamp 0
transform 1 0 1830 0 1 730
box -6 -8 26 248
use FILL  FILL_0__997_
timestamp 0
transform -1 0 2790 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__998_
timestamp 0
transform 1 0 2250 0 1 730
box -6 -8 26 248
use FILL  FILL_0__999_
timestamp 0
transform -1 0 2570 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1000_
timestamp 0
transform 1 0 1370 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1001_
timestamp 0
transform -1 0 1370 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1002_
timestamp 0
transform 1 0 2930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1003_
timestamp 0
transform -1 0 1470 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1004_
timestamp 0
transform -1 0 1750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1005_
timestamp 0
transform 1 0 1790 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1006_
timestamp 0
transform -1 0 1390 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1007_
timestamp 0
transform 1 0 1590 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1008_
timestamp 0
transform -1 0 1250 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1009_
timestamp 0
transform -1 0 890 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1010_
timestamp 0
transform 1 0 2450 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1011_
timestamp 0
transform 1 0 2550 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1012_
timestamp 0
transform 1 0 1970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1013_
timestamp 0
transform 1 0 2550 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1014_
timestamp 0
transform 1 0 2290 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1015_
timestamp 0
transform -1 0 2330 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1016_
timestamp 0
transform 1 0 1010 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1017_
timestamp 0
transform -1 0 750 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1018_
timestamp 0
transform -1 0 1230 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1019_
timestamp 0
transform -1 0 1330 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1020_
timestamp 0
transform -1 0 970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1021_
timestamp 0
transform -1 0 1470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1022_
timestamp 0
transform -1 0 30 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1023_
timestamp 0
transform -1 0 1270 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1024_
timestamp 0
transform -1 0 30 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1025_
timestamp 0
transform 1 0 390 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1026_
timestamp 0
transform -1 0 1630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1027_
timestamp 0
transform -1 0 1110 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1028_
timestamp 0
transform -1 0 550 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1029_
timestamp 0
transform 1 0 670 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1030_
timestamp 0
transform -1 0 1530 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1031_
timestamp 0
transform -1 0 130 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1032_
timestamp 0
transform 1 0 250 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1033_
timestamp 0
transform -1 0 270 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1034_
timestamp 0
transform 1 0 2810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1035_
timestamp 0
transform 1 0 2710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1036_
timestamp 0
transform -1 0 2210 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1037_
timestamp 0
transform -1 0 2190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1038_
timestamp 0
transform 1 0 2490 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1039_
timestamp 0
transform 1 0 2430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1040_
timestamp 0
transform -1 0 2310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1041_
timestamp 0
transform 1 0 2030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1042_
timestamp 0
transform -1 0 1450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1043_
timestamp 0
transform -1 0 1810 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1044_
timestamp 0
transform -1 0 1910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1045_
timestamp 0
transform -1 0 1530 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1046_
timestamp 0
transform -1 0 690 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1047_
timestamp 0
transform 1 0 390 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1048_
timestamp 0
transform 1 0 810 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1049_
timestamp 0
transform 1 0 1650 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1050_
timestamp 0
transform 1 0 1090 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1051_
timestamp 0
transform -1 0 30 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1052_
timestamp 0
transform 1 0 150 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1053_
timestamp 0
transform 1 0 290 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1054_
timestamp 0
transform -1 0 550 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1055_
timestamp 0
transform 1 0 850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1056_
timestamp 0
transform -1 0 1530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1057_
timestamp 0
transform 1 0 1070 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1058_
timestamp 0
transform -1 0 1390 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1059_
timestamp 0
transform -1 0 2450 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1060_
timestamp 0
transform 1 0 1310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1061_
timestamp 0
transform -1 0 1250 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1062_
timestamp 0
transform -1 0 970 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1063_
timestamp 0
transform -1 0 750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1064_
timestamp 0
transform 1 0 710 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1065_
timestamp 0
transform -1 0 1410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1066_
timestamp 0
transform 1 0 1090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1067_
timestamp 0
transform 1 0 1450 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1068_
timestamp 0
transform 1 0 850 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1069_
timestamp 0
transform -1 0 730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1070_
timestamp 0
transform 1 0 110 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1071_
timestamp 0
transform -1 0 590 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1072_
timestamp 0
transform -1 0 450 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1073_
timestamp 0
transform -1 0 310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1074_
timestamp 0
transform -1 0 1870 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1075_
timestamp 0
transform -1 0 1850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1076_
timestamp 0
transform -1 0 2230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1077_
timestamp 0
transform -1 0 2250 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1078_
timestamp 0
transform 1 0 2110 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1079_
timestamp 0
transform 1 0 1670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1080_
timestamp 0
transform -1 0 2090 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1081_
timestamp 0
transform 1 0 1930 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1082_
timestamp 0
transform -1 0 1550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1083_
timestamp 0
transform 1 0 2070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1084_
timestamp 0
transform -1 0 1990 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1085_
timestamp 0
transform -1 0 1950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1086_
timestamp 0
transform -1 0 590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1087_
timestamp 0
transform -1 0 30 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1088_
timestamp 0
transform 1 0 430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1089_
timestamp 0
transform -1 0 590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1090_
timestamp 0
transform 1 0 710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1091_
timestamp 0
transform 1 0 150 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1092_
timestamp 0
transform -1 0 170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1093_
timestamp 0
transform -1 0 970 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1094_
timestamp 0
transform 1 0 290 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1095_
timestamp 0
transform -1 0 30 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1096_
timestamp 0
transform 1 0 570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1097_
timestamp 0
transform -1 0 3670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1098_
timestamp 0
transform -1 0 2190 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1099_
timestamp 0
transform -1 0 2050 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1100_
timestamp 0
transform 1 0 1910 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1101_
timestamp 0
transform -1 0 1790 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1102_
timestamp 0
transform -1 0 1010 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1103_
timestamp 0
transform 1 0 850 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1104_
timestamp 0
transform 1 0 430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1105_
timestamp 0
transform 1 0 290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1106_
timestamp 0
transform 1 0 1130 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1107_
timestamp 0
transform 1 0 710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1108_
timestamp 0
transform 1 0 1150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1109_
timestamp 0
transform -1 0 1430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1110_
timestamp 0
transform -1 0 730 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1111_
timestamp 0
transform -1 0 170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1112_
timestamp 0
transform -1 0 450 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1113_
timestamp 0
transform -1 0 1190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1114_
timestamp 0
transform 1 0 1430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1115_
timestamp 0
transform 1 0 690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1116_
timestamp 0
transform 1 0 1190 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1117_
timestamp 0
transform -1 0 590 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1118_
timestamp 0
transform -1 0 290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1119_
timestamp 0
transform 1 0 1050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1120_
timestamp 0
transform -1 0 950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1121_
timestamp 0
transform 1 0 810 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1122_
timestamp 0
transform -1 0 310 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1123_
timestamp 0
transform -1 0 690 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1124_
timestamp 0
transform -1 0 570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1125_
timestamp 0
transform -1 0 450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1126_
timestamp 0
transform 1 0 2290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1127_
timestamp 0
transform -1 0 1750 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1128_
timestamp 0
transform 1 0 1830 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1129_
timestamp 0
transform 1 0 2130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1130_
timestamp 0
transform 1 0 1970 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1131_
timestamp 0
transform -1 0 2090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1132_
timestamp 0
transform 1 0 2190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1133_
timestamp 0
transform -1 0 1610 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1134_
timestamp 0
transform 1 0 2850 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1135_
timestamp 0
transform 1 0 1850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1136_
timestamp 0
transform -1 0 2010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1137_
timestamp 0
transform -1 0 1730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1138_
timestamp 0
transform -1 0 30 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1139_
timestamp 0
transform -1 0 170 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1140_
timestamp 0
transform -1 0 610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1141_
timestamp 0
transform -1 0 310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1142_
timestamp 0
transform -1 0 170 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1143_
timestamp 0
transform 1 0 150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1144_
timestamp 0
transform -1 0 30 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1145_
timestamp 0
transform 1 0 150 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1146_
timestamp 0
transform -1 0 30 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1147_
timestamp 0
transform -1 0 30 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1148_
timestamp 0
transform 1 0 290 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1149_
timestamp 0
transform 1 0 150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1150_
timestamp 0
transform -1 0 2350 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1151_
timestamp 0
transform -1 0 1370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1152_
timestamp 0
transform -1 0 1690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1153_
timestamp 0
transform -1 0 1350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1154_
timestamp 0
transform -1 0 1410 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1155_
timestamp 0
transform 1 0 1530 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1156_
timestamp 0
transform 1 0 1270 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1157_
timestamp 0
transform -1 0 1090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1158_
timestamp 0
transform -1 0 1230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1159_
timestamp 0
transform -1 0 1670 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1160_
timestamp 0
transform -1 0 1150 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1161_
timestamp 0
transform -1 0 970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1162_
timestamp 0
transform 1 0 710 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1163_
timestamp 0
transform -1 0 30 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1164_
timestamp 0
transform -1 0 30 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1165_
timestamp 0
transform -1 0 1010 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1166_
timestamp 0
transform -1 0 1230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1167_
timestamp 0
transform 1 0 830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1168_
timestamp 0
transform 1 0 430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1169_
timestamp 0
transform 1 0 990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1170_
timestamp 0
transform -1 0 450 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1171_
timestamp 0
transform 1 0 290 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1172_
timestamp 0
transform 1 0 570 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1173_
timestamp 0
transform 1 0 990 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1174_
timestamp 0
transform 1 0 1410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1175_
timestamp 0
transform 1 0 850 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1176_
timestamp 0
transform 1 0 1130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1177_
timestamp 0
transform 1 0 1830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1178_
timestamp 0
transform 1 0 1970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1179_
timestamp 0
transform -1 0 2550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1180_
timestamp 0
transform -1 0 30 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1181_
timestamp 0
transform -1 0 1730 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1182_
timestamp 0
transform -1 0 2410 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1183_
timestamp 0
transform 1 0 1830 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1184_
timestamp 0
transform 1 0 1930 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1185_
timestamp 0
transform -1 0 1990 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1186_
timestamp 0
transform -1 0 1670 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1187_
timestamp 0
transform 1 0 1890 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1188_
timestamp 0
transform 1 0 2170 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1189_
timestamp 0
transform -1 0 1590 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1190_
timestamp 0
transform -1 0 2050 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1191_
timestamp 0
transform -1 0 1450 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1192_
timestamp 0
transform -1 0 970 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1193_
timestamp 0
transform -1 0 830 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1194_
timestamp 0
transform -1 0 450 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1195_
timestamp 0
transform 1 0 110 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1196_
timestamp 0
transform -1 0 590 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1197_
timestamp 0
transform 1 0 850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1198_
timestamp 0
transform -1 0 1010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1199_
timestamp 0
transform 1 0 1550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1200_
timestamp 0
transform 1 0 1270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1201_
timestamp 0
transform 1 0 1690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1202_
timestamp 0
transform -1 0 1310 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1203_
timestamp 0
transform 1 0 2110 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1204_
timestamp 0
transform 1 0 3190 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1205_
timestamp 0
transform -1 0 2450 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1206_
timestamp 0
transform -1 0 3050 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1207_
timestamp 0
transform 1 0 2670 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1208_
timestamp 0
transform 1 0 2690 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1209_
timestamp 0
transform -1 0 2850 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1210_
timestamp 0
transform 1 0 2970 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1211_
timestamp 0
transform -1 0 1810 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1212_
timestamp 0
transform -1 0 1170 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1213_
timestamp 0
transform -1 0 1070 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1214_
timestamp 0
transform 1 0 950 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1215_
timestamp 0
transform -1 0 590 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1216_
timestamp 0
transform 1 0 390 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1217_
timestamp 0
transform 1 0 810 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1218_
timestamp 0
transform 1 0 1290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1219_
timestamp 0
transform 1 0 1610 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1220_
timestamp 0
transform -1 0 2250 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1221_
timestamp 0
transform 1 0 2330 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1222_
timestamp 0
transform 1 0 2870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1223_
timestamp 0
transform -1 0 2570 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1224_
timestamp 0
transform 1 0 2750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1225_
timestamp 0
transform -1 0 2790 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1226_
timestamp 0
transform -1 0 3050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1227_
timestamp 0
transform 1 0 2930 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1228_
timestamp 0
transform -1 0 2990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1229_
timestamp 0
transform 1 0 3030 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1230_
timestamp 0
transform 1 0 3230 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1231_
timestamp 0
transform 1 0 1930 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1232_
timestamp 0
transform 1 0 2030 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1233_
timestamp 0
transform -1 0 2490 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1234_
timestamp 0
transform 1 0 1190 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1235_
timestamp 0
transform 1 0 1330 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1236_
timestamp 0
transform -1 0 270 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1237_
timestamp 0
transform 1 0 530 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1238_
timestamp 0
transform 1 0 670 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1239_
timestamp 0
transform 1 0 1970 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1240_
timestamp 0
transform -1 0 2090 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1241_
timestamp 0
transform 1 0 1690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1242_
timestamp 0
transform 1 0 2170 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1243_
timestamp 0
transform -1 0 2650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1244_
timestamp 0
transform -1 0 1290 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1245_
timestamp 0
transform -1 0 850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1246_
timestamp 0
transform -1 0 450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1247_
timestamp 0
transform 1 0 2370 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1248_
timestamp 0
transform -1 0 1370 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1249_
timestamp 0
transform -1 0 2270 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1250_
timestamp 0
transform -1 0 2070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1251_
timestamp 0
transform 1 0 1990 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1252_
timestamp 0
transform -1 0 1750 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1253_
timestamp 0
transform -1 0 1230 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1254_
timestamp 0
transform 1 0 2110 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1255_
timestamp 0
transform 1 0 1870 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1256_
timestamp 0
transform -1 0 1610 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1257_
timestamp 0
transform -1 0 950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1258_
timestamp 0
transform 1 0 150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1259_
timestamp 0
transform 1 0 1990 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1260_
timestamp 0
transform -1 0 1850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1261_
timestamp 0
transform -1 0 1870 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1262_
timestamp 0
transform -1 0 2410 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1263_
timestamp 0
transform -1 0 2130 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1264_
timestamp 0
transform -1 0 1610 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1265_
timestamp 0
transform -1 0 1270 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1266_
timestamp 0
transform 1 0 1730 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1267_
timestamp 0
transform 1 0 2530 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1268_
timestamp 0
transform -1 0 1370 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1269_
timestamp 0
transform -1 0 1130 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1270_
timestamp 0
transform 1 0 850 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1271_
timestamp 0
transform -1 0 430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1272_
timestamp 0
transform 1 0 1710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1273_
timestamp 0
transform 1 0 1450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1274_
timestamp 0
transform 1 0 1650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1275_
timestamp 0
transform -1 0 1350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1276_
timestamp 0
transform -1 0 310 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1277_
timestamp 0
transform -1 0 810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1278_
timestamp 0
transform 1 0 1610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1279_
timestamp 0
transform 1 0 1470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1280_
timestamp 0
transform 1 0 570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1281_
timestamp 0
transform -1 0 170 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1282_
timestamp 0
transform 1 0 970 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1283_
timestamp 0
transform 1 0 810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1284_
timestamp 0
transform -1 0 430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1285_
timestamp 0
transform -1 0 430 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1286_
timestamp 0
transform -1 0 30 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1287_
timestamp 0
transform -1 0 30 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1288_
timestamp 0
transform -1 0 710 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1289_
timestamp 0
transform -1 0 30 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1290_
timestamp 0
transform -1 0 150 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1291_
timestamp 0
transform 1 0 150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1292_
timestamp 0
transform -1 0 1090 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1293_
timestamp 0
transform 1 0 290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1294_
timestamp 0
transform -1 0 290 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1295_
timestamp 0
transform -1 0 790 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1296_
timestamp 0
transform 1 0 290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1297_
timestamp 0
transform -1 0 310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1298_
timestamp 0
transform -1 0 930 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1299_
timestamp 0
transform -1 0 30 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1300_
timestamp 0
transform -1 0 30 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1301_
timestamp 0
transform 1 0 810 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1302_
timestamp 0
transform -1 0 730 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1303_
timestamp 0
transform 1 0 290 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1304_
timestamp 0
transform 1 0 150 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1305_
timestamp 0
transform 1 0 570 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1306_
timestamp 0
transform 1 0 950 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1307_
timestamp 0
transform 1 0 1130 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1308_
timestamp 0
transform -1 0 450 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1309_
timestamp 0
transform 1 0 710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1310_
timestamp 0
transform 1 0 1090 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1311_
timestamp 0
transform 1 0 2270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1312_
timestamp 0
transform 1 0 2370 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1313_
timestamp 0
transform 1 0 2110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1314_
timestamp 0
transform 1 0 1830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1315_
timestamp 0
transform 1 0 1430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1316_
timestamp 0
transform 1 0 1550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1317_
timestamp 0
transform 1 0 1930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1318_
timestamp 0
transform 1 0 2070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1319_
timestamp 0
transform 1 0 2350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1320_
timestamp 0
transform -1 0 2270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1321_
timestamp 0
transform -1 0 2110 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1322_
timestamp 0
transform -1 0 2430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1323_
timestamp 0
transform 1 0 2470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1324_
timestamp 0
transform 1 0 3430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1325_
timestamp 0
transform -1 0 3310 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1326_
timestamp 0
transform 1 0 3230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1327_
timestamp 0
transform 1 0 3370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1328_
timestamp 0
transform -1 0 3670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1329_
timestamp 0
transform -1 0 3530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1330_
timestamp 0
transform 1 0 3510 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1331_
timestamp 0
transform 1 0 3370 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1332_
timestamp 0
transform 1 0 2730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1333_
timestamp 0
transform -1 0 2810 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1334_
timestamp 0
transform 1 0 3430 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1335_
timestamp 0
transform 1 0 2890 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1336_
timestamp 0
transform 1 0 430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1337_
timestamp 0
transform 1 0 570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1338_
timestamp 0
transform -1 0 1470 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1339_
timestamp 0
transform 1 0 150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1340_
timestamp 0
transform 1 0 430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1341_
timestamp 0
transform -1 0 1330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1342_
timestamp 0
transform 1 0 810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1343_
timestamp 0
transform -1 0 1450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1344_
timestamp 0
transform -1 0 1470 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1345_
timestamp 0
transform 1 0 1050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1346_
timestamp 0
transform 1 0 1170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1347_
timestamp 0
transform 1 0 910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1348_
timestamp 0
transform -1 0 970 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1349_
timestamp 0
transform 1 0 1090 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1350_
timestamp 0
transform -1 0 690 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1351_
timestamp 0
transform 1 0 690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1352_
timestamp 0
transform -1 0 310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1353_
timestamp 0
transform -1 0 170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1354_
timestamp 0
transform 1 0 2050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1355_
timestamp 0
transform 1 0 2090 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1356_
timestamp 0
transform -1 0 2450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1357_
timestamp 0
transform -1 0 3090 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1358_
timestamp 0
transform -1 0 2330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1359_
timestamp 0
transform 1 0 2690 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1360_
timestamp 0
transform 1 0 2190 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1361_
timestamp 0
transform -1 0 1970 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1362_
timestamp 0
transform 1 0 3230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1363_
timestamp 0
transform -1 0 2190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1364_
timestamp 0
transform 1 0 2250 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1365_
timestamp 0
transform -1 0 1790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1366_
timestamp 0
transform 1 0 1650 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1367_
timestamp 0
transform -1 0 1930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1368_
timestamp 0
transform -1 0 1830 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1369_
timestamp 0
transform -1 0 1410 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1370_
timestamp 0
transform -1 0 1530 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1371_
timestamp 0
transform -1 0 30 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1372_
timestamp 0
transform -1 0 30 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1373_
timestamp 0
transform 1 0 690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1374_
timestamp 0
transform -1 0 570 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1375_
timestamp 0
transform -1 0 430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1376_
timestamp 0
transform -1 0 150 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1377_
timestamp 0
transform -1 0 550 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1378_
timestamp 0
transform -1 0 570 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1379_
timestamp 0
transform -1 0 150 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1380_
timestamp 0
transform 1 0 390 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1381_
timestamp 0
transform 1 0 710 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1382_
timestamp 0
transform 1 0 410 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1383_
timestamp 0
transform -1 0 650 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1384_
timestamp 0
transform -1 0 270 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1385_
timestamp 0
transform -1 0 30 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1386_
timestamp 0
transform -1 0 30 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1387_
timestamp 0
transform 1 0 150 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1388_
timestamp 0
transform 1 0 430 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1389_
timestamp 0
transform 1 0 1050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1390_
timestamp 0
transform 1 0 810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1391_
timestamp 0
transform 1 0 570 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1392_
timestamp 0
transform 1 0 290 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1393_
timestamp 0
transform 1 0 670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1394_
timestamp 0
transform 1 0 1190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1395_
timestamp 0
transform 1 0 910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1396_
timestamp 0
transform -1 0 550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1397_
timestamp 0
transform 1 0 1090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1398_
timestamp 0
transform 1 0 1930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1399_
timestamp 0
transform 1 0 2490 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1400_
timestamp 0
transform -1 0 2550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1401_
timestamp 0
transform -1 0 1010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1402_
timestamp 0
transform 1 0 850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1403_
timestamp 0
transform 1 0 1250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1404_
timestamp 0
transform -1 0 1070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1405_
timestamp 0
transform -1 0 1830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1406_
timestamp 0
transform 1 0 2670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1407_
timestamp 0
transform 1 0 2750 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1408_
timestamp 0
transform 1 0 3150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1409_
timestamp 0
transform 1 0 3570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1410_
timestamp 0
transform 1 0 3290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1411_
timestamp 0
transform 1 0 3430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1412_
timestamp 0
transform -1 0 2910 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1413_
timestamp 0
transform 1 0 2830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1414_
timestamp 0
transform 1 0 3910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1415_
timestamp 0
transform 1 0 2330 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1416_
timestamp 0
transform 1 0 2410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1417_
timestamp 0
transform 1 0 2550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1418_
timestamp 0
transform 1 0 810 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1419_
timestamp 0
transform -1 0 590 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1420_
timestamp 0
transform -1 0 30 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1421_
timestamp 0
transform -1 0 1570 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1422_
timestamp 0
transform 1 0 1670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1423_
timestamp 0
transform 1 0 2170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1424_
timestamp 0
transform 1 0 2290 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1425_
timestamp 0
transform 1 0 2050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1426_
timestamp 0
transform -1 0 1930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1427_
timestamp 0
transform -1 0 1790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1428_
timestamp 0
transform 1 0 2410 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1429_
timestamp 0
transform 1 0 2290 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1430_
timestamp 0
transform -1 0 2170 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1431_
timestamp 0
transform 1 0 1370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1432_
timestamp 0
transform 1 0 1330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1433_
timestamp 0
transform 1 0 2530 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1434_
timestamp 0
transform 1 0 2690 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1435_
timestamp 0
transform 1 0 2730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1436_
timestamp 0
transform 1 0 3310 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1437_
timestamp 0
transform 1 0 2630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1438_
timestamp 0
transform -1 0 2550 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1439_
timestamp 0
transform -1 0 2590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1440_
timestamp 0
transform 1 0 2430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1441_
timestamp 0
transform -1 0 2570 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1442_
timestamp 0
transform -1 0 2310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1443_
timestamp 0
transform 1 0 1890 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1444_
timestamp 0
transform -1 0 1230 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1445_
timestamp 0
transform -1 0 1370 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1446_
timestamp 0
transform -1 0 730 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1447_
timestamp 0
transform -1 0 590 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1448_
timestamp 0
transform -1 0 1630 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1449_
timestamp 0
transform 1 0 1490 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1450_
timestamp 0
transform -1 0 1770 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1451_
timestamp 0
transform -1 0 830 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1452_
timestamp 0
transform -1 0 30 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1453_
timestamp 0
transform 1 0 270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1454_
timestamp 0
transform -1 0 1230 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1455_
timestamp 0
transform -1 0 970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1456_
timestamp 0
transform 1 0 1090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1457_
timestamp 0
transform -1 0 830 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1458_
timestamp 0
transform -1 0 310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1459_
timestamp 0
transform -1 0 170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1460_
timestamp 0
transform 1 0 150 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1461_
timestamp 0
transform -1 0 450 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1462_
timestamp 0
transform 1 0 670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1463_
timestamp 0
transform -1 0 1150 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1464_
timestamp 0
transform 1 0 1190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1465_
timestamp 0
transform 1 0 850 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1466_
timestamp 0
transform 1 0 990 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1467_
timestamp 0
transform 1 0 1250 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1468_
timestamp 0
transform -1 0 1570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1469_
timestamp 0
transform 1 0 2470 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1470_
timestamp 0
transform -1 0 2230 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1471_
timestamp 0
transform -1 0 2630 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1472_
timestamp 0
transform -1 0 2890 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1473_
timestamp 0
transform -1 0 2770 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1474_
timestamp 0
transform 1 0 2810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1475_
timestamp 0
transform 1 0 3310 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1476_
timestamp 0
transform -1 0 2910 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1477_
timestamp 0
transform 1 0 3110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1478_
timestamp 0
transform 1 0 3250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1479_
timestamp 0
transform 1 0 3590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1480_
timestamp 0
transform -1 0 3190 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1481_
timestamp 0
transform -1 0 3030 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1482_
timestamp 0
transform 1 0 4070 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1483_
timestamp 0
transform -1 0 2570 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1484_
timestamp 0
transform -1 0 3370 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1485_
timestamp 0
transform 1 0 3330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1486_
timestamp 0
transform 1 0 2910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1487_
timestamp 0
transform -1 0 2030 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1488_
timestamp 0
transform -1 0 1250 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1489_
timestamp 0
transform 1 0 1090 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1490_
timestamp 0
transform 1 0 2750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1491_
timestamp 0
transform -1 0 3090 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1492_
timestamp 0
transform 1 0 2850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1493_
timestamp 0
transform -1 0 2670 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1494_
timestamp 0
transform -1 0 2830 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1495_
timestamp 0
transform 1 0 2930 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1496_
timestamp 0
transform 1 0 3170 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1497_
timestamp 0
transform -1 0 3450 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1498_
timestamp 0
transform 1 0 3010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1499_
timestamp 0
transform -1 0 3150 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1500_
timestamp 0
transform -1 0 3770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1501_
timestamp 0
transform 1 0 4110 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1502_
timestamp 0
transform 1 0 3990 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1503_
timestamp 0
transform 1 0 4390 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1504_
timestamp 0
transform -1 0 3890 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1505_
timestamp 0
transform -1 0 3610 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1506_
timestamp 0
transform -1 0 3750 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1507_
timestamp 0
transform 1 0 3310 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1508_
timestamp 0
transform -1 0 1770 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1509_
timestamp 0
transform -1 0 3190 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1510_
timestamp 0
transform -1 0 1490 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1511_
timestamp 0
transform 1 0 950 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1512_
timestamp 0
transform 1 0 1990 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1513_
timestamp 0
transform -1 0 1630 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1514_
timestamp 0
transform 1 0 1330 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1515_
timestamp 0
transform 1 0 1630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1516_
timestamp 0
transform -1 0 1870 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1517_
timestamp 0
transform -1 0 1910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1518_
timestamp 0
transform -1 0 1790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1519_
timestamp 0
transform 1 0 1490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1520_
timestamp 0
transform 1 0 290 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1521_
timestamp 0
transform 1 0 430 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1522_
timestamp 0
transform 1 0 2030 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1523_
timestamp 0
transform -1 0 2610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1524_
timestamp 0
transform 1 0 3110 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1525_
timestamp 0
transform 1 0 2970 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1526_
timestamp 0
transform -1 0 2970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1527_
timestamp 0
transform 1 0 3050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1528_
timestamp 0
transform 1 0 3190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1529_
timestamp 0
transform 1 0 2610 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1530_
timestamp 0
transform -1 0 3130 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1531_
timestamp 0
transform 1 0 2170 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1532_
timestamp 0
transform -1 0 2450 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1533_
timestamp 0
transform -1 0 2310 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1534_
timestamp 0
transform 1 0 2730 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1535_
timestamp 0
transform 1 0 2870 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1536_
timestamp 0
transform 1 0 3270 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1537_
timestamp 0
transform 1 0 2170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1538_
timestamp 0
transform -1 0 2310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1539_
timestamp 0
transform -1 0 2890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1540_
timestamp 0
transform -1 0 2510 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1541_
timestamp 0
transform 1 0 3530 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1542_
timestamp 0
transform 1 0 3970 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1543_
timestamp 0
transform 1 0 3870 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1544_
timestamp 0
transform 1 0 3890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1545_
timestamp 0
transform -1 0 4270 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1546_
timestamp 0
transform -1 0 3710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1547_
timestamp 0
transform 1 0 3770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1548_
timestamp 0
transform 1 0 4090 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1549_
timestamp 0
transform -1 0 3390 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1550_
timestamp 0
transform -1 0 3470 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1551_
timestamp 0
transform -1 0 3290 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1552_
timestamp 0
transform -1 0 3150 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1553_
timestamp 0
transform 1 0 2870 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1554_
timestamp 0
transform -1 0 2250 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1555_
timestamp 0
transform -1 0 2750 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1556_
timestamp 0
transform -1 0 2370 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1557_
timestamp 0
transform -1 0 2110 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1558_
timestamp 0
transform 1 0 2530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1559_
timestamp 0
transform -1 0 2650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1560_
timestamp 0
transform 1 0 2790 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1561_
timestamp 0
transform 1 0 2910 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1562_
timestamp 0
transform 1 0 2390 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1563_
timestamp 0
transform -1 0 2970 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1564_
timestamp 0
transform 1 0 2650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1565_
timestamp 0
transform 1 0 3130 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1566_
timestamp 0
transform 1 0 3010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1567_
timestamp 0
transform -1 0 2610 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1568_
timestamp 0
transform 1 0 2970 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1569_
timestamp 0
transform 1 0 3150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1570_
timestamp 0
transform 1 0 3290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1571_
timestamp 0
transform -1 0 2870 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1572_
timestamp 0
transform 1 0 3250 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1573_
timestamp 0
transform -1 0 2730 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1574_
timestamp 0
transform 1 0 2770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1575_
timestamp 0
transform 1 0 3390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1576_
timestamp 0
transform 1 0 3670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1577_
timestamp 0
transform 1 0 4010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1578_
timestamp 0
transform -1 0 3730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1579_
timestamp 0
transform 1 0 1690 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1580_
timestamp 0
transform 1 0 1550 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1581_
timestamp 0
transform 1 0 1710 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1582_
timestamp 0
transform -1 0 3750 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1583_
timestamp 0
transform 1 0 3590 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1584_
timestamp 0
transform -1 0 3470 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1585_
timestamp 0
transform 1 0 3370 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1586_
timestamp 0
transform -1 0 3570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1587_
timestamp 0
transform -1 0 3830 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1588_
timestamp 0
transform 1 0 3630 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1589_
timestamp 0
transform -1 0 3770 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1590_
timestamp 0
transform -1 0 3390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1591_
timestamp 0
transform 1 0 3530 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1592_
timestamp 0
transform 1 0 2990 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1593_
timestamp 0
transform -1 0 3570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1594_
timestamp 0
transform -1 0 3450 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1595_
timestamp 0
transform 1 0 3170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1596_
timestamp 0
transform -1 0 3050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1597_
timestamp 0
transform -1 0 2930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1598_
timestamp 0
transform 1 0 3030 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__1599_
timestamp 0
transform 1 0 2590 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1600_
timestamp 0
transform -1 0 2790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1601_
timestamp 0
transform 1 0 3110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1602_
timestamp 0
transform -1 0 3410 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1603_
timestamp 0
transform 1 0 3510 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1604_
timestamp 0
transform 1 0 3530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1605_
timestamp 0
transform 1 0 3650 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1606_
timestamp 0
transform -1 0 3350 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1607_
timestamp 0
transform -1 0 2730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1608_
timestamp 0
transform 1 0 3930 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1609_
timestamp 0
transform 1 0 3790 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1610_
timestamp 0
transform 1 0 1830 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1611_
timestamp 0
transform 1 0 2490 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1612_
timestamp 0
transform -1 0 3590 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1613_
timestamp 0
transform -1 0 3450 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1614_
timestamp 0
transform 1 0 3290 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1615_
timestamp 0
transform -1 0 3410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1616_
timestamp 0
transform -1 0 3230 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1617_
timestamp 0
transform -1 0 3230 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1618_
timestamp 0
transform -1 0 3290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1619_
timestamp 0
transform -1 0 3310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__1620_
timestamp 0
transform -1 0 3290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1621_
timestamp 0
transform 1 0 3330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1622_
timestamp 0
transform 1 0 3470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1623_
timestamp 0
transform 1 0 3710 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1624_
timestamp 0
transform -1 0 3610 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1625_
timestamp 0
transform -1 0 3390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1626_
timestamp 0
transform -1 0 2870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1627_
timestamp 0
transform -1 0 3010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1628_
timestamp 0
transform -1 0 3510 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1629_
timestamp 0
transform 1 0 3350 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1630_
timestamp 0
transform -1 0 3150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1631_
timestamp 0
transform 1 0 2490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1632_
timestamp 0
transform 1 0 2210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1633_
timestamp 0
transform 1 0 2630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1634_
timestamp 0
transform -1 0 3350 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1635_
timestamp 0
transform 1 0 2630 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1636_
timestamp 0
transform 1 0 2890 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1637_
timestamp 0
transform -1 0 3070 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1638_
timestamp 0
transform -1 0 3810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1639_
timestamp 0
transform 1 0 3510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1640_
timestamp 0
transform 1 0 3610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1641_
timestamp 0
transform 1 0 3650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1642_
timestamp 0
transform 1 0 2390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1643_
timestamp 0
transform 1 0 2770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1644_
timestamp 0
transform 1 0 2910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1645_
timestamp 0
transform 1 0 3190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1646_
timestamp 0
transform 1 0 3050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1647_
timestamp 0
transform 1 0 3310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1648_
timestamp 0
transform -1 0 3710 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1649_
timestamp 0
transform 1 0 4690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1650_
timestamp 0
transform 1 0 4550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1651_
timestamp 0
transform 1 0 5070 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1652_
timestamp 0
transform 1 0 4930 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1653_
timestamp 0
transform 1 0 4550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1654_
timestamp 0
transform -1 0 4690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1655_
timestamp 0
transform 1 0 4950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1656_
timestamp 0
transform 1 0 4810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1657_
timestamp 0
transform 1 0 5570 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1658_
timestamp 0
transform 1 0 5430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__1659_
timestamp 0
transform 1 0 4930 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1660_
timestamp 0
transform -1 0 5070 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1661_
timestamp 0
transform 1 0 5210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1662_
timestamp 0
transform 1 0 5070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1663_
timestamp 0
transform 1 0 4990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1664_
timestamp 0
transform -1 0 4870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1692_
timestamp 0
transform 1 0 5330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1693_
timestamp 0
transform 1 0 5430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1694_
timestamp 0
transform 1 0 5430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1695_
timestamp 0
transform -1 0 5570 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1696_
timestamp 0
transform 1 0 5610 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1697_
timestamp 0
transform -1 0 5230 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1698_
timestamp 0
transform -1 0 5330 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1699_
timestamp 0
transform -1 0 5130 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1700_
timestamp 0
transform -1 0 4430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1701_
timestamp 0
transform -1 0 4530 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1702_
timestamp 0
transform 1 0 4530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1703_
timestamp 0
transform 1 0 5510 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__1704_
timestamp 0
transform 1 0 4750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1705_
timestamp 0
transform 1 0 4370 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1706_
timestamp 0
transform -1 0 4710 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1707_
timestamp 0
transform 1 0 4830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1708_
timestamp 0
transform -1 0 4650 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1709_
timestamp 0
transform 1 0 4690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1710_
timestamp 0
transform 1 0 5190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1711_
timestamp 0
transform 1 0 5050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1712_
timestamp 0
transform -1 0 5290 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1713_
timestamp 0
transform -1 0 5250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1714_
timestamp 0
transform 1 0 5270 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1715_
timestamp 0
transform 1 0 5510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1716_
timestamp 0
transform -1 0 5430 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1717_
timestamp 0
transform 1 0 5430 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1718_
timestamp 0
transform -1 0 4870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1719_
timestamp 0
transform -1 0 5170 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1720_
timestamp 0
transform -1 0 5390 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1721_
timestamp 0
transform -1 0 4450 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1722_
timestamp 0
transform -1 0 4390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1723_
timestamp 0
transform 1 0 4210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1724_
timestamp 0
transform 1 0 4050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1725_
timestamp 0
transform -1 0 4170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1726_
timestamp 0
transform 1 0 4270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1727_
timestamp 0
transform 1 0 4290 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1728_
timestamp 0
transform 1 0 3450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1729_
timestamp 0
transform -1 0 3430 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1730_
timestamp 0
transform -1 0 3570 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1731_
timestamp 0
transform 1 0 3650 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1732_
timestamp 0
transform -1 0 3810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1733_
timestamp 0
transform 1 0 3950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1734_
timestamp 0
transform -1 0 5070 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1735_
timestamp 0
transform -1 0 4930 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1736_
timestamp 0
transform 1 0 4830 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1737_
timestamp 0
transform 1 0 4550 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1738_
timestamp 0
transform 1 0 4990 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1739_
timestamp 0
transform 1 0 5090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1740_
timestamp 0
transform 1 0 4950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1741_
timestamp 0
transform 1 0 4750 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1742_
timestamp 0
transform -1 0 4070 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1743_
timestamp 0
transform 1 0 3910 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1744_
timestamp 0
transform -1 0 3810 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1745_
timestamp 0
transform 1 0 3850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1746_
timestamp 0
transform -1 0 3710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1747_
timestamp 0
transform 1 0 4190 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1748_
timestamp 0
transform -1 0 4130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1749_
timestamp 0
transform -1 0 4650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1750_
timestamp 0
transform 1 0 3830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1751_
timestamp 0
transform -1 0 3950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1752_
timestamp 0
transform -1 0 3890 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1753_
timestamp 0
transform -1 0 4150 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1754_
timestamp 0
transform 1 0 3990 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1755_
timestamp 0
transform 1 0 4070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1756_
timestamp 0
transform -1 0 3570 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1757_
timestamp 0
transform 1 0 3850 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1758_
timestamp 0
transform 1 0 4270 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1759_
timestamp 0
transform -1 0 4650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1760_
timestamp 0
transform 1 0 4470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1761_
timestamp 0
transform -1 0 4370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1762_
timestamp 0
transform -1 0 4150 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1763_
timestamp 0
transform -1 0 4010 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1764_
timestamp 0
transform -1 0 3990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1765_
timestamp 0
transform 1 0 4230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1766_
timestamp 0
transform 1 0 4130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1767_
timestamp 0
transform 1 0 4410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1768_
timestamp 0
transform -1 0 4070 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1769_
timestamp 0
transform 1 0 4670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1770_
timestamp 0
transform -1 0 4410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1771_
timestamp 0
transform -1 0 4330 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1772_
timestamp 0
transform -1 0 4450 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1773_
timestamp 0
transform -1 0 4270 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1774_
timestamp 0
transform 1 0 4530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1775_
timestamp 0
transform -1 0 4490 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1776_
timestamp 0
transform 1 0 4610 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1777_
timestamp 0
transform 1 0 4910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1778_
timestamp 0
transform 1 0 4770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1779_
timestamp 0
transform 1 0 4750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1780_
timestamp 0
transform 1 0 4510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1781_
timestamp 0
transform -1 0 4210 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1782_
timestamp 0
transform 1 0 4290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1783_
timestamp 0
transform -1 0 2790 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1784_
timestamp 0
transform -1 0 3570 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1785_
timestamp 0
transform -1 0 3670 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1786_
timestamp 0
transform -1 0 4170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1787_
timestamp 0
transform 1 0 4330 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1788_
timestamp 0
transform 1 0 4990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1789_
timestamp 0
transform 1 0 4850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1790_
timestamp 0
transform 1 0 5090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1791_
timestamp 0
transform 1 0 5550 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1792_
timestamp 0
transform 1 0 5510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1793_
timestamp 0
transform 1 0 5350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1794_
timestamp 0
transform 1 0 5350 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1795_
timestamp 0
transform -1 0 5230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1796_
timestamp 0
transform 1 0 5470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1797_
timestamp 0
transform -1 0 5350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1798_
timestamp 0
transform 1 0 4570 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1799_
timestamp 0
transform 1 0 4710 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1800_
timestamp 0
transform 1 0 4170 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1801_
timestamp 0
transform -1 0 3950 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1802_
timestamp 0
transform -1 0 3810 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1803_
timestamp 0
transform 1 0 3670 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1804_
timestamp 0
transform 1 0 3790 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1805_
timestamp 0
transform -1 0 4330 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1806_
timestamp 0
transform 1 0 4350 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1807_
timestamp 0
transform 1 0 4230 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1808_
timestamp 0
transform -1 0 4670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1809_
timestamp 0
transform -1 0 4810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1810_
timestamp 0
transform -1 0 4890 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1811_
timestamp 0
transform -1 0 4770 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1812_
timestamp 0
transform 1 0 4590 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1813_
timestamp 0
transform 1 0 5050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1814_
timestamp 0
transform -1 0 4930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1815_
timestamp 0
transform 1 0 4870 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1816_
timestamp 0
transform 1 0 5010 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1817_
timestamp 0
transform 1 0 5230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1818_
timestamp 0
transform 1 0 5090 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1819_
timestamp 0
transform -1 0 4430 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1820_
timestamp 0
transform 1 0 4470 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1821_
timestamp 0
transform -1 0 4890 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1822_
timestamp 0
transform 1 0 4750 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1823_
timestamp 0
transform -1 0 4070 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1824_
timestamp 0
transform 1 0 4970 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1825_
timestamp 0
transform 1 0 4850 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1826_
timestamp 0
transform -1 0 5350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1827_
timestamp 0
transform -1 0 5190 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1828_
timestamp 0
transform 1 0 5010 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1829_
timestamp 0
transform 1 0 5190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1830_
timestamp 0
transform 1 0 4950 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1831_
timestamp 0
transform 1 0 5050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1832_
timestamp 0
transform 1 0 5190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1833_
timestamp 0
transform 1 0 5490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1834_
timestamp 0
transform 1 0 5530 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1835_
timestamp 0
transform -1 0 4550 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1836_
timestamp 0
transform 1 0 4610 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1837_
timestamp 0
transform -1 0 5630 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1838_
timestamp 0
transform -1 0 4670 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1839_
timestamp 0
transform 1 0 4290 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1840_
timestamp 0
transform -1 0 5630 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1841_
timestamp 0
transform 1 0 4790 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1842_
timestamp 0
transform 1 0 5570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1843_
timestamp 0
transform 1 0 5470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1844_
timestamp 0
transform 1 0 4850 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1845_
timestamp 0
transform 1 0 5170 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1846_
timestamp 0
transform 1 0 5470 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1847_
timestamp 0
transform -1 0 5350 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1848_
timestamp 0
transform -1 0 5530 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1849_
timestamp 0
transform 1 0 5210 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1850_
timestamp 0
transform 1 0 5570 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1851_
timestamp 0
transform -1 0 5450 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1852_
timestamp 0
transform -1 0 5350 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1853_
timestamp 0
transform -1 0 4950 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1854_
timestamp 0
transform 1 0 5390 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1855_
timestamp 0
transform -1 0 5070 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1856_
timestamp 0
transform -1 0 4430 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1857_
timestamp 0
transform -1 0 3910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1858_
timestamp 0
transform -1 0 3950 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1859_
timestamp 0
transform 1 0 3990 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1860_
timestamp 0
transform 1 0 4050 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1861_
timestamp 0
transform -1 0 4170 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1862_
timestamp 0
transform -1 0 4130 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1863_
timestamp 0
transform -1 0 3870 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1864_
timestamp 0
transform -1 0 5210 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1865_
timestamp 0
transform -1 0 5490 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1866_
timestamp 0
transform 1 0 4350 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1867_
timestamp 0
transform -1 0 3930 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1868_
timestamp 0
transform 1 0 4450 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1869_
timestamp 0
transform -1 0 5310 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1870_
timestamp 0
transform -1 0 4850 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1871_
timestamp 0
transform -1 0 5130 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1872_
timestamp 0
transform -1 0 4710 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1873_
timestamp 0
transform -1 0 4950 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1874_
timestamp 0
transform 1 0 5490 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1875_
timestamp 0
transform 1 0 5250 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1876_
timestamp 0
transform -1 0 5050 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1877_
timestamp 0
transform -1 0 4570 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1878_
timestamp 0
transform -1 0 3850 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1879_
timestamp 0
transform -1 0 3790 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1880_
timestamp 0
transform -1 0 5630 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1881_
timestamp 0
transform 1 0 5490 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1882_
timestamp 0
transform -1 0 5370 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1883_
timestamp 0
transform -1 0 5250 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1884_
timestamp 0
transform -1 0 5130 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1885_
timestamp 0
transform 1 0 5370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1886_
timestamp 0
transform -1 0 4730 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1887_
timestamp 0
transform -1 0 4630 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1888_
timestamp 0
transform -1 0 4490 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1889_
timestamp 0
transform 1 0 4230 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1890_
timestamp 0
transform -1 0 3710 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1891_
timestamp 0
transform -1 0 4110 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1892_
timestamp 0
transform -1 0 3590 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1893_
timestamp 0
transform -1 0 3470 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1894_
timestamp 0
transform -1 0 2650 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1895_
timestamp 0
transform -1 0 2630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1896_
timestamp 0
transform -1 0 30 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1897_
timestamp 0
transform 1 0 2650 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1898_
timestamp 0
transform -1 0 3130 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1899_
timestamp 0
transform 1 0 3530 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1900_
timestamp 0
transform -1 0 3250 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1901_
timestamp 0
transform -1 0 3670 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1902_
timestamp 0
transform -1 0 3990 0 -1 250
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert0
timestamp 0
transform -1 0 2370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert1
timestamp 0
transform -1 0 2490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert2
timestamp 0
transform 1 0 4050 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert3
timestamp 0
transform 1 0 4510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert4
timestamp 0
transform -1 0 3770 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert5
timestamp 0
transform 1 0 1730 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert6
timestamp 0
transform -1 0 1610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert7
timestamp 0
transform 1 0 3710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert8
timestamp 0
transform -1 0 4690 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert9
timestamp 0
transform 1 0 5030 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert10
timestamp 0
transform -1 0 5210 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert11
timestamp 0
transform 1 0 5490 0 -1 250
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert17
timestamp 0
transform -1 0 3890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert18
timestamp 0
transform 1 0 3990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert19
timestamp 0
transform 1 0 5110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert20
timestamp 0
transform 1 0 5310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert21
timestamp 0
transform 1 0 2350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert22
timestamp 0
transform 1 0 5550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert23
timestamp 0
transform -1 0 2250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert24
timestamp 0
transform 1 0 2990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert25
timestamp 0
transform 1 0 2670 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert26
timestamp 0
transform 1 0 1610 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert27
timestamp 0
transform -1 0 3490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert28
timestamp 0
transform -1 0 1490 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert29
timestamp 0
transform -1 0 5410 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert30
timestamp 0
transform 1 0 5150 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert31
timestamp 0
transform 1 0 4750 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert32
timestamp 0
transform 1 0 4950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert12
timestamp 0
transform 1 0 4050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert13
timestamp 0
transform -1 0 4070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert14
timestamp 0
transform 1 0 3490 0 1 5530
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert15
timestamp 0
transform -1 0 3830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert16
timestamp 0
transform 1 0 4370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__927_
timestamp 0
transform -1 0 4290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__928_
timestamp 0
transform 1 0 3810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__929_
timestamp 0
transform -1 0 3870 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__930_
timestamp 0
transform 1 0 3970 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__931_
timestamp 0
transform 1 0 4170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__932_
timestamp 0
transform -1 0 2870 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__933_
timestamp 0
transform 1 0 4370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__934_
timestamp 0
transform -1 0 4630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__935_
timestamp 0
transform 1 0 5550 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__936_
timestamp 0
transform 1 0 4490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__937_
timestamp 0
transform 1 0 4810 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__938_
timestamp 0
transform -1 0 4990 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__939_
timestamp 0
transform -1 0 4850 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__940_
timestamp 0
transform -1 0 4090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__941_
timestamp 0
transform -1 0 3630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__942_
timestamp 0
transform -1 0 4050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__943_
timestamp 0
transform -1 0 4330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__944_
timestamp 0
transform -1 0 3670 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__945_
timestamp 0
transform -1 0 3990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__946_
timestamp 0
transform 1 0 5090 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__947_
timestamp 0
transform 1 0 4950 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__948_
timestamp 0
transform 1 0 4670 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__949_
timestamp 0
transform 1 0 4510 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__950_
timestamp 0
transform -1 0 4250 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__951_
timestamp 0
transform 1 0 4410 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__952_
timestamp 0
transform 1 0 4550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__953_
timestamp 0
transform 1 0 4490 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__954_
timestamp 0
transform 1 0 4970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__955_
timestamp 0
transform 1 0 5090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__956_
timestamp 0
transform 1 0 5350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__957_
timestamp 0
transform 1 0 5210 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__958_
timestamp 0
transform 1 0 5570 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__959_
timestamp 0
transform -1 0 5530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__960_
timestamp 0
transform 1 0 4170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__961_
timestamp 0
transform -1 0 4850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__962_
timestamp 0
transform 1 0 4690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__963_
timestamp 0
transform -1 0 5210 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__964_
timestamp 0
transform 1 0 4330 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__965_
timestamp 0
transform 1 0 4450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__966_
timestamp 0
transform 1 0 4310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__967_
timestamp 0
transform -1 0 4450 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__968_
timestamp 0
transform -1 0 4090 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__969_
timestamp 0
transform -1 0 4210 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__970_
timestamp 0
transform 1 0 5210 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__971_
timestamp 0
transform -1 0 4330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__972_
timestamp 0
transform -1 0 4450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__973_
timestamp 0
transform -1 0 5370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__974_
timestamp 0
transform 1 0 4190 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__975_
timestamp 0
transform -1 0 4330 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__976_
timestamp 0
transform -1 0 5350 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__977_
timestamp 0
transform -1 0 5450 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__978_
timestamp 0
transform 1 0 5490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__979_
timestamp 0
transform -1 0 5250 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__980_
timestamp 0
transform 1 0 4970 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__981_
timestamp 0
transform -1 0 5110 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__982_
timestamp 0
transform 1 0 4610 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__983_
timestamp 0
transform -1 0 4150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__984_
timestamp 0
transform -1 0 4270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__985_
timestamp 0
transform -1 0 3210 0 1 730
box -6 -8 26 248
use FILL  FILL_1__986_
timestamp 0
transform 1 0 5310 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__987_
timestamp 0
transform 1 0 5170 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__988_
timestamp 0
transform -1 0 3070 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__989_
timestamp 0
transform -1 0 2710 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__990_
timestamp 0
transform 1 0 2470 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__991_
timestamp 0
transform 1 0 2450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__992_
timestamp 0
transform 1 0 2590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__993_
timestamp 0
transform 1 0 2130 0 1 250
box -6 -8 26 248
use FILL  FILL_1__994_
timestamp 0
transform -1 0 2350 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__995_
timestamp 0
transform -1 0 1530 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__996_
timestamp 0
transform 1 0 1850 0 1 730
box -6 -8 26 248
use FILL  FILL_1__997_
timestamp 0
transform -1 0 2810 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__998_
timestamp 0
transform 1 0 2270 0 1 730
box -6 -8 26 248
use FILL  FILL_1__999_
timestamp 0
transform -1 0 2590 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1000_
timestamp 0
transform 1 0 1390 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1001_
timestamp 0
transform -1 0 1390 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1002_
timestamp 0
transform 1 0 2950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1003_
timestamp 0
transform -1 0 1490 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1004_
timestamp 0
transform -1 0 1770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1005_
timestamp 0
transform 1 0 1810 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1006_
timestamp 0
transform -1 0 1410 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1007_
timestamp 0
transform 1 0 1610 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1008_
timestamp 0
transform -1 0 1270 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1009_
timestamp 0
transform -1 0 910 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1010_
timestamp 0
transform 1 0 2470 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1011_
timestamp 0
transform 1 0 2570 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1012_
timestamp 0
transform 1 0 1990 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1013_
timestamp 0
transform 1 0 2570 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1014_
timestamp 0
transform 1 0 2310 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1015_
timestamp 0
transform -1 0 2350 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1016_
timestamp 0
transform 1 0 1030 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1017_
timestamp 0
transform -1 0 770 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1018_
timestamp 0
transform -1 0 1250 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1019_
timestamp 0
transform -1 0 1350 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1020_
timestamp 0
transform -1 0 990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1021_
timestamp 0
transform -1 0 1490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1022_
timestamp 0
transform -1 0 50 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1023_
timestamp 0
transform -1 0 1290 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1024_
timestamp 0
transform -1 0 50 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1025_
timestamp 0
transform 1 0 410 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1026_
timestamp 0
transform -1 0 1650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1027_
timestamp 0
transform -1 0 1130 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1028_
timestamp 0
transform -1 0 570 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1029_
timestamp 0
transform 1 0 690 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1030_
timestamp 0
transform -1 0 1550 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1031_
timestamp 0
transform -1 0 150 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1032_
timestamp 0
transform 1 0 270 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1033_
timestamp 0
transform -1 0 290 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1034_
timestamp 0
transform 1 0 2830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1035_
timestamp 0
transform 1 0 2730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1036_
timestamp 0
transform -1 0 2230 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1037_
timestamp 0
transform -1 0 2210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1038_
timestamp 0
transform 1 0 2510 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1039_
timestamp 0
transform 1 0 2450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1040_
timestamp 0
transform -1 0 2330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1041_
timestamp 0
transform 1 0 2050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1042_
timestamp 0
transform -1 0 1470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1043_
timestamp 0
transform -1 0 1830 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1044_
timestamp 0
transform -1 0 1930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1045_
timestamp 0
transform -1 0 1550 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1046_
timestamp 0
transform -1 0 710 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1047_
timestamp 0
transform 1 0 410 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1048_
timestamp 0
transform 1 0 830 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1049_
timestamp 0
transform 1 0 1670 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1050_
timestamp 0
transform 1 0 1110 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1051_
timestamp 0
transform -1 0 50 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1052_
timestamp 0
transform 1 0 170 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1053_
timestamp 0
transform 1 0 310 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1054_
timestamp 0
transform -1 0 570 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1055_
timestamp 0
transform 1 0 870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1056_
timestamp 0
transform -1 0 1550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1057_
timestamp 0
transform 1 0 1090 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1058_
timestamp 0
transform -1 0 1410 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1059_
timestamp 0
transform -1 0 2470 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1060_
timestamp 0
transform 1 0 1330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1061_
timestamp 0
transform -1 0 1270 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1062_
timestamp 0
transform -1 0 990 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1063_
timestamp 0
transform -1 0 770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1064_
timestamp 0
transform 1 0 730 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1065_
timestamp 0
transform -1 0 1430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1066_
timestamp 0
transform 1 0 1110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1067_
timestamp 0
transform 1 0 1470 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1068_
timestamp 0
transform 1 0 870 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1069_
timestamp 0
transform -1 0 750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1070_
timestamp 0
transform 1 0 130 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1071_
timestamp 0
transform -1 0 610 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1072_
timestamp 0
transform -1 0 470 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1073_
timestamp 0
transform -1 0 330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1074_
timestamp 0
transform -1 0 1890 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1075_
timestamp 0
transform -1 0 1870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1076_
timestamp 0
transform -1 0 2250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1077_
timestamp 0
transform -1 0 2270 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1078_
timestamp 0
transform 1 0 2130 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1079_
timestamp 0
transform 1 0 1690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1080_
timestamp 0
transform -1 0 2110 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1081_
timestamp 0
transform 1 0 1950 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1082_
timestamp 0
transform -1 0 1570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1083_
timestamp 0
transform 1 0 2090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1084_
timestamp 0
transform -1 0 2010 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1085_
timestamp 0
transform -1 0 1970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1086_
timestamp 0
transform -1 0 610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1087_
timestamp 0
transform -1 0 50 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1088_
timestamp 0
transform 1 0 450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1089_
timestamp 0
transform -1 0 610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1090_
timestamp 0
transform 1 0 730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1091_
timestamp 0
transform 1 0 170 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1092_
timestamp 0
transform -1 0 190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1093_
timestamp 0
transform -1 0 990 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1094_
timestamp 0
transform 1 0 310 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1095_
timestamp 0
transform -1 0 50 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1096_
timestamp 0
transform 1 0 590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1097_
timestamp 0
transform -1 0 3690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1098_
timestamp 0
transform -1 0 2210 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1099_
timestamp 0
transform -1 0 2070 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1100_
timestamp 0
transform 1 0 1930 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1101_
timestamp 0
transform -1 0 1810 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1102_
timestamp 0
transform -1 0 1030 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1103_
timestamp 0
transform 1 0 870 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1104_
timestamp 0
transform 1 0 450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1105_
timestamp 0
transform 1 0 310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1106_
timestamp 0
transform 1 0 1150 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1107_
timestamp 0
transform 1 0 730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1108_
timestamp 0
transform 1 0 1170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1109_
timestamp 0
transform -1 0 1450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1110_
timestamp 0
transform -1 0 750 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1111_
timestamp 0
transform -1 0 190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1112_
timestamp 0
transform -1 0 470 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1113_
timestamp 0
transform -1 0 1210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1114_
timestamp 0
transform 1 0 1450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1115_
timestamp 0
transform 1 0 710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1116_
timestamp 0
transform 1 0 1210 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1117_
timestamp 0
transform -1 0 610 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1118_
timestamp 0
transform -1 0 310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1119_
timestamp 0
transform 1 0 1070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1120_
timestamp 0
transform -1 0 970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1121_
timestamp 0
transform 1 0 830 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1122_
timestamp 0
transform -1 0 330 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1123_
timestamp 0
transform -1 0 710 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1124_
timestamp 0
transform -1 0 590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1125_
timestamp 0
transform -1 0 470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1126_
timestamp 0
transform 1 0 2310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1127_
timestamp 0
transform -1 0 1770 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1128_
timestamp 0
transform 1 0 1850 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1129_
timestamp 0
transform 1 0 2150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1130_
timestamp 0
transform 1 0 1990 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1131_
timestamp 0
transform -1 0 2110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1132_
timestamp 0
transform 1 0 2210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1133_
timestamp 0
transform -1 0 1630 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1134_
timestamp 0
transform 1 0 2870 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1135_
timestamp 0
transform 1 0 1870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1136_
timestamp 0
transform -1 0 2030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1137_
timestamp 0
transform -1 0 1750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1138_
timestamp 0
transform -1 0 50 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1139_
timestamp 0
transform -1 0 190 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1140_
timestamp 0
transform -1 0 630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1141_
timestamp 0
transform -1 0 330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1142_
timestamp 0
transform -1 0 190 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1143_
timestamp 0
transform 1 0 170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1144_
timestamp 0
transform -1 0 50 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1145_
timestamp 0
transform 1 0 170 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1146_
timestamp 0
transform -1 0 50 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1147_
timestamp 0
transform -1 0 50 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1148_
timestamp 0
transform 1 0 310 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1149_
timestamp 0
transform 1 0 170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1150_
timestamp 0
transform -1 0 2370 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1151_
timestamp 0
transform -1 0 1390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1152_
timestamp 0
transform -1 0 1710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1153_
timestamp 0
transform -1 0 1370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1154_
timestamp 0
transform -1 0 1430 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1155_
timestamp 0
transform 1 0 1550 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1156_
timestamp 0
transform 1 0 1290 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1157_
timestamp 0
transform -1 0 1110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1158_
timestamp 0
transform -1 0 1250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1159_
timestamp 0
transform -1 0 1690 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1160_
timestamp 0
transform -1 0 1170 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1161_
timestamp 0
transform -1 0 990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1162_
timestamp 0
transform 1 0 730 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1163_
timestamp 0
transform -1 0 50 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1164_
timestamp 0
transform -1 0 50 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1165_
timestamp 0
transform -1 0 1030 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1166_
timestamp 0
transform -1 0 1250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1167_
timestamp 0
transform 1 0 850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1168_
timestamp 0
transform 1 0 450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1169_
timestamp 0
transform 1 0 1010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1170_
timestamp 0
transform -1 0 470 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1171_
timestamp 0
transform 1 0 310 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1172_
timestamp 0
transform 1 0 590 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1173_
timestamp 0
transform 1 0 1010 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1174_
timestamp 0
transform 1 0 1430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1175_
timestamp 0
transform 1 0 870 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1176_
timestamp 0
transform 1 0 1150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1177_
timestamp 0
transform 1 0 1850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1178_
timestamp 0
transform 1 0 1990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1179_
timestamp 0
transform -1 0 2570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1180_
timestamp 0
transform -1 0 50 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1181_
timestamp 0
transform -1 0 1750 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1182_
timestamp 0
transform -1 0 2430 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1183_
timestamp 0
transform 1 0 1850 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1184_
timestamp 0
transform 1 0 1950 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1185_
timestamp 0
transform -1 0 2010 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1186_
timestamp 0
transform -1 0 1690 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1187_
timestamp 0
transform 1 0 1910 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1188_
timestamp 0
transform 1 0 2190 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1189_
timestamp 0
transform -1 0 1610 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1190_
timestamp 0
transform -1 0 2070 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1191_
timestamp 0
transform -1 0 1470 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1192_
timestamp 0
transform -1 0 990 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1193_
timestamp 0
transform -1 0 850 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1194_
timestamp 0
transform -1 0 470 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1195_
timestamp 0
transform 1 0 130 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1196_
timestamp 0
transform -1 0 610 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1197_
timestamp 0
transform 1 0 870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1198_
timestamp 0
transform -1 0 1030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1199_
timestamp 0
transform 1 0 1570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1200_
timestamp 0
transform 1 0 1290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1201_
timestamp 0
transform 1 0 1710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1202_
timestamp 0
transform -1 0 1330 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1203_
timestamp 0
transform 1 0 2130 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1204_
timestamp 0
transform 1 0 3210 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1205_
timestamp 0
transform -1 0 2470 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1206_
timestamp 0
transform -1 0 3070 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1207_
timestamp 0
transform 1 0 2690 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1208_
timestamp 0
transform 1 0 2710 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1209_
timestamp 0
transform -1 0 2870 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1210_
timestamp 0
transform 1 0 2990 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1211_
timestamp 0
transform -1 0 1830 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1212_
timestamp 0
transform -1 0 1190 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1213_
timestamp 0
transform -1 0 1090 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1214_
timestamp 0
transform 1 0 970 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1215_
timestamp 0
transform -1 0 610 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1216_
timestamp 0
transform 1 0 410 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1217_
timestamp 0
transform 1 0 830 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1218_
timestamp 0
transform 1 0 1310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1219_
timestamp 0
transform 1 0 1630 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1220_
timestamp 0
transform -1 0 2270 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1221_
timestamp 0
transform 1 0 2350 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1222_
timestamp 0
transform 1 0 2890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1223_
timestamp 0
transform -1 0 2590 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1224_
timestamp 0
transform 1 0 2770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1225_
timestamp 0
transform -1 0 2810 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1226_
timestamp 0
transform -1 0 3070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1227_
timestamp 0
transform 1 0 2950 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1228_
timestamp 0
transform -1 0 3010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1229_
timestamp 0
transform 1 0 3050 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1230_
timestamp 0
transform 1 0 3250 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1231_
timestamp 0
transform 1 0 1950 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1232_
timestamp 0
transform 1 0 2050 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1233_
timestamp 0
transform -1 0 2510 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1234_
timestamp 0
transform 1 0 1210 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1235_
timestamp 0
transform 1 0 1350 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1236_
timestamp 0
transform -1 0 290 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1237_
timestamp 0
transform 1 0 550 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1238_
timestamp 0
transform 1 0 690 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1239_
timestamp 0
transform 1 0 1990 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1240_
timestamp 0
transform -1 0 2110 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1241_
timestamp 0
transform 1 0 1710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1242_
timestamp 0
transform 1 0 2190 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1243_
timestamp 0
transform -1 0 2670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1244_
timestamp 0
transform -1 0 1310 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1245_
timestamp 0
transform -1 0 870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1246_
timestamp 0
transform -1 0 470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1247_
timestamp 0
transform 1 0 2390 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1248_
timestamp 0
transform -1 0 1390 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1249_
timestamp 0
transform -1 0 2290 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1250_
timestamp 0
transform -1 0 2090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1251_
timestamp 0
transform 1 0 2010 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1252_
timestamp 0
transform -1 0 1770 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1253_
timestamp 0
transform -1 0 1250 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1254_
timestamp 0
transform 1 0 2130 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1255_
timestamp 0
transform 1 0 1890 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1256_
timestamp 0
transform -1 0 1630 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1257_
timestamp 0
transform -1 0 970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1258_
timestamp 0
transform 1 0 170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1259_
timestamp 0
transform 1 0 2010 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1260_
timestamp 0
transform -1 0 1870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1261_
timestamp 0
transform -1 0 1890 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1262_
timestamp 0
transform -1 0 2430 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1263_
timestamp 0
transform -1 0 2150 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1264_
timestamp 0
transform -1 0 1630 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1265_
timestamp 0
transform -1 0 1290 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1266_
timestamp 0
transform 1 0 1750 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1267_
timestamp 0
transform 1 0 2550 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1268_
timestamp 0
transform -1 0 1390 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1269_
timestamp 0
transform -1 0 1150 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1270_
timestamp 0
transform 1 0 870 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1271_
timestamp 0
transform -1 0 450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1272_
timestamp 0
transform 1 0 1730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1273_
timestamp 0
transform 1 0 1470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1274_
timestamp 0
transform 1 0 1670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1275_
timestamp 0
transform -1 0 1370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1276_
timestamp 0
transform -1 0 330 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1277_
timestamp 0
transform -1 0 830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1278_
timestamp 0
transform 1 0 1630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1279_
timestamp 0
transform 1 0 1490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1280_
timestamp 0
transform 1 0 590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1281_
timestamp 0
transform -1 0 190 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1282_
timestamp 0
transform 1 0 990 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1283_
timestamp 0
transform 1 0 830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1284_
timestamp 0
transform -1 0 450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1285_
timestamp 0
transform -1 0 450 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1286_
timestamp 0
transform -1 0 50 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1287_
timestamp 0
transform -1 0 50 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1288_
timestamp 0
transform -1 0 730 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1289_
timestamp 0
transform -1 0 50 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1290_
timestamp 0
transform -1 0 170 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1291_
timestamp 0
transform 1 0 170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1292_
timestamp 0
transform -1 0 1110 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1293_
timestamp 0
transform 1 0 310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1294_
timestamp 0
transform -1 0 310 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1295_
timestamp 0
transform -1 0 810 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1296_
timestamp 0
transform 1 0 310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1297_
timestamp 0
transform -1 0 330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1298_
timestamp 0
transform -1 0 950 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1299_
timestamp 0
transform -1 0 50 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1300_
timestamp 0
transform -1 0 50 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1301_
timestamp 0
transform 1 0 830 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1302_
timestamp 0
transform -1 0 750 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1303_
timestamp 0
transform 1 0 310 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1304_
timestamp 0
transform 1 0 170 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1305_
timestamp 0
transform 1 0 590 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1306_
timestamp 0
transform 1 0 970 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1307_
timestamp 0
transform 1 0 1150 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1308_
timestamp 0
transform -1 0 470 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1309_
timestamp 0
transform 1 0 730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1310_
timestamp 0
transform 1 0 1110 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1311_
timestamp 0
transform 1 0 2290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1312_
timestamp 0
transform 1 0 2390 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1313_
timestamp 0
transform 1 0 2130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1314_
timestamp 0
transform 1 0 1850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1315_
timestamp 0
transform 1 0 1450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1316_
timestamp 0
transform 1 0 1570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1317_
timestamp 0
transform 1 0 1950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1318_
timestamp 0
transform 1 0 2090 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1319_
timestamp 0
transform 1 0 2370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1320_
timestamp 0
transform -1 0 2290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1321_
timestamp 0
transform -1 0 2130 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1322_
timestamp 0
transform -1 0 2450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1323_
timestamp 0
transform 1 0 2490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1324_
timestamp 0
transform 1 0 3450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1325_
timestamp 0
transform -1 0 3330 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1326_
timestamp 0
transform 1 0 3250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1327_
timestamp 0
transform 1 0 3390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1328_
timestamp 0
transform -1 0 3690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1329_
timestamp 0
transform -1 0 3550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1330_
timestamp 0
transform 1 0 3530 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1331_
timestamp 0
transform 1 0 3390 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1332_
timestamp 0
transform 1 0 2750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1333_
timestamp 0
transform -1 0 2830 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1334_
timestamp 0
transform 1 0 3450 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1335_
timestamp 0
transform 1 0 2910 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1336_
timestamp 0
transform 1 0 450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1337_
timestamp 0
transform 1 0 590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1338_
timestamp 0
transform -1 0 1490 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1339_
timestamp 0
transform 1 0 170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1340_
timestamp 0
transform 1 0 450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1341_
timestamp 0
transform -1 0 1350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1342_
timestamp 0
transform 1 0 830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1343_
timestamp 0
transform -1 0 1470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1344_
timestamp 0
transform -1 0 1490 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1345_
timestamp 0
transform 1 0 1070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1346_
timestamp 0
transform 1 0 1190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1347_
timestamp 0
transform 1 0 930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1348_
timestamp 0
transform -1 0 990 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1349_
timestamp 0
transform 1 0 1110 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1350_
timestamp 0
transform -1 0 710 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1351_
timestamp 0
transform 1 0 710 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1352_
timestamp 0
transform -1 0 330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1353_
timestamp 0
transform -1 0 190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1354_
timestamp 0
transform 1 0 2070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1355_
timestamp 0
transform 1 0 2110 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1356_
timestamp 0
transform -1 0 2470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1357_
timestamp 0
transform -1 0 3110 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1358_
timestamp 0
transform -1 0 2350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1359_
timestamp 0
transform 1 0 2710 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1360_
timestamp 0
transform 1 0 2210 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1361_
timestamp 0
transform -1 0 1990 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1362_
timestamp 0
transform 1 0 3250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1363_
timestamp 0
transform -1 0 2210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1364_
timestamp 0
transform 1 0 2270 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1365_
timestamp 0
transform -1 0 1810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1366_
timestamp 0
transform 1 0 1670 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1367_
timestamp 0
transform -1 0 1950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1368_
timestamp 0
transform -1 0 1850 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1369_
timestamp 0
transform -1 0 1430 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1370_
timestamp 0
transform -1 0 1550 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1371_
timestamp 0
transform -1 0 50 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1372_
timestamp 0
transform -1 0 50 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1373_
timestamp 0
transform 1 0 710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1374_
timestamp 0
transform -1 0 590 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1375_
timestamp 0
transform -1 0 450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1376_
timestamp 0
transform -1 0 170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1377_
timestamp 0
transform -1 0 570 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1378_
timestamp 0
transform -1 0 590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1379_
timestamp 0
transform -1 0 170 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1380_
timestamp 0
transform 1 0 410 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1381_
timestamp 0
transform 1 0 730 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1382_
timestamp 0
transform 1 0 430 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1383_
timestamp 0
transform -1 0 670 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1384_
timestamp 0
transform -1 0 290 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1385_
timestamp 0
transform -1 0 50 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1386_
timestamp 0
transform -1 0 50 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1387_
timestamp 0
transform 1 0 170 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1388_
timestamp 0
transform 1 0 450 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1389_
timestamp 0
transform 1 0 1070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1390_
timestamp 0
transform 1 0 830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1391_
timestamp 0
transform 1 0 590 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1392_
timestamp 0
transform 1 0 310 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1393_
timestamp 0
transform 1 0 690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1394_
timestamp 0
transform 1 0 1210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1395_
timestamp 0
transform 1 0 930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1396_
timestamp 0
transform -1 0 570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1397_
timestamp 0
transform 1 0 1110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1398_
timestamp 0
transform 1 0 1950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1399_
timestamp 0
transform 1 0 2510 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1400_
timestamp 0
transform -1 0 2570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1401_
timestamp 0
transform -1 0 1030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1402_
timestamp 0
transform 1 0 870 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1403_
timestamp 0
transform 1 0 1270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1404_
timestamp 0
transform -1 0 1090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1405_
timestamp 0
transform -1 0 1850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1406_
timestamp 0
transform 1 0 2690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1407_
timestamp 0
transform 1 0 2770 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1408_
timestamp 0
transform 1 0 3170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1409_
timestamp 0
transform 1 0 3590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1410_
timestamp 0
transform 1 0 3310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1411_
timestamp 0
transform 1 0 3450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1412_
timestamp 0
transform -1 0 2930 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1413_
timestamp 0
transform 1 0 2850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1414_
timestamp 0
transform 1 0 3930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1415_
timestamp 0
transform 1 0 2350 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1416_
timestamp 0
transform 1 0 2430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1417_
timestamp 0
transform 1 0 2570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1418_
timestamp 0
transform 1 0 830 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1419_
timestamp 0
transform -1 0 610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1420_
timestamp 0
transform -1 0 50 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1421_
timestamp 0
transform -1 0 1590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1422_
timestamp 0
transform 1 0 1690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1423_
timestamp 0
transform 1 0 2190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1424_
timestamp 0
transform 1 0 2310 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1425_
timestamp 0
transform 1 0 2070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1426_
timestamp 0
transform -1 0 1950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1427_
timestamp 0
transform -1 0 1810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1428_
timestamp 0
transform 1 0 2430 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1429_
timestamp 0
transform 1 0 2310 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1430_
timestamp 0
transform -1 0 2190 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1431_
timestamp 0
transform 1 0 1390 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1432_
timestamp 0
transform 1 0 1350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1433_
timestamp 0
transform 1 0 2550 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1434_
timestamp 0
transform 1 0 2710 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1435_
timestamp 0
transform 1 0 2750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1436_
timestamp 0
transform 1 0 3330 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1437_
timestamp 0
transform 1 0 2650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1438_
timestamp 0
transform -1 0 2570 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1439_
timestamp 0
transform -1 0 2610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1440_
timestamp 0
transform 1 0 2450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1441_
timestamp 0
transform -1 0 2590 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1442_
timestamp 0
transform -1 0 2330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1443_
timestamp 0
transform 1 0 1910 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1444_
timestamp 0
transform -1 0 1250 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1445_
timestamp 0
transform -1 0 1390 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1446_
timestamp 0
transform -1 0 750 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1447_
timestamp 0
transform -1 0 610 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1448_
timestamp 0
transform -1 0 1650 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1449_
timestamp 0
transform 1 0 1510 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1450_
timestamp 0
transform -1 0 1790 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1451_
timestamp 0
transform -1 0 850 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1452_
timestamp 0
transform -1 0 50 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1453_
timestamp 0
transform 1 0 290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1454_
timestamp 0
transform -1 0 1250 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1455_
timestamp 0
transform -1 0 990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1456_
timestamp 0
transform 1 0 1110 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1457_
timestamp 0
transform -1 0 850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1458_
timestamp 0
transform -1 0 330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1459_
timestamp 0
transform -1 0 190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1460_
timestamp 0
transform 1 0 170 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1461_
timestamp 0
transform -1 0 470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1462_
timestamp 0
transform 1 0 690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1463_
timestamp 0
transform -1 0 1170 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1464_
timestamp 0
transform 1 0 1210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1465_
timestamp 0
transform 1 0 870 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1466_
timestamp 0
transform 1 0 1010 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1467_
timestamp 0
transform 1 0 1270 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1468_
timestamp 0
transform -1 0 1590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1469_
timestamp 0
transform 1 0 2490 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1470_
timestamp 0
transform -1 0 2250 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1471_
timestamp 0
transform -1 0 2650 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1472_
timestamp 0
transform -1 0 2910 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1473_
timestamp 0
transform -1 0 2790 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1474_
timestamp 0
transform 1 0 2830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1475_
timestamp 0
transform 1 0 3330 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1476_
timestamp 0
transform -1 0 2930 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1477_
timestamp 0
transform 1 0 3130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1478_
timestamp 0
transform 1 0 3270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1479_
timestamp 0
transform 1 0 3610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1480_
timestamp 0
transform -1 0 3210 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1481_
timestamp 0
transform -1 0 3050 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1482_
timestamp 0
transform 1 0 4090 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1483_
timestamp 0
transform -1 0 2590 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1484_
timestamp 0
transform -1 0 3390 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1485_
timestamp 0
transform 1 0 3350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1486_
timestamp 0
transform 1 0 2930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1487_
timestamp 0
transform -1 0 2050 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1488_
timestamp 0
transform -1 0 1270 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1489_
timestamp 0
transform 1 0 1110 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1490_
timestamp 0
transform 1 0 2770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1491_
timestamp 0
transform -1 0 3110 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1492_
timestamp 0
transform 1 0 2870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1493_
timestamp 0
transform -1 0 2690 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1494_
timestamp 0
transform -1 0 2850 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1495_
timestamp 0
transform 1 0 2950 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1496_
timestamp 0
transform 1 0 3190 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1497_
timestamp 0
transform -1 0 3470 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1498_
timestamp 0
transform 1 0 3030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1499_
timestamp 0
transform -1 0 3170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1500_
timestamp 0
transform -1 0 3790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1501_
timestamp 0
transform 1 0 4130 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1502_
timestamp 0
transform 1 0 4010 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1503_
timestamp 0
transform 1 0 4410 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1504_
timestamp 0
transform -1 0 3910 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1505_
timestamp 0
transform -1 0 3630 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1506_
timestamp 0
transform -1 0 3770 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1507_
timestamp 0
transform 1 0 3330 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1508_
timestamp 0
transform -1 0 1790 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1509_
timestamp 0
transform -1 0 3210 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1510_
timestamp 0
transform -1 0 1510 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1511_
timestamp 0
transform 1 0 970 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1512_
timestamp 0
transform 1 0 2010 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1513_
timestamp 0
transform -1 0 1650 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1514_
timestamp 0
transform 1 0 1350 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1515_
timestamp 0
transform 1 0 1650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1516_
timestamp 0
transform -1 0 1890 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1517_
timestamp 0
transform -1 0 1930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1518_
timestamp 0
transform -1 0 1810 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1519_
timestamp 0
transform 1 0 1510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1520_
timestamp 0
transform 1 0 310 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1521_
timestamp 0
transform 1 0 450 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1522_
timestamp 0
transform 1 0 2050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1523_
timestamp 0
transform -1 0 2630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1524_
timestamp 0
transform 1 0 3130 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1525_
timestamp 0
transform 1 0 2990 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1526_
timestamp 0
transform -1 0 2990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1527_
timestamp 0
transform 1 0 3070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1528_
timestamp 0
transform 1 0 3210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1529_
timestamp 0
transform 1 0 2630 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1530_
timestamp 0
transform -1 0 3150 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1531_
timestamp 0
transform 1 0 2190 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1532_
timestamp 0
transform -1 0 2470 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1533_
timestamp 0
transform -1 0 2330 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1534_
timestamp 0
transform 1 0 2750 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1535_
timestamp 0
transform 1 0 2890 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1536_
timestamp 0
transform 1 0 3290 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1537_
timestamp 0
transform 1 0 2190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1538_
timestamp 0
transform -1 0 2330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1539_
timestamp 0
transform -1 0 2910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1540_
timestamp 0
transform -1 0 2530 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1541_
timestamp 0
transform 1 0 3550 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1542_
timestamp 0
transform 1 0 3990 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1543_
timestamp 0
transform 1 0 3890 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1544_
timestamp 0
transform 1 0 3910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1545_
timestamp 0
transform -1 0 4290 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1546_
timestamp 0
transform -1 0 3730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1547_
timestamp 0
transform 1 0 3790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1548_
timestamp 0
transform 1 0 4110 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1549_
timestamp 0
transform -1 0 3410 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1550_
timestamp 0
transform -1 0 3490 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1551_
timestamp 0
transform -1 0 3310 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1552_
timestamp 0
transform -1 0 3170 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1553_
timestamp 0
transform 1 0 2890 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1554_
timestamp 0
transform -1 0 2270 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1555_
timestamp 0
transform -1 0 2770 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1556_
timestamp 0
transform -1 0 2390 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1557_
timestamp 0
transform -1 0 2130 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1558_
timestamp 0
transform 1 0 2550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1559_
timestamp 0
transform -1 0 2670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1560_
timestamp 0
transform 1 0 2810 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1561_
timestamp 0
transform 1 0 2930 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1562_
timestamp 0
transform 1 0 2410 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1563_
timestamp 0
transform -1 0 2990 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1564_
timestamp 0
transform 1 0 2670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1565_
timestamp 0
transform 1 0 3150 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1566_
timestamp 0
transform 1 0 3030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1567_
timestamp 0
transform -1 0 2630 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1568_
timestamp 0
transform 1 0 2990 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1569_
timestamp 0
transform 1 0 3170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1570_
timestamp 0
transform 1 0 3310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1571_
timestamp 0
transform -1 0 2890 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1572_
timestamp 0
transform 1 0 3270 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1573_
timestamp 0
transform -1 0 2750 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1574_
timestamp 0
transform 1 0 2790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1575_
timestamp 0
transform 1 0 3410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1576_
timestamp 0
transform 1 0 3690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1577_
timestamp 0
transform 1 0 4030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1578_
timestamp 0
transform -1 0 3750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1579_
timestamp 0
transform 1 0 1710 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1580_
timestamp 0
transform 1 0 1570 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1581_
timestamp 0
transform 1 0 1730 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1582_
timestamp 0
transform -1 0 3770 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1583_
timestamp 0
transform 1 0 3610 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1584_
timestamp 0
transform -1 0 3490 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1585_
timestamp 0
transform 1 0 3390 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1586_
timestamp 0
transform -1 0 3590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1587_
timestamp 0
transform -1 0 3850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1588_
timestamp 0
transform 1 0 3650 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1589_
timestamp 0
transform -1 0 3790 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1590_
timestamp 0
transform -1 0 3410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1591_
timestamp 0
transform 1 0 3550 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1592_
timestamp 0
transform 1 0 3010 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1593_
timestamp 0
transform -1 0 3590 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1594_
timestamp 0
transform -1 0 3470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1595_
timestamp 0
transform 1 0 3190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1596_
timestamp 0
transform -1 0 3070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1597_
timestamp 0
transform -1 0 2950 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1598_
timestamp 0
transform 1 0 3050 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__1599_
timestamp 0
transform 1 0 2610 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1600_
timestamp 0
transform -1 0 2810 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1601_
timestamp 0
transform 1 0 3130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1602_
timestamp 0
transform -1 0 3430 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1603_
timestamp 0
transform 1 0 3530 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1604_
timestamp 0
transform 1 0 3550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1605_
timestamp 0
transform 1 0 3670 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1606_
timestamp 0
transform -1 0 3370 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1607_
timestamp 0
transform -1 0 2750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1608_
timestamp 0
transform 1 0 3950 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1609_
timestamp 0
transform 1 0 3810 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1610_
timestamp 0
transform 1 0 1850 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1611_
timestamp 0
transform 1 0 2510 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1612_
timestamp 0
transform -1 0 3610 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1613_
timestamp 0
transform -1 0 3470 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1614_
timestamp 0
transform 1 0 3310 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1615_
timestamp 0
transform -1 0 3430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1616_
timestamp 0
transform -1 0 3250 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1617_
timestamp 0
transform -1 0 3250 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1618_
timestamp 0
transform -1 0 3310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1619_
timestamp 0
transform -1 0 3330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__1620_
timestamp 0
transform -1 0 3310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1621_
timestamp 0
transform 1 0 3350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1622_
timestamp 0
transform 1 0 3490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1623_
timestamp 0
transform 1 0 3730 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1624_
timestamp 0
transform -1 0 3630 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1625_
timestamp 0
transform -1 0 3410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1626_
timestamp 0
transform -1 0 2890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1627_
timestamp 0
transform -1 0 3030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1628_
timestamp 0
transform -1 0 3530 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1629_
timestamp 0
transform 1 0 3370 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1630_
timestamp 0
transform -1 0 3170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1631_
timestamp 0
transform 1 0 2510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1632_
timestamp 0
transform 1 0 2230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1633_
timestamp 0
transform 1 0 2650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1634_
timestamp 0
transform -1 0 3370 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1635_
timestamp 0
transform 1 0 2650 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1636_
timestamp 0
transform 1 0 2910 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1637_
timestamp 0
transform -1 0 3090 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1638_
timestamp 0
transform -1 0 3830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1639_
timestamp 0
transform 1 0 3530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1640_
timestamp 0
transform 1 0 3630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1641_
timestamp 0
transform 1 0 3670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1642_
timestamp 0
transform 1 0 2410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1643_
timestamp 0
transform 1 0 2790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1644_
timestamp 0
transform 1 0 2930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1645_
timestamp 0
transform 1 0 3210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1646_
timestamp 0
transform 1 0 3070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1647_
timestamp 0
transform 1 0 3330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1648_
timestamp 0
transform -1 0 3730 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1649_
timestamp 0
transform 1 0 4710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1650_
timestamp 0
transform 1 0 4570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1651_
timestamp 0
transform 1 0 5090 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1652_
timestamp 0
transform 1 0 4950 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1653_
timestamp 0
transform 1 0 4570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1654_
timestamp 0
transform -1 0 4710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1655_
timestamp 0
transform 1 0 4970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1656_
timestamp 0
transform 1 0 4830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1657_
timestamp 0
transform 1 0 5590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1658_
timestamp 0
transform 1 0 5450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__1659_
timestamp 0
transform 1 0 4950 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1660_
timestamp 0
transform -1 0 5090 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__1661_
timestamp 0
transform 1 0 5230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1662_
timestamp 0
transform 1 0 5090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1663_
timestamp 0
transform 1 0 5010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1664_
timestamp 0
transform -1 0 4890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__1692_
timestamp 0
transform 1 0 5350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1693_
timestamp 0
transform 1 0 5450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__1694_
timestamp 0
transform 1 0 5450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1695_
timestamp 0
transform -1 0 5590 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1696_
timestamp 0
transform 1 0 5630 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1697_
timestamp 0
transform -1 0 5250 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1698_
timestamp 0
transform -1 0 5350 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1699_
timestamp 0
transform -1 0 5150 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1700_
timestamp 0
transform -1 0 4450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1701_
timestamp 0
transform -1 0 4550 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1702_
timestamp 0
transform 1 0 4550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1703_
timestamp 0
transform 1 0 5530 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__1704_
timestamp 0
transform 1 0 4770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1705_
timestamp 0
transform 1 0 4390 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1706_
timestamp 0
transform -1 0 4730 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1707_
timestamp 0
transform 1 0 4850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1708_
timestamp 0
transform -1 0 4670 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1709_
timestamp 0
transform 1 0 4710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1710_
timestamp 0
transform 1 0 5210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1711_
timestamp 0
transform 1 0 5070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1712_
timestamp 0
transform -1 0 5310 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1713_
timestamp 0
transform -1 0 5270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1714_
timestamp 0
transform 1 0 5290 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1715_
timestamp 0
transform 1 0 5530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1716_
timestamp 0
transform -1 0 5450 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1717_
timestamp 0
transform 1 0 5450 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1718_
timestamp 0
transform -1 0 4890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1719_
timestamp 0
transform -1 0 5190 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1720_
timestamp 0
transform -1 0 5410 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1721_
timestamp 0
transform -1 0 4470 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1722_
timestamp 0
transform -1 0 4410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1723_
timestamp 0
transform 1 0 4230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1724_
timestamp 0
transform 1 0 4070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1725_
timestamp 0
transform -1 0 4190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1726_
timestamp 0
transform 1 0 4290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1727_
timestamp 0
transform 1 0 4310 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1728_
timestamp 0
transform 1 0 3470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1729_
timestamp 0
transform -1 0 3450 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1730_
timestamp 0
transform -1 0 3590 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1731_
timestamp 0
transform 1 0 3670 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1732_
timestamp 0
transform -1 0 3830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1733_
timestamp 0
transform 1 0 3970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1734_
timestamp 0
transform -1 0 5090 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1735_
timestamp 0
transform -1 0 4950 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1736_
timestamp 0
transform 1 0 4850 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1737_
timestamp 0
transform 1 0 4570 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1738_
timestamp 0
transform 1 0 5010 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1739_
timestamp 0
transform 1 0 5110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1740_
timestamp 0
transform 1 0 4970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1741_
timestamp 0
transform 1 0 4770 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__1742_
timestamp 0
transform -1 0 4090 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1743_
timestamp 0
transform 1 0 3930 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1744_
timestamp 0
transform -1 0 3830 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1745_
timestamp 0
transform 1 0 3870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1746_
timestamp 0
transform -1 0 3730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1747_
timestamp 0
transform 1 0 4210 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1748_
timestamp 0
transform -1 0 4150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1749_
timestamp 0
transform -1 0 4670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1750_
timestamp 0
transform 1 0 3850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1751_
timestamp 0
transform -1 0 3970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__1752_
timestamp 0
transform -1 0 3910 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1753_
timestamp 0
transform -1 0 4170 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1754_
timestamp 0
transform 1 0 4010 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1755_
timestamp 0
transform 1 0 4090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1756_
timestamp 0
transform -1 0 3590 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1757_
timestamp 0
transform 1 0 3870 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1758_
timestamp 0
transform 1 0 4290 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1759_
timestamp 0
transform -1 0 4670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1760_
timestamp 0
transform 1 0 4490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1761_
timestamp 0
transform -1 0 4390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1762_
timestamp 0
transform -1 0 4170 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1763_
timestamp 0
transform -1 0 4030 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1764_
timestamp 0
transform -1 0 4010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1765_
timestamp 0
transform 1 0 4250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1766_
timestamp 0
transform 1 0 4150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1767_
timestamp 0
transform 1 0 4430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1768_
timestamp 0
transform -1 0 4090 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1769_
timestamp 0
transform 1 0 4690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1770_
timestamp 0
transform -1 0 4430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1771_
timestamp 0
transform -1 0 4350 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1772_
timestamp 0
transform -1 0 4470 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1773_
timestamp 0
transform -1 0 4290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1774_
timestamp 0
transform 1 0 4550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1775_
timestamp 0
transform -1 0 4510 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1776_
timestamp 0
transform 1 0 4630 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1777_
timestamp 0
transform 1 0 4930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1778_
timestamp 0
transform 1 0 4790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1779_
timestamp 0
transform 1 0 4770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1780_
timestamp 0
transform 1 0 4530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1781_
timestamp 0
transform -1 0 4230 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1782_
timestamp 0
transform 1 0 4310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1783_
timestamp 0
transform -1 0 2810 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1784_
timestamp 0
transform -1 0 3590 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1785_
timestamp 0
transform -1 0 3690 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1786_
timestamp 0
transform -1 0 4190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1787_
timestamp 0
transform 1 0 4350 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1788_
timestamp 0
transform 1 0 5010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1789_
timestamp 0
transform 1 0 4870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1790_
timestamp 0
transform 1 0 5110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1791_
timestamp 0
transform 1 0 5570 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1792_
timestamp 0
transform 1 0 5530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1793_
timestamp 0
transform 1 0 5370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1794_
timestamp 0
transform 1 0 5370 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1795_
timestamp 0
transform -1 0 5250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1796_
timestamp 0
transform 1 0 5490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1797_
timestamp 0
transform -1 0 5370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1798_
timestamp 0
transform 1 0 4590 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1799_
timestamp 0
transform 1 0 4730 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1800_
timestamp 0
transform 1 0 4190 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1801_
timestamp 0
transform -1 0 3970 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1802_
timestamp 0
transform -1 0 3830 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1803_
timestamp 0
transform 1 0 3690 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1804_
timestamp 0
transform 1 0 3810 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1805_
timestamp 0
transform -1 0 4350 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1806_
timestamp 0
transform 1 0 4370 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1807_
timestamp 0
transform 1 0 4250 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1808_
timestamp 0
transform -1 0 4690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1809_
timestamp 0
transform -1 0 4830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1810_
timestamp 0
transform -1 0 4910 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1811_
timestamp 0
transform -1 0 4790 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1812_
timestamp 0
transform 1 0 4610 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1813_
timestamp 0
transform 1 0 5070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1814_
timestamp 0
transform -1 0 4950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1815_
timestamp 0
transform 1 0 4890 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1816_
timestamp 0
transform 1 0 5030 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1817_
timestamp 0
transform 1 0 5250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1818_
timestamp 0
transform 1 0 5110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1819_
timestamp 0
transform -1 0 4450 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1820_
timestamp 0
transform 1 0 4490 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1821_
timestamp 0
transform -1 0 4910 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1822_
timestamp 0
transform 1 0 4770 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1823_
timestamp 0
transform -1 0 4090 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1824_
timestamp 0
transform 1 0 4990 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1825_
timestamp 0
transform 1 0 4870 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1826_
timestamp 0
transform -1 0 5370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1827_
timestamp 0
transform -1 0 5210 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1828_
timestamp 0
transform 1 0 5030 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1829_
timestamp 0
transform 1 0 5210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1830_
timestamp 0
transform 1 0 4970 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1831_
timestamp 0
transform 1 0 5070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1832_
timestamp 0
transform 1 0 5210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__1833_
timestamp 0
transform 1 0 5510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1834_
timestamp 0
transform 1 0 5550 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__1835_
timestamp 0
transform -1 0 4570 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1836_
timestamp 0
transform 1 0 4630 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1837_
timestamp 0
transform -1 0 5650 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1838_
timestamp 0
transform -1 0 4690 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1839_
timestamp 0
transform 1 0 4310 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1840_
timestamp 0
transform -1 0 5650 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1841_
timestamp 0
transform 1 0 4810 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1842_
timestamp 0
transform 1 0 5590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__1843_
timestamp 0
transform 1 0 5490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__1844_
timestamp 0
transform 1 0 4870 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1845_
timestamp 0
transform 1 0 5190 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1846_
timestamp 0
transform 1 0 5490 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1847_
timestamp 0
transform -1 0 5370 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__1848_
timestamp 0
transform -1 0 5550 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__1849_
timestamp 0
transform 1 0 5230 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1850_
timestamp 0
transform 1 0 5590 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1851_
timestamp 0
transform -1 0 5470 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1852_
timestamp 0
transform -1 0 5370 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1853_
timestamp 0
transform -1 0 4970 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1854_
timestamp 0
transform 1 0 5410 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1855_
timestamp 0
transform -1 0 5090 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1856_
timestamp 0
transform -1 0 4450 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1857_
timestamp 0
transform -1 0 3930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1858_
timestamp 0
transform -1 0 3970 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1859_
timestamp 0
transform 1 0 4010 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1860_
timestamp 0
transform 1 0 4070 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1861_
timestamp 0
transform -1 0 4190 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1862_
timestamp 0
transform -1 0 4150 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1863_
timestamp 0
transform -1 0 3890 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1864_
timestamp 0
transform -1 0 5230 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1865_
timestamp 0
transform -1 0 5510 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1866_
timestamp 0
transform 1 0 4370 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1867_
timestamp 0
transform -1 0 3950 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1868_
timestamp 0
transform 1 0 4470 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1869_
timestamp 0
transform -1 0 5330 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1870_
timestamp 0
transform -1 0 4870 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1871_
timestamp 0
transform -1 0 5150 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1872_
timestamp 0
transform -1 0 4730 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1873_
timestamp 0
transform -1 0 4970 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1874_
timestamp 0
transform 1 0 5510 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1875_
timestamp 0
transform 1 0 5270 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__1876_
timestamp 0
transform -1 0 5070 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1877_
timestamp 0
transform -1 0 4590 0 1 730
box -6 -8 26 248
use FILL  FILL_1__1878_
timestamp 0
transform -1 0 3870 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1879_
timestamp 0
transform -1 0 3810 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1880_
timestamp 0
transform -1 0 5650 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1881_
timestamp 0
transform 1 0 5510 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1882_
timestamp 0
transform -1 0 5390 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1883_
timestamp 0
transform -1 0 5270 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1884_
timestamp 0
transform -1 0 5150 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__1885_
timestamp 0
transform 1 0 5390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__1886_
timestamp 0
transform -1 0 4750 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1887_
timestamp 0
transform -1 0 4650 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1888_
timestamp 0
transform -1 0 4510 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1889_
timestamp 0
transform 1 0 4250 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1890_
timestamp 0
transform -1 0 3730 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1891_
timestamp 0
transform -1 0 4130 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1892_
timestamp 0
transform -1 0 3610 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1893_
timestamp 0
transform -1 0 3490 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1894_
timestamp 0
transform -1 0 2670 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__1895_
timestamp 0
transform -1 0 2650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__1896_
timestamp 0
transform -1 0 50 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__1897_
timestamp 0
transform 1 0 2670 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1898_
timestamp 0
transform -1 0 3150 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1899_
timestamp 0
transform 1 0 3550 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1900_
timestamp 0
transform -1 0 3270 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__1901_
timestamp 0
transform -1 0 3690 0 1 250
box -6 -8 26 248
use FILL  FILL_1__1902_
timestamp 0
transform -1 0 4010 0 -1 250
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert0
timestamp 0
transform -1 0 2390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert1
timestamp 0
transform -1 0 2510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert2
timestamp 0
transform 1 0 4070 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert3
timestamp 0
transform 1 0 4530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert4
timestamp 0
transform -1 0 3790 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert5
timestamp 0
transform 1 0 1750 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert6
timestamp 0
transform -1 0 1630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert7
timestamp 0
transform 1 0 3730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert8
timestamp 0
transform -1 0 4710 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert9
timestamp 0
transform 1 0 5050 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert10
timestamp 0
transform -1 0 5230 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert11
timestamp 0
transform 1 0 5510 0 -1 250
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert17
timestamp 0
transform -1 0 3910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert18
timestamp 0
transform 1 0 4010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert19
timestamp 0
transform 1 0 5130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert20
timestamp 0
transform 1 0 5330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert21
timestamp 0
transform 1 0 2370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert22
timestamp 0
transform 1 0 5570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert23
timestamp 0
transform -1 0 2270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert24
timestamp 0
transform 1 0 3010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert25
timestamp 0
transform 1 0 2690 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert26
timestamp 0
transform 1 0 1630 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert27
timestamp 0
transform -1 0 3510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert28
timestamp 0
transform -1 0 1510 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert29
timestamp 0
transform -1 0 5430 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert30
timestamp 0
transform 1 0 5170 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert31
timestamp 0
transform 1 0 4770 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert32
timestamp 0
transform 1 0 4970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert12
timestamp 0
transform 1 0 4070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert13
timestamp 0
transform -1 0 4090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert14
timestamp 0
transform 1 0 3510 0 1 5530
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert15
timestamp 0
transform -1 0 3850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert16
timestamp 0
transform 1 0 4390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__1492_
timestamp 0
transform 1 0 2890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert32
timestamp 0
transform 1 0 4990 0 -1 2650
box -6 -8 26 248
<< labels >>
flabel metal1 s 5723 2 5783 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal3 s 5056 5816 5064 5824 3 FreeSans 16 90 0 0 ABCmd_i[7]
port 2 nsew
flabel metal3 s 5096 5816 5104 5824 3 FreeSans 16 90 0 0 ABCmd_i[6]
port 3 nsew
flabel metal3 s 5276 5816 5284 5824 3 FreeSans 16 90 0 0 ABCmd_i[5]
port 4 nsew
flabel metal3 s 5476 5816 5484 5824 3 FreeSans 16 90 0 0 ABCmd_i[4]
port 5 nsew
flabel metal3 s 5516 5816 5524 5824 3 FreeSans 16 90 0 0 ABCmd_i[3]
port 6 nsew
flabel metal2 s 5757 1797 5763 1803 3 FreeSans 16 0 0 0 ABCmd_i[2]
port 7 nsew
flabel metal2 s 5757 2757 5763 2763 3 FreeSans 16 0 0 0 ABCmd_i[1]
port 8 nsew
flabel metal2 s 5757 2797 5763 2803 3 FreeSans 16 0 0 0 ABCmd_i[0]
port 9 nsew
flabel metal3 s 3716 -24 3724 -16 7 FreeSans 16 270 0 0 ACC_o[7]
port 10 nsew
flabel metal3 s 3636 -24 3644 -16 7 FreeSans 16 270 0 0 ACC_o[6]
port 11 nsew
flabel metal3 s 3596 -24 3604 -16 7 FreeSans 16 270 0 0 ACC_o[5]
port 12 nsew
flabel metal3 s 3176 -24 3184 -16 7 FreeSans 16 270 0 0 ACC_o[4]
port 13 nsew
flabel metal3 s 2716 -24 2724 -16 7 FreeSans 16 270 0 0 ACC_o[3]
port 14 nsew
flabel metal2 s -23 3717 -17 3723 7 FreeSans 16 0 0 0 ACC_o[2]
port 15 nsew
flabel metal2 s -23 2797 -17 2803 7 FreeSans 16 0 0 0 ACC_o[1]
port 16 nsew
flabel metal2 s -23 2757 -17 2763 7 FreeSans 16 0 0 0 ACC_o[0]
port 17 nsew
flabel metal3 s 4036 -24 4044 -16 7 FreeSans 16 270 0 0 Done_o
port 18 nsew
flabel metal3 s 4116 5816 4124 5824 3 FreeSans 16 90 0 0 LoadA_i
port 19 nsew
flabel metal3 s 4856 5816 4864 5824 3 FreeSans 16 90 0 0 LoadB_i
port 20 nsew
flabel metal3 s 5016 5816 5024 5824 3 FreeSans 16 90 0 0 LoadCmd_i
port 21 nsew
flabel metal3 s 3616 5816 3624 5824 3 FreeSans 16 90 0 0 clk
port 22 nsew
flabel metal3 s 5556 5816 5564 5824 3 FreeSans 16 90 0 0 reset
port 23 nsew
<< properties >>
string FIXED_BBOX -40 -40 5760 5820
<< end >>
