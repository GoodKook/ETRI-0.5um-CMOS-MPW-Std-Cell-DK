magic
tech scmos
magscale 1 6
timestamp 1721857824
<< nwell >>
rect -36 581 142 815
<< ntransistor >>
rect 50 41 62 101
<< ptransistor >>
rect 50 677 62 737
<< ndiffusion >>
rect 44 41 50 101
rect 62 41 68 101
<< pdiffusion >>
rect 44 677 50 737
rect 62 677 68 737
<< ndcontact >>
rect 8 41 44 101
rect 68 41 104 101
<< pdcontact >>
rect 8 677 44 737
rect 68 677 104 737
<< psubstratepcontact >>
rect -18 -19 123 17
<< nsubstratencontact >>
rect -18 761 123 797
<< polysilicon >>
rect 50 737 62 749
rect 50 665 62 677
rect 50 101 62 113
rect 50 29 62 41
<< metal1 >>
rect -18 797 123 803
rect -18 755 123 761
rect -18 17 123 23
rect -18 -25 123 -19
<< end >>
